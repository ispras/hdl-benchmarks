//
// Conformal-LEC Version 15.10-d003 ( 23-Apr-2015) ( 64 bit executable)
//
module top ( 
    n0 , 
    n1 , 
    n2 , 
    n3 , 
    n4 , 
    n5 , 
    n6 , 
    n7 , 
    n8 , 
    n9 , 
    n10 , 
    n11 , 
    n12 , 
    n13 , 
    n14 , 
    n15 , 
    n16 , 
    n17 , 
    n18 , 
    n19 , 
    n20 , 
    n21 , 
    n22 , 
    n23 , 
    n24 , 
    n25 , 
    n26 , 
    n27 , 
    n28 , 
    n29 , 
    n30 , 
    n31 , 
    n32 , 
    n33 , 
    n34 , 
    n35 , 
    n36 , 
    n37 , 
    n38 , 
    n39 , 
    n40 , 
    n41 , 
    n42 , 
    n43 , 
    n44 , 
    n45 , 
    n46 , 
    n47 , 
    n48 , 
    n49 , 
    n50 , 
    n51 , 
    n52 , 
    n53 , 
    n54 , 
    n55 , 
    n56 , 
    n57 , 
    n58 , 
    n59 , 
    n60 , 
    n61 , 
    n62 , 
    n63 , 
    n64 , 
    n65 , 
    n66 , 
    n67 , 
    n68 , 
    n69 , 
    n70 , 
    n71 , 
    n72 , 
    n73 , 
    n74 , 
    n75 , 
    n76 , 
    n77 , 
    n78 , 
    n79 , 
    n80 , 
    n81 , 
    n82 , 
    n83 , 
    n84 , 
    n85 , 
    n86 , 
    n87 , 
    n88 , 
    n89 , 
    n90 , 
    n91 , 
    n92 , 
    n93 , 
    n94 , 
    n95 , 
    n96 , 
    n97 , 
    n98 , 
    n99 , 
    n100 , 
    n101 , 
    n102 , 
    n103 , 
    n104 , 
    n105 , 
    n106 , 
    n107 , 
    n108 , 
    n109 , 
    n110 , 
    n111 , 
    n112 , 
    n113 , 
    n114 , 
    n115 , 
    n116 , 
    n117 , 
    n118 , 
    n119 , 
    n120 , 
    n121 , 
    n122 , 
    n123 , 
    n124 , 
    n125 , 
    n126 , 
    n127 , 
    n128 , 
    n129 , 
    n130 , 
    n131 , 
    n132 , 
    n133 , 
    n134 , 
    n135 , 
    n136 , 
    n137 , 
    n138 , 
    n139 , 
    n140 , 
    n141 , 
    n142 , 
    n143 , 
    n144 , 
    n145 , 
    n146 , 
    n147 , 
    n148 , 
    n149 , 
    n150 , 
    n151 , 
    n152 , 
    n153 , 
    n154 , 
    n155 , 
    n156 , 
    n157 , 
    n158 , 
    n159 , 
    n160 , 
    n161 , 
    n162 , 
    n163 , 
    n164 , 
    n165 , 
    n166 , 
    n167 , 
    n168 , 
    n169 , 
    n170 , 
    n171 , 
    n172 , 
    n173 , 
    n174 , 
    n175 , 
    n176 , 
    n177 , 
    n178 , 
    n179 , 
    n180 , 
    n181 , 
    n182 , 
    n183 , 
    n184 , 
    n185 , 
    n186 , 
    n187 , 
    n188 , 
    n189 , 
    n190 , 
    n191 , 
    n192 , 
    n193 , 
    n194 , 
    n195 , 
    n196 , 
    n197 , 
    n198 , 
    n199 , 
    n200 , 
    n201 , 
    n202 , 
    n203 , 
    n204 , 
    n205 , 
    n206 , 
    n207 , 
    n208 , 
    n209 , 
    n210 , 
    n211 , 
    n212 , 
    n213 , 
    n214 , 
    n215 , 
    n216 , 
    n217 , 
    n218 , 
    n219 , 
    n220 , 
    n221 , 
    n222 , 
    n223 , 
    n224 , 
    n225 , 
    n226 , 
    n227 , 
    n228 , 
    n229 , 
    n230 , 
    n231 , 
    n232 , 
    n233 , 
    n234 , 
    n235 , 
    n236 , 
    n237 , 
    n238 , 
    n239 , 
    n240 , 
    n241 , 
    n242 , 
    n243 , 
    n244 , 
    n245 , 
    n246 , 
    n247 , 
    n248 , 
    n249 , 
    n250 , 
    n251 , 
    n252 , 
    n253 , 
    n254 , 
    n255 , 
    n256 , 
    n257 , 
    n258 , 
    n259 , 
    n260 , 
    n261 , 
    n262 , 
    n263 , 
    n264 , 
    n265 , 
    n266 , 
    n267 , 
    n268 , 
    n269 , 
    n270 , 
    n271 , 
    n272 , 
    n273 , 
    n274 , 
    n275 , 
    n276 , 
    n277 , 
    n278 , 
    n279 , 
    n280 , 
    n281 , 
    n282 , 
    n283 , 
    n284 , 
    n285 , 
    n286 , 
    n287 , 
    n288 , 
    n289 , 
    n290 , 
    n291 , 
    n292 , 
    n293 , 
    n294 , 
    n295 , 
    n296 , 
    n297 , 
    n298 , 
    n299 , 
    n300 , 
    n301 , 
    n302 , 
    n303 , 
    n304 , 
    n305 , 
    n306 , 
    n307 , 
    n308 , 
    n309 , 
    n310 , 
    n311 , 
    n312 , 
    n313 , 
    n314 , 
    n315 , 
    n316 , 
    n317 , 
    n318 , 
    n319 , 
    n320 , 
    n321 , 
    n322 , 
    n323 , 
    n324 , 
    n325 , 
    n326 , 
    n327 , 
    n328 , 
    n329 , 
    n330 , 
    n331 , 
    n332 , 
    n333 , 
    n334 , 
    n335 , 
    n336 , 
    n337 , 
    n338 , 
    n339 , 
    n340 , 
    n341 , 
    n342 , 
    n343 , 
    n344 , 
    n345 , 
    n346 , 
    n347 , 
    n348 , 
    n349 , 
    n350 , 
    n351 , 
    n352 , 
    n353 , 
    n354 , 
    n355 , 
    n356 , 
    n357 , 
    n358 , 
    n359 , 
    n360 , 
    n361 , 
    n362 , 
    n363 , 
    n364 , 
    n365 , 
    n366 , 
    n367 , 
    n368 , 
    n369 , 
    n370 , 
    n371 , 
    n372 , 
    n373 , 
    n374 , 
    n375 , 
    n376 , 
    n377 , 
    n378 , 
    n379 , 
    n380 , 
    n381 , 
    n382 , 
    n383 , 
    n384 , 
    n385 , 
    n386 , 
    n387 , 
    n388 , 
    n389 , 
    n390 , 
    n391 , 
    n392 , 
    n393 , 
    n394 , 
    n395 , 
    n396 , 
    n397 , 
    n398 , 
    n399 , 
    n400 , 
    n401 , 
    n402 , 
    n403 , 
    n404 , 
    n405 , 
    n406 , 
    n407 , 
    n408 , 
    n409 , 
    n410 , 
    n411 , 
    n412 , 
    n413 , 
    n414 , 
    n415 , 
    n416 , 
    n417 , 
    n418 , 
    n419 , 
    n420 , 
    n421 , 
    n422 , 
    n423 , 
    n424 , 
    n425 , 
    n426 , 
    n427 , 
    n428 , 
    n429 , 
    n430 , 
    n431 , 
    n432 , 
    n433 , 
    n434 , 
    n435 , 
    n436 , 
    n437 , 
    n438 , 
    n439 , 
    n440 , 
    n441 , 
    n442 , 
    n443 , 
    n444 , 
    n445 , 
    n446 , 
    n447 , 
    n448 , 
    n449 , 
    n450 , 
    n451 , 
    n452 , 
    n453 , 
    n454 , 
    n455 , 
    n456 , 
    n457 , 
    n458 , 
    n459 , 
    n460 , 
    n461 , 
    n462 , 
    n463 , 
    n464 , 
    n465 , 
    n466 , 
    n467 , 
    n468 , 
    n469 , 
    n470 , 
    n471 , 
    n472 , 
    n473 , 
    n474 , 
    n475 , 
    n476 , 
    n477 , 
    n478 , 
    n479 , 
    n480 , 
    n481 , 
    n482 , 
    n483 , 
    n484 , 
    n485 , 
    n486 , 
    n487 , 
    n488 , 
    n489 , 
    n490 , 
    n491 , 
    n492 , 
    n493 , 
    n494 , 
    n495 , 
    n496 , 
    n497 , 
    n498 , 
    n499 , 
    n500 , 
    n501 , 
    n502 , 
    n503 , 
    n504 , 
    n505 , 
    n506 , 
    n507 , 
    n508 , 
    n509 , 
    n510 , 
    n511 , 
    n512 , 
    n513 , 
    n514 , 
    n515 , 
    n516 , 
    n517 , 
    n518 , 
    n519 , 
    n520 , 
    n521 , 
    n522 , 
    n523 , 
    n524 , 
    n525 , 
    n526 , 
    n527 , 
    n528 , 
    n529 , 
    n530 , 
    n531 , 
    n532 , 
    n533 , 
    n534 , 
    n535 , 
    n536 , 
    n537 , 
    n538 , 
    n539 , 
    n540 , 
    n541 , 
    n542 , 
    n543 , 
    n544 , 
    n545 , 
    n546 , 
    n547 , 
    n548 , 
    n549 , 
    n550 , 
    n551 , 
    n552 , 
    n553 , 
    n554 , 
    n555 , 
    n556 , 
    n557 , 
    n558 , 
    n559 , 
    n560 , 
    n561 , 
    n562 , 
    n563 , 
    n564 , 
    n565 , 
    n566 , 
    n567 , 
    n568 , 
    n569 , 
    n570 , 
    n571 , 
    n572 , 
    n573 , 
    n574 , 
    n575 , 
    n576 , 
    n577 , 
    n578 , 
    n579 , 
    n580 , 
    n581 , 
    n582 , 
    n583 , 
    n584 , 
    n585 , 
    n586 , 
    n587 , 
    n588 , 
    n589 , 
    n590 , 
    n591 , 
    n592 , 
    n593 , 
    n594 , 
    n595 , 
    n596 , 
    n597 , 
    n598 , 
    n599 , 
    n600 , 
    n601 , 
    n602 , 
    n603 , 
    n604 , 
    n605 , 
    n606 , 
    n607 , 
    n608 , 
    n609 , 
    n610 , 
    n611 , 
    n612 , 
    n613 , 
    n614 , 
    n615 , 
    n616 , 
    n617 , 
    n618 , 
    n619 , 
    n620 , 
    n621 , 
    n622 , 
    n623 , 
    n624 , 
    n625 , 
    n626 , 
    n627 , 
    n628 , 
    n629 , 
    n630 , 
    n631 , 
    n632 , 
    n633 , 
    n634 , 
    n635 , 
    n636 , 
    n637 , 
    n638 , 
    n639 , 
    n640 , 
    n641 , 
    n642 , 
    n643 , 
    n644 , 
    n645 , 
    n646 , 
    n647 , 
    n648 , 
    n649 , 
    n650 , 
    n651 , 
    n652 , 
    n653 , 
    n654 , 
    n655 , 
    n656 , 
    n657 , 
    n658 , 
    n659 , 
    n660 , 
    n661 , 
    n662 , 
    n663 , 
    n664 , 
    n665 , 
    n666 , 
    n667 , 
    n668 , 
    n669 , 
    n670 , 
    n671 , 
    n672 , 
    n673 , 
    n674 , 
    n675 , 
    n676 , 
    n677 , 
    n678 , 
    n679 , 
    n680 , 
    n681 , 
    n682 , 
    n683 , 
    n684 , 
    n685 , 
    n686 , 
    n687 , 
    n688 , 
    n689 , 
    n690 , 
    n691 , 
    n692 , 
    n693 , 
    n694 , 
    n695 , 
    n696 , 
    n697 , 
    n698 , 
    n699 , 
    n700 , 
    n701 , 
    n702 , 
    n703 , 
    n704 , 
    n705 , 
    n706 , 
    n707 , 
    n708 , 
    n709 , 
    n710 , 
    n711 , 
    n712 , 
    n713 , 
    n714 , 
    n715 , 
    n716 , 
    n717 , 
    n718 , 
    n719 , 
    n720 , 
    n721 , 
    n722 , 
    n723 , 
    n724 , 
    n725 , 
    n726 , 
    n727 , 
    n728 , 
    n729 , 
    n730 , 
    n731 , 
    n732 , 
    n733 , 
    n734 , 
    n735 , 
    n736 , 
    n737 , 
    n738 , 
    n739 , 
    n740 , 
    n741 , 
    n742 , 
    n743 , 
    n744 , 
    n745 , 
    n746 , 
    n747 , 
    n748 , 
    n749 , 
    n750 , 
    n751 , 
    n752 , 
    n753 , 
    n754 , 
    n755 , 
    n756 , 
    n757 , 
    n758 , 
    n759 , 
    n760 , 
    n761 , 
    n762 , 
    n763 , 
    n764 , 
    n765 , 
    n766 , 
    n767 , 
    n768 , 
    n769 , 
    n770 , 
    n771 , 
    n772 , 
    n773 , 
    n774 , 
    n775 , 
    n776 , 
    n777 , 
    n778 , 
    n779 , 
    n780 , 
    n781 , 
    n782 , 
    n783 , 
    n784 , 
    n785 , 
    n786 , 
    n787 , 
    n788 , 
    n789 , 
    n790 , 
    n791 , 
    n792 , 
    n793 , 
    n794 , 
    n795 , 
    n796 , 
    n797 , 
    n798 , 
    n799 , 
    n800 , 
    n801 , 
    n802 , 
    n803 , 
    n804 , 
    n805 , 
    n806 , 
    n807 , 
    n808 , 
    n809 , 
    n810 , 
    n811 , 
    n812 , 
    n813 , 
    n814 , 
    n815 , 
    n816 , 
    n817 , 
    n818 , 
    n819 , 
    n820 , 
    n821 , 
    n822 , 
    n823 , 
    n824 , 
    n825 , 
    n826 , 
    n827 , 
    n828 , 
    n829 , 
    n830 , 
    n831 , 
    n832 , 
    n833 , 
    n834 , 
    n835 , 
    n836 , 
    n837 , 
    n838 , 
    n839 , 
    n840 , 
    n841 , 
    n842 , 
    n843 , 
    n844 , 
    n845 , 
    n846 , 
    n847 , 
    n848 , 
    n849 , 
    n850 , 
    n851 , 
    n852 , 
    n853 , 
    n854 , 
    n855 , 
    n856 , 
    n857 , 
    n858 , 
    n859 , 
    n860 , 
    n861 , 
    n862 , 
    n863 , 
    n864 , 
    n865 , 
    n866 , 
    n867 , 
    n868 , 
    n869 , 
    n870 , 
    n871 , 
    n872 , 
    n873 , 
    n874 , 
    n875 , 
    n876 , 
    n877 , 
    n878 , 
    n879 , 
    n880 , 
    n881 , 
    n882 , 
    n883 , 
    n884 , 
    n885 , 
    n886 , 
    n887 , 
    n888 , 
    n889 , 
    n890 , 
    n891 , 
    n892 , 
    n893 , 
    n894 , 
    n895 , 
    n896 , 
    n897 , 
    n898 , 
    n899 , 
    n900 , 
    n901 , 
    n902 , 
    n903 , 
    n904 , 
    n905 , 
    n906 , 
    n907 , 
    n908 , 
    n909 , 
    n910 , 
    n911 , 
    n912 , 
    n913 , 
    n914 , 
    n915 , 
    n916 , 
    n917 , 
    n918 , 
    n919 , 
    n920 , 
    n921 , 
    n922 , 
    n923 , 
    n924 , 
    n925 , 
    n926 , 
    n927 , 
    n928 , 
    n929 , 
    n930 , 
    n931 , 
    n932 , 
    n933 , 
    n934 , 
    n935 , 
    n936 , 
    n937 , 
    n938 , 
    n939 , 
    n940 , 
    n941 , 
    n942 , 
    n943 , 
    n944 , 
    n945 , 
    n946 , 
    n947 , 
    n948 , 
    n949 , 
    n950 , 
    n951 , 
    n952 , 
    n953 , 
    n954 , 
    n955 , 
    n956 , 
    n957 , 
    n958 , 
    n959 , 
    n960 , 
    n961 , 
    n962 , 
    n963 , 
    n964 , 
    n965 , 
    n966 , 
    n967 , 
    n968 , 
    n969 , 
    n970 , 
    n971 , 
    n972 , 
    n973 , 
    n974 , 
    n975 , 
    n976 , 
    n977 , 
    n978 , 
    n979 , 
    n980 , 
    n981 , 
    n982 , 
    n983 , 
    n984 , 
    n985 , 
    n986 , 
    n987 , 
    n988 , 
    n989 , 
    n990 , 
    n991 , 
    n992 , 
    n993 , 
    n994 , 
    n995 , 
    n996 , 
    n997 , 
    n998 , 
    n999 , 
    n1000 , 
    n1001 , 
    n1002 , 
    n1003 , 
    n1004 , 
    n1005 , 
    n1006 , 
    n1007 , 
    n1008 , 
    n1009 , 
    n1010 , 
    n1011 , 
    n1012 , 
    n1013 , 
    n1014 , 
    n1015 , 
    n1016 , 
    n1017 , 
    n1018 , 
    n1019 , 
    n1020 , 
    n1021 , 
    n1022 , 
    n1023 , 
    n1024 , 
    n1025 , 
    n1026 , 
    n1027 , 
    n1028 , 
    n1029 , 
    n1030 , 
    n1031 , 
    n1032 , 
    n1033 , 
    n1034 , 
    n1035 , 
    n1036 , 
    n1037 , 
    n1038 , 
    n1039 , 
    n1040 , 
    n1041 , 
    n1042 , 
    n1043 , 
    n1044 , 
    n1045 , 
    n1046 , 
    n1047 , 
    n1048 , 
    n1049 , 
    n1050 , 
    n1051 , 
    n1052 , 
    n1053 , 
    n1054 , 
    n1055 , 
    n1056 , 
    n1057 , 
    n1058 , 
    n1059 , 
    n1060 , 
    n1061 , 
    n1062 , 
    n1063 , 
    n1064 , 
    n1065 , 
    n1066 , 
    n1067 , 
    n1068 , 
    n1069 , 
    n1070 , 
    n1071 , 
    n1072 , 
    n1073 , 
    n1074 , 
    n1075 , 
    n1076 , 
    n1077 , 
    n1078 , 
    n1079 , 
    n1080 , 
    n1081 , 
    n1082 , 
    n1083 , 
    n1084 , 
    n1085 , 
    n1086 , 
    n1087 , 
    n1088 , 
    n1089 , 
    n1090 , 
    n1091 , 
    n1092 , 
    n1093 , 
    n1094 , 
    n1095 , 
    n1096 , 
    n1097 , 
    n1098 , 
    n1099 , 
    n1100 , 
    n1101 , 
    n1102 , 
    n1103 , 
    n1104 , 
    n1105 , 
    n1106 , 
    n1107 , 
    n1108 , 
    n1109 , 
    n1110 , 
    n1111 , 
    n1112 , 
    n1113 , 
    n1114 , 
    n1115 , 
    n1116 , 
    n1117 , 
    n1118 , 
    n1119 , 
    n1120 , 
    n1121 , 
    n1122 , 
    n1123 , 
    n1124 , 
    n1125 , 
    n1126 , 
    n1127 , 
    n1128 , 
    n1129 , 
    n1130 , 
    n1131 , 
    n1132 , 
    n1133 , 
    n1134 , 
    n1135 , 
    n1136 , 
    n1137 , 
    n1138 , 
    n1139 , 
    n1140 , 
    n1141 , 
    n1142 , 
    n1143 , 
    n1144 , 
    n1145 , 
    n1146 , 
    n1147 , 
    n1148 , 
    n1149 , 
    n1150 , 
    n1151 , 
    n1152 , 
    n1153 , 
    n1154 , 
    n1155 , 
    n1156 , 
    n1157 , 
    n1158 , 
    n1159 , 
    n1160 , 
    n1161 , 
    n1162 , 
    n1163 , 
    n1164 , 
    n1165 , 
    n1166 , 
    n1167 , 
    n1168 , 
    n1169 , 
    n1170 , 
    n1171 , 
    n1172 , 
    n1173 , 
    n1174 , 
    n1175 , 
    n1176 , 
    n1177 , 
    n1178 , 
    n1179 , 
    n1180 , 
    n1181 , 
    n1182 , 
    n1183 , 
    n1184 , 
    n1185 , 
    n1186 , 
    n1187 , 
    n1188 , 
    n1189 , 
    n1190 , 
    n1191 , 
    n1192 , 
    n1193 , 
    n1194 , 
    n1195 , 
    n1196 , 
    n1197 , 
    n1198 , 
    n1199 , 
    n1200 , 
    n1201 , 
    n1202 , 
    n1203 , 
    n1204 , 
    n1205 , 
    n1206 , 
    n1207 , 
    n1208 , 
    n1209 , 
    n1210 , 
    n1211 , 
    n1212 , 
    n1213 , 
    n1214 , 
    n1215 , 
    n1216 , 
    n1217 , 
    n1218 , 
    n1219 , 
    n1220 , 
    n1221 , 
    n1222 , 
    n1223 , 
    n1224 , 
    n1225 , 
    n1226 , 
    n1227 , 
    n1228 , 
    n1229 , 
    n1230 , 
    n1231 , 
    n1232 , 
    n1233 , 
    n1234 , 
    n1235 , 
    n1236 , 
    n1237 , 
    n1238 , 
    n1239 , 
    n1240 , 
    n1241 , 
    n1242 , 
    n1243 , 
    n1244 , 
    n1245 , 
    n1246 , 
    n1247 , 
    n1248 , 
    n1249 , 
    n1250 , 
    n1251 , 
    n1252 , 
    n1253 , 
    n1254 , 
    n1255 , 
    n1256 , 
    n1257 , 
    n1258 , 
    n1259 , 
    n1260 , 
    n1261 , 
    n1262 , 
    n1263 , 
    n1264 , 
    n1265 , 
    n1266 , 
    n1267 , 
    n1268 , 
    n1269 , 
    n1270 , 
    n1271 , 
    n1272 , 
    n1273 , 
    n1274 , 
    n1275 , 
    n1276 , 
    n1277 , 
    n1278 , 
    n1279 , 
    n1280 , 
    n1281 , 
    n1282 , 
    n1283 , 
    n1284 , 
    n1285 , 
    n1286 , 
    n1287 , 
    n1288 , 
    n1289 , 
    n1290 , 
    n1291 , 
    n1292 , 
    n1293 , 
    n1294 , 
    n1295 , 
    n1296 , 
    n1297 , 
    n1298 , 
    n1299 , 
    n1300 , 
    n1301 , 
    n1302 , 
    n1303 , 
    n1304 , 
    n1305 , 
    n1306 , 
    n1307 , 
    n1308 , 
    n1309 , 
    n1310 , 
    n1311 , 
    n1312 , 
    n1313 , 
    n1314 , 
    n1315 , 
    n1316 , 
    n1317 , 
    n1318 , 
    n1319 , 
    n1320 , 
    n1321 , 
    n1322 , 
    n1323 , 
    n1324 , 
    n1325 , 
    n1326 , 
    n1327 , 
    n1328 , 
    n1329 , 
    n1330 , 
    n1331 , 
    n1332 , 
    n1333 , 
    n1334 , 
    n1335 , 
    n1336 , 
    n1337 , 
    n1338 , 
    n1339 , 
    n1340 , 
    n1341 , 
    n1342 , 
    n1343 , 
    n1344 , 
    n1345 , 
    n1346 , 
    n1347 , 
    n1348 , 
    n1349 , 
    n1350 , 
    n1351 , 
    n1352 , 
    n1353 , 
    n1354 , 
    n1355 , 
    n1356 , 
    n1357 , 
    n1358 , 
    n1359 , 
    n1360 , 
    n1361 , 
    n1362 , 
    n1363 , 
    n1364 , 
    n1365 , 
    n1366 , 
    n1367 , 
    n1368 , 
    n1369 , 
    n1370 , 
    n1371 , 
    n1372 , 
    n1373 , 
    n1374 , 
    n1375 , 
    n1376 , 
    n1377 , 
    n1378 , 
    n1379 , 
    n1380 , 
    n1381 , 
    n1382 , 
    n1383 , 
    n1384 , 
    n1385 , 
    n1386 , 
    n1387 , 
    n1388 , 
    n1389 , 
    n1390 , 
    n1391 , 
    n1392 , 
    n1393 , 
    n1394 , 
    n1395 , 
    n1396 , 
    n1397 , 
    n1398 , 
    n1399 , 
    n1400 , 
    n1401 , 
    n1402 , 
    n1403 , 
    n1404 , 
    n1405 , 
    n1406 , 
    n1407 , 
    n1408 , 
    n1409 , 
    n1410 , 
    n1411 , 
    n1412 , 
    n1413 , 
    n1414 , 
    n1415 , 
    n1416 , 
    n1417 , 
    n1418 , 
    n1419 , 
    n1420 , 
    n1421 , 
    n1422 , 
    n1423 , 
    n1424 , 
    n1425 , 
    n1426 , 
    n1427 , 
    n1428 , 
    n1429 , 
    n1430 , 
    n1431 , 
    n1432 , 
    n1433 , 
    n1434 , 
    n1435 , 
    n1436 , 
    n1437 , 
    n1438 , 
    n1439 , 
    n1440 , 
    n1441 , 
    n1442 , 
    n1443 , 
    n1444 , 
    n1445 , 
    n1446 , 
    n1447 , 
    n1448 , 
    n1449 , 
    n1450 , 
    n1451 , 
    n1452 , 
    n1453 , 
    n1454 , 
    n1455 , 
    n1456 , 
    n1457 , 
    n1458 , 
    n1459 , 
    n1460 , 
    n1461 , 
    n1462 , 
    n1463 , 
    n1464 , 
    n1465 , 
    n1466 , 
    n1467 , 
    n1468 , 
    n1469 , 
    n1470 , 
    n1471 , 
    n1472 , 
    n1473 , 
    n1474 , 
    n1475 , 
    n1476 , 
    n1477 , 
    n1478 , 
    n1479 , 
    n1480 , 
    n1481 , 
    n1482 , 
    n1483 , 
    n1484 , 
    n1485 , 
    n1486 , 
    n1487 , 
    n1488 , 
    n1489 , 
    n1490 , 
    n1491 , 
    n1492 , 
    n1493 , 
    n1494 , 
    n1495 , 
    n1496 , 
    n1497 , 
    n1498 , 
    n1499 , 
    n1500 , 
    n1501 , 
    n1502 , 
    n1503 , 
    n1504 , 
    n1505 , 
    n1506 , 
    n1507 , 
    n1508 , 
    n1509 , 
    n1510 , 
    n1511 , 
    n1512 , 
    n1513 , 
    n1514 , 
    n1515 , 
    n1516 , 
    n1517 , 
    n1518 , 
    n1519 , 
    n1520 , 
    n1521 , 
    n1522 , 
    n1523 , 
    n1524 , 
    n1525 , 
    n1526 , 
    n1527 , 
    n1528 , 
    n1529 , 
    n1530 , 
    n1531 , 
    n1532 , 
    n1533 , 
    n1534 , 
    n1535 , 
    n1536 , 
    n1537 , 
    n1538 , 
    n1539 , 
    n1540 , 
    n1541 , 
    n1542 , 
    n1543 , 
    n1544 , 
    n1545 , 
    n1546 , 
    n1547 , 
    n1548 , 
    n1549 , 
    n1550 , 
    n1551 , 
    n1552 , 
    n1553 , 
    n1554 , 
    n1555 , 
    n1556 , 
    n1557 , 
    n1558 , 
    n1559 , 
    n1560 , 
    n1561 , 
    n1562 , 
    n1563 , 
    n1564 , 
    n1565 , 
    n1566 , 
    n1567 , 
    n1568 , 
    n1569 , 
    n1570 , 
    n1571 , 
    n1572 , 
    n1573 , 
    n1574 , 
    n1575 , 
    n1576 , 
    n1577 , 
    n1578 , 
    n1579 , 
    n1580 , 
    n1581 , 
    n1582 , 
    n1583 , 
    n1584 , 
    n1585 , 
    n1586 , 
    n1587 , 
    n1588 , 
    n1589 , 
    n1590 , 
    n1591 , 
    n1592 , 
    n1593 , 
    n1594 , 
    n1595 , 
    n1596 , 
    n1597 , 
    n1598 , 
    n1599 , 
    n1600 , 
    n1601 , 
    n1602 , 
    n1603 , 
    n1604 , 
    n1605 , 
    n1606 , 
    n1607 , 
    n1608 , 
    n1609 , 
    n1610 , 
    n1611 , 
    n1612 , 
    n1613 , 
    n1614 , 
    n1615 , 
    n1616 , 
    n1617 , 
    n1618 , 
    n1619 , 
    n1620 , 
    n1621 , 
    n1622 , 
    n1623 , 
    n1624 , 
    n1625 , 
    n1626 , 
    n1627 , 
    n1628 , 
    n1629 , 
    n1630 , 
    n1631 , 
    n1632 , 
    n1633 , 
    n1634 , 
    n1635 , 
    n1636 , 
    n1637 , 
    n1638 , 
    n1639 , 
    n1640 , 
    n1641 , 
    n1642 , 
    n1643 , 
    n1644 , 
    n1645 , 
    n1646 , 
    n1647 , 
    n1648 , 
    n1649 , 
    n1650 , 
    n1651 , 
    n1652 , 
    n1653 , 
    n1654 , 
    n1655 , 
    n1656 , 
    n1657 , 
    n1658 , 
    n1659 , 
    n1660 , 
    n1661 , 
    n1662 , 
    n1663 , 
    n1664 , 
    n1665 , 
    n1666 , 
    n1667 , 
    n1668 , 
    n1669 , 
    n1670 , 
    n1671 , 
    n1672 , 
    n1673 , 
    n1674 , 
    n1675 , 
    n1676 , 
    n1677 , 
    n1678 , 
    n1679 , 
    n1680 , 
    n1681 , 
    n1682 , 
    n1683 , 
    n1684 , 
    n1685 , 
    n1686 , 
    n1687 , 
    n1688 , 
    n1689 , 
    n1690 , 
    n1691 , 
    n1692 , 
    n1693 , 
    n1694 , 
    n1695 , 
    n1696 , 
    n1697 , 
    n1698 , 
    n1699 , 
    n1700 , 
    n1701 , 
    n1702 , 
    n1703 , 
    n1704 , 
    n1705 , 
    n1706 , 
    n1707 , 
    n1708 , 
    n1709 , 
    n1710 , 
    n1711 , 
    n1712 , 
    n1713 , 
    n1714 , 
    n1715 , 
    n1716 , 
    n1717 , 
    n1718 , 
    n1719 , 
    n1720 , 
    n1721 , 
    n1722 , 
    n1723 , 
    n1724 , 
    n1725 , 
    n1726 , 
    n1727 , 
    n1728 , 
    n1729 , 
    n1730 , 
    n1731 , 
    n1732 , 
    n1733 , 
    n1734 , 
    n1735 , 
    n1736 , 
    n1737 , 
    n1738 , 
    n1739 , 
    n1740 , 
    n1741 , 
    n1742 , 
    n1743 , 
    n1744 , 
    n1745 , 
    n1746 , 
    n1747 , 
    n1748 , 
    n1749 , 
    n1750 , 
    n1751 , 
    n1752 , 
    n1753 , 
    n1754 , 
    n1755 , 
    n1756 , 
    n1757 , 
    n1758 , 
    n1759 , 
    n1760 , 
    n1761 , 
    n1762 , 
    n1763 , 
    n1764 , 
    n1765 , 
    n1766 , 
    n1767 , 
    n1768 , 
    n1769 , 
    n1770 , 
    n1771 , 
    n1772 , 
    n1773 , 
    n1774 , 
    n1775 , 
    n1776 , 
    n1777 , 
    n1778 , 
    n1779 , 
    n1780 , 
    n1781 , 
    n1782 , 
    n1783 , 
    n1784 , 
    n1785 , 
    n1786 , 
    n1787 , 
    n1788 , 
    n1789 , 
    n1790 , 
    n1791 , 
    n1792 , 
    n1793 , 
    n1794 , 
    n1795 , 
    n1796 , 
    n1797 , 
    n1798 , 
    n1799 , 
    n1800 , 
    n1801 , 
    n1802 , 
    n1803 , 
    n1804 , 
    n1805 , 
    n1806 , 
    n1807 , 
    n1808 , 
    n1809 , 
    n1810 , 
    n1811 , 
    n1812 , 
    n1813 , 
    n1814 , 
    n1815 , 
    n1816 , 
    n1817 , 
    n1818 , 
    n1819 , 
    n1820 , 
    n1821 , 
    n1822 , 
    n1823 , 
    n1824 , 
    n1825 , 
    n1826 , 
    n1827 , 
    n1828 , 
    n1829 , 
    n1830 , 
    n1831 , 
    n1832 , 
    n1833 , 
    n1834 , 
    n1835 , 
    n1836 , 
    n1837 , 
    n1838 , 
    n1839 , 
    n1840 , 
    n1841 , 
    n1842 , 
    n1843 , 
    n1844 , 
    n1845 , 
    n1846 , 
    n1847 , 
    n1848 , 
    n1849 , 
    n1850 , 
    n1851 , 
    n1852 , 
    n1853 , 
    n1854 , 
    n1855 , 
    n1856 , 
    n1857 , 
    n1858 , 
    n1859 , 
    n1860 , 
    n1861 , 
    n1862 , 
    n1863 , 
    n1864 , 
    n1865 , 
    n1866 , 
    n1867 , 
    n1868 , 
    n1869 , 
    n1870 , 
    n1871 , 
    n1872 , 
    n1873 , 
    n1874 , 
    n1875 , 
    n1876 , 
    n1877 , 
    n1878 , 
    n1879 , 
    n1880 , 
    n1881 , 
    n1882 , 
    n1883 , 
    n1884 , 
    n1885 , 
    n1886 , 
    n1887 , 
    n1888 , 
    n1889 , 
    n1890 , 
    n1891 , 
    n1892 , 
    n1893 , 
    n1894 , 
    n1895 , 
    n1896 , 
    n1897 , 
    n1898 , 
    n1899 , 
    n1900 , 
    n1901 , 
    n1902 , 
    n1903 , 
    n1904 , 
    n1905 , 
    n1906 , 
    n1907 , 
    n1908 , 
    n1909 , 
    n1910 , 
    n1911 , 
    n1912 , 
    n1913 , 
    n1914 , 
    n1915 , 
    n1916 , 
    n1917 , 
    n1918 , 
    n1919 , 
    n1920 , 
    n1921 , 
    n1922 , 
    n1923 , 
    n1924 , 
    n1925 , 
    n1926 , 
    n1927 , 
    n1928 , 
    n1929 , 
    n1930 , 
    n1931 , 
    n1932 , 
    n1933 , 
    n1934 , 
    n1935 , 
    n1936 , 
    n1937 , 
    n1938 , 
    n1939 , 
    n1940 , 
    n1941 , 
    n1942 , 
    n1943 , 
    n1944 , 
    n1945 , 
    n1946 , 
    n1947 , 
    n1948 , 
    n1949 , 
    n1950 , 
    n1951 , 
    n1952 , 
    n1953 , 
    n1954 , 
    n1955 , 
    n1956 , 
    n1957 , 
    n1958 , 
    n1959 , 
    n1960 , 
    n1961 , 
    n1962 , 
    n1963 , 
    n1964 , 
    n1965 , 
    n1966 , 
    n1967 , 
    n1968 , 
    n1969 , 
    n1970 , 
    n1971 , 
    n1972 , 
    n1973 , 
    n1974 , 
    n1975 , 
    n1976 , 
    n1977 , 
    n1978 , 
    n1979 , 
    n1980 , 
    n1981 , 
    n1982 , 
    n1983 , 
    n1984 , 
    n1985 , 
    n1986 , 
    n1987 , 
    n1988 , 
    n1989 , 
    n1990 , 
    n1991 , 
    n1992 , 
    n1993 , 
    n1994 , 
    n1995 , 
    n1996 , 
    n1997 , 
    n1998 , 
    n1999 , 
    n2000 , 
    n2001 , 
    n2002 , 
    n2003 , 
    n2004 , 
    n2005 , 
    n2006 , 
    n2007 , 
    n2008 , 
    n2009 , 
    n2010 , 
    n2011 , 
    n2012 , 
    n2013 , 
    n2014 , 
    n2015 , 
    n2016 , 
    n2017 , 
    n2018 , 
    n2019 , 
    n2020 , 
    n2021 , 
    n2022 , 
    n2023 , 
    n2024 , 
    n2025 , 
    n2026 , 
    n2027 , 
    n2028 , 
    n2029 , 
    n2030 , 
    n2031 , 
    n2032 , 
    n2033 , 
    n2034 , 
    n2035 , 
    n2036 , 
    n2037 , 
    n2038 , 
    n2039 , 
    n2040 , 
    n2041 , 
    n2042 , 
    n2043 , 
    n2044 , 
    n2045 , 
    n2046 , 
    n2047 , 
    n2048 , 
    n2049 , 
    n2050 , 
    n2051 , 
    n2052 , 
    n2053 , 
    n2054 , 
    n2055 , 
    n2056 , 
    n2057 , 
    n2058 , 
    n2059 , 
    n2060 , 
    n2061 , 
    n2062 , 
    n2063 , 
    n2064 , 
    n2065 , 
    n2066 , 
    n2067 , 
    n2068 , 
    n2069 , 
    n2070 , 
    n2071 , 
    n2072 , 
    n2073 , 
    n2074 , 
    n2075 , 
    n2076 , 
    n2077 , 
    n2078 , 
    n2079 , 
    n2080 , 
    n2081 , 
    n2082 , 
    n2083 , 
    n2084 , 
    n2085 , 
    n2086 , 
    n2087 , 
    n2088 , 
    n2089 , 
    n2090 , 
    n2091 , 
    n2092 , 
    n2093 , 
    n2094 , 
    n2095 , 
    n2096 , 
    n2097 , 
    n2098 , 
    n2099 , 
    n2100 , 
    n2101 , 
    n2102 , 
    n2103 , 
    n2104 , 
    n2105 , 
    n2106 , 
    n2107 , 
    n2108 , 
    n2109 , 
    n2110 , 
    n2111 , 
    n2112 , 
    n2113 , 
    n2114 , 
    n2115 , 
    n2116 , 
    n2117 , 
    n2118 , 
    n2119 , 
    n2120 , 
    n2121 , 
    n2122 , 
    n2123 , 
    n2124 , 
    n2125 , 
    n2126 , 
    n2127 , 
    n2128 , 
    n2129 , 
    n2130 , 
    n2131 , 
    n2132 , 
    n2133 , 
    n2134 , 
    n2135 , 
    n2136 , 
    n2137 , 
    n2138 , 
    n2139 , 
    n2140 , 
    n2141 , 
    n2142 , 
    n2143 , 
    n2144 , 
    n2145 , 
    n2146 , 
    n2147 , 
    n2148 , 
    n2149 , 
    n2150 , 
    n2151 , 
    n2152 , 
    n2153 , 
    n2154 , 
    n2155 , 
    n2156 , 
    n2157 , 
    n2158 , 
    n2159 , 
    n2160 , 
    n2161 , 
    n2162 , 
    n2163 , 
    n2164 , 
    n2165 , 
    n2166 , 
    n2167 , 
    n2168 , 
    n2169 , 
    n2170 , 
    n2171 , 
    n2172 , 
    n2173 , 
    n2174 , 
    n2175 , 
    n2176 , 
    n2177 , 
    n2178 , 
    n2179 , 
    n2180 , 
    n2181 , 
    n2182 , 
    n2183 , 
    n2184 , 
    n2185 , 
    n2186 , 
    n2187 , 
    n2188 , 
    n2189 , 
    n2190 , 
    n2191 , 
    n2192 , 
    n2193 , 
    n2194 , 
    n2195 , 
    n2196 , 
    n2197 , 
    n2198 , 
    n2199 , 
    n2200 , 
    n2201 , 
    n2202 , 
    n2203 , 
    n2204 , 
    n2205 , 
    n2206 , 
    n2207 , 
    n2208 , 
    n2209 , 
    n2210 , 
    n2211 , 
    n2212 , 
    n2213 , 
    n2214 , 
    n2215 , 
    n2216 , 
    n2217 , 
    n2218 , 
    n2219 , 
    n2220 , 
    n2221 , 
    n2222 , 
    n2223 , 
    n2224 , 
    n2225 , 
    n2226 , 
    n2227 , 
    n2228 , 
    n2229 , 
    n2230 , 
    n2231 , 
    n2232 , 
    n2233 , 
    n2234 , 
    n2235 , 
    n2236 , 
    n2237 , 
    n2238 , 
    n2239 , 
    n2240 , 
    n2241 , 
    n2242 , 
    n2243 , 
    n2244 , 
    n2245 , 
    n2246 , 
    n2247 , 
    n2248 , 
    n2249 , 
    n2250 , 
    n2251 , 
    n2252 , 
    n2253 , 
    n2254 , 
    n2255 , 
    n2256 , 
    n2257 , 
    n2258 , 
    n2259 , 
    n2260 , 
    n2261 , 
    n2262 , 
    n2263 , 
    n2264 , 
    n2265 , 
    n2266 , 
    n2267 , 
    n2268 , 
    n2269 , 
    n2270 , 
    n2271 , 
    n2272 , 
    n2273 , 
    n2274 , 
    n2275 , 
    n2276 , 
    n2277 , 
    n2278 , 
    n2279 , 
    n2280 , 
    n2281 , 
    n2282 , 
    n2283 , 
    n2284 , 
    n2285 , 
    n2286 , 
    n2287 , 
    n2288 , 
    n2289 , 
    n2290 , 
    n2291 , 
    n2292 , 
    n2293 , 
    n2294 , 
    n2295 , 
    n2296 , 
    n2297 , 
    n2298 , 
    n2299 , 
    n2300 , 
    n2301 , 
    n2302 , 
    n2303 , 
    n2304 , 
    n2305 , 
    n2306 , 
    n2307 , 
    n2308 , 
    n2309 , 
    n2310 , 
    n2311 , 
    n2312 , 
    n2313 , 
    n2314 , 
    n2315 , 
    n2316 , 
    n2317 , 
    n2318 , 
    n2319 , 
    n2320 , 
    n2321 , 
    n2322 , 
    n2323 , 
    n2324 , 
    n2325 , 
    n2326 , 
    n2327 , 
    n2328 , 
    n2329 , 
    n2330 , 
    n2331 , 
    n2332 , 
    n2333 , 
    n2334 , 
    n2335 , 
    n2336 , 
    n2337 , 
    n2338 , 
    n2339 , 
    n2340 , 
    n2341 , 
    n2342 , 
    n2343 , 
    n2344 , 
    n2345 , 
    n2346 , 
    n2347 , 
    n2348 , 
    n2349 , 
    n2350 , 
    n2351 , 
    n2352 , 
    n2353 , 
    n2354 , 
    n2355 , 
    n2356 , 
    n2357 , 
    n2358 , 
    n2359 , 
    n2360 , 
    n2361 , 
    n2362 , 
    n2363 , 
    n2364 , 
    n2365 , 
    n2366 , 
    n2367 , 
    n2368 , 
    n2369 , 
    n2370 , 
    n2371 , 
    n2372 , 
    n2373 , 
    n2374 , 
    n2375 , 
    n2376 , 
    n2377 , 
    n2378 , 
    n2379 , 
    n2380 , 
    n2381 , 
    n2382 , 
    n2383 , 
    n2384 , 
    n2385 , 
    n2386 , 
    n2387 , 
    n2388 , 
    n2389 , 
    n2390 , 
    n2391 , 
    n2392 , 
    n2393 , 
    n2394 , 
    n2395 , 
    n2396 , 
    n2397 , 
    n2398 , 
    n2399 , 
    n2400 , 
    n2401 , 
    n2402 , 
    n2403 , 
    n2404 , 
    n2405 , 
    n2406 , 
    n2407 , 
    n2408 , 
    n2409 , 
    n2410 , 
    n2411 , 
    n2412 , 
    n2413 , 
    n2414 , 
    n2415 , 
    n2416 , 
    n2417 , 
    n2418 , 
    n2419 , 
    n2420 , 
    n2421 , 
    n2422 , 
    n2423 , 
    n2424 , 
    n2425 , 
    n2426 , 
    n2427 , 
    n2428 , 
    n2429 , 
    n2430 , 
    n2431 , 
    n2432 , 
    n2433 , 
    n2434 , 
    n2435 , 
    n2436 , 
    n2437 , 
    n2438 , 
    n2439 , 
    n2440 , 
    n2441 , 
    n2442 , 
    n2443 , 
    n2444 , 
    n2445 , 
    n2446 , 
    n2447 , 
    n2448 , 
    n2449 , 
    n2450 , 
    n2451 , 
    n2452 , 
    n2453 , 
    n2454 , 
    n2455 , 
    n2456 , 
    n2457 , 
    n2458 , 
    n2459 , 
    n2460 , 
    n2461 , 
    n2462 , 
    n2463 , 
    n2464 , 
    n2465 , 
    n2466 , 
    n2467 , 
    n2468 , 
    n2469 , 
    n2470 , 
    n2471 , 
    n2472 , 
    n2473 , 
    n2474 , 
    n2475 , 
    n2476 , 
    n2477 , 
    n2478 , 
    n2479 , 
    n2480 , 
    n2481 , 
    n2482 , 
    n2483 , 
    n2484 , 
    n2485 , 
    n2486 , 
    n2487 , 
    n2488 , 
    n2489 , 
    n2490 , 
    n2491 , 
    n2492 , 
    n2493 , 
    n2494 , 
    n2495 , 
    n2496 , 
    n2497 , 
    n2498 , 
    n2499 , 
    n2500 , 
    n2501 , 
    n2502 , 
    n2503 , 
    n2504 , 
    n2505 , 
    n2506 , 
    n2507 , 
    n2508 , 
    n2509 , 
    n2510 , 
    n2511 , 
    n2512 , 
    n2513 , 
    n2514 , 
    n2515 , 
    n2516 , 
    n2517 , 
    n2518 , 
    n2519 , 
    n2520 , 
    n2521 , 
    n2522 , 
    n2523 , 
    n2524 , 
    n2525 , 
    n2526 , 
    n2527 , 
    n2528 , 
    n2529 , 
    n2530 , 
    n2531 , 
    n2532 , 
    n2533 , 
    n2534 , 
    n2535 , 
    n2536 , 
    n2537 , 
    n2538 , 
    n2539 , 
    n2540 , 
    n2541 , 
    n2542 , 
    n2543 , 
    n2544 , 
    n2545 , 
    n2546 , 
    n2547 , 
    n2548 , 
    n2549 , 
    n2550 , 
    n2551 , 
    n2552 , 
    n2553 , 
    n2554 , 
    n2555 , 
    n2556 , 
    n2557 , 
    n2558 , 
    n2559 , 
    n2560 , 
    n2561 , 
    n2562 , 
    n2563 , 
    n2564 , 
    n2565 , 
    n2566 , 
    n2567 , 
    n2568 , 
    n2569 , 
    n2570 , 
    n2571 , 
    n2572 , 
    n2573 , 
    n2574 , 
    n2575 , 
    n2576 , 
    n2577 , 
    n2578 , 
    n2579 , 
    n2580 , 
    n2581 , 
    n2582 , 
    n2583 , 
    n2584 , 
    n2585 , 
    n2586 , 
    n2587 , 
    n2588 , 
    n2589 , 
    n2590 , 
    n2591 , 
    n2592 , 
    n2593 , 
    n2594 , 
    n2595 , 
    n2596 , 
    n2597 , 
    n2598 , 
    n2599 , 
    n2600 , 
    n2601 , 
    n2602 , 
    n2603 , 
    n2604 , 
    n2605 , 
    n2606 , 
    n2607 , 
    n2608 , 
    n2609 , 
    n2610 , 
    n2611 , 
    n2612 , 
    n2613 , 
    n2614 , 
    n2615 , 
    n2616 , 
    n2617 , 
    n2618 , 
    n2619 , 
    n2620 , 
    n2621 , 
    n2622 , 
    n2623 , 
    n2624 , 
    n2625 , 
    n2626 , 
    n2627 , 
    n2628 , 
    n2629 , 
    n2630 , 
    n2631 , 
    n2632 , 
    n2633 , 
    n2634 , 
    n2635 , 
    n2636 , 
    n2637 , 
    n2638 , 
    n2639 , 
    n2640 , 
    n2641 , 
    n2642 , 
    n2643 , 
    n2644 , 
    n2645 , 
    n2646 , 
    n2647 , 
    n2648 , 
    n2649 , 
    n2650 , 
    n2651 , 
    n2652 , 
    n2653 , 
    n2654 , 
    n2655 , 
    n2656 , 
    n2657 , 
    n2658 , 
    n2659 , 
    n2660 , 
    n2661 , 
    n2662 , 
    n2663 , 
    n2664 , 
    n2665 , 
    n2666 , 
    n2667 , 
    n2668 , 
    n2669 , 
    n2670 , 
    n2671 , 
    n2672 , 
    n2673 , 
    n2674 , 
    n2675 , 
    n2676 , 
    n2677 , 
    n2678 , 
    n2679 , 
    n2680 , 
    n2681 , 
    n2682 , 
    n2683 , 
    n2684 , 
    n2685 , 
    n2686 , 
    n2687 , 
    n2688 , 
    n2689 , 
    n2690 , 
    n2691 , 
    n2692 , 
    n2693 , 
    n2694 , 
    n2695 , 
    n2696 , 
    n2697 , 
    n2698 , 
    n2699 , 
    n2700 , 
    n2701 , 
    n2702 , 
    n2703 , 
    n2704 , 
    n2705 , 
    n2706 , 
    n2707 , 
    n2708 , 
    n2709 , 
    n2710 , 
    n2711 , 
    n2712 , 
    n2713 , 
    n2714 , 
    n2715 , 
    n2716 , 
    n2717 , 
    n2718 , 
    n2719 , 
    n2720 , 
    n2721 , 
    n2722 , 
    n2723 , 
    n2724 , 
    n2725 , 
    n2726 , 
    n2727 , 
    n2728 , 
    n2729 , 
    n2730 , 
    n2731 , 
    n2732 , 
    n2733 , 
    n2734 , 
    n2735 , 
    n2736 , 
    n2737 , 
    n2738 , 
    n2739 , 
    n2740 , 
    n2741 , 
    n2742 , 
    n2743 , 
    n2744 , 
    n2745 , 
    n2746 , 
    n2747 , 
    n2748 , 
    n2749 , 
    n2750 , 
    n2751 , 
    n2752 , 
    n2753 , 
    n2754 , 
    n2755 , 
    n2756 , 
    n2757 , 
    n2758 , 
    n2759 , 
    n2760 , 
    n2761 , 
    n2762 , 
    n2763 , 
    n2764 , 
    n2765 , 
    n2766 , 
    n2767 , 
    n2768 , 
    n2769 , 
    n2770 , 
    n2771 , 
    n2772 , 
    n2773 , 
    n2774 , 
    n2775 , 
    n2776 , 
    n2777 , 
    n2778 , 
    n2779 , 
    n2780 , 
    n2781 , 
    n2782 , 
    n2783 , 
    n2784 , 
    n2785 , 
    n2786 , 
    n2787 , 
    n2788 , 
    n2789 , 
    n2790 , 
    n2791 , 
    n2792 , 
    n2793 , 
    n2794 , 
    n2795 , 
    n2796 , 
    n2797 , 
    n2798 , 
    n2799 , 
    n2800 , 
    n2801 , 
    n2802 , 
    n2803 , 
    n2804 , 
    n2805 , 
    n2806 , 
    n2807 , 
    n2808 , 
    n2809 , 
    n2810 , 
    n2811 , 
    n2812 , 
    n2813 , 
    n2814 , 
    n2815 , 
    n2816 , 
    n2817 , 
    n2818 , 
    n2819 , 
    n2820 , 
    n2821 , 
    n2822 , 
    n2823 , 
    n2824 , 
    n2825 , 
    n2826 , 
    n2827 , 
    n2828 , 
    n2829 , 
    n2830 , 
    n2831 , 
    n2832 , 
    n2833 , 
    n2834 , 
    n2835 , 
    n2836 , 
    n2837 , 
    n2838 , 
    n2839 , 
    n2840 , 
    n2841 , 
    n2842 , 
    n2843 , 
    n2844 , 
    n2845 , 
    n2846 , 
    n2847 , 
    n2848 , 
    n2849 , 
    n2850 , 
    n2851 , 
    n2852 , 
    n2853 , 
    n2854 , 
    n2855 , 
    n2856 , 
    n2857 , 
    n2858 , 
    n2859 , 
    n2860 , 
    n2861 , 
    n2862 , 
    n2863 , 
    n2864 , 
    n2865 , 
    n2866 , 
    n2867 , 
    n2868 , 
    n2869 , 
    n2870 , 
    n2871 , 
    n2872 , 
    n2873 , 
    n2874 , 
    n2875 , 
    n2876 , 
    n2877 , 
    n2878 , 
    n2879 , 
    n2880 , 
    n2881 , 
    n2882 , 
    n2883 , 
    n2884 , 
    n2885 , 
    n2886 , 
    n2887 , 
    n2888 , 
    n2889 , 
    n2890 , 
    n2891 , 
    n2892 , 
    n2893 , 
    n2894 , 
    n2895 , 
    n2896 , 
    n2897 , 
    n2898 , 
    n2899 , 
    n2900 , 
    n2901 , 
    n2902 , 
    n2903 , 
    n2904 , 
    n2905 , 
    n2906 , 
    n2907 , 
    n2908 , 
    n2909 , 
    n2910 , 
    n2911 , 
    n2912 , 
    n2913 , 
    n2914 , 
    n2915 , 
    n2916 , 
    n2917 , 
    n2918 , 
    n2919 , 
    n2920 , 
    n2921 , 
    n2922 , 
    n2923 , 
    n2924 , 
    n2925 , 
    n2926 , 
    n2927 , 
    n2928 , 
    n2929 , 
    n2930 , 
    n2931 , 
    n2932 , 
    n2933 , 
    n2934 , 
    n2935 , 
    n2936 , 
    n2937 , 
    n2938 , 
    n2939 , 
    n2940 , 
    n2941 , 
    n2942 , 
    n2943 , 
    n2944 , 
    n2945 , 
    n2946 , 
    n2947 , 
    n2948 , 
    n2949 , 
    n2950 , 
    n2951 , 
    n2952 , 
    n2953 , 
    n2954 , 
    n2955 , 
    n2956 , 
    n2957 , 
    n2958 , 
    n2959 , 
    n2960 , 
    n2961 , 
    n2962 , 
    n2963 , 
    n2964 , 
    n2965 , 
    n2966 , 
    n2967 , 
    n2968 , 
    n2969 , 
    n2970 , 
    n2971 , 
    n2972 , 
    n2973 , 
    n2974 , 
    n2975 , 
    n2976 , 
    n2977 , 
    n2978 , 
    n2979 , 
    n2980 , 
    n2981 , 
    n2982 , 
    n2983 , 
    n2984 , 
    n2985 , 
    n2986 , 
    n2987 , 
    n2988 , 
    n2989 , 
    n2990 , 
    n2991 , 
    n2992 , 
    n2993 , 
    n2994 , 
    n2995 , 
    n2996 , 
    n2997 , 
    n2998 , 
    n2999 , 
    n3000 , 
    n3001 , 
    n3002 , 
    n3003 , 
    n3004 , 
    n3005 , 
    n3006 , 
    n3007 , 
    n3008 , 
    n3009 , 
    n3010 , 
    n3011 , 
    n3012 , 
    n3013 , 
    n3014 , 
    n3015 , 
    n3016 , 
    n3017 , 
    n3018 , 
    n3019 , 
    n3020 , 
    n3021 , 
    n3022 , 
    n3023 , 
    n3024 , 
    n3025 , 
    n3026 , 
    n3027 , 
    n3028 , 
    n3029 , 
    n3030 , 
    n3031 , 
    n3032 , 
    n3033 , 
    n3034 , 
    n3035 , 
    n3036 , 
    n3037 , 
    n3038 , 
    n3039 , 
    n3040 , 
    n3041 , 
    n3042 , 
    n3043 , 
    n3044 , 
    n3045 , 
    n3046 , 
    n3047 , 
    n3048 , 
    n3049 , 
    n3050 , 
    n3051 , 
    n3052 , 
    n3053 , 
    n3054 , 
    n3055 , 
    n3056 , 
    n3057 , 
    n3058 , 
    n3059 , 
    n3060 , 
    n3061 , 
    n3062 , 
    n3063 , 
    n3064 , 
    n3065 , 
    n3066 , 
    n3067 , 
    n3068 , 
    n3069 , 
    n3070 , 
    n3071 , 
    n3072 , 
    n3073 , 
    n3074 , 
    n3075 , 
    n3076 , 
    n3077 , 
    n3078 , 
    n3079 , 
    n3080 , 
    n3081 , 
    n3082 , 
    n3083 , 
    n3084 , 
    n3085 , 
    n3086 , 
    n3087 , 
    n3088 , 
    n3089 , 
    n3090 , 
    n3091 , 
    n3092 , 
    n3093 , 
    n3094 , 
    n3095 , 
    n3096 , 
    n3097 , 
    n3098 , 
    n3099 , 
    n3100 , 
    n3101 , 
    n3102 , 
    n3103 , 
    n3104 , 
    n3105 , 
    n3106 , 
    n3107 , 
    n3108 , 
    n3109 , 
    n3110 , 
    n3111 , 
    n3112 , 
    n3113 , 
    n3114 , 
    n3115 , 
    n3116 , 
    n3117 , 
    n3118 , 
    n3119 , 
    n3120 , 
    n3121 , 
    n3122 , 
    n3123 , 
    n3124 , 
    n3125 , 
    n3126 , 
    n3127 , 
    n3128 , 
    n3129 , 
    n3130 , 
    n3131 , 
    n3132 , 
    n3133 , 
    n3134 , 
    n3135 , 
    n3136 , 
    n3137 , 
    n3138 , 
    n3139 , 
    n3140 , 
    n3141 , 
    n3142 , 
    n3143 , 
    n3144 , 
    n3145 , 
    n3146 , 
    n3147 , 
    n3148 , 
    n3149 , 
    n3150 , 
    n3151 , 
    n3152 , 
    n3153 , 
    n3154 , 
    n3155 , 
    n3156 , 
    n3157 , 
    n3158 , 
    n3159 , 
    n3160 , 
    n3161 , 
    n3162 , 
    n3163 , 
    n3164 , 
    n3165 , 
    n3166 , 
    n3167 , 
    n3168 , 
    n3169 , 
    n3170 , 
    n3171 , 
    n3172 , 
    n3173 , 
    n3174 , 
    n3175 , 
    n3176 , 
    n3177 , 
    n3178 , 
    n3179 , 
    n3180 , 
    n3181 , 
    n3182 , 
    n3183 , 
    n3184 , 
    n3185 , 
    n3186 , 
    n3187 , 
    n3188 , 
    n3189 , 
    n3190 , 
    n3191 , 
    n3192 , 
    n3193 , 
    n3194 , 
    n3195 , 
    n3196 , 
    n3197 , 
    n3198 , 
    n3199 , 
    n3200 , 
    n3201 , 
    n3202 , 
    n3203 , 
    n3204 , 
    n3205 , 
    n3206 , 
    n3207 , 
    n3208 , 
    n3209 , 
    n3210 , 
    n3211 , 
    n3212 , 
    n3213 , 
    n3214 , 
    n3215 , 
    n3216 , 
    n3217 , 
    n3218 , 
    n3219 , 
    n3220 , 
    n3221 , 
    n3222 , 
    n3223 , 
    n3224 , 
    n3225 , 
    n3226 , 
    n3227 , 
    n3228 , 
    n3229 , 
    n3230 , 
    n3231 , 
    n3232 , 
    n3233 , 
    n3234 , 
    n3235 , 
    n3236 , 
    n3237 , 
    n3238 , 
    n3239 , 
    n3240 , 
    n3241 , 
    n3242 , 
    n3243 , 
    n3244 , 
    n3245 , 
    n3246 , 
    n3247 , 
    n3248 , 
    n3249 , 
    n3250 , 
    n3251 , 
    n3252 , 
    n3253 , 
    n3254 , 
    n3255 , 
    n3256 , 
    n3257 , 
    n3258 , 
    n3259 , 
    n3260 , 
    n3261 , 
    n3262 , 
    n3263 , 
    n3264 , 
    n3265 , 
    n3266 , 
    n3267 , 
    n3268 , 
    n3269 , 
    n3270 , 
    n3271 , 
    n3272 , 
    n3273 , 
    n3274 , 
    n3275 , 
    n3276 , 
    n3277 , 
    n3278 , 
    n3279 , 
    n3280 , 
    n3281 , 
    n3282 , 
    n3283 , 
    n3284 , 
    n3285 , 
    n3286 , 
    n3287 , 
    n3288 , 
    n3289 , 
    n3290 , 
    n3291 , 
    n3292 , 
    n3293 , 
    n3294 , 
    n3295 , 
    n3296 , 
    n3297 , 
    n3298 , 
    n3299 , 
    n3300 , 
    n3301 , 
    n3302 , 
    n3303 , 
    n3304 , 
    n3305 , 
    n3306 , 
    n3307 , 
    n3308 , 
    n3309 , 
    n3310 , 
    n3311 , 
    n3312 , 
    n3313 , 
    n3314 , 
    n3315 , 
    n3316 , 
    n3317 , 
    n3318 , 
    n3319 , 
    n3320 , 
    n3321 , 
    n3322 , 
    n3323 , 
    n3324 , 
    n3325 , 
    n3326 , 
    n3327 , 
    n3328 , 
    n3329 , 
    n3330 , 
    n3331 , 
    n3332 , 
    n3333 , 
    n3334 , 
    n3335 , 
    n3336 , 
    n3337 , 
    n3338 , 
    n3339 , 
    n3340 , 
    n3341 , 
    n3342 , 
    n3343 , 
    n3344 , 
    n3345 , 
    n3346 , 
    n3347 , 
    n3348 , 
    n3349 , 
    n3350 , 
    n3351 , 
    n3352 , 
    n3353 , 
    n3354 , 
    n3355 , 
    n3356 , 
    n3357 , 
    n3358 , 
    n3359 , 
    n3360 , 
    n3361 , 
    n3362 , 
    n3363 , 
    n3364 , 
    n3365 , 
    n3366 , 
    n3367 , 
    n3368 , 
    n3369 , 
    n3370 , 
    n3371 , 
    n3372 , 
    n3373 , 
    n3374 , 
    n3375 , 
    n3376 , 
    n3377 , 
    n3378 , 
    n3379 , 
    n3380 , 
    n3381 , 
    n3382 , 
    n3383 , 
    n3384 , 
    n3385 , 
    n3386 , 
    n3387 , 
    n3388 , 
    n3389 , 
    n3390 , 
    n3391 , 
    n3392 , 
    n3393 , 
    n3394 , 
    n3395 , 
    n3396 , 
    n3397 , 
    n3398 , 
    n3399 , 
    n3400 , 
    n3401 , 
    n3402 , 
    n3403 , 
    n3404 , 
    n3405 , 
    n3406 , 
    n3407 , 
    n3408 , 
    n3409 , 
    n3410 , 
    n3411 , 
    n3412 , 
    n3413 , 
    n3414 , 
    n3415 , 
    n3416 , 
    n3417 , 
    n3418 , 
    n3419 , 
    n3420 , 
    n3421 , 
    n3422 , 
    n3423 , 
    n3424 , 
    n3425 , 
    n3426 , 
    n3427 , 
    n3428 , 
    n3429 , 
    n3430 , 
    n3431 , 
    n3432 , 
    n3433 , 
    n3434 , 
    n3435 , 
    n3436 , 
    n3437 , 
    n3438 , 
    n3439 , 
    n3440 , 
    n3441 , 
    n3442 , 
    n3443 , 
    n3444 , 
    n3445 , 
    n3446 , 
    n3447 , 
    n3448 , 
    n3449 , 
    n3450 , 
    n3451 , 
    n3452 , 
    n3453 , 
    n3454 , 
    n3455 , 
    n3456 , 
    n3457 , 
    n3458 , 
    n3459 , 
    n3460 , 
    n3461 , 
    n3462 , 
    n3463 , 
    n3464 , 
    n3465 , 
    n3466 , 
    n3467 , 
    n3468 , 
    n3469 , 
    n3470 , 
    n3471 , 
    n3472 , 
    n3473 , 
    n3474 , 
    n3475 , 
    n3476 , 
    n3477 , 
    n3478 , 
    n3479 , 
    n3480 , 
    n3481 , 
    n3482 , 
    n3483 , 
    n3484 , 
    n3485 , 
    n3486 , 
    n3487 , 
    n3488 , 
    n3489 , 
    n3490 , 
    n3491 , 
    n3492 , 
    n3493 , 
    n3494 , 
    n3495 , 
    n3496 , 
    n3497 , 
    n3498 , 
    n3499 , 
    n3500 , 
    n3501 , 
    n3502 , 
    n3503 , 
    n3504 , 
    n3505 , 
    n3506 , 
    n3507 , 
    n3508 , 
    n3509 , 
    n3510 , 
    n3511 , 
    n3512 , 
    n3513 , 
    n3514 , 
    n3515 , 
    n3516 , 
    n3517 , 
    n3518 , 
    n3519 , 
    n3520 , 
    n3521 , 
    n3522 , 
    n3523 , 
    n3524 , 
    n3525 , 
    n3526 , 
    n3527 , 
    n3528 , 
    n3529 , 
    n3530 , 
    n3531 , 
    n3532 , 
    n3533 , 
    n3534 , 
    n3535 , 
    n3536 , 
    n3537 , 
    n3538 , 
    n3539 , 
    n3540 , 
    n3541 , 
    n3542 , 
    n3543 , 
    n3544 , 
    n3545 , 
    n3546 , 
    n3547 , 
    n3548 , 
    n3549 , 
    n3550 , 
    n3551 , 
    n3552 , 
    n3553 , 
    n3554 , 
    n3555 , 
    n3556 , 
    n3557 , 
    n3558 , 
    n3559 , 
    n3560 , 
    n3561 , 
    n3562 , 
    n3563 , 
    n3564 , 
    n3565 , 
    n3566 , 
    n3567 , 
    n3568 , 
    n3569 , 
    n3570 , 
    n3571 , 
    n3572 , 
    n3573 , 
    n3574 , 
    n3575 , 
    n3576 , 
    n3577 , 
    n3578 , 
    n3579 , 
    n3580 , 
    n3581 , 
    n3582 , 
    n3583 , 
    n3584 , 
    n3585 , 
    n3586 , 
    n3587 , 
    n3588 , 
    n3589 , 
    n3590 , 
    n3591 , 
    n3592 , 
    n3593 , 
    n3594 , 
    n3595 , 
    n3596 , 
    n3597 , 
    n3598 , 
    n3599 , 
    n3600 , 
    n3601 , 
    n3602 , 
    n3603 , 
    n3604 , 
    n3605 , 
    n3606 , 
    n3607 , 
    n3608 , 
    n3609 , 
    n3610 , 
    n3611 , 
    n3612 , 
    n3613 , 
    n3614 , 
    n3615 , 
    n3616 , 
    n3617 , 
    n3618 , 
    n3619 , 
    n3620 , 
    n3621 , 
    n3622 , 
    n3623 , 
    n3624 , 
    n3625 , 
    n3626 , 
    n3627 , 
    n3628 , 
    n3629 , 
    n3630 , 
    n3631 , 
    n3632 , 
    n3633 , 
    n3634 , 
    n3635 , 
    n3636 , 
    n3637 , 
    n3638 , 
    n3639 , 
    n3640 , 
    n3641 , 
    n3642 , 
    n3643 , 
    n3644 , 
    n3645 , 
    n3646 , 
    n3647 , 
    n3648 , 
    n3649 , 
    n3650 , 
    n3651 , 
    n3652 , 
    n3653 , 
    n3654 , 
    n3655 , 
    n3656 , 
    n3657 , 
    n3658 , 
    n3659 , 
    n3660 , 
    n3661 , 
    n3662 , 
    n3663 , 
    n3664 , 
    n3665 , 
    n3666 , 
    n3667 , 
    n3668 , 
    n3669 , 
    n3670 , 
    n3671 , 
    n3672 , 
    n3673 , 
    n3674 , 
    n3675 , 
    n3676 , 
    n3677 , 
    n3678 , 
    n3679 , 
    n3680 , 
    n3681 , 
    n3682 , 
    n3683 , 
    n3684 , 
    n3685 , 
    n3686 , 
    n3687 , 
    n3688 , 
    n3689 , 
    n3690 , 
    n3691 , 
    n3692 , 
    n3693 , 
    n3694 , 
    n3695 , 
    n3696 , 
    n3697 , 
    n3698 , 
    n3699 , 
    n3700 , 
    n3701 , 
    n3702 , 
    n3703 , 
    n3704 , 
    n3705 , 
    n3706 , 
    n3707 , 
    n3708 , 
    n3709 , 
    n3710 , 
    n3711 , 
    n3712 , 
    n3713 , 
    n3714 , 
    n3715 , 
    n3716 , 
    n3717 , 
    n3718 , 
    n3719 , 
    n3720 , 
    n3721 , 
    n3722 , 
    n3723 , 
    n3724 , 
    n3725 , 
    n3726 , 
    n3727 , 
    n3728 , 
    n3729 , 
    n3730 , 
    n3731 , 
    n3732 , 
    n3733 , 
    n3734 , 
    n3735 , 
    n3736 , 
    n3737 , 
    n3738 , 
    n3739 , 
    n3740 , 
    n3741 , 
    n3742 , 
    n3743 , 
    n3744 , 
    n3745 , 
    n3746 , 
    n3747 , 
    n3748 , 
    n3749 , 
    n3750 , 
    n3751 , 
    n3752 , 
    n3753 , 
    n3754 , 
    n3755 , 
    n3756 , 
    n3757 , 
    n3758 , 
    n3759 , 
    n3760 , 
    n3761 , 
    n3762 , 
    n3763 , 
    n3764 , 
    n3765 , 
    n3766 , 
    n3767 , 
    n3768 , 
    n3769 , 
    n3770 , 
    n3771 , 
    n3772 , 
    n3773 , 
    n3774 , 
    n3775 , 
    n3776 , 
    n3777 , 
    n3778 , 
    n3779 , 
    n3780 , 
    n3781 , 
    n3782 , 
    n3783 , 
    n3784 , 
    n3785 , 
    n3786 , 
    n3787 , 
    n3788 , 
    n3789 , 
    n3790 , 
    n3791 , 
    n3792 , 
    n3793 , 
    n3794 , 
    n3795 , 
    n3796 , 
    n3797 , 
    n3798 , 
    n3799 , 
    n3800 , 
    n3801 , 
    n3802 , 
    n3803 , 
    n3804 , 
    n3805 , 
    n3806 , 
    n3807 , 
    n3808 , 
    n3809 , 
    n3810 , 
    n3811 , 
    n3812 , 
    n3813 , 
    n3814 , 
    n3815 , 
    n3816 , 
    n3817 , 
    n3818 , 
    n3819 , 
    n3820 , 
    n3821 , 
    n3822 , 
    n3823 , 
    n3824 , 
    n3825 , 
    n3826 , 
    n3827 , 
    n3828 , 
    n3829 , 
    n3830 , 
    n3831 , 
    n3832 , 
    n3833 , 
    n3834 , 
    n3835 , 
    n3836 , 
    n3837 , 
    n3838 , 
    n3839 , 
    n3840 , 
    n3841 , 
    n3842 , 
    n3843 , 
    n3844 , 
    n3845 , 
    n3846 , 
    n3847 , 
    n3848 , 
    n3849 , 
    n3850 , 
    n3851 , 
    n3852 , 
    n3853 , 
    n3854 , 
    n3855 , 
    n3856 , 
    n3857 , 
    n3858 , 
    n3859 , 
    n3860 , 
    n3861 , 
    n3862 , 
    n3863 , 
    n3864 , 
    n3865 , 
    n3866 , 
    n3867 , 
    n3868 , 
    n3869 , 
    n3870 , 
    n3871 , 
    n3872 , 
    n3873 , 
    n3874 , 
    n3875 , 
    n3876 , 
    n3877 , 
    n3878 , 
    n3879 , 
    n3880 , 
    n3881 , 
    n3882 , 
    n3883 , 
    n3884 , 
    n3885 , 
    n3886 , 
    n3887 , 
    n3888 , 
    n3889 , 
    n3890 , 
    n3891 , 
    n3892 , 
    n3893 , 
    n3894 , 
    n3895 , 
    n3896 , 
    n3897 , 
    n3898 , 
    n3899 , 
    n3900 , 
    n3901 , 
    n3902 , 
    n3903 , 
    n3904 , 
    n3905 , 
    n3906 , 
    n3907 , 
    n3908 , 
    n3909 , 
    n3910 , 
    n3911 , 
    n3912 , 
    n3913 , 
    n3914 , 
    n3915 , 
    n3916 , 
    n3917 , 
    n3918 , 
    n3919 , 
    n3920 , 
    n3921 , 
    n3922 , 
    n3923 , 
    n3924 , 
    n3925 , 
    n3926 , 
    n3927 , 
    n3928 , 
    n3929 , 
    n3930 , 
    n3931 , 
    n3932 , 
    n3933 , 
    n3934 , 
    n3935 , 
    n3936 , 
    n3937 , 
    n3938 , 
    n3939 , 
    n3940 , 
    n3941 , 
    n3942 , 
    n3943 , 
    n3944 , 
    n3945 , 
    n3946 , 
    n3947 , 
    n3948 , 
    n3949 , 
    n3950 , 
    n3951 , 
    n3952 , 
    n3953 , 
    n3954 , 
    n3955 , 
    n3956 , 
    n3957 , 
    n3958 , 
    n3959 , 
    n3960 , 
    n3961 , 
    n3962 , 
    n3963 , 
    n3964 , 
    n3965 , 
    n3966 , 
    n3967 , 
    n3968 , 
    n3969 , 
    n3970 , 
    n3971 , 
    n3972 , 
    n3973 , 
    n3974 , 
    n3975 , 
    n3976 , 
    n3977 , 
    n3978 , 
    n3979 , 
    n3980 , 
    n3981 , 
    n3982 , 
    n3983 , 
    n3984 , 
    n3985 , 
    n3986 , 
    n3987 , 
    n3988 , 
    n3989 , 
    n3990 , 
    n3991 , 
    n3992 , 
    n3993 , 
    n3994 , 
    n3995 , 
    n3996 , 
    n3997 , 
    n3998 , 
    n3999 , 
    n4000 , 
    n4001 , 
    n4002 , 
    n4003 , 
    n4004 , 
    n4005 , 
    n4006 , 
    n4007 , 
    n4008 , 
    n4009 , 
    n4010 , 
    n4011 , 
    n4012 , 
    n4013 , 
    n4014 , 
    n4015 , 
    n4016 , 
    n4017 , 
    n4018 , 
    n4019 , 
    n4020 , 
    n4021 , 
    n4022 , 
    n4023 , 
    n4024 , 
    n4025 , 
    n4026 , 
    n4027 , 
    n4028 , 
    n4029 , 
    n4030 , 
    n4031 , 
    n4032 , 
    n4033 , 
    n4034 , 
    n4035 , 
    n4036 , 
    n4037 , 
    n4038 , 
    n4039 , 
    n4040 , 
    n4041 , 
    n4042 , 
    n4043 , 
    n4044 , 
    n4045 , 
    n4046 , 
    n4047 , 
    n4048 , 
    n4049 , 
    n4050 , 
    n4051 , 
    n4052 , 
    n4053 , 
    n4054 , 
    n4055 , 
    n4056 , 
    n4057 , 
    n4058 , 
    n4059 , 
    n4060 , 
    n4061 , 
    n4062 , 
    n4063 , 
    n4064 , 
    n4065 , 
    n4066 , 
    n4067 , 
    n4068 , 
    n4069 , 
    n4070 , 
    n4071 , 
    n4072 , 
    n4073 , 
    n4074 , 
    n4075 , 
    n4076 , 
    n4077 , 
    n4078 , 
    n4079 , 
    n4080 , 
    n4081 , 
    n4082 , 
    n4083 , 
    n4084 , 
    n4085 , 
    n4086 , 
    n4087 , 
    n4088 , 
    n4089 , 
    n4090 , 
    n4091 , 
    n4092 , 
    n4093 , 
    n4094 , 
    n4095 , 
    n4096 , 
    n4097 , 
    n4098 , 
    n4099 , 
    n4100 , 
    n4101 , 
    n4102 , 
    n4103 , 
    n4104 , 
    n4105 , 
    n4106 , 
    n4107 , 
    n4108 , 
    n4109 , 
    n4110 , 
    n4111 , 
    n4112 , 
    n4113 , 
    n4114 , 
    n4115 , 
    n4116 , 
    n4117 , 
    n4118 , 
    n4119 , 
    n4120 , 
    n4121 , 
    n4122 , 
    n4123 , 
    n4124 , 
    n4125 , 
    n4126 , 
    n4127 , 
    n4128 , 
    n4129 , 
    n4130 , 
    n4131 , 
    n4132 , 
    n4133 , 
    n4134 , 
    n4135 , 
    n4136 , 
    n4137 , 
    n4138 , 
    n4139 , 
    n4140 , 
    n4141 , 
    n4142 , 
    n4143 , 
    n4144 , 
    n4145 , 
    n4146 , 
    n4147 , 
    n4148 , 
    n4149 , 
    n4150 , 
    n4151 , 
    n4152 , 
    n4153 , 
    n4154 , 
    n4155 , 
    n4156 , 
    n4157 , 
    n4158 , 
    n4159 , 
    n4160 , 
    n4161 , 
    n4162 , 
    n4163 , 
    n4164 , 
    n4165 , 
    n4166 , 
    n4167 , 
    n4168 , 
    n4169 , 
    n4170 , 
    n4171 , 
    n4172 , 
    n4173 , 
    n4174 , 
    n4175 , 
    n4176 , 
    n4177 , 
    n4178 , 
    n4179 , 
    n4180 , 
    n4181 , 
    n4182 , 
    n4183 , 
    n4184 , 
    n4185 , 
    n4186 , 
    n4187 , 
    n4188 , 
    n4189 , 
    n4190 , 
    n4191 , 
    n4192 , 
    n4193 , 
    n4194 , 
    n4195 , 
    n4196 , 
    n4197 , 
    n4198 , 
    n4199 , 
    n4200 , 
    n4201 , 
    n4202 , 
    n4203 , 
    n4204 , 
    n4205 , 
    n4206 , 
    n4207 , 
    n4208 , 
    n4209 , 
    n4210 , 
    n4211 , 
    n4212 , 
    n4213 , 
    n4214 , 
    n4215 , 
    n4216 , 
    n4217 , 
    n4218 , 
    n4219 , 
    n4220 , 
    n4221 , 
    n4222 , 
    n4223 , 
    n4224 , 
    n4225 , 
    n4226 , 
    n4227 , 
    n4228 , 
    n4229 , 
    n4230 , 
    n4231 , 
    n4232 , 
    n4233 , 
    n4234 , 
    n4235 , 
    n4236 , 
    n4237 , 
    n4238 , 
    n4239 , 
    n4240 , 
    n4241 , 
    n4242 , 
    n4243 , 
    n4244 , 
    n4245 , 
    n4246 , 
    n4247 , 
    n4248 , 
    n4249 , 
    n4250 , 
    n4251 , 
    n4252 , 
    n4253 , 
    n4254 , 
    n4255 , 
    n4256 , 
    n4257 , 
    n4258 , 
    n4259 , 
    n4260 , 
    n4261 , 
    n4262 , 
    n4263 , 
    n4264 , 
    n4265 , 
    n4266 , 
    n4267 , 
    n4268 , 
    n4269 , 
    n4270 , 
    n4271 , 
    n4272 , 
    n4273 , 
    n4274 , 
    n4275 , 
    n4276 , 
    n4277 , 
    n4278 , 
    n4279 , 
    n4280 , 
    n4281 , 
    n4282 , 
    n4283 , 
    n4284 , 
    n4285 , 
    n4286 , 
    n4287 , 
    n4288 , 
    n4289 , 
    n4290 , 
    n4291 , 
    n4292 , 
    n4293 , 
    n4294 , 
    n4295 , 
    n4296 , 
    n4297 , 
    n4298 , 
    n4299 , 
    n4300 , 
    n4301 , 
    n4302 , 
    n4303 , 
    n4304 , 
    n4305 , 
    n4306 , 
    n4307 , 
    n4308 , 
    n4309 , 
    n4310 , 
    n4311 , 
    n4312 , 
    n4313 , 
    n4314 , 
    n4315 , 
    n4316 , 
    n4317 , 
    n4318 , 
    n4319 , 
    n4320 , 
    n4321 , 
    n4322 , 
    n4323 , 
    n4324 , 
    n4325 , 
    n4326 , 
    n4327 , 
    n4328 , 
    n4329 , 
    n4330 , 
    n4331 , 
    n4332 , 
    n4333 , 
    n4334 , 
    n4335 , 
    n4336 , 
    n4337 , 
    n4338 , 
    n4339 , 
    n4340 , 
    n4341 , 
    n4342 , 
    n4343 , 
    n4344 , 
    n4345 , 
    n4346 , 
    n4347 , 
    n4348 , 
    n4349 , 
    n4350 , 
    n4351 , 
    n4352 , 
    n4353 , 
    n4354 , 
    n4355 , 
    n4356 , 
    n4357 , 
    n4358 , 
    n4359 , 
    n4360 , 
    n4361 , 
    n4362 , 
    n4363 , 
    n4364 , 
    n4365 , 
    n4366 , 
    n4367 , 
    n4368 , 
    n4369 , 
    n4370 , 
    n4371 , 
    n4372 , 
    n4373 , 
    n4374 , 
    n4375 , 
    n4376 , 
    n4377 , 
    n4378 , 
    n4379 , 
    n4380 , 
    n4381 , 
    n4382 , 
    n4383 , 
    n4384 , 
    n4385 , 
    n4386 , 
    n4387 , 
    n4388 , 
    n4389 , 
    n4390 , 
    n4391 , 
    n4392 , 
    n4393 , 
    n4394 , 
    n4395 , 
    n4396 , 
    n4397 , 
    n4398 , 
    n4399 , 
    n4400 , 
    n4401 , 
    n4402 , 
    n4403 , 
    n4404 , 
    n4405 , 
    n4406 , 
    n4407 , 
    n4408 , 
    n4409 , 
    n4410 , 
    n4411 , 
    n4412 , 
    n4413 , 
    n4414 , 
    n4415 , 
    n4416 , 
    n4417 , 
    n4418 , 
    n4419 , 
    n4420 , 
    n4421 , 
    n4422 , 
    n4423 , 
    n4424 , 
    n4425 , 
    n4426 , 
    n4427 , 
    n4428 , 
    n4429 , 
    n4430 , 
    n4431 , 
    n4432 , 
    n4433 , 
    n4434 , 
    n4435 , 
    n4436 , 
    n4437 , 
    n4438 , 
    n4439 , 
    n4440 , 
    n4441 , 
    n4442 , 
    n4443 , 
    n4444 , 
    n4445 , 
    n4446 , 
    n4447 , 
    n4448 , 
    n4449 , 
    n4450 , 
    n4451 , 
    n4452 , 
    n4453 , 
    n4454 , 
    n4455 , 
    n4456 , 
    n4457 , 
    n4458 , 
    n4459 , 
    n4460 , 
    n4461 , 
    n4462 , 
    n4463 , 
    n4464 , 
    n4465 , 
    n4466 , 
    n4467 , 
    n4468 , 
    n4469 , 
    n4470 , 
    n4471 , 
    n4472 , 
    n4473 , 
    n4474 , 
    n4475 , 
    n4476 , 
    n4477 , 
    n4478 , 
    n4479 , 
    n4480 , 
    n4481 , 
    n4482 , 
    n4483 , 
    n4484 , 
    n4485 , 
    n4486 , 
    n4487 , 
    n4488 , 
    n4489 , 
    n4490 , 
    n4491 , 
    n4492 , 
    n4493 , 
    n4494 , 
    n4495 , 
    n4496 , 
    n4497 , 
    n4498 , 
    n4499 , 
    n4500 , 
    n4501 , 
    n4502 , 
    n4503 , 
    n4504 , 
    n4505 , 
    n4506 , 
    n4507 , 
    n4508 , 
    n4509 , 
    n4510 , 
    n4511 , 
    n4512 , 
    n4513 , 
    n4514 , 
    n4515 , 
    n4516 , 
    n4517 , 
    n4518 , 
    n4519 , 
    n4520 , 
    n4521 , 
    n4522 , 
    n4523 , 
    n4524 , 
    n4525 , 
    n4526 , 
    n4527 , 
    n4528 , 
    n4529 , 
    n4530 , 
    n4531 , 
    n4532 , 
    n4533 , 
    n4534 , 
    n4535 , 
    n4536 , 
    n4537 , 
    n4538 , 
    n4539 , 
    n4540 , 
    n4541 , 
    n4542 , 
    n4543 , 
    n4544 , 
    n4545 , 
    n4546 , 
    n4547 , 
    n4548 , 
    n4549 , 
    n4550 , 
    n4551 , 
    n4552 , 
    n4553 , 
    n4554 , 
    n4555 , 
    n4556 , 
    n4557 , 
    n4558 , 
    n4559 , 
    n4560 , 
    n4561 , 
    n4562 , 
    n4563 , 
    n4564 , 
    n4565 , 
    n4566 , 
    n4567 , 
    n4568 , 
    n4569 , 
    n4570 , 
    n4571 , 
    n4572 , 
    n4573 , 
    n4574 , 
    n4575 , 
    n4576 , 
    n4577 , 
    n4578 , 
    n4579 , 
    n4580 , 
    n4581 , 
    n4582 , 
    n4583 , 
    n4584 , 
    n4585 , 
    n4586 , 
    n4587 , 
    n4588 , 
    n4589 , 
    n4590 , 
    n4591 , 
    n4592 , 
    n4593 , 
    n4594 , 
    n4595 , 
    n4596 , 
    n4597 , 
    n4598 , 
    n4599 , 
    n4600 , 
    n4601 , 
    n4602 , 
    n4603 , 
    n4604 , 
    n4605 , 
    n4606 , 
    n4607 , 
    n4608 , 
    n4609 , 
    n4610 , 
    n4611 , 
    n4612 , 
    n4613 , 
    n4614 , 
    n4615 , 
    n4616 , 
    n4617 , 
    n4618 , 
    n4619 , 
    n4620 , 
    n4621 , 
    n4622 , 
    n4623 , 
    n4624 , 
    n4625 , 
    n4626 , 
    n4627 , 
    n4628 , 
    n4629 , 
    n4630 , 
    n4631 , 
    n4632 , 
    n4633 , 
    n4634 , 
    n4635 , 
    n4636 , 
    n4637 , 
    n4638 , 
    n4639 , 
    n4640 , 
    n4641 , 
    n4642 , 
    n4643 , 
    n4644 , 
    n4645 , 
    n4646 , 
    n4647 , 
    n4648 , 
    n4649 , 
    n4650 , 
    n4651 , 
    n4652 , 
    n4653 , 
    n4654 , 
    n4655 , 
    n4656 , 
    n4657 , 
    n4658 , 
    n4659 , 
    n4660 , 
    n4661 , 
    n4662 , 
    n4663 , 
    n4664 , 
    n4665 , 
    n4666 , 
    n4667 , 
    n4668 , 
    n4669 , 
    n4670 , 
    n4671 , 
    n4672 , 
    n4673 , 
    n4674 , 
    n4675 , 
    n4676 , 
    n4677 , 
    n4678 , 
    n4679 , 
    n4680 , 
    n4681 , 
    n4682 , 
    n4683 , 
    n4684 , 
    n4685 , 
    n4686 , 
    n4687 , 
    n4688 , 
    n4689 , 
    n4690 , 
    n4691 , 
    n4692 , 
    n4693 , 
    n4694 , 
    n4695 , 
    n4696 , 
    n4697 , 
    n4698 , 
    n4699 , 
    n4700 , 
    n4701 , 
    n4702 , 
    n4703 , 
    n4704 , 
    n4705 , 
    n4706 , 
    n4707 , 
    n4708 , 
    n4709 , 
    n4710 , 
    n4711 , 
    n4712 , 
    n4713 , 
    n4714 , 
    n4715 , 
    n4716 , 
    n4717 , 
    n4718 , 
    n4719 , 
    n4720 , 
    n4721 , 
    n4722 , 
    n4723 , 
    n4724 , 
    n4725 , 
    n4726 , 
    n4727 , 
    n4728 , 
    n4729 , 
    n4730 , 
    n4731 , 
    n4732 , 
    n4733 , 
    n4734 , 
    n4735 , 
    n4736 , 
    n4737 , 
    n4738 , 
    n4739 , 
    n4740 , 
    n4741 , 
    n4742 , 
    n4743 , 
    n4744 , 
    n4745 , 
    n4746 , 
    n4747 , 
    n4748 , 
    n4749 , 
    n4750 , 
    n4751 , 
    n4752 , 
    n4753 , 
    n4754 , 
    n4755 , 
    n4756 , 
    n4757 , 
    n4758 , 
    n4759 , 
    n4760 , 
    n4761 , 
    n4762 , 
    n4763 , 
    n4764 , 
    n4765 , 
    n4766 , 
    n4767 , 
    n4768 , 
    n4769 , 
    n4770 , 
    n4771 , 
    n4772 , 
    n4773 , 
    n4774 , 
    n4775 , 
    n4776 , 
    n4777 , 
    n4778 , 
    n4779 , 
    n4780 , 
    n4781 , 
    n4782 , 
    n4783 , 
    n4784 , 
    n4785 , 
    n4786 , 
    n4787 , 
    n4788 , 
    n4789 , 
    n4790 , 
    n4791 , 
    n4792 , 
    n4793 , 
    n4794 , 
    n4795 , 
    n4796 , 
    n4797 , 
    n4798 , 
    n4799 , 
    n4800 , 
    n4801 , 
    n4802 , 
    n4803 , 
    n4804 , 
    n4805 , 
    n4806 , 
    n4807 , 
    n4808 , 
    n4809 , 
    n4810 , 
    n4811 , 
    n4812 , 
    n4813 , 
    n4814 , 
    n4815 , 
    n4816 , 
    n4817 , 
    n4818 , 
    n4819 , 
    n4820 , 
    n4821 , 
    n4822 , 
    n4823 , 
    n4824 , 
    n4825 , 
    n4826 , 
    n4827 , 
    n4828 , 
    n4829 , 
    n4830 , 
    n4831 , 
    n4832 , 
    n4833 , 
    n4834 , 
    n4835 , 
    n4836 , 
    n4837 , 
    n4838 , 
    n4839 , 
    n4840 , 
    n4841 , 
    n4842 , 
    n4843 , 
    n4844 , 
    n4845 , 
    n4846 , 
    n4847 , 
    n4848 , 
    n4849 , 
    n4850 , 
    n4851 , 
    n4852 , 
    n4853 , 
    n4854 , 
    n4855 , 
    n4856 , 
    n4857 , 
    n4858 , 
    n4859 , 
    n4860 , 
    n4861 , 
    n4862 , 
    n4863 , 
    n4864 , 
    n4865 , 
    n4866 , 
    n4867 , 
    n4868 , 
    n4869 , 
    n4870 , 
    n4871 , 
    n4872 , 
    n4873 , 
    n4874 , 
    n4875 , 
    n4876 , 
    n4877 , 
    n4878 , 
    n4879 , 
    n4880 , 
    n4881 , 
    n4882 , 
    n4883 , 
    n4884 , 
    n4885 , 
    n4886 , 
    n4887 , 
    n4888 , 
    n4889 , 
    n4890 , 
    n4891 , 
    n4892 , 
    n4893 , 
    n4894 , 
    n4895 , 
    n4896 , 
    n4897 , 
    n4898 , 
    n4899 , 
    n4900 , 
    n4901 , 
    n4902 , 
    n4903 , 
    n4904 , 
    n4905 , 
    n4906 , 
    n4907 , 
    n4908 , 
    n4909 , 
    n4910 , 
    n4911 , 
    n4912 , 
    n4913 , 
    n4914 , 
    n4915 , 
    n4916 , 
    n4917 , 
    n4918 , 
    n4919 , 
    n4920 , 
    n4921 , 
    n4922 , 
    n4923 , 
    n4924 , 
    n4925 , 
    n4926 , 
    n4927 , 
    n4928 , 
    n4929 , 
    n4930 , 
    n4931 , 
    n4932 , 
    n4933 , 
    n4934 , 
    n4935 , 
    n4936 , 
    n4937 , 
    n4938 , 
    n4939 , 
    n4940 , 
    n4941 , 
    n4942 , 
    n4943 , 
    n4944 , 
    n4945 , 
    n4946 , 
    n4947 , 
    n4948 , 
    n4949 , 
    n4950 , 
    n4951 , 
    n4952 , 
    n4953 , 
    n4954 , 
    n4955 , 
    n4956 , 
    n4957 , 
    n4958 , 
    n4959 , 
    n4960 , 
    n4961 , 
    n4962 , 
    n4963 , 
    n4964 , 
    n4965 , 
    n4966 , 
    n4967 , 
    n4968 , 
    n4969 , 
    n4970 , 
    n4971 , 
    n4972 , 
    n4973 , 
    n4974 , 
    n4975 , 
    n4976 , 
    n4977 , 
    n4978 , 
    n4979 , 
    n4980 , 
    n4981 , 
    n4982 , 
    n4983 , 
    n4984 , 
    n4985 , 
    n4986 , 
    n4987 , 
    n4988 , 
    n4989 , 
    n4990 , 
    n4991 , 
    n4992 , 
    n4993 , 
    n4994 , 
    n4995 , 
    n4996 , 
    n4997 , 
    n4998 , 
    n4999 , 
    n5000 , 
    n5001 , 
    n5002 , 
    n5003 , 
    n5004 , 
    n5005 , 
    n5006 , 
    n5007 );
input  n0 , 
    n1 , 
    n2 , 
    n3 , 
    n4 , 
    n5 , 
    n6 , 
    n7 , 
    n8 , 
    n9 , 
    n10 , 
    n11 , 
    n12 , 
    n13 , 
    n14 , 
    n15 , 
    n16 , 
    n17 , 
    n18 , 
    n19 , 
    n20 , 
    n21 , 
    n22 , 
    n23 , 
    n24 , 
    n25 , 
    n26 , 
    n27 , 
    n28 , 
    n29 , 
    n30 , 
    n31 , 
    n32 , 
    n33 , 
    n34 , 
    n35 , 
    n36 , 
    n37 , 
    n38 , 
    n39 , 
    n40 , 
    n41 , 
    n42 , 
    n43 , 
    n44 , 
    n45 , 
    n46 , 
    n47 , 
    n48 , 
    n49 , 
    n50 , 
    n51 , 
    n52 , 
    n53 , 
    n54 , 
    n55 , 
    n56 , 
    n57 , 
    n58 , 
    n59 , 
    n60 , 
    n61 , 
    n62 , 
    n63 , 
    n64 , 
    n65 , 
    n66 , 
    n67 , 
    n68 , 
    n69 , 
    n70 , 
    n71 , 
    n72 , 
    n73 , 
    n74 , 
    n75 , 
    n76 , 
    n77 , 
    n78 , 
    n79 , 
    n80 , 
    n81 , 
    n82 , 
    n83 , 
    n84 , 
    n85 , 
    n86 , 
    n87 , 
    n88 , 
    n89 , 
    n90 , 
    n91 , 
    n92 , 
    n93 , 
    n94 , 
    n95 , 
    n96 , 
    n97 , 
    n98 , 
    n99 , 
    n100 , 
    n101 , 
    n102 , 
    n103 , 
    n104 , 
    n105 , 
    n106 , 
    n107 , 
    n108 , 
    n109 , 
    n110 , 
    n111 , 
    n112 , 
    n113 , 
    n114 , 
    n115 , 
    n116 , 
    n117 , 
    n118 , 
    n119 , 
    n120 , 
    n121 , 
    n122 , 
    n123 , 
    n124 , 
    n125 , 
    n126 , 
    n127 , 
    n128 , 
    n129 , 
    n130 , 
    n131 , 
    n132 , 
    n133 , 
    n134 , 
    n135 , 
    n136 , 
    n137 , 
    n138 , 
    n139 , 
    n140 , 
    n141 , 
    n142 , 
    n143 , 
    n144 , 
    n145 , 
    n146 , 
    n147 , 
    n148 , 
    n149 , 
    n150 , 
    n151 , 
    n152 , 
    n153 , 
    n154 , 
    n155 , 
    n156 , 
    n157 , 
    n158 , 
    n159 , 
    n160 , 
    n161 , 
    n162 , 
    n163 , 
    n164 , 
    n165 , 
    n166 , 
    n167 , 
    n168 , 
    n169 , 
    n170 , 
    n171 , 
    n172 , 
    n173 , 
    n174 , 
    n175 , 
    n176 , 
    n177 , 
    n178 , 
    n179 , 
    n180 , 
    n181 , 
    n182 , 
    n183 , 
    n184 , 
    n185 , 
    n186 , 
    n187 , 
    n188 , 
    n189 , 
    n190 , 
    n191 , 
    n192 , 
    n193 , 
    n194 , 
    n195 , 
    n196 , 
    n197 , 
    n198 , 
    n199 , 
    n200 , 
    n201 , 
    n202 , 
    n203 , 
    n204 , 
    n205 , 
    n206 , 
    n207 , 
    n208 , 
    n209 , 
    n210 , 
    n211 , 
    n212 , 
    n213 , 
    n214 , 
    n215 , 
    n216 , 
    n217 , 
    n218 , 
    n219 , 
    n220 , 
    n221 , 
    n222 , 
    n223 , 
    n224 , 
    n225 , 
    n226 , 
    n227 , 
    n228 , 
    n229 , 
    n230 , 
    n231 , 
    n232 , 
    n233 , 
    n234 , 
    n235 , 
    n236 , 
    n237 , 
    n238 , 
    n239 , 
    n240 , 
    n241 , 
    n242 , 
    n243 , 
    n244 , 
    n245 , 
    n246 , 
    n247 , 
    n248 , 
    n249 , 
    n250 , 
    n251 , 
    n252 , 
    n253 , 
    n254 , 
    n255 , 
    n256 , 
    n257 , 
    n258 , 
    n259 , 
    n260 , 
    n261 , 
    n262 , 
    n263 , 
    n264 , 
    n265 , 
    n266 , 
    n267 , 
    n268 , 
    n269 , 
    n270 , 
    n271 , 
    n272 , 
    n273 , 
    n274 , 
    n275 , 
    n276 , 
    n277 , 
    n278 , 
    n279 , 
    n280 , 
    n281 , 
    n282 , 
    n283 , 
    n284 , 
    n285 , 
    n286 , 
    n287 , 
    n288 , 
    n289 , 
    n290 , 
    n291 , 
    n292 , 
    n293 , 
    n294 , 
    n295 , 
    n296 , 
    n297 , 
    n298 , 
    n299 , 
    n300 , 
    n301 , 
    n302 , 
    n303 , 
    n304 , 
    n305 , 
    n306 , 
    n307 , 
    n308 , 
    n309 , 
    n310 , 
    n311 , 
    n312 , 
    n313 , 
    n314 , 
    n315 , 
    n316 , 
    n317 , 
    n318 , 
    n319 , 
    n320 , 
    n321 , 
    n322 , 
    n323 , 
    n324 , 
    n325 , 
    n326 , 
    n327 , 
    n328 , 
    n329 , 
    n330 , 
    n331 , 
    n332 , 
    n333 , 
    n334 , 
    n335 , 
    n336 , 
    n337 , 
    n338 , 
    n339 , 
    n340 , 
    n341 , 
    n342 , 
    n343 , 
    n344 , 
    n345 , 
    n346 , 
    n347 , 
    n348 , 
    n349 , 
    n350 , 
    n351 , 
    n352 , 
    n353 , 
    n354 , 
    n355 , 
    n356 , 
    n357 , 
    n358 , 
    n359 , 
    n360 , 
    n361 , 
    n362 , 
    n363 , 
    n364 , 
    n365 , 
    n366 , 
    n367 , 
    n368 , 
    n369 , 
    n370 , 
    n371 , 
    n372 , 
    n373 , 
    n374 , 
    n375 , 
    n376 , 
    n377 , 
    n378 , 
    n379 , 
    n380 , 
    n381 , 
    n382 , 
    n383 , 
    n384 , 
    n385 , 
    n386 , 
    n387 , 
    n388 , 
    n389 , 
    n390 , 
    n391 , 
    n392 , 
    n393 , 
    n394 , 
    n395 , 
    n396 , 
    n397 , 
    n398 , 
    n399 , 
    n400 , 
    n401 , 
    n402 , 
    n403 , 
    n404 , 
    n405 , 
    n406 , 
    n407 , 
    n408 , 
    n409 , 
    n410 , 
    n411 , 
    n412 , 
    n413 , 
    n414 , 
    n415 , 
    n416 , 
    n417 , 
    n418 , 
    n419 , 
    n420 , 
    n421 , 
    n422 , 
    n423 , 
    n424 , 
    n425 , 
    n426 , 
    n427 , 
    n428 , 
    n429 , 
    n430 , 
    n431 , 
    n432 , 
    n433 , 
    n434 , 
    n435 , 
    n436 , 
    n437 , 
    n438 , 
    n439 , 
    n440 , 
    n441 , 
    n442 , 
    n443 , 
    n444 , 
    n445 , 
    n446 , 
    n447 , 
    n448 , 
    n449 , 
    n450 , 
    n451 , 
    n452 , 
    n453 , 
    n454 , 
    n455 , 
    n456 , 
    n457 , 
    n458 , 
    n459 , 
    n460 , 
    n461 , 
    n462 , 
    n463 , 
    n464 , 
    n465 , 
    n466 , 
    n467 , 
    n468 , 
    n469 , 
    n470 , 
    n471 , 
    n472 , 
    n473 , 
    n474 , 
    n475 , 
    n476 , 
    n477 , 
    n478 , 
    n479 , 
    n480 , 
    n481 , 
    n482 , 
    n483 , 
    n484 , 
    n485 , 
    n486 , 
    n487 , 
    n488 , 
    n489 , 
    n490 , 
    n491 , 
    n492 , 
    n493 , 
    n494 , 
    n495 , 
    n496 , 
    n497 , 
    n498 , 
    n499 , 
    n500 , 
    n501 , 
    n502 , 
    n503 , 
    n504 , 
    n505 , 
    n506 , 
    n507 , 
    n508 , 
    n509 , 
    n510 , 
    n511 , 
    n512 , 
    n513 , 
    n514 , 
    n515 , 
    n516 , 
    n517 , 
    n518 , 
    n519 , 
    n520 , 
    n521 , 
    n522 , 
    n523 , 
    n524 , 
    n525 , 
    n526 , 
    n527 , 
    n528 , 
    n529 , 
    n530 , 
    n531 , 
    n532 , 
    n533 , 
    n534 , 
    n535 , 
    n536 , 
    n537 , 
    n538 , 
    n539 , 
    n540 , 
    n541 , 
    n542 , 
    n543 , 
    n544 , 
    n545 , 
    n546 , 
    n547 , 
    n548 , 
    n549 , 
    n550 , 
    n551 , 
    n552 , 
    n553 , 
    n554 , 
    n555 , 
    n556 , 
    n557 , 
    n558 , 
    n559 , 
    n560 , 
    n561 , 
    n562 , 
    n563 , 
    n564 , 
    n565 , 
    n566 , 
    n567 , 
    n568 , 
    n569 , 
    n570 , 
    n571 , 
    n572 , 
    n573 , 
    n574 , 
    n575 , 
    n576 , 
    n577 , 
    n578 , 
    n579 , 
    n580 , 
    n581 , 
    n582 , 
    n583 , 
    n584 , 
    n585 , 
    n586 , 
    n587 , 
    n588 , 
    n589 , 
    n590 , 
    n591 , 
    n592 , 
    n593 , 
    n594 , 
    n595 , 
    n596 , 
    n597 , 
    n598 , 
    n599 , 
    n600 , 
    n601 , 
    n602 , 
    n603 , 
    n604 , 
    n605 , 
    n606 , 
    n607 , 
    n608 , 
    n609 , 
    n610 , 
    n611 , 
    n612 , 
    n613 , 
    n614 , 
    n615 , 
    n616 , 
    n617 , 
    n618 , 
    n619 , 
    n620 , 
    n621 , 
    n622 , 
    n623 , 
    n624 , 
    n625 , 
    n626 , 
    n627 , 
    n628 , 
    n629 , 
    n630 , 
    n631 , 
    n632 , 
    n633 , 
    n634 , 
    n635 , 
    n636 , 
    n637 , 
    n638 , 
    n639 , 
    n640 , 
    n641 , 
    n642 , 
    n643 , 
    n644 , 
    n645 , 
    n646 , 
    n647 , 
    n648 , 
    n649 , 
    n650 , 
    n651 , 
    n652 , 
    n653 , 
    n654 , 
    n655 , 
    n656 , 
    n657 , 
    n658 , 
    n659 , 
    n660 , 
    n661 , 
    n662 , 
    n663 , 
    n664 , 
    n665 , 
    n666 , 
    n667 , 
    n668 , 
    n669 , 
    n670 , 
    n671 , 
    n672 , 
    n673 , 
    n674 , 
    n675 , 
    n676 , 
    n677 , 
    n678 , 
    n679 , 
    n680 , 
    n681 , 
    n682 , 
    n683 , 
    n684 , 
    n685 , 
    n686 , 
    n687 , 
    n688 , 
    n689 , 
    n690 , 
    n691 , 
    n692 , 
    n693 , 
    n694 , 
    n695 , 
    n696 , 
    n697 , 
    n698 , 
    n699 , 
    n700 , 
    n701 , 
    n702 , 
    n703 , 
    n704 , 
    n705 , 
    n706 , 
    n707 , 
    n708 , 
    n709 , 
    n710 , 
    n711 , 
    n712 , 
    n713 , 
    n714 , 
    n715 , 
    n716 , 
    n717 , 
    n718 , 
    n719 , 
    n720 , 
    n721 , 
    n722 , 
    n723 , 
    n724 , 
    n725 , 
    n726 , 
    n727 , 
    n728 , 
    n729 , 
    n730 , 
    n731 , 
    n732 , 
    n733 , 
    n734 , 
    n735 , 
    n736 , 
    n737 , 
    n738 , 
    n739 , 
    n740 , 
    n741 , 
    n742 , 
    n743 , 
    n744 , 
    n745 , 
    n746 , 
    n747 , 
    n748 , 
    n749 , 
    n750 , 
    n751 , 
    n752 , 
    n753 , 
    n754 , 
    n755 , 
    n756 , 
    n757 , 
    n758 , 
    n759 , 
    n760 , 
    n761 , 
    n762 , 
    n763 , 
    n764 , 
    n765 , 
    n766 , 
    n767 , 
    n768 , 
    n769 , 
    n770 , 
    n771 , 
    n772 , 
    n773 , 
    n774 , 
    n775 , 
    n776 , 
    n777 , 
    n778 , 
    n779 , 
    n780 , 
    n781 , 
    n782 , 
    n783 , 
    n784 , 
    n785 , 
    n786 , 
    n787 , 
    n788 , 
    n789 , 
    n790 , 
    n791 , 
    n792 , 
    n793 , 
    n794 , 
    n795 , 
    n796 , 
    n797 , 
    n798 , 
    n799 , 
    n800 , 
    n801 , 
    n802 , 
    n803 , 
    n804 , 
    n805 , 
    n806 , 
    n807 , 
    n808 , 
    n809 , 
    n810 , 
    n811 , 
    n812 , 
    n813 , 
    n814 , 
    n815 , 
    n816 , 
    n817 , 
    n818 , 
    n819 , 
    n820 , 
    n821 , 
    n822 , 
    n823 , 
    n824 , 
    n825 , 
    n826 , 
    n827 , 
    n828 , 
    n829 , 
    n830 , 
    n831 , 
    n832 , 
    n833 , 
    n834 , 
    n835 , 
    n836 , 
    n837 , 
    n838 , 
    n839 , 
    n840 , 
    n841 , 
    n842 , 
    n843 , 
    n844 , 
    n845 , 
    n846 , 
    n847 , 
    n848 , 
    n849 , 
    n850 , 
    n851 , 
    n852 , 
    n853 , 
    n854 , 
    n855 , 
    n856 , 
    n857 , 
    n858 , 
    n859 , 
    n860 , 
    n861 , 
    n862 , 
    n863 , 
    n864 , 
    n865 , 
    n866 , 
    n867 , 
    n868 , 
    n869 , 
    n870 , 
    n871 , 
    n872 , 
    n873 , 
    n874 , 
    n875 , 
    n876 , 
    n877 , 
    n878 , 
    n879 , 
    n880 , 
    n881 , 
    n882 , 
    n883 , 
    n884 , 
    n885 , 
    n886 , 
    n887 , 
    n888 , 
    n889 , 
    n890 , 
    n891 , 
    n892 , 
    n893 , 
    n894 , 
    n895 , 
    n896 , 
    n897 , 
    n898 , 
    n899 , 
    n900 , 
    n901 , 
    n902 , 
    n903 , 
    n904 , 
    n905 , 
    n906 , 
    n907 , 
    n908 , 
    n909 , 
    n910 , 
    n911 , 
    n912 , 
    n913 , 
    n914 , 
    n915 , 
    n916 , 
    n917 , 
    n918 , 
    n919 , 
    n920 , 
    n921 , 
    n922 , 
    n923 , 
    n924 , 
    n925 , 
    n926 , 
    n927 , 
    n928 , 
    n929 , 
    n930 , 
    n931 , 
    n932 , 
    n933 , 
    n934 , 
    n935 , 
    n936 , 
    n937 , 
    n938 , 
    n939 , 
    n940 , 
    n941 , 
    n942 , 
    n943 , 
    n944 , 
    n945 , 
    n946 , 
    n947 , 
    n948 , 
    n949 , 
    n950 , 
    n951 , 
    n952 , 
    n953 , 
    n954 , 
    n955 , 
    n956 , 
    n957 , 
    n958 , 
    n959 , 
    n960 , 
    n961 , 
    n962 , 
    n963 , 
    n964 , 
    n965 , 
    n966 , 
    n967 , 
    n968 , 
    n969 , 
    n970 , 
    n971 , 
    n972 , 
    n973 , 
    n974 , 
    n975 , 
    n976 , 
    n977 , 
    n978 , 
    n979 , 
    n980 , 
    n981 , 
    n982 , 
    n983 , 
    n984 , 
    n985 , 
    n986 , 
    n987 , 
    n988 , 
    n989 , 
    n990 , 
    n991 , 
    n992 , 
    n993 , 
    n994 , 
    n995 , 
    n996 , 
    n997 , 
    n998 , 
    n999 , 
    n1000 , 
    n1001 , 
    n1002 , 
    n1003 , 
    n1004 , 
    n1005 , 
    n1006 , 
    n1007 , 
    n1008 , 
    n1009 , 
    n1010 , 
    n1011 , 
    n1012 , 
    n1013 , 
    n1014 , 
    n1015 , 
    n1016 , 
    n1017 , 
    n1018 , 
    n1019 , 
    n1020 , 
    n1021 , 
    n1022 , 
    n1023 , 
    n1024 , 
    n1025 , 
    n1026 , 
    n1027 , 
    n1028 , 
    n1029 , 
    n1030 , 
    n1031 , 
    n1032 , 
    n1033 , 
    n1034 , 
    n1035 , 
    n1036 , 
    n1037 , 
    n1038 , 
    n1039 , 
    n1040 , 
    n1041 , 
    n1042 , 
    n1043 , 
    n1044 , 
    n1045 , 
    n1046 , 
    n1047 , 
    n1048 , 
    n1049 , 
    n1050 , 
    n1051 , 
    n1052 , 
    n1053 , 
    n1054 , 
    n1055 , 
    n1056 , 
    n1057 , 
    n1058 , 
    n1059 , 
    n1060 , 
    n1061 , 
    n1062 , 
    n1063 , 
    n1064 , 
    n1065 , 
    n1066 , 
    n1067 , 
    n1068 , 
    n1069 , 
    n1070 , 
    n1071 , 
    n1072 , 
    n1073 , 
    n1074 , 
    n1075 , 
    n1076 , 
    n1077 , 
    n1078 , 
    n1079 , 
    n1080 , 
    n1081 , 
    n1082 , 
    n1083 , 
    n1084 , 
    n1085 , 
    n1086 , 
    n1087 , 
    n1088 , 
    n1089 , 
    n1090 , 
    n1091 , 
    n1092 , 
    n1093 , 
    n1094 , 
    n1095 , 
    n1096 , 
    n1097 , 
    n1098 , 
    n1099 , 
    n1100 , 
    n1101 , 
    n1102 , 
    n1103 , 
    n1104 , 
    n1105 , 
    n1106 , 
    n1107 , 
    n1108 , 
    n1109 , 
    n1110 , 
    n1111 , 
    n1112 , 
    n1113 , 
    n1114 , 
    n1115 , 
    n1116 , 
    n1117 , 
    n1118 , 
    n1119 , 
    n1120 , 
    n1121 , 
    n1122 , 
    n1123 , 
    n1124 , 
    n1125 , 
    n1126 , 
    n1127 , 
    n1128 , 
    n1129 , 
    n1130 , 
    n1131 , 
    n1132 , 
    n1133 , 
    n1134 , 
    n1135 , 
    n1136 , 
    n1137 , 
    n1138 , 
    n1139 , 
    n1140 , 
    n1141 , 
    n1142 , 
    n1143 , 
    n1144 , 
    n1145 , 
    n1146 , 
    n1147 , 
    n1148 , 
    n1149 , 
    n1150 , 
    n1151 , 
    n1152 , 
    n1153 , 
    n1154 , 
    n1155 , 
    n1156 , 
    n1157 , 
    n1158 , 
    n1159 , 
    n1160 , 
    n1161 , 
    n1162 , 
    n1163 , 
    n1164 , 
    n1165 , 
    n1166 , 
    n1167 , 
    n1168 , 
    n1169 , 
    n1170 , 
    n1171 , 
    n1172 , 
    n1173 , 
    n1174 , 
    n1175 , 
    n1176 , 
    n1177 , 
    n1178 , 
    n1179 , 
    n1180 , 
    n1181 , 
    n1182 , 
    n1183 , 
    n1184 , 
    n1185 , 
    n1186 , 
    n1187 , 
    n1188 , 
    n1189 , 
    n1190 , 
    n1191 , 
    n1192 , 
    n1193 , 
    n1194 , 
    n1195 , 
    n1196 , 
    n1197 , 
    n1198 , 
    n1199 , 
    n1200 , 
    n1201 , 
    n1202 , 
    n1203 , 
    n1204 , 
    n1205 , 
    n1206 , 
    n1207 , 
    n1208 , 
    n1209 , 
    n1210 , 
    n1211 , 
    n1212 , 
    n1213 , 
    n1214 , 
    n1215 , 
    n1216 , 
    n1217 , 
    n1218 , 
    n1219 , 
    n1220 , 
    n1221 , 
    n1222 , 
    n1223 , 
    n1224 , 
    n1225 , 
    n1226 , 
    n1227 , 
    n1228 , 
    n1229 , 
    n1230 , 
    n1231 , 
    n1232 , 
    n1233 , 
    n1234 , 
    n1235 , 
    n1236 , 
    n1237 , 
    n1238 , 
    n1239 , 
    n1240 , 
    n1241 , 
    n1242 , 
    n1243 , 
    n1244 , 
    n1245 , 
    n1246 , 
    n1247 , 
    n1248 , 
    n1249 , 
    n1250 , 
    n1251 , 
    n1252 , 
    n1253 , 
    n1254 , 
    n1255 , 
    n1256 , 
    n1257 , 
    n1258 , 
    n1259 , 
    n1260 , 
    n1261 , 
    n1262 , 
    n1263 , 
    n1264 , 
    n1265 , 
    n1266 , 
    n1267 , 
    n1268 , 
    n1269 , 
    n1270 , 
    n1271 , 
    n1272 , 
    n1273 , 
    n1274 , 
    n1275 , 
    n1276 , 
    n1277 , 
    n1278 , 
    n1279 , 
    n1280 , 
    n1281 , 
    n1282 , 
    n1283 , 
    n1284 , 
    n1285 , 
    n1286 , 
    n1287 , 
    n1288 , 
    n1289 , 
    n1290 , 
    n1291 , 
    n1292 , 
    n1293 , 
    n1294 , 
    n1295 , 
    n1296 , 
    n1297 , 
    n1298 , 
    n1299 , 
    n1300 , 
    n1301 , 
    n1302 , 
    n1303 , 
    n1304 , 
    n1305 , 
    n1306 , 
    n1307 , 
    n1308 , 
    n1309 , 
    n1310 , 
    n1311 , 
    n1312 , 
    n1313 , 
    n1314 , 
    n1315 , 
    n1316 , 
    n1317 , 
    n1318 , 
    n1319 , 
    n1320 , 
    n1321 , 
    n1322 , 
    n1323 , 
    n1324 , 
    n1325 , 
    n1326 , 
    n1327 , 
    n1328 , 
    n1329 , 
    n1330 , 
    n1331 , 
    n1332 , 
    n1333 , 
    n1334 , 
    n1335 , 
    n1336 , 
    n1337 , 
    n1338 , 
    n1339 , 
    n1340 , 
    n1341 , 
    n1342 , 
    n1343 , 
    n1344 , 
    n1345 , 
    n1346 , 
    n1347 , 
    n1348 , 
    n1349 , 
    n1350 , 
    n1351 , 
    n1352 , 
    n1353 , 
    n1354 , 
    n1355 , 
    n1356 , 
    n1357 , 
    n1358 , 
    n1359 , 
    n1360 , 
    n1361 , 
    n1362 , 
    n1363 , 
    n1364 , 
    n1365 , 
    n1366 , 
    n1367 , 
    n1368 , 
    n1369 , 
    n1370 , 
    n1371 , 
    n1372 , 
    n1373 , 
    n1374 , 
    n1375 , 
    n1376 , 
    n1377 , 
    n1378 , 
    n1379 , 
    n1380 , 
    n1381 , 
    n1382 , 
    n1383 , 
    n1384 , 
    n1385 , 
    n1386 , 
    n1387 , 
    n1388 , 
    n1389 , 
    n1390 , 
    n1391 , 
    n1392 , 
    n1393 , 
    n1394 , 
    n1395 , 
    n1396 , 
    n1397 , 
    n1398 , 
    n1399 , 
    n1400 , 
    n1401 , 
    n1402 , 
    n1403 , 
    n1404 , 
    n1405 , 
    n1406 , 
    n1407 , 
    n1408 , 
    n1409 , 
    n1410 , 
    n1411 , 
    n1412 , 
    n1413 , 
    n1414 , 
    n1415 , 
    n1416 , 
    n1417 , 
    n1418 , 
    n1419 , 
    n1420 , 
    n1421 , 
    n1422 , 
    n1423 , 
    n1424 , 
    n1425 , 
    n1426 , 
    n1427 , 
    n1428 , 
    n1429 , 
    n1430 , 
    n1431 , 
    n1432 , 
    n1433 , 
    n1434 , 
    n1435 , 
    n1436 , 
    n1437 , 
    n1438 , 
    n1439 , 
    n1440 , 
    n1441 , 
    n1442 , 
    n1443 , 
    n1444 , 
    n1445 , 
    n1446 , 
    n1447 , 
    n1448 , 
    n1449 , 
    n1450 , 
    n1451 , 
    n1452 , 
    n1453 , 
    n1454 , 
    n1455 , 
    n1456 , 
    n1457 , 
    n1458 , 
    n1459 , 
    n1460 , 
    n1461 , 
    n1462 , 
    n1463 , 
    n1464 , 
    n1465 , 
    n1466 , 
    n1467 , 
    n1468 , 
    n1469 , 
    n1470 , 
    n1471 , 
    n1472 , 
    n1473 , 
    n1474 , 
    n1475 , 
    n1476 , 
    n1477 , 
    n1478 , 
    n1479 , 
    n1480 , 
    n1481 , 
    n1482 , 
    n1483 , 
    n1484 , 
    n1485 , 
    n1486 , 
    n1487 , 
    n1488 , 
    n1489 , 
    n1490 , 
    n1491 , 
    n1492 , 
    n1493 , 
    n1494 , 
    n1495 , 
    n1496 , 
    n1497 , 
    n1498 , 
    n1499 , 
    n1500 , 
    n1501 , 
    n1502 , 
    n1503 , 
    n1504 , 
    n1505 , 
    n1506 , 
    n1507 , 
    n1508 , 
    n1509 , 
    n1510 , 
    n1511 , 
    n1512 , 
    n1513 , 
    n1514 , 
    n1515 , 
    n1516 , 
    n1517 , 
    n1518 , 
    n1519 , 
    n1520 , 
    n1521 , 
    n1522 , 
    n1523 , 
    n1524 , 
    n1525 , 
    n1526 , 
    n1527 , 
    n1528 , 
    n1529 , 
    n1530 , 
    n1531 , 
    n1532 , 
    n1533 , 
    n1534 , 
    n1535 , 
    n1536 , 
    n1537 , 
    n1538 , 
    n1539 , 
    n1540 , 
    n1541 , 
    n1542 , 
    n1543 , 
    n1544 , 
    n1545 , 
    n1546 , 
    n1547 , 
    n1548 , 
    n1549 , 
    n1550 , 
    n1551 , 
    n1552 , 
    n1553 , 
    n1554 , 
    n1555 , 
    n1556 , 
    n1557 , 
    n1558 , 
    n1559 , 
    n1560 , 
    n1561 , 
    n1562 , 
    n1563 , 
    n1564 , 
    n1565 , 
    n1566 , 
    n1567 , 
    n1568 , 
    n1569 , 
    n1570 , 
    n1571 , 
    n1572 , 
    n1573 , 
    n1574 , 
    n1575 , 
    n1576 , 
    n1577 , 
    n1578 , 
    n1579 , 
    n1580 , 
    n1581 , 
    n1582 , 
    n1583 , 
    n1584 , 
    n1585 , 
    n1586 , 
    n1587 , 
    n1588 , 
    n1589 , 
    n1590 , 
    n1591 , 
    n1592 , 
    n1593 , 
    n1594 , 
    n1595 , 
    n1596 , 
    n1597 , 
    n1598 , 
    n1599 , 
    n1600 , 
    n1601 , 
    n1602 , 
    n1603 , 
    n1604 , 
    n1605 , 
    n1606 , 
    n1607 , 
    n1608 , 
    n1609 , 
    n1610 , 
    n1611 , 
    n1612 , 
    n1613 , 
    n1614 , 
    n1615 , 
    n1616 , 
    n1617 , 
    n1618 , 
    n1619 , 
    n1620 , 
    n1621 , 
    n1622 , 
    n1623 , 
    n1624 , 
    n1625 , 
    n1626 , 
    n1627 , 
    n1628 , 
    n1629 , 
    n1630 , 
    n1631 , 
    n1632 , 
    n1633 , 
    n1634 , 
    n1635 , 
    n1636 , 
    n1637 , 
    n1638 , 
    n1639 , 
    n1640 , 
    n1641 , 
    n1642 , 
    n1643 , 
    n1644 , 
    n1645 , 
    n1646 , 
    n1647 , 
    n1648 , 
    n1649 , 
    n1650 , 
    n1651 , 
    n1652 , 
    n1653 , 
    n1654 , 
    n1655 , 
    n1656 , 
    n1657 , 
    n1658 , 
    n1659 , 
    n1660 , 
    n1661 , 
    n1662 , 
    n1663 , 
    n1664 , 
    n1665 , 
    n1666 , 
    n1667 , 
    n1668 , 
    n1669 , 
    n1670 , 
    n1671 , 
    n1672 , 
    n1673 , 
    n1674 , 
    n1675 , 
    n1676 , 
    n1677 , 
    n1678 , 
    n1679 , 
    n1680 , 
    n1681 , 
    n1682 , 
    n1683 , 
    n1684 , 
    n1685 , 
    n1686 , 
    n1687 , 
    n1688 , 
    n1689 , 
    n1690 , 
    n1691 , 
    n1692 , 
    n1693 , 
    n1694 , 
    n1695 , 
    n1696 , 
    n1697 , 
    n1698 , 
    n1699 , 
    n1700 , 
    n1701 , 
    n1702 , 
    n1703 , 
    n1704 , 
    n1705 , 
    n1706 , 
    n1707 , 
    n1708 , 
    n1709 , 
    n1710 , 
    n1711 , 
    n1712 , 
    n1713 , 
    n1714 , 
    n1715 , 
    n1716 , 
    n1717 , 
    n1718 , 
    n1719 , 
    n1720 , 
    n1721 , 
    n1722 , 
    n1723 , 
    n1724 , 
    n1725 , 
    n1726 , 
    n1727 , 
    n1728 , 
    n1729 , 
    n1730 , 
    n1731 , 
    n1732 , 
    n1733 , 
    n1734 , 
    n1735 , 
    n1736 , 
    n1737 , 
    n1738 , 
    n1739 , 
    n1740 , 
    n1741 , 
    n1742 , 
    n1743 , 
    n1744 , 
    n1745 , 
    n1746 , 
    n1747 , 
    n1748 , 
    n1749 , 
    n1750 , 
    n1751 , 
    n1752 , 
    n1753 , 
    n1754 , 
    n1755 , 
    n1756 , 
    n1757 , 
    n1758 , 
    n1759 , 
    n1760 , 
    n1761 , 
    n1762 , 
    n1763 , 
    n1764 , 
    n1765 , 
    n1766 , 
    n1767 , 
    n1768 , 
    n1769 , 
    n1770 , 
    n1771 , 
    n1772 , 
    n1773 , 
    n1774 , 
    n1775 , 
    n1776 , 
    n1777 , 
    n1778 , 
    n1779 , 
    n1780 , 
    n1781 , 
    n1782 , 
    n1783 , 
    n1784 , 
    n1785 , 
    n1786 , 
    n1787 , 
    n1788 , 
    n1789 , 
    n1790 , 
    n1791 , 
    n1792 , 
    n1793 , 
    n1794 , 
    n1795 , 
    n1796 , 
    n1797 , 
    n1798 , 
    n1799 , 
    n1800 , 
    n1801 , 
    n1802 , 
    n1803 , 
    n1804 , 
    n1805 , 
    n1806 , 
    n1807 , 
    n1808 , 
    n1809 , 
    n1810 , 
    n1811 , 
    n1812 , 
    n1813 , 
    n1814 , 
    n1815 , 
    n1816 , 
    n1817 , 
    n1818 , 
    n1819 , 
    n1820 , 
    n1821 , 
    n1822 , 
    n1823 , 
    n1824 , 
    n1825 , 
    n1826 , 
    n1827 , 
    n1828 , 
    n1829 , 
    n1830 , 
    n1831 , 
    n1832 , 
    n1833 , 
    n1834 , 
    n1835 , 
    n1836 , 
    n1837 , 
    n1838 , 
    n1839 , 
    n1840 , 
    n1841 , 
    n1842 , 
    n1843 , 
    n1844 , 
    n1845 , 
    n1846 , 
    n1847 , 
    n1848 , 
    n1849 , 
    n1850 , 
    n1851 , 
    n1852 , 
    n1853 , 
    n1854 , 
    n1855 , 
    n1856 , 
    n1857 , 
    n1858 , 
    n1859 , 
    n1860 , 
    n1861 , 
    n1862 , 
    n1863 , 
    n1864 , 
    n1865 , 
    n1866 , 
    n1867 , 
    n1868 , 
    n1869 , 
    n1870 , 
    n1871 , 
    n1872 , 
    n1873 , 
    n1874 , 
    n1875 , 
    n1876 , 
    n1877 , 
    n1878 , 
    n1879 , 
    n1880 , 
    n1881 , 
    n1882 , 
    n1883 , 
    n1884 , 
    n1885 , 
    n1886 , 
    n1887 , 
    n1888 , 
    n1889 , 
    n1890 , 
    n1891 , 
    n1892 , 
    n1893 , 
    n1894 , 
    n1895 , 
    n1896 , 
    n1897 , 
    n1898 , 
    n1899 , 
    n1900 , 
    n1901 , 
    n1902 , 
    n1903 , 
    n1904 , 
    n1905 , 
    n1906 , 
    n1907 , 
    n1908 , 
    n1909 , 
    n1910 , 
    n1911 , 
    n1912 , 
    n1913 , 
    n1914 , 
    n1915 , 
    n1916 , 
    n1917 , 
    n1918 , 
    n1919 , 
    n1920 , 
    n1921 , 
    n1922 , 
    n1923 , 
    n1924 , 
    n1925 , 
    n1926 , 
    n1927 , 
    n1928 , 
    n1929 , 
    n1930 , 
    n1931 , 
    n1932 , 
    n1933 , 
    n1934 , 
    n1935 , 
    n1936 , 
    n1937 , 
    n1938 , 
    n1939 , 
    n1940 , 
    n1941 , 
    n1942 , 
    n1943 , 
    n1944 , 
    n1945 , 
    n1946 , 
    n1947 , 
    n1948 , 
    n1949 , 
    n1950 , 
    n1951 , 
    n1952 , 
    n1953 , 
    n1954 , 
    n1955 , 
    n1956 , 
    n1957 , 
    n1958 , 
    n1959 , 
    n1960 , 
    n1961 , 
    n1962 , 
    n1963 , 
    n1964 , 
    n1965 , 
    n1966 , 
    n1967 , 
    n1968 , 
    n1969 , 
    n1970 , 
    n1971 , 
    n1972 , 
    n1973 , 
    n1974 , 
    n1975 , 
    n1976 , 
    n1977 , 
    n1978 , 
    n1979 , 
    n1980 , 
    n1981 , 
    n1982 , 
    n1983 , 
    n1984 , 
    n1985 , 
    n1986 , 
    n1987 , 
    n1988 , 
    n1989 , 
    n1990 , 
    n1991 , 
    n1992 , 
    n1993 , 
    n1994 , 
    n1995 , 
    n1996 , 
    n1997 , 
    n1998 , 
    n1999 , 
    n2000 , 
    n2001 , 
    n2002 , 
    n2003 , 
    n2004 , 
    n2005 , 
    n2006 , 
    n2007 , 
    n2008 , 
    n2009 , 
    n2010 , 
    n2011 , 
    n2012 , 
    n2013 , 
    n2014 , 
    n2015 , 
    n2016 , 
    n2017 , 
    n2018 , 
    n2019 , 
    n2020 , 
    n2021 , 
    n2022 , 
    n2023 , 
    n2024 , 
    n2025 , 
    n2026 , 
    n2027 , 
    n2028 , 
    n2029 , 
    n2030 , 
    n2031 , 
    n2032 , 
    n2033 , 
    n2034 , 
    n2035 , 
    n2036 , 
    n2037 , 
    n2038 , 
    n2039 , 
    n2040 , 
    n2041 , 
    n2042 , 
    n2043 , 
    n2044 , 
    n2045 , 
    n2046 , 
    n2047 , 
    n2048 , 
    n2049 , 
    n2050 , 
    n2051 , 
    n2052 , 
    n2053 , 
    n2054 , 
    n2055 , 
    n2056 , 
    n2057 , 
    n2058 , 
    n2059 , 
    n2060 , 
    n2061 , 
    n2062 , 
    n2063 , 
    n2064 , 
    n2065 , 
    n2066 , 
    n2067 , 
    n2068 , 
    n2069 , 
    n2070 , 
    n2071 , 
    n2072 , 
    n2073 , 
    n2074 , 
    n2075 , 
    n2076 , 
    n2077 , 
    n2078 , 
    n2079 , 
    n2080 , 
    n2081 , 
    n2082 , 
    n2083 , 
    n2084 , 
    n2085 , 
    n2086 , 
    n2087 , 
    n2088 , 
    n2089 , 
    n2090 , 
    n2091 , 
    n2092 , 
    n2093 , 
    n2094 , 
    n2095 , 
    n2096 , 
    n2097 , 
    n2098 , 
    n2099 , 
    n2100 , 
    n2101 , 
    n2102 , 
    n2103 , 
    n2104 , 
    n2105 , 
    n2106 , 
    n2107 , 
    n2108 , 
    n2109 , 
    n2110 , 
    n2111 , 
    n2112 , 
    n2113 , 
    n2114 , 
    n2115 , 
    n2116 , 
    n2117 , 
    n2118 , 
    n2119 , 
    n2120 , 
    n2121 , 
    n2122 , 
    n2123 , 
    n2124 , 
    n2125 , 
    n2126 , 
    n2127 , 
    n2128 , 
    n2129 , 
    n2130 , 
    n2131 , 
    n2132 , 
    n2133 , 
    n2134 , 
    n2135 , 
    n2136 , 
    n2137 , 
    n2138 , 
    n2139 , 
    n2140 , 
    n2141 , 
    n2142 , 
    n2143 , 
    n2144 , 
    n2145 , 
    n2146 , 
    n2147 , 
    n2148 , 
    n2149 , 
    n2150 , 
    n2151 , 
    n2152 , 
    n2153 , 
    n2154 , 
    n2155 , 
    n2156 , 
    n2157 , 
    n2158 , 
    n2159 , 
    n2160 , 
    n2161 , 
    n2162 , 
    n2163 , 
    n2164 , 
    n2165 , 
    n2166 , 
    n2167 , 
    n2168 , 
    n2169 , 
    n2170 , 
    n2171 , 
    n2172 , 
    n2173 , 
    n2174 , 
    n2175 , 
    n2176 , 
    n2177 , 
    n2178 , 
    n2179 , 
    n2180 , 
    n2181 , 
    n2182 , 
    n2183 , 
    n2184 , 
    n2185 , 
    n2186 , 
    n2187 , 
    n2188 , 
    n2189 , 
    n2190 , 
    n2191 , 
    n2192 , 
    n2193 , 
    n2194 , 
    n2195 , 
    n2196 , 
    n2197 , 
    n2198 , 
    n2199 , 
    n2200 , 
    n2201 , 
    n2202 , 
    n2203 , 
    n2204 , 
    n2205 , 
    n2206 , 
    n2207 , 
    n2208 , 
    n2209 , 
    n2210 , 
    n2211 , 
    n2212 , 
    n2213 , 
    n2214 , 
    n2215 , 
    n2216 , 
    n2217 , 
    n2218 , 
    n2219 , 
    n2220 , 
    n2221 , 
    n2222 , 
    n2223 , 
    n2224 , 
    n2225 , 
    n2226 , 
    n2227 , 
    n2228 , 
    n2229 , 
    n2230 , 
    n2231 , 
    n2232 , 
    n2233 , 
    n2234 , 
    n2235 , 
    n2236 , 
    n2237 , 
    n2238 , 
    n2239 , 
    n2240 , 
    n2241 , 
    n2242 , 
    n2243 , 
    n2244 , 
    n2245 , 
    n2246 , 
    n2247 , 
    n2248 , 
    n2249 , 
    n2250 , 
    n2251 , 
    n2252 , 
    n2253 , 
    n2254 , 
    n2255 , 
    n2256 , 
    n2257 , 
    n2258 , 
    n2259 , 
    n2260 , 
    n2261 , 
    n2262 , 
    n2263 , 
    n2264 , 
    n2265 , 
    n2266 , 
    n2267 , 
    n2268 , 
    n2269 , 
    n2270 , 
    n2271 , 
    n2272 , 
    n2273 , 
    n2274 , 
    n2275 , 
    n2276 , 
    n2277 , 
    n2278 , 
    n2279 , 
    n2280 , 
    n2281 ;
output n2282 , 
    n2283 , 
    n2284 , 
    n2285 , 
    n2286 , 
    n2287 , 
    n2288 , 
    n2289 , 
    n2290 , 
    n2291 , 
    n2292 , 
    n2293 , 
    n2294 , 
    n2295 , 
    n2296 , 
    n2297 , 
    n2298 , 
    n2299 , 
    n2300 , 
    n2301 , 
    n2302 , 
    n2303 , 
    n2304 , 
    n2305 , 
    n2306 , 
    n2307 , 
    n2308 , 
    n2309 , 
    n2310 , 
    n2311 , 
    n2312 , 
    n2313 , 
    n2314 , 
    n2315 , 
    n2316 , 
    n2317 , 
    n2318 , 
    n2319 , 
    n2320 , 
    n2321 , 
    n2322 , 
    n2323 , 
    n2324 , 
    n2325 , 
    n2326 , 
    n2327 , 
    n2328 , 
    n2329 , 
    n2330 , 
    n2331 , 
    n2332 , 
    n2333 , 
    n2334 , 
    n2335 , 
    n2336 , 
    n2337 , 
    n2338 , 
    n2339 , 
    n2340 , 
    n2341 , 
    n2342 , 
    n2343 , 
    n2344 , 
    n2345 , 
    n2346 , 
    n2347 , 
    n2348 , 
    n2349 , 
    n2350 , 
    n2351 , 
    n2352 , 
    n2353 , 
    n2354 , 
    n2355 , 
    n2356 , 
    n2357 , 
    n2358 , 
    n2359 , 
    n2360 , 
    n2361 , 
    n2362 , 
    n2363 , 
    n2364 , 
    n2365 , 
    n2366 , 
    n2367 , 
    n2368 , 
    n2369 , 
    n2370 , 
    n2371 , 
    n2372 , 
    n2373 , 
    n2374 , 
    n2375 , 
    n2376 , 
    n2377 , 
    n2378 , 
    n2379 , 
    n2380 , 
    n2381 , 
    n2382 , 
    n2383 , 
    n2384 , 
    n2385 , 
    n2386 , 
    n2387 , 
    n2388 , 
    n2389 , 
    n2390 , 
    n2391 , 
    n2392 , 
    n2393 , 
    n2394 , 
    n2395 , 
    n2396 , 
    n2397 , 
    n2398 , 
    n2399 , 
    n2400 , 
    n2401 , 
    n2402 , 
    n2403 , 
    n2404 , 
    n2405 , 
    n2406 , 
    n2407 , 
    n2408 , 
    n2409 , 
    n2410 , 
    n2411 , 
    n2412 , 
    n2413 , 
    n2414 , 
    n2415 , 
    n2416 , 
    n2417 , 
    n2418 , 
    n2419 , 
    n2420 , 
    n2421 , 
    n2422 , 
    n2423 , 
    n2424 , 
    n2425 , 
    n2426 , 
    n2427 , 
    n2428 , 
    n2429 , 
    n2430 , 
    n2431 , 
    n2432 , 
    n2433 , 
    n2434 , 
    n2435 , 
    n2436 , 
    n2437 , 
    n2438 , 
    n2439 , 
    n2440 , 
    n2441 , 
    n2442 , 
    n2443 , 
    n2444 , 
    n2445 , 
    n2446 , 
    n2447 , 
    n2448 , 
    n2449 , 
    n2450 , 
    n2451 , 
    n2452 , 
    n2453 , 
    n2454 , 
    n2455 , 
    n2456 , 
    n2457 , 
    n2458 , 
    n2459 , 
    n2460 , 
    n2461 , 
    n2462 , 
    n2463 , 
    n2464 , 
    n2465 , 
    n2466 , 
    n2467 , 
    n2468 , 
    n2469 , 
    n2470 , 
    n2471 , 
    n2472 , 
    n2473 , 
    n2474 , 
    n2475 , 
    n2476 , 
    n2477 , 
    n2478 , 
    n2479 , 
    n2480 , 
    n2481 , 
    n2482 , 
    n2483 , 
    n2484 , 
    n2485 , 
    n2486 , 
    n2487 , 
    n2488 , 
    n2489 , 
    n2490 , 
    n2491 , 
    n2492 , 
    n2493 , 
    n2494 , 
    n2495 , 
    n2496 , 
    n2497 , 
    n2498 , 
    n2499 , 
    n2500 , 
    n2501 , 
    n2502 , 
    n2503 , 
    n2504 , 
    n2505 , 
    n2506 , 
    n2507 , 
    n2508 , 
    n2509 , 
    n2510 , 
    n2511 , 
    n2512 , 
    n2513 , 
    n2514 , 
    n2515 , 
    n2516 , 
    n2517 , 
    n2518 , 
    n2519 , 
    n2520 , 
    n2521 , 
    n2522 , 
    n2523 , 
    n2524 , 
    n2525 , 
    n2526 , 
    n2527 , 
    n2528 , 
    n2529 , 
    n2530 , 
    n2531 , 
    n2532 , 
    n2533 , 
    n2534 , 
    n2535 , 
    n2536 , 
    n2537 , 
    n2538 , 
    n2539 , 
    n2540 , 
    n2541 , 
    n2542 , 
    n2543 , 
    n2544 , 
    n2545 , 
    n2546 , 
    n2547 , 
    n2548 , 
    n2549 , 
    n2550 , 
    n2551 , 
    n2552 , 
    n2553 , 
    n2554 , 
    n2555 , 
    n2556 , 
    n2557 , 
    n2558 , 
    n2559 , 
    n2560 , 
    n2561 , 
    n2562 , 
    n2563 , 
    n2564 , 
    n2565 , 
    n2566 , 
    n2567 , 
    n2568 , 
    n2569 , 
    n2570 , 
    n2571 , 
    n2572 , 
    n2573 , 
    n2574 , 
    n2575 , 
    n2576 , 
    n2577 , 
    n2578 , 
    n2579 , 
    n2580 , 
    n2581 , 
    n2582 , 
    n2583 , 
    n2584 , 
    n2585 , 
    n2586 , 
    n2587 , 
    n2588 , 
    n2589 , 
    n2590 , 
    n2591 , 
    n2592 , 
    n2593 , 
    n2594 , 
    n2595 , 
    n2596 , 
    n2597 , 
    n2598 , 
    n2599 , 
    n2600 , 
    n2601 , 
    n2602 , 
    n2603 , 
    n2604 , 
    n2605 , 
    n2606 , 
    n2607 , 
    n2608 , 
    n2609 , 
    n2610 , 
    n2611 , 
    n2612 , 
    n2613 , 
    n2614 , 
    n2615 , 
    n2616 , 
    n2617 , 
    n2618 , 
    n2619 , 
    n2620 , 
    n2621 , 
    n2622 , 
    n2623 , 
    n2624 , 
    n2625 , 
    n2626 , 
    n2627 , 
    n2628 , 
    n2629 , 
    n2630 , 
    n2631 , 
    n2632 , 
    n2633 , 
    n2634 , 
    n2635 , 
    n2636 , 
    n2637 , 
    n2638 , 
    n2639 , 
    n2640 , 
    n2641 , 
    n2642 , 
    n2643 , 
    n2644 , 
    n2645 , 
    n2646 , 
    n2647 , 
    n2648 , 
    n2649 , 
    n2650 , 
    n2651 , 
    n2652 , 
    n2653 , 
    n2654 , 
    n2655 , 
    n2656 , 
    n2657 , 
    n2658 , 
    n2659 , 
    n2660 , 
    n2661 , 
    n2662 , 
    n2663 , 
    n2664 , 
    n2665 , 
    n2666 , 
    n2667 , 
    n2668 , 
    n2669 , 
    n2670 , 
    n2671 , 
    n2672 , 
    n2673 , 
    n2674 , 
    n2675 , 
    n2676 , 
    n2677 , 
    n2678 , 
    n2679 , 
    n2680 , 
    n2681 , 
    n2682 , 
    n2683 , 
    n2684 , 
    n2685 , 
    n2686 , 
    n2687 , 
    n2688 , 
    n2689 , 
    n2690 , 
    n2691 , 
    n2692 , 
    n2693 , 
    n2694 , 
    n2695 , 
    n2696 , 
    n2697 , 
    n2698 , 
    n2699 , 
    n2700 , 
    n2701 , 
    n2702 , 
    n2703 , 
    n2704 , 
    n2705 , 
    n2706 , 
    n2707 , 
    n2708 , 
    n2709 , 
    n2710 , 
    n2711 , 
    n2712 , 
    n2713 , 
    n2714 , 
    n2715 , 
    n2716 , 
    n2717 , 
    n2718 , 
    n2719 , 
    n2720 , 
    n2721 , 
    n2722 , 
    n2723 , 
    n2724 , 
    n2725 , 
    n2726 , 
    n2727 , 
    n2728 , 
    n2729 , 
    n2730 , 
    n2731 , 
    n2732 , 
    n2733 , 
    n2734 , 
    n2735 , 
    n2736 , 
    n2737 , 
    n2738 , 
    n2739 , 
    n2740 , 
    n2741 , 
    n2742 , 
    n2743 , 
    n2744 , 
    n2745 , 
    n2746 , 
    n2747 , 
    n2748 , 
    n2749 , 
    n2750 , 
    n2751 , 
    n2752 , 
    n2753 , 
    n2754 , 
    n2755 , 
    n2756 , 
    n2757 , 
    n2758 , 
    n2759 , 
    n2760 , 
    n2761 , 
    n2762 , 
    n2763 , 
    n2764 , 
    n2765 , 
    n2766 , 
    n2767 , 
    n2768 , 
    n2769 , 
    n2770 , 
    n2771 , 
    n2772 , 
    n2773 , 
    n2774 , 
    n2775 , 
    n2776 , 
    n2777 , 
    n2778 , 
    n2779 , 
    n2780 , 
    n2781 , 
    n2782 , 
    n2783 , 
    n2784 , 
    n2785 , 
    n2786 , 
    n2787 , 
    n2788 , 
    n2789 , 
    n2790 , 
    n2791 , 
    n2792 , 
    n2793 , 
    n2794 , 
    n2795 , 
    n2796 , 
    n2797 , 
    n2798 , 
    n2799 , 
    n2800 , 
    n2801 , 
    n2802 , 
    n2803 , 
    n2804 , 
    n2805 , 
    n2806 , 
    n2807 , 
    n2808 , 
    n2809 , 
    n2810 , 
    n2811 , 
    n2812 , 
    n2813 , 
    n2814 , 
    n2815 , 
    n2816 , 
    n2817 , 
    n2818 , 
    n2819 , 
    n2820 , 
    n2821 , 
    n2822 , 
    n2823 , 
    n2824 , 
    n2825 , 
    n2826 , 
    n2827 , 
    n2828 , 
    n2829 , 
    n2830 , 
    n2831 , 
    n2832 , 
    n2833 , 
    n2834 , 
    n2835 , 
    n2836 , 
    n2837 , 
    n2838 , 
    n2839 , 
    n2840 , 
    n2841 , 
    n2842 , 
    n2843 , 
    n2844 , 
    n2845 , 
    n2846 , 
    n2847 , 
    n2848 , 
    n2849 , 
    n2850 , 
    n2851 , 
    n2852 , 
    n2853 , 
    n2854 , 
    n2855 , 
    n2856 , 
    n2857 , 
    n2858 , 
    n2859 , 
    n2860 , 
    n2861 , 
    n2862 , 
    n2863 , 
    n2864 , 
    n2865 , 
    n2866 , 
    n2867 , 
    n2868 , 
    n2869 , 
    n2870 , 
    n2871 , 
    n2872 , 
    n2873 , 
    n2874 , 
    n2875 , 
    n2876 , 
    n2877 , 
    n2878 , 
    n2879 , 
    n2880 , 
    n2881 , 
    n2882 , 
    n2883 , 
    n2884 , 
    n2885 , 
    n2886 , 
    n2887 , 
    n2888 , 
    n2889 , 
    n2890 , 
    n2891 , 
    n2892 , 
    n2893 , 
    n2894 , 
    n2895 , 
    n2896 , 
    n2897 , 
    n2898 , 
    n2899 , 
    n2900 , 
    n2901 , 
    n2902 , 
    n2903 , 
    n2904 , 
    n2905 , 
    n2906 , 
    n2907 , 
    n2908 , 
    n2909 , 
    n2910 , 
    n2911 , 
    n2912 , 
    n2913 , 
    n2914 , 
    n2915 , 
    n2916 , 
    n2917 , 
    n2918 , 
    n2919 , 
    n2920 , 
    n2921 , 
    n2922 , 
    n2923 , 
    n2924 , 
    n2925 , 
    n2926 , 
    n2927 , 
    n2928 , 
    n2929 , 
    n2930 , 
    n2931 , 
    n2932 , 
    n2933 , 
    n2934 , 
    n2935 , 
    n2936 , 
    n2937 , 
    n2938 , 
    n2939 , 
    n2940 , 
    n2941 , 
    n2942 , 
    n2943 , 
    n2944 , 
    n2945 , 
    n2946 , 
    n2947 , 
    n2948 , 
    n2949 , 
    n2950 , 
    n2951 , 
    n2952 , 
    n2953 , 
    n2954 , 
    n2955 , 
    n2956 , 
    n2957 , 
    n2958 , 
    n2959 , 
    n2960 , 
    n2961 , 
    n2962 , 
    n2963 , 
    n2964 , 
    n2965 , 
    n2966 , 
    n2967 , 
    n2968 , 
    n2969 , 
    n2970 , 
    n2971 , 
    n2972 , 
    n2973 , 
    n2974 , 
    n2975 , 
    n2976 , 
    n2977 , 
    n2978 , 
    n2979 , 
    n2980 , 
    n2981 , 
    n2982 , 
    n2983 , 
    n2984 , 
    n2985 , 
    n2986 , 
    n2987 , 
    n2988 , 
    n2989 , 
    n2990 , 
    n2991 , 
    n2992 , 
    n2993 , 
    n2994 , 
    n2995 , 
    n2996 , 
    n2997 , 
    n2998 , 
    n2999 , 
    n3000 , 
    n3001 , 
    n3002 , 
    n3003 , 
    n3004 , 
    n3005 , 
    n3006 , 
    n3007 , 
    n3008 , 
    n3009 , 
    n3010 , 
    n3011 , 
    n3012 , 
    n3013 , 
    n3014 , 
    n3015 , 
    n3016 , 
    n3017 , 
    n3018 , 
    n3019 , 
    n3020 , 
    n3021 , 
    n3022 , 
    n3023 , 
    n3024 , 
    n3025 , 
    n3026 , 
    n3027 , 
    n3028 , 
    n3029 , 
    n3030 , 
    n3031 , 
    n3032 , 
    n3033 , 
    n3034 , 
    n3035 , 
    n3036 , 
    n3037 , 
    n3038 , 
    n3039 , 
    n3040 , 
    n3041 , 
    n3042 , 
    n3043 , 
    n3044 , 
    n3045 , 
    n3046 , 
    n3047 , 
    n3048 , 
    n3049 , 
    n3050 , 
    n3051 , 
    n3052 , 
    n3053 , 
    n3054 , 
    n3055 , 
    n3056 , 
    n3057 , 
    n3058 , 
    n3059 , 
    n3060 , 
    n3061 , 
    n3062 , 
    n3063 , 
    n3064 , 
    n3065 , 
    n3066 , 
    n3067 , 
    n3068 , 
    n3069 , 
    n3070 , 
    n3071 , 
    n3072 , 
    n3073 , 
    n3074 , 
    n3075 , 
    n3076 , 
    n3077 , 
    n3078 , 
    n3079 , 
    n3080 , 
    n3081 , 
    n3082 , 
    n3083 , 
    n3084 , 
    n3085 , 
    n3086 , 
    n3087 , 
    n3088 , 
    n3089 , 
    n3090 , 
    n3091 , 
    n3092 , 
    n3093 , 
    n3094 , 
    n3095 , 
    n3096 , 
    n3097 , 
    n3098 , 
    n3099 , 
    n3100 , 
    n3101 , 
    n3102 , 
    n3103 , 
    n3104 , 
    n3105 , 
    n3106 , 
    n3107 , 
    n3108 , 
    n3109 , 
    n3110 , 
    n3111 , 
    n3112 , 
    n3113 , 
    n3114 , 
    n3115 , 
    n3116 , 
    n3117 , 
    n3118 , 
    n3119 , 
    n3120 , 
    n3121 , 
    n3122 , 
    n3123 , 
    n3124 , 
    n3125 , 
    n3126 , 
    n3127 , 
    n3128 , 
    n3129 , 
    n3130 , 
    n3131 , 
    n3132 , 
    n3133 , 
    n3134 , 
    n3135 , 
    n3136 , 
    n3137 , 
    n3138 , 
    n3139 , 
    n3140 , 
    n3141 , 
    n3142 , 
    n3143 , 
    n3144 , 
    n3145 , 
    n3146 , 
    n3147 , 
    n3148 , 
    n3149 , 
    n3150 , 
    n3151 , 
    n3152 , 
    n3153 , 
    n3154 , 
    n3155 , 
    n3156 , 
    n3157 , 
    n3158 , 
    n3159 , 
    n3160 , 
    n3161 , 
    n3162 , 
    n3163 , 
    n3164 , 
    n3165 , 
    n3166 , 
    n3167 , 
    n3168 , 
    n3169 , 
    n3170 , 
    n3171 , 
    n3172 , 
    n3173 , 
    n3174 , 
    n3175 , 
    n3176 , 
    n3177 , 
    n3178 , 
    n3179 , 
    n3180 , 
    n3181 , 
    n3182 , 
    n3183 , 
    n3184 , 
    n3185 , 
    n3186 , 
    n3187 , 
    n3188 , 
    n3189 , 
    n3190 , 
    n3191 , 
    n3192 , 
    n3193 , 
    n3194 , 
    n3195 , 
    n3196 , 
    n3197 , 
    n3198 , 
    n3199 , 
    n3200 , 
    n3201 , 
    n3202 , 
    n3203 , 
    n3204 , 
    n3205 , 
    n3206 , 
    n3207 , 
    n3208 , 
    n3209 , 
    n3210 , 
    n3211 , 
    n3212 , 
    n3213 , 
    n3214 , 
    n3215 , 
    n3216 , 
    n3217 , 
    n3218 , 
    n3219 , 
    n3220 , 
    n3221 , 
    n3222 , 
    n3223 , 
    n3224 , 
    n3225 , 
    n3226 , 
    n3227 , 
    n3228 , 
    n3229 , 
    n3230 , 
    n3231 , 
    n3232 , 
    n3233 , 
    n3234 , 
    n3235 , 
    n3236 , 
    n3237 , 
    n3238 , 
    n3239 , 
    n3240 , 
    n3241 , 
    n3242 , 
    n3243 , 
    n3244 , 
    n3245 , 
    n3246 , 
    n3247 , 
    n3248 , 
    n3249 , 
    n3250 , 
    n3251 , 
    n3252 , 
    n3253 , 
    n3254 , 
    n3255 , 
    n3256 , 
    n3257 , 
    n3258 , 
    n3259 , 
    n3260 , 
    n3261 , 
    n3262 , 
    n3263 , 
    n3264 , 
    n3265 , 
    n3266 , 
    n3267 , 
    n3268 , 
    n3269 , 
    n3270 , 
    n3271 , 
    n3272 , 
    n3273 , 
    n3274 , 
    n3275 , 
    n3276 , 
    n3277 , 
    n3278 , 
    n3279 , 
    n3280 , 
    n3281 , 
    n3282 , 
    n3283 , 
    n3284 , 
    n3285 , 
    n3286 , 
    n3287 , 
    n3288 , 
    n3289 , 
    n3290 , 
    n3291 , 
    n3292 , 
    n3293 , 
    n3294 , 
    n3295 , 
    n3296 , 
    n3297 , 
    n3298 , 
    n3299 , 
    n3300 , 
    n3301 , 
    n3302 , 
    n3303 , 
    n3304 , 
    n3305 , 
    n3306 , 
    n3307 , 
    n3308 , 
    n3309 , 
    n3310 , 
    n3311 , 
    n3312 , 
    n3313 , 
    n3314 , 
    n3315 , 
    n3316 , 
    n3317 , 
    n3318 , 
    n3319 , 
    n3320 , 
    n3321 , 
    n3322 , 
    n3323 , 
    n3324 , 
    n3325 , 
    n3326 , 
    n3327 , 
    n3328 , 
    n3329 , 
    n3330 , 
    n3331 , 
    n3332 , 
    n3333 , 
    n3334 , 
    n3335 , 
    n3336 , 
    n3337 , 
    n3338 , 
    n3339 , 
    n3340 , 
    n3341 , 
    n3342 , 
    n3343 , 
    n3344 , 
    n3345 , 
    n3346 , 
    n3347 , 
    n3348 , 
    n3349 , 
    n3350 , 
    n3351 , 
    n3352 , 
    n3353 , 
    n3354 , 
    n3355 , 
    n3356 , 
    n3357 , 
    n3358 , 
    n3359 , 
    n3360 , 
    n3361 , 
    n3362 , 
    n3363 , 
    n3364 , 
    n3365 , 
    n3366 , 
    n3367 , 
    n3368 , 
    n3369 , 
    n3370 , 
    n3371 , 
    n3372 , 
    n3373 , 
    n3374 , 
    n3375 , 
    n3376 , 
    n3377 , 
    n3378 , 
    n3379 , 
    n3380 , 
    n3381 , 
    n3382 , 
    n3383 , 
    n3384 , 
    n3385 , 
    n3386 , 
    n3387 , 
    n3388 , 
    n3389 , 
    n3390 , 
    n3391 , 
    n3392 , 
    n3393 , 
    n3394 , 
    n3395 , 
    n3396 , 
    n3397 , 
    n3398 , 
    n3399 , 
    n3400 , 
    n3401 , 
    n3402 , 
    n3403 , 
    n3404 , 
    n3405 , 
    n3406 , 
    n3407 , 
    n3408 , 
    n3409 , 
    n3410 , 
    n3411 , 
    n3412 , 
    n3413 , 
    n3414 , 
    n3415 , 
    n3416 , 
    n3417 , 
    n3418 , 
    n3419 , 
    n3420 , 
    n3421 , 
    n3422 , 
    n3423 , 
    n3424 , 
    n3425 , 
    n3426 , 
    n3427 , 
    n3428 , 
    n3429 , 
    n3430 , 
    n3431 , 
    n3432 , 
    n3433 , 
    n3434 , 
    n3435 , 
    n3436 , 
    n3437 , 
    n3438 , 
    n3439 , 
    n3440 , 
    n3441 , 
    n3442 , 
    n3443 , 
    n3444 , 
    n3445 , 
    n3446 , 
    n3447 , 
    n3448 , 
    n3449 , 
    n3450 , 
    n3451 , 
    n3452 , 
    n3453 , 
    n3454 , 
    n3455 , 
    n3456 , 
    n3457 , 
    n3458 , 
    n3459 , 
    n3460 , 
    n3461 , 
    n3462 , 
    n3463 , 
    n3464 , 
    n3465 , 
    n3466 , 
    n3467 , 
    n3468 , 
    n3469 , 
    n3470 , 
    n3471 , 
    n3472 , 
    n3473 , 
    n3474 , 
    n3475 , 
    n3476 , 
    n3477 , 
    n3478 , 
    n3479 , 
    n3480 , 
    n3481 , 
    n3482 , 
    n3483 , 
    n3484 , 
    n3485 , 
    n3486 , 
    n3487 , 
    n3488 , 
    n3489 , 
    n3490 , 
    n3491 , 
    n3492 , 
    n3493 , 
    n3494 , 
    n3495 , 
    n3496 , 
    n3497 , 
    n3498 , 
    n3499 , 
    n3500 , 
    n3501 , 
    n3502 , 
    n3503 , 
    n3504 , 
    n3505 , 
    n3506 , 
    n3507 , 
    n3508 , 
    n3509 , 
    n3510 , 
    n3511 , 
    n3512 , 
    n3513 , 
    n3514 , 
    n3515 , 
    n3516 , 
    n3517 , 
    n3518 , 
    n3519 , 
    n3520 , 
    n3521 , 
    n3522 , 
    n3523 , 
    n3524 , 
    n3525 , 
    n3526 , 
    n3527 , 
    n3528 , 
    n3529 , 
    n3530 , 
    n3531 , 
    n3532 , 
    n3533 , 
    n3534 , 
    n3535 , 
    n3536 , 
    n3537 , 
    n3538 , 
    n3539 , 
    n3540 , 
    n3541 , 
    n3542 , 
    n3543 , 
    n3544 , 
    n3545 , 
    n3546 , 
    n3547 , 
    n3548 , 
    n3549 , 
    n3550 , 
    n3551 , 
    n3552 , 
    n3553 , 
    n3554 , 
    n3555 , 
    n3556 , 
    n3557 , 
    n3558 , 
    n3559 , 
    n3560 , 
    n3561 , 
    n3562 , 
    n3563 , 
    n3564 , 
    n3565 , 
    n3566 , 
    n3567 , 
    n3568 , 
    n3569 , 
    n3570 , 
    n3571 , 
    n3572 , 
    n3573 , 
    n3574 , 
    n3575 , 
    n3576 , 
    n3577 , 
    n3578 , 
    n3579 , 
    n3580 , 
    n3581 , 
    n3582 , 
    n3583 , 
    n3584 , 
    n3585 , 
    n3586 , 
    n3587 , 
    n3588 , 
    n3589 , 
    n3590 , 
    n3591 , 
    n3592 , 
    n3593 , 
    n3594 , 
    n3595 , 
    n3596 , 
    n3597 , 
    n3598 , 
    n3599 , 
    n3600 , 
    n3601 , 
    n3602 , 
    n3603 , 
    n3604 , 
    n3605 , 
    n3606 , 
    n3607 , 
    n3608 , 
    n3609 , 
    n3610 , 
    n3611 , 
    n3612 , 
    n3613 , 
    n3614 , 
    n3615 , 
    n3616 , 
    n3617 , 
    n3618 , 
    n3619 , 
    n3620 , 
    n3621 , 
    n3622 , 
    n3623 , 
    n3624 , 
    n3625 , 
    n3626 , 
    n3627 , 
    n3628 , 
    n3629 , 
    n3630 , 
    n3631 , 
    n3632 , 
    n3633 , 
    n3634 , 
    n3635 , 
    n3636 , 
    n3637 , 
    n3638 , 
    n3639 , 
    n3640 , 
    n3641 , 
    n3642 , 
    n3643 , 
    n3644 , 
    n3645 , 
    n3646 , 
    n3647 , 
    n3648 , 
    n3649 , 
    n3650 , 
    n3651 , 
    n3652 , 
    n3653 , 
    n3654 , 
    n3655 , 
    n3656 , 
    n3657 , 
    n3658 , 
    n3659 , 
    n3660 , 
    n3661 , 
    n3662 , 
    n3663 , 
    n3664 , 
    n3665 , 
    n3666 , 
    n3667 , 
    n3668 , 
    n3669 , 
    n3670 , 
    n3671 , 
    n3672 , 
    n3673 , 
    n3674 , 
    n3675 , 
    n3676 , 
    n3677 , 
    n3678 , 
    n3679 , 
    n3680 , 
    n3681 , 
    n3682 , 
    n3683 , 
    n3684 , 
    n3685 , 
    n3686 , 
    n3687 , 
    n3688 , 
    n3689 , 
    n3690 , 
    n3691 , 
    n3692 , 
    n3693 , 
    n3694 , 
    n3695 , 
    n3696 , 
    n3697 , 
    n3698 , 
    n3699 , 
    n3700 , 
    n3701 , 
    n3702 , 
    n3703 , 
    n3704 , 
    n3705 , 
    n3706 , 
    n3707 , 
    n3708 , 
    n3709 , 
    n3710 , 
    n3711 , 
    n3712 , 
    n3713 , 
    n3714 , 
    n3715 , 
    n3716 , 
    n3717 , 
    n3718 , 
    n3719 , 
    n3720 , 
    n3721 , 
    n3722 , 
    n3723 , 
    n3724 , 
    n3725 , 
    n3726 , 
    n3727 , 
    n3728 , 
    n3729 , 
    n3730 , 
    n3731 , 
    n3732 , 
    n3733 , 
    n3734 , 
    n3735 , 
    n3736 , 
    n3737 , 
    n3738 , 
    n3739 , 
    n3740 , 
    n3741 , 
    n3742 , 
    n3743 , 
    n3744 , 
    n3745 , 
    n3746 , 
    n3747 , 
    n3748 , 
    n3749 , 
    n3750 , 
    n3751 , 
    n3752 , 
    n3753 , 
    n3754 , 
    n3755 , 
    n3756 , 
    n3757 , 
    n3758 , 
    n3759 , 
    n3760 , 
    n3761 , 
    n3762 , 
    n3763 , 
    n3764 , 
    n3765 , 
    n3766 , 
    n3767 , 
    n3768 , 
    n3769 , 
    n3770 , 
    n3771 , 
    n3772 , 
    n3773 , 
    n3774 , 
    n3775 , 
    n3776 , 
    n3777 , 
    n3778 , 
    n3779 , 
    n3780 , 
    n3781 , 
    n3782 , 
    n3783 , 
    n3784 , 
    n3785 , 
    n3786 , 
    n3787 , 
    n3788 , 
    n3789 , 
    n3790 , 
    n3791 , 
    n3792 , 
    n3793 , 
    n3794 , 
    n3795 , 
    n3796 , 
    n3797 , 
    n3798 , 
    n3799 , 
    n3800 , 
    n3801 , 
    n3802 , 
    n3803 , 
    n3804 , 
    n3805 , 
    n3806 , 
    n3807 , 
    n3808 , 
    n3809 , 
    n3810 , 
    n3811 , 
    n3812 , 
    n3813 , 
    n3814 , 
    n3815 , 
    n3816 , 
    n3817 , 
    n3818 , 
    n3819 , 
    n3820 , 
    n3821 , 
    n3822 , 
    n3823 , 
    n3824 , 
    n3825 , 
    n3826 , 
    n3827 , 
    n3828 , 
    n3829 , 
    n3830 , 
    n3831 , 
    n3832 , 
    n3833 , 
    n3834 , 
    n3835 , 
    n3836 , 
    n3837 , 
    n3838 , 
    n3839 , 
    n3840 , 
    n3841 , 
    n3842 , 
    n3843 , 
    n3844 , 
    n3845 , 
    n3846 , 
    n3847 , 
    n3848 , 
    n3849 , 
    n3850 , 
    n3851 , 
    n3852 , 
    n3853 , 
    n3854 , 
    n3855 , 
    n3856 , 
    n3857 , 
    n3858 , 
    n3859 , 
    n3860 , 
    n3861 , 
    n3862 , 
    n3863 , 
    n3864 , 
    n3865 , 
    n3866 , 
    n3867 , 
    n3868 , 
    n3869 , 
    n3870 , 
    n3871 , 
    n3872 , 
    n3873 , 
    n3874 , 
    n3875 , 
    n3876 , 
    n3877 , 
    n3878 , 
    n3879 , 
    n3880 , 
    n3881 , 
    n3882 , 
    n3883 , 
    n3884 , 
    n3885 , 
    n3886 , 
    n3887 , 
    n3888 , 
    n3889 , 
    n3890 , 
    n3891 , 
    n3892 , 
    n3893 , 
    n3894 , 
    n3895 , 
    n3896 , 
    n3897 , 
    n3898 , 
    n3899 , 
    n3900 , 
    n3901 , 
    n3902 , 
    n3903 , 
    n3904 , 
    n3905 , 
    n3906 , 
    n3907 , 
    n3908 , 
    n3909 , 
    n3910 , 
    n3911 , 
    n3912 , 
    n3913 , 
    n3914 , 
    n3915 , 
    n3916 , 
    n3917 , 
    n3918 , 
    n3919 , 
    n3920 , 
    n3921 , 
    n3922 , 
    n3923 , 
    n3924 , 
    n3925 , 
    n3926 , 
    n3927 , 
    n3928 , 
    n3929 , 
    n3930 , 
    n3931 , 
    n3932 , 
    n3933 , 
    n3934 , 
    n3935 , 
    n3936 , 
    n3937 , 
    n3938 , 
    n3939 , 
    n3940 , 
    n3941 , 
    n3942 , 
    n3943 , 
    n3944 , 
    n3945 , 
    n3946 , 
    n3947 , 
    n3948 , 
    n3949 , 
    n3950 , 
    n3951 , 
    n3952 , 
    n3953 , 
    n3954 , 
    n3955 , 
    n3956 , 
    n3957 , 
    n3958 , 
    n3959 , 
    n3960 , 
    n3961 , 
    n3962 , 
    n3963 , 
    n3964 , 
    n3965 , 
    n3966 , 
    n3967 , 
    n3968 , 
    n3969 , 
    n3970 , 
    n3971 , 
    n3972 , 
    n3973 , 
    n3974 , 
    n3975 , 
    n3976 , 
    n3977 , 
    n3978 , 
    n3979 , 
    n3980 , 
    n3981 , 
    n3982 , 
    n3983 , 
    n3984 , 
    n3985 , 
    n3986 , 
    n3987 , 
    n3988 , 
    n3989 , 
    n3990 , 
    n3991 , 
    n3992 , 
    n3993 , 
    n3994 , 
    n3995 , 
    n3996 , 
    n3997 , 
    n3998 , 
    n3999 , 
    n4000 , 
    n4001 , 
    n4002 , 
    n4003 , 
    n4004 , 
    n4005 , 
    n4006 , 
    n4007 , 
    n4008 , 
    n4009 , 
    n4010 , 
    n4011 , 
    n4012 , 
    n4013 , 
    n4014 , 
    n4015 , 
    n4016 , 
    n4017 , 
    n4018 , 
    n4019 , 
    n4020 , 
    n4021 , 
    n4022 , 
    n4023 , 
    n4024 , 
    n4025 , 
    n4026 , 
    n4027 , 
    n4028 , 
    n4029 , 
    n4030 , 
    n4031 , 
    n4032 , 
    n4033 , 
    n4034 , 
    n4035 , 
    n4036 , 
    n4037 , 
    n4038 , 
    n4039 , 
    n4040 , 
    n4041 , 
    n4042 , 
    n4043 , 
    n4044 , 
    n4045 , 
    n4046 , 
    n4047 , 
    n4048 , 
    n4049 , 
    n4050 , 
    n4051 , 
    n4052 , 
    n4053 , 
    n4054 , 
    n4055 , 
    n4056 , 
    n4057 , 
    n4058 , 
    n4059 , 
    n4060 , 
    n4061 , 
    n4062 , 
    n4063 , 
    n4064 , 
    n4065 , 
    n4066 , 
    n4067 , 
    n4068 , 
    n4069 , 
    n4070 , 
    n4071 , 
    n4072 , 
    n4073 , 
    n4074 , 
    n4075 , 
    n4076 , 
    n4077 , 
    n4078 , 
    n4079 , 
    n4080 , 
    n4081 , 
    n4082 , 
    n4083 , 
    n4084 , 
    n4085 , 
    n4086 , 
    n4087 , 
    n4088 , 
    n4089 , 
    n4090 , 
    n4091 , 
    n4092 , 
    n4093 , 
    n4094 , 
    n4095 , 
    n4096 , 
    n4097 , 
    n4098 , 
    n4099 , 
    n4100 , 
    n4101 , 
    n4102 , 
    n4103 , 
    n4104 , 
    n4105 , 
    n4106 , 
    n4107 , 
    n4108 , 
    n4109 , 
    n4110 , 
    n4111 , 
    n4112 , 
    n4113 , 
    n4114 , 
    n4115 , 
    n4116 , 
    n4117 , 
    n4118 , 
    n4119 , 
    n4120 , 
    n4121 , 
    n4122 , 
    n4123 , 
    n4124 , 
    n4125 , 
    n4126 , 
    n4127 , 
    n4128 , 
    n4129 , 
    n4130 , 
    n4131 , 
    n4132 , 
    n4133 , 
    n4134 , 
    n4135 , 
    n4136 , 
    n4137 , 
    n4138 , 
    n4139 , 
    n4140 , 
    n4141 , 
    n4142 , 
    n4143 , 
    n4144 , 
    n4145 , 
    n4146 , 
    n4147 , 
    n4148 , 
    n4149 , 
    n4150 , 
    n4151 , 
    n4152 , 
    n4153 , 
    n4154 , 
    n4155 , 
    n4156 , 
    n4157 , 
    n4158 , 
    n4159 , 
    n4160 , 
    n4161 , 
    n4162 , 
    n4163 , 
    n4164 , 
    n4165 , 
    n4166 , 
    n4167 , 
    n4168 , 
    n4169 , 
    n4170 , 
    n4171 , 
    n4172 , 
    n4173 , 
    n4174 , 
    n4175 , 
    n4176 , 
    n4177 , 
    n4178 , 
    n4179 , 
    n4180 , 
    n4181 , 
    n4182 , 
    n4183 , 
    n4184 , 
    n4185 , 
    n4186 , 
    n4187 , 
    n4188 , 
    n4189 , 
    n4190 , 
    n4191 , 
    n4192 , 
    n4193 , 
    n4194 , 
    n4195 , 
    n4196 , 
    n4197 , 
    n4198 , 
    n4199 , 
    n4200 , 
    n4201 , 
    n4202 , 
    n4203 , 
    n4204 , 
    n4205 , 
    n4206 , 
    n4207 , 
    n4208 , 
    n4209 , 
    n4210 , 
    n4211 , 
    n4212 , 
    n4213 , 
    n4214 , 
    n4215 , 
    n4216 , 
    n4217 , 
    n4218 , 
    n4219 , 
    n4220 , 
    n4221 , 
    n4222 , 
    n4223 , 
    n4224 , 
    n4225 , 
    n4226 , 
    n4227 , 
    n4228 , 
    n4229 , 
    n4230 , 
    n4231 , 
    n4232 , 
    n4233 , 
    n4234 , 
    n4235 , 
    n4236 , 
    n4237 , 
    n4238 , 
    n4239 , 
    n4240 , 
    n4241 , 
    n4242 , 
    n4243 , 
    n4244 , 
    n4245 , 
    n4246 , 
    n4247 , 
    n4248 , 
    n4249 , 
    n4250 , 
    n4251 , 
    n4252 , 
    n4253 , 
    n4254 , 
    n4255 , 
    n4256 , 
    n4257 , 
    n4258 , 
    n4259 , 
    n4260 , 
    n4261 , 
    n4262 , 
    n4263 , 
    n4264 , 
    n4265 , 
    n4266 , 
    n4267 , 
    n4268 , 
    n4269 , 
    n4270 , 
    n4271 , 
    n4272 , 
    n4273 , 
    n4274 , 
    n4275 , 
    n4276 , 
    n4277 , 
    n4278 , 
    n4279 , 
    n4280 , 
    n4281 , 
    n4282 , 
    n4283 , 
    n4284 , 
    n4285 , 
    n4286 , 
    n4287 , 
    n4288 , 
    n4289 , 
    n4290 , 
    n4291 , 
    n4292 , 
    n4293 , 
    n4294 , 
    n4295 , 
    n4296 , 
    n4297 , 
    n4298 , 
    n4299 , 
    n4300 , 
    n4301 , 
    n4302 , 
    n4303 , 
    n4304 , 
    n4305 , 
    n4306 , 
    n4307 , 
    n4308 , 
    n4309 , 
    n4310 , 
    n4311 , 
    n4312 , 
    n4313 , 
    n4314 , 
    n4315 , 
    n4316 , 
    n4317 , 
    n4318 , 
    n4319 , 
    n4320 , 
    n4321 , 
    n4322 , 
    n4323 , 
    n4324 , 
    n4325 , 
    n4326 , 
    n4327 , 
    n4328 , 
    n4329 , 
    n4330 , 
    n4331 , 
    n4332 , 
    n4333 , 
    n4334 , 
    n4335 , 
    n4336 , 
    n4337 , 
    n4338 , 
    n4339 , 
    n4340 , 
    n4341 , 
    n4342 , 
    n4343 , 
    n4344 , 
    n4345 , 
    n4346 , 
    n4347 , 
    n4348 , 
    n4349 , 
    n4350 , 
    n4351 , 
    n4352 , 
    n4353 , 
    n4354 , 
    n4355 , 
    n4356 , 
    n4357 , 
    n4358 , 
    n4359 , 
    n4360 , 
    n4361 , 
    n4362 , 
    n4363 , 
    n4364 , 
    n4365 , 
    n4366 , 
    n4367 , 
    n4368 , 
    n4369 , 
    n4370 , 
    n4371 , 
    n4372 , 
    n4373 , 
    n4374 , 
    n4375 , 
    n4376 , 
    n4377 , 
    n4378 , 
    n4379 , 
    n4380 , 
    n4381 , 
    n4382 , 
    n4383 , 
    n4384 , 
    n4385 , 
    n4386 , 
    n4387 , 
    n4388 , 
    n4389 , 
    n4390 , 
    n4391 , 
    n4392 , 
    n4393 , 
    n4394 , 
    n4395 , 
    n4396 , 
    n4397 , 
    n4398 , 
    n4399 , 
    n4400 , 
    n4401 , 
    n4402 , 
    n4403 , 
    n4404 , 
    n4405 , 
    n4406 , 
    n4407 , 
    n4408 , 
    n4409 , 
    n4410 , 
    n4411 , 
    n4412 , 
    n4413 , 
    n4414 , 
    n4415 , 
    n4416 , 
    n4417 , 
    n4418 , 
    n4419 , 
    n4420 , 
    n4421 , 
    n4422 , 
    n4423 , 
    n4424 , 
    n4425 , 
    n4426 , 
    n4427 , 
    n4428 , 
    n4429 , 
    n4430 , 
    n4431 , 
    n4432 , 
    n4433 , 
    n4434 , 
    n4435 , 
    n4436 , 
    n4437 , 
    n4438 , 
    n4439 , 
    n4440 , 
    n4441 , 
    n4442 , 
    n4443 , 
    n4444 , 
    n4445 , 
    n4446 , 
    n4447 , 
    n4448 , 
    n4449 , 
    n4450 , 
    n4451 , 
    n4452 , 
    n4453 , 
    n4454 , 
    n4455 , 
    n4456 , 
    n4457 , 
    n4458 , 
    n4459 , 
    n4460 , 
    n4461 , 
    n4462 , 
    n4463 , 
    n4464 , 
    n4465 , 
    n4466 , 
    n4467 , 
    n4468 , 
    n4469 , 
    n4470 , 
    n4471 , 
    n4472 , 
    n4473 , 
    n4474 , 
    n4475 , 
    n4476 , 
    n4477 , 
    n4478 , 
    n4479 , 
    n4480 , 
    n4481 , 
    n4482 , 
    n4483 , 
    n4484 , 
    n4485 , 
    n4486 , 
    n4487 , 
    n4488 , 
    n4489 , 
    n4490 , 
    n4491 , 
    n4492 , 
    n4493 , 
    n4494 , 
    n4495 , 
    n4496 , 
    n4497 , 
    n4498 , 
    n4499 , 
    n4500 , 
    n4501 , 
    n4502 , 
    n4503 , 
    n4504 , 
    n4505 , 
    n4506 , 
    n4507 , 
    n4508 , 
    n4509 , 
    n4510 , 
    n4511 , 
    n4512 , 
    n4513 , 
    n4514 , 
    n4515 , 
    n4516 , 
    n4517 , 
    n4518 , 
    n4519 , 
    n4520 , 
    n4521 , 
    n4522 , 
    n4523 , 
    n4524 , 
    n4525 , 
    n4526 , 
    n4527 , 
    n4528 , 
    n4529 , 
    n4530 , 
    n4531 , 
    n4532 , 
    n4533 , 
    n4534 , 
    n4535 , 
    n4536 , 
    n4537 , 
    n4538 , 
    n4539 , 
    n4540 , 
    n4541 , 
    n4542 , 
    n4543 , 
    n4544 , 
    n4545 , 
    n4546 , 
    n4547 , 
    n4548 , 
    n4549 , 
    n4550 , 
    n4551 , 
    n4552 , 
    n4553 , 
    n4554 , 
    n4555 , 
    n4556 , 
    n4557 , 
    n4558 , 
    n4559 , 
    n4560 , 
    n4561 , 
    n4562 , 
    n4563 , 
    n4564 , 
    n4565 , 
    n4566 , 
    n4567 , 
    n4568 , 
    n4569 , 
    n4570 , 
    n4571 , 
    n4572 , 
    n4573 , 
    n4574 , 
    n4575 , 
    n4576 , 
    n4577 , 
    n4578 , 
    n4579 , 
    n4580 , 
    n4581 , 
    n4582 , 
    n4583 , 
    n4584 , 
    n4585 , 
    n4586 , 
    n4587 , 
    n4588 , 
    n4589 , 
    n4590 , 
    n4591 , 
    n4592 , 
    n4593 , 
    n4594 , 
    n4595 , 
    n4596 , 
    n4597 , 
    n4598 , 
    n4599 , 
    n4600 , 
    n4601 , 
    n4602 , 
    n4603 , 
    n4604 , 
    n4605 , 
    n4606 , 
    n4607 , 
    n4608 , 
    n4609 , 
    n4610 , 
    n4611 , 
    n4612 , 
    n4613 , 
    n4614 , 
    n4615 , 
    n4616 , 
    n4617 , 
    n4618 , 
    n4619 , 
    n4620 , 
    n4621 , 
    n4622 , 
    n4623 , 
    n4624 , 
    n4625 , 
    n4626 , 
    n4627 , 
    n4628 , 
    n4629 , 
    n4630 , 
    n4631 , 
    n4632 , 
    n4633 , 
    n4634 , 
    n4635 , 
    n4636 , 
    n4637 , 
    n4638 , 
    n4639 , 
    n4640 , 
    n4641 , 
    n4642 , 
    n4643 , 
    n4644 , 
    n4645 , 
    n4646 , 
    n4647 , 
    n4648 , 
    n4649 , 
    n4650 , 
    n4651 , 
    n4652 , 
    n4653 , 
    n4654 , 
    n4655 , 
    n4656 , 
    n4657 , 
    n4658 , 
    n4659 , 
    n4660 , 
    n4661 , 
    n4662 , 
    n4663 , 
    n4664 , 
    n4665 , 
    n4666 , 
    n4667 , 
    n4668 , 
    n4669 , 
    n4670 , 
    n4671 , 
    n4672 , 
    n4673 , 
    n4674 , 
    n4675 , 
    n4676 , 
    n4677 , 
    n4678 , 
    n4679 , 
    n4680 , 
    n4681 , 
    n4682 , 
    n4683 , 
    n4684 , 
    n4685 , 
    n4686 , 
    n4687 , 
    n4688 , 
    n4689 , 
    n4690 , 
    n4691 , 
    n4692 , 
    n4693 , 
    n4694 , 
    n4695 , 
    n4696 , 
    n4697 , 
    n4698 , 
    n4699 , 
    n4700 , 
    n4701 , 
    n4702 , 
    n4703 , 
    n4704 , 
    n4705 , 
    n4706 , 
    n4707 , 
    n4708 , 
    n4709 , 
    n4710 , 
    n4711 , 
    n4712 , 
    n4713 , 
    n4714 , 
    n4715 , 
    n4716 , 
    n4717 , 
    n4718 , 
    n4719 , 
    n4720 , 
    n4721 , 
    n4722 , 
    n4723 , 
    n4724 , 
    n4725 , 
    n4726 , 
    n4727 , 
    n4728 , 
    n4729 , 
    n4730 , 
    n4731 , 
    n4732 , 
    n4733 , 
    n4734 , 
    n4735 , 
    n4736 , 
    n4737 , 
    n4738 , 
    n4739 , 
    n4740 , 
    n4741 , 
    n4742 , 
    n4743 , 
    n4744 , 
    n4745 , 
    n4746 , 
    n4747 , 
    n4748 , 
    n4749 , 
    n4750 , 
    n4751 , 
    n4752 , 
    n4753 , 
    n4754 , 
    n4755 , 
    n4756 , 
    n4757 , 
    n4758 , 
    n4759 , 
    n4760 , 
    n4761 , 
    n4762 , 
    n4763 , 
    n4764 , 
    n4765 , 
    n4766 , 
    n4767 , 
    n4768 , 
    n4769 , 
    n4770 , 
    n4771 , 
    n4772 , 
    n4773 , 
    n4774 , 
    n4775 , 
    n4776 , 
    n4777 , 
    n4778 , 
    n4779 , 
    n4780 , 
    n4781 , 
    n4782 , 
    n4783 , 
    n4784 , 
    n4785 , 
    n4786 , 
    n4787 , 
    n4788 , 
    n4789 , 
    n4790 , 
    n4791 , 
    n4792 , 
    n4793 , 
    n4794 , 
    n4795 , 
    n4796 , 
    n4797 , 
    n4798 , 
    n4799 , 
    n4800 , 
    n4801 , 
    n4802 , 
    n4803 , 
    n4804 , 
    n4805 , 
    n4806 , 
    n4807 , 
    n4808 , 
    n4809 , 
    n4810 , 
    n4811 , 
    n4812 , 
    n4813 , 
    n4814 , 
    n4815 , 
    n4816 , 
    n4817 , 
    n4818 , 
    n4819 , 
    n4820 , 
    n4821 , 
    n4822 , 
    n4823 , 
    n4824 , 
    n4825 , 
    n4826 , 
    n4827 , 
    n4828 , 
    n4829 , 
    n4830 , 
    n4831 , 
    n4832 , 
    n4833 , 
    n4834 , 
    n4835 , 
    n4836 , 
    n4837 , 
    n4838 , 
    n4839 , 
    n4840 , 
    n4841 , 
    n4842 , 
    n4843 , 
    n4844 , 
    n4845 , 
    n4846 , 
    n4847 , 
    n4848 , 
    n4849 , 
    n4850 , 
    n4851 , 
    n4852 , 
    n4853 , 
    n4854 , 
    n4855 , 
    n4856 , 
    n4857 , 
    n4858 , 
    n4859 , 
    n4860 , 
    n4861 , 
    n4862 , 
    n4863 , 
    n4864 , 
    n4865 , 
    n4866 , 
    n4867 , 
    n4868 , 
    n4869 , 
    n4870 , 
    n4871 , 
    n4872 , 
    n4873 , 
    n4874 , 
    n4875 , 
    n4876 , 
    n4877 , 
    n4878 , 
    n4879 , 
    n4880 , 
    n4881 , 
    n4882 , 
    n4883 , 
    n4884 , 
    n4885 , 
    n4886 , 
    n4887 , 
    n4888 , 
    n4889 , 
    n4890 , 
    n4891 , 
    n4892 , 
    n4893 , 
    n4894 , 
    n4895 , 
    n4896 , 
    n4897 , 
    n4898 , 
    n4899 , 
    n4900 , 
    n4901 , 
    n4902 , 
    n4903 , 
    n4904 , 
    n4905 , 
    n4906 , 
    n4907 , 
    n4908 , 
    n4909 , 
    n4910 , 
    n4911 , 
    n4912 , 
    n4913 , 
    n4914 , 
    n4915 , 
    n4916 , 
    n4917 , 
    n4918 , 
    n4919 , 
    n4920 , 
    n4921 , 
    n4922 , 
    n4923 , 
    n4924 , 
    n4925 , 
    n4926 , 
    n4927 , 
    n4928 , 
    n4929 , 
    n4930 , 
    n4931 , 
    n4932 , 
    n4933 , 
    n4934 , 
    n4935 , 
    n4936 , 
    n4937 , 
    n4938 , 
    n4939 , 
    n4940 , 
    n4941 , 
    n4942 , 
    n4943 , 
    n4944 , 
    n4945 , 
    n4946 , 
    n4947 , 
    n4948 , 
    n4949 , 
    n4950 , 
    n4951 , 
    n4952 , 
    n4953 , 
    n4954 , 
    n4955 , 
    n4956 , 
    n4957 , 
    n4958 , 
    n4959 , 
    n4960 , 
    n4961 , 
    n4962 , 
    n4963 , 
    n4964 , 
    n4965 , 
    n4966 , 
    n4967 , 
    n4968 , 
    n4969 , 
    n4970 , 
    n4971 , 
    n4972 , 
    n4973 , 
    n4974 , 
    n4975 , 
    n4976 , 
    n4977 , 
    n4978 , 
    n4979 , 
    n4980 , 
    n4981 , 
    n4982 , 
    n4983 , 
    n4984 , 
    n4985 , 
    n4986 , 
    n4987 , 
    n4988 , 
    n4989 , 
    n4990 , 
    n4991 , 
    n4992 , 
    n4993 , 
    n4994 , 
    n4995 , 
    n4996 , 
    n4997 , 
    n4998 , 
    n4999 , 
    n5000 , 
    n5001 , 
    n5002 , 
    n5003 , 
    n5004 , 
    n5005 , 
    n5006 , 
    n5007 ;

wire 
    RI19a22f70_2797 , 
    RI1754a798_67 , 
    RI19ad04a8_2209 , 
    RI19a23e70_2789 , 
    RI1754c610_2 , 
    RI19a23510_2794 , 
    RI19a859b8_2755 , 
    RI17534808_603 , 
    RI173f4d68_1562 , 
    RI173ac078_1917 , 
    RI17516358_697 , 
    RI1753aa78_586 , 
    RI19aad828_2471 , 
    RI17491398_1028 , 
    RI19ac0a40_2326 , 
    RI1751df18_673 , 
    RI173c95b0_1774 , 
    RI17340030_2129 , 
    RI174125e8_1418 , 
    RI19a8ffa8_2683 , 
    RI17465bf8_1240 , 
    RI19ac0680_2328 , 
    RI174ae8d0_885 , 
    RI1733be90_2149 , 
    RI173c9268_1775 , 
    RI173ff808_1510 , 
    RI173b67d0_1866 , 
    RI1752e610_622 , 
    RI1749baf0_977 , 
    RI19ab9a38_2383 , 
    RI173d4068_1722 , 
    RI1738b378_2077 , 
    RI1744bb40_1367 , 
    RI19a9c5f0_2595 , 
    RI17470350_1189 , 
    RI19acb828_2243 , 
    RI174b9460_834 , 
    RI173dd410_1677 , 
    RI173cee48_1747 , 
    RI17345580_2103 , 
    RI17446938_1392 , 
    RI19a8c498_2709 , 
    RI1746b148_1214 , 
    RI19abd890_2354 , 
    RI174b3e20_859 , 
    RI173ec398_1604 , 
    RI173a36a8_1959 , 
    RI1747e900_1119 , 
    RI19acf1d0_2217 , 
    RI17510160_716 , 
    RI19aa05b0_2566 , 
    RI17488680_1071 , 
    RI173895f0_2086 , 
    RI1740b9a0_1451 , 
    RI173c2cb0_1806 , 
    RI17339730_2161 , 
    RI174a7fd0_917 , 
    RI19ab3138_2431 , 
    RI19a95048_2647 , 
    RI1752a308_635 , 
    RI173ee468_1594 , 
    RI173a5778_1949 , 
    RI17493120_1019 , 
    RI19a9f548_2574 , 
    RI1748a750_1061 , 
    RI19ace168_2224 , 
    RI17513a18_705 , 
    RI173cd750_1754 , 
    RI173441d0_2109 , 
    RI17445588_1398 , 
    RI19a8dfc8_2697 , 
    RI17469d98_1220 , 
    RI19abeda8_2342 , 
    RI174b2a70_865 , 
    RI173bee58_1825 , 
    RI173f9250_1541 , 
    RI173b0560_1896 , 
    RI17389938_2085 , 
    RI19aadb70_2470 , 
    RI17524b60_652 , 
    RI19aab938_2485 , 
    RI17495880_1007 , 
    RI173e1268_1658 , 
    RI17398578_2013 , 
    RI17459088_1302 , 
    RI19a93d88_2655 , 
    RI1747d898_1124 , 
    RI19ac40a0_2299 , 
    RI174ce388_769 , 
    RI19a9e030_2584 , 
    RI1748be48_1054 , 
    RI173feae8_1514 , 
    RI173b5ab0_1870 , 
    RI173c0208_1819 , 
    RI19aa7c48_2511 , 
    RI1749add0_981 , 
    RI19a88e38_2732 , 
    RI1752d170_626 , 
    RI19a9bfd8_2598 , 
    RI1746f978_1192 , 
    RI1733b800_2151 , 
    RI173c4d80_1796 , 
    RI1740da70_1441 , 
    RI19ac21b0_2313 , 
    RI174aa0a0_907 , 
    RI19a91e98_2669 , 
    RI174613c8_1262 , 
    RI17399298_2009 , 
    RI173e1f88_1654 , 
    RI17459da8_1298 , 
    RI19a86c00_2747 , 
    RI174cf828_765 , 
    RI19aa5740_2526 , 
    RI1747e5b8_1120 , 
    RI173fda80_1519 , 
    RI173bc068_1839 , 
    RI17404d58_1484 , 
    RI17332ae8_2194 , 
    RI19ab5d48_2410 , 
    RI174a1040_951 , 
    RI173ad0e0_1912 , 
    RI173e7820_1627 , 
    RI1739e7e8_1983 , 
    RI1745f2f8_1272 , 
    RI19aa1d20_2554 , 
    RI17483b08_1094 , 
    RI19a82d30_2774 , 
    RI17508ac8_739 , 
    RI19a876c8_2742 , 
    RI174d1208_760 , 
    RI173d46f8_1720 , 
    RI1738ba08_2075 , 
    RI1744c1d0_1365 , 
    RI19a9ca28_2593 , 
    RI174709e0_1187 , 
    RI19acbc60_2241 , 
    RI174b9eb0_832 , 
    RI173a8f40_1932 , 
    RI173f1c30_1577 , 
    RI174b75e8_842 , 
    RI19ab0870_2450 , 
    RI1748df18_1044 , 
    RI19ac1d78_2315 , 
    RI175191c0_688 , 
    RI19abe6a0_2346 , 
    RI174b1d50_869 , 
    RI173db9d0_1685 , 
    RI17392ce0_2040 , 
    RI174534a8_1330 , 
    RI19ac7700_2274 , 
    RI174c5850_796 , 
    RI19a97820_2629 , 
    RI17478000_1151 , 
    RI174146b8_1408 , 
    RI17407170_1473 , 
    RI173be480_1828 , 
    RI17334f00_2183 , 
    RI174a3458_940 , 
    RI19ab4dd0_2417 , 
    RI1738ca70_2070 , 
    RI173c6b08_1787 , 
    RI1733d588_2142 , 
    RI1740f7f8_1432 , 
    RI19a90cc8_2677 , 
    RI17463150_1253 , 
    RI19ac1148_2322 , 
    RI174abe28_898 , 
    RI19aa48b8_2533 , 
    RI17480688_1110 , 
    RI19a85c10_2754 , 
    RI175019d0_755 , 
    RI173e4058_1644 , 
    RI1739b368_1999 , 
    RI1745be78_1288 , 
    RI19ab5f28_2409 , 
    RI174a1388_950 , 
    RI173f6460_1555 , 
    RI173ad770_1910 , 
    RI1752f060_620 , 
    RI19ab3c00_2425 , 
    RI17520330_666 , 
    RI19aac6d0_2480 , 
    RI17492a90_1021 , 
    RI173caca8_1767 , 
    RI17341728_2122 , 
    RI17413ce0_1411 , 
    RI19abf4b0_2338 , 
    RI174affc8_878 , 
    RI19a8e8b0_2693 , 
    RI174672f0_1233 , 
    RI19aac838_2479 , 
    RI17492dd8_1020 , 
    RI173e81f8_1624 , 
    RI1739f1c0_1980 , 
    RI1745fcd0_1269 , 
    RI19aa2248_2551 , 
    RI174844e0_1091 , 
    RI19a83438_2771 , 
    RI17509a40_736 , 
    RI174046c8_1486 , 
    RI17405730_1481 , 
    RI173bca40_1836 , 
    RI173334c0_2191 , 
    RI174a1a18_948 , 
    RI19ab63d8_2407 , 
    RI173a2cd0_1962 , 
    RI173dcd80_1679 , 
    RI17394090_2034 , 
    RI17454858_1324 , 
    RI19ac5e28_2285 , 
    RI174c7740_790 , 
    RI19a96038_2640 , 
    RI174793b0_1145 , 
    RI173fa2b8_1536 , 
    RI173b15c8_1891 , 
    RI17394db0_2030 , 
    RI19aa9d90_2497 , 
    RI174968e8_1002 , 
    RI19a9cc08_2592 , 
    RI17526528_647 , 
    RI19aa0358_2567 , 
    RI17488338_1072 , 
    RI19acef78_2218 , 
    RI1750fc38_717 , 
    RI173a3360_1960 , 
    RI173ec050_1605 , 
    RI1747c4e8_1130 , 
    RI19ac6080_2284 , 
    RI174c7c68_789 , 
    RI173ceb00_1748 , 
    RI17345238_2104 , 
    RI174465f0_1393 , 
    RI19abd6b0_2355 , 
    RI174b3ad8_860 , 
    RI19a8c240_2710 , 
    RI1746ae00_1215 , 
    RI19a8a2d8_2723 , 
    RI1746f630_1193 , 
    RI175361d0_598 , 
    RI1740d3e0_1443 , 
    RI173c46f0_1798 , 
    RI1733b170_2153 , 
    RI174a9a10_909 , 
    RI19ab1ef0_2440 , 
    RI173d3690_1725 , 
    RI1738a9a0_2080 , 
    RI1744b168_1370 , 
    RI19acb300_2246 , 
    RI174b8650_837 , 
    RI175385e8_592 , 
    RI17539218_590 , 
    RI17539e48_588 , 
    RI17537fd0_593 , 
    RI17536770_597 , 
    RI175379b8_594 , 
    RI17539830_589 , 
    RI174118c8_1422 , 
    RI173eda90_1597 , 
    RI17403318_1492 , 
    RI173ba628_1847 , 
    RI175342e0_604 , 
    RI19ab73c8_2400 , 
    RI1749f600_959 , 
    RI1744f650_1349 , 
    RI19a99f80_2612 , 
    RI17473e60_1171 , 
    RI19ac96e0_2259 , 
    RI174bf658_815 , 
    RI173d7b78_1704 , 
    RI1738ee88_2059 , 
    RI17400f00_1503 , 
    RI173f2608_1574 , 
    RI173a9918_1929 , 
    RI174be1b8_819 , 
    RI19aae7a0_2465 , 
    RI1748ec38_1040 , 
    RI19a23330_2795 , 
    RI1751a138_685 , 
    RI173ad428_1911 , 
    RI173e7b68_1626 , 
    RI1739eb30_1982 , 
    RI1745f640_1271 , 
    RI19a82f88_2773 , 
    RI17508ff0_738 , 
    RI19aa1f00_2553 , 
    RI17483e50_1093 , 
    RI173ffe98_1508 , 
    RI174050a0_1483 , 
    RI173bc3b0_1838 , 
    RI17332e30_2193 , 
    RI173e5750_1637 , 
    RI173f4048_1566 , 
    RI173ab358_1921 , 
    RI1750b408_731 , 
    RI19abcfa8_2359 , 
    RI1751ca78_677 , 
    RI19aad300_2474 , 
    RI17490678_1032 , 
    RI1744e5e8_1354 , 
    RI19acb120_2247 , 
    RI174bd768_821 , 
    RI19a9bd80_2599 , 
    RI17472df8_1176 , 
    RI173d6b10_1709 , 
    RI1738de20_2064 , 
    RI17497950_997 , 
    RI173eeaf8_1592 , 
    RI173a5e08_1947 , 
    RI19acc200_2238 , 
    RI17514468_703 , 
    RI19a9d400_2589 , 
    RI1748ade0_1059 , 
    RI173b2630_1886 , 
    RI173b6e60_1864 , 
    RI1740c030_1449 , 
    RI173c3340_1804 , 
    RI17339dc0_2159 , 
    RI19ab0ff0_2446 , 
    RI174a8660_915 , 
    RI1738cdb8_2069 , 
    RI173c7198_1785 , 
    RI1733dc18_2140 , 
    RI1740fe88_1430 , 
    RI19a90f20_2676 , 
    RI174637e0_1251 , 
    RI19ac12b0_2321 , 
    RI174ac4b8_896 , 
    RI173e43a0_1643 , 
    RI1739b6b0_1998 , 
    RI1745c1c0_1287 , 
    RI19a85e68_2753 , 
    RI17501ef8_754 , 
    RI19aa4a98_2532 , 
    RI174809d0_1109 , 
    RI173e4a30_1641 , 
    RI173f39b8_1568 , 
    RI173aacc8_1923 , 
    RI17502420_753 , 
    RI19a23150_2796 , 
    RI1751c028_679 , 
    RI19aaf628_2458 , 
    RI1748ffe8_1034 , 
    RI173c8200_1780 , 
    RI1733ec80_2135 , 
    RI17410ef0_1425 , 
    RI19ac1b98_2316 , 
    RI174ad520_891 , 
    RI19a919e8_2671 , 
    RI17464848_1246 , 
    RI173f6af0_1553 , 
    RI17404038_1488 , 
    RI173bb348_1843 , 
    RI17535780_600 , 
    RI174a0320_955 , 
    RI19ab7da0_2396 , 
    RI173f53f8_1560 , 
    RI173e6b00_1631 , 
    RI1739dac8_1987 , 
    RI1745e5d8_1276 , 
    RI19a84e00_2760 , 
    RI17507628_743 , 
    RI19aa3aa8_2540 , 
    RI17482de8_1098 , 
    RI173a3018_1961 , 
    RI173dd0c8_1678 , 
    RI173943d8_2033 , 
    RI17454ba0_1323 , 
    RI19a96290_2639 , 
    RI174796f8_1144 , 
    RI173b1910_1890 , 
    RI173fa600_1535 , 
    RI173971c8_2019 , 
    RI19a9e6c0_2581 , 
    RI17526a50_646 , 
    RI19aa9f70_2496 , 
    RI17496c30_1001 , 
    RI174a2dc8_942 , 
    RI173cf190_1746 , 
    RI173458c8_2102 , 
    RI17446c80_1391 , 
    RI19a8c6f0_2708 , 
    RI1746b490_1213 , 
    RI19abd9f8_2353 , 
    RI174b4168_858 , 
    RI173dd758_1676 , 
    RI173a39f0_1958 , 
    RI173ec6e0_1603 , 
    RI17480d18_1108 , 
    RI19acf428_2216 , 
    RI17510688_715 , 
    RI19aa0790_2565 , 
    RI174889c8_1070 , 
    RI1733c1d8_2148 , 
    RI173cb680_1764 , 
    RI173b6b18_1865 , 
    RI173ffb50_1509 , 
    RI1752eb38_621 , 
    RI1749be38_976 , 
    RI19ab9c18_2382 , 
    RI173d43b0_1721 , 
    RI1738b6c0_2076 , 
    RI1744be88_1366 , 
    RI19a9c848_2594 , 
    RI17470698_1188 , 
    RI19acba08_2242 , 
    RI174b9988_833 , 
    RI17450d48_1342 , 
    RI17408520_1467 , 
    RI173bf830_1822 , 
    RI173362b0_2177 , 
    RI174a4808_934 , 
    RI19ab34f8_2429 , 
    RI173ce470_1750 , 
    RI1744b7f8_1368 , 
    RI173c5410_1794 , 
    RI1740e100_1439 , 
    RI19a922d0_2667 , 
    RI17461a58_1260 , 
    RI19ac25e8_2311 , 
    RI174aa730_905 , 
    RI173e2960_1651 , 
    RI17399c70_2006 , 
    RI1745a780_1295 , 
    RI19a87218_2744 , 
    RI174d07a0_762 , 
    RI19aa5fb0_2523 , 
    RI1747ef90_1117 , 
    RI173ce128_1751 , 
    RI17344860_2107 , 
    RI17445c18_1396 , 
    RI19a8bbb0_2713 , 
    RI1746a428_1218 , 
    RI19abd188_2358 , 
    RI174b3100_863 , 
    RI173bf1a0_1824 , 
    RI19aabb90_2484 , 
    RI17495bc8_1006 , 
    RI19aaf448_2459 , 
    RI17525088_651 , 
    RI173f9598_1540 , 
    RI173b08a8_1895 , 
    RI1738bd50_2074 , 
    RI173fee30_1513 , 
    RI173b5df8_1869 , 
    RI173c2620_1808 , 
    RI1749b118_980 , 
    RI19aa7e28_2510 , 
    RI19a89e28_2725 , 
    RI1752d698_625 , 
    RI173a7500_1940 , 
    RI173988c0_2012 , 
    RI173e15b0_1657 , 
    RI174593d0_1301 , 
    RI19a93fe0_2654 , 
    RI1747dbe0_1123 , 
    RI19ac4280_2298 , 
    RI174ce8b0_768 , 
    RI17459a60_1299 , 
    RI17398f50_2010 , 
    RI173e1c40_1655 , 
    RI19a869a8_2748 , 
    RI174cf300_766 , 
    RI19aa5560_2527 , 
    RI1747e270_1121 , 
    RI173d3348_1726 , 
    RI1738a658_2081 , 
    RI1744ae20_1371 , 
    RI19abbe50_2368 , 
    RI174b8308_838 , 
    RI19ac4460_2297 , 
    RI174cedd8_767 , 
    RI173efea8_1586 , 
    RI17403660_1491 , 
    RI173ba970_1846 , 
    RI1749f948_958 , 
    RI19ab7530_2399 , 
    RI19a8fd50_2684 , 
    RI17465568_1242 , 
    RI1744f998_1348 , 
    RI19a9a160_2611 , 
    RI174741a8_1170 , 
    RI19ac9938_2258 , 
    RI174bfb80_814 , 
    RI173d7ec0_1703 , 
    RI1738f1d0_2058 , 
    RI17460d38_1264 , 
    RI17409f60_1459 , 
    RI173c1270_1814 , 
    RI17337cf0_2169 , 
    RI174a6590_925 , 
    RI19ab2148_2439 , 
    RI19aaa510_2493 , 
    RI17497608_998 , 
    RI173eca28_1602 , 
    RI173a3d38_1957 , 
    RI17483130_1097 , 
    RI19acf680_2215 , 
    RI17510bb0_714 , 
    RI19aa0970_2564 , 
    RI17488d10_1069 , 
    RI17335c20_2179 , 
    RI1745d570_1281 , 
    RI173d71a0_1707 , 
    RI1738e4b0_2062 , 
    RI1744ec78_1352 , 
    RI19a99698_2616 , 
    RI17473488_1174 , 
    RI19ac90c8_2262 , 
    RI174be6e0_818 , 
    RI173f4390_1565 , 
    RI173ab6a0_1920 , 
    RI1750ecc0_720 , 
    RI19abe2e0_2348 , 
    RI1751cfa0_676 , 
    RI19aad468_2473 , 
    RI174909c0_1031 , 
    RI19aa3238_2544 , 
    RI174820c8_1102 , 
    RI173d74e8_1706 , 
    RI1738e7f8_2061 , 
    RI1744efc0_1351 , 
    RI19ac92a8_2261 , 
    RI174bec08_817 , 
    RI19a998f0_2615 , 
    RI174737d0_1173 , 
    RI173f4a20_1563 , 
    RI173abd30_1918 , 
    RI17512aa0_708 , 
    RI19abf690_2337 , 
    RI1751d9f0_674 , 
    RI19aad648_2472 , 
    RI17491050_1029 , 
    RI173ddaa0_1675 , 
    RI174018d8_1500 , 
    RI173b8be8_1855 , 
    RI175319a0_612 , 
    RI1749dbc0_967 , 
    RI19ab8b38_2390 , 
    RI19a23678_2793 , 
    RI1751ab88_683 , 
    RI1744fce0_1347 , 
    RI173c98f8_1773 , 
    RI17340378_2128 , 
    RI17412930_1417 , 
    RI19a90188_2682 , 
    RI17465f40_1239 , 
    RI19ac0860_2327 , 
    RI174aec18_884 , 
    RI173e7190_1629 , 
    RI1739e158_1985 , 
    RI1745ec68_1274 , 
    RI19aa3c88_2539 , 
    RI17483478_1096 , 
    RI19a85058_2759 , 
    RI17508078_741 , 
    RI173cc6e8_1759 , 
    RI17343168_2114 , 
    RI17415720_1403 , 
    RI19a8d410_2702 , 
    RI17468d30_1225 , 
    RI19abe4c0_2347 , 
    RI174b1a08_870 , 
    RI1740fb40_1431 , 
    RI173f7ea0_1547 , 
    RI173af1b0_1902 , 
    RI1733d8d0_2141 , 
    RI19aa5a88_2525 , 
    RI17522c70_658 , 
    RI19aaac18_2490 , 
    RI174944d0_1013 , 
    RI17444ef8_1400 , 
    RI173dc060_1683 , 
    RI17393370_2038 , 
    RI17453b38_1328 , 
    RI19ac7b38_2272 , 
    RI174c62a0_794 , 
    RI19a97dc0_2627 , 
    RI17478690_1149 , 
    RI17447ce8_1386 , 
    RI17407800_1471 , 
    RI173beb10_1826 , 
    RI17335590_2181 , 
    RI174a3ae8_938 , 
    RI19ab52f8_2415 , 
    RI173d8f28_1698 , 
    RI17390238_2053 , 
    RI17450a00_1343 , 
    RI19a98630_2623 , 
    RI17475210_1165 , 
    RI19ac81c8_2269 , 
    RI174c1548_809 , 
    RI19ab4380_2422 , 
    RI174a5f00_927 , 
    RI173fac90_1533 , 
    RI173b1fa0_1888 , 
    RI1739b9f8_1997 , 
    RI19aa12d0_2559 , 
    RI175274a0_644 , 
    RI19aaa330_2494 , 
    RI174972c0_999 , 
    RI173cf820_1744 , 
    RI17345f58_2100 , 
    RI17447310_1389 , 
    RI19abddb8_2351 , 
    RI174b47f8_856 , 
    RI19a8cb28_2706 , 
    RI1746bb20_1211 , 
    RI19abcdc8_2360 , 
    RI174b6580_847 , 
    RI173e0200_1663 , 
    RI17397510_2018 , 
    RI17458020_1307 , 
    RI19ac3290_2305 , 
    RI174cc9c0_774 , 
    RI19a93068_2661 , 
    RI1747c830_1129 , 
    RI174c8be0_786 , 
    RI173dfeb8_1664 , 
    RI17401c20_1499 , 
    RI173b8f30_1854 , 
    RI17531ec8_611 , 
    RI1749df08_966 , 
    RI19ab8d90_2389 , 
    RI17453160_1331 , 
    RI17408868_1466 , 
    RI173bfb78_1821 , 
    RI173365f8_2176 , 
    RI174a4b50_933 , 
    RI19ab36d8_2428 , 
    RI173f9c28_1538 , 
    RI173eb330_1609 , 
    RI173a2640_1964 , 
    RI17475558_1164 , 
    RI19a9fae8_2571 , 
    RI17487618_1076 , 
    RI19ace870_2221 , 
    RI1750e798_721 , 
    RI173a7848_1939 , 
    RI17398c08_2011 , 
    RI173e18f8_1656 , 
    RI17459718_1300 , 
    RI19a94238_2653 , 
    RI1747df28_1122 , 
    RI174a9d58_908 , 
    RI173f0880_1583 , 
    RI173a7b90_1938 , 
    RI19aafad8_2456 , 
    RI1748cb68_1050 , 
    RI19a85508_2757 , 
    RI175172d0_694 , 
    RI17340a08_2126 , 
    RI173f8f08_1542 , 
    RI17404380_1487 , 
    RI173bb690_1842 , 
    RI17535ca8_599 , 
    RI174a0668_954 , 
    RI19ab7f80_2395 , 
    RI173d8be0_1699 , 
    RI1738fef0_2054 , 
    RI174506b8_1344 , 
    RI19a983d8_2624 , 
    RI17474ec8_1166 , 
    RI19ac7f70_2270 , 
    RI174c1020_810 , 
    RI173e2618_1652 , 
    RI17399928_2007 , 
    RI1745a438_1296 , 
    RI19a86fc0_2745 , 
    RI174d0278_763 , 
    RI19aa5dd0_2524 , 
    RI1747ec48_1118 , 
    RI173d39d8_1724 , 
    RI173c50c8_1795 , 
    RI1733bb48_2150 , 
    RI1740ddb8_1440 , 
    RI19ac2390_2312 , 
    RI174aa3e8_906 , 
    RI19a920f0_2668 , 
    RI17461710_1261 , 
    RI17335f68_2178 , 
    RI173b0bf0_1894 , 
    RI173f98e0_1539 , 
    RI1738e168_2063 , 
    RI19a981f8_2625 , 
    RI175255b0_650 , 
    RI19aa9688_2500 , 
    RI17495f10_1005 , 
    RI17344ba8_2106 , 
    RI17445f60_1395 , 
    RI19abd2f0_2357 , 
    RI174b3448_862 , 
    RI19a8be08_2712 , 
    RI1746a770_1217 , 
    RI173d2cb8_1728 , 
    RI17411f58_1420 , 
    RI173c4060_1800 , 
    RI1740cd50_1445 , 
    RI1733aae0_2155 , 
    RI174a9380_911 , 
    RI19ab1860_2442 , 
    RI173c39d0_1802 , 
    RI173fe110_1517 , 
    RI173b50d8_1873 , 
    RI173b95c0_1852 , 
    RI19a88460_2736 , 
    RI1752c1f8_629 , 
    RI19aa71f8_2515 , 
    RI1749a3f8_984 , 
    RI173d2970_1729 , 
    RI17389c80_2084 , 
    RI1744a448_1374 , 
    RI19a89888_2727 , 
    RI1746ec58_1196 , 
    RI19abb5e0_2372 , 
    RI174b7930_841 , 
    RI19a23858_2792 , 
    RI1751b0b0_682 , 
    RI173915e8_2047 , 
    RI173cb9c8_1763 , 
    RI17342448_2118 , 
    RI17414a00_1407 , 
    RI19a8f210_2689 , 
    RI17468010_1229 , 
    RI19abfc30_2334 , 
    RI174b0ce8_874 , 
    RI173e8f18_1620 , 
    RI1739fee0_1976 , 
    RI174609f0_1265 , 
    RI19aa2e78_2546 , 
    RI17485200_1087 , 
    RI19a83f78_2766 , 
    RI1750aee0_732 , 
    RI173e9f80_1615 , 
    RI173db340_1687 , 
    RI17392650_2042 , 
    RI17452e18_1332 , 
    RI19ac74a8_2275 , 
    RI174c4e00_798 , 
    RI19a976b8_2630 , 
    RI17477628_1154 , 
    RI173f8878_1544 , 
    RI173afb88_1899 , 
    RI17344518_2108 , 
    RI19aaa858_2492 , 
    RI17523be8_655 , 
    RI19aab410_2487 , 
    RI17494ea8_1010 , 
    RI19abaa28_2376 , 
    RI174b68c8_846 , 
    RI173a0228_1975 , 
    RI1740bce8_1450 , 
    RI173c2ff8_1805 , 
    RI17339a78_2160 , 
    RI19ab0e10_2447 , 
    RI174a8318_916 , 
    RI173e0548_1662 , 
    RI17397858_2017 , 
    RI17458368_1306 , 
    RI19ac34e8_2304 , 
    RI174ccee8_773 , 
    RI19a932c0_2660 , 
    RI1747cb78_1128 , 
    RI173b1c58_1889 , 
    RI174098d0_1461 , 
    RI173c0be0_1816 , 
    RI17337660_2171 , 
    RI1745c508_1286 , 
    RI173f6e38_1552 , 
    RI173ae148_1907 , 
    RI17332458_2196 , 
    RI19aaca18_2478 , 
    RI17493468_1018 , 
    RI19ab6cc0_2403 , 
    RI175212a8_663 , 
    RI173cb338_1765 , 
    RI17341db8_2120 , 
    RI17414370_1409 , 
    RI19a8efb8_2690 , 
    RI17467980_1231 , 
    RI19abfa50_2335 , 
    RI174b0658_876 , 
    RI19a831e0_2772 , 
    RI17509518_737 , 
    RI173d95b8_1696 , 
    RI173908c8_2051 , 
    RI17451090_1341 , 
    RI19ac8330_2268 , 
    RI174c1f98_807 , 
    RI19a98888_2622 , 
    RI174758a0_1163 , 
    RI19ab54d8_2414 , 
    RI17520858_665 , 
    RI173f67a8_1554 , 
    RI173adab8_1909 , 
    RI17532918_609 , 
    RI17411238_1424 , 
    RI173e9260_1619 , 
    RI17402c88_1494 , 
    RI173b9f98_1849 , 
    RI17533890_606 , 
    RI1749ef70_961 , 
    RI19ab7008_2402 , 
    RI17400870_1505 , 
    RI173c6478_1789 , 
    RI1733cef8_2144 , 
    RI1740f168_1434 , 
    RI19ac30b0_2306 , 
    RI174ab798_900 , 
    RI19a92e10_2662 , 
    RI17462ac0_1255 , 
    RI173acd98_1913 , 
    RI173e74d8_1628 , 
    RI1739e4a0_1984 , 
    RI1745efb0_1273 , 
    RI19aa3ee0_2538 , 
    RI174837c0_1095 , 
    RI19a852b0_2758 , 
    RI175085a0_740 , 
    RI173fb668_1530 , 
    RI17404a10_1485 , 
    RI173bbd20_1840 , 
    RI173327a0_2195 , 
    RI174a0cf8_952 , 
    RI19ab5a00_2411 , 
    RI1733f9a0_2131 , 
    RI173c8f20_1776 , 
    RI17411c10_1421 , 
    RI19ac04a0_2329 , 
    RI174ae240_887 , 
    RI173c6e50_1786 , 
    RI173b6488_1867 , 
    RI173ff4c0_1511 , 
    RI1752e0e8_623 , 
    RI1749b7a8_978 , 
    RI19ab98d0_2384 , 
    RI173d3d20_1723 , 
    RI1738b030_2078 , 
    RI19acb648_2244 , 
    RI174b8f38_835 , 
    RI19a9c398_2596 , 
    RI17470008_1190 , 
    RI173f22c0_1575 , 
    RI174039a8_1490 , 
    RI173bacb8_1845 , 
    RI17534d30_602 , 
    RI1749fc90_957 , 
    RI19ab7878_2398 , 
    RI173e6470_1633 , 
    RI1739d438_1989 , 
    RI1745df48_1278 , 
    RI19a84950_2762 , 
    RI17506bd8_745 , 
    RI19aa3580_2542 , 
    RI17482758_1100 , 
    RI173f9f70_1537 , 
    RI173b1280_1892 , 
    RI17392998_2041 , 
    RI19a9b420_2603 , 
    RI17526000_648 , 
    RI19aa9bb0_2498 , 
    RI174965a0_1003 , 
    RI173dca38_1680 , 
    RI17393d48_2035 , 
    RI17454510_1325 , 
    RI19a95de0_2641 , 
    RI17479068_1146 , 
    RI174c7218_791 , 
    RI19ac5bd0_2286 , 
    RI173ebd08_1606 , 
    RI1747a0d0_1141 , 
    RI19aa0100_2568 , 
    RI17487ff0_1073 , 
    RI19aced20_2219 , 
    RI1750f710_718 , 
    RI173ce7b8_1749 , 
    RI17344ef0_2105 , 
    RI174462a8_1394 , 
    RI19a8bfe8_2711 , 
    RI1746aab8_1216 , 
    RI19abd4d0_2356 , 
    RI174b3790_861 , 
    RI173cd408_1755 , 
    RI17343e88_2110 , 
    RI17445240_1399 , 
    RI19a8dd70_2698 , 
    RI17469a50_1221 , 
    RI19abebc8_2343 , 
    RI174b2728_866 , 
    RI173f8bc0_1543 , 
    RI173afed0_1898 , 
    RI17346930_2097 , 
    RI19aac388_2481 , 
    RI17524110_654 , 
    RI19aab5f0_2486 , 
    RI174951f0_1009 , 
    RI173dc6f0_1681 , 
    RI17393a00_2036 , 
    RI174541c8_1326 , 
    RI19a95b88_2642 , 
    RI17478d20_1147 , 
    RI19ac5978_2287 , 
    RI174c6cf0_792 , 
    RI17407e90_1469 , 
    RI1744c518_1364 , 
    RI19ab5820_2412 , 
    RI174a4178_936 , 
    RI17332110_2197 , 
    RI1740b658_1452 , 
    RI173c2968_1807 , 
    RI19ab2f58_2432 , 
    RI174a7c88_918 , 
    RI173393e8_2162 , 
    RI19a93518_2659 , 
    RI17529de0_636 , 
    RI173a5430_1950 , 
    RI173ee120_1595 , 
    RI17490d08_1030 , 
    RI19a9f368_2575 , 
    RI1748a408_1062 , 
    RI19acdf10_2225 , 
    RI175134f0_706 , 
    RI19a87470_2743 , 
    RI174d0cc8_761 , 
    RI173f18e8_1578 , 
    RI173a8bf8_1933 , 
    RI174b51d0_853 , 
    RI19ab0528_2451 , 
    RI1748dbd0_1045 , 
    RI19ab3a20_2426 , 
    RI17518c98_689 , 
    RI174122a0_1419 , 
    RI173be138_1829 , 
    RI17406e28_1474 , 
    RI17334bb8_2184 , 
    RI19ab4bf0_2418 , 
    RI174a3110_941 , 
    RI1738c728_2071 , 
    RI173c67c0_1788 , 
    RI1733d240_2143 , 
    RI1740f4b0_1433 , 
    RI19a90a70_2678 , 
    RI17462e08_1254 , 
    RI19ac0f68_2323 , 
    RI174abae0_899 , 
    RI173e3d10_1645 , 
    RI1739b020_2000 , 
    RI1745bb30_1289 , 
    RI175014a8_756 , 
    RI19aa46d8_2534 , 
    RI17480340_1111 , 
    RI173e50c0_1639 , 
    RI173d6480_1711 , 
    RI1738d790_2066 , 
    RI1744df58_1356 , 
    RI19acadd8_2249 , 
    RI174bcd18_823 , 
    RI19a9b8d0_2601 , 
    RI17472768_1178 , 
    RI17400bb8_1504 , 
    RI173f1f78_1576 , 
    RI173a9288_1931 , 
    RI174ba3d8_831 , 
    RI19ab0a50_2449 , 
    RI1748e260_1043 , 
    RI19ad0238_2210 , 
    RI175196e8_687 , 
    RI173eb678_1608 , 
    RI173ba2e0_1848 , 
    RI17402fd0_1493 , 
    RI17533db8_605 , 
    RI1749f2b8_960 , 
    RI19ab71e8_2401 , 
    RI17411580_1423 , 
    RI173d7830_1705 , 
    RI1738eb40_2060 , 
    RI1744f308_1350 , 
    RI19ac9500_2260 , 
    RI174bf130_816 , 
    RI19a99d28_2613 , 
    RI17473b18_1172 , 
    RI173b0218_1897 , 
    RI173ee7b0_1593 , 
    RI173a5ac0_1948 , 
    RI17495538_1008 , 
    RI19ace3c0_2223 , 
    RI17513f40_704 , 
    RI19a9f728_2573 , 
    RI1748aa98_1060 , 
    RI173e5408_1638 , 
    RI173f3d00_1567 , 
    RI173ab010_1922 , 
    RI17507b50_742 , 
    RI19aaf790_2457 , 
    RI17490330_1033 , 
    RI19a83b40_2768 , 
    RI1751c550_678 , 
    RI1744e2a0_1355 , 
    RI173d67c8_1710 , 
    RI1738dad8_2065 , 
    RI19acaf40_2248 , 
    RI174bd240_822 , 
    RI19a9bb28_2600 , 
    RI17472ab0_1177 , 
    RI1744b4b0_1369 , 
    RI1744e930_1353 , 
    RI174081d8_1468 , 
    RI173bf4e8_1823 , 
    RI174a44c0_935 , 
    RI19ab3318_2430 , 
    RI173f50b0_1561 , 
    RI173e67b8_1632 , 
    RI1739d780_1988 , 
    RI1745e290_1277 , 
    RI19a84ba8_2761 , 
    RI17507100_744 , 
    RI19aa38c8_2541 , 
    RI17482aa0_1099 , 
    RI173f46d8_1564 , 
    RI17403cf0_1489 , 
    RI173bb000_1844 , 
    RI17535258_601 , 
    RI1749ffd8_956 , 
    RI19ab7a58_2397 , 
    RI173e22d0_1653 , 
    RI173f3670_1569 , 
    RI173aa980_1924 , 
    RI174cfd50_764 , 
    RI19a23c18_2790 , 
    RI1751bb00_680 , 
    RI19aaf268_2460 , 
    RI1748fca0_1035 , 
    RI173c7eb8_1781 , 
    RI1733e938_2136 , 
    RI17410ba8_1426 , 
    RI19a91808_2672 , 
    RI17464500_1247 , 
    RI19ac1a30_2317 , 
    RI174ad1d8_892 , 
    RI173e0f20_1659 , 
    RI17398230_2014 , 
    RI17458d40_1303 , 
    RI19ac3d58_2300 , 
    RI174cde60_770 , 
    RI19a93ba8_2656 , 
    RI1747d550_1125 , 
    RI174a09b0_953 , 
    RI173fe7a0_1515 , 
    RI173b5768_1871 , 
    RI173bddf0_1830 , 
    RI19a88be0_2733 , 
    RI1752cc48_627 , 
    RI19aa7a68_2512 , 
    RI1749aa88_982 , 
    RI173ac708_1915 , 
    RI1751d4c8_675 , 
    RI19ac36c8_2303 , 
    RI1751e968_671 , 
    RI19aadfa8_2468 , 
    RI17491a28_1026 , 
    RI173e2ff0_1649 , 
    RI1739a300_2004 , 
    RI1745ae10_1293 , 
    RI19aa62f8_2521 , 
    RI1747f620_1115 , 
    RI173c5aa0_1792 , 
    RI1733c520_2147 , 
    RI1740e790_1437 , 
    RI19a92708_2665 , 
    RI174620e8_1258 , 
    RI19ac2a98_2309 , 
    RI174aadc0_903 , 
    RI173d9900_1695 , 
    RI17390c10_2050 , 
    RI19ac8510_2267 , 
    RI174c24c0_806 , 
    RI19a98ae0_2621 , 
    RI17475be8_1162 , 
    RI174513d8_1340 , 
    RI173413e0_2123 , 
    RI17337318_2172 , 
    RI1745a0f0_1297 , 
    RI174a5bb8_928 , 
    RI19ab4038_2423 , 
    RI173c0898_1817 , 
    RI17409588_1462 , 
    RI173f1258_1580 , 
    RI173a8568_1935 , 
    RI174b09a0_875 , 
    RI19a94df0_2648 , 
    RI17518248_691 , 
    RI19ab01e0_2453 , 
    RI1748d540_1047 , 
    RI173c5758_1793 , 
    RI1740e448_1438 , 
    RI19a92528_2666 , 
    RI17461da0_1259 , 
    RI19ac2840_2310 , 
    RI174aaa78_904 , 
    RI173e2ca8_1650 , 
    RI17399fb8_2005 , 
    RI1745aac8_1294 , 
    RI19aa6190_2522 , 
    RI1747f2d8_1116 , 
    RI17336940_2175 , 
    RI173c43a8_1799 , 
    RI173c4a38_1797 , 
    RI173ff178_1512 , 
    RI173b6140_1868 , 
    RI1752dbc0_624 , 
    RI1749b460_979 , 
    RI19ab96f0_2385 , 
    RI1738ace8_2079 , 
    RI19acb4e0_2245 , 
    RI174b8a10_836 , 
    RI19a9c1b8_2597 , 
    RI1746fcc0_1191 , 
    RI1739c3d0_1994 , 
    RI1745cee0_1283 , 
    RI19a864f8_2750 , 
    RI17503398_750 , 
    RI19aa5218_2529 , 
    RI174816f0_1105 , 
    RI17402940_1495 , 
    RI173b9c50_1850 , 
    RI17533368_607 , 
    RI173e6e48_1630 , 
    RI19ab9498_2386 , 
    RI1749ec28_962 , 
    RI19a838e8_2769 , 
    RI1750a490_734 , 
    RI173d9f90_1693 , 
    RI173912a0_2048 , 
    RI17451a68_1338 , 
    RI19a98f90_2619 , 
    RI17476278_1160 , 
    RI19ac89c0_2265 , 
    RI174c2f10_804 , 
    RI173f74c8_1550 , 
    RI173ae7d8_1905 , 
    RI17336c88_2174 , 
    RI19aacdd8_2476 , 
    RI17493af8_1016 , 
    RI19ab9df8_2381 , 
    RI17521cf8_661 , 
    RI173b2978_1885 , 
    RI17485548_1086 , 
    RI19a9e8a0_2580 , 
    RI17489058_1068 , 
    RI19acd358_2230 , 
    RI175110d8_713 , 
    RI173ecd70_1601 , 
    RI173a4080_1956 , 
    RI17477970_1153 , 
    RI1740a2a8_1458 , 
    RI173c15b8_1813 , 
    RI17338038_2168 , 
    RI174a68d8_924 , 
    RI19ab2328_2438 , 
    RI17406108_1478 , 
    RI173aeb20_1904 , 
    RI173f7810_1549 , 
    RI173390a0_2163 , 
    RI19aad120_2475 , 
    RI17493e40_1015 , 
    RI19abba90_2370 , 
    RI17522220_660 , 
    RI173cc058_1761 , 
    RI17342ad8_2116 , 
    RI17415090_1405 , 
    RI19a8cd80_2705 , 
    RI174686a0_1227 , 
    RI19abdf98_2350 , 
    RI174b1378_872 , 
    RI19abb298_2373 , 
    RI174b72a0_843 , 
    RI173e46e8_1642 , 
    RI1740c6c0_1447 , 
    RI1733a450_2157 , 
    RI174a8cf0_913 , 
    RI19ab1518_2444 , 
    RI17391fc0_2044 , 
    RI173cc3a0_1760 , 
    RI17342e20_2115 , 
    RI174153d8_1404 , 
    RI19a8cfd8_2704 , 
    RI174689e8_1226 , 
    RI19abe100_2349 , 
    RI174b16c0_871 , 
    RI173a0f48_1971 , 
    RI173e9c38_1616 , 
    RI174658b0_1241 , 
    RI19acfd88_2212 , 
    RI1750c380_728 , 
    RI19aa0f10_2561 , 
    RI17485f20_1083 , 
    RI173ea958_1612 , 
    RI173fa948_1534 , 
    RI1744a100_1375 , 
    RI19a8e220_2696 , 
    RI17466918_1236 , 
    RI173d8208_1702 , 
    RI1738f518_2057 , 
    RI19ac9b90_2257 , 
    RI174c00a8_813 , 
    RI19a9a3b8_2610 , 
    RI174744f0_1169 , 
    RI173f5740_1559 , 
    RI173aca50_1914 , 
    RI17520d80_664 , 
    RI19aae110_2467 , 
    RI17491d70_1025 , 
    RI19ac4f28_2292 , 
    RI1751ee90_670 , 
    RI19aa8bc0_2505 , 
    RI174989b8_992 , 
    RI173a50e8_1951 , 
    RI173eddd8_1596 , 
    RI1748e8f0_1041 , 
    RI19acdcb8_2226 , 
    RI17512fc8_707 , 
    RI19a9f188_2576 , 
    RI1748a0c0_1063 , 
    RI17512578_709 , 
    RI1740afc8_1454 , 
    RI173c22d8_1809 , 
    RI17338d58_2164 , 
    RI19ab2d78_2433 , 
    RI174a75f8_920 , 
    RI173c5de8_1791 , 
    RI1733c868_2146 , 
    RI1740ead8_1436 , 
    RI19ac2cf0_2308 , 
    RI174ab108_902 , 
    RI19a92960_2664 , 
    RI17462430_1257 , 
    RI173e3338_1648 , 
    RI1739a648_2003 , 
    RI1745b158_1292 , 
    RI19a87920_2741 , 
    RI17500530_759 , 
    RI19aa6640_2520 , 
    RI1747f968_1114 , 
    RI173f5a88_1558 , 
    RI17524638_653 , 
    RI19aae458_2466 , 
    RI174920b8_1024 , 
    RI19ac6878_2281 , 
    RI1751f3b8_669 , 
    RI17450028_1346 , 
    RI19ac9de8_2256 , 
    RI174c05d0_812 , 
    RI19a9a610_2609 , 
    RI17474838_1168 , 
    RI173d8550_1701 , 
    RI1738f860_2056 , 
    RI173ca960_1768 , 
    RI17413998_1412 , 
    RI19abf2d0_2339 , 
    RI174afc80_879 , 
    RI19a8e6d0_2694 , 
    RI17466fa8_1234 , 
    RI173ca618_1769 , 
    RI17341098_2124 , 
    RI17413650_1413 , 
    RI19abf0f0_2340 , 
    RI174af938_880 , 
    RI19a8e478_2695 , 
    RI17466c60_1235 , 
    RI173e7eb0_1625 , 
    RI1739ee78_1981 , 
    RI1745f988_1270 , 
    RI19aa2068_2552 , 
    RI17484198_1092 , 
    RI17406450_1477 , 
    RI173f7b58_1548 , 
    RI173aee68_1903 , 
    RI1733b4b8_2152 , 
    RI19aaaa38_2491 , 
    RI17494188_1014 , 
    RI19aa4318_2536 , 
    RI17522748_659 , 
    RI19ab29b8_2435 , 
    RI174a6f68_922 , 
    RI173fc388_1526 , 
    RI173b3350_1882 , 
    RI173a71b8_1941 , 
    RI19a90368_2681 , 
    RI17529390_638 , 
    RI19aa8878_2506 , 
    RI17498670_993 , 
    RI173d0bd0_1738 , 
    RI17347308_2094 , 
    RI174486c0_1383 , 
    RI19a8af08_2718 , 
    RI1746ced0_1205 , 
    RI19abc8a0_2363 , 
    RI174b5ba8_850 , 
    RI1739ca60_1992 , 
    RI173e5a98_1636 , 
    RI19a841d0_2765 , 
    RI17503de8_748 , 
    RI19aa3058_2545 , 
    RI17481d80_1103 , 
    RI173eaca0_1611 , 
    RI173dc3a8_1682 , 
    RI173936b8_2037 , 
    RI17453e80_1327 , 
    RI19ac7d90_2271 , 
    RI174c67c8_793 , 
    RI19a98018_2626 , 
    RI174789d8_1148 , 
    RI173406c0_2127 , 
    RI17450370_1345 , 
    RI19aca040_2255 , 
    RI174c0af8_811 , 
    RI19a9a868_2608 , 
    RI17474b80_1167 , 
    RI173d8898_1700 , 
    RI1738fba8_2055 , 
    RI173a22f8_1965 , 
    RI173eafe8_1610 , 
    RI17473140_1175 , 
    RI19a9f908_2572 , 
    RI174872d0_1077 , 
    RI19ace618_2222 , 
    RI1750e270_722 , 
    RI173fb320_1531 , 
    RI1740ca08_1446 , 
    RI173c3d18_1801 , 
    RI1733a798_2156 , 
    RI174a9038_912 , 
    RI19ab16f8_2443 , 
    RI173c3688_1803 , 
    RI173fddc8_1518 , 
    RI173b4d90_1874 , 
    RI173b71a8_1863 , 
    RI19a88208_2737 , 
    RI1752bcd0_630 , 
    RI19aa7090_2516 , 
    RI1749a0b0_985 , 
    RI173d22e0_1731 , 
    RI173892a8_2087 , 
    RI17449db8_1376 , 
    RI19a89720_2728 , 
    RI1746e5c8_1198 , 
    RI173daff8_1688 , 
    RI17392308_2043 , 
    RI17452ad0_1333 , 
    RI19ac7250_2276 , 
    RI174c48d8_799 , 
    RI19a97460_2631 , 
    RI174772e0_1155 , 
    RI173f8530_1545 , 
    RI173af840_1900 , 
    RI17342100_2119 , 
    RI19aa8f80_2503 , 
    RI175236c0_656 , 
    RI19aab0c8_2488 , 
    RI17494b60_1011 , 
    RI173e8bd0_1621 , 
    RI1739fb98_1977 , 
    RI174606a8_1266 , 
    RI19aa2c20_2547 , 
    RI17484eb8_1088 , 
    RI19a83d20_2767 , 
    RI1750a9b8_733 , 
    RI173caff0_1766 , 
    RI17341a70_2121 , 
    RI17414028_1410 , 
    RI19a8ed60_2691 , 
    RI17467638_1232 , 
    RI19abf870_2336 , 
    RI174b0310_877 , 
    RI174053e8_1482 , 
    RI173a6e70_1942 , 
    RI173a1fb0_1966 , 
    RI17470d28_1186 , 
    RI19aa19d8_2555 , 
    RI17486f88_1078 , 
    RI19a82b50_2775 , 
    RI1750dd48_723 , 
    RI173f0538_1584 , 
    RI19acd100_2231 , 
    RI17516da8_695 , 
    RI19a9e468_2582 , 
    RI1748c820_1051 , 
    RI174a7940_919 , 
    RI173d3000_1727 , 
    RI1738a310_2082 , 
    RI1744aad8_1372 , 
    RI19abbc70_2369 , 
    RI174b7fc0_839 , 
    RI19a8a080_2724 , 
    RI1746f2e8_1194 , 
    RI17457cd8_1308 , 
    RI17409240_1463 , 
    RI173c0550_1818 , 
    RI17336fd0_2173 , 
    RI174a5870_929 , 
    RI19ab3de0_2424 , 
    RI173f6118_1556 , 
    RI1752b7a8_631 , 
    RI19ab2508_2437 , 
    RI1751fe08_667 , 
    RI19aac040_2482 , 
    RI17492748_1022 , 
    RI173db688_1686 , 
    RI173b88a0_1856 , 
    RI17401590_1501 , 
    RI17531478_613 , 
    RI1749d878_968 , 
    RI19ab8958_2391 , 
    RI1751a660_684 , 
    RI19a88028_2738 , 
    RI1752b280_632 , 
    RI19aa6d48_2517 , 
    RI17499a20_987 , 
    RI173fd738_1520 , 
    RI173b4700_1876 , 
    RI173b4a48_1875 , 
    RI173d1f98_1732 , 
    RI173599e0_2088 , 
    RI17449a70_1377 , 
    RI19a894c8_2729 , 
    RI1746e280_1199 , 
    RI19abaf50_2374 , 
    RI174b6f58_844 , 
    RI19abcbe8_2361 , 
    RI174b6238_848 , 
    RI173dfb70_1665 , 
    RI17396e80_2020 , 
    RI17457648_1310 , 
    RI19a95930_2643 , 
    RI1747c1a0_1131 , 
    RI19ac5720_2288 , 
    RI174cbf70_776 , 
    RI17390f58_2049 , 
    RI173e8888_1622 , 
    RI1739f850_1978 , 
    RI17460360_1267 , 
    RI19aa27e8_2549 , 
    RI17484b70_1089 , 
    RI173cf4d8_1745 , 
    RI17345c10_2101 , 
    RI17446fc8_1390 , 
    RI19a8c948_2707 , 
    RI1746b7d8_1212 , 
    RI19abdbd8_2352 , 
    RI174b44b0_857 , 
    RI173995e0_2008 , 
    RI19a9fcc8_2570 , 
    RI17526f78_645 , 
    RI19aaa150_2495 , 
    RI17496f78_1000 , 
    RI173358d8_2180 , 
    RI17409c18_1460 , 
    RI173c0f28_1815 , 
    RI173379a8_2170 , 
    RI1745e920_1275 , 
    RI174a6248_926 , 
    RI19ab4560_2421 , 
    RI19a8faf8_2685 , 
    RI17465220_1243 , 
    RI1740a5f0_1457 , 
    RI173fc040_1527 , 
    RI173b3008_1883 , 
    RI173a4da0_1952 , 
    RI19aa8530_2507 , 
    RI17498328_994 , 
    RI19a8eb08_2692 , 
    RI17528e68_639 , 
    RI173d0888_1739 , 
    RI17346fc0_2095 , 
    RI17448378_1384 , 
    RI19a8acb0_2719 , 
    RI1746cb88_1206 , 
    RI19abc6c0_2364 , 
    RI174b5860_851 , 
    RI1733fce8_2130 , 
    RI173eee40_1591 , 
    RI173964a8_2023 , 
    RI173cdde0_1752 , 
    RI174001e0_1507 , 
    RI173b74f0_1862 , 
    RI1752f588_619 , 
    RI1749c4c8_974 , 
    RI19aba050_2380 , 
    RI173d1c50_1733 , 
    RI17359698_2089 , 
    RI17449728_1378 , 
    RI19a89270_2730 , 
    RI1746df38_1200 , 
    RI19abad70_2375 , 
    RI174b6c10_845 , 
    RI173fd3f0_1521 , 
    RI173b43b8_1877 , 
    RI19a87dd0_2739 , 
    RI1752ad58_633 , 
    RI19aa6b68_2518 , 
    RI174996d8_988 , 
    RI173c9f88_1771 , 
    RI17412fc0_1415 , 
    RI19ac0d88_2324 , 
    RI174af2a8_882 , 
    RI19a90818_2679 , 
    RI174665d0_1237 , 
    RI173ddde8_1674 , 
    RI173950f8_2029 , 
    RI174558c0_1319 , 
    RI19a96bf0_2635 , 
    RI1747a418_1140 , 
    RI19ac69e0_2280 , 
    RI174c9108_785 , 
    RI173c8bd8_1777 , 
    RI1733f658_2132 , 
    RI19ac0338_2330 , 
    RI174adef8_888 , 
    RI17454ee8_1322 , 
    RI17455578_1320 , 
    RI17408bb0_1465 , 
    RI173bfec0_1820 , 
    RI174a4e98_932 , 
    RI19ab3840_2427 , 
    RI17394720_2032 , 
    RI19a964e8_2638 , 
    RI17479a40_1143 , 
    RI19ac63c8_2283 , 
    RI174c8190_788 , 
    RI173d6e58_1708 , 
    RI173b8210_1858 , 
    RI17530a28_615 , 
    RI1749d1e8_970 , 
    RI19ab82c8_2394 , 
    RI1739a990_2002 , 
    RI173e3680_1647 , 
    RI1745b4a0_1291 , 
    RI19a87b78_2740 , 
    RI17500a58_758 , 
    RI19aa6988_2519 , 
    RI1747fcb0_1113 , 
    RI173b0f38_1893 , 
    RI17390580_2052 , 
    RI19a99ad0_2614 , 
    RI17525ad8_649 , 
    RI19aa9868_2499 , 
    RI17496258_1004 , 
    RI19aa7540_2514 , 
    RI17523198_657 , 
    RI17455230_1321 , 
    RI19acd5b0_2229 , 
    RI17511600_712 , 
    RI17395ad0_2026 , 
    RI173de7c0_1671 , 
    RI17456298_1316 , 
    RI19a946e8_2651 , 
    RI1747adf0_1137 , 
    RI19ac4910_2295 , 
    RI174ca080_782 , 
    RI1744a790_1373 , 
    RI1749cb58_972 , 
    RI19aba578_2378 , 
    RI173a1290_1970 , 
    RI17467cc8_1230 , 
    RI19aa10f0_2560 , 
    RI17486268_1082 , 
    RI19acffe0_2211 , 
    RI1750c8a8_727 , 
    RI174458d0_1397 , 
    RI174074b8_1472 , 
    RI173be7c8_1827 , 
    RI19ab5118_2416 , 
    RI174a37a0_939 , 
    RI17335248_2182 , 
    RI1733f310_2133 , 
    RI19a9e288_2583 , 
    RI1748c4d8_1052 , 
    RI19a96998_2636 , 
    RI1752a830_634 , 
    RI173ac3c0_1916 , 
    RI17519c10_686 , 
    RI19aadd50_2469 , 
    RI174916e0_1027 , 
    RI19ac1f58_2314 , 
    RI1751e440_672 , 
    RI17406ae0_1475 , 
    RI17405a78_1480 , 
    RI173bcd88_1835 , 
    RI17333808_2190 , 
    RI174a1d60_947 , 
    RI19ab65b8_2406 , 
    RI173e8540_1623 , 
    RI1739f508_1979 , 
    RI17460018_1268 , 
    RI19aa24a0_2550 , 
    RI17484828_1090 , 
    RI19a83690_2770 , 
    RI17509f68_735 , 
    RI175373a0_595 , 
    RI1753a460_587 , 
    RI19abe808_2345 , 
    RI174b2098_868 , 
    RI173dbd18_1684 , 
    RI17393028_2039 , 
    RI174537f0_1329 , 
    RI19a97b68_2628 , 
    RI17478348_1150 , 
    RI19ac7958_2273 , 
    RI174c5d78_795 , 
    RI19ab6090_2408 , 
    RI174a16d0_949 , 
    RI1744c860_1363 , 
    RI19acbe40_2240 , 
    RI174ba900_830 , 
    RI19a9ce60_2591 , 
    RI17471070_1185 , 
    RI173d4d88_1718 , 
    RI1738c098_2073 , 
    RI173c9c40_1772 , 
    RI17412c78_1416 , 
    RI19ac0ba8_2325 , 
    RI174aef60_883 , 
    RI19a905c0_2680 , 
    RI17466288_1238 , 
    RI173d4a40_1719 , 
    RI173b7ec8_1859 , 
    RI17530500_616 , 
    RI1749cea0_971 , 
    RI19aba8c0_2377 , 
    RI173d5418_1716 , 
    RI1744cef0_1361 , 
    RI19a9aac0_2607 , 
    RI17471700_1183 , 
    RI19aca298_2254 , 
    RI174bb350_828 , 
    RI173df198_1668 , 
    RI19a9b1c8_2604 , 
    RI174720d8_1180 , 
    RI19aca9a0_2251 , 
    RI174bc2c8_825 , 
    RI173d5df0_1713 , 
    RI1738d100_2068 , 
    RI1744d8c8_1358 , 
    RI173a4710_1954 , 
    RI173deb08_1670 , 
    RI17395e18_2025 , 
    RI174565e0_1315 , 
    RI19ac4b68_2294 , 
    RI174ca5a8_781 , 
    RI19a94940_2650 , 
    RI1747b138_1136 , 
    RI173cfb68_1743 , 
    RI1744d238_1360 , 
    RI17461080_1263 , 
    RI173a08b8_1973 , 
    RI173e95a8_1618 , 
    RI19acf8d8_2214 , 
    RI1750b930_730 , 
    RI19aa0b50_2563 , 
    RI17485890_1085 , 
    RI173bdaa8_1831 , 
    RI17406798_1476 , 
    RI17334528_2186 , 
    RI174a2a80_943 , 
    RI19ab48a8_2419 , 
    RI173c8548_1779 , 
    RI1733efc8_2134 , 
    RI19a8f648_2687 , 
    RI17464b90_1245 , 
    RI19abff78_2332 , 
    RI174ad868_890 , 
    RI19a8f8a0_2686 , 
    RI17464ed8_1244 , 
    RI19ac0158_2331 , 
    RI174adbb0_889 , 
    RI173c8890_1778 , 
    RI173e6128_1634 , 
    RI1739d0f0_1990 , 
    RI1745dc00_1279 , 
    RI19aa3418_2543 , 
    RI17482410_1101 , 
    RI19a846f8_2763 , 
    RI175066b0_746 , 
    RI1744d580_1359 , 
    RI173d5760_1715 , 
    RI19aca4f0_2253 , 
    RI174bb878_827 , 
    RI19a9ad18_2606 , 
    RI17471a48_1182 , 
    RI19ac5108_2291 , 
    RI174caff8_779 , 
    RI173ea2c8_1614 , 
    RI173a15d8_1969 , 
    RI1746a0e0_1219 , 
    RI19aa1438_2558 , 
    RI174865b0_1081 , 
    RI19a82538_2778 , 
    RI1750cdd0_726 , 
    RI173ccd78_1757 , 
    RI173437f8_2112 , 
    RI17444bb0_1401 , 
    RI19a8d8c0_2700 , 
    RI174693c0_1223 , 
    RI17394a68_2031 , 
    RI19ac6620_2282 , 
    RI174c86b8_787 , 
    RI19a96740_2637 , 
    RI17479d88_1142 , 
    RI173a4a58_1953 , 
    RI173ed748_1598 , 
    RI1748c190_1053 , 
    RI19a9efa8_2577 , 
    RI17489a30_1065 , 
    RI19acda60_2227 , 
    RI17512050_710 , 
    RI173d0540_1740 , 
    RI17346c78_2096 , 
    RI17448030_1385 , 
    RI19a8aad0_2720 , 
    RI1746c840_1207 , 
    RI19abc4e0_2365 , 
    RI174b5518_852 , 
    RI19ac1670_2319 , 
    RI174acb48_894 , 
    RI173cfeb0_1742 , 
    RI173465e8_2098 , 
    RI174479a0_1387 , 
    RI19a8a878_2721 , 
    RI1746c1b0_1209 , 
    RI19abc378_2366 , 
    RI174b4e88_854 , 
    RI173fb9b0_1529 , 
    RI173a0570_1974 , 
    RI19a8b958_2714 , 
    RI17528418_641 , 
    RI19aa8080_2509 , 
    RI17497c98_996 , 
    RI173a7ed8_1937 , 
    RI173fafd8_1532 , 
    RI173b22e8_1887 , 
    RI1739de10_1986 , 
    RI19aa29c8_2548 , 
    RI175279c8_643 , 
    RI173fe458_1516 , 
    RI173b5420_1872 , 
    RI173bb9d8_1841 , 
    RI19a88a00_2734 , 
    RI1752c720_628 , 
    RI19aa7888_2513 , 
    RI1749a740_983 , 
    RI17389fc8_2083 , 
    RI19abb748_2371 , 
    RI174b7c78_840 , 
    RI19a89bd0_2726 , 
    RI1746efa0_1195 , 
    RI173efb60_1587 , 
    RI19accc50_2233 , 
    RI17515e30_698 , 
    RI17457990_1309 , 
    RI1740d098_1444 , 
    RI1733ae28_2154 , 
    RI174a96c8_910 , 
    RI19ab1ba8_2441 , 
    RI1740d728_1442 , 
    RI173bd760_1832 , 
    RI173341e0_2187 , 
    RI174a2738_944 , 
    RI19ab4740_2420 , 
    RI173fbcf8_1528 , 
    RI173b2cc0_1884 , 
    RI173a2988_1963 , 
    RI19aa81e8_2508 , 
    RI17497fe0_995 , 
    RI19a8d230_2703 , 
    RI17528940_640 , 
    RI173e98f0_1617 , 
    RI173a0c00_1972 , 
    RI17463498_1252 , 
    RI19acfb30_2213 , 
    RI1750be58_729 , 
    RI19aa0d30_2562 , 
    RI17485bd8_1084 , 
    RI173f15a0_1579 , 
    RI173a88b0_1934 , 
    RI174b2db8_864 , 
    RI19aa40c0_2537 , 
    RI17518770_690 , 
    RI19ab03c0_2452 , 
    RI1748d888_1046 , 
    RI173d2628_1730 , 
    RI173b7b80_1860 , 
    RI1752ffd8_617 , 
    RI1746e910_1197 , 
    RI174a5528_930 , 
    RI19accea8_2232 , 
    RI17516880_696 , 
    RI173f01f0_1585 , 
    RI173fd0a8_1522 , 
    RI173b4070_1878 , 
    RI19aa9430_2501 , 
    RI17499390_989 , 
    RI173d1908_1734 , 
    RI17359350_2090 , 
    RI174493e0_1379 , 
    RI19a89018_2731 , 
    RI1746dbf0_1201 , 
    RI17514990_702 , 
    RI19a9ed50_2578 , 
    RI174896e8_1066 , 
    RI173bc6f8_1837 , 
    RI17487960_1075 , 
    RI173df4e0_1667 , 
    RI173967f0_2022 , 
    RI17456fb8_1312 , 
    RI19a954f8_2645 , 
    RI1747bb10_1133 , 
    RI19ac52e8_2290 , 
    RI174cb520_778 , 
    RI174bdc90_820 , 
    RI1740ac80_1455 , 
    RI173c1f90_1810 , 
    RI17338a10_2165 , 
    RI174a72b0_921 , 
    RI19ab2b98_2434 , 
    RI19ac6e18_2278 , 
    RI174c3e88_801 , 
    RI173a8220_1936 , 
    RI173f0f10_1581 , 
    RI174ae588_886 , 
    RI19a887a8_2735 , 
    RI17517d20_692 , 
    RI19ab0000_2454 , 
    RI1748d1f8_1048 , 
    RI17457300_1311 , 
    RI19a8b4a8_2716 , 
    RI1746d560_1203 , 
    RI173d1278_1736 , 
    RI17358cc0_2092 , 
    RI17448d50_1381 , 
    RI19abef88_2341 , 
    RI174af5f0_881 , 
    RI1740ee20_1435 , 
    RI173d50d0_1717 , 
    RI1738c3e0_2072 , 
    RI1744cba8_1362 , 
    RI19acc020_2239 , 
    RI174bae28_829 , 
    RI19a9d1a8_2590 , 
    RI174713b8_1184 , 
    RI173d0f18_1737 , 
    RI17347650_2093 , 
    RI17448a08_1382 , 
    RI19abca80_2362 , 
    RI174b5ef0_849 , 
    RI19a8b250_2717 , 
    RI1746d218_1204 , 
    RI19acc5c0_2236 , 
    RI17514eb8_701 , 
    RI173e0890_1661 , 
    RI17397ba0_2016 , 
    RI174586b0_1305 , 
    RI19ac3920_2302 , 
    RI174cd410_772 , 
    RI19a936f8_2658 , 
    RI1747cec0_1127 , 
    RI17530f50_614 , 
    RI173f2950_1573 , 
    RI173a9c60_1928 , 
    RI174c1a70_808 , 
    RI19aae980_2464 , 
    RI1748ef80_1039 , 
    RI173f2c98_1572 , 
    RI19a97028_2633 , 
    RI17476c50_1157 , 
    RI173da968_1690 , 
    RI17391c78_2045 , 
    RI17452440_1335 , 
    RI19ac6ff8_2277 , 
    RI174c43b0_800 , 
    RI173da620_1691 , 
    RI17391930_2046 , 
    RI174520f8_1336 , 
    RI19ac8e70_2263 , 
    RI174c3960_802 , 
    RI19a99440_2617 , 
    RI17476908_1158 , 
    RI17405dc0_1479 , 
    RI173bd0d0_1834 , 
    RI17333b50_2189 , 
    RI17408ef8_1464 , 
    RI19ab6900_2405 , 
    RI174a20a8_946 , 
    RI19acc818_2235 , 
    RI175153e0_700 , 
    RI17397ee8_2015 , 
    RI173e0bd8_1660 , 
    RI174589f8_1304 , 
    RI19ac3b00_2301 , 
    RI174cd938_771 , 
    RI19a93950_2657 , 
    RI1747d208_1126 , 
    RI17410860_1427 , 
    RI17401f68_1498 , 
    RI173b9278_1853 , 
    RI175323f0_610 , 
    RI1749e250_965 , 
    RI19ab8f70_2388 , 
    RI173d9270_1697 , 
    RI173a1c68_1967 , 
    RI173f81e8_1546 , 
    RI173af4f8_1901 , 
    RI19aaad80_2489 , 
    RI17494818_1012 , 
    RI173cca30_1758 , 
    RI173434b0_2113 , 
    RI17415a68_1402 , 
    RI19a8d668_2701 , 
    RI17469078_1224 , 
    RI173d5aa8_1714 , 
    RI19aca748_2252 , 
    RI174bbda0_826 , 
    RI19a9af70_2605 , 
    RI17471d90_1181 , 
    RI173f2fe0_1571 , 
    RI173aa2f0_1926 , 
    RI19aaeea8_2462 , 
    RI1748f610_1037 , 
    RI19a9d9a0_2587 , 
    RI1748b470_1057 , 
    RI17499d68_986 , 
    RI19aabcf8_2483 , 
    RI17492400_1023 , 
    RI173a9fa8_1927 , 
    RI174c5328_797 , 
    RI19aaeb60_2463 , 
    RI1748f2c8_1038 , 
    RI173c74e0_1784 , 
    RI1733df60_2139 , 
    RI174101d0_1429 , 
    RI19ac1490_2320 , 
    RI174ac800_895 , 
    RI19a91100_2675 , 
    RI17463b28_1250 , 
    RI174025f8_1496 , 
    RI173b9908_1851 , 
    RI17532e40_608 , 
    RI19ab92b8_2387 , 
    RI1749e8e0_963 , 
    RI173dacb0_1689 , 
    RI17452788_1334 , 
    RI19a97208_2632 , 
    RI17476f98_1156 , 
    RI173ca2d0_1770 , 
    RI17340d50_2125 , 
    RI17413308_1414 , 
    RI173a95d0_1930 , 
    RI173c6130_1790 , 
    RI1733cbb0_2145 , 
    RI19a92bb8_2663 , 
    RI17462778_1256 , 
    RI19ac2f48_2307 , 
    RI174ab450_901 , 
    RI19aba398_2379 , 
    RI1749c810_973 , 
    RI173de130_1673 , 
    RI17395440_2028 , 
    RI17455c08_1318 , 
    RI19ac6bc0_2279 , 
    RI174c9630_784 , 
    RI19a96e48_2634 , 
    RI1747a760_1139 , 
    RI173d01f8_1741 , 
    RI17400528_1506 , 
    RI173b7838_1861 , 
    RI1752fab0_618 , 
    RI173ef188_1590 , 
    RI173a6498_1945 , 
    RI1749c180_975 , 
    RI173fcd60_1523 , 
    RI173b3d28_1879 , 
    RI173ade00_1908 , 
    RI19aa90e8_2502 , 
    RI17499048_990 , 
    RI173cd0c0_1756 , 
    RI17343b40_2111 , 
    RI19a8db18_2699 , 
    RI17469708_1222 , 
    RI19abe9e8_2344 , 
    RI174b23e0_867 , 
    RI19a82970_2776 , 
    RI1750d820_724 , 
    RI19aa17f8_2556 , 
    RI17486c40_1079 , 
    RI1739c088_1995 , 
    RI1745cb98_1284 , 
    RI19a86318_2751 , 
    RI17502e70_751 , 
    RI19aa4ed0_2530 , 
    RI174813a8_1106 , 
    RI173df828_1666 , 
    RI17396b38_2021 , 
    RI19a95750_2644 , 
    RI1747be58_1132 , 
    RI19ac5540_2289 , 
    RI174cba48_777 , 
    RI173ef4d0_1589 , 
    RI173a67e0_1944 , 
    RI1749e598_964 , 
    RI19a9dbf8_2586 , 
    RI1748b7b8_1056 , 
    RI173da2d8_1692 , 
    RI17451db0_1337 , 
    RI19ac8c18_2264 , 
    RI174c3438_803 , 
    RI19a991e8_2618 , 
    RI174765c0_1159 , 
    RI173d9c48_1694 , 
    RI17451720_1339 , 
    RI19ac8768_2266 , 
    RI174c29e8_805 , 
    RI19a98d38_2620 , 
    RI17475f30_1161 , 
    RI173f7180_1551 , 
    RI173ae490_1906 , 
    RI17334870_2185 , 
    RI19aacbf8_2477 , 
    RI174937b0_1017 , 
    RI19ab8778_2392 , 
    RI175217d0_662 , 
    RI173f5dd0_1557 , 
    RI17527ef0_642 , 
    RI19ab0c30_2448 , 
    RI1751f8e0_668 , 
    RI173ef818_1588 , 
    RI173a6b28_1943 , 
    RI19acc9f8_2234 , 
    RI17515908_699 , 
    RI19a9de50_2585 , 
    RI1748bb00_1055 , 
    RI173f3328_1570 , 
    RI173aa638_1925 , 
    RI174cc498_775 , 
    RI19aaf088_2461 , 
    RI1748f958_1036 , 
    RI19a23a38_2791 , 
    RI1751b5d8_681 , 
    RI173c7b70_1782 , 
    RI1733e5f0_2137 , 
    RI19ac1850_2318 , 
    RI174ace90_893 , 
    RI19a915b0_2673 , 
    RI174641b8_1248 , 
    RI173cbd10_1762 , 
    RI17342790_2117 , 
    RI17414d48_1406 , 
    RI19a8f3f0_2688 , 
    RI17468358_1228 , 
    RI19abfd98_2333 , 
    RI174b1030_873 , 
    RI174022b0_1497 , 
    RI17333178_2192 , 
    RI17456c70_1313 , 
    RI173eb9c0_1607 , 
    RI17477cb8_1152 , 
    RI19a9ff20_2569 , 
    RI17487ca8_1074 , 
    RI19aceac8_2220 , 
    RI1750f1e8_719 , 
    RI1740c378_1448 , 
    RI173cda98_1753 , 
    RI19ab11d0_2445 , 
    RI174a89a8_914 , 
    RI1733a108_2158 , 
    RI173a6150_1946 , 
    RI19acc3e0_2237 , 
    RI19a9d658_2588 , 
    RI1748b128_1058 , 
    RI173f0bc8_1582 , 
    RI174ac170_897 , 
    RI19a86de0_2746 , 
    RI175177f8_693 , 
    RI19aafcb8_2455 , 
    RI1748ceb0_1049 , 
    RI19a85760_2756 , 
    RI17500f80_757 , 
    RI17407b48_1470 , 
    RI19ab5640_2413 , 
    RI174a3e30_937 , 
    RI173bd418_1833 , 
    RI17333e98_2188 , 
    RI1740b310_1453 , 
    RI174a23f0_945 , 
    RI19ab6ae0_2404 , 
    RI19a8a530_2722 , 
    RI1746be68_1210 , 
    RI19abc198_2367 , 
    RI174b4b40_855 , 
    RI173462a0_2099 , 
    RI17447658_1388 , 
    RI173de478_1672 , 
    RI173ed0b8_1600 , 
    RI173a43c8_1955 , 
    RI19a9eaf8_2579 , 
    RI174893a0_1067 , 
    RI173c7828_1783 , 
    RI1733e2a8_2138 , 
    RI17410518_1428 , 
    RI19a91358_2674 , 
    RI17463e70_1249 , 
    RI1739c718_1993 , 
    RI1745d228_1282 , 
    RI19aa53f8_2528 , 
    RI17481a38_1104 , 
    RI19a86750_2749 , 
    RI175038c0_749 , 
    RI19ac46b8_2296 , 
    RI174c9b58_783 , 
    RI19a94b98_2649 , 
    RI1747b480_1135 , 
    RI17395788_2027 , 
    RI17455f50_1317 , 
    RI19a94490_2652 , 
    RI1747aaa8_1138 , 
    RI1748e5a8_1042 , 
    RI173c1900_1812 , 
    RI17338380_2167 , 
    RI174a6c20_923 , 
    RI19ab2670_2436 , 
    RI173dee50_1669 , 
    RI17396160_2024 , 
    RI17456928_1314 , 
    RI19ac4dc0_2293 , 
    RI174caad0_780 , 
    RI1739acd8_2001 , 
    RI173e39c8_1646 , 
    RI1745b7e8_1290 , 
    RI19aa44f8_2535 , 
    RI1747fff8_1112 , 
    RI173b8558_1857 , 
    RI17401248_1502 , 
    RI1749d530_969 , 
    RI19ab8430_2393 , 
    RI19a860c0_2752 , 
    RI17502948_752 , 
    RI19aa4cf0_2531 , 
    RI17481060_1107 , 
    RI173e4d78_1640 , 
    RI1739bd40_1996 , 
    RI1745c850_1285 , 
    RI173d6138_1712 , 
    RI1738d448_2067 , 
    RI1744dc10_1357 , 
    RI19a9b678_2602 , 
    RI17472420_1179 , 
    RI19acabf8_2250 , 
    RI174bc7f0_824 , 
    RI173ed400_1599 , 
    RI17489d78_1064 , 
    RI19acd808_2228 , 
    RI17511b28_711 , 
    RI19a952a0_2646 , 
    RI1747b7c8_1134 , 
    RI174a51e0_931 , 
    RI1740a938_1456 , 
    RI173c1c48_1811 , 
    RI173386c8_2166 , 
    RI17359008_2091 , 
    RI173fc6d0_1525 , 
    RI173b3698_1881 , 
    RI19a91c40_2670 , 
    RI175298b8_637 , 
    RI173e5de0_1635 , 
    RI1739cda8_1991 , 
    RI1745d8b8_1280 , 
    RI19a843b0_2764 , 
    RI17506188_747 , 
    RI173d15c0_1735 , 
    RI173fca18_1524 , 
    RI173b39e0_1880 , 
    RI173ab9e8_1919 , 
    RI19aa8da0_2504 , 
    RI17498d00_991 , 
    RI19a8b700_2715 , 
    RI1746d8a8_1202 , 
    RI173ea610_1613 , 
    RI173a1920_1968 , 
    RI1746c4f8_1208 , 
    RI19a82790_2777 , 
    RI1750d2f8_725 , 
    RI19aa1618_2557 , 
    RI174868f8_1080 , 
    RI17449098_1380 , 
    RI1754a6a8_69 , 
    RI1754a720_68 , 
    RI1754a630_70 , 
    RI1754bad0_26 , 
    RI1754a5b8_71 , 
    RI17538c00_591 , 
    RI19a25298_2780 , 
    RI1754b788_33 , 
    RI1754b878_31 , 
    RI1754c430_6 , 
    RI17536d88_596 , 
    RI1754b800_32 , 
    RI1754b530_38 , 
    RI19a822e0_2779 , 
    RI19ad0700_2208 , 
    RI1754bcb0_22 , 
    RI19a24ed8_2782 , 
    RI19a250b8_2781 , 
    RI1754be18_19 , 
    RI1754b350_42 , 
    RI1754c250_10 , 
    RI1754b1e8_45 , 
    RI19a24320_2787 , 
    RI19a24578_2786 , 
    RI1754b5a8_37 , 
    RI19ad21b8_2198 , 
    RI1754c160_12 , 
    RI1754a900_64 , 
    RI19a24c80_2783 , 
    RI1754bf08_17 , 
    RI1754ac48_57 , 
    RI1754bf80_16 , 
    RI1754bc38_23 , 
    RI19a240c8_2788 , 
    RI1754c070_14 , 
    RI1754b3c8_41 , 
    RI1754af18_51 , 
    RI1754b080_48 , 
    RI1754af90_50 , 
    RI1754bda0_20 , 
    RI1754aea0_52 , 
    RI1754b260_44 , 
    RI19ad0bb0_2206 , 
    RI19a24a28_2784 , 
    RI1754ae28_53 , 
    RI1754a888_65 , 
    RI1754bbc0_24 , 
    RI19ad0e08_2205 , 
    RI1754a810_66 , 
    RI1754b440_40 , 
    RI1754adb0_54 , 
    RI1754c3b8_7 , 
    RI19ad1060_2204 , 
    RI1754ba58_27 , 
    RI1754c340_8 , 
    RI1754aa68_61 , 
    RI1754ad38_55 , 
    RI19ad12b8_2203 , 
    RI1754be90_18 , 
    RI1754c2c8_9 , 
    RI1754c1d8_11 , 
    RI19a247d0_2785 , 
    RI1754b170_46 , 
    RI1754aae0_60 , 
    RI1754acc0_56 , 
    RI1754a978_63 , 
    RI19ad1588_2202 , 
    RI1754b620_36 , 
    RI1754bd28_21 , 
    RI1754b9e0_28 , 
    RI1754bb48_25 , 
    RI1754ab58_59 , 
    RI1754abd0_58 , 
    RI1754b2d8_43 , 
    RI1754c598_3 , 
    RI19ad1858_2201 , 
    RI1754b4b8_39 , 
    RI1754b0f8_47 , 
    RI1754c0e8_13 , 
    RI1754bff8_15 , 
    RI1754b698_35 , 
    RI19ad1c18_2200 , 
    RI1754c520_4 , 
    RI1754b968_29 , 
    RI19ad1ee8_2199 , 
    RI1754b008_49 , 
    RI1754c4a8_5 , 
    RI1754b710_34 , 
    RI1754a9f0_62 , 
    RI1754b8f0_30 , 
    RI19ad0958_2207 , 
    R_147ef_11ce6748 , 
    R_5f38_10569f58 , 
    R_13287_11ce6b08 , 
    R_c94b_102f7608 , 
    R_20a_1204ce78 , 
    R_12f29_10571bb8 , 
    R_13a43_13a1dec8 , 
    R_1474d_1056fbd8 , 
    R_14493_12657988 , 
    R_11fd1_11ce17e8 , 
    R_14705_1264d248 , 
    R_105_f8cc2b8 , 
    R_13cb9_11ce3c28 , 
    R_138ee_13309fa8 , 
    R_129dc_11543018 , 
    R_10bcf_11ce1ba8 , 
    R_13b6e_13a1e648 , 
    R_14840_13a13ec8 , 
    R_13482_10563838 , 
    R_12d08_12650088 , 
    R_10303_12b42dd8 , 
    R_1437c_1056ac78 , 
    R_87e9_1056cd98 , 
    R_a30d_13320588 , 
    R_144a2_133222e8 , 
    R_1236b_13a1c8e8 , 
    R_1396e_105627f8 , 
    R_9ba7_10567258 , 
    R_1f3_13797a68 , 
    R_11c_13796528 , 
    R_7a_1331e148 , 
    R_117c9_1264ba88 , 
    R_13b3f_1153ed38 , 
    R_11abc_1264c2a8 , 
    R_20d_137962a8 , 
    R_207_1265a548 , 
    R_14828_1207a118 , 
    R_148eb_105aa7d8 , 
    R_f3a4_10568bf8 , 
    R_1b6_13799d68 , 
    R_13429_1207f4d8 , 
    R_14506_1056e878 , 
    R_159_12b3d158 , 
    R_108_105aaeb8 , 
    R_102_13794cc8 , 
    R_b1_12053638 , 
    R_54_13309d28 , 
    R_145d8_12b3ae58 , 
    R_1278a_12083718 , 
    R_13640_11cdeae8 , 
    R_f706_11542578 , 
    R_dc82_1153ebf8 , 
    R_1491b_1265ef08 , 
    R_14a05_10569738 , 
    R_13fc5_102eac28 , 
    R_1405a_115415d8 , 
    R_136b3_126461c8 , 
    R_1a0_132f9c88 , 
    R_16f_1265bee8 , 
    R_1480d_105a9dd8 , 
    R_61_13304288 , 
    R_e082_13798fa8 , 
    R_10c7d_12082bd8 , 
    R_14793_1379e188 , 
    R_11ee1_102f4688 , 
    R_128ba_12b27758 , 
    R_70_120513d8 , 
    R_129f0_12049bd8 , 
    R_117e7_102f5588 , 
    R_fee6_13309e68 , 
    R_148f7_132f3ce8 , 
    R_1362d_11ce39a8 , 
    R_10693_126510c8 , 
    R_11998_12656808 , 
    R_143ec_11537df8 , 
    R_138e8_1264afe8 , 
    R_12650_12649b48 , 
    R_137a1_105b63f8 , 
    R_13afd_120772d8 , 
    R_1490c_1264a7c8 , 
    R_105e5_13306f88 , 
    R_12e2b_132fa868 , 
    R_144e7_12b38e78 , 
    R_143e4_11cddf08 , 
    R_1324a_1264c348 , 
    R_1215a_11542ed8 , 
    R_f685_11541678 , 
    R_149ba_102ecb68 , 
    R_135dc_12646088 , 
    R_1476c_11cd7928 , 
    R_146bd_11537998 , 
    R_1df_12b39378 , 
    R_13ee8_133069e8 , 
    R_130_1265ac28 , 
    R_65_12047c98 , 
    R_13d75_1330d6a8 , 
    R_13933_12081198 , 
    R_133b5_12648388 , 
    R_125a0_13311488 , 
    R_8c_1379a808 , 
    R_eadc_1207ead8 , 
    R_134c7_126487e8 , 
    R_11df5_1056e9b8 , 
    R_144d5_102f8aa8 , 
    R_12b2a_102eed28 , 
    R_143d2_11538898 , 
    R_1462c_102f8508 , 
    R_13269_11543658 , 
    R_f4_1331e0a8 , 
    R_d7_132fde28 , 
    R_238_1204ec78 , 
    R_21b_1265e508 , 
    R_12f3d_12b38b58 , 
    R_112f1_1153c858 , 
    R_f09_f8c93d8 , 
    R_1487c_11cd99a8 , 
    R_c08f_1207cb98 , 
    R_923a_13a1ab88 , 
    R_14042_102f2108 , 
    R_143e8_102f3b48 , 
    R_c2e7_13a19e68 , 
    R_c175_12045118 , 
    R_1450f_102f8b48 , 
    R_12b14_12077238 , 
    R_149e4_13a1c528 , 
    R_12a04_11ce2968 , 
    R_145ed_13a14e68 , 
    R_13884_13796488 , 
    R_13b0b_1330a688 , 
    R_b5a4_102f4868 , 
    R_14584_1056ec38 , 
    R_13cee_12653148 , 
    R_10bed_12080ab8 , 
    R_117f0_102ef4a8 , 
    R_10a2a_133048c8 , 
    R_1be_137995e8 , 
    R_151_12b448b8 , 
    R_ef06_10563c98 , 
    R_f9d4_1056b178 , 
    R_e88a_13a13a68 , 
    R_13c67_102f38c8 , 
    R_128eb_10568dd8 , 
    R_12eaf_f8c3118 , 
    R_204_12039778 , 
    R_14951_1265ebe8 , 
    R_149c3_11ce5348 , 
    R_1ad_12b28e78 , 
    R_13f99_102f0da8 , 
    R_162_12b25e58 , 
    R_12003_11cdf628 , 
    R_10b_11539478 , 
    R_ff_1203c6f8 , 
    R_1484f_1153ea18 , 
    R_a8_12b425b8 , 
    R_5d_13312068 , 
    R_210_12043bd8 , 
    R_13d84_102f4188 , 
    R_142e1_10568658 , 
    R_10f30_11cd9ae8 , 
    R_1293d_12b43d78 , 
    R_10b34_1056da18 , 
    R_11a07_102eb4e8 , 
    R_145b1_12082db8 , 
    R_12c96_13a190a8 , 
    R_d3b0_10565958 , 
    R_13f2c_102f4b88 , 
    R_fb8a_13a18608 , 
    R_130d5_13319c88 , 
    R_13f89_102f36e8 , 
    R_146ff_13a1a4a8 , 
    R_10ccb_1264f868 , 
    R_124c3_1056f138 , 
    R_10786_102f2568 , 
    R_12a16_10568e78 , 
    R_10726_102ef408 , 
    R_137d3_12656da8 , 
    R_13863_11cddb48 , 
    R_14993_102f27e8 , 
    R_bab1_1264a2c8 , 
    R_1451e_10565818 , 
    R_12a46_126515c8 , 
    R_e7da_102f3508 , 
    R_12756_13a1f0e8 , 
    R_c4_13797ba8 , 
    R_128da_1207ec18 , 
    R_c282_12076838 , 
    R_1272e_1056cbb8 , 
    R_14a5f_120797b8 , 
    R_14448_12663648 , 
    R_c2_12048058 , 
    R_1372d_11ce2aa8 , 
    R_f878_1207c7d8 , 
    R_13a76_13797888 , 
    R_13a17_13796b68 , 
    R_1cb_12044ad8 , 
    R_14462_12b3f8b8 , 
    R_6021_1379bd48 , 
    R_144_13795128 , 
    R_1383e_105671b8 , 
    R_147ab_1056a6d8 , 
    R_c6_1330e0a8 , 
    R_249_12654368 , 
    R_1305a_13796ca8 , 
    R_12e4b_13307348 , 
    R_14a38_137a1e28 , 
    R_d1de_11cd9ea8 , 
    R_138e2_11cd83c8 , 
    R_13e62_1056dab8 , 
    R_114a7_1331d748 , 
    R_12f53_13319648 , 
    R_f8a4_11543a18 , 
    R_11ec3_13a157c8 , 
    R_12c06_11cdac68 , 
    R_12be8_12649788 , 
    R_136c6_11cdc6a8 , 
    R_1482e_13a1a228 , 
    R_10ba7_115431f8 , 
    R_89f2_11545098 , 
    R_11953_1153c538 , 
    R_9e64_11ce48a8 , 
    R_e77d_11ce3ea8 , 
    R_1091c_13a1a2c8 , 
    R_114ec_12650628 , 
    R_1286a_11cdcd88 , 
    R_10d6d_1265db08 , 
    R_1228f_1331f0e8 , 
    R_1c5_126590a8 , 
    R_14490_132f7d48 , 
    R_1a1_1264a408 , 
    R_976e_12056398 , 
    R_6845_12648ec8 , 
    R_16e_1379a3a8 , 
    R_14a_12657528 , 
    R_12718_10566fd8 , 
    R_145c9_12075438 , 
    R_c0_132fa5e8 , 
    R_9c_12655f48 , 
    R_d230_102edec8 , 
    R_69_12658888 , 
    R_13097_11ce5b68 , 
    R_11051_1264a5e8 , 
    R_145f0_11536818 , 
    R_13ccd_132f9288 , 
    R_e0_12661ac8 , 
    R_22f_1331df68 , 
    R_12a2a_11cd9f48 , 
    R_10a54_11540458 , 
    R_d027_13795628 , 
    R_144d2_105677f8 , 
    R_14638_11cd9228 , 
    R_1454b_10568338 , 
    R_147fe_1265bb28 , 
    R_e861_12650448 , 
    R_c03c_137931e8 , 
    R_13574_102f97c8 , 
    R_10e6d_102ec0c8 , 
    R_c8_1331c348 , 
    R_247_12b3bad8 , 
    R_77_126636e8 , 
    R_13a50_1056bb78 , 
    R_129a5_11543798 , 
    R_ef35_102f6d48 , 
    R_1028c_137951c8 , 
    R_1348b_12051838 , 
    R_11f8b_11cdc428 , 
    R_1452d_f8c5878 , 
    R_12a3b_12650308 , 
    R_13fd5_12079d58 , 
    R_dd89_13302de8 , 
    R_13dcc_102f7ec8 , 
    R_14822_102f5768 , 
    R_baf1_12084e38 , 
    R_1315c_11ce75a8 , 
    R_df0e_12654d68 , 
    R_efea_11cdc248 , 
    R_fe90_13a14a08 , 
    R_1453c_102ec208 , 
    R_aaa7_102edba8 , 
    R_13c4e_13a1c988 , 
    R_f758_13a13d88 , 
    R_1485e_12b38f18 , 
    R_ece9_1264c488 , 
    R_14a35_12037f18 , 
    R_1190c_102ecfc8 , 
    R_12810_12650d08 , 
    R_f016_12044df8 , 
    R_1494e_13a14f08 , 
    R_14344_1264eaa8 , 
    R_10e_1265af48 , 
    R_13f62_12075758 , 
    R_fc_133201c8 , 
    R_1378e_11cdd8c8 , 
    R_147eb_120847f8 , 
    R_13331_13308ec8 , 
    R_213_12654f48 , 
    R_146ae_1265dc48 , 
    R_201_1153b138 , 
    R_11d47_f8cc0d8 , 
    R_c820_13a19328 , 
    R_edbe_132fbd08 , 
    R_be_132f4148 , 
    R_a1_12043c78 , 
    R_131b9_102f29c8 , 
    R_12eb9_1153f738 , 
    R_146e1_1153fb98 , 
    R_1487f_13a173e8 , 
    R_13fb4_11544af8 , 
    R_1446b_10568798 , 
    R_ef60_1264cf28 , 
    R_1463b_1207bd38 , 
    R_13166_1153aff8 , 
    R_10a4b_10565bd8 , 
    R_14599_12080c98 , 
    R_10b18_12080018 , 
    R_7254_12055078 , 
    R_db04_1207b3d8 , 
    R_149f9_10570cb8 , 
    R_14a4a_1265d608 , 
    R_14796_1264b808 , 
    R_120d3_1379f3a8 , 
    R_119cb_102f2068 , 
    R_12acb_10565458 , 
    R_145b4_12083358 , 
    R_11ae9_12651528 , 
    R_13af6_f8ce6f8 , 
    R_13451_102f0128 , 
    R_ef8c_1204e098 , 
    R_ca_12b3e058 , 
    R_245_f8c5ff8 , 
    R_af_12b2a8b8 , 
    R_10e57_11544eb8 , 
    R_b243_f8c5698 , 
    R_13633_13a13248 , 
    R_11c97_10562078 , 
    R_13838_102f5e48 , 
    R_efb7_13a1bc68 , 
    R_d4db_10566038 , 
    R_10bc8_11ce66a8 , 
    R_c9c0_102eee68 , 
    R_13608_10563798 , 
    R_8f_12b299b8 , 
    R_59_133089c8 , 
    R_134f1_102ebf88 , 
    R_10499_1331e828 , 
    R_14424_102f8f08 , 
    R_1d6_133209e8 , 
    R_ebe2_13a18568 , 
    R_139_12b44ef8 , 
    R_97_13792c48 , 
    R_144ed_105660d8 , 
    R_120c8_11541d58 , 
    R_11736_11cde408 , 
    R_149a8_13317528 , 
    R_1450c_1056eff8 , 
    R_147d9_120828b8 , 
    R_11ea5_1264a9a8 , 
    R_11425_1207c918 , 
    R_d53e_1207c2d8 , 
    R_14787_12b352b8 , 
    R_13cf3_10571078 , 
    R_13f36_1330ebe8 , 
    R_d00d_102ee968 , 
    R_a1e6_11cde368 , 
    R_13f77_13a19648 , 
    R_118_132f5f48 , 
    R_13688_120832b8 , 
    R_1f7_105a9978 , 
    R_f630_1056b858 , 
    R_136a1_1153fa58 , 
    R_1b7_126577a8 , 
    R_158_12b27938 , 
    R_ec_1330a868 , 
    R_223_f8c32f8 , 
    R_133bf_11543338 , 
    R_f2a8_102f47c8 , 
    R_e112_12076e78 , 
    R_12b72_1056c6b8 , 
    R_2f00_102f3d28 , 
    R_14819_1331de28 , 
    R_e809_13313c48 , 
    R_14358_11cd8788 , 
    R_1473e_11543b58 , 
    R_139c7_102ed1a8 , 
    R_13d65_12036a78 , 
    R_12c10_102ea548 , 
    R_13870_11ce5e88 , 
    R_dede_13a16448 , 
    R_12c49_12b27438 , 
    R_1192b_12645e08 , 
    R_bd66_126533c8 , 
    R_13fa2_1379f6c8 , 
    R_13407_1056df18 , 
    R_118b0_1204acb8 , 
    R_13c3e_126496e8 , 
    R_1438a_11cda268 , 
    R_11e51_102fa268 , 
    R_102b9_132f6588 , 
    R_d9_1330dec8 , 
    R_bc_13799c28 , 
    R_236_13795f88 , 
    R_ffee_1264d568 , 
    R_10ea9_102f8788 , 
    R_14852_13a154a8 , 
    R_e696_11cdce28 , 
    R_1ae_1203c3d8 , 
    R_1457e_133027e8 , 
    R_161_12656c68 , 
    R_127_12b3cc58 , 
    R_ea26_1265a4a8 , 
    R_1e8_11539298 , 
    R_139e4_102f59e8 , 
    R_1477b_1204f218 , 
    R_1459c_12056a78 , 
    R_1336e_11545138 , 
    R_108cd_102f7ce8 , 
    R_13b4f_13305c28 , 
    R_1a2_12b423d8 , 
    R_16d_12664c28 , 
    R_14656_11ce6ce8 , 
    R_827e_1207e998 , 
    R_11ab0_1204a358 , 
    R_144ab_12b39af8 , 
    R_144c3_12080338 , 
    R_12794_102f5b28 , 
    R_13149_102f7888 , 
    R_144e4_12b28838 , 
    R_13e_12660da8 , 
    R_123_1330d888 , 
    R_e7_137956c8 , 
    R_cc_12038918 , 
    R_137c7_102f79c8 , 
    R_243_13796d48 , 
    R_13795_13795588 , 
    R_228_10570c18 , 
    R_13f01_1056e2d8 , 
    R_13d8e_11cd77e8 , 
    R_1ec_12039ef8 , 
    R_f175_13a17ca8 , 
    R_1d1_126540e8 , 
    R_14409_12b434b8 , 
    R_138b2_102f06c8 , 
    R_14653_1207e0d8 , 
    R_13044_102f7a68 , 
    R_13133_13a1ae08 , 
    R_10b8f_1265ad68 , 
    R_12e35_12b3b858 , 
    R_12df0_12050bb8 , 
    R_fc88_1207be78 , 
    R_13804_102ef548 , 
    R_13b68_137a1ba8 , 
    R_134_13312b68 , 
    R_14990_1331ae08 , 
    R_1db_12043db8 , 
    R_ccdc_102f6488 , 
    R_1494b_11ce61a8 , 
    R_12c39_10562ed8 , 
    R_131c2_11ce4b28 , 
    R_12d97_126626a8 , 
    R_12d59_12b26b78 , 
    R_1352d_13315188 , 
    R_12c4f_13321d48 , 
    R_1343e_10562d98 , 
    R_1345b_102fa088 , 
    R_1167d_115410d8 , 
    R_14008_1264dec8 , 
    R_11bc8_11544e18 , 
    R_13c9a_1207e178 , 
    R_148be_12b27f78 , 
    R_14360_105ad078 , 
    R_13aa3_12078138 , 
    R_116da_13a1a7c8 , 
    R_14732_102f5448 , 
    R_cec6_132f3608 , 
    R_133dc_13a1ea08 , 
    R_14942_f8c5058 , 
    R_13a0f_10563018 , 
    R_bd10_f8ce978 , 
    R_12da1_12647528 , 
    R_12af5_12052418 , 
    R_13cf9_13a1c0c8 , 
    R_13658_12646628 , 
    R_149bd_1204adf8 , 
    R_13233_11cde908 , 
    R_12585_1207a898 , 
    R_118e9_10564a58 , 
    R_1359a_13a18928 , 
    R_12451_13a1d568 , 
    R_dcbb_1265bf88 , 
    R_f424_13a1b948 , 
    R_1226a_11cdef48 , 
    R_14641_13a12d48 , 
    R_1257c_11ce4448 , 
    R_e309_120806f8 , 
    R_11ccc_13314be8 , 
    R_146c0_13a15908 , 
    R_14843_13a196e8 , 
    R_11d00_1207f9d8 , 
    R_14a1d_13a14c88 , 
    R_13d54_11ce00c8 , 
    R_135b5_132fdd88 , 
    R_d40b_10569058 , 
    R_145f9_102ee148 , 
    R_14882_1056d838 , 
    R_101a4_f8c2ad8 , 
    R_13abf_13a15188 , 
    R_eab3_126509e8 , 
    R_8296_13322608 , 
    R_6d_12036618 , 
    R_50_12b3c118 , 
    R_11b19_102ee508 , 
    R_de1d_13a193c8 , 
    R_14477_11cdcc48 , 
    R_1195d_12038198 , 
    R_14527_102eb6c8 , 
    R_be8c_126504e8 , 
    R_11e87_12b3c398 , 
    R_14a02_13309aa8 , 
    R_12b_1203e6d8 , 
    R_f1_13799ea8 , 
    R_21e_126608a8 , 
    R_1e4_12b28338 , 
    R_115ff_13304148 , 
    R_10d8e_1264cfc8 , 
    R_11500_12083c18 , 
    R_c4bc_137945e8 , 
    R_1465c_10568f18 , 
    R_133e6_11cd9048 , 
    R_7c4f_11ce4a88 , 
    R_11f78_12b2c118 , 
    R_1013a_132f59a8 , 
    R_149e1_105b62b8 , 
    R_150_1330cac8 , 
    R_111_12b3e238 , 
    R_f9_1204ba78 , 
    R_ba_1331bc68 , 
    R_4b_1264c028 , 
    R_216_1204a038 , 
    R_13733_f8d0098 , 
    R_1fe_120539f8 , 
    R_146de_12648748 , 
    R_1bf_1265cd48 , 
    R_74_1331da68 , 
    R_f5c3_1264d108 , 
    R_f1f7_120367f8 , 
    R_e338_13301ac8 , 
    R_1486d_1056e558 , 
    R_13e2d_12047fb8 , 
    R_12344_137a0de8 , 
    R_14729_10570178 , 
    R_13364_105717f8 , 
    R_11160_1153e298 , 
    R_10a01_11cde228 , 
    R_13c6f_12041658 , 
    R_148c4_10568978 , 
    R_11c81_132f7348 , 
    R_10ec5_11cdb028 , 
    R_14441_12659008 , 
    R_cbab_105a9a18 , 
    R_1238a_126482e8 , 
    R_a6_12660448 , 
    R_12b36_11ce6428 , 
    R_dc46_10566498 , 
    R_11f_137936e8 , 
    R_ce_12055fd8 , 
    R_241_132fd748 , 
    R_147f8_1207ccd8 , 
    R_1f0_13798a08 , 
    R_1467d_1056bcb8 , 
    R_14668_11546178 , 
    R_132cc_1153edd8 , 
    R_136ba_11ce37c8 , 
    R_12c23_102f1d48 , 
    R_106be_1264edc8 , 
    R_11bde_10564878 , 
    R_11a1a_11cd9a48 , 
    R_9548_11ce6ba8 , 
    R_f451_11542438 , 
    R_119b7_105663f8 , 
    R_142e5_102f2388 , 
    R_147e4_13a19dc8 , 
    R_d862_12661348 , 
    R_d940_13a19d28 , 
    R_eb8c_13a19288 , 
    R_1175e_11cda088 , 
    R_146f9_11ce4768 , 
    R_14551_102eae08 , 
    R_14578_12b3a6d8 , 
    R_1467a_13a13568 , 
    R_1130e_1056bfd8 , 
    R_1493f_1056d3d8 , 
    R_14948_102f76a8 , 
    R_10230_1153d1b8 , 
    R_f4d1_13a17848 , 
    R_14772_11cda8a8 , 
    R_1466e_1203e138 , 
    R_14999_120382d8 , 
    R_9d72_102f18e8 , 
    R_eeaf_10566f38 , 
    R_13083_12b3ff98 , 
    R_e288_11541fd8 , 
    R_13969_102ea408 , 
    R_13825_1264d928 , 
    R_134a8_13a13c48 , 
    R_fcde_115390b8 , 
    R_14566_102f6988 , 
    R_f5eb_11544558 , 
    R_12318_102ec348 , 
    R_d2c9_11cd9408 , 
    R_16c_132f7ca8 , 
    R_d894_1056f778 , 
    R_12323_102ec8e8 , 
    R_1a3_13303108 , 
    R_118ba_13307ac8 , 
    R_12704_10562938 , 
    R_148c7_1264d888 , 
    R_148bb_12661d48 , 
    R_1221a_13a1d248 , 
    R_135b0_12651348 , 
    R_1470e_10562898 , 
    R_efa_1207d1d8 , 
    R_ce1e_102f95e8 , 
    R_126e3_105b5c78 , 
    R_14026_102ecd48 , 
    R_11e36_102ed608 , 
    R_11515_12039318 , 
    R_108e3_1056dd38 , 
    R_128f4_1207aa78 , 
    R_147ae_1207ce18 , 
    R_12235_12650e48 , 
    R_12183_12052eb8 , 
    R_14647_102f04e8 , 
    R_13aef_11cdd968 , 
    R_1249f_102f9368 , 
    R_f34d_13a18ec8 , 
    R_12c3f_f8cfd78 , 
    R_13d5d_1153d4d8 , 
    R_12126_102ef228 , 
    R_ad_12b3b358 , 
    R_92_13312d48 , 
    R_113db_f8cb4f8 , 
    R_10d98_f8c6318 , 
    R_1481f_1264dce8 , 
    R_ad98_102f3aa8 , 
    R_55_132f50e8 , 
    R_102d5_f8ced38 , 
    R_144ae_11545ef8 , 
    R_a3e0_12655308 , 
    R_5dbf_13a15f48 , 
    R_e2_1203f858 , 
    R_22d_1379de68 , 
    R_135c4_105b5bd8 , 
    R_13cff_13a16308 , 
    R_12692_102eb8a8 , 
    R_13375_13794a48 , 
    R_12f6a_10562438 , 
    R_128c4_102ea5e8 , 
    R_122f0_12650f88 , 
    R_14855_12056f78 , 
    R_14885_13795a88 , 
    R_bb92_11ce0ca8 , 
    R_8b04_1265cf28 , 
    R_e71c_115426b8 , 
    R_14a23_120545d8 , 
    R_149_1330f408 , 
    R_b8_13305048 , 
    R_1c6_1379cce8 , 
    R_e13d_102eb448 , 
    R_14617_11ce2f08 , 
    R_13557_11545778 , 
    R_148cd_12082c78 , 
    R_11768_1264ffe8 , 
    R_12503_11cdd008 , 
    R_1239d_1330d1a8 , 
    R_1448c_105662b8 , 
    R_160_f8c0d78 , 
    R_143_13795e48 , 
    R_1252c_102f1208 , 
    R_1cc_f8cc858 , 
    R_149de_11cde7c8 , 
    R_1af_12b40678 , 
    R_a28f_11ce5708 , 
    R_f7ae_11ce57a8 , 
    R_1243d_10571118 , 
    R_d0df_126478e8 , 
    R_1498d_1153fe18 , 
    R_10350_11cda6c8 , 
    R_103a6_10569878 , 
    R_128b0_1056c118 , 
    R_14936_10561e98 , 
    R_10d1b_11cd7748 , 
    R_ed92_102eea08 , 
    R_145d2_11cdb208 , 
    R_109f6_1153ca38 , 
    R_cc46_1207b298 , 
    R_11006_126501c8 , 
    R_188_1265c348 , 
    R_187_12b25d18 , 
    R_12f_1379dbe8 , 
    R_db_12663f08 , 
    R_84_12652ce8 , 
    R_81_12042a58 , 
    R_234_12b43af8 , 
    R_1e0_133037e8 , 
    R_13ed7_1207ad98 , 
    R_189_f8c6458 , 
    R_186_126553a8 , 
    R_157_132f7a28 , 
    R_d0_105aa238 , 
    R_23f_13307848 , 
    R_11399_12b3c1b8 , 
    R_1b8_11537358 , 
    R_f82c_f8cdc58 , 
    R_d9ca_10562bb8 , 
    R_145f6_f8c3398 , 
    R_1449c_11ce71e8 , 
    R_13850_13a1fe08 , 
    R_135e3_13306da8 , 
    R_ec0b_132fa368 , 
    R_147e0_13a12fc8 , 
    R_13add_132ff728 , 
    R_f65b_12084578 , 
    R_10cb4_11cdf9e8 , 
    R_18a_133173e8 , 
    R_185_12042cd8 , 
    R_134d0_12651028 , 
    R_144f3_102f3fa8 , 
    R_12dd1_f8c52d8 , 
    R_135a9_10567938 , 
    R_11b39_102ec988 , 
    R_1386a_102ebda8 , 
    R_14747_12042b98 , 
    R_148d0_137a0a28 , 
    R_11f4d_137986e8 , 
    R_13d05_12081378 , 
    R_f56e_102f2608 , 
    R_62_12b26498 , 
    R_10e0b_1056abd8 , 
    R_ba73_1264c8e8 , 
    R_14888_12653288 , 
    R_fc34_1379c428 , 
    R_18b_12663fa8 , 
    R_184_1153acd8 , 
    R_119d5_1331dc48 , 
    R_122b5_13305688 , 
    R_e051_12649f08 , 
    R_ca0a_10567438 , 
    R_10a84_115427f8 , 
    R_668e_10563f18 , 
    R_14539_102f7108 , 
    R_c3d6_11cdb7a8 , 
    R_11703_132fa728 , 
    R_1472f_105708f8 , 
    R_1307a_11cdc1a8 , 
    R_fdae_1153d258 , 
    R_13ac5_102ee3c8 , 
    R_120bd_1153ff58 , 
    R_13f6e_12649dc8 , 
    R_1177b_1207fbb8 , 
    R_f804_1379efe8 , 
    R_111d5_13a17c08 , 
    R_14750_13304008 , 
    R_137d9_12055e98 , 
    R_87_132ffa48 , 
    R_7e_137949a8 , 
    R_f140_1056f598 , 
    R_d43f_12079678 , 
    R_11900_1056f6d8 , 
    R_18c_12660e48 , 
    R_c969_1330f9a8 , 
    R_183_126587e8 , 
    R_11093_102f60c8 , 
    R_f31e_120770f8 , 
    R_f06_1265f728 , 
    R_d5cf_102f5128 , 
    R_10874_12037838 , 
    R_11324_13a1f228 , 
    R_13621_120823b8 , 
    R_120dd_f8cdcf8 , 
    R_148d3_12049a98 , 
    R_13e42_12648888 , 
    R_144c0_12078db8 , 
    R_12978_13316d08 , 
    R_11b5e_13a1b088 , 
    R_13025_13a1ef08 , 
    R_e615_12084bb8 , 
    R_149b7_102ea4a8 , 
    R_1497e_1207ef38 , 
    R_11fee_12b2a3b8 , 
    R_11b_12b43198 , 
    R_5e_126647c8 , 
    R_1f4_1265d108 , 
    R_1445f_13792888 , 
    R_13981_13798aa8 , 
    R_14569_11cdbfc8 , 
    R_114_12b3e4b8 , 
    R_f6_12664188 , 
    R_9f_12054d58 , 
    R_66_13308068 , 
    R_219_1203c338 , 
    R_132a5_12654868 , 
    R_f9aa_11cdd5a8 , 
    R_1fb_126610c8 , 
    R_1a4_13798648 , 
    R_16b_1331a2c8 , 
    R_9a_12658568 , 
    R_13c54_102f6e88 , 
    R_14933_1207e5d8 , 
    R_a6b7_1264b588 , 
    R_10fad_13a15548 , 
    R_18d_13321a28 , 
    R_182_13315cc8 , 
    R_14a58_102f65c8 , 
    R_c8f6_132f4a08 , 
    R_1458d_13a17ac8 , 
    R_126d9_11545598 , 
    R_10942_102f85a8 , 
    R_14a32_12654ea8 , 
    R_b7bc_12b28798 , 
    R_1389f_11cda3a8 , 
    R_14602_102ed7e8 , 
    R_100bf_1330b9e8 , 
    R_112eb_115386b8 , 
    R_146d5_105b59f8 , 
    R_1206a_1207c878 , 
    R_e2de_1264ce88 , 
    R_13b3a_11cddaa8 , 
    R_13739_10563bf8 , 
    R_148d6_11cd86e8 , 
    R_1319d_11544918 , 
    R_12f7f_12077eb8 , 
    R_1242c_f8cda78 , 
    R_14483_12054fd8 , 
    R_14456_102ea728 , 
    R_6b42_120790d8 , 
    R_1186d_f8cbb38 , 
    R_147d3_12648e28 , 
    R_11add_1056c4d8 , 
    R_13c18_1264df68 , 
    R_13e19_132f7c08 , 
    R_b6_1265e148 , 
    R_13bb8_1265edc8 , 
    R_146a8_12050118 , 
    R_18e_12043ef8 , 
    R_181_12647a28 , 
    R_b677_12083178 , 
    R_1176f_1379f8a8 , 
    R_11d7b_102f2d88 , 
    R_145bd_1207cff8 , 
    R_13bae_105700d8 , 
    R_10fed_1330ad68 , 
    R_1479f_11cde4a8 , 
    R_71_1265e8c8 , 
    R_3ca5_102eebe8 , 
    R_14769_1056b718 , 
    R_139ba_11ce35e8 , 
    R_ccf5_13a128e8 , 
    R_13964_1207def8 , 
    R_13920_133128e8 , 
    R_13b74_11cd8dc8 , 
    R_13e6d_11cd90e8 , 
    R_13ae8_11545db8 , 
    R_e946_13796668 , 
    R_12db3_10562b18 , 
    R_7b5f_1264bc68 , 
    R_139f5_132fc348 , 
    R_cd6e_10562a78 , 
    R_13626_12077cd8 , 
    R_148dc_102f3c88 , 
    R_11db0_13302748 , 
    R_1470b_115413f8 , 
    R_fd8e_120835d8 , 
    R_142aa_102f2a68 , 
    R_1267b_1056b538 , 
    R_10df7_1264ae08 , 
    R_b753_102ebe48 , 
    R_14a47_102eeb48 , 
    R_12f94_1379c068 , 
    R_f3d0_1264e3c8 , 
    R_13cd6_10565638 , 
    R_123b1_12b3e378 , 
    R_144cf_f8c96f8 , 
    R_13d0c_102f6168 , 
    R_13c61_12081d78 , 
    R_134f6_11ce6608 , 
    R_112c2_12b294b8 , 
    R_11922_1056c898 , 
    R_11971_1207dbd8 , 
    R_138_1265b308 , 
    R_d2_12654c28 , 
    R_23d_12656088 , 
    R_8a_1379cba8 , 
    R_38ad_12048418 , 
    R_7b_12651de8 , 
    R_13889_10564918 , 
    R_13188_12079c18 , 
    R_13b8c_13a15728 , 
    R_947f_1056eaf8 , 
    R_1d7_12649648 , 
    R_149db_102f1668 , 
    R_ac1d_120826d8 , 
    R_13a06_105668f8 , 
    R_18f_132fc988 , 
    R_180_1265fea8 , 
    R_10e36_11ce6d88 , 
    R_136a7_12035cb8 , 
    R_148df_13a1d608 , 
    R_1380f_12080838 , 
    R_1485b_1265a688 , 
    R_14930_102f1a28 , 
    R_10044_102f1c08 , 
    R_d2a3_1207bbf8 , 
    R_1c0_1203c0b8 , 
    R_14f_12b25778 , 
    R_8472_126654e8 , 
    R_1483d_11ce0d48 , 
    R_12b67_11cdf3a8 , 
    R_11346_12655448 , 
    R_13893_12084d98 , 
    R_103f0_1207ecb8 , 
    R_1308d_1379eea8 , 
    R_f8ce_102f10c8 , 
    R_13f82_11543978 , 
    R_12359_133022e8 , 
    R_12cd3_13a1f728 , 
    R_13546_1153efb8 , 
    R_143b6_115408b8 , 
    R_148e5_10568518 , 
    R_10a79_11545278 , 
    R_1368d_102f3be8 , 
    R_14002_12047518 , 
    R_febc_1207caf8 , 
    R_14987_10571d98 , 
    R_14894_126569e8 , 
    R_13e23_102f1708 , 
    R_12304_10569e18 , 
    R_12daa_f8cc218 , 
    R_1289e_13316128 , 
    R_146ea_132fd6a8 , 
    R_104_12b414d8 , 
    R_e9_12055a78 , 
    R_226_12652568 , 
    R_20b_12656bc8 , 
    R_1484c_1056c078 , 
    R_149fc_12077a58 , 
    R_143f0_120442b8 , 
    R_107_1203f538 , 
    R_208_12b260d8 , 
    R_1d2_1203ce78 , 
    R_1442a_102f6668 , 
    R_13d_1379c568 , 
    R_134be_13a19148 , 
    R_145cf_13304328 , 
    R_12fa4_1153e0b8 , 
    R_1053d_12079858 , 
    R_ee_f8c86b8 , 
    R_221_12652888 , 
    R_13eb5_132f7ac8 , 
    R_190_133178e8 , 
    R_17f_115396f8 , 
    R_137af_11ce6e28 , 
    R_1455a_102ed748 , 
    R_10db8_102f74c8 , 
    R_ab_1264cde8 , 
    R_1187e_12077698 , 
    R_5a_126653a8 , 
    R_7e57_13a1a188 , 
    R_146ed_1153a238 , 
    R_1b0_12b29918 , 
    R_15f_1265f188 , 
    R_138b8_1264a368 , 
    R_13bd6_102f9188 , 
    R_14a17_102f0ee8 , 
    R_143a6_133121a8 , 
    R_11f57_12649328 , 
    R_14972_13302608 , 
    R_10701_1207f1b8 , 
    R_14503_1203e3b8 , 
    R_a4_12b36e98 , 
    R_6a_12b40178 , 
    R_aeba_105624d8 , 
    R_1379b_11ce6ec8 , 
    R_134e2_13a1e3c8 , 
    R_10973_12663008 , 
    R_11c66_102f7ba8 , 
    R_1325f_126468a8 , 
    R_1327d_10570d58 , 
    R_13417_102f3968 , 
    R_101_1264f048 , 
    R_95_133017a8 , 
    R_20e_1265e788 , 
    R_13c59_105b5638 , 
    R_13ca1_12652f68 , 
    R_1481c_11cdb988 , 
    R_14611_11545458 , 
    R_12fae_102f7388 , 
    R_1469f_1207d138 , 
    R_142dd_13314828 , 
    R_1279d_12079fd8 , 
    R_12646_1056b2b8 , 
    R_11486_102ee788 , 
    R_13389_1207fb18 , 
    R_1492d_11ce64c8 , 
    R_12d46_12648928 , 
    R_145b7_12b3d5b8 , 
    R_b211_12048c38 , 
    R_143aa_13795c68 , 
    R_1110c_11cdc928 , 
    R_1a5_12b3c618 , 
    R_16a_137a1248 , 
    R_df67_1207b8d8 , 
    R_124f6_1264f2c8 , 
    R_12b54_102f2248 , 
    R_d7dc_13a17de8 , 
    R_1247b_11ce4808 , 
    R_149ea_11540598 , 
    R_10a_12b30678 , 
    R_13c77_13a1cc08 , 
    R_205_12653dc8 , 
    R_14753_1264efa8 , 
    R_191_12043d18 , 
    R_17e_132f8568 , 
    R_11c4b_13a15c28 , 
    R_13208_11542758 , 
    R_e0ad_133021a8 , 
    R_11a3f_12b3e9b8 , 
    R_1230e_f8cb598 , 
    R_eee_1056adb8 , 
    R_14444_12648108 , 
    R_1dc_11538d98 , 
    R_12b7a_1264f188 , 
    R_133_13313888 , 
    R_147b1_105b5a98 , 
    R_f116_11ce1068 , 
    R_13a5c_1379a268 , 
    R_14340_12078458 , 
    R_e522_1330ed28 , 
    R_146f0_1153da78 , 
    R_136f4_12649148 , 
    R_119e8_1153e798 , 
    R_1391b_12b277f8 , 
    R_fd37_120394f8 , 
    R_1461d_11539dd8 , 
    R_ee50_102eb9e8 , 
    R_dd_132f61c8 , 
    R_232_105afa58 , 
    R_4c_12652b08 , 
    R_135a0_1153f0f8 , 
    R_125d0_12b3f6d8 , 
    R_b4_13302988 , 
    R_51_13309648 , 
    R_f925_12048b98 , 
    R_14034_f8cf198 , 
    R_123e9_f8c0eb8 , 
    R_14726_1203bc58 , 
    R_10894_1153ad78 , 
    R_1b9_1379b7a8 , 
    R_156_137927e8 , 
    R_1471a_1379da08 , 
    R_13d4e_11544f58 , 
    R_112ae_115429d8 , 
    R_dcb0_10564e18 , 
    R_13ae3_12083498 , 
    R_11a90_13a1ba88 , 
    R_13f1a_10566998 , 
    R_fdd5_1264d068 , 
    R_13acb_13a17988 , 
    R_ef1_13a16ee8 , 
    R_145e1_12b40d58 , 
    R_14915_102f7748 , 
    R_ed3c_120760b8 , 
    R_13cdc_11542398 , 
    R_f544_102f5d08 , 
    R_147e7_13793fa8 , 
    R_e4_133095a8 , 
    R_8d_1153d078 , 
    R_78_12044178 , 
    R_22b_12b3b538 , 
    R_128ff_105b6178 , 
    R_148ac_102f0f88 , 
    R_1e9_133208a8 , 
    R_192_12b44a98 , 
    R_17d_12661f28 , 
    R_12b83_13305e08 , 
    R_fbb3_10567078 , 
    R_126_12660588 , 
    R_cfc6_1264a868 , 
    R_1492a_13a1e1e8 , 
    R_116bb_1207d6d8 , 
    R_144d8_1330d9c8 , 
    R_e6f2_102ecc08 , 
    R_14a14_1207bdd8 , 
    R_10f70_11544a58 , 
    R_119fa_1207f2f8 , 
    R_cef5_1265b6c8 , 
    R_115b3_12082458 , 
    R_211_1265c028 , 
    R_146cc_11542618 , 
    R_fe_120448f8 , 
    R_119df_1056bad8 , 
    R_13787_11ce21e8 , 
    R_147dd_11ce6068 , 
    R_14695_11cdf8a8 , 
    R_149b1_102fa128 , 
    R_110af_1379aee8 , 
    R_14560_1330b3a8 , 
    R_143ff_11cdca68 , 
    R_d4_12654a48 , 
    R_23b_13799408 , 
    R_1c7_132fc0c8 , 
    R_148_105aacd8 , 
    R_13d6d_13a17668 , 
    R_ce64_1056f9f8 , 
    R_14474_13307a28 , 
    R_12bde_102f62a8 , 
    R_1436a_102eefa8 , 
    R_14957_11540db8 , 
    R_b634_11cdc068 , 
    R_1460e_11ce2dc8 , 
    R_f24f_11ce2fa8 , 
    R_13763_105679d8 , 
    R_f0b2_102f7f68 , 
    R_14620_11ce6108 , 
    R_131f5_12084618 , 
    R_1490f_12651e88 , 
    R_136cc_1264fcc8 , 
    R_f227_1207a398 , 
    R_13959_1153f918 , 
    R_142cf_12659aa8 , 
    R_f6b2_11cdfb28 , 
    R_1ed_1203f5d8 , 
    R_a2f6_11cdb3e8 , 
    R_fc5e_13a18888 , 
    R_122_12663d28 , 
    R_13f67_12083b78 , 
    R_13740_11cdb348 , 
    R_146c9_1153fd78 , 
    R_145db_13a12b68 , 
    R_101ae_13a1fae8 , 
    R_bb03_12b29ff8 , 
    R_1101b_12045f38 , 
    R_12bfd_10564b98 , 
    R_121a5_1056a138 , 
    R_127df_1330a728 , 
    R_11617_105656d8 , 
    R_13f90_12080518 , 
    R_13be9_12662388 , 
    R_12760_1331ab88 , 
    R_126bb_10563b58 , 
    R_147c6_12081cd8 , 
    R_21c_12b41398 , 
    R_13b33_102f0588 , 
    R_1f8_132f5fe8 , 
    R_11d2f_105665d8 , 
    R_1227d_1265f2c8 , 
    R_11a35_102f44a8 , 
    R_1479c_1056c758 , 
    R_116e4_12659828 , 
    R_14662_1207ceb8 , 
    R_14515_12079ad8 , 
    R_117_12650c68 , 
    R_115ca_11ce5fc8 , 
    R_f3_1379bde8 , 
    R_e229_102ecca8 , 
    R_202_12b3f098 , 
    R_1e5_1203a218 , 
    R_12a_1331fea8 , 
    R_10d_1330bda8 , 
    R_135d6_1056fef8 , 
    R_14918_13a1d888 , 
    R_1452a_10564378 , 
    R_14984_1056bc18 , 
    R_1cd_1265c8e8 , 
    R_eb34_11cda628 , 
    R_125ac_11ce4308 , 
    R_193_f8c7cb8 , 
    R_1216d_1264d7e8 , 
    R_17c_132fe648 , 
    R_142_13792ce8 , 
    R_cdb8_102f4f48 , 
    R_144bd_11cdeb88 , 
    R_131ae_1056bd58 , 
    R_14909_1379f768 , 
    R_14924_12b3adb8 , 
    R_102a2_12b41e38 , 
    R_13aa8_120525f8 , 
    R_d3ca_102ef7c8 , 
    R_1459f_120792b8 , 
    R_120b3_12b407b8 , 
    R_127a7_105683d8 , 
    R_14545_1056b218 , 
    R_12056_1204f178 , 
    R_11f2a_10563ab8 , 
    R_e021_12b26718 , 
    R_f377_1056d1f8 , 
    R_127ca_13a16da8 , 
    R_14689_120838f8 , 
    R_11be7_1207a6b8 , 
    R_139a1_1264c668 , 
    R_14536_12b42978 , 
    R_13c2d_11cdd828 , 
    R_14906_11544ff8 , 
    R_11a5d_132f52c8 , 
    R_ca63_1331c8e8 , 
    R_14714_102f77e8 , 
    R_14799_137933c8 , 
    R_1390f_13a14828 , 
    R_1234f_12083858 , 
    R_142c6_12081738 , 
    R_127ae_12b3ccf8 , 
    R_13590_12079a38 , 
    R_148b8_102eaa48 , 
    R_5735_137a0988 , 
    R_1a6_12038698 , 
    R_169_1203e458 , 
    R_127c1_12082638 , 
    R_1288a_137a1ec8 , 
    R_1488e_102f6708 , 
    R_113b9_1264ea08 , 
    R_1430f_11cd8fa8 , 
    R_f97f_13304dc8 , 
    R_104fa_120761f8 , 
    R_119ae_11cdfa88 , 
    R_12c78_1207ca58 , 
    R_d606_11ce46c8 , 
    R_146a5_102f90e8 , 
    R_14900_120781d8 , 
    R_1374f_13a16808 , 
    R_ff3c_11ce1f68 , 
    R_e834_10564238 , 
    R_14a5e_105aa4b8 , 
    R_13465_13316bc8 , 
    R_13d25_11540b38 , 
    R_56_13308248 , 
    R_ef7_1153e838 , 
    R_13193_102ec7a8 , 
    R_132f1_13a145a8 , 
    R_1291e_1056ee18 , 
    R_14921_105640f8 , 
    R_1371a_12083fd8 , 
    R_14837_132f32e8 , 
    R_13a37_12b3d338 , 
    R_dad2_1379c6a8 , 
    R_1495d_12b43878 , 
    R_149f3_12b27c58 , 
    R_107c6_1203f998 , 
    R_1456c_12b437d8 , 
    R_11888_13794868 , 
    R_13b62_13a13428 , 
    R_1360f_10563158 , 
    R_1b1_12657ac8 , 
    R_10844_1153e1f8 , 
    R_194_1331d4c8 , 
    R_17b_1265ea08 , 
    R_15e_126544a8 , 
    R_be25_102ec028 , 
    R_148fd_102eb768 , 
    R_14683_13a1d9c8 , 
    R_a069_12080298 , 
    R_1233a_13a143c8 , 
    R_6e_13304b48 , 
    R_1334f_1204e598 , 
    R_121e7_1207ff78 , 
    R_12bb7_102f3e68 , 
    R_12bcc_12652608 , 
    R_f783_13797b08 , 
    R_14680_12076fb8 , 
    R_13d2b_12085338 , 
    R_11bbe_1153de38 , 
    R_148e8_1264bda8 , 
    R_148fa_102f5948 , 
    R_149d8_132fc168 , 
    R_148ee_120808d8 , 
    R_148f4_11cd8468 , 
    R_ff98_12b41618 , 
    R_13bc3_102f8d28 , 
    R_12b1f_120564d8 , 
    R_c961_12080f18 , 
    R_214_12655588 , 
    R_dff5_102ed9c8 , 
    R_13d49_13a16bc8 , 
    R_fb_1379f808 , 
    R_12958_102f1848 , 
    R_12220_1379e908 , 
    R_144de_12076798 , 
    R_c6d1_10566178 , 
    R_11547_1264cc08 , 
    R_138ac_102eb128 , 
    R_12853_105b58b8 , 
    R_1f1_12655268 , 
    R_11e_12b29b98 , 
    R_13d30_1207b658 , 
    R_b2_105aa0f8 , 
    R_d5a1_105690f8 , 
    R_c700_13304788 , 
    R_a359_12662888 , 
    R_1449f_12055898 , 
    R_14587_10565ef8 , 
    R_14759_1056e378 , 
    R_1385d_1056ab38 , 
    R_1401f_132fb588 , 
    R_1245b_12658f68 , 
    R_fe3a_11cdb168 , 
    R_a47d_13a18f68 , 
    R_145ea_1056c438 , 
    R_99a4_102f5bc8 , 
    R_1491e_12661528 , 
    R_1c1_126618e8 , 
    R_b180_12039a98 , 
    R_14e_12b29e18 , 
    R_13b1f_12052c38 , 
    R_146e4_f8cb638 , 
    R_14581_10571b18 , 
    R_1354d_12040078 , 
    R_13508_120842f8 , 
    R_148d9_13a14d28 , 
    R_149c0_102ed068 , 
    R_1477e_10568fb8 , 
    R_14735_105680b8 , 
    R_13d35_11ce1108 , 
    R_4d49_102f8dc8 , 
    R_133aa_11545b38 , 
    R_14518_102f67a8 , 
    R_bf1d_1153d618 , 
    R_a9_1204d4b8 , 
    R_14702_12b3d0b8 , 
    R_1431c_11cde188 , 
    R_9323_1331d068 , 
    R_14a2f_12075ed8 , 
    R_1e1_13321ca8 , 
    R_12e_105af9b8 , 
    R_9d_1379c9c8 , 
    R_12caa_126508a8 , 
    R_115df_10566c18 , 
    R_144fd_102f1b68 , 
    R_127f1_12b2a098 , 
    R_137eb_12082138 , 
    R_11b9a_12b3f278 , 
    R_1483a_12081f58 , 
    R_7d2b_11ce4948 , 
    R_13a49_102f8e68 , 
    R_1493c_11cdc568 , 
    R_14a3e_102ed428 , 
    R_195_12045cb8 , 
    R_14489_12b3fe58 , 
    R_17a_1330dc48 , 
    R_1066b_1264a228 , 
    R_139b5_11536318 , 
    R_12775_126513e8 , 
    R_13d43_13a1c168 , 
    R_13e78_1056a598 , 
    R_90_f8cccb8 , 
    R_75_12b443b8 , 
    R_14816_10565db8 , 
    R_e4c7_10571398 , 
    R_14354_13317348 , 
    R_146c3_12b3bfd8 , 
    R_db95_12b2ff98 , 
    R_b45b_11ce7508 , 
    R_145de_1056b5d8 , 
    R_13c7d_1056d798 , 
    R_c7c0_102ed4c8 , 
    R_1ff_13315c28 , 
    R_1361a_102f01c8 , 
    R_110_1204b938 , 
    R_10c17_13a13888 , 
    R_d6_1264b1c8 , 
    R_239_12b2a958 , 
    R_144a8_115369f8 , 
    R_12516_13305188 , 
    R_14699_10567e38 , 
    R_12de4_12045b18 , 
    R_10fd9_11ce1928 , 
    R_145c6_13a1cb68 , 
    R_147c3_13a177a8 , 
    R_1313e_1207a1b8 , 
    R_e9a6_1153dcf8 , 
    R_123a6_12077418 , 
    R_e669_1056eb98 , 
    R_eea5_13793c88 , 
    R_8e12_f8c7538 , 
    R_11a2c_12b3f1d8 , 
    R_bc89_12664548 , 
    R_b132_13300a88 , 
    R_14626_102f4ae8 , 
    R_125c9_11ce5c08 , 
    R_14891_1265e0a8 , 
    R_13ba9_1056f4f8 , 
    R_11299_1056a4f8 , 
    R_1395f_1207ba18 , 
    R_1085f_13312a28 , 
    R_c642_12b41b18 , 
    R_1445c_f8ce478 , 
    R_14981_12b3f598 , 
    R_148e2_12650b28 , 
    R_988f_13a1e968 , 
    R_962b_105647d8 , 
    R_124a7_12079498 , 
    R_fe64_1153f378 , 
    R_11f16_102eb088 , 
    R_13e03_1379bf28 , 
    R_14927_11cdf808 , 
    R_1ba_1330eb48 , 
    R_14471_13793be8 , 
    R_121fd_11ce3048 , 
    R_14499_1207a9d8 , 
    R_155_12b43f58 , 
    R_98_12048af8 , 
    R_e916_105699b8 , 
    R_e1ea_1056b998 , 
    R_11af3_13793788 , 
    R_13bcf_12650948 , 
    R_10070_12077e18 , 
    R_f2f6_126613e8 , 
    R_104a3_11542d98 , 
    R_149ae_10565138 , 
    R_1430b_1204c8d8 , 
    R_ede8_1056dfb8 , 
    R_13495_13a1e008 , 
    R_df_132f6808 , 
    R_230_12664a48 , 
    R_136ac_102eacc8 , 
    R_dd20_137974c8 , 
    R_14741_132f2c08 , 
    R_137c1_11543dd8 , 
    R_14364_11ce6568 , 
    R_11d60_132fc8e8 , 
    R_14a44_105b60d8 , 
    R_13749_11543518 , 
    R_854a_1207fed8 , 
    R_14a11_12045a78 , 
    R_1a7_12659b48 , 
    R_168_105b3158 , 
    R_f03_13a17208 , 
    R_1274c_12653fa8 , 
    R_147b7_12079df8 , 
    R_a2_1379e228 , 
    R_63_f8c7b78 , 
    R_13c49_102ecac8 , 
    R_d68f_12078a98 , 
    R_148f1_11cde688 , 
    R_196_11536778 , 
    R_179_13301c08 , 
    R_11c1b_120757f8 , 
    R_1181a_10565098 , 
    R_14912_13300628 , 
    R_10c93_13310768 , 
    R_147f2_10571618 , 
    R_c832_12075f78 , 
    R_14530_11540778 , 
    R_e8ba_11ce3b88 , 
    R_14903_11ce50c8 , 
    R_14629_115412b8 , 
    R_11966_10562118 , 
    R_f8fa_105b4d78 , 
    R_1d8_1331f5e8 , 
    R_1281b_1207f6b8 , 
    R_137_1331a7c8 , 
    R_5f_12b428d8 , 
    R_12288_126495a8 , 
    R_a469_13a14648 , 
    R_130cc_13a17348 , 
    R_136e6_11cdcb08 , 
    R_d806_102f5a88 , 
    R_fd98_12052d78 , 
    R_144b4_1153eab8 , 
    R_1482b_12b3b3f8 , 
    R_13858_12081e18 , 
    R_1d3_1265ae08 , 
    R_13c_1265b1c8 , 
    R_14596_12048558 , 
    R_eb_1153bf98 , 
    R_224_12b29698 , 
    R_13d3c_132f70c8 , 
    R_c353_102f31e8 , 
    R_1092e_13a140a8 , 
    R_1018e_10563478 , 
    R_12875_1153eb58 , 
    R_13693_13795448 , 
    R_123bb_11ce7008 , 
    R_dfc9_12647208 , 
    R_da6d_12082098 , 
    R_1198e_1153d758 , 
    R_149ff_1264c848 , 
    R_1180e_12648248 , 
    R_12535_126604e8 , 
    R_12780_10568b58 , 
    R_9dc0_102f6f28 , 
    R_c4a7_1330a908 , 
    R_11bfb_12649968 , 
    R_13fe4_105622f8 , 
    R_12e0c_13797388 , 
    R_1454e_11ce1c48 , 
    R_14069_1153db18 , 
    R_10c0e_120464d8 , 
    R_13c1f_f8c8938 , 
    R_d910_1056e418 , 
    R_cfae_13a15368 , 
    R_10806_1264d608 , 
    R_13706_13319b48 , 
    R_12e21_1330cb68 , 
    R_f8_12665808 , 
    R_67_105aac38 , 
    R_217_105b3fb8 , 
    R_12a8e_1264ef08 , 
    R_e5ea_115436f8 , 
    R_14858_10571c58 , 
    R_111b8_102ebbc8 , 
    R_12ba4_12b28ab8 , 
    R_108f1_102f35a8 , 
    R_138a5_1264e468 , 
    R_131ff_13a1eaa8 , 
    R_11448_11ce41c8 , 
    R_11534_13a13ce8 , 
    R_12d1d_1207c238 , 
    R_134e8_13a1e8c8 , 
    R_b82e_1153c2b8 , 
    R_11572_11ce43a8 , 
    R_14897_1265c988 , 
    R_125fa_1265b128 , 
    R_b95d_102f8008 , 
    R_14436_10570718 , 
    R_f951_132fcde8 , 
    R_10246_1056ae58 , 
    R_12041_11ce0ac8 , 
    R_138cd_1153e018 , 
    R_1b2_12660f88 , 
    R_197_1379a768 , 
    R_121dd_12659328 , 
    R_178_12658d88 , 
    R_15d_133195a8 , 
    R_13f24_13318428 , 
    R_146f6_132fbc68 , 
    R_b880_12083d58 , 
    R_12ab4_132f57c8 , 
    R_ed14_133110c8 , 
    R_144f0_132ff0e8 , 
    R_10aa5_12053f98 , 
    R_1290a_11ce1388 , 
    R_9d4e_11cddbe8 , 
    R_e6_12b344f8 , 
    R_b0_12b3f458 , 
    R_229_126659e8 , 
    R_12b3f_105b6538 , 
    R_1f5_1203e958 , 
    R_f624_1265b808 , 
    R_14711_11ce2828 , 
    R_fe05_102f9548 , 
    R_1118b_11cdb8e8 , 
    R_1c8_f8c6b38 , 
    R_147_12b38c98 , 
    R_11a_1204b438 , 
    R_14778_13a1f688 , 
    R_137fd_11544418 , 
    R_f0_13795d08 , 
    R_c3_132ff188 , 
    R_21f_1265a2c8 , 
    R_12e60_132f3a68 , 
    R_4a02_12646e48 , 
    R_c5_12657e88 , 
    R_132ae_1056ef58 , 
    R_d400_133126a8 , 
    R_128a8_f8c9978 , 
    R_ecbd_12040a78 , 
    R_146ba_11cd8c88 , 
    R_ea59_102f5088 , 
    R_1183a_1204a498 , 
    R_13d1f_1207ddb8 , 
    R_136e0_11ce7148 , 
    R_ddb7_12078b38 , 
    R_14575_13307c08 , 
    R_14864_13a1b768 , 
    R_1471d_12040bb8 , 
    R_11237_1056f958 , 
    R_13fee_12663288 , 
    R_c1_1204fd58 , 
    R_14632_11cd85a8 , 
    R_4d_12662d88 , 
    R_b895_1264a4a8 , 
    R_11b87_12648b08 , 
    R_111c4_12076658 , 
    R_a534_12b3d018 , 
    R_11805_12b41578 , 
    R_c901_126603a8 , 
    R_13bde_13a1bbc8 , 
    R_149b4_10564d78 , 
    R_c7_126589c8 , 
    R_248_1331ef08 , 
    R_5b_12655088 , 
    R_13720_102f3f08 , 
    R_b9b1_1056c9d8 , 
    R_f1cc_10567ed8 , 
    R_cd0b_11542f78 , 
    R_1497b_11cdfda8 , 
    R_12d6f_13799b88 , 
    R_14305_120844d8 , 
    R_145ae_102efe08 , 
    R_147d6_12b27b18 , 
    R_13dc3_11cdbf28 , 
    R_dc22_1153d438 , 
    R_5970_11cdbe88 , 
    R_113_1265c528 , 
    R_82_f8cbc78 , 
    R_1fc_12050078 , 
    R_b00a_1153e658 , 
    R_1346e_10567bb8 , 
    R_1dd_12b395f8 , 
    R_10390_1207ed58 , 
    R_12cf4_13310ee8 , 
    R_10675_1203cab8 , 
    R_1399b_1264c3e8 , 
    R_132_120518d8 , 
    R_d8_12b3c938 , 
    R_237_105a9fb8 , 
    R_d4b2_1265bda8 , 
    R_14453_12649d28 , 
    R_10e2c_102ecde8 , 
    R_52_13799868 , 
    R_143dc_120824f8 , 
    R_13ebe_11ce4128 , 
    R_14053_102f21a8 , 
    R_10960_133050e8 , 
    R_1037b_1264a048 , 
    R_7fe6_12b3f638 , 
    R_12685_11cdf088 , 
    R_135e9_11ce0de8 , 
    R_bf_1379fa88 , 
    R_85_12b41898 , 
    R_149d5_11541358 , 
    R_13f4d_10561fd8 , 
    R_d0f1_1056a1d8 , 
    R_a3f3_12646da8 , 
    R_1311d_13a131a8 , 
    R_1026e_11541ad8 , 
    R_139de_13310588 , 
    R_144cc_11ce23c8 , 
    R_1403a_1331cc08 , 
    R_1ce_12656628 , 
    R_198_12b3fdb8 , 
    R_d37f_1379a1c8 , 
    R_177_1330de28 , 
    R_141_12b3cf78 , 
    R_14500_102f92c8 , 
    R_c9_12b28fb8 , 
    R_246_1203df58 , 
    R_93_12659be8 , 
    R_72_132fe788 , 
    R_125bf_105685b8 , 
    R_1a8_137a0d48 , 
    R_147a5_1264a728 , 
    R_167_1204f678 , 
    R_7f_105ac998 , 
    R_149f0_13a1fea8 , 
    R_12210_13793aa8 , 
    R_13db7_11ce11a8 , 
    R_100e9_132f3ec8 , 
    R_5362_13a18108 , 
    R_124d7_13a18e28 , 
    R_14a55_133001c8 , 
    R_12419_1153d398 , 
    R_108b6_1264e0a8 , 
    R_10d4d_11cded68 , 
    R_1464a_13a15b88 , 
    R_c7f2_11cdc748 , 
    R_13c83_11544698 , 
    R_1489a_f8c6c78 , 
    R_125b6_12040b18 , 
    R_c00b_12079718 , 
    R_eeb_13a13608 , 
    R_f088_1330ba88 , 
    R_1365e_1207b838 , 
    R_fa81_12052198 , 
    R_145f3_13a14788 , 
    R_10995_102f3148 , 
    R_123f8_13a13388 , 
    R_6358_1204fe98 , 
    R_14763_11ce4c68 , 
    R_1433c_12077c38 , 
    R_dde7_13a141e8 , 
    R_13ef9_1204a858 , 
    R_14810_1056db58 , 
    R_13fdc_102f15c8 , 
    R_d995_11ce0fc8 , 
    R_117fc_12056078 , 
    R_8d57_11ce53e8 , 
    R_11bb4_12b39cd8 , 
    R_13b97_1207a438 , 
    R_14068_11cdc108 , 
    R_1335a_105b5ef8 , 
    R_1043d_13a1c5c8 , 
    R_128cf_11cdabc8 , 
    R_1219b_1207a938 , 
    R_10dce_105631f8 , 
    R_bbfa_10564418 , 
    R_11864_12b44318 , 
    R_12435_11ce4088 , 
    R_a7_1265a5e8 , 
    R_111f4_11cdf6c8 , 
    R_135cf_1207eb78 , 
    R_102ef_1153c218 , 
    R_12ca0_11ce0668 , 
    R_1c2_1330f228 , 
    R_c6f4_12056438 , 
    R_1404f_12b3e738 , 
    R_ee7b_1379a628 , 
    R_127e9_f8c8078 , 
    R_14d_1203cbf8 , 
    R_bd_1203f3f8 , 
    R_48_13301848 , 
    R_10afa_13a15d68 , 
    R_ed66_11ce3368 , 
    R_13a92_102f0bc8 , 
    R_e9fb_12646268 , 
    R_10d30_12084078 , 
    R_149ab_1153d7f8 , 
    R_88_13300d08 , 
    R_6b_105aaff8 , 
    R_11c31_115418f8 , 
    R_13677_102f9868 , 
    R_133f2_1379f088 , 
    R_13edf_120837b8 , 
    R_d399_137980a8 , 
    R_1446e_1207d958 , 
    R_1382d_1207d9f8 , 
    R_cb_1331fa48 , 
    R_244_1264c708 , 
    R_12dc8_13a1f548 , 
    R_12299_1265d1a8 , 
    R_1474a_12076dd8 , 
    R_13844_12663aa8 , 
    R_13c11_1153d578 , 
    R_14650_1056f278 , 
    R_146fc_12647848 , 
    R_10f84_1207bab8 , 
    R_131cc_12b272f8 , 
    R_1451b_10567cf8 , 
    R_14390_10567c58 , 
    R_13754_12082318 , 
    R_1bb_12664868 , 
    R_154_1204e1d8 , 
    R_14831_1264f408 , 
    R_7c_105b1cb8 , 
    R_f1a0_12075938 , 
    R_e9d0_1153f558 , 
    R_f0eb_102f7568 , 
    R_fb0c_1331a368 , 
    R_1397b_1331b268 , 
    R_e589_1379bb68 , 
    R_1381a_120547b8 , 
    R_1463e_105703f8 , 
    R_12e76_11cd9908 , 
    R_199_132fb3a8 , 
    R_176_12b265d8 , 
    R_125_13798008 , 
    R_11ad2_102ed108 , 
    R_1ea_1265a868 , 
    R_10764_11cd9548 , 
    R_14563_1264d6a8 , 
    R_12c1a_102f0268 , 
    R_146d2_1203a998 , 
    R_147bd_102f9048 , 
    R_fa57_1207f398 , 
    R_c5a3_120849d8 , 
    R_11dc9_f8c9b58 , 
    R_11d95_1153f198 , 
    R_1329b_11cd95e8 , 
    R_14861_f8c41f8 , 
    R_1064a_10561f38 , 
    R_ce07_f8c8f78 , 
    R_14720_11ce07a8 , 
    R_13ca7_12078098 , 
    R_147f5_1207a078 , 
    R_142d3_12036758 , 
    R_13dee_12083a38 , 
    R_ec91_126490a8 , 
    R_13421_11544c38 , 
    R_cf92_11cdfee8 , 
    R_4c49_13a1d748 , 
    R_114d1_13307de8 , 
    R_cff7_12076bf8 , 
    R_142ff_11ce1b08 , 
    R_139c0_13a1e5a8 , 
    R_143cc_1056e738 , 
    R_ba4e_13a1d388 , 
    R_12485_105b6358 , 
    R_11f0c_13a1aea8 , 
    R_14867_12054b78 , 
    R_137b5_10569cd8 , 
    R_11d1b_12649288 , 
    R_13d7b_102f56c8 , 
    R_14a2c_102f12a8 , 
    R_14608_13a155e8 , 
    R_144c9_10571578 , 
    R_fc0a_11541858 , 
    R_144fa_120775f8 , 
    R_129_1331c988 , 
    R_13561_1330d068 , 
    R_e1_12661708 , 
    R_1299a_1207b158 , 
    R_1489d_105686f8 , 
    R_22e_132f2ac8 , 
    R_6d01_102f72e8 , 
    R_ffc3_12656e48 , 
    R_1496f_102f9908 , 
    R_1e6_13792a68 , 
    R_14760_11ce3868 , 
    R_d2d1_13793468 , 
    R_12145_1207b978 , 
    R_f5_11537038 , 
    R_bb_13799cc8 , 
    R_21a_1265b088 , 
    R_14975_11541998 , 
    R_147c0_11ce20a8 , 
    R_13b7f_1153a198 , 
    R_13615_12084c58 , 
    R_14a29_10571438 , 
    R_13526_102f49a8 , 
    R_11215_12075b18 , 
    R_10e4c_13a169e8 , 
    R_13d97_105651d8 , 
    R_1b3_1379b348 , 
    R_13fab_11538758 , 
    R_10ff9_105aad78 , 
    R_145c0_11cd7f68 , 
    R_145fc_120476f8 , 
    R_15c_137992c8 , 
    R_67bc_13311028 , 
    R_efc2_11cdefe8 , 
    R_145cc_132f8388 , 
    R_ae_1379c1a8 , 
    R_1263c_11cdf768 , 
    R_57_126522e8 , 
    R_14659_1264e1e8 , 
    R_13899_133075c8 , 
    R_125e5_13311348 , 
    R_113fb_11ce7288 , 
    R_11e0e_102f4908 , 
    R_11270_12b29a58 , 
    R_f61a_13305cc8 , 
    R_1499f_133198c8 , 
    R_121_13795808 , 
    R_106_12b25a98 , 
    R_1458a_102eb268 , 
    R_126cf_13a19788 , 
    R_209_1379cb08 , 
    R_1ee_12656268 , 
    R_12c5a_102ef688 , 
    R_1270e_11cdb708 , 
    R_e437_102f2c48 , 
    R_147cf_11ce5168 , 
    R_e233_1056d338 , 
    R_13bbe_11ce55c8 , 
    R_11e6b_1207d458 , 
    R_13f0b_12b42f18 , 
    R_103_12b41c58 , 
    R_cd_12b39a58 , 
    R_242_12654688 , 
    R_20c_12b43c38 , 
    R_11ce5_1379e048 , 
    R_ef4_1056dc98 , 
    R_11823_13a15fe8 , 
    R_130b8_13a12988 , 
    R_12baf_12648ba8 , 
    R_119a4_102f3288 , 
    R_f4e5_1264b308 , 
    R_12c6f_11cdea48 , 
    R_1473b_102fa308 , 
    R_8b_132f8608 , 
    R_11467_105659f8 , 
    R_11b4a_11ce1568 , 
    R_137f7_12077878 , 
    R_e5b5_1153d938 , 
    R_14775_13a1bda8 , 
    R_14671_1264ab88 , 
    R_14066_12084258 , 
    R_13954_12076518 , 
    R_de4d_12b26538 , 
    R_149f6_11cda308 , 
    R_aff6_102f4a48 , 
    R_d75d_1207c0f8 , 
    R_10f46_12081ff8 , 
    R_c50b_11cdd3c8 , 
    R_136ed_12082ef8 , 
    R_101d1_1056e198 , 
    R_1a9_12037658 , 
    R_166_120507f8 , 
    R_9b_12b3b178 , 
    R_bb16_12650268 , 
    R_1265a_105635b8 , 
    R_b802_1265dba8 , 
    R_131ea_102f4cc8 , 
    R_14a0e_10570e98 , 
    R_19a_12662068 , 
    R_175_12b3fc78 , 
    R_109_12b2c7f8 , 
    R_206_105b5b38 , 
    R_146b4_1153fcd8 , 
    R_11e21_11cd9e08 , 
    R_104ba_f8c7218 , 
    R_13fbc_11541218 , 
    R_144ba_102f8c88 , 
    R_11622_102ed388 , 
    R_13c02_12b29198 , 
    R_13ba3_105626b8 , 
    R_ff0f_12081918 , 
    R_123d6_11541e98 , 
    R_fd64_102f3328 , 
    R_14486_102ef728 , 
    R_13776_1379fd08 , 
    R_14665_132f5ae8 , 
    R_10098_13793968 , 
    R_11072_13a1ed28 , 
    R_14554_10565778 , 
    R_137a8_1056b678 , 
    R_11b55_12649a08 , 
    R_14411_12663508 , 
    R_84a7_12b40fd8 , 
    R_133fc_1153ee78 , 
    R_da_1331b088 , 
    R_a0_1379b2a8 , 
    R_235_1264d4c8 , 
    R_1333b_11542c58 , 
    R_132e7_11ce28c8 , 
    R_1357d_1153feb8 , 
    R_14644_1056d978 , 
    R_100_1265f0e8 , 
    R_79_137a1388 , 
    R_e0d7_126556c8 , 
    R_11b42_1264b6c8 , 
    R_20f_12b28018 , 
    R_f4db_1207bfb8 , 
    R_1193e_13a19968 , 
    R_138d5_1379b848 , 
    R_13e4c_1207f118 , 
    R_13a7e_102f6ac8 , 
    R_12d79_102ee468 , 
    R_116a8_12084398 , 
    R_116_1265f868 , 
    R_148a3_11cdecc8 , 
    R_13273_13a1a688 , 
    R_1f9_1379ddc8 , 
    R_1025b_1330bee8 , 
    R_122e8_12b39878 , 
    R_11ba2_11544738 , 
    R_12521_1056c258 , 
    R_e8e6_f8cf4b8 , 
    R_8cd2_1264ac28 , 
    R_11a11_126477a8 , 
    R_143c6_120850b8 , 
    R_13e99_12039e58 , 
    R_1466b_13306808 , 
    R_14465_1207a758 , 
    R_134b3_102f3468 , 
    R_11fe7_1330c3e8 , 
    R_1258d_13a14dc8 , 
    R_14677_105712f8 , 
    R_1367d_102eb628 , 
    R_1e2_12663c88 , 
    R_b9_12661848 , 
    R_12d_12660268 , 
    R_f47c_1153ded8 , 
    R_1468c_13a1aae8 , 
    R_145ba_120815f8 , 
    R_14790_11cd9cc8 , 
    R_14419_12048f58 , 
    R_13bb3_1207b6f8 , 
    R_1046b_105688d8 , 
    R_1232e_13314008 , 
    R_1170d_1264c528 , 
    R_14a41_1056fa98 , 
    R_14459_11cd92c8 , 
    R_14480_11cdcf68 , 
    R_13a88_11ce3f48 , 
    R_c8f0_102f0d08 , 
    R_134ff_1056bf38 , 
    R_aac5_13a18748 , 
    R_14509_13a1e148 , 
    R_cebc_12039d18 , 
    R_135bd_12081058 , 
    R_147ba_12078ef8 , 
    R_f4a6_105654f8 , 
    R_1182e_13a19aa8 , 
    R_142eb_11cdec28 , 
    R_13bf5_10568ab8 , 
    R_12093_12077058 , 
    R_13dac_13a15688 , 
    R_dc51_13304f08 , 
    R_13e8f_1264a0e8 , 
    R_13c89_12b39f58 , 
    R_f0be_102f1de8 , 
    R_9373_10563e78 , 
    R_11a48_13a195a8 , 
    R_f3f9_1153f9b8 , 
    R_1d4_12b42fb8 , 
    R_e3f1_12b25bd8 , 
    R_13c27_13309b48 , 
    R_240_105ab4f8 , 
    R_cf_13311a28 , 
    R_13c38_1204a3f8 , 
    R_13b_13300f88 , 
    R_11ef6_11cd7888 , 
    R_135c9_11ce6888 , 
    R_116d1_1153d898 , 
    R_149d2_12080158 , 
    R_ba5b_12b403f8 , 
    R_ea84_1330ca28 , 
    R_f59a_11ce3908 , 
    R_1496c_1331e968 , 
    R_12bd5_11ce3fe8 , 
    R_1253e_105b6678 , 
    R_14873_11cd79c8 , 
    R_149a5_132ff868 , 
    R_14512_11540bd8 , 
    R_14756_10565318 , 
    R_1c9_13313a68 , 
    R_d09b_12660948 , 
    R_203_12050cf8 , 
    R_10c_12038058 , 
    R_146_12b42298 , 
    R_136c1_12b276b8 , 
    R_1480a_12649e68 , 
    R_1d9_1379e7c8 , 
    R_13e84_1056ad18 , 
    R_1021c_1056fc78 , 
    R_136_132fe6e8 , 
    R_145ff_102ef2c8 , 
    R_19b_12b28dd8 , 
    R_1031a_11540e58 , 
    R_1f2_11538438 , 
    R_13114_102f3648 , 
    R_ec36_12042af8 , 
    R_222_133189c8 , 
    R_6f_12b3a458 , 
    R_96_1203c838 , 
    R_ed_1203deb8 , 
    R_11d_1204c838 , 
    R_174_13318928 , 
    R_119f1_13316588 , 
    R_1486a_13a1d428 , 
    R_11717_1207d778 , 
    R_14781_115447d8 , 
    R_13995_12038738 , 
    R_e4f5_12049598 , 
    R_74a9_12645d68 , 
    R_10208_12038558 , 
    R_145ab_12b3f9f8 , 
    R_227_1331e508 , 
    R_e8_133028e8 , 
    R_13809_1153faf8 , 
    R_f732_12649008 , 
    R_14524_137968e8 , 
    R_146d8_11cd94a8 , 
    R_14064_1264d2e8 , 
    R_12dfa_11cd88c8 , 
    R_135ef_102f0a88 , 
    R_10ee5_12047798 , 
    R_14548_120493b8 , 
    R_11030_11cdbca8 , 
    R_1400f_13a1a368 , 
    R_f051_1264e6e8 , 
    R_de7c_102eafe8 , 
    R_13538_120754d8 , 
    R_13e56_12b297d8 , 
    R_84eb_1331c2a8 , 
    R_1498a_1207e3f8 , 
    R_148a6_115459f8 , 
    R_212_1330bd08 , 
    R_fd_13307d48 , 
    R_144a5_13a1c028 , 
    R_10110_120369d8 , 
    R_12b5e_12651208 , 
    R_149ed_13303428 , 
    R_144db_12078598 , 
    R_bf9f_11cd9b88 , 
    R_14017_f8c20d8 , 
    R_13a3d_f8ca918 , 
    R_13b2d_120830d8 , 
    R_8e_132f37e8 , 
    R_12aeb_120810f8 , 
    R_a23e_11ce5ca8 , 
    R_12ce9_12081c38 , 
    R_f00_1207c058 , 
    R_c1fe_1264be48 , 
    R_f2d2_11cdf948 , 
    R_14385_12044c18 , 
    R_143c0_1265fb88 , 
    R_14496_13a1c668 , 
    R_14738_12b28bf8 , 
    R_cab9_102f99a8 , 
    R_1255c_f8c61d8 , 
    R_143ba_11cde868 , 
    R_147c9_13a18ce8 , 
    R_13311_13a198c8 , 
    R_147a2_102f2ce8 , 
    R_fbe0_13a1b628 , 
    R_dcc6_12664ae8 , 
    R_103cf_12085158 , 
    R_13909_1204f5d8 , 
    R_1197b_115433d8 , 
    R_144e1_13a1f4a8 , 
    R_145a2_11cd7ce8 , 
    R_12d50_120851f8 , 
    R_12380_10563338 , 
    R_107a7_1379f9e8 , 
    R_10e8a_102ea688 , 
    R_122fb_13a17708 , 
    R_12aa7_12037798 , 
    R_12107_1264d428 , 
    R_14533_1330c8e8 , 
    R_14542_120759d8 , 
    R_4276_102effe8 , 
    R_1478d_115453b8 , 
    R_130c1_11542258 , 
    R_13ff8_102f9fe8 , 
    R_1aa_13795268 , 
    R_116b1_13a159a8 , 
    R_1bc_126536e8 , 
    R_b76e_1153c8f8 , 
    R_4e_13792e28 , 
    R_60_12b44bd8 , 
    R_a5_13311668 , 
    R_b7_1379f948 , 
    R_153_13793288 , 
    R_165_13306948 , 
    R_f9fe_102f9408 , 
    R_14431_12080478 , 
    R_1c3_12047158 , 
    R_64_f8c1bd8 , 
    R_14c_120387d8 , 
    R_12471_102f7068 , 
    R_148c1_13316f88 , 
    R_11433_1265f048 , 
    R_13ce2_1264aa48 , 
    R_121bd_115449b8 , 
    R_14813_10566d58 , 
    R_147fb_102f83c8 , 
    R_146ab_12051658 , 
    R_12c65_1264cb68 , 
    R_e2b4_f8c0f58 , 
    R_10c61_120805b8 , 
    R_10f1d_10566df8 , 
    R_10de4_1379b5c8 , 
    R_ae51_105ab098 , 
    R_146f3_12659d28 , 
    R_d03f_126484c8 , 
    R_9fe2_11543fb8 , 
    R_10b79_12657028 , 
    R_64c2_12662748 , 
    R_139d0_102f1fc8 , 
    R_13639_1207f578 , 
    R_1b4_12654728 , 
    R_1cf_133184c8 , 
    R_e214_1207ae38 , 
    R_140_12665448 , 
    R_15b_f8c0378 , 
    R_1435c_13304d28 , 
    R_10745_12056898 , 
    R_1044f_120557f8 , 
    R_10824_11ce3188 , 
    R_13820_12b41438 , 
    R_69b8_11cdc888 , 
    R_124b9_1056d658 , 
    R_143f4_102edd88 , 
    R_142f5_1264a908 , 
    R_76_f8ca198 , 
    R_ac_12660a88 , 
    R_1269b_11cd9368 , 
    R_147b4_120766f8 , 
    R_14834_13a16a88 , 
    R_12e88_102f8a08 , 
    R_f021_102ec168 , 
    R_f6dd_13a163a8 , 
    R_145e4_126463a8 , 
    R_14723_1264db08 , 
    R_173_f8c3438 , 
    R_19c_12b40218 , 
    R_11142_10562f78 , 
    R_23e_1265bc68 , 
    R_d1_13311f28 , 
    R_13512_12080dd8 , 
    R_7859_11cdaee8 , 
    R_14593_115458b8 , 
    R_148a9_12647ac8 , 
    R_10577_11545318 , 
    R_133ca_1203e098 , 
    R_13b92_13a14be8 , 
    R_10efd_102ec3e8 , 
    R_f0b_1153f4b8 , 
    R_12e15_10568018 , 
    R_200_12b29eb8 , 
    R_21d_137a03e8 , 
    R_f2_12652ec8 , 
    R_10f_12b3e5f8 , 
    R_ca13_11ce4628 , 
    R_14966_11546218 , 
    R_13ad8_1203a358 , 
    R_12d8d_105b5db8 , 
    R_10165_1264cac8 , 
    R_1337f_13a12c08 , 
    R_53_f8c2a38 , 
    R_149c9_132f4fa8 , 
    R_10aae_1207c558 , 
    R_13aad_11541a38 , 
    R_12362_10563dd8 , 
    R_5c4e_1056ced8 , 
    R_130f5_1056a098 , 
    R_12a7c_11cdde68 , 
    R_14415_12b2a318 , 
    R_1488b_13a189c8 , 
    R_14062_1204cf18 , 
    R_14784_11cd8508 , 
    R_1032f_10570f38 , 
    R_9bdf_102ee5a8 , 
    R_13bf0_1331c528 , 
    R_11b90_11ce0208 , 
    R_149cf_13a17b68 , 
    R_12021_11ce25a8 , 
    R_1de_12056d98 , 
    R_49_1331f4a8 , 
    R_131_105ab3b8 , 
    R_1462f_13794688 , 
    R_10628_1203d2d8 , 
    R_122bf_10570038 , 
    R_11387_11540d18 , 
    R_11fa6_13306308 , 
    R_85b5_120819b8 , 
    R_142ef_102eec88 , 
    R_1434c_102f13e8 , 
    R_22c_1379b708 , 
    R_5c_137944a8 , 
    R_e3_1203e778 , 
    R_b948_1153a5f8 , 
    R_e169_11cd7a68 , 
    R_d051_11536ef8 , 
    R_10e01_120551b8 , 
    R_233_12b392d8 , 
    R_68_12b283d8 , 
    R_dc_13300768 , 
    R_13bfb_13316a88 , 
    R_10ad6_10565598 , 
    R_14870_10570538 , 
    R_12260_13a1b268 , 
    R_d661_1265cfc8 , 
    R_14572_11cd9d68 , 
    R_130ff_12078318 , 
    R_a98a_11cdaf88 , 
    R_14978_12b321f8 , 
    R_14a1a_115445f8 , 
    R_14a26_13792568 , 
    R_b327_12648568 , 
    R_108fb_105b5e58 , 
    R_1440d_11544238 , 
    R_10cff_13a1dc48 , 
    R_139ae_11cd8b48 , 
    R_14338_11cda808 , 
    R_106b3_13a16088 , 
    R_c4f8_11ce12e8 , 
    R_215_1265b948 , 
    R_fa_133070c8 , 
    R_11b68_1264ec88 , 
    R_129b1_1056f098 , 
    R_13670_10564558 , 
    R_1439c_11cdd148 , 
    R_107e6_11cdbc08 , 
    R_f279_13a1acc8 , 
    R_12ed9_102edf68 , 
    R_12bc1_13a1f048 , 
    R_13b19_12b2ba38 , 
    R_e361_120812d8 , 
    R_bef9_11ce0528 , 
    R_13ce8_120793f8 , 
    R_a235_12084a78 , 
    R_14521_1264f228 , 
    R_13cad_13a1edc8 , 
    R_148af_11540098 , 
    R_10968_13304968 , 
    R_13fcb_102f0c68 , 
    R_11645_13304e68 , 
    R_bf09_1056b498 , 
    R_12553_13310308 , 
    R_145d5_132fa228 , 
    R_146a2_1207bf18 , 
    R_136fc_12076018 , 
    R_149a2_1264d1a8 , 
    R_12b9a_13a14968 , 
    R_137cc_10569af8 , 
    R_c5ef_12081238 , 
    R_1184d_11cd9188 , 
    R_13c8f_102ed568 , 
    R_109bf_1379c248 , 
    R_14326_13301528 , 
    R_11123_12045258 , 
    R_e197_11ce3228 , 
    R_172_126656c8 , 
    R_19d_132ffb88 , 
    R_c306_f8c5418 , 
    R_b5_133157c8 , 
    R_13902_13799ae8 , 
    R_14348_1056c398 , 
    R_1457b_102f5628 , 
    R_14766_105674d8 , 
    R_d2c1_12036e38 , 
    R_1f6_1330dce8 , 
    R_10c28_12080e78 , 
    R_119_133166c8 , 
    R_1300e_12646bc8 , 
    R_13129_10567b18 , 
    R_1394d_1056f318 , 
    R_14846_13798b48 , 
    R_146cf_1379e868 , 
    R_10019_11542118 , 
    R_fb35_132fb4e8 , 
    R_11a23_126506c8 , 
    R_9aae_1056dbf8 , 
    R_14468_1264aea8 , 
    R_7aaf_f8c22b8 , 
    R_b5af_1264e508 , 
    R_13f11_11cd7b08 , 
    R_e6c6_12075cf8 , 
    R_14374_102f0768 , 
    R_14605_13a182e8 , 
    R_13de4_102f94a8 , 
    R_102c2_1264ed28 , 
    R_91_13799548 , 
    R_135f5_11cda4e8 , 
    R_14807_1331e288 , 
    R_14a08_11cdc388 , 
    R_cb44_12b3ee18 , 
    R_13a63_11544198 , 
    R_109ca_1264cd48 , 
    R_12e41_10569198 , 
    R_e46a_13a181a8 , 
    R_12963_13a1afe8 , 
    R_14a5a_12b42158 , 
    R_13e38_1207efd8 , 
    R_144ea_1264f5e8 , 
    R_11668_137a1d88 , 
    R_13ec7_11540318 , 
    R_ff67_13799688 , 
    R_13b27_102eb588 , 
    R_fa2a_1056e0f8 , 
    R_145a5_132f4dc8 , 
    R_14060_13a15ae8 , 
    R_164_12b27118 , 
    R_104d9_120779b8 , 
    R_1ab_f8c2998 , 
    R_23c_13319328 , 
    R_bbdf_133063a8 , 
    R_d3_12659968 , 
    R_cc7b_13a1b128 , 
    R_12ffe_1331cd48 , 
    R_1323e_126561c8 , 
    R_1207f_133190a8 , 
    R_10f99_126549a8 , 
    R_913d_12646b28 , 
    R_c3ee_102f6848 , 
    R_13b12_13a1a728 , 
    R_10a0c_11cdf1c8 , 
    R_13974_13a19008 , 
    R_13602_126635a8 , 
    R_124e1_11cdb668 , 
    R_142d7_12b30d58 , 
    R_14960_105b5598 , 
    R_f86d_120385f8 , 
    R_148a0_12b38ab8 , 
    R_e63f_f8cb9f8 , 
    R_12741_105642d8 , 
    R_684e_1056aa98 , 
    R_13b04_12081558 , 
    R_1453f_11ce2328 , 
    R_148b5_1207f898 , 
    R_1499c_12080658 , 
    R_128e2_12647668 , 
    R_13345_11ce0988 , 
    R_cd4f_102f2f68 , 
    R_13dd3_1204cd38 , 
    R_13ea4_11ce0708 , 
    R_f16b_11cda448 , 
    R_139fe_1153e5b8 , 
    R_12eed_102ee1e8 , 
    R_13479_13306b28 , 
    R_1135b_1056d158 , 
    R_131a5_1153dc58 , 
    R_14744_1264b3a8 , 
    R_144c6_1056d5b8 , 
    R_13109_f8c4798 , 
    R_137bb_10564058 , 
    R_146db_1056a818 , 
    R_119c2_13a1a548 , 
    R_eb5e_1056d018 , 
    R_b0d7_1153e3d8 , 
    R_13b9e_12083038 , 
    R_1116a_13a15868 , 
    R_12a65_10564c38 , 
    R_14969_11cdb2a8 , 
    R_1464d_12075618 , 
    R_e3c5_12080a18 , 
    R_1469c_120511f8 , 
    R_d50f_12663828 , 
    R_137f0_12079358 , 
    R_11593_1207a258 , 
    R_14350_1207d8b8 , 
    R_cbe2_11536a98 , 
    R_110ed_10563d38 , 
    R_1125d_102f86e8 , 
    R_13c09_11ce4268 , 
    R_135fc_13795948 , 
    R_14557_11cdcec8 , 
    R_112_13312248 , 
    R_1fd_133221a8 , 
    R_9e_11539838 , 
    R_143b2_11cddd28 , 
    R_12fec_102efea8 , 
    R_c4d7_13a1f408 , 
    R_1398e_13320bc8 , 
    R_12894_11ce1428 , 
    R_b6f4_102f9ea8 , 
    R_fcb3_12649be8 , 
    R_12375_1207edf8 , 
    R_146b1_102ed248 , 
    R_11b11_11545818 , 
    R_58_13317a28 , 
    R_73_12b3e0f8 , 
    R_bd7c_11ce2be8 , 
    R_12fd8_10565278 , 
    R_14876_12054678 , 
    R_138da_1153dbb8 , 
    R_14825_12647168 , 
    R_14a4d_12646ee8 , 
    R_124_1203edb8 , 
    R_15a_f8c6958 , 
    R_1b5_1331afe8 , 
    R_1eb_12038d78 , 
    R_1475d_11546038 , 
    R_171_105aa5f8 , 
    R_106ea_102f6528 , 
    R_19e_1331e788 , 
    R_11a86_1204ffd8 , 
    R_fad7_102f5ee8 , 
    R_e21e_1056b7b8 , 
    R_12933_11cd7c48 , 
    R_6c_12040938 , 
    R_99_12b27618 , 
    R_1353d_1153d9d8 , 
    R_b283_1330acc8 , 
    R_143ae_13a1cca8 , 
    R_14801_11540c78 , 
    R_149e7_10568298 , 
    R_14708_1203c018 , 
    R_14450_13a17028 , 
    R_128_12b43b98 , 
    R_145_1265aa48 , 
    R_1ca_1265ff48 , 
    R_1e7_12b3d798 , 
    R_7741_13a16128 , 
    R_da39_12b40718 , 
    R_e38d_12651168 , 
    R_12fc4_11544878 , 
    R_145e7_11544058 , 
    R_1465f_105676b8 , 
    R_10fc1_12078638 , 
    R_704f_11ce4da8 , 
    R_13a8d_13318108 , 
    R_145c3_1264da68 , 
    R_faad_13a1fd68 , 
    R_12738_10570678 , 
    R_11935_13a1ff48 , 
    R_11720_1330eaa8 , 
    R_d16a_11ce5de8 , 
    R_13e0d_13a1b4e8 , 
    R_1447d_11ce3a48 , 
    R_152_12b3c4d8 , 
    R_105ba_13306bc8 , 
    R_b1aa_12649468 , 
    R_1bd_12653be8 , 
    R_14a50_13a161c8 , 
    R_13a83_10567a78 , 
    R_123c2_13797108 , 
    R_144b7_13305d68 , 
    R_13814_137926a8 , 
    R_12cbd_13a14328 , 
    R_11bab_120768d8 , 
    R_c07e_13a18b08 , 
    R_142f9_11545e58 , 
    R_1478a_12652928 , 
    R_14a3b_11ce2d28 , 
    R_c3a2_13a19508 , 
    R_aa_126535a8 , 
    R_146e7_10566538 , 
    R_138fb_12082778 , 
    R_13988_133186a8 , 
    R_13c43_1264cca8 , 
    R_14590_132f3b08 , 
    R_110cf_137940e8 , 
    R_13326_12648d88 , 
    R_13153_10567118 , 
    R_1405e_f8c95b8 , 
    R_1051f_13793b48 , 
    R_f518_12075bb8 , 
    R_143a2_12079038 , 
    R_147a8_12657de8 , 
    R_13cb3_102f6fc8 , 
    R_10c3d_f8c5b98 , 
    R_e7ab_1264f7c8 , 
    R_13449_12077378 , 
    R_14403_12b29418 , 
    R_148b2_132fc708 , 
    R_1468f_10562cf8 , 
    R_f7_13309828 , 
    R_13f54_102f4e08 , 
    R_218_12050258 , 
    R_83_1379cd88 , 
    R_12f16_137a0b68 , 
    R_10598_102ead68 , 
    R_10365_12051478 , 
    R_13ab4_13a12ca8 , 
    R_13393_10568a18 , 
    R_13683_1207cf58 , 
    R_13a_105ac2b8 , 
    R_127d5_11cdf268 , 
    R_11917_11ce1248 , 
    R_1d5_1265e468 , 
    R_12e98_1204e778 , 
    R_b3_12655ea8 , 
    R_149cc_10564cd8 , 
    R_134d9_10565f98 , 
    R_fd0b_102ec488 , 
    R_af25_133136a8 , 
    R_11948_12b288d8 , 
    R_149c6_1207b018 , 
    R_14b_12b28a18 , 
    R_1c4_12652e28 , 
    R_10199_13a1f368 , 
    R_80_12055438 , 
    R_10b70_f8cd438 , 
    R_10cdf_115401d8 , 
    R_11a66_1207dc78 , 
    R_132fc_13307708 , 
    R_8c7b_12076b58 , 
    R_1495a_1207a2f8 , 
    R_1201a_10570218 , 
    R_132d6_11ce0348 , 
    R_14963_13304be8 , 
    R_1285e_11545c78 , 
    R_130de_102f58a8 , 
    R_fb5f_13a1e288 , 
    R_13ecf_1207c5f8 , 
    R_1456f_13a1f5e8 , 
    R_ea_1331a9a8 , 
    R_120_12b400d8 , 
    R_13eac_11ce2a08 , 
    R_12568_1056b0d8 , 
    R_e3ba_1207df98 , 
    R_dcf2_12085298 , 
    R_1ef_f8c2cb8 , 
    R_225_12b3a318 , 
    R_f7da_1204e9f8 , 
    R_f857_13a13748 , 
    R_1461a_13301988 , 
    R_146b7_13a15228 , 
    R_1384a_126503a8 , 
    R_c8e7_105b6498 , 
    R_86_137a1a68 , 
    R_a3_126621a8 , 
    R_f862_13a1a908 , 
    R_10ab7_102f7b08 , 
    R_11890_102eb308 , 
    R_df3c_120774b8 , 
    R_1369b_1330c2a8 , 
    R_12e03_132ff368 , 
    R_1356b_102f5da8 , 
    R_10e42_1207e718 , 
    R_10f59_f8c2c18 , 
    R_127b6_12b412f8 , 
    R_120e7_12b44818 , 
    R_12492_1265b9e8 , 
    R_10d12_13792b08 , 
    R_130ae_12044b78 , 
    R_13652_11ce1ce8 , 
    R_117a7_12080fb8 , 
    R_14674_13a13ba8 , 
    R_11306_11540638 , 
    R_d5_126617a8 , 
    R_de_1265ce88 , 
    R_12c_1379b488 , 
    R_135_f8c6f98 , 
    R_1da_12664b88 , 
    R_1e3_1153c498 , 
    R_122dd_13a1b6c8 , 
    R_231_1379a6c8 , 
    R_23a_12660b28 , 
    R_1240e_13a150e8 , 
    R_14686_13a137e8 , 
    R_146c6_f8cf918 , 
    R_13f5b_1207c738 , 
    R_ebb7_102efd68 , 
    R_1447a_105697d8 , 
    R_13c95_12650ee8 , 
    R_11de0_12083cb8 , 
    R_11552_12648c48 , 
    R_11cb2_1207ab18 , 
    R_14849_11ce0028 , 
    R_13f45_13a134c8 , 
    R_13726_12084f78 , 
    R_121f2_102f30a8 , 
    R_ef_1379b0c8 , 
    R_163_12b38a18 , 
    R_1ac_12b29558 , 
    R_220_12b25638 , 
    R_14623_13a12a28 , 
    R_1393a_11ce3408 , 
    R_139ea_11cd8828 , 
    R_cf49_11541718 , 
    R_b889_1056a458 , 
    R_1349f_1204fdf8 , 
    R_170_120440d8 , 
    R_19f_133087e8 , 
    R_a9d8_102f22e8 , 
    R_7d_12660308 , 
    R_1460b_10569a58 , 
    R_11983_13318568 , 
    R_a6e4_13314648 , 
    R_144b1_1207b478 , 
    R_14614_12664f48 , 
    R_139d7_132fda68 , 
    R_ec64_11ce6248 , 
    R_12d32_115454f8 , 
    R_82bb_1204a678 , 
    R_1472c_13a139c8 , 
    R_144f7_10565e58 , 
    R_10dad_12082f98 , 
    R_b05c_1330b4e8 , 
    R_13ef1_105714d8 , 
    R_14635_12b3b038 , 
    R_117b5_1056fdb8 , 
    R_14692_11cdf128 , 
    R_13f_1203dd78 , 
    R_1055c_105672f8 , 
    R_1d0_12040258 , 
    R_13aba_1265cde8 , 
    R_131e1_102f2ec8 , 
    R_eb07_1153ef18 , 
    R_9c9a_1056c578 , 
    R_10605_11545d18 , 
    R_13a97_12079218 , 
    R_1331b_102efc28 , 
    R_14879_11ce58e8 , 
    R_14996_102eb3a8 , 
    R_1405c_11ce34a8 , 
    R_14945_1056e238 , 
    R_b65f_11cdba28 , 
    R_13f3e_13a1e508 , 
    R_dbc0_132fb9e8 , 
    R_1351c_13797068 , 
    R_14804_120788b8 , 
    R_14a0b_133206c8 , 
    R_89_126595a8 , 
    R_13c33_11ce3688 , 
    R_4f_12b44d18 , 
    R_cb5a_12b256d8 , 
    R_13b85_10571258 , 
    R_138f4_1330a9a8 , 
    R_ee1a_1264fae8 , 
    R_10411_102f8828 , 
    R_14331_1056be98 , 
    R_14717_1153a378 , 
    R_94_1330ee68 , 
    R_e5_1153cfd8 , 
    R_22a_12b43698 , 
    R_cba1_13a16e48 , 
    R_129d1_12047978 , 
    R_143d8_11cdc2e8 , 
    R_13070_1264b268 , 
    R_12915_1056d518 , 
    R_12942_11cdd0a8 , 
    R_145a8_12662608 , 
    R_fda2_1264e328 , 
    R_ee25_13a16588 , 
    R_13a1f_11cde2c8 , 
    R_1432d_11cdddc8 , 
    R_13be3_12036bb8 , 
    R_fe10_13a14468 , 
    R_12610_1204bcf8 , 
    R_13701_11cdc608 , 
    R_12597_105711b8 , 
    R_1441d_12035d58 , 
    R_1443c_137979c8 , 
    R_139a7_11ce70a8 , 
    R_13ad3_1056bdf8 , 
    R_143e0_102efcc8 , 
    R_147cc_13315ae8 , 
    R_1444b_11cdad08 , 
    R_12631_12036c58 , 
    R_13dda_102f4fe8 , 
    R_efd_13a14fa8 , 
    R_14954_12054358 , 
    R_1287f_115422f8 , 
    R_1169f_102f8968 , 
    R_13a2b_1264b628 , 
    R_11285_102f9e08 , 
    R_12548_1056ce38 , 
    R_1173e_12649fa8 , 
    R_10b51_13a18a68 , 
    R_148ca_13a18c48 , 
    R_12c82_102f0448 , 
    R_13b79_11543d38 , 
    R_14057_f8cd618 , 
    R_a2e4_1056c618 , 
    R_101e6_1330c7a8 , 
    R_13a56_f8c0a58 , 
    R_d6bc_13a1ca28 , 
    R_4a_1265e648 , 
    R_115_13316c68 , 
    R_1224c_12b3d478 , 
    R_1fa_1265d388 , 
    R_eeda_11cd81e8 , 
    R_1455d_11cd9fe8 , 
    R_1402e_1264dc48 , 
    R_c753_12039098 , 
    R_1283c_13a1da68 , 
    R_aeda_13a1d6a8 , 
    R_14939_1379f448 , 
    R_14a20_13a13e28 , 
    R_13a9d_12081698 , 
    R_117c0_11ce3e08 , 
    R_114e1_132f28e8 , 
    R_1476f_132fb768;
wire n203077 , n203078 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , 
     n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , 
     n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , 
     n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , 
     n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , 
     n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , 
     n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , 
     n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , 
     n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , 
     n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , 
     n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , 
     n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , 
     n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , 
     n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , 
     n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , 
     n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , 
     n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , 
     n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , 
     n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , 
     n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , 
     n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , 
     n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , 
     n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , 
     n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , 
     n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , 
     n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , 
     n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , 
     n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , 
     n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , 
     n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , 
     n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , 
     n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , 
     n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , 
     n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , 
     n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , 
     n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , 
     n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , 
     n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , 
     n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , 
     n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , 
     n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , 
     n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , 
     n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , 
     n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , 
     n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , 
     n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , 
     n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , 
     n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , 
     n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , 
     n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , 
     n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , 
     n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , 
     n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , 
     n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , 
     n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , 
     n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , 
     n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , 
     n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , 
     n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , 
     n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , 
     n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , 
     n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , 
     n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , 
     n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , 
     n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , 
     n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , 
     n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , 
     n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , 
     n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , 
     n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , 
     n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , 
     n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , 
     n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , 
     n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , 
     n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , 
     n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , 
     n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , 
     n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , 
     n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , 
     n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , 
     n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , 
     n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , 
     n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , 
     n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , 
     n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , 
     n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , 
     n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , 
     n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , 
     n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , 
     n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , 
     n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , 
     n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , 
     n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , 
     n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , 
     n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , 
     n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , 
     n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , 
     n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , 
     n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , 
     n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , 
     n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , 
     n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , 
     n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , 
     n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , 
     n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , 
     n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , 
     n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , 
     n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , 
     n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , 
     n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , 
     n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , 
     n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , 
     n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , 
     n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , 
     n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , 
     n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , 
     n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , 
     n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n204252 , n204253 , n204254 , n204255 , 
     n204256 , n204257 , n204258 , n204259 , n204260 , n204261 , n204262 , n204263 , n204264 , n204265 , 
     n204266 , n204267 , n204268 , n204269 , n204270 , n204271 , n204272 , n204273 , n204274 , n204275 , 
     n204276 , n204277 , n204278 , n204279 , n204280 , n204281 , n204282 , n204283 , n204284 , n204285 , 
     n204286 , n204287 , n204288 , n204289 , n204290 , n204291 , n204292 , n204293 , n204294 , n204295 , 
     n204296 , n204297 , n204298 , n204299 , n204300 , n204301 , n204302 , n204303 , n204304 , n204305 , 
     n204306 , n204307 , n204308 , n204309 , n204310 , n204311 , n204312 , n204313 , n204314 , n204315 , 
     n204316 , n204317 , n204318 , n204319 , n204320 , n204321 , n204322 , n204323 , n204324 , n204325 , 
     n204326 , n204327 , n204328 , n204329 , n204330 , n204331 , n204332 , n204333 , n204334 , n204335 , 
     n204336 , n204337 , n204338 , n204339 , n204340 , n204341 , n204342 , n204343 , n204344 , n204345 , 
     n204346 , n204347 , n204348 , n204349 , n204350 , n204351 , n204352 , n204353 , n204354 , n204355 , 
     n204356 , n204357 , n204358 , n204359 , n204360 , n204361 , n204362 , n204363 , n204364 , n204365 , 
     n204366 , n204367 , n204368 , n204369 , n204370 , n204371 , n204372 , n204373 , n204374 , n204375 , 
     n204376 , n204377 , n204378 , n204379 , n204380 , n204381 , n204382 , n204383 , n204384 , n204385 , 
     n204386 , n204387 , n204388 , n204389 , n204390 , n204391 , n204392 , n204393 , n204394 , n204395 , 
     n204396 , n204397 , n204398 , n204399 , n204400 , n204401 , n204402 , n204403 , n204404 , n204405 , 
     n204406 , n204407 , n204408 , n204409 , n204410 , n204411 , n204412 , n204413 , n204414 , n204415 , 
     n204416 , n204417 , n204418 , n204419 , n204420 , n204421 , n204422 , n204423 , n204424 , n204425 , 
     n204426 , n204427 , n204428 , n204429 , n204430 , n204431 , n204432 , n204433 , n204434 , n204435 , 
     n204436 , n204437 , n204438 , n204439 , n204440 , n204441 , n204442 , n204443 , n204444 , n204445 , 
     n204446 , n204447 , n204448 , n204449 , n204450 , n204451 , n204452 , n204453 , n204454 , n204455 , 
     n204456 , n204457 , n204458 , n204459 , n204460 , n204461 , n204462 , n204463 , n204464 , n204465 , 
     n204466 , n204467 , n204468 , n204469 , n204470 , n204471 , n204472 , n204473 , n204474 , n204475 , 
     n204476 , n204477 , n204478 , n204479 , n204480 , n204481 , n204482 , n204483 , n204484 , n204485 , 
     n204486 , n204487 , n204488 , n204489 , n204490 , n204491 , n204492 , n204493 , n204494 , n204495 , 
     n204496 , n204497 , n204498 , n204499 , n204500 , n204501 , n204502 , n204503 , n204504 , n204505 , 
     n204506 , n204507 , n204508 , n204509 , n204510 , n204511 , n204512 , n204513 , n204514 , n204515 , 
     n204516 , n204517 , n204518 , n204519 , n204520 , n204521 , n204522 , n204523 , n204524 , n204525 , 
     n204526 , n204527 , n204528 , n204529 , n204530 , n204531 , n204532 , n204533 , n204534 , n204535 , 
     n204536 , n204537 , n204538 , n204539 , n204540 , n204541 , n204542 , n204543 , n204544 , n204545 , 
     n204546 , n204547 , n204548 , n204549 , n204550 , n204551 , n204552 , n204553 , n204554 , n204555 , 
     n204556 , n204557 , n204558 , n204559 , n204560 , n204561 , n204562 , n204563 , n204564 , n204565 , 
     n204566 , n204567 , n204568 , n204569 , n204570 , n204571 , n204572 , n204573 , n204574 , n204575 , 
     n204576 , n204577 , n204578 , n204579 , n204580 , n204581 , n204582 , n204583 , n204584 , n204585 , 
     n204586 , n204587 , n204588 , n204589 , n204590 , n204591 , n204592 , n204593 , n204594 , n204595 , 
     n204596 , n204597 , n204598 , n204599 , n204600 , n204601 , n204602 , n204603 , n204604 , n204605 , 
     n204606 , n204607 , n204608 , n204609 , n204610 , n204611 , n204612 , n204613 , n204614 , n204615 , 
     n204616 , n204617 , n204618 , n204619 , n204620 , n204621 , n204622 , n204623 , n204624 , n204625 , 
     n204626 , n204627 , n204628 , n204629 , n204630 , n204631 , n204632 , n204633 , n204634 , n204635 , 
     n204636 , n204637 , n204638 , n204639 , n204640 , n204641 , n204642 , n204643 , n204644 , n204645 , 
     n204646 , n204647 , n204648 , n204649 , n204650 , n204651 , n204652 , n204653 , n204654 , n204655 , 
     n204656 , n204657 , n204658 , n204659 , n204660 , n204661 , n204662 , n204663 , n204664 , n204665 , 
     n204666 , n204667 , n204668 , n204669 , n204670 , n204671 , n204672 , n204673 , n204674 , n204675 , 
     n204676 , n204677 , n204678 , n204679 , n204680 , n204681 , n204682 , n204683 , n204684 , n204685 , 
     n204686 , n204687 , n204688 , n204689 , n204690 , n204691 , n204692 , n204693 , n204694 , n204695 , 
     n204696 , n204697 , n204698 , n204699 , n204700 , n204701 , n204702 , n204703 , n204704 , n204705 , 
     n204706 , n204707 , n204708 , n204709 , n204710 , n204711 , n204712 , n204713 , n204714 , n204715 , 
     n204716 , n204717 , n204718 , n204719 , n204720 , n204721 , n204722 , n204723 , n204724 , n204725 , 
     n204726 , n204727 , n204728 , n204729 , n204730 , n204731 , n204732 , n204733 , n204734 , n204735 , 
     n204736 , n204737 , n204738 , n204739 , n204740 , n204741 , n204742 , n204743 , n204744 , n204745 , 
     n204746 , n204747 , n204748 , n204749 , n204750 , n204751 , n204752 , n204753 , n204754 , n204755 , 
     n204756 , n204757 , n204758 , n204759 , n204760 , n204761 , n204762 , n204763 , n204764 , n204765 , 
     n204766 , n204767 , n204768 , n204769 , n204770 , n204771 , n204772 , n204773 , n204774 , n204775 , 
     n204776 , n204777 , n204778 , n204779 , n204780 , n204781 , n204782 , n204783 , n204784 , n204785 , 
     n204786 , n204787 , n204788 , n204789 , n204790 , n204791 , n204792 , n204793 , n204794 , n204795 , 
     n204796 , n204797 , n204798 , n204799 , n204800 , n204801 , n204802 , n204803 , n204804 , n204805 , 
     n204806 , n204807 , n204808 , n204809 , n204810 , n204811 , n204812 , n204813 , n204814 , n204815 , 
     n204816 , n204817 , n204818 , n204819 , n204820 , n204821 , n204822 , n204823 , n204824 , n204825 , 
     n204826 , n204827 , n204828 , n204829 , n204830 , n204831 , n204832 , n204833 , n204834 , n204835 , 
     n204836 , n204837 , n204838 , n204839 , n204840 , n204841 , n204842 , n204843 , n204844 , n204845 , 
     n204846 , n204847 , n204848 , n204849 , n204850 , n204851 , n204852 , n204853 , n204854 , n204855 , 
     n204856 , n204857 , n204858 , n204859 , n204860 , n204861 , n204862 , n204863 , n204864 , n204865 , 
     n204866 , n204867 , n204868 , n204869 , n204870 , n204871 , n204872 , n204873 , n204874 , n204875 , 
     n204876 , n204877 , n204878 , n204879 , n204880 , n204881 , n204882 , n204883 , n204884 , n204885 , 
     n204886 , n204887 , n204888 , n204889 , n204890 , n204891 , n204892 , n204893 , n204894 , n204895 , 
     n204896 , n204897 , n204898 , n204899 , n204900 , n204901 , n204902 , n204903 , n204904 , n204905 , 
     n204906 , n204907 , n204908 , n204909 , n204910 , n204911 , n204912 , n204913 , n204914 , n204915 , 
     n204916 , n204917 , n204918 , n204919 , n204920 , n204921 , n204922 , n204923 , n204924 , n204925 , 
     n204926 , n204927 , n204928 , n204929 , n204930 , n204931 , n204932 , n204933 , n204934 , n204935 , 
     n204936 , n204937 , n204938 , n204939 , n204940 , n204941 , n204942 , n204943 , n204944 , n204945 , 
     n204946 , n204947 , n204948 , n204949 , n204950 , n204951 , n204952 , n204953 , n204954 , n204955 , 
     n204956 , n204957 , n204958 , n204959 , n204960 , n204961 , n204962 , n204963 , n204964 , n204965 , 
     n204966 , n204967 , n204968 , n204969 , n204970 , n204971 , n204972 , n204973 , n204974 , n204975 , 
     n204976 , n204977 , n204978 , n204979 , n204980 , n204981 , n204982 , n204983 , n204984 , n204985 , 
     n204986 , n204987 , n204988 , n204989 , n204990 , n204991 , n204992 , n204993 , n204994 , n204995 , 
     n204996 , n204997 , n204998 , n204999 , n205000 , n205001 , n205002 , n205003 , n205004 , n205005 , 
     n205006 , n205007 , n205008 , n205009 , n205010 , n205011 , n205012 , n205013 , n205014 , n205015 , 
     n205016 , n205017 , n205018 , n205019 , n205020 , n205021 , n205022 , n205023 , n205024 , n205025 , 
     n205026 , n205027 , n205028 , n205029 , n205030 , n205031 , n205032 , n205033 , n205034 , n205035 , 
     n205036 , n205037 , n205038 , n205039 , n205040 , n205041 , n205042 , n205043 , n205044 , n205045 , 
     n205046 , n205047 , n205048 , n205049 , n205050 , n205051 , n205052 , n205053 , n205054 , n205055 , 
     n205056 , n205057 , n205058 , n205059 , n205060 , n205061 , n205062 , n205063 , n205064 , n205065 , 
     n205066 , n205067 , n205068 , n205069 , n205070 , n205071 , n205072 , n205073 , n205074 , n205075 , 
     n205076 , n205077 , n205078 , n205079 , n205080 , n205081 , n205082 , n205083 , n205084 , n205085 , 
     n205086 , n205087 , n205088 , n205089 , n205090 , n205091 , n205092 , n205093 , n205094 , n205095 , 
     n205096 , n205097 , n205098 , n205099 , n205100 , n205101 , n205102 , n205103 , n205104 , n205105 , 
     n205106 , n205107 , n205108 , n205109 , n205110 , n205111 , n205112 , n205113 , n205114 , n205115 , 
     n205116 , n205117 , n205118 , n205119 , n205120 , n205121 , n205122 , n205123 , n205124 , n205125 , 
     n205126 , n205127 , n205128 , n205129 , n205130 , n205131 , n205132 , n205133 , n205134 , n205135 , 
     n205136 , n205137 , n205138 , n205139 , n205140 , n205141 , n205142 , n205143 , n205144 , n205145 , 
     n205146 , n205147 , n205148 , n205149 , n205150 , n205151 , n205152 , n205153 , n205154 , n205155 , 
     n205156 , n205157 , n205158 , n205159 , n205160 , n205161 , n205162 , n205163 , n205164 , n205165 , 
     n205166 , n205167 , n205168 , n205169 , n205170 , n205171 , n205172 , n205173 , n205174 , n205175 , 
     n205176 , n205177 , n205178 , n205179 , n205180 , n205181 , n205182 , n205183 , n205184 , n205185 , 
     n205186 , n205187 , n205188 , n205189 , n205190 , n205191 , n205192 , n205193 , n205194 , n205195 , 
     n205196 , n205197 , n205198 , n205199 , n205200 , n205201 , n205202 , n205203 , n205204 , n205205 , 
     n205206 , n205207 , n205208 , n205209 , n205210 , n205211 , n205212 , n205213 , n205214 , n205215 , 
     n205216 , n205217 , n205218 , n205219 , n205220 , n205221 , n205222 , n205223 , n205224 , n205225 , 
     n205226 , n205227 , n205228 , n205229 , n205230 , n205231 , n205232 , n205233 , n205234 , n205235 , 
     n205236 , n205237 , n205238 , n205239 , n205240 , n205241 , n205242 , n205243 , n205244 , n205245 , 
     n205246 , n205247 , n205248 , n205249 , n205250 , n205251 , n205252 , n205253 , n205254 , n205255 , 
     n205256 , n205257 , n205258 , n205259 , n205260 , n205261 , n205262 , n205263 , n205264 , n205265 , 
     n205266 , n205267 , n205268 , n205269 , n205270 , n205271 , n205272 , n205273 , n205274 , n205275 , 
     n205276 , n205277 , n205278 , n205279 , n205280 , n205281 , n205282 , n205283 , n205284 , n205285 , 
     n205286 , n205287 , n205288 , n205289 , n205290 , n205291 , n205292 , n205293 , n205294 , n205295 , 
     n205296 , n205297 , n205298 , n205299 , n205300 , n205301 , n205302 , n205303 , n205304 , n205305 , 
     n205306 , n205307 , n205308 , n205309 , n205310 , n205311 , n205312 , n205313 , n205314 , n205315 , 
     n205316 , n205317 , n205318 , n205319 , n205320 , n205321 , n205322 , n205323 , n205324 , n205325 , 
     n205326 , n205327 , n205328 , n205329 , n205330 , n205331 , n205332 , n205333 , n205334 , n205335 , 
     n205336 , n205337 , n205338 , n205339 , n205340 , n205341 , n205342 , n205343 , n205344 , n205345 , 
     n205346 , n205347 , n205348 , n205349 , n205350 , n205351 , n205352 , n205353 , n205354 , n205355 , 
     n205356 , n205357 , n205358 , n205359 , n205360 , n205361 , n205362 , n205363 , n205364 , n205365 , 
     n205366 , n205367 , n205368 , n205369 , n205370 , n205371 , n205372 , n205373 , n205374 , n205375 , 
     n205376 , n205377 , n205378 , n205379 , n205380 , n205381 , n205382 , n205383 , n205384 , n205385 , 
     n205386 , n205387 , n205388 , n205389 , n205390 , n205391 , n205392 , n205393 , n205394 , n205395 , 
     n205396 , n205397 , n205398 , n205399 , n205400 , n205401 , n205402 , n205403 , n205404 , n205405 , 
     n205406 , n205407 , n205408 , n205409 , n205410 , n205411 , n205412 , n205413 , n205414 , n205415 , 
     n205416 , n205417 , n205418 , n205419 , n205420 , n205421 , n205422 , n205423 , n205424 , n205425 , 
     n205426 , n205427 , n27667 , n27668 , n27669 , n27670 , n205432 , n205433 , n205434 , n205435 , 
     n205436 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n205445 , 
     n205446 , n27686 , n27687 , n27688 , n27689 , n205451 , n27691 , n205453 , n27693 , n27694 , 
     n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n205464 , n27704 , 
     n205466 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , 
     n205476 , n27716 , n205478 , n27718 , n205480 , n27720 , n27721 , n27722 , n27723 , n27724 , 
     n27725 , n27726 , n27727 , n27728 , n205490 , n27730 , n205492 , n27732 , n27733 , n27734 , 
     n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n205504 , n27744 , 
     n205506 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , 
     n205516 , n27756 , n205518 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , 
     n27765 , n27766 , n27767 , n27768 , n27769 , n205531 , n27771 , n205533 , n27773 , n27774 , 
     n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n205543 , n27783 , n205545 , 
     n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , 
     n27795 , n27796 , n27797 , n205559 , n27799 , n205561 , n27801 , n27802 , n27803 , n27804 , 
     n27805 , n27806 , n27807 , n27808 , n27809 , n205571 , n27811 , n205573 , n27813 , n27814 , 
     n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n205583 , n27823 , n205585 , 
     n27825 , n205587 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , 
     n27835 , n205597 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , 
     n27845 , n27846 , n27847 , n27848 , n205610 , n27850 , n205612 , n27852 , n27853 , n27854 , 
     n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n205622 , n27862 , n205624 , n27864 , 
     n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , 
     n27875 , n27876 , n205638 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , 
     n27885 , n27886 , n27887 , n205649 , n27889 , n205651 , n27891 , n27892 , n27893 , n27894 , 
     n27895 , n27896 , n27897 , n27898 , n27899 , n205661 , n27901 , n205663 , n27903 , n27904 , 
     n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n205673 , n27913 , n205675 , 
     n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , 
     n205686 , n27926 , n205688 , n27928 , n205690 , n27930 , n27931 , n27932 , n27933 , n27934 , 
     n27935 , n27936 , n27937 , n27938 , n205700 , n27940 , n205702 , n27942 , n27943 , n27944 , 
     n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , 
     n205716 , n27956 , n205718 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , 
     n27965 , n27966 , n205728 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , 
     n27975 , n27976 , n27977 , n205739 , n27979 , n205741 , n27981 , n205743 , n27983 , n27984 , 
     n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n205753 , n27993 , n205755 , 
     n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , 
     n205766 , n28006 , n205768 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , 
     n28015 , n28016 , n28017 , n205779 , n28019 , n205781 , n28021 , n28022 , n28023 , n28024 , 
     n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n205795 , 
     n28035 , n205797 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , 
     n28045 , n205807 , n28047 , n205809 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , 
     n28055 , n28056 , n28057 , n205819 , n28059 , n205821 , n28061 , n205823 , n28063 , n28064 , 
     n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n205833 , n28073 , n205835 , 
     n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , 
     n205846 , n28086 , n205848 , n28088 , n205850 , n28090 , n28091 , n28092 , n28093 , n28094 , 
     n28095 , n28096 , n28097 , n28098 , n205860 , n28100 , n28101 , n28102 , n28103 , n28104 , 
     n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n205875 , 
     n28115 , n205877 , n28117 , n205879 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , 
     n28125 , n28126 , n28127 , n205889 , n28129 , n205891 , n28131 , n28132 , n28133 , n28134 , 
     n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n205902 , n28142 , n28143 , n28144 , 
     n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n205912 , n28152 , n205914 , n28154 , 
     n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , 
     n205926 , n28166 , n205928 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , 
     n28175 , n28176 , n205938 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , 
     n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n205952 , n28192 , n205954 , n28194 , 
     n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n205964 , n28204 , 
     n205966 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , 
     n28215 , n205977 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , 
     n28225 , n28226 , n205988 , n28228 , n205990 , n28230 , n28231 , n28232 , n28233 , n28234 , 
     n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n206002 , n28242 , n206004 , n28244 , 
     n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n206014 , n28254 , 
     n206016 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , 
     n28265 , n28266 , n28267 , n206029 , n28269 , n206031 , n28271 , n206033 , n28273 , n28274 , 
     n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n206043 , n28283 , n206045 , 
     n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , 
     n206056 , n28296 , n206058 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , 
     n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , 
     n28315 , n28316 , n28317 , n206079 , n28319 , n206081 , n28321 , n28322 , n28323 , n28324 , 
     n28325 , n28326 , n28327 , n28328 , n28329 , n206091 , n28331 , n206093 , n28333 , n28334 , 
     n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , 
     n206106 , n28346 , n206108 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , 
     n28355 , n28356 , n28357 , n206119 , n28359 , n206121 , n28361 , n28362 , n28363 , n28364 , 
     n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n206132 , n28372 , n206134 , n28374 , 
     n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n206144 , n28384 , 
     n206146 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , 
     n28395 , n28396 , n206158 , n28398 , n206160 , n28400 , n28401 , n28402 , n28403 , n28404 , 
     n28405 , n28406 , n28407 , n28408 , n206170 , n28410 , n206172 , n28412 , n28413 , n28414 , 
     n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n206185 , 
     n28425 , n28426 , n28427 , n28428 , n206190 , n28430 , n206192 , n28432 , n28433 , n28434 , 
     n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n206202 , n28442 , n206204 , n28444 , 
     n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , 
     n206216 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , 
     n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n206232 , n28472 , n206234 , n28474 , 
     n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , 
     n206246 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , 
     n28495 , n206257 , n28497 , n206259 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , 
     n28505 , n28506 , n28507 , n28508 , n28509 , n206271 , n28511 , n206273 , n28513 , n28514 , 
     n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , 
     n206286 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , 
     n28535 , n206297 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , 
     n28545 , n206307 , n28547 , n206309 , n28549 , n206311 , n28551 , n28552 , n28553 , n28554 , 
     n28555 , n28556 , n28557 , n28558 , n28559 , n206321 , n28561 , n206323 , n28563 , n28564 , 
     n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n206335 , 
     n28575 , n206337 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , 
     n28585 , n206347 , n28587 , n206349 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , 
     n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , 
     n28605 , n28606 , n28607 , n206369 , n28609 , n206371 , n28611 , n28612 , n28613 , n28614 , 
     n28615 , n28616 , n28617 , n28618 , n28619 , n206381 , n28621 , n28622 , n28623 , n28624 , 
     n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , 
     n28635 , n206397 , n28637 , n206399 , n28639 , n206401 , n28641 , n28642 , n28643 , n28644 , 
     n28645 , n28646 , n28647 , n28648 , n28649 , n206411 , n28651 , n206413 , n28653 , n28654 , 
     n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n206425 , 
     n28665 , n206427 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , 
     n28675 , n206437 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , 
     n28685 , n28686 , n28687 , n28688 , n28689 , n206451 , n28691 , n28692 , n206454 , n28694 , 
     n206456 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , 
     n206466 , n28706 , n206468 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , 
     n28715 , n28716 , n28717 , n206479 , n28719 , n206481 , n28721 , n28722 , n28723 , n28724 , 
     n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n206493 , n28733 , n206495 , 
     n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , 
     n28745 , n28746 , n28747 , n206509 , n28749 , n206511 , n28751 , n206513 , n28753 , n28754 , 
     n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n206523 , n28763 , n206525 , 
     n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n206535 , 
     n28775 , n206537 , n28777 , n206539 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , 
     n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n206552 , n28792 , n206554 , n28794 , 
     n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n206564 , n28804 , 
     n206566 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , 
     n28815 , n28816 , n28817 , n28818 , n28819 , n206581 , n28821 , n28822 , n28823 , n28824 , 
     n28825 , n28826 , n28827 , n28828 , n28829 , n206591 , n28831 , n206593 , n28833 , n28834 , 
     n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n206605 , 
     n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , 
     n28855 , n28856 , n206618 , n28858 , n206620 , n28860 , n28861 , n28862 , n28863 , n28864 , 
     n28865 , n28866 , n28867 , n28868 , n206630 , n28870 , n206632 , n28872 , n28873 , n28874 , 
     n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n206645 , 
     n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , 
     n206656 , n28896 , n206658 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , 
     n28905 , n28906 , n28907 , n206669 , n28909 , n206671 , n28911 , n28912 , n28913 , n28914 , 
     n28915 , n28916 , n28917 , n28918 , n28919 , n206681 , n28921 , n206683 , n28923 , n28924 , 
     n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , 
     n28935 , n28936 , n28937 , n28938 , n28939 , n206701 , n28941 , n28942 , n28943 , n28944 , 
     n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , 
     n28955 , n28956 , n28957 , n28958 , n28959 , n206721 , n28961 , n206723 , n28963 , n28964 , 
     n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , 
     n206736 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , 
     n28985 , n206747 , n28987 , n206749 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , 
     n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n206763 , n29003 , n206765 , 
     n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , 
     n29015 , n206777 , n29017 , n206779 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , 
     n29025 , n29026 , n29027 , n206789 , n29029 , n206791 , n29031 , n29032 , n29033 , n29034 , 
     n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n206803 , n29043 , n206805 , 
     n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n206815 , 
     n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , 
     n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n206832 , n29072 , n29073 , n29074 , 
     n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , 
     n206846 , n29086 , n206848 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , 
     n29095 , n206857 , n29097 , n206859 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , 
     n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n206875 , 
     n29115 , n206877 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , 
     n29125 , n206887 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , 
     n29135 , n29136 , n29137 , n29138 , n206900 , n29140 , n206902 , n29142 , n29143 , n29144 , 
     n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n206914 , n29154 , 
     n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , 
     n29165 , n29166 , n206928 , n29168 , n206930 , n29170 , n29171 , n29172 , n29173 , n29174 , 
     n29175 , n29176 , n29177 , n29178 , n206940 , n29180 , n206942 , n29182 , n29183 , n29184 , 
     n29185 , n29186 , n29187 , n29188 , n29189 , n206951 , n29191 , n206953 , n29193 , n29194 , 
     n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n206963 , n29203 , n206965 , 
     n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , 
     n206976 , n29216 , n206978 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , 
     n29225 , n29226 , n206988 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , 
     n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n207002 , n29242 , n29243 , n29244 , 
     n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n207012 , n29252 , n29253 , n29254 , 
     n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n207023 , n29263 , n207025 , 
     n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , 
     n29275 , n29276 , n29277 , n29278 , n207040 , n29280 , n29281 , n207043 , n29283 , n207045 , 
     n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , 
     n29295 , n29296 , n29297 , n207059 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , 
     n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n207072 , n29312 , n207074 , n29314 , 
     n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n207084 , n29324 , 
     n207086 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , 
     n29335 , n29336 , n207098 , n29338 , n207100 , n29340 , n29341 , n29342 , n29343 , n29344 , 
     n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n207114 , n29354 , 
     n207116 , n29356 , n207118 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , 
     n29365 , n29366 , n207128 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , 
     n29375 , n29376 , n29377 , n207139 , n29379 , n207141 , n29381 , n29382 , n29383 , n29384 , 
     n29385 , n29386 , n29387 , n29388 , n29389 , n207151 , n29391 , n207153 , n29393 , n29394 , 
     n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n207164 , n29404 , 
     n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n207173 , n29413 , n207175 , 
     n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , 
     n29425 , n29426 , n29427 , n29428 , n207190 , n29430 , n207192 , n29432 , n29433 , n29434 , 
     n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n207202 , n29442 , n29443 , n29444 , 
     n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n207214 , n29454 , 
     n207216 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , 
     n207226 , n29466 , n207228 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , 
     n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n207242 , n29482 , n207244 , n29484 , 
     n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n207254 , n29494 , 
     n207256 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , 
     n29505 , n29506 , n29507 , n29508 , n29509 , n207271 , n29511 , n207273 , n29513 , n29514 , 
     n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n207285 , 
     n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , 
     n207296 , n29536 , n207298 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , 
     n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n207313 , n29553 , n207315 , 
     n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n207325 , 
     n29565 , n207327 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , 
     n29575 , n29576 , n207338 , n29578 , n207340 , n29580 , n29581 , n29582 , n29583 , n29584 , 
     n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n207355 , 
     n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , 
     n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , 
     n207376 , n207377 , n29617 , n29618 , n207380 , n29620 , n207382 , n29622 , n29623 , n29624 , 
     n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n207392 , n29632 , n207394 , n29634 , 
     n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , 
     n29645 , n207407 , n29647 , n207409 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , 
     n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n207422 , n29662 , n29663 , n29664 , 
     n29665 , n29666 , n29667 , n29668 , n207430 , n29670 , n29671 , n29672 , n29673 , n29674 , 
     n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , 
     n207446 , n29686 , n207448 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , 
     n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n207464 , n29704 , 
     n207466 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , 
     n29715 , n207477 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , 
     n29725 , n29726 , n29727 , n29728 , n29729 , n207491 , n29731 , n207493 , n29733 , n207495 , 
     n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n207504 , n29744 , 
     n207506 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , 
     n207516 , n29756 , n29757 , n207519 , n29759 , n207521 , n29761 , n29762 , n29763 , n29764 , 
     n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n207533 , n29773 , n207535 , 
     n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n207545 , 
     n29785 , n207547 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , 
     n29795 , n29796 , n29797 , n29798 , n207560 , n29800 , n29801 , n29802 , n207564 , n29804 , 
     n29805 , n207567 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , 
     n29815 , n29816 , n29817 , n207579 , n29819 , n207581 , n29821 , n29822 , n29823 , n29824 , 
     n29825 , n29826 , n29827 , n29828 , n29829 , n207591 , n29831 , n207593 , n29833 , n29834 , 
     n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , 
     n29845 , n207607 , n29847 , n207609 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , 
     n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n207625 , 
     n29865 , n207627 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , 
     n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , 
     n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , 
     n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n207662 , n29902 , n207664 , n29904 , 
     n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n207675 , 
     n29915 , n207677 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , 
     n29925 , n207687 , n29927 , n207689 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , 
     n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n207704 , n29944 , 
     n207706 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , 
     n207716 , n29956 , n207718 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , 
     n29965 , n29966 , n207728 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , 
     n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , 
     n29985 , n207747 , n29987 , n207749 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , 
     n29995 , n29996 , n29997 , n207759 , n29999 , n207761 , n30001 , n30002 , n30003 , n30004 , 
     n30005 , n30006 , n30007 , n30008 , n30009 , n207771 , n30011 , n30012 , n30013 , n30014 , 
     n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n207783 , n30023 , n207785 , 
     n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , 
     n207796 , n30036 , n207798 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , 
     n30045 , n207807 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , 
     n30055 , n30056 , n207818 , n30058 , n207820 , n30060 , n30061 , n30062 , n30063 , n30064 , 
     n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , 
     n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n207842 , n30082 , n207844 , n30084 , 
     n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n207853 , n30093 , n207855 , 
     n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , 
     n207866 , n30106 , n207868 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , 
     n30115 , n30116 , n207878 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , 
     n30125 , n30126 , n30127 , n30128 , n30129 , n207891 , n30131 , n207893 , n30133 , n30134 , 
     n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n207903 , n30143 , n207905 , 
     n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , 
     n30155 , n30156 , n207918 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , 
     n30165 , n30166 , n30167 , n30168 , n207930 , n30170 , n207932 , n30172 , n30173 , n30174 , 
     n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n207942 , n30182 , n207944 , n30184 , 
     n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , 
     n30195 , n30196 , n30197 , n30198 , n207960 , n30200 , n207962 , n30202 , n30203 , n30204 , 
     n30205 , n30206 , n30207 , n30208 , n30209 , n207971 , n30211 , n30212 , n30213 , n30214 , 
     n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , 
     n207986 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , 
     n30235 , n207997 , n30237 , n207999 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , 
     n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , 
     n30255 , n208017 , n30257 , n30258 , n30259 , n30260 , n30261 , n208023 , n30263 , n208025 , 
     n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n208035 , 
     n30275 , n208037 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , 
     n30285 , n208047 , n30287 , n208049 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , 
     n30295 , n30296 , n208058 , n30298 , n208060 , n30300 , n30301 , n30302 , n30303 , n30304 , 
     n30305 , n30306 , n30307 , n30308 , n30309 , n208071 , n30311 , n208073 , n30313 , n208075 , 
     n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n208085 , 
     n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , 
     n30335 , n30336 , n30337 , n30338 , n208100 , n30340 , n208102 , n30342 , n30343 , n30344 , 
     n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , 
     n208116 , n30356 , n208118 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , 
     n30365 , n30366 , n208128 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , 
     n30375 , n30376 , n30377 , n30378 , n30379 , n208141 , n30381 , n208143 , n30383 , n30384 , 
     n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n208154 , n30394 , 
     n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n208165 , 
     n30405 , n208167 , n30407 , n208169 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , 
     n30415 , n30416 , n30417 , n208179 , n30419 , n208181 , n30421 , n30422 , n30423 , n30424 , 
     n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , 
     n208196 , n30436 , n208198 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , 
     n30445 , n30446 , n30447 , n30448 , n208210 , n30450 , n208212 , n30452 , n30453 , n30454 , 
     n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , 
     n30465 , n208227 , n30467 , n208229 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , 
     n30475 , n30476 , n30477 , n208239 , n30479 , n208241 , n30481 , n30482 , n30483 , n30484 , 
     n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , 
     n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n208263 , n30503 , n208265 , 
     n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n208274 , n30514 , 
     n208276 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , 
     n30525 , n30526 , n30527 , n208289 , n30529 , n208291 , n30531 , n30532 , n30533 , n30534 , 
     n30535 , n30536 , n30537 , n30538 , n30539 , n208301 , n30541 , n208303 , n30543 , n30544 , 
     n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , 
     n30555 , n30556 , n30557 , n30558 , n208320 , n30560 , n30561 , n30562 , n30563 , n30564 , 
     n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , 
     n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , 
     n30585 , n30586 , n30587 , n208349 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , 
     n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , 
     n30605 , n30606 , n30607 , n30608 , n208370 , n30610 , n30611 , n30612 , n30613 , n30614 , 
     n30615 , n30616 , n30617 , n30618 , n208380 , n30620 , n208382 , n30622 , n30623 , n30624 , 
     n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , 
     n208396 , n30636 , n208398 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , 
     n30645 , n208407 , n30647 , n208409 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , 
     n30655 , n30656 , n30657 , n208419 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , 
     n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , 
     n30675 , n30676 , n30677 , n30678 , n30679 , n208441 , n30681 , n208443 , n30683 , n208445 , 
     n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , 
     n30695 , n30696 , n30697 , n208459 , n30699 , n208461 , n30701 , n30702 , n30703 , n30704 , 
     n30705 , n30706 , n30707 , n30708 , n208470 , n30710 , n30711 , n30712 , n30713 , n30714 , 
     n30715 , n30716 , n30717 , n30718 , n30719 , n208481 , n30721 , n30722 , n30723 , n30724 , 
     n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , 
     n30735 , n208497 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , 
     n208506 , n208507 , n30747 , n30748 , n30749 , n208511 , n30751 , n208513 , n30753 , n30754 , 
     n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , 
     n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n208533 , n30773 , n208535 , 
     n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n208545 , 
     n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n208553 , n30793 , n30794 , 
     n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n208565 , 
     n30805 , n208567 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , 
     n30815 , n208577 , n30817 , n208579 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , 
     n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , 
     n208596 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , 
     n30845 , n30846 , n30847 , n30848 , n208610 , n30850 , n208612 , n30852 , n30853 , n30854 , 
     n30855 , n30856 , n30857 , n30858 , n30859 , n208621 , n30861 , n208623 , n30863 , n30864 , 
     n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , 
     n208636 , n30876 , n30877 , n30878 , n30879 , n208641 , n30881 , n208643 , n30883 , n30884 , 
     n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n208653 , n30893 , n208655 , 
     n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , 
     n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n208672 , n30912 , n30913 , n30914 , 
     n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , 
     n30925 , n208687 , n30927 , n208689 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , 
     n30935 , n30936 , n30937 , n208699 , n30939 , n208701 , n30941 , n30942 , n30943 , n30944 , 
     n30945 , n30946 , n30947 , n30948 , n208710 , n30950 , n30951 , n30952 , n30953 , n30954 , 
     n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n208725 , 
     n30965 , n208727 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , 
     n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , 
     n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n208753 , n30993 , n208755 , 
     n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , 
     n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , 
     n208776 , n31016 , n208778 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , 
     n31025 , n31026 , n31027 , n31028 , n208790 , n31030 , n208792 , n31032 , n31033 , n31034 , 
     n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , 
     n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , 
     n31055 , n208817 , n31057 , n208819 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , 
     n31065 , n31066 , n31067 , n208829 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , 
     n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n208843 , n31083 , n31084 , 
     n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n208853 , n31093 , n208855 , 
     n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , 
     n31105 , n208867 , n31107 , n208869 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , 
     n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n208883 , n31123 , n208885 , 
     n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , 
     n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n208904 , n31144 , 
     n208906 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , 
     n208916 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , 
     n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n208934 , n31174 , 
     n208936 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n208944 , n31184 , 
     n208946 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , 
     n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , 
     n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , 
     n31215 , n31216 , n31217 , n31218 , n208980 , n31220 , n208982 , n31222 , n31223 , n31224 , 
     n31225 , n31226 , n31227 , n31228 , n31229 , n208991 , n31231 , n31232 , n31233 , n31234 , 
     n31235 , n31236 , n31237 , n208999 , n31239 , n209001 , n31241 , n31242 , n31243 , n31244 , 
     n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , 
     n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , 
     n31265 , n31266 , n31267 , n31268 , n31269 , n209031 , n31271 , n209033 , n31273 , n31274 , 
     n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n209045 , 
     n31285 , n209047 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , 
     n31295 , n31296 , n31297 , n31298 , n31299 , n209061 , n31301 , n209063 , n31303 , n31304 , 
     n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , 
     n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , 
     n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , 
     n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , 
     n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n209114 , n31354 , 
     n31355 , n31356 , n31357 , n209119 , n31359 , n209121 , n31361 , n31362 , n31363 , n31364 , 
     n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , 
     n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n209145 , 
     n209146 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n209153 , n31393 , n31394 , 
     n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , 
     n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , 
     n209176 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , 
     n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , 
     n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , 
     n31445 , n209207 , n31447 , n209209 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , 
     n31455 , n209217 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , 
     n31465 , n31466 , n209228 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , 
     n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n209242 , n31482 , n31483 , n31484 , 
     n31485 , n31486 , n31487 , n31488 , n31489 , n209251 , n31491 , n31492 , n31493 , n31494 , 
     n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , 
     n31505 , n31506 , n31507 , n31508 , n209270 , n31510 , n31511 , n31512 , n31513 , n31514 , 
     n31515 , n31516 , n31517 , n31518 , n209280 , n31520 , n209282 , n31522 , n31523 , n31524 , 
     n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , 
     n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n209302 , n31542 , n31543 , n31544 , 
     n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n209312 , n31552 , n31553 , n31554 , 
     n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , 
     n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n209335 , 
     n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , 
     n31585 , n209347 , n31587 , n209349 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , 
     n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n209363 , n31603 , n209365 , 
     n31605 , n209367 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , 
     n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n209385 , 
     n31625 , n31626 , n209388 , n31628 , n209390 , n31630 , n31631 , n31632 , n31633 , n31634 , 
     n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , 
     n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , 
     n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , 
     n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n209435 , 
     n31675 , n209437 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , 
     n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , 
     n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , 
     n209466 , n31706 , n209468 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , 
     n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , 
     n31725 , n31726 , n31727 , n31728 , n209490 , n31730 , n31731 , n31732 , n31733 , n31734 , 
     n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n209502 , n31742 , n209504 , n31744 , 
     n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , 
     n209516 , n31756 , n209518 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , 
     n31765 , n31766 , n209528 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , 
     n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , 
     n209546 , n31786 , n209548 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , 
     n31795 , n31796 , n31797 , n31798 , n31799 , n209561 , n31801 , n31802 , n31803 , n31804 , 
     n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , 
     n31815 , n31816 , n31817 , n209579 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , 
     n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , 
     n31835 , n209597 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , 
     n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , 
     n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n209624 , n31864 , 
     n209626 , n31866 , n209628 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , 
     n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , 
     n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , 
     n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n209662 , n31902 , n31903 , n31904 , 
     n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n209673 , n31913 , n209675 , 
     n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , 
     n31925 , n31926 , n31927 , n31928 , n209690 , n209691 , n31931 , n31932 , n31933 , n31934 , 
     n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n209703 , n31943 , n209705 , 
     n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , 
     n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n209722 , n31962 , n209724 , n31964 , 
     n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n209733 , n31973 , n209735 , 
     n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n209743 , n31983 , n31984 , 
     n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , 
     n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , 
     n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , 
     n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n209785 , 
     n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , 
     n209796 , n32036 , n209798 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , 
     n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , 
     n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , 
     n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , 
     n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n209844 , n32084 , 
     n209846 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , 
     n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , 
     n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n209873 , n32113 , n209875 , 
     n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n209884 , n32124 , 
     n209886 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n209894 , n32134 , 
     n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , 
     n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , 
     n32155 , n32156 , n32157 , n32158 , n32159 , n209921 , n32161 , n32162 , n32163 , n32164 , 
     n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , 
     n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n209942 , n32182 , n32183 , n32184 , 
     n32185 , n32186 , n32187 , n32188 , n32189 , n209951 , n32191 , n209953 , n32193 , n32194 , 
     n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n209965 , 
     n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , 
     n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , 
     n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , 
     n32235 , n32236 , n32237 , n32238 , n210000 , n32240 , n210002 , n32242 , n32243 , n32244 , 
     n32245 , n32246 , n32247 , n32248 , n32249 , n210011 , n32251 , n32252 , n32253 , n32254 , 
     n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , 
     n32265 , n32266 , n32267 , n210029 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , 
     n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n210044 , n32284 , 
     n210046 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , 
     n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , 
     n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , 
     n210076 , n32316 , n210078 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , 
     n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , 
     n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , 
     n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , 
     n32355 , n32356 , n210118 , n32358 , n210120 , n32360 , n32361 , n32362 , n32363 , n32364 , 
     n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n210135 , 
     n32375 , n210137 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , 
     n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n210154 , n32394 , 
     n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , 
     n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , 
     n32415 , n32416 , n210178 , n32418 , n210180 , n32420 , n32421 , n32422 , n32423 , n32424 , 
     n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , 
     n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , 
     n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n210212 , n32452 , n210214 , n32454 , 
     n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , 
     n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , 
     n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , 
     n210246 , n210247 , n32487 , n210249 , n210250 , n32490 , n210252 , n210253 , n32493 , n32494 , 
     n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n210262 , n32502 , n210264 , n32504 , 
     n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , 
     n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , 
     n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , 
     n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , 
     n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , 
     n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , 
     n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , 
     n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , 
     n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , 
     n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n210364 , n32604 , 
     n210366 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , 
     n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , 
     n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , 
     n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , 
     n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , 
     n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , 
     n32665 , n32666 , n32667 , n210429 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , 
     n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , 
     n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , 
     n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , 
     n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , 
     n32715 , n32716 , n32717 , n32718 , n210480 , n32720 , n32721 , n32722 , n32723 , n32724 , 
     n32725 , n32726 , n32727 , n210489 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , 
     n32735 , n32736 , n210498 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , 
     n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , 
     n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , 
     n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n210533 , n32773 , n32774 , 
     n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , 
     n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n210555 , 
     n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n210564 , n32804 , 
     n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , 
     n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , 
     n32825 , n210587 , n32827 , n210589 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , 
     n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , 
     n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , 
     n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , 
     n32865 , n32866 , n210628 , n210629 , n32869 , n210631 , n210632 , n32872 , n32873 , n32874 , 
     n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , 
     n32885 , n32886 , n32887 , n210649 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , 
     n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , 
     n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , 
     n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , 
     n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , 
     n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , 
     n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , 
     n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , 
     n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , 
     n32975 , n210737 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , 
     n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , 
     n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , 
     n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , 
     n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , 
     n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , 
     n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , 
     n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , 
     n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , 
     n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , 
     n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , 
     n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , 
     n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , 
     n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , 
     n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , 
     n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , 
     n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , 
     n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , 
     n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , 
     n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , 
     n33175 , n33176 , n33177 , n33178 , n210940 , n210941 , n33181 , n33182 , n33183 , n33184 , 
     n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n210953 , n33193 , n33194 , 
     n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , 
     n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , 
     n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , 
     n33225 , n33226 , n210988 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , 
     n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , 
     n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , 
     n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , 
     n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , 
     n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , 
     n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , 
     n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , 
     n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , 
     n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , 
     n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , 
     n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , 
     n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , 
     n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , 
     n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , 
     n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n211144 , n33384 , 
     n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , 
     n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , 
     n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , 
     n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , 
     n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , 
     n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , 
     n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , 
     n33455 , n33456 , n33457 , n211219 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , 
     n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , 
     n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , 
     n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , 
     n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , 
     n33505 , n33506 , n33507 , n33508 , n211270 , n211271 , n33511 , n33512 , n33513 , n33514 , 
     n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , 
     n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , 
     n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n211302 , n33542 , n33543 , n33544 , 
     n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , 
     n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , 
     n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , 
     n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , 
     n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , 
     n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , 
     n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , 
     n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , 
     n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , 
     n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , 
     n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , 
     n33655 , n33656 , n33657 , n211419 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , 
     n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , 
     n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , 
     n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , 
     n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , 
     n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , 
     n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , 
     n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , 
     n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , 
     n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , 
     n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , 
     n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , 
     n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n211543 , n211544 , n33784 , 
     n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , 
     n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , 
     n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , 
     n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , 
     n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , 
     n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , 
     n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , 
     n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , 
     n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , 
     n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , 
     n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , 
     n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , 
     n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , 
     n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , 
     n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , 
     n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , 
     n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , 
     n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , 
     n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , 
     n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , 
     n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , 
     n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , 
     n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , 
     n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , 
     n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , 
     n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , 
     n211806 , n211807 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , 
     n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , 
     n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , 
     n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , 
     n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , 
     n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , 
     n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , 
     n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , 
     n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , 
     n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , 
     n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , 
     n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , 
     n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , 
     n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , 
     n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , 
     n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , 
     n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , 
     n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , 
     n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , 
     n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , 
     n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , 
     n212016 , n212017 , n34257 , n212019 , n212020 , n34260 , n34261 , n34262 , n34263 , n34264 , 
     n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , 
     n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , 
     n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , 
     n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , 
     n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , 
     n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , 
     n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , 
     n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , 
     n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , 
     n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , 
     n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , 
     n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , 
     n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , 
     n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , 
     n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , 
     n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , 
     n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , 
     n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , 
     n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , 
     n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , 
     n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , 
     n34475 , n34476 , n34477 , n34478 , n212240 , n212241 , n34481 , n34482 , n34483 , n34484 , 
     n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , 
     n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , 
     n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , 
     n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , 
     n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , 
     n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , 
     n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , 
     n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , 
     n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , 
     n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , 
     n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , 
     n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , 
     n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , 
     n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , 
     n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , 
     n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , 
     n34645 , n34646 , n34647 , n212409 , n212410 , n34650 , n34651 , n34652 , n34653 , n34654 , 
     n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , 
     n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , 
     n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , 
     n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , 
     n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , 
     n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , 
     n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , 
     n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , 
     n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , 
     n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , 
     n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , 
     n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , 
     n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , 
     n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , 
     n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , 
     n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , 
     n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , 
     n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , 
     n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n212602 , n212603 , n34843 , n34844 , 
     n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , 
     n34855 , n34856 , n34857 , n34858 , n34859 , n212621 , n212622 , n212623 , n212624 , n34864 , 
     n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , 
     n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , 
     n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , 
     n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , 
     n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , 
     n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , 
     n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , 
     n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , 
     n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , 
     n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , 
     n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , 
     n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , 
     n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , 
     n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , 
     n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , 
     n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , 
     n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , 
     n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , 
     n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , 
     n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , 
     n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n212834 , n212835 , 
     n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , 
     n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , 
     n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , 
     n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , 
     n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , 
     n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , 
     n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , 
     n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , 
     n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , 
     n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , 
     n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , 
     n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , 
     n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , 
     n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , 
     n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , 
     n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , 
     n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , 
     n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , 
     n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , 
     n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , 
     n35275 , n35276 , n213038 , n213039 , n35279 , n213041 , n213042 , n35282 , n35283 , n35284 , 
     n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , 
     n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , 
     n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , 
     n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , 
     n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , 
     n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , 
     n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , 
     n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , 
     n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , 
     n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , 
     n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , 
     n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , 
     n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , 
     n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , 
     n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , 
     n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , 
     n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , 
     n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n213223 , n213224 , n35464 , 
     n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , 
     n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , 
     n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , 
     n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , 
     n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , 
     n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , 
     n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , 
     n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , 
     n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , 
     n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , 
     n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , 
     n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , 
     n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , 
     n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n213362 , n213363 , n35603 , n35604 , 
     n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , 
     n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , 
     n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , 
     n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n213405 , 
     n213406 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , 
     n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , 
     n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , 
     n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , 
     n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , 
     n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , 
     n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , 
     n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , 
     n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , 
     n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , 
     n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , 
     n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , 
     n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , 
     n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , 
     n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , 
     n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , 
     n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , 
     n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , 
     n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , 
     n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , 
     n35845 , n213607 , n213608 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , 
     n35855 , n35856 , n35857 , n35858 , n213620 , n213621 , n35861 , n35862 , n35863 , n35864 , 
     n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , 
     n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , 
     n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , 
     n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , 
     n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , 
     n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , 
     n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , 
     n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , 
     n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , 
     n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , 
     n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , 
     n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , 
     n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , 
     n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , 
     n36005 , n36006 , n213768 , n213769 , n36009 , n36010 , n36011 , n213773 , n213774 , n36014 , 
     n213776 , n213777 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , 
     n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , 
     n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , 
     n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , 
     n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , 
     n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , 
     n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , 
     n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , 
     n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , 
     n36105 , n213867 , n213868 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , 
     n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , 
     n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , 
     n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , 
     n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , 
     n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n213924 , n213925 , 
     n36165 , n213927 , n213928 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n213935 , 
     n213936 , n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , 
     n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , 
     n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , 
     n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , 
     n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , 
     n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , 
     n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , 
     n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , 
     n36255 , n214017 , n214018 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , 
     n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , 
     n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , 
     n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , 
     n36295 , n36296 , n214058 , n214059 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , 
     n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , 
     n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , 
     n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , 
     n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , 
     n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , 
     n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , 
     n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , 
     n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , 
     n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , 
     n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , 
     n214166 , n214167 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , 
     n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , 
     n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , 
     n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , 
     n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , 
     n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , 
     n36465 , n36466 , n36467 , n214229 , n214230 , n36470 , n214232 , n214233 , n36473 , n214235 , 
     n214236 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , 
     n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , 
     n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , 
     n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , 
     n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , 
     n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , 
     n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , 
     n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , 
     n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , 
     n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , 
     n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , 
     n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , 
     n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , 
     n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , 
     n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , 
     n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , 
     n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , 
     n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , 
     n36655 , n36656 , n36657 , n214419 , n214420 , n36660 , n214422 , n36662 , n36663 , n36664 , 
     n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , 
     n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , 
     n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , 
     n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , 
     n36705 , n214467 , n214468 , n36708 , n36709 , n36710 , n214472 , n214473 , n36713 , n36714 , 
     n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , 
     n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , 
     n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , 
     n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , 
     n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , 
     n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , 
     n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , 
     n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , 
     n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , 
     n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , 
     n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , 
     n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , 
     n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , 
     n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , 
     n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , 
     n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , 
     n36875 , n36876 , n36877 , n214639 , n214640 , n36880 , n36881 , n36882 , n36883 , n36884 , 
     n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , 
     n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , 
     n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , 
     n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , 
     n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , 
     n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , 
     n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n214712 , n214713 , n36953 , n214715 , 
     n214716 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , 
     n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , 
     n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , 
     n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , 
     n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , 
     n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , 
     n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , 
     n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , 
     n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , 
     n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , 
     n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , 
     n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , 
     n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , 
     n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , 
     n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , 
     n37105 , n37106 , n37107 , n214869 , n214870 , n37110 , n37111 , n37112 , n37113 , n37114 , 
     n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , 
     n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , 
     n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , 
     n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , 
     n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , 
     n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , 
     n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , 
     n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , 
     n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , 
     n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n214974 , n214975 , 
     n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , 
     n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , 
     n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , 
     n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , 
     n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , 
     n37265 , n37266 , n37267 , n37268 , n37269 , n215031 , n215032 , n37272 , n37273 , n37274 , 
     n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , 
     n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , 
     n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , 
     n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , 
     n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , 
     n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , 
     n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , n215105 , 
     n215106 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , 
     n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , 
     n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , 
     n37375 , n37376 , n37377 , n215139 , n215140 , n37380 , n215142 , n215143 , n37383 , n37384 , 
     n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , 
     n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , 
     n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , 
     n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , 
     n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , 
     n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , 
     n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , 
     n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , 
     n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , 
     n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , 
     n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , n215255 , 
     n215256 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , 
     n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , 
     n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , 
     n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , 
     n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , 
     n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , 
     n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , 
     n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , 
     n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , 
     n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , 
     n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , 
     n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , 
     n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , 
     n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , 
     n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , 
     n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , 
     n215416 , n215417 , n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , 
     n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , 
     n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , 
     n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , 
     n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , 
     n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , 
     n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , 
     n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , 
     n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , 
     n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , 
     n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , 
     n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , 
     n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , 
     n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , 
     n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , 
     n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , 
     n37815 , n37816 , n37817 , n215579 , n215580 , n37820 , n37821 , n37822 , n37823 , n37824 , 
     n37825 , n215587 , n215588 , n215589 , n215590 , n37830 , n37831 , n37832 , n37833 , n37834 , 
     n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , 
     n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , 
     n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , 
     n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , 
     n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , 
     n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , n37893 , n37894 , 
     n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , 
     n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , 
     n37915 , n37916 , n37917 , n37918 , n215680 , n215681 , n37921 , n37922 , n37923 , n37924 , 
     n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , 
     n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , 
     n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , 
     n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , 
     n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , 
     n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , 
     n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , 
     n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , 
     n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , 
     n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , 
     n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , 
     n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , n215802 , n215803 , n38043 , n38044 , 
     n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , 
     n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , 
     n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , 
     n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , 
     n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , 
     n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , 
     n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , 
     n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , 
     n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , 
     n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , 
     n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , 
     n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , 
     n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , 
     n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , 
     n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , n215954 , n215955 , 
     n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , 
     n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , 
     n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , 
     n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , 
     n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , 
     n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , 
     n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , 
     n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , 
     n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , 
     n38285 , n38286 , n38287 , n216049 , n216050 , n38290 , n216052 , n216053 , n38293 , n38294 , 
     n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , 
     n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , 
     n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , 
     n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , 
     n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , 
     n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , 
     n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , 
     n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , n38371 , n38372 , n38373 , n38374 , 
     n38375 , n216137 , n216138 , n38378 , n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , 
     n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , 
     n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , 
     n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , 
     n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , 
     n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , 
     n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , 
     n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , n38451 , n216213 , n216214 , n38454 , 
     n216216 , n216217 , n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , n216224 , n216225 , 
     n216226 , n216227 , n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , 
     n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , 
     n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , 
     n38495 , n38496 , n38497 , n38498 , n38499 , n216261 , n216262 , n38502 , n38503 , n38504 , 
     n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , 
     n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , 
     n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , 
     n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , 
     n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , 
     n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , 
     n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , 
     n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , 
     n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , n38591 , n38592 , n38593 , n38594 , 
     n38595 , n38596 , n38597 , n216359 , n216360 , n38600 , n38601 , n38602 , n38603 , n38604 , 
     n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , n38611 , n38612 , n38613 , n38614 , 
     n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , n38621 , n38622 , n38623 , n38624 , 
     n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , n38631 , n38632 , n38633 , n38634 , 
     n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , n38641 , n38642 , n38643 , n38644 , 
     n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , n38651 , n216413 , n216414 , n38654 , 
     n216416 , n216417 , n38657 , n38658 , n38659 , n38660 , n38661 , n38662 , n38663 , n38664 , 
     n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , n38671 , n38672 , n38673 , n38674 , 
     n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , n38681 , n38682 , n38683 , n38684 , 
     n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , n38691 , n38692 , n38693 , n38694 , 
     n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , n38701 , n38702 , n38703 , n38704 , 
     n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , n38711 , n38712 , n38713 , n38714 , 
     n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , n38721 , n38722 , n38723 , n38724 , 
     n38725 , n38726 , n38727 , n38728 , n216490 , n216491 , n38731 , n216493 , n216494 , n38734 , 
     n216496 , n216497 , n38737 , n38738 , n38739 , n38740 , n38741 , n38742 , n38743 , n38744 , 
     n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , n38751 , n38752 , n38753 , n38754 , 
     n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , n38761 , n38762 , n38763 , n38764 , 
     n38765 , n38766 , n38767 , n38768 , n38769 , n38770 , n38771 , n38772 , n38773 , n38774 , 
     n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , n38781 , n38782 , n38783 , n38784 , 
     n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , n38791 , n38792 , n38793 , n38794 , 
     n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , n38801 , n38802 , n38803 , n38804 , 
     n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , n38811 , n38812 , n38813 , n38814 , 
     n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , n38821 , n38822 , n38823 , n216585 , 
     n216586 , n38826 , n38827 , n38828 , n38829 , n38830 , n38831 , n38832 , n38833 , n38834 , 
     n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , n216602 , n216603 , n38843 , n38844 , 
     n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , n38851 , n38852 , n38853 , n38854 , 
     n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , n38861 , n38862 , n38863 , n38864 , 
     n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , n38871 , n38872 , n38873 , n38874 , 
     n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , n38881 , n38882 , n38883 , n38884 , 
     n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , n38891 , n38892 , n216654 , n216655 , 
     n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , n38903 , n38904 , 
     n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , n38911 , n38912 , n38913 , n38914 , 
     n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , n38921 , n38922 , n38923 , n38924 , 
     n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , n38931 , n38932 , n38933 , n38934 , 
     n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , n38941 , n38942 , n38943 , n38944 , 
     n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , n38951 , n38952 , n38953 , n38954 , 
     n216716 , n216717 , n38957 , n38958 , n38959 , n38960 , n38961 , n38962 , n38963 , n38964 , 
     n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , n38971 , n38972 , n38973 , n38974 , 
     n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , n38981 , n38982 , n38983 , n38984 , 
     n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , n38991 , n38992 , n38993 , n38994 , 
     n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , n39001 , n39002 , n39003 , n39004 , 
     n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , n39011 , n39012 , n39013 , n39014 , 
     n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , n39021 , n39022 , n39023 , n39024 , 
     n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , n39031 , n39032 , n39033 , n39034 , 
     n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , n39041 , n39042 , n39043 , n39044 , 
     n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , n39051 , n39052 , n39053 , n39054 , 
     n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , n39061 , n39062 , n39063 , n39064 , 
     n39065 , n39066 , n39067 , n39068 , n216830 , n216831 , n39071 , n39072 , n39073 , n39074 , 
     n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , n39081 , n39082 , n39083 , n39084 , 
     n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , n39091 , n39092 , n39093 , n39094 , 
     n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , n39101 , n39102 , n39103 , n39104 , 
     n39105 , n216867 , n216868 , n39108 , n39109 , n39110 , n39111 , n39112 , n39113 , n39114 , 
     n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , n39121 , n39122 , n39123 , n39124 , 
     n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , n39131 , n39132 , n39133 , n39134 , 
     n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , n39141 , n39142 , n39143 , n39144 , 
     n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , n39153 , n39154 , 
     n39155 , n39156 , n39157 , n216919 , n216920 , n39160 , n39161 , n39162 , n39163 , n39164 , 
     n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , n39171 , n39172 , n39173 , n39174 , 
     n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , n39181 , n39182 , n39183 , n39184 , 
     n39185 , n39186 , n216948 , n216949 , n39189 , n216951 , n216952 , n39192 , n39193 , n39194 , 
     n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , n39201 , n39202 , n39203 , n39204 , 
     n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , n39211 , n39212 , n39213 , n39214 , 
     n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , n39221 , n39222 , n39223 , n216985 , 
     n216986 , n39226 , n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , n39233 , n39234 , 
     n39235 , n216997 , n216998 , n216999 , n217000 , n39240 , n217002 , n217003 , n39243 , n39244 , 
     n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , n39251 , n39252 , n39253 , n39254 , 
     n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , n39261 , n39262 , n39263 , n39264 , 
     n39265 , n39266 , n39267 , n39268 , n39269 , n39270 , n39271 , n39272 , n39273 , n39274 , 
     n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , n39281 , n39282 , n39283 , n39284 , 
     n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , n39291 , n39292 , n39293 , n217055 , 
     n217056 , n39296 , n39297 , n39298 , n39299 , n39300 , n39301 , n39302 , n39303 , n39304 , 
     n39305 , n39306 , n39307 , n39308 , n39309 , n217071 , n217072 , n39312 , n39313 , n39314 , 
     n39315 , n39316 , n39317 , n39318 , n39319 , n39320 , n39321 , n39322 , n39323 , n39324 , 
     n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , n39331 , n39332 , n39333 , n39334 , 
     n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , n39341 , n39342 , n39343 , n39344 , 
     n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , n217112 , n217113 , n39353 , n217115 , 
     n39355 , n217117 , n217118 , n39358 , n39359 , n39360 , n39361 , n39362 , n39363 , n39364 , 
     n39365 , n39366 , n39367 , n39368 , n39369 , n39370 , n39371 , n39372 , n39373 , n39374 , 
     n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , n39381 , n39382 , n39383 , n39384 , 
     n39385 , n39386 , n39387 , n39388 , n39389 , n39390 , n39391 , n39392 , n39393 , n39394 , 
     n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , n39401 , n39402 , n39403 , n39404 , 
     n39405 , n39406 , n39407 , n39408 , n39409 , n39410 , n39411 , n39412 , n39413 , n39414 , 
     n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , n39421 , n39422 , n39423 , n39424 , 
     n39425 , n39426 , n39427 , n39428 , n217190 , n217191 , n39431 , n39432 , n39433 , n39434 , 
     n39435 , n39436 , n39437 , n39438 , n39439 , n39440 , n39441 , n39442 , n39443 , n39444 , 
     n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , n39451 , n39452 , n39453 , n39454 , 
     n39455 , n39456 , n39457 , n39458 , n39459 , n39460 , n39461 , n39462 , n39463 , n39464 , 
     n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , n39471 , n39472 , n39473 , n39474 , 
     n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , n39481 , n217243 , n217244 , n39484 , 
     n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , n39491 , n39492 , n39493 , n39494 , 
     n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , n39501 , n39502 , n39503 , n39504 , 
     n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , n39511 , n39512 , n39513 , n39514 , 
     n39515 , n39516 , n39517 , n39518 , n39519 , n39520 , n39521 , n39522 , n39523 , n39524 , 
     n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , n39531 , n39532 , n39533 , n39534 , 
     n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , n39541 , n39542 , n39543 , n39544 , 
     n39545 , n39546 , n39547 , n39548 , n39549 , n39550 , n39551 , n39552 , n39553 , n39554 , 
     n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , n39561 , n39562 , n39563 , n39564 , 
     n39565 , n39566 , n217328 , n217329 , n39569 , n39570 , n39571 , n39572 , n39573 , n39574 , 
     n217336 , n217337 , n217338 , n217339 , n39579 , n39580 , n39581 , n39582 , n39583 , n39584 , 
     n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , n39591 , n39592 , n39593 , n39594 , 
     n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , n39601 , n39602 , n39603 , n39604 , 
     n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , n39611 , n39612 , n39613 , n39614 , 
     n39615 , n39616 , n39617 , n39618 , n39619 , n39620 , n39621 , n39622 , n39623 , n39624 , 
     n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , n39631 , n39632 , n39633 , n39634 , 
     n39635 , n39636 , n39637 , n39638 , n39639 , n39640 , n39641 , n39642 , n39643 , n39644 , 
     n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , n39651 , n39652 , n39653 , n39654 , 
     n39655 , n39656 , n39657 , n39658 , n39659 , n217421 , n217422 , n39662 , n39663 , n39664 , 
     n39665 , n39666 , n39667 , n39668 , n39669 , n39670 , n39671 , n39672 , n39673 , n39674 , 
     n39675 , n39676 , n39677 , n39678 , n39679 , n39680 , n39681 , n39682 , n39683 , n39684 , 
     n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , n39691 , n39692 , n39693 , n39694 , 
     n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , n39701 , n39702 , n39703 , n39704 , 
     n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , n39711 , n39712 , n217474 , n217475 , 
     n39715 , n217477 , n217478 , n39718 , n39719 , n39720 , n39721 , n39722 , n39723 , n39724 , 
     n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , n39731 , n39732 , n39733 , n39734 , 
     n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , n39741 , n39742 , n39743 , n39744 , 
     n39745 , n39746 , n39747 , n39748 , n39749 , n217511 , n217512 , n39752 , n217514 , n217515 , 
     n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , n39761 , n39762 , n39763 , n39764 , 
     n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , n39771 , n39772 , n39773 , n39774 , 
     n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , n39781 , n39782 , n39783 , n39784 , 
     n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , n39791 , n39792 , n39793 , n39794 , 
     n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , n39801 , n39802 , n39803 , n39804 , 
     n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , n39811 , n39812 , n39813 , n39814 , 
     n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , n39821 , n39822 , n39823 , n217585 , 
     n217586 , n39826 , n217588 , n217589 , n39829 , n39830 , n39831 , n39832 , n39833 , n39834 , 
     n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , n39841 , n39842 , n39843 , n39844 , 
     n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , n39851 , n39852 , n39853 , n39854 , 
     n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , n39861 , n39862 , n39863 , n39864 , 
     n39865 , n39866 , n39867 , n39868 , n39869 , n39870 , n39871 , n39872 , n39873 , n39874 , 
     n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , n39881 , n39882 , n39883 , n39884 , 
     n39885 , n39886 , n39887 , n39888 , n39889 , n217651 , n217652 , n39892 , n39893 , n39894 , 
     n39895 , n39896 , n39897 , n39898 , n39899 , n39900 , n39901 , n39902 , n39903 , n39904 , 
     n39905 , n39906 , n39907 , n39908 , n39909 , n39910 , n39911 , n39912 , n39913 , n39914 , 
     n39915 , n39916 , n39917 , n39918 , n39919 , n39920 , n39921 , n39922 , n39923 , n39924 , 
     n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , n39931 , n39932 , n39933 , n39934 , 
     n39935 , n39936 , n39937 , n39938 , n39939 , n39940 , n39941 , n39942 , n39943 , n39944 , 
     n39945 , n39946 , n39947 , n39948 , n39949 , n39950 , n39951 , n39952 , n39953 , n39954 , 
     n39955 , n217717 , n217718 , n39958 , n39959 , n39960 , n39961 , n39962 , n39963 , n39964 , 
     n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , n39971 , n39972 , n39973 , n39974 , 
     n39975 , n39976 , n39977 , n39978 , n39979 , n39980 , n39981 , n39982 , n39983 , n39984 , 
     n39985 , n39986 , n39987 , n39988 , n39989 , n39990 , n39991 , n39992 , n39993 , n39994 , 
     n39995 , n39996 , n39997 , n39998 , n39999 , n40000 , n40001 , n40002 , n40003 , n40004 , 
     n40005 , n40006 , n40007 , n40008 , n40009 , n40010 , n40011 , n40012 , n40013 , n40014 , 
     n40015 , n40016 , n40017 , n40018 , n40019 , n40020 , n40021 , n40022 , n40023 , n40024 , 
     n40025 , n40026 , n40027 , n40028 , n40029 , n40030 , n40031 , n40032 , n40033 , n40034 , 
     n40035 , n40036 , n40037 , n40038 , n40039 , n40040 , n40041 , n40042 , n40043 , n40044 , 
     n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , n40051 , n40052 , n40053 , n40054 , 
     n217816 , n217817 , n40057 , n217819 , n217820 , n40060 , n40061 , n40062 , n40063 , n40064 , 
     n40065 , n40066 , n40067 , n40068 , n40069 , n40070 , n40071 , n40072 , n217834 , n217835 , 
     n40075 , n40076 , n40077 , n40078 , n40079 , n40080 , n40081 , n40082 , n40083 , n40084 , 
     n40085 , n40086 , n40087 , n40088 , n40089 , n40090 , n40091 , n40092 , n40093 , n40094 , 
     n40095 , n40096 , n40097 , n40098 , n40099 , n40100 , n40101 , n40102 , n40103 , n40104 , 
     n40105 , n40106 , n40107 , n40108 , n40109 , n40110 , n40111 , n40112 , n40113 , n40114 , 
     n40115 , n40116 , n40117 , n40118 , n40119 , n40120 , n40121 , n40122 , n217884 , n217885 , 
     n40125 , n40126 , n40127 , n40128 , n40129 , n40130 , n40131 , n40132 , n40133 , n40134 , 
     n40135 , n40136 , n40137 , n40138 , n40139 , n40140 , n40141 , n40142 , n40143 , n40144 , 
     n40145 , n40146 , n40147 , n40148 , n40149 , n40150 , n40151 , n40152 , n40153 , n40154 , 
     n40155 , n40156 , n40157 , n40158 , n40159 , n40160 , n40161 , n40162 , n40163 , n40164 , 
     n40165 , n40166 , n40167 , n40168 , n40169 , n40170 , n40171 , n40172 , n217934 , n217935 , 
     n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , n40181 , n40182 , n40183 , n40184 , 
     n40185 , n40186 , n40187 , n40188 , n40189 , n40190 , n40191 , n40192 , n40193 , n40194 , 
     n40195 , n40196 , n40197 , n40198 , n40199 , n40200 , n40201 , n40202 , n40203 , n40204 , 
     n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , n40211 , n40212 , n40213 , n40214 , 
     n40215 , n40216 , n40217 , n40218 , n40219 , n217981 , n217982 , n40222 , n40223 , n40224 , 
     n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , n40231 , n40232 , n40233 , n40234 , 
     n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , n40241 , n40242 , n40243 , n40244 , 
     n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , n40251 , n40252 , n40253 , n40254 , 
     n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , n40261 , n40262 , n218024 , n218025 , 
     n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , n40271 , n40272 , n40273 , n40274 , 
     n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , n40281 , n40282 , n40283 , n40284 , 
     n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , n40291 , n40292 , n40293 , n40294 , 
     n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , n40301 , n40302 , n40303 , n40304 , 
     n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , n40311 , n40312 , n40313 , n40314 , 
     n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , n40321 , n40322 , n218084 , n218085 , 
     n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , n40331 , n40332 , n40333 , n40334 , 
     n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , n40341 , n40342 , n40343 , n40344 , 
     n40345 , n40346 , n40347 , n40348 , n40349 , n40350 , n40351 , n40352 , n40353 , n40354 , 
     n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , n40361 , n40362 , n40363 , n40364 , 
     n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , n40371 , n40372 , n40373 , n40374 , 
     n40375 , n40376 , n40377 , n40378 , n40379 , n40380 , n40381 , n40382 , n40383 , n40384 , 
     n40385 , n218147 , n218148 , n40388 , n40389 , n40390 , n40391 , n40392 , n40393 , n40394 , 
     n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , n40401 , n40402 , n40403 , n40404 , 
     n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , n40411 , n40412 , n40413 , n40414 , 
     n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , n40421 , n40422 , n40423 , n40424 , 
     n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , n40431 , n40432 , n40433 , n40434 , 
     n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , n218202 , n218203 , n40443 , n40444 , 
     n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , n40451 , n40452 , n40453 , n40454 , 
     n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , n40461 , n40462 , n40463 , n40464 , 
     n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , n40471 , n40472 , n40473 , n40474 , 
     n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , n40481 , n40482 , n40483 , n40484 , 
     n40485 , n40486 , n40487 , n40488 , n40489 , n40490 , n40491 , n40492 , n40493 , n40494 , 
     n40495 , n40496 , n40497 , n40498 , n40499 , n40500 , n40501 , n40502 , n40503 , n40504 , 
     n40505 , n40506 , n40507 , n40508 , n40509 , n40510 , n40511 , n40512 , n40513 , n40514 , 
     n40515 , n40516 , n40517 , n40518 , n40519 , n218281 , n218282 , n40522 , n40523 , n40524 , 
     n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , n40531 , n218293 , n218294 , n40534 , 
     n40535 , n218297 , n218298 , n40538 , n218300 , n218301 , n40541 , n40542 , n40543 , n40544 , 
     n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , n40551 , n40552 , n40553 , n40554 , 
     n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , n40561 , n40562 , n40563 , n40564 , 
     n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , n40571 , n40572 , n40573 , n40574 , 
     n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , n40581 , n40582 , n40583 , n40584 , 
     n40585 , n40586 , n40587 , n40588 , n40589 , n218351 , n218352 , n40592 , n40593 , n40594 , 
     n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , n40601 , n40602 , n40603 , n218365 , 
     n218366 , n40606 , n40607 , n40608 , n218370 , n218371 , n40611 , n40612 , n40613 , n40614 , 
     n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , n40621 , n40622 , n40623 , n40624 , 
     n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , n40631 , n40632 , n40633 , n40634 , 
     n218396 , n218397 , n40637 , n40638 , n40639 , n40640 , n40641 , n218403 , n218404 , n218405 , 
     n218406 , n40646 , n40647 , n40648 , n40649 , n40650 , n40651 , n40652 , n40653 , n40654 , 
     n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , n40661 , n40662 , n40663 , n40664 , 
     n40665 , n40666 , n40667 , n40668 , n40669 , n218431 , n218432 , n40672 , n40673 , n40674 , 
     n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , n40681 , n40682 , n40683 , n40684 , 
     n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , n40691 , n40692 , n40693 , n40694 , 
     n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , n40701 , n40702 , n40703 , n40704 , 
     n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , n40711 , n40712 , n40713 , n40714 , 
     n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , n40721 , n218483 , n218484 , n40724 , 
     n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , n40731 , n40732 , n40733 , n40734 , 
     n40735 , n40736 , n40737 , n40738 , n40739 , n40740 , n40741 , n40742 , n40743 , n40744 , 
     n40745 , n40746 , n40747 , n40748 , n40749 , n218511 , n218512 , n40752 , n40753 , n40754 , 
     n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , n40761 , n40762 , n40763 , n40764 , 
     n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , n40771 , n40772 , n40773 , n40774 , 
     n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , n218542 , n218543 , n40783 , n218545 , 
     n218546 , n40786 , n40787 , n40788 , n40789 , n40790 , n40791 , n40792 , n40793 , n40794 , 
     n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , n40801 , n40802 , n40803 , n40804 , 
     n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , n40811 , n40812 , n40813 , n40814 , 
     n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , n40821 , n40822 , n40823 , n40824 , 
     n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , n40831 , n40832 , n40833 , n40834 , 
     n218596 , n218597 , n40837 , n40838 , n40839 , n40840 , n40841 , n40842 , n40843 , n40844 , 
     n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , n40851 , n40852 , n40853 , n40854 , 
     n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , n40861 , n40862 , n218624 , n218625 , 
     n40865 , n40866 , n40867 , n40868 , n40869 , n40870 , n40871 , n40872 , n40873 , n40874 , 
     n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , n40881 , n40882 , n40883 , n40884 , 
     n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , n40891 , n40892 , n40893 , n218655 , 
     n218656 , n40896 , n40897 , n40898 , n40899 , n40900 , n40901 , n40902 , n40903 , n40904 , 
     n40905 , n40906 , n40907 , n40908 , n40909 , n40910 , n40911 , n40912 , n40913 , n40914 , 
     n40915 , n40916 , n40917 , n40918 , n218680 , n218681 , n40921 , n40922 , n40923 , n40924 , 
     n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , n40931 , n40932 , n40933 , n40934 , 
     n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , n40941 , n40942 , n40943 , n40944 , 
     n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , n40951 , n40952 , n40953 , n40954 , 
     n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , n40961 , n40962 , n40963 , n40964 , 
     n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , n218732 , n218733 , n40973 , n40974 , 
     n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , n40981 , n40982 , n40983 , n218745 , 
     n218746 , n40986 , n218748 , n218749 , n40989 , n40990 , n40991 , n40992 , n40993 , n40994 , 
     n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , n41001 , n41002 , n41003 , n41004 , 
     n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , n41011 , n41012 , n218774 , n218775 , 
     n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , n41021 , n41022 , n41023 , n41024 , 
     n218786 , n218787 , n41027 , n41028 , n41029 , n41030 , n41031 , n41032 , n41033 , n41034 , 
     n41035 , n41036 , n41037 , n41038 , n41039 , n41040 , n41041 , n41042 , n41043 , n41044 , 
     n41045 , n41046 , n41047 , n41048 , n41049 , n41050 , n41051 , n41052 , n41053 , n41054 , 
     n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , n41061 , n41062 , n41063 , n41064 , 
     n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , n41071 , n218833 , n218834 , n41074 , 
     n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , n41081 , n41082 , n41083 , n41084 , 
     n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , n41091 , n41092 , n41093 , n41094 , 
     n41095 , n41096 , n41097 , n41098 , n41099 , n41100 , n41101 , n41102 , n218864 , n218865 , 
     n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , n41111 , n41112 , n41113 , n41114 , 
     n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , n41121 , n41122 , n41123 , n41124 , 
     n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , n41131 , n41132 , n41133 , n218895 , 
     n218896 , n41136 , n41137 , n41138 , n41139 , n41140 , n41141 , n41142 , n41143 , n41144 , 
     n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , n41151 , n41152 , n41153 , n41154 , 
     n41155 , n218917 , n218918 , n41158 , n41159 , n41160 , n41161 , n41162 , n41163 , n41164 , 
     n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , n41171 , n41172 , n41173 , n218935 , 
     n218936 , n41176 , n218938 , n218939 , n41179 , n41180 , n41181 , n41182 , n41183 , n41184 , 
     n41185 , n41186 , n41187 , n41188 , n41189 , n41190 , n41191 , n41192 , n41193 , n41194 , 
     n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , n41201 , n41202 , n41203 , n41204 , 
     n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , n41211 , n41212 , n41213 , n41214 , 
     n41215 , n41216 , n41217 , n41218 , n41219 , n218981 , n218982 , n41222 , n218984 , n218985 , 
     n41225 , n41226 , n41227 , n41228 , n41229 , n41230 , n41231 , n41232 , n41233 , n41234 , 
     n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , n41241 , n41242 , n41243 , n41244 , 
     n41245 , n41246 , n41247 , n219009 , n219010 , n41250 , n41251 , n41252 , n41253 , n41254 , 
     n41255 , n41256 , n41257 , n41258 , n41259 , n219021 , n219022 , n41262 , n41263 , n41264 , 
     n41265 , n41266 , n41267 , n41268 , n41269 , n41270 , n41271 , n41272 , n41273 , n41274 , 
     n41275 , n41276 , n41277 , n41278 , n41279 , n41280 , n41281 , n41282 , n41283 , n41284 , 
     n41285 , n41286 , n41287 , n41288 , n41289 , n41290 , n219052 , n219053 , n41293 , n41294 , 
     n41295 , n41296 , n41297 , n41298 , n41299 , n41300 , n41301 , n41302 , n41303 , n41304 , 
     n41305 , n41306 , n41307 , n41308 , n41309 , n41310 , n41311 , n41312 , n41313 , n41314 , 
     n41315 , n41316 , n41317 , n41318 , n41319 , n41320 , n41321 , n41322 , n219084 , n219085 , 
     n41325 , n41326 , n41327 , n41328 , n41329 , n41330 , n41331 , n41332 , n219094 , n219095 , 
     n41335 , n41336 , n41337 , n41338 , n41339 , n41340 , n41341 , n41342 , n41343 , n41344 , 
     n41345 , n41346 , n41347 , n219109 , n219110 , n41350 , n41351 , n219113 , n41353 , n219115 , 
     n219116 , n41356 , n41357 , n41358 , n41359 , n41360 , n41361 , n41362 , n41363 , n41364 , 
     n41365 , n41366 , n41367 , n41368 , n41369 , n41370 , n41371 , n41372 , n41373 , n41374 , 
     n41375 , n41376 , n41377 , n41378 , n41379 , n41380 , n41381 , n41382 , n41383 , n41384 , 
     n41385 , n41386 , n41387 , n41388 , n41389 , n41390 , n41391 , n41392 , n41393 , n41394 , 
     n41395 , n219157 , n219158 , n41398 , n41399 , n41400 , n41401 , n41402 , n41403 , n41404 , 
     n41405 , n41406 , n41407 , n219169 , n219170 , n41410 , n41411 , n41412 , n41413 , n41414 , 
     n41415 , n41416 , n41417 , n41418 , n41419 , n41420 , n41421 , n41422 , n41423 , n41424 , 
     n41425 , n41426 , n41427 , n41428 , n41429 , n41430 , n41431 , n41432 , n41433 , n41434 , 
     n41435 , n41436 , n41437 , n41438 , n219200 , n219201 , n41441 , n41442 , n41443 , n41444 , 
     n41445 , n41446 , n41447 , n41448 , n41449 , n41450 , n41451 , n41452 , n41453 , n219215 , 
     n219216 , n41456 , n41457 , n219219 , n219220 , n41460 , n41461 , n41462 , n41463 , n41464 , 
     n41465 , n41466 , n41467 , n41468 , n41469 , n41470 , n41471 , n41472 , n41473 , n41474 , 
     n41475 , n41476 , n41477 , n41478 , n41479 , n41480 , n41481 , n41482 , n41483 , n41484 , 
     n41485 , n41486 , n41487 , n41488 , n41489 , n41490 , n41491 , n41492 , n41493 , n41494 , 
     n41495 , n41496 , n41497 , n41498 , n41499 , n41500 , n41501 , n41502 , n41503 , n41504 , 
     n41505 , n41506 , n41507 , n219269 , n219270 , n41510 , n41511 , n41512 , n41513 , n41514 , 
     n41515 , n41516 , n41517 , n41518 , n41519 , n41520 , n41521 , n41522 , n41523 , n41524 , 
     n41525 , n41526 , n41527 , n41528 , n41529 , n41530 , n41531 , n41532 , n41533 , n41534 , 
     n41535 , n41536 , n41537 , n41538 , n41539 , n41540 , n41541 , n41542 , n41543 , n41544 , 
     n41545 , n41546 , n41547 , n41548 , n41549 , n219311 , n219312 , n41552 , n219314 , n219315 , 
     n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , n41561 , n41562 , n41563 , n41564 , 
     n41565 , n41566 , n219328 , n219329 , n41569 , n41570 , n41571 , n41572 , n41573 , n41574 , 
     n41575 , n41576 , n41577 , n41578 , n41579 , n41580 , n41581 , n41582 , n41583 , n41584 , 
     n41585 , n41586 , n41587 , n41588 , n41589 , n41590 , n41591 , n41592 , n41593 , n41594 , 
     n219356 , n219357 , n41597 , n219359 , n219360 , n41600 , n41601 , n41602 , n41603 , n41604 , 
     n41605 , n41606 , n41607 , n41608 , n41609 , n41610 , n41611 , n41612 , n41613 , n41614 , 
     n41615 , n41616 , n41617 , n41618 , n41619 , n41620 , n41621 , n41622 , n41623 , n41624 , 
     n41625 , n41626 , n41627 , n41628 , n41629 , n41630 , n41631 , n41632 , n41633 , n41634 , 
     n219396 , n219397 , n41637 , n41638 , n41639 , n41640 , n41641 , n41642 , n41643 , n41644 , 
     n41645 , n41646 , n41647 , n41648 , n41649 , n41650 , n41651 , n41652 , n41653 , n41654 , 
     n41655 , n41656 , n41657 , n41658 , n41659 , n41660 , n41661 , n41662 , n41663 , n41664 , 
     n41665 , n41666 , n41667 , n41668 , n219430 , n219431 , n41671 , n41672 , n41673 , n41674 , 
     n41675 , n41676 , n41677 , n41678 , n41679 , n41680 , n41681 , n41682 , n41683 , n41684 , 
     n41685 , n41686 , n41687 , n41688 , n41689 , n41690 , n41691 , n41692 , n41693 , n41694 , 
     n41695 , n219457 , n219458 , n41698 , n41699 , n41700 , n41701 , n41702 , n41703 , n41704 , 
     n41705 , n41706 , n41707 , n219469 , n219470 , n41710 , n41711 , n41712 , n41713 , n41714 , 
     n41715 , n41716 , n41717 , n41718 , n41719 , n219481 , n219482 , n41722 , n41723 , n41724 , 
     n41725 , n41726 , n41727 , n41728 , n41729 , n41730 , n41731 , n41732 , n41733 , n41734 , 
     n41735 , n41736 , n41737 , n41738 , n41739 , n41740 , n41741 , n41742 , n41743 , n41744 , 
     n41745 , n41746 , n41747 , n219509 , n219510 , n41750 , n41751 , n41752 , n41753 , n41754 , 
     n41755 , n41756 , n41757 , n41758 , n41759 , n41760 , n41761 , n41762 , n41763 , n41764 , 
     n41765 , n41766 , n41767 , n41768 , n41769 , n41770 , n41771 , n41772 , n41773 , n41774 , 
     n41775 , n219537 , n219538 , n41778 , n41779 , n41780 , n41781 , n41782 , n41783 , n41784 , 
     n41785 , n41786 , n41787 , n41788 , n41789 , n41790 , n41791 , n41792 , n41793 , n41794 , 
     n41795 , n41796 , n41797 , n41798 , n41799 , n41800 , n41801 , n41802 , n41803 , n41804 , 
     n41805 , n41806 , n41807 , n41808 , n41809 , n41810 , n41811 , n41812 , n41813 , n41814 , 
     n41815 , n41816 , n41817 , n41818 , n41819 , n41820 , n41821 , n41822 , n219584 , n219585 , 
     n41825 , n41826 , n41827 , n41828 , n41829 , n41830 , n41831 , n41832 , n219594 , n219595 , 
     n41835 , n41836 , n41837 , n41838 , n41839 , n41840 , n41841 , n41842 , n41843 , n41844 , 
     n41845 , n41846 , n41847 , n41848 , n41849 , n41850 , n41851 , n41852 , n41853 , n41854 , 
     n41855 , n41856 , n41857 , n41858 , n41859 , n41860 , n219622 , n219623 , n41863 , n219625 , 
     n219626 , n41866 , n41867 , n41868 , n41869 , n41870 , n41871 , n41872 , n41873 , n41874 , 
     n41875 , n41876 , n41877 , n41878 , n41879 , n41880 , n41881 , n41882 , n41883 , n41884 , 
     n41885 , n41886 , n41887 , n41888 , n219650 , n219651 , n41891 , n41892 , n41893 , n41894 , 
     n41895 , n41896 , n41897 , n41898 , n41899 , n41900 , n219662 , n219663 , n41903 , n41904 , 
     n41905 , n41906 , n41907 , n41908 , n41909 , n41910 , n41911 , n41912 , n219674 , n219675 , 
     n41915 , n41916 , n41917 , n41918 , n41919 , n41920 , n41921 , n41922 , n41923 , n41924 , 
     n41925 , n41926 , n41927 , n41928 , n41929 , n41930 , n41931 , n41932 , n41933 , n41934 , 
     n41935 , n41936 , n41937 , n41938 , n41939 , n219701 , n219702 , n41942 , n41943 , n41944 , 
     n41945 , n41946 , n41947 , n41948 , n41949 , n41950 , n41951 , n41952 , n41953 , n41954 , 
     n219716 , n219717 , n41957 , n41958 , n41959 , n41960 , n41961 , n41962 , n41963 , n41964 , 
     n41965 , n41966 , n219728 , n219729 , n41969 , n41970 , n41971 , n41972 , n41973 , n41974 , 
     n41975 , n41976 , n41977 , n41978 , n41979 , n41980 , n41981 , n41982 , n41983 , n41984 , 
     n41985 , n41986 , n41987 , n41988 , n41989 , n41990 , n41991 , n41992 , n41993 , n41994 , 
     n41995 , n41996 , n41997 , n219759 , n219760 , n42000 , n42001 , n42002 , n42003 , n42004 , 
     n42005 , n42006 , n42007 , n42008 , n42009 , n42010 , n42011 , n42012 , n219774 , n219775 , 
     n42015 , n42016 , n42017 , n42018 , n42019 , n42020 , n42021 , n42022 , n42023 , n42024 , 
     n42025 , n42026 , n42027 , n42028 , n42029 , n42030 , n42031 , n42032 , n42033 , n42034 , 
     n42035 , n42036 , n42037 , n42038 , n42039 , n42040 , n42041 , n42042 , n42043 , n42044 , 
     n42045 , n42046 , n42047 , n42048 , n42049 , n42050 , n42051 , n42052 , n42053 , n219815 , 
     n219816 , n42056 , n42057 , n42058 , n42059 , n42060 , n42061 , n219823 , n219824 , n42064 , 
     n42065 , n219827 , n219828 , n42068 , n42069 , n42070 , n42071 , n42072 , n42073 , n42074 , 
     n42075 , n42076 , n42077 , n42078 , n219840 , n219841 , n42081 , n42082 , n42083 , n42084 , 
     n42085 , n42086 , n42087 , n42088 , n219850 , n219851 , n42091 , n42092 , n42093 , n42094 , 
     n42095 , n42096 , n42097 , n42098 , n42099 , n42100 , n42101 , n42102 , n219864 , n219865 , 
     n42105 , n219867 , n219868 , n42108 , n42109 , n42110 , n42111 , n42112 , n42113 , n42114 , 
     n42115 , n42116 , n42117 , n42118 , n42119 , n219881 , n219882 , n42122 , n42123 , n42124 , 
     n42125 , n42126 , n42127 , n42128 , n219890 , n219891 , n42131 , n42132 , n42133 , n42134 , 
     n42135 , n42136 , n42137 , n42138 , n42139 , n42140 , n219902 , n219903 , n42143 , n219905 , 
     n219906 , n42146 , n42147 , n42148 , n42149 , n42150 , n42151 , n219913 , n219914 , n42154 , 
     n42155 , n42156 , n42157 , n42158 , n42159 , n42160 , n42161 , n42162 , n42163 , n42164 , 
     n42165 , n219927 , n219928 , n42168 , n42169 , n42170 , n42171 , n42172 , n42173 , n42174 , 
     n42175 , n42176 , n42177 , n42178 , n42179 , n42180 , n42181 , n42182 , n42183 , n42184 , 
     n42185 , n42186 , n42187 , n42188 , n42189 , n42190 , n42191 , n42192 , n42193 , n42194 , 
     n42195 , n42196 , n219958 , n219959 , n42199 , n42200 , n42201 , n42202 , n42203 , n42204 , 
     n42205 , n42206 , n42207 , n42208 , n219970 , n219971 , n42211 , n219973 , n219974 , n42214 , 
     n219976 , n219977 , n42217 , n219979 , n219980 , n42220 , n219982 , n219983 , n42223 , n42224 , 
     n42225 , n42226 , n42227 , n42228 , n42229 , n42230 , n219992 , n219993 , n42233 , n42234 , 
     n42235 , n42236 , n42237 , n42238 , n42239 , n42240 , n42241 , n42242 , n220004 , n220005 , 
     n42245 , n42246 , n42247 , n42248 , n42249 , n42250 , n42251 , n42252 , n42253 , n42254 , 
     n42255 , n42256 , n42257 , n42258 , n42259 , n42260 , n42261 , n42262 , n42263 , n42264 , 
     n42265 , n42266 , n42267 , n42268 , n42269 , n42270 , n42271 , n42272 , n42273 , n220035 , 
     n220036 , n42276 , n42277 , n42278 , n42279 , n42280 , n42281 , n42282 , n42283 , n42284 , 
     n42285 , n220047 , n220048 , n42288 , n42289 , n42290 , n42291 , n42292 , n42293 , n42294 , 
     n42295 , n42296 , n42297 , n42298 , n42299 , n42300 , n42301 , n42302 , n42303 , n42304 , 
     n42305 , n42306 , n42307 , n42308 , n42309 , n42310 , n42311 , n42312 , n220074 , n220075 , 
     n42315 , n42316 , n42317 , n42318 , n42319 , n42320 , n42321 , n42322 , n42323 , n42324 , 
     n42325 , n42326 , n42327 , n220089 , n220090 , n42330 , n42331 , n42332 , n42333 , n42334 , 
     n42335 , n42336 , n42337 , n42338 , n42339 , n42340 , n42341 , n42342 , n42343 , n42344 , 
     n42345 , n42346 , n42347 , n42348 , n42349 , n42350 , n42351 , n42352 , n220114 , n220115 , 
     n42355 , n42356 , n42357 , n42358 , n42359 , n42360 , n42361 , n42362 , n42363 , n42364 , 
     n220126 , n220127 , n42367 , n42368 , n42369 , n42370 , n42371 , n42372 , n42373 , n42374 , 
     n42375 , n42376 , n42377 , n42378 , n42379 , n42380 , n42381 , n42382 , n42383 , n220145 , 
     n220146 , n42386 , n42387 , n42388 , n42389 , n42390 , n42391 , n220153 , n220154 , n42394 , 
     n220156 , n220157 , n42397 , n42398 , n42399 , n42400 , n42401 , n42402 , n42403 , n42404 , 
     n220166 , n220167 , n42407 , n42408 , n42409 , n42410 , n42411 , n42412 , n42413 , n42414 , 
     n42415 , n42416 , n220178 , n220179 , n42419 , n42420 , n42421 , n42422 , n42423 , n42424 , 
     n220186 , n220187 , n42427 , n42428 , n42429 , n42430 , n42431 , n42432 , n42433 , n42434 , 
     n42435 , n42436 , n220198 , n220199 , n42439 , n220201 , n220202 , n42442 , n42443 , n42444 , 
     n42445 , n42446 , n42447 , n42448 , n42449 , n42450 , n42451 , n220213 , n220214 , n42454 , 
     n42455 , n42456 , n42457 , n42458 , n42459 , n42460 , n42461 , n42462 , n42463 , n220225 , 
     n220226 , n42466 , n42467 , n42468 , n42469 , n42470 , n42471 , n42472 , n42473 , n42474 , 
     n42475 , n220237 , n220238 , n42478 , n42479 , n42480 , n42481 , n42482 , n42483 , n42484 , 
     n42485 , n42486 , n42487 , n220249 , n220250 , n42490 , n42491 , n42492 , n42493 , n42494 , 
     n42495 , n42496 , n42497 , n42498 , n42499 , n42500 , n42501 , n42502 , n42503 , n42504 , 
     n42505 , n42506 , n42507 , n42508 , n42509 , n42510 , n42511 , n42512 , n220274 , n220275 , 
     n42515 , n220277 , n220278 , n42518 , n42519 , n42520 , n42521 , n42522 , n42523 , n42524 , 
     n42525 , n42526 , n42527 , n220289 , n220290 , n42530 , n42531 , n42532 , n42533 , n42534 , 
     n42535 , n42536 , n42537 , n42538 , n42539 , n42540 , n42541 , n42542 , n42543 , n42544 , 
     n42545 , n42546 , n42547 , n42548 , n42549 , n42550 , n42551 , n42552 , n42553 , n42554 , 
     n42555 , n42556 , n42557 , n42558 , n220320 , n220321 , n42561 , n42562 , n42563 , n42564 , 
     n42565 , n42566 , n220328 , n220329 , n42569 , n220331 , n220332 , n42572 , n42573 , n42574 , 
     n42575 , n42576 , n42577 , n42578 , n42579 , n42580 , n42581 , n220343 , n220344 , n42584 , 
     n220346 , n220347 , n42587 , n42588 , n42589 , n42590 , n42591 , n42592 , n42593 , n42594 , 
     n42595 , n42596 , n42597 , n42598 , n42599 , n42600 , n42601 , n42602 , n42603 , n42604 , 
     n42605 , n42606 , n42607 , n42608 , n42609 , n42610 , n42611 , n42612 , n42613 , n42614 , 
     n42615 , n42616 , n42617 , n42618 , n42619 , n42620 , n42621 , n42622 , n42623 , n42624 , 
     n42625 , n42626 , n42627 , n42628 , n42629 , n42630 , n42631 , n42632 , n42633 , n42634 , 
     n42635 , n42636 , n42637 , n42638 , n220400 , n220401 , n42641 , n42642 , n42643 , n42644 , 
     n42645 , n42646 , n42647 , n42648 , n42649 , n42650 , n220412 , n220413 , n42653 , n42654 , 
     n42655 , n42656 , n42657 , n42658 , n220420 , n220421 , n42661 , n220423 , n220424 , n42664 , 
     n42665 , n42666 , n42667 , n42668 , n42669 , n42670 , n220432 , n220433 , n220434 , n220435 , 
     n42675 , n42676 , n42677 , n42678 , n42679 , n42680 , n42681 , n42682 , n42683 , n42684 , 
     n42685 , n220447 , n220448 , n42688 , n42689 , n42690 , n42691 , n42692 , n42693 , n42694 , 
     n220456 , n220457 , n42697 , n220459 , n220460 , n42700 , n42701 , n42702 , n42703 , n42704 , 
     n42705 , n220467 , n220468 , n42708 , n42709 , n220471 , n220472 , n42712 , n42713 , n42714 , 
     n42715 , n42716 , n42717 , n42718 , n220480 , n220481 , n42721 , n42722 , n42723 , n42724 , 
     n42725 , n42726 , n42727 , n42728 , n42729 , n42730 , n220492 , n220493 , n42733 , n42734 , 
     n42735 , n42736 , n42737 , n42738 , n42739 , n42740 , n42741 , n42742 , n220504 , n220505 , 
     n42745 , n42746 , n42747 , n42748 , n42749 , n42750 , n42751 , n42752 , n42753 , n42754 , 
     n42755 , n42756 , n220518 , n220519 , n42759 , n42760 , n42761 , n42762 , n42763 , n42764 , 
     n42765 , n42766 , n220528 , n220529 , n42769 , n220531 , n220532 , n42772 , n220534 , n220535 , 
     n42775 , n42776 , n42777 , n42778 , n42779 , n42780 , n220542 , n220543 , n42783 , n220545 , 
     n220546 , n42786 , n42787 , n42788 , n42789 , n42790 , n42791 , n42792 , n42793 , n42794 , 
     n42795 , n220557 , n220558 , n42798 , n220560 , n220561 , n42801 , n42802 , n42803 , n42804 , 
     n42805 , n42806 , n220568 , n220569 , n42809 , n42810 , n42811 , n42812 , n220574 , n220575 , 
     n42815 , n220577 , n220578 , n42818 , n42819 , n42820 , n42821 , n42822 , n42823 , n42824 , 
     n42825 , n42826 , n42827 , n220589 , n220590 , n42830 , n42831 , n42832 , n42833 , n42834 , 
     n42835 , n42836 , n42837 , n42838 , n42839 , n220601 , n220602 , n42842 , n42843 , n42844 , 
     n42845 , n42846 , n42847 , n42848 , n42849 , n42850 , n42851 , n220613 , n220614 , n42854 , 
     n220616 , n220617 , n42857 , n220619 , n220620 , n42860 , n220622 , n220623 , n42863 , n42864 , 
     n42865 , n42866 , n42867 , n42868 , n220630 , n220631 , n42871 , n42872 , n42873 , n42874 , 
     n42875 , n42876 , n42877 , n42878 , n42879 , n42880 , n220642 , n220643 , n42883 , n42884 , 
     n42885 , n42886 , n42887 , n42888 , n42889 , n42890 , n220652 , n220653 , n42893 , n220655 , 
     n220656 , n42896 , n42897 , n42898 , n42899 , n42900 , n42901 , n42902 , n42903 , n42904 , 
     n42905 , n220667 , n220668 , n42908 , n42909 , n42910 , n42911 , n42912 , n42913 , n42914 , 
     n42915 , n42916 , n42917 , n220679 , n220680 , n42920 , n42921 , n42922 , n42923 , n42924 , 
     n42925 , n42926 , n42927 , n220689 , n220690 , n42930 , n42931 , n42932 , n42933 , n42934 , 
     n42935 , n42936 , n42937 , n42938 , n42939 , n42940 , n42941 , n42942 , n42943 , n42944 , 
     n42945 , n42946 , n42947 , n42948 , n42949 , n42950 , n42951 , n42952 , n220714 , n220715 , 
     n42955 , n42956 , n42957 , n42958 , n42959 , n42960 , n42961 , n42962 , n42963 , n220725 , 
     n220726 , n42966 , n42967 , n42968 , n42969 , n42970 , n42971 , n42972 , n42973 , n42974 , 
     n42975 , n220737 , n220738 , n42978 , n42979 , n42980 , n42981 , n42982 , n42983 , n42984 , 
     n42985 , n42986 , n42987 , n220749 , n220750 , n42990 , n42991 , n42992 , n42993 , n42994 , 
     n42995 , n42996 , n42997 , n42998 , n42999 , n220761 , n220762 , n43002 , n43003 , n43004 , 
     n43005 , n43006 , n43007 , n220769 , n220770 , n43010 , n43011 , n43012 , n43013 , n43014 , 
     n43015 , n43016 , n43017 , n220779 , n220780 , n43020 , n43021 , n43022 , n43023 , n43024 , 
     n43025 , n43026 , n43027 , n43028 , n43029 , n43030 , n220792 , n220793 , n43033 , n43034 , 
     n43035 , n43036 , n43037 , n43038 , n43039 , n43040 , n43041 , n43042 , n220804 , n220805 , 
     n43045 , n43046 , n43047 , n43048 , n43049 , n43050 , n43051 , n43052 , n220814 , n220815 , 
     n43055 , n43056 , n43057 , n43058 , n43059 , n43060 , n43061 , n43062 , n43063 , n43064 , 
     n220826 , n220827 , n43067 , n43068 , n43069 , n43070 , n43071 , n43072 , n43073 , n43074 , 
     n220836 , n220837 , n43077 , n43078 , n43079 , n43080 , n43081 , n43082 , n220844 , n220845 , 
     n43085 , n43086 , n43087 , n43088 , n220850 , n220851 , n43091 , n43092 , n43093 , n43094 , 
     n43095 , n43096 , n43097 , n43098 , n43099 , n43100 , n43101 , n220863 , n220864 , n43104 , 
     n43105 , n43106 , n220868 , n220869 , n43109 , n43110 , n43111 , n43112 , n43113 , n43114 , 
     n43115 , n43116 , n220878 , n220879 , n43119 , n43120 , n43121 , n43122 , n43123 , n43124 , 
     n220886 , n220887 , n43127 , n220889 , n220890 , n43130 , n220892 , n220893 , n43133 , n220895 , 
     n220896 , n43136 , n43137 , n43138 , n43139 , n43140 , n43141 , n43142 , n43143 , n220905 , 
     n220906 , n43146 , n43147 , n43148 , n43149 , n43150 , n43151 , n43152 , n43153 , n43154 , 
     n43155 , n220917 , n220918 , n43158 , n43159 , n43160 , n43161 , n43162 , n43163 , n43164 , 
     n43165 , n43166 , n43167 , n220929 , n220930 , n43170 , n220932 , n220933 , n43173 , n43174 , 
     n43175 , n43176 , n43177 , n43178 , n43179 , n43180 , n43181 , n43182 , n220944 , n220945 , 
     n43185 , n43186 , n43187 , n43188 , n43189 , n43190 , n220952 , n220953 , n43193 , n43194 , 
     n43195 , n43196 , n43197 , n43198 , n43199 , n43200 , n43201 , n43202 , n220964 , n220965 , 
     n43205 , n43206 , n43207 , n43208 , n43209 , n43210 , n43211 , n43212 , n43213 , n43214 , 
     n220976 , n220977 , n43217 , n43218 , n43219 , n43220 , n43221 , n43222 , n220984 , n220985 , 
     n43225 , n43226 , n43227 , n43228 , n43229 , n43230 , n43231 , n220993 , n220994 , n43234 , 
     n43235 , n43236 , n43237 , n43238 , n43239 , n43240 , n43241 , n43242 , n43243 , n43244 , 
     n221006 , n221007 , n43247 , n43248 , n43249 , n43250 , n43251 , n43252 , n221014 , n221015 , 
     n43255 , n43256 , n43257 , n43258 , n43259 , n43260 , n43261 , n43262 , n43263 , n43264 , 
     n43265 , n43266 , n43267 , n43268 , n43269 , n43270 , n43271 , n43272 , n43273 , n43274 , 
     n43275 , n43276 , n43277 , n43278 , n43279 , n43280 , n43281 , n43282 , n43283 , n43284 , 
     n43285 , n43286 , n43287 , n221049 , n221050 , n43290 , n43291 , n43292 , n43293 , n43294 , 
     n43295 , n43296 , n43297 , n43298 , n43299 , n221061 , n221062 , n43302 , n43303 , n43304 , 
     n43305 , n43306 , n43307 , n221069 , n221070 , n43310 , n43311 , n43312 , n43313 , n43314 , 
     n43315 , n43316 , n43317 , n43318 , n43319 , n221081 , n221082 , n43322 , n43323 , n43324 , 
     n43325 , n43326 , n43327 , n43328 , n43329 , n221091 , n221092 , n43332 , n221094 , n221095 , 
     n43335 , n43336 , n43337 , n43338 , n43339 , n43340 , n43341 , n43342 , n43343 , n43344 , 
     n221106 , n221107 , n43347 , n43348 , n43349 , n43350 , n43351 , n43352 , n43353 , n221115 , 
     n221116 , n221117 , n221118 , n43358 , n221120 , n221121 , n43361 , n43362 , n43363 , n43364 , 
     n43365 , n43366 , n221128 , n221129 , n43369 , n43370 , n43371 , n43372 , n43373 , n43374 , 
     n43375 , n43376 , n221138 , n221139 , n43379 , n43380 , n43381 , n43382 , n43383 , n43384 , 
     n43385 , n43386 , n221148 , n221149 , n43389 , n43390 , n43391 , n43392 , n221154 , n221155 , 
     n43395 , n43396 , n43397 , n43398 , n43399 , n43400 , n43401 , n43402 , n43403 , n43404 , 
     n221166 , n221167 , n43407 , n43408 , n43409 , n43410 , n43411 , n43412 , n43413 , n43414 , 
     n43415 , n43416 , n221178 , n221179 , n43419 , n43420 , n43421 , n43422 , n43423 , n43424 , 
     n43425 , n43426 , n43427 , n43428 , n221190 , n221191 , n43431 , n43432 , n43433 , n43434 , 
     n221196 , n221197 , n43437 , n43438 , n43439 , n43440 , n43441 , n43442 , n221204 , n221205 , 
     n43445 , n43446 , n43447 , n43448 , n43449 , n43450 , n43451 , n43452 , n43453 , n43454 , 
     n43455 , n43456 , n43457 , n43458 , n43459 , n43460 , n43461 , n43462 , n43463 , n43464 , 
     n43465 , n43466 , n43467 , n43468 , n43469 , n43470 , n221232 , n221233 , n43473 , n43474 , 
     n43475 , n43476 , n43477 , n43478 , n43479 , n43480 , n43481 , n43482 , n43483 , n43484 , 
     n43485 , n43486 , n43487 , n43488 , n43489 , n43490 , n43491 , n43492 , n43493 , n43494 , 
     n43495 , n43496 , n43497 , n43498 , n43499 , n43500 , n43501 , n221263 , n221264 , n43504 , 
     n43505 , n43506 , n43507 , n43508 , n43509 , n221271 , n221272 , n43512 , n43513 , n43514 , 
     n43515 , n43516 , n43517 , n221279 , n221280 , n221281 , n221282 , n43522 , n43523 , n43524 , 
     n43525 , n43526 , n43527 , n43528 , n43529 , n221291 , n221292 , n43532 , n43533 , n43534 , 
     n43535 , n43536 , n43537 , n43538 , n43539 , n43540 , n43541 , n221303 , n221304 , n43544 , 
     n43545 , n43546 , n43547 , n43548 , n43549 , n43550 , n221312 , n221313 , n43553 , n43554 , 
     n43555 , n43556 , n43557 , n43558 , n221320 , n221321 , n43561 , n221323 , n221324 , n43564 , 
     n43565 , n43566 , n43567 , n43568 , n43569 , n43570 , n43571 , n43572 , n43573 , n221335 , 
     n221336 , n43576 , n43577 , n221339 , n221340 , n43580 , n43581 , n43582 , n43583 , n43584 , 
     n43585 , n43586 , n43587 , n43588 , n43589 , n43590 , n43591 , n221353 , n221354 , n43594 , 
     n43595 , n43596 , n43597 , n43598 , n43599 , n43600 , n221362 , n221363 , n43603 , n221365 , 
     n221366 , n43606 , n221368 , n221369 , n43609 , n43610 , n43611 , n43612 , n43613 , n43614 , 
     n43615 , n43616 , n221378 , n221379 , n43619 , n43620 , n43621 , n43622 , n43623 , n43624 , 
     n43625 , n43626 , n43627 , n43628 , n221390 , n221391 , n43631 , n43632 , n43633 , n43634 , 
     n43635 , n43636 , n43637 , n43638 , n43639 , n43640 , n221402 , n221403 , n43643 , n43644 , 
     n43645 , n221407 , n221408 , n43648 , n43649 , n43650 , n43651 , n43652 , n43653 , n43654 , 
     n43655 , n43656 , n43657 , n221419 , n221420 , n43660 , n43661 , n43662 , n43663 , n43664 , 
     n43665 , n43666 , n43667 , n43668 , n43669 , n221431 , n221432 , n43672 , n221434 , n221435 , 
     n43675 , n221437 , n221438 , n43678 , n43679 , n43680 , n43681 , n43682 , n43683 , n43684 , 
     n43685 , n221447 , n221448 , n43688 , n43689 , n43690 , n43691 , n43692 , n43693 , n43694 , 
     n43695 , n43696 , n43697 , n221459 , n221460 , n43700 , n221462 , n221463 , n43703 , n43704 , 
     n43705 , n43706 , n43707 , n43708 , n43709 , n43710 , n43711 , n43712 , n43713 , n43714 , 
     n43715 , n43716 , n221478 , n221479 , n43719 , n43720 , n43721 , n43722 , n43723 , n43724 , 
     n43725 , n43726 , n43727 , n43728 , n43729 , n221491 , n221492 , n43732 , n43733 , n43734 , 
     n43735 , n43736 , n43737 , n43738 , n43739 , n43740 , n221502 , n221503 , n43743 , n43744 , 
     n43745 , n43746 , n43747 , n43748 , n43749 , n43750 , n43751 , n43752 , n221514 , n221515 , 
     n43755 , n43756 , n43757 , n43758 , n43759 , n221521 , n221522 , n43762 , n43763 , n43764 , 
     n43765 , n43766 , n43767 , n43768 , n43769 , n43770 , n43771 , n43772 , n43773 , n221535 , 
     n221536 , n221537 , n221538 , n43778 , n43779 , n43780 , n43781 , n221543 , n221544 , n43784 , 
     n221546 , n221547 , n43787 , n43788 , n43789 , n43790 , n43791 , n43792 , n221554 , n221555 , 
     n43795 , n43796 , n43797 , n43798 , n43799 , n43800 , n43801 , n43802 , n43803 , n43804 , 
     n221566 , n221567 , n43807 , n43808 , n43809 , n43810 , n43811 , n43812 , n43813 , n43814 , 
     n43815 , n43816 , n221578 , n221579 , n43819 , n43820 , n43821 , n43822 , n43823 , n43824 , 
     n43825 , n43826 , n43827 , n43828 , n221590 , n221591 , n43831 , n43832 , n43833 , n43834 , 
     n221596 , n221597 , n43837 , n43838 , n43839 , n43840 , n43841 , n43842 , n221604 , n221605 , 
     n43845 , n43846 , n43847 , n43848 , n43849 , n43850 , n43851 , n43852 , n221614 , n221615 , 
     n43855 , n43856 , n43857 , n43858 , n43859 , n43860 , n43861 , n43862 , n221624 , n221625 , 
     n43865 , n43866 , n221628 , n221629 , n43869 , n43870 , n43871 , n43872 , n43873 , n43874 , 
     n43875 , n43876 , n43877 , n43878 , n43879 , n221641 , n221642 , n43882 , n221644 , n221645 , 
     n43885 , n43886 , n43887 , n43888 , n43889 , n43890 , n221652 , n221653 , n43893 , n43894 , 
     n43895 , n43896 , n221658 , n221659 , n43899 , n43900 , n43901 , n43902 , n43903 , n43904 , 
     n43905 , n43906 , n221668 , n221669 , n43909 , n43910 , n43911 , n43912 , n43913 , n43914 , 
     n43915 , n43916 , n43917 , n43918 , n221680 , n221681 , n43921 , n43922 , n43923 , n43924 , 
     n43925 , n43926 , n43927 , n43928 , n43929 , n43930 , n221692 , n221693 , n43933 , n43934 , 
     n43935 , n43936 , n43937 , n43938 , n43939 , n43940 , n221702 , n221703 , n43943 , n43944 , 
     n43945 , n43946 , n43947 , n43948 , n43949 , n43950 , n43951 , n43952 , n221714 , n221715 , 
     n43955 , n43956 , n43957 , n43958 , n43959 , n43960 , n43961 , n43962 , n43963 , n43964 , 
     n221726 , n221727 , n43967 , n43968 , n43969 , n43970 , n43971 , n43972 , n43973 , n43974 , 
     n43975 , n43976 , n221738 , n221739 , n43979 , n43980 , n43981 , n43982 , n43983 , n43984 , 
     n43985 , n43986 , n43987 , n43988 , n43989 , n43990 , n43991 , n43992 , n43993 , n43994 , 
     n43995 , n43996 , n43997 , n43998 , n43999 , n221761 , n221762 , n44002 , n44003 , n44004 , 
     n44005 , n44006 , n44007 , n221769 , n221770 , n44010 , n44011 , n44012 , n44013 , n221775 , 
     n221776 , n44016 , n221778 , n221779 , n44019 , n44020 , n44021 , n44022 , n221784 , n221785 , 
     n221786 , n221787 , n44027 , n44028 , n44029 , n44030 , n44031 , n44032 , n221794 , n221795 , 
     n44035 , n44036 , n44037 , n44038 , n44039 , n44040 , n44041 , n44042 , n221804 , n221805 , 
     n44045 , n221807 , n221808 , n44048 , n44049 , n44050 , n44051 , n44052 , n44053 , n221815 , 
     n221816 , n44056 , n44057 , n44058 , n44059 , n44060 , n44061 , n221823 , n221824 , n44064 , 
     n221826 , n221827 , n44067 , n44068 , n44069 , n44070 , n44071 , n44072 , n44073 , n44074 , 
     n221836 , n221837 , n44077 , n44078 , n44079 , n44080 , n221842 , n221843 , n44083 , n44084 , 
     n44085 , n44086 , n44087 , n44088 , n44089 , n44090 , n221852 , n221853 , n44093 , n44094 , 
     n44095 , n44096 , n44097 , n44098 , n44099 , n44100 , n44101 , n44102 , n221864 , n221865 , 
     n44105 , n44106 , n44107 , n44108 , n44109 , n44110 , n221872 , n221873 , n44113 , n44114 , 
     n44115 , n44116 , n44117 , n44118 , n221880 , n221881 , n44121 , n221883 , n221884 , n44124 , 
     n44125 , n44126 , n44127 , n44128 , n44129 , n221891 , n221892 , n44132 , n44133 , n44134 , 
     n44135 , n44136 , n44137 , n44138 , n44139 , n44140 , n44141 , n44142 , n44143 , n44144 , 
     n44145 , n44146 , n44147 , n44148 , n44149 , n44150 , n44151 , n44152 , n44153 , n44154 , 
     n221916 , n221917 , n44157 , n44158 , n44159 , n44160 , n44161 , n44162 , n44163 , n44164 , 
     n44165 , n44166 , n221928 , n221929 , n44169 , n44170 , n44171 , n44172 , n44173 , n44174 , 
     n44175 , n44176 , n44177 , n44178 , n221940 , n221941 , n44181 , n44182 , n44183 , n44184 , 
     n44185 , n44186 , n44187 , n44188 , n221950 , n221951 , n44191 , n44192 , n44193 , n44194 , 
     n44195 , n44196 , n221958 , n221959 , n44199 , n44200 , n44201 , n44202 , n44203 , n44204 , 
     n44205 , n44206 , n44207 , n44208 , n221970 , n221971 , n44211 , n44212 , n44213 , n44214 , 
     n44215 , n44216 , n221978 , n221979 , n44219 , n221981 , n221982 , n44222 , n44223 , n44224 , 
     n44225 , n44226 , n44227 , n44228 , n44229 , n44230 , n44231 , n221993 , n221994 , n44234 , 
     n44235 , n44236 , n44237 , n44238 , n44239 , n222001 , n222002 , n44242 , n44243 , n44244 , 
     n44245 , n44246 , n44247 , n44248 , n44249 , n222011 , n222012 , n44252 , n222014 , n222015 , 
     n44255 , n222017 , n222018 , n44258 , n44259 , n44260 , n44261 , n222023 , n222024 , n44264 , 
     n222026 , n222027 , n44267 , n44268 , n44269 , n44270 , n222032 , n222033 , n44273 , n44274 , 
     n44275 , n44276 , n44277 , n44278 , n44279 , n44280 , n44281 , n44282 , n222044 , n222045 , 
     n44285 , n44286 , n44287 , n44288 , n44289 , n44290 , n44291 , n44292 , n222054 , n222055 , 
     n44295 , n222057 , n222058 , n44298 , n222060 , n222061 , n44301 , n44302 , n44303 , n44304 , 
     n44305 , n44306 , n44307 , n44308 , n44309 , n44310 , n222072 , n222073 , n44313 , n44314 , 
     n44315 , n44316 , n44317 , n44318 , n222080 , n222081 , n44321 , n44322 , n44323 , n44324 , 
     n44325 , n44326 , n44327 , n44328 , n222090 , n222091 , n44331 , n44332 , n44333 , n44334 , 
     n44335 , n44336 , n44337 , n44338 , n44339 , n44340 , n222102 , n222103 , n44343 , n44344 , 
     n44345 , n44346 , n44347 , n44348 , n44349 , n44350 , n44351 , n44352 , n44353 , n44354 , 
     n222116 , n222117 , n44357 , n44358 , n44359 , n44360 , n222122 , n222123 , n44363 , n222125 , 
     n222126 , n44366 , n44367 , n44368 , n44369 , n44370 , n44371 , n222133 , n222134 , n44374 , 
     n222136 , n222137 , n44377 , n44378 , n44379 , n44380 , n44381 , n44382 , n44383 , n44384 , 
     n222146 , n222147 , n44387 , n44388 , n44389 , n44390 , n44391 , n44392 , n44393 , n44394 , 
     n44395 , n44396 , n222158 , n222159 , n44399 , n222161 , n222162 , n44402 , n44403 , n44404 , 
     n44405 , n44406 , n44407 , n44408 , n44409 , n44410 , n44411 , n44412 , n44413 , n222175 , 
     n222176 , n44416 , n44417 , n44418 , n44419 , n44420 , n44421 , n222183 , n222184 , n44424 , 
     n44425 , n44426 , n44427 , n222189 , n222190 , n44430 , n44431 , n44432 , n44433 , n44434 , 
     n44435 , n44436 , n44437 , n44438 , n44439 , n222201 , n222202 , n44442 , n222204 , n222205 , 
     n44445 , n44446 , n44447 , n44448 , n44449 , n44450 , n44451 , n44452 , n44453 , n44454 , 
     n222216 , n222217 , n44457 , n44458 , n44459 , n44460 , n44461 , n44462 , n44463 , n44464 , 
     n44465 , n44466 , n222228 , n222229 , n44469 , n44470 , n44471 , n44472 , n44473 , n44474 , 
     n44475 , n44476 , n44477 , n44478 , n222240 , n222241 , n44481 , n44482 , n44483 , n44484 , 
     n44485 , n44486 , n222248 , n222249 , n44489 , n222251 , n222252 , n44492 , n44493 , n44494 , 
     n44495 , n44496 , n44497 , n44498 , n44499 , n44500 , n44501 , n44502 , n44503 , n222265 , 
     n222266 , n44506 , n44507 , n222269 , n222270 , n44510 , n44511 , n44512 , n44513 , n44514 , 
     n44515 , n44516 , n44517 , n44518 , n44519 , n222281 , n222282 , n44522 , n44523 , n44524 , 
     n44525 , n44526 , n44527 , n44528 , n44529 , n44530 , n44531 , n222293 , n222294 , n44534 , 
     n44535 , n44536 , n44537 , n44538 , n44539 , n222301 , n222302 , n44542 , n222304 , n222305 , 
     n44545 , n44546 , n44547 , n44548 , n44549 , n44550 , n44551 , n44552 , n222314 , n222315 , 
     n44555 , n44556 , n44557 , n44558 , n44559 , n44560 , n44561 , n44562 , n222324 , n222325 , 
     n44565 , n222327 , n222328 , n44568 , n44569 , n44570 , n44571 , n44572 , n44573 , n44574 , 
     n44575 , n44576 , n44577 , n222339 , n222340 , n44580 , n44581 , n44582 , n44583 , n44584 , 
     n44585 , n44586 , n44587 , n222349 , n222350 , n44590 , n44591 , n44592 , n44593 , n44594 , 
     n44595 , n222357 , n222358 , n44598 , n44599 , n44600 , n44601 , n44602 , n44603 , n44604 , 
     n44605 , n222367 , n222368 , n44608 , n222370 , n222371 , n44611 , n44612 , n44613 , n44614 , 
     n44615 , n44616 , n44617 , n44618 , n44619 , n44620 , n222382 , n222383 , n44623 , n44624 , 
     n44625 , n44626 , n44627 , n44628 , n44629 , n44630 , n222392 , n222393 , n44633 , n44634 , 
     n222396 , n222397 , n44637 , n44638 , n44639 , n44640 , n222402 , n222403 , n44643 , n44644 , 
     n44645 , n44646 , n44647 , n44648 , n44649 , n44650 , n222412 , n222413 , n44653 , n44654 , 
     n44655 , n44656 , n44657 , n222419 , n222420 , n44660 , n44661 , n44662 , n44663 , n44664 , 
     n44665 , n44666 , n44667 , n222429 , n222430 , n44670 , n44671 , n44672 , n44673 , n222435 , 
     n222436 , n44676 , n44677 , n222439 , n222440 , n44680 , n222442 , n222443 , n44683 , n44684 , 
     n44685 , n44686 , n44687 , n44688 , n44689 , n44690 , n44691 , n44692 , n222454 , n222455 , 
     n44695 , n44696 , n44697 , n44698 , n44699 , n44700 , n222462 , n222463 , n44703 , n44704 , 
     n44705 , n44706 , n44707 , n44708 , n222470 , n222471 , n44711 , n44712 , n44713 , n44714 , 
     n44715 , n44716 , n222478 , n222479 , n44719 , n44720 , n44721 , n44722 , n44723 , n44724 , 
     n222486 , n222487 , n44727 , n44728 , n44729 , n44730 , n44731 , n44732 , n44733 , n44734 , 
     n222496 , n222497 , n44737 , n44738 , n44739 , n44740 , n44741 , n44742 , n222504 , n222505 , 
     n44745 , n44746 , n44747 , n44748 , n44749 , n44750 , n222512 , n222513 , n44753 , n44754 , 
     n44755 , n44756 , n44757 , n44758 , n44759 , n44760 , n44761 , n44762 , n222524 , n222525 , 
     n44765 , n44766 , n44767 , n44768 , n44769 , n222531 , n222532 , n222533 , n222534 , n44774 , 
     n222536 , n222537 , n44777 , n44778 , n44779 , n44780 , n44781 , n44782 , n44783 , n44784 , 
     n44785 , n44786 , n222548 , n222549 , n44789 , n44790 , n44791 , n44792 , n44793 , n44794 , 
     n222556 , n222557 , n44797 , n44798 , n44799 , n44800 , n44801 , n44802 , n44803 , n44804 , 
     n222566 , n222567 , n44807 , n44808 , n44809 , n44810 , n44811 , n44812 , n44813 , n44814 , 
     n222576 , n222577 , n44817 , n222579 , n222580 , n44820 , n222582 , n222583 , n44823 , n222585 , 
     n222586 , n44826 , n222588 , n222589 , n44829 , n44830 , n44831 , n44832 , n44833 , n44834 , 
     n222596 , n222597 , n44837 , n222599 , n222600 , n44840 , n222602 , n222603 , n44843 , n44844 , 
     n44845 , n44846 , n44847 , n44848 , n44849 , n44850 , n44851 , n44852 , n222614 , n222615 , 
     n44855 , n44856 , n44857 , n44858 , n44859 , n44860 , n222622 , n222623 , n44863 , n222625 , 
     n222626 , n44866 , n222628 , n222629 , n44869 , n222631 , n222632 , n44872 , n44873 , n44874 , 
     n44875 , n44876 , n44877 , n44878 , n44879 , n44880 , n44881 , n222643 , n222644 , n44884 , 
     n44885 , n44886 , n44887 , n44888 , n44889 , n44890 , n44891 , n44892 , n44893 , n222655 , 
     n222656 , n44896 , n44897 , n44898 , n44899 , n44900 , n44901 , n44902 , n44903 , n44904 , 
     n44905 , n222667 , n222668 , n44908 , n44909 , n44910 , n44911 , n44912 , n44913 , n44914 , 
     n44915 , n44916 , n44917 , n222679 , n222680 , n44920 , n44921 , n44922 , n44923 , n44924 , 
     n44925 , n222687 , n222688 , n44928 , n44929 , n44930 , n44931 , n44932 , n44933 , n44934 , 
     n44935 , n44936 , n44937 , n222699 , n222700 , n44940 , n44941 , n44942 , n44943 , n44944 , 
     n44945 , n44946 , n44947 , n222709 , n222710 , n44950 , n44951 , n44952 , n44953 , n44954 , 
     n44955 , n222717 , n222718 , n44958 , n222720 , n222721 , n44961 , n44962 , n44963 , n44964 , 
     n44965 , n44966 , n222728 , n222729 , n44969 , n44970 , n44971 , n44972 , n44973 , n44974 , 
     n44975 , n44976 , n44977 , n44978 , n222740 , n222741 , n44981 , n44982 , n44983 , n44984 , 
     n44985 , n44986 , n44987 , n44988 , n44989 , n44990 , n222752 , n222753 , n44993 , n44994 , 
     n44995 , n44996 , n44997 , n44998 , n44999 , n222761 , n222762 , n45002 , n45003 , n45004 , 
     n45005 , n45006 , n45007 , n45008 , n45009 , n45010 , n45011 , n222773 , n222774 , n45014 , 
     n45015 , n45016 , n45017 , n45018 , n45019 , n45020 , n222782 , n222783 , n45023 , n45024 , 
     n45025 , n45026 , n45027 , n45028 , n222790 , n222791 , n45031 , n222793 , n222794 , n45034 , 
     n222796 , n222797 , n45037 , n45038 , n45039 , n45040 , n45041 , n45042 , n45043 , n45044 , 
     n45045 , n45046 , n222808 , n222809 , n45049 , n45050 , n45051 , n45052 , n222814 , n222815 , 
     n45055 , n222817 , n222818 , n45058 , n222820 , n45060 , n45061 , n45062 , n45063 , n45064 , 
     n45065 , n222827 , n222828 , n45068 , n45069 , n45070 , n45071 , n45072 , n45073 , n45074 , 
     n45075 , n45076 , n45077 , n222839 , n222840 , n45080 , n45081 , n45082 , n45083 , n45084 , 
     n45085 , n45086 , n45087 , n45088 , n45089 , n222851 , n222852 , n45092 , n45093 , n45094 , 
     n45095 , n45096 , n45097 , n222859 , n222860 , n45100 , n45101 , n45102 , n45103 , n222865 , 
     n222866 , n45106 , n45107 , n45108 , n45109 , n45110 , n45111 , n45112 , n45113 , n45114 , 
     n45115 , n222877 , n222878 , n45118 , n45119 , n45120 , n45121 , n222883 , n222884 , n45124 , 
     n222886 , n222887 , n45127 , n45128 , n45129 , n45130 , n45131 , n45132 , n45133 , n45134 , 
     n45135 , n45136 , n222898 , n222899 , n45139 , n45140 , n45141 , n45142 , n45143 , n45144 , 
     n45145 , n45146 , n222908 , n222909 , n45149 , n222911 , n222912 , n45152 , n45153 , n45154 , 
     n45155 , n45156 , n45157 , n45158 , n45159 , n222921 , n222922 , n45162 , n45163 , n45164 , 
     n45165 , n45166 , n45167 , n222929 , n222930 , n45170 , n45171 , n45172 , n45173 , n45174 , 
     n45175 , n45176 , n45177 , n222939 , n222940 , n45180 , n45181 , n45182 , n45183 , n45184 , 
     n45185 , n45186 , n45187 , n222949 , n222950 , n45190 , n45191 , n45192 , n45193 , n45194 , 
     n45195 , n45196 , n45197 , n45198 , n45199 , n222961 , n222962 , n45202 , n45203 , n45204 , 
     n45205 , n45206 , n45207 , n222969 , n222970 , n45210 , n45211 , n45212 , n45213 , n45214 , 
     n45215 , n45216 , n45217 , n45218 , n45219 , n222981 , n222982 , n45222 , n45223 , n45224 , 
     n45225 , n45226 , n45227 , n45228 , n45229 , n45230 , n45231 , n222993 , n222994 , n45234 , 
     n222996 , n222997 , n45237 , n45238 , n45239 , n45240 , n45241 , n45242 , n223004 , n223005 , 
     n45245 , n45246 , n45247 , n45248 , n45249 , n45250 , n45251 , n45252 , n45253 , n223015 , 
     n223016 , n45256 , n223018 , n223019 , n45259 , n45260 , n45261 , n45262 , n45263 , n45264 , 
     n223026 , n223027 , n45267 , n45268 , n45269 , n45270 , n45271 , n45272 , n223034 , n223035 , 
     n45275 , n45276 , n45277 , n45278 , n45279 , n45280 , n45281 , n45282 , n45283 , n45284 , 
     n45285 , n45286 , n223048 , n223049 , n45289 , n45290 , n45291 , n45292 , n45293 , n45294 , 
     n223056 , n223057 , n45297 , n45298 , n45299 , n45300 , n45301 , n45302 , n223064 , n223065 , 
     n45305 , n45306 , n45307 , n45308 , n45309 , n45310 , n45311 , n45312 , n45313 , n45314 , 
     n223076 , n223077 , n45317 , n45318 , n45319 , n45320 , n45321 , n45322 , n45323 , n45324 , 
     n45325 , n45326 , n223088 , n223089 , n45329 , n45330 , n45331 , n45332 , n45333 , n45334 , 
     n45335 , n45336 , n223098 , n223099 , n45339 , n45340 , n45341 , n45342 , n223104 , n223105 , 
     n45345 , n223107 , n223108 , n45348 , n223110 , n223111 , n45351 , n45352 , n45353 , n45354 , 
     n223116 , n223117 , n45357 , n45358 , n45359 , n45360 , n45361 , n45362 , n223124 , n223125 , 
     n45365 , n45366 , n45367 , n45368 , n45369 , n45370 , n45371 , n45372 , n45373 , n45374 , 
     n223136 , n223137 , n45377 , n223139 , n223140 , n45380 , n45381 , n45382 , n45383 , n45384 , 
     n45385 , n45386 , n45387 , n45388 , n45389 , n45390 , n223152 , n223153 , n45393 , n223155 , 
     n223156 , n45396 , n45397 , n45398 , n45399 , n45400 , n45401 , n223163 , n223164 , n45404 , 
     n223166 , n223167 , n45407 , n45408 , n45409 , n45410 , n223172 , n223173 , n45413 , n45414 , 
     n45415 , n45416 , n45417 , n45418 , n45419 , n45420 , n45421 , n45422 , n223184 , n223185 , 
     n45425 , n45426 , n45427 , n45428 , n223190 , n223191 , n45431 , n223193 , n223194 , n45434 , 
     n45435 , n45436 , n45437 , n45438 , n45439 , n45440 , n45441 , n45442 , n45443 , n223205 , 
     n223206 , n45446 , n45447 , n223209 , n223210 , n45450 , n45451 , n45452 , n45453 , n45454 , 
     n45455 , n45456 , n45457 , n45458 , n223220 , n223221 , n45461 , n45462 , n45463 , n45464 , 
     n45465 , n45466 , n45467 , n45468 , n223230 , n223231 , n45471 , n45472 , n45473 , n45474 , 
     n45475 , n45476 , n45477 , n45478 , n223240 , n223241 , n45481 , n45482 , n45483 , n45484 , 
     n45485 , n45486 , n45487 , n45488 , n45489 , n45490 , n223252 , n223253 , n45493 , n223255 , 
     n223256 , n45496 , n45497 , n45498 , n45499 , n45500 , n45501 , n45502 , n45503 , n223265 , 
     n223266 , n45506 , n45507 , n45508 , n45509 , n223271 , n223272 , n45512 , n45513 , n45514 , 
     n45515 , n45516 , n45517 , n45518 , n45519 , n45520 , n45521 , n223283 , n223284 , n45524 , 
     n223286 , n223287 , n45527 , n45528 , n45529 , n45530 , n45531 , n45532 , n45533 , n45534 , 
     n45535 , n45536 , n223298 , n223299 , n45539 , n45540 , n45541 , n45542 , n45543 , n45544 , 
     n45545 , n45546 , n45547 , n45548 , n223310 , n223311 , n45551 , n223313 , n223314 , n45554 , 
     n45555 , n45556 , n45557 , n45558 , n45559 , n223321 , n223322 , n45562 , n45563 , n45564 , 
     n45565 , n45566 , n45567 , n223329 , n223330 , n45570 , n45571 , n45572 , n45573 , n45574 , 
     n45575 , n223337 , n223338 , n45578 , n45579 , n45580 , n45581 , n45582 , n45583 , n45584 , 
     n45585 , n45586 , n45587 , n45588 , n45589 , n45590 , n45591 , n45592 , n45593 , n223355 , 
     n223356 , n45596 , n45597 , n45598 , n45599 , n45600 , n45601 , n45602 , n45603 , n45604 , 
     n45605 , n45606 , n223368 , n223369 , n45609 , n45610 , n45611 , n45612 , n45613 , n45614 , 
     n45615 , n45616 , n45617 , n45618 , n45619 , n223381 , n223382 , n45622 , n45623 , n45624 , 
     n45625 , n45626 , n45627 , n45628 , n45629 , n45630 , n45631 , n223393 , n223394 , n45634 , 
     n223396 , n223397 , n45637 , n223399 , n223400 , n45640 , n45641 , n45642 , n45643 , n45644 , 
     n45645 , n223407 , n223408 , n45648 , n45649 , n45650 , n45651 , n45652 , n45653 , n223415 , 
     n223416 , n45656 , n45657 , n45658 , n45659 , n223421 , n223422 , n45662 , n223424 , n223425 , 
     n45665 , n45666 , n45667 , n45668 , n45669 , n45670 , n45671 , n45672 , n45673 , n45674 , 
     n223436 , n223437 , n45677 , n45678 , n45679 , n45680 , n45681 , n45682 , n223444 , n223445 , 
     n45685 , n45686 , n45687 , n45688 , n45689 , n45690 , n45691 , n45692 , n223454 , n223455 , 
     n45695 , n45696 , n45697 , n45698 , n45699 , n45700 , n45701 , n45702 , n223464 , n223465 , 
     n45705 , n223467 , n223468 , n45708 , n45709 , n45710 , n45711 , n223473 , n223474 , n45714 , 
     n45715 , n45716 , n45717 , n45718 , n45719 , n45720 , n45721 , n45722 , n45723 , n223485 , 
     n223486 , n45726 , n45727 , n45728 , n45729 , n45730 , n45731 , n45732 , n45733 , n45734 , 
     n45735 , n223497 , n223498 , n45738 , n45739 , n45740 , n45741 , n223503 , n223504 , n45744 , 
     n223506 , n223507 , n45747 , n223509 , n223510 , n45750 , n45751 , n45752 , n45753 , n45754 , 
     n45755 , n45756 , n45757 , n223519 , n223520 , n45760 , n45761 , n45762 , n45763 , n45764 , 
     n45765 , n45766 , n45767 , n223529 , n223530 , n45770 , n45771 , n45772 , n45773 , n223535 , 
     n223536 , n45776 , n45777 , n45778 , n45779 , n45780 , n45781 , n45782 , n45783 , n45784 , 
     n223546 , n223547 , n45787 , n45788 , n45789 , n45790 , n45791 , n45792 , n45793 , n45794 , 
     n45795 , n45796 , n223558 , n223559 , n45799 , n223561 , n223562 , n45802 , n45803 , n45804 , 
     n45805 , n45806 , n45807 , n45808 , n45809 , n45810 , n45811 , n223573 , n223574 , n45814 , 
     n45815 , n45816 , n45817 , n45818 , n45819 , n45820 , n45821 , n223583 , n223584 , n45824 , 
     n45825 , n45826 , n45827 , n45828 , n45829 , n45830 , n45831 , n45832 , n45833 , n223595 , 
     n223596 , n45836 , n45837 , n45838 , n45839 , n45840 , n45841 , n223603 , n223604 , n45844 , 
     n45845 , n45846 , n45847 , n45848 , n45849 , n45850 , n45851 , n223613 , n223614 , n45854 , 
     n45855 , n45856 , n45857 , n45858 , n45859 , n223621 , n223622 , n45862 , n45863 , n45864 , 
     n45865 , n223627 , n223628 , n45868 , n223630 , n223631 , n45871 , n45872 , n45873 , n45874 , 
     n45875 , n45876 , n45877 , n45878 , n45879 , n45880 , n223642 , n223643 , n45883 , n45884 , 
     n45885 , n45886 , n45887 , n45888 , n223650 , n223651 , n45891 , n223653 , n223654 , n45894 , 
     n45895 , n45896 , n45897 , n45898 , n45899 , n223661 , n223662 , n45902 , n45903 , n45904 , 
     n45905 , n45906 , n45907 , n223669 , n223670 , n45910 , n45911 , n45912 , n45913 , n45914 , 
     n45915 , n45916 , n45917 , n223679 , n223680 , n45920 , n45921 , n45922 , n45923 , n45924 , 
     n45925 , n45926 , n45927 , n45928 , n45929 , n223691 , n223692 , n45932 , n45933 , n45934 , 
     n45935 , n45936 , n45937 , n223699 , n223700 , n45940 , n45941 , n45942 , n45943 , n45944 , 
     n45945 , n45946 , n45947 , n45948 , n45949 , n223711 , n223712 , n45952 , n45953 , n45954 , 
     n45955 , n45956 , n45957 , n223719 , n223720 , n45960 , n45961 , n45962 , n45963 , n45964 , 
     n45965 , n223727 , n223728 , n45968 , n223730 , n223731 , n45971 , n45972 , n45973 , n45974 , 
     n223736 , n223737 , n45977 , n45978 , n45979 , n45980 , n45981 , n45982 , n45983 , n45984 , 
     n223746 , n223747 , n45987 , n45988 , n45989 , n45990 , n223752 , n223753 , n45993 , n45994 , 
     n45995 , n45996 , n45997 , n45998 , n45999 , n46000 , n46001 , n46002 , n223764 , n223765 , 
     n46005 , n46006 , n46007 , n46008 , n46009 , n46010 , n46011 , n46012 , n46013 , n223775 , 
     n223776 , n46016 , n46017 , n46018 , n46019 , n46020 , n46021 , n46022 , n223784 , n223785 , 
     n46025 , n46026 , n46027 , n46028 , n223790 , n223791 , n46031 , n223793 , n46033 , n46034 , 
     n46035 , n46036 , n46037 , n46038 , n46039 , n46040 , n46041 , n46042 , n223804 , n223805 , 
     n46045 , n46046 , n46047 , n46048 , n223810 , n223811 , n46051 , n46052 , n46053 , n46054 , 
     n223816 , n223817 , n46057 , n46058 , n46059 , n46060 , n46061 , n46062 , n46063 , n46064 , 
     n223826 , n223827 , n46067 , n46068 , n46069 , n46070 , n46071 , n46072 , n46073 , n46074 , 
     n223836 , n223837 , n46077 , n223839 , n223840 , n46080 , n46081 , n46082 , n46083 , n46084 , 
     n46085 , n223847 , n223848 , n46088 , n223850 , n223851 , n46091 , n46092 , n46093 , n46094 , 
     n46095 , n46096 , n223858 , n223859 , n46099 , n46100 , n46101 , n46102 , n46103 , n46104 , 
     n46105 , n46106 , n223868 , n223869 , n46109 , n46110 , n46111 , n46112 , n46113 , n46114 , 
     n46115 , n46116 , n46117 , n46118 , n223880 , n223881 , n46121 , n46122 , n46123 , n46124 , 
     n223886 , n223887 , n46127 , n223889 , n223890 , n46130 , n223892 , n223893 , n46133 , n46134 , 
     n46135 , n46136 , n46137 , n46138 , n46139 , n46140 , n46141 , n46142 , n223904 , n223905 , 
     n46145 , n46146 , n46147 , n46148 , n223910 , n223911 , n46151 , n46152 , n46153 , n46154 , 
     n46155 , n46156 , n46157 , n46158 , n223920 , n223921 , n46161 , n223923 , n223924 , n46164 , 
     n46165 , n46166 , n46167 , n46168 , n46169 , n46170 , n46171 , n46172 , n46173 , n46174 , 
     n46175 , n46176 , n223938 , n223939 , n46179 , n46180 , n46181 , n46182 , n46183 , n46184 , 
     n46185 , n46186 , n46187 , n46188 , n223950 , n223951 , n46191 , n46192 , n46193 , n46194 , 
     n46195 , n46196 , n46197 , n46198 , n46199 , n46200 , n46201 , n46202 , n46203 , n46204 , 
     n223966 , n223967 , n46207 , n223969 , n223970 , n46210 , n46211 , n46212 , n46213 , n46214 , 
     n46215 , n223977 , n223978 , n46218 , n46219 , n46220 , n46221 , n46222 , n46223 , n223985 , 
     n223986 , n46226 , n46227 , n46228 , n46229 , n223991 , n46231 , n46232 , n46233 , n46234 , 
     n46235 , n46236 , n46237 , n46238 , n224000 , n224001 , n46241 , n224003 , n224004 , n46244 , 
     n46245 , n46246 , n46247 , n46248 , n46249 , n224011 , n224012 , n46252 , n46253 , n46254 , 
     n46255 , n46256 , n46257 , n46258 , n46259 , n224021 , n224022 , n46262 , n224024 , n224025 , 
     n46265 , n46266 , n46267 , n46268 , n46269 , n46270 , n46271 , n46272 , n224034 , n224035 , 
     n46275 , n46276 , n46277 , n46278 , n46279 , n46280 , n224042 , n224043 , n46283 , n224045 , 
     n224046 , n46286 , n46287 , n46288 , n46289 , n46290 , n46291 , n224053 , n224054 , n46294 , 
     n46295 , n46296 , n46297 , n224059 , n224060 , n46300 , n224062 , n224063 , n46303 , n46304 , 
     n46305 , n46306 , n224068 , n224069 , n46309 , n46310 , n46311 , n46312 , n46313 , n46314 , 
     n224076 , n224077 , n46317 , n46318 , n46319 , n46320 , n46321 , n46322 , n224084 , n224085 , 
     n46325 , n46326 , n46327 , n46328 , n224090 , n224091 , n46331 , n224093 , n224094 , n46334 , 
     n46335 , n46336 , n46337 , n224099 , n224100 , n46340 , n46341 , n46342 , n46343 , n46344 , 
     n46345 , n224107 , n224108 , n46348 , n46349 , n46350 , n46351 , n46352 , n46353 , n224115 , 
     n224116 , n46356 , n224118 , n224119 , n46359 , n224121 , n224122 , n46362 , n46363 , n46364 , 
     n46365 , n46366 , n46367 , n224129 , n224130 , n46370 , n46371 , n46372 , n46373 , n46374 , 
     n46375 , n224137 , n224138 , n46378 , n224140 , n224141 , n46381 , n46382 , n46383 , n46384 , 
     n46385 , n46386 , n224148 , n224149 , n46389 , n46390 , n46391 , n46392 , n46393 , n46394 , 
     n46395 , n46396 , n46397 , n46398 , n224160 , n224161 , n46401 , n46402 , n46403 , n46404 , 
     n46405 , n46406 , n46407 , n46408 , n224170 , n224171 , n46411 , n46412 , n46413 , n46414 , 
     n46415 , n46416 , n46417 , n224179 , n224180 , n46420 , n224182 , n224183 , n46423 , n46424 , 
     n46425 , n46426 , n46427 , n46428 , n46429 , n46430 , n46431 , n46432 , n46433 , n46434 , 
     n224196 , n224197 , n46437 , n46438 , n46439 , n46440 , n46441 , n46442 , n46443 , n46444 , 
     n224206 , n224207 , n46447 , n46448 , n46449 , n46450 , n46451 , n46452 , n224214 , n224215 , 
     n46455 , n224217 , n224218 , n46458 , n46459 , n46460 , n46461 , n46462 , n46463 , n224225 , 
     n224226 , n46466 , n46467 , n46468 , n46469 , n46470 , n46471 , n224233 , n224234 , n46474 , 
     n224236 , n224237 , n46477 , n46478 , n46479 , n46480 , n46481 , n46482 , n46483 , n224245 , 
     n224246 , n46486 , n224248 , n224249 , n46489 , n46490 , n46491 , n46492 , n224254 , n224255 , 
     n46495 , n46496 , n46497 , n46498 , n46499 , n46500 , n46501 , n46502 , n224264 , n224265 , 
     n46505 , n46506 , n46507 , n46508 , n46509 , n46510 , n224272 , n224273 , n46513 , n46514 , 
     n46515 , n46516 , n46517 , n46518 , n224280 , n224281 , n46521 , n46522 , n46523 , n46524 , 
     n46525 , n46526 , n46527 , n46528 , n46529 , n46530 , n224292 , n224293 , n46533 , n46534 , 
     n46535 , n46536 , n224298 , n224299 , n46539 , n46540 , n46541 , n46542 , n46543 , n46544 , 
     n224306 , n224307 , n46547 , n46548 , n46549 , n46550 , n46551 , n46552 , n224314 , n224315 , 
     n46555 , n46556 , n46557 , n46558 , n46559 , n46560 , n224322 , n224323 , n46563 , n46564 , 
     n46565 , n46566 , n46567 , n46568 , n224330 , n224331 , n46571 , n46572 , n46573 , n46574 , 
     n46575 , n46576 , n46577 , n46578 , n46579 , n46580 , n224342 , n224343 , n46583 , n46584 , 
     n46585 , n46586 , n46587 , n46588 , n224350 , n224351 , n46591 , n46592 , n46593 , n46594 , 
     n46595 , n46596 , n46597 , n46598 , n224360 , n224361 , n46601 , n224363 , n224364 , n46604 , 
     n46605 , n46606 , n46607 , n224369 , n224370 , n46610 , n224372 , n224373 , n46613 , n46614 , 
     n46615 , n46616 , n46617 , n46618 , n224380 , n224381 , n46621 , n224383 , n46623 , n46624 , 
     n46625 , n46626 , n46627 , n46628 , n46629 , n46630 , n46631 , n46632 , n46633 , n46634 , 
     n224396 , n224397 , n46637 , n46638 , n46639 , n46640 , n224402 , n224403 , n46643 , n46644 , 
     n46645 , n46646 , n46647 , n46648 , n46649 , n46650 , n224412 , n224413 , n46653 , n224415 , 
     n224416 , n46656 , n46657 , n46658 , n46659 , n46660 , n46661 , n46662 , n46663 , n46664 , 
     n46665 , n224427 , n224428 , n46668 , n46669 , n46670 , n46671 , n46672 , n46673 , n224435 , 
     n224436 , n46676 , n46677 , n46678 , n46679 , n46680 , n46681 , n224443 , n224444 , n46684 , 
     n46685 , n46686 , n46687 , n224449 , n224450 , n46690 , n224452 , n224453 , n46693 , n46694 , 
     n46695 , n46696 , n46697 , n46698 , n46699 , n46700 , n224462 , n224463 , n46703 , n46704 , 
     n46705 , n46706 , n46707 , n46708 , n46709 , n46710 , n224472 , n224473 , n46713 , n46714 , 
     n46715 , n46716 , n224478 , n224479 , n46719 , n46720 , n46721 , n46722 , n46723 , n46724 , 
     n46725 , n46726 , n46727 , n46728 , n224490 , n224491 , n46731 , n46732 , n46733 , n46734 , 
     n46735 , n46736 , n46737 , n46738 , n46739 , n46740 , n224502 , n224503 , n46743 , n46744 , 
     n46745 , n46746 , n46747 , n46748 , n224510 , n224511 , n46751 , n46752 , n46753 , n46754 , 
     n46755 , n46756 , n46757 , n46758 , n224520 , n224521 , n46761 , n46762 , n46763 , n46764 , 
     n46765 , n46766 , n46767 , n224529 , n224530 , n46770 , n46771 , n46772 , n46773 , n224535 , 
     n224536 , n46776 , n46777 , n46778 , n46779 , n46780 , n46781 , n46782 , n46783 , n46784 , 
     n46785 , n224547 , n224548 , n46788 , n46789 , n46790 , n46791 , n46792 , n46793 , n224555 , 
     n224556 , n46796 , n46797 , n224559 , n224560 , n46800 , n46801 , n46802 , n46803 , n46804 , 
     n46805 , n46806 , n46807 , n224569 , n224570 , n46810 , n46811 , n46812 , n46813 , n46814 , 
     n46815 , n46816 , n46817 , n46818 , n46819 , n224581 , n224582 , n46822 , n46823 , n46824 , 
     n46825 , n46826 , n46827 , n46828 , n46829 , n46830 , n46831 , n46832 , n46833 , n224595 , 
     n224596 , n46836 , n46837 , n46838 , n46839 , n46840 , n46841 , n46842 , n46843 , n224605 , 
     n224606 , n46846 , n224608 , n224609 , n46849 , n46850 , n46851 , n46852 , n46853 , n46854 , 
     n46855 , n46856 , n46857 , n46858 , n224620 , n224621 , n46861 , n224623 , n224624 , n46864 , 
     n224626 , n224627 , n46867 , n46868 , n46869 , n46870 , n46871 , n46872 , n224634 , n224635 , 
     n46875 , n46876 , n46877 , n46878 , n46879 , n46880 , n224642 , n224643 , n46883 , n46884 , 
     n46885 , n46886 , n46887 , n46888 , n46889 , n46890 , n46891 , n46892 , n46893 , n46894 , 
     n224656 , n224657 , n46897 , n224659 , n224660 , n46900 , n46901 , n46902 , n46903 , n46904 , 
     n46905 , n224667 , n224668 , n46908 , n46909 , n46910 , n46911 , n224673 , n224674 , n46914 , 
     n46915 , n46916 , n46917 , n46918 , n46919 , n46920 , n46921 , n46922 , n46923 , n224685 , 
     n224686 , n46926 , n46927 , n46928 , n46929 , n224691 , n224692 , n46932 , n46933 , n46934 , 
     n46935 , n46936 , n46937 , n224699 , n224700 , n46940 , n46941 , n46942 , n46943 , n46944 , 
     n46945 , n224707 , n224708 , n46948 , n46949 , n46950 , n46951 , n46952 , n46953 , n224715 , 
     n224716 , n46956 , n46957 , n46958 , n46959 , n46960 , n46961 , n224723 , n224724 , n46964 , 
     n46965 , n46966 , n46967 , n46968 , n46969 , n46970 , n46971 , n46972 , n46973 , n224735 , 
     n224736 , n46976 , n46977 , n46978 , n46979 , n46980 , n46981 , n46982 , n46983 , n46984 , 
     n46985 , n224747 , n224748 , n46988 , n46989 , n46990 , n46991 , n46992 , n46993 , n46994 , 
     n46995 , n224757 , n224758 , n224759 , n224760 , n47000 , n224762 , n224763 , n47003 , n47004 , 
     n47005 , n47006 , n224768 , n224769 , n47009 , n47010 , n47011 , n47012 , n47013 , n47014 , 
     n224776 , n224777 , n47017 , n47018 , n47019 , n47020 , n47021 , n47022 , n47023 , n47024 , 
     n47025 , n47026 , n224788 , n224789 , n47029 , n47030 , n47031 , n47032 , n47033 , n47034 , 
     n47035 , n47036 , n47037 , n47038 , n224800 , n224801 , n47041 , n224803 , n224804 , n47044 , 
     n224806 , n224807 , n47047 , n47048 , n47049 , n47050 , n47051 , n47052 , n224814 , n224815 , 
     n47055 , n47056 , n47057 , n47058 , n224820 , n224821 , n47061 , n47062 , n47063 , n47064 , 
     n47065 , n47066 , n47067 , n47068 , n47069 , n47070 , n224832 , n224833 , n47073 , n47074 , 
     n47075 , n47076 , n47077 , n47078 , n224840 , n224841 , n47081 , n224843 , n224844 , n47084 , 
     n47085 , n47086 , n47087 , n47088 , n224850 , n224851 , n47091 , n224853 , n224854 , n47094 , 
     n224856 , n224857 , n224858 , n224859 , n47099 , n47100 , n47101 , n47102 , n47103 , n224865 , 
     n224866 , n47106 , n47107 , n47108 , n47109 , n47110 , n47111 , n47112 , n224874 , n224875 , 
     n47115 , n224877 , n224878 , n47118 , n47119 , n47120 , n47121 , n224883 , n224884 , n47124 , 
     n47125 , n47126 , n47127 , n47128 , n47129 , n47130 , n47131 , n224893 , n224894 , n47134 , 
     n47135 , n47136 , n47137 , n47138 , n47139 , n47140 , n47141 , n224903 , n224904 , n47144 , 
     n47145 , n47146 , n47147 , n47148 , n47149 , n224911 , n224912 , n47152 , n224914 , n224915 , 
     n47155 , n47156 , n47157 , n47158 , n47159 , n47160 , n47161 , n47162 , n224924 , n224925 , 
     n47165 , n47166 , n47167 , n47168 , n47169 , n47170 , n47171 , n47172 , n47173 , n47174 , 
     n47175 , n224937 , n224938 , n47178 , n47179 , n47180 , n47181 , n47182 , n47183 , n47184 , 
     n224946 , n224947 , n47187 , n224949 , n224950 , n47190 , n47191 , n47192 , n47193 , n47194 , 
     n47195 , n47196 , n47197 , n224959 , n224960 , n47200 , n47201 , n47202 , n47203 , n47204 , 
     n47205 , n224967 , n224968 , n47208 , n224970 , n224971 , n47211 , n47212 , n47213 , n47214 , 
     n47215 , n47216 , n47217 , n47218 , n224980 , n224981 , n224982 , n224983 , n47223 , n47224 , 
     n47225 , n47226 , n47227 , n47228 , n224990 , n224991 , n47231 , n224993 , n224994 , n47234 , 
     n47235 , n47236 , n47237 , n224999 , n225000 , n47240 , n225002 , n225003 , n47243 , n47244 , 
     n47245 , n47246 , n47247 , n47248 , n47249 , n47250 , n225012 , n225013 , n47253 , n47254 , 
     n47255 , n47256 , n47257 , n47258 , n225020 , n225021 , n47261 , n47262 , n47263 , n47264 , 
     n225026 , n225027 , n47267 , n47268 , n47269 , n47270 , n225032 , n225033 , n47273 , n47274 , 
     n47275 , n47276 , n225038 , n225039 , n47279 , n47280 , n47281 , n47282 , n225044 , n225045 , 
     n47285 , n47286 , n47287 , n47288 , n47289 , n47290 , n225052 , n225053 , n47293 , n47294 , 
     n47295 , n47296 , n47297 , n47298 , n225060 , n225061 , n47301 , n47302 , n47303 , n47304 , 
     n47305 , n47306 , n47307 , n47308 , n47309 , n47310 , n47311 , n47312 , n47313 , n225075 , 
     n225076 , n47316 , n47317 , n47318 , n47319 , n47320 , n47321 , n225083 , n225084 , n47324 , 
     n225086 , n225087 , n47327 , n225089 , n225090 , n47330 , n47331 , n47332 , n47333 , n47334 , 
     n47335 , n47336 , n47337 , n47338 , n47339 , n225101 , n225102 , n47342 , n225104 , n225105 , 
     n47345 , n47346 , n47347 , n225109 , n225110 , n225111 , n225112 , n47352 , n47353 , n47354 , 
     n47355 , n47356 , n47357 , n225119 , n225120 , n47360 , n47361 , n47362 , n47363 , n47364 , 
     n47365 , n225127 , n225128 , n47368 , n47369 , n47370 , n47371 , n47372 , n47373 , n47374 , 
     n47375 , n225137 , n225138 , n47378 , n47379 , n47380 , n47381 , n225143 , n225144 , n47384 , 
     n225146 , n225147 , n47387 , n47388 , n47389 , n47390 , n47391 , n47392 , n225154 , n225155 , 
     n47395 , n225157 , n225158 , n47398 , n47399 , n47400 , n47401 , n47402 , n47403 , n225165 , 
     n225166 , n47406 , n47407 , n47408 , n47409 , n47410 , n47411 , n47412 , n47413 , n225175 , 
     n225176 , n225177 , n225178 , n47418 , n47419 , n47420 , n47421 , n47422 , n47423 , n225185 , 
     n225186 , n47426 , n47427 , n47428 , n47429 , n47430 , n47431 , n47432 , n47433 , n47434 , 
     n47435 , n47436 , n47437 , n225199 , n225200 , n47440 , n47441 , n47442 , n47443 , n47444 , 
     n47445 , n47446 , n47447 , n225209 , n225210 , n47450 , n47451 , n47452 , n47453 , n47454 , 
     n47455 , n225217 , n225218 , n47458 , n47459 , n47460 , n47461 , n225223 , n225224 , n47464 , 
     n47465 , n47466 , n47467 , n225229 , n225230 , n47470 , n225232 , n225233 , n47473 , n47474 , 
     n47475 , n47476 , n47477 , n225239 , n225240 , n47480 , n47481 , n225243 , n225244 , n47484 , 
     n47485 , n47486 , n47487 , n47488 , n47489 , n225251 , n225252 , n47492 , n47493 , n47494 , 
     n47495 , n225257 , n225258 , n47498 , n47499 , n47500 , n47501 , n225263 , n225264 , n47504 , 
     n47505 , n47506 , n47507 , n225269 , n225270 , n47510 , n47511 , n47512 , n47513 , n47514 , 
     n47515 , n47516 , n47517 , n225279 , n225280 , n47520 , n225282 , n47522 , n225284 , n225285 , 
     n47525 , n47526 , n47527 , n47528 , n47529 , n47530 , n47531 , n47532 , n47533 , n47534 , 
     n47535 , n225297 , n225298 , n47538 , n47539 , n225301 , n225302 , n47542 , n47543 , n47544 , 
     n47545 , n47546 , n47547 , n225309 , n225310 , n47550 , n47551 , n47552 , n47553 , n47554 , 
     n47555 , n47556 , n47557 , n225319 , n225320 , n47560 , n47561 , n47562 , n47563 , n47564 , 
     n47565 , n47566 , n225328 , n225329 , n225330 , n225331 , n47571 , n47572 , n47573 , n47574 , 
     n47575 , n47576 , n47577 , n47578 , n225340 , n225341 , n47581 , n225343 , n225344 , n47584 , 
     n47585 , n47586 , n47587 , n47588 , n47589 , n225351 , n225352 , n47592 , n47593 , n47594 , 
     n47595 , n47596 , n47597 , n225359 , n225360 , n47600 , n47601 , n47602 , n47603 , n47604 , 
     n47605 , n47606 , n47607 , n47608 , n47609 , n225371 , n225372 , n47612 , n47613 , n47614 , 
     n47615 , n47616 , n47617 , n225379 , n225380 , n47620 , n225382 , n225383 , n47623 , n47624 , 
     n47625 , n47626 , n225388 , n225389 , n47629 , n47630 , n47631 , n47632 , n47633 , n47634 , 
     n47635 , n47636 , n47637 , n47638 , n47639 , n47640 , n47641 , n225403 , n225404 , n47644 , 
     n47645 , n47646 , n47647 , n47648 , n47649 , n47650 , n47651 , n225413 , n225414 , n47654 , 
     n47655 , n47656 , n47657 , n47658 , n47659 , n47660 , n47661 , n225423 , n225424 , n47664 , 
     n47665 , n47666 , n47667 , n225429 , n225430 , n47670 , n47671 , n47672 , n47673 , n225435 , 
     n225436 , n47676 , n225438 , n225439 , n47679 , n47680 , n47681 , n47682 , n47683 , n47684 , 
     n225446 , n225447 , n47687 , n47688 , n47689 , n225451 , n225452 , n47692 , n47693 , n47694 , 
     n47695 , n47696 , n47697 , n225459 , n225460 , n47700 , n47701 , n47702 , n47703 , n47704 , 
     n47705 , n225467 , n225468 , n47708 , n47709 , n47710 , n47711 , n225473 , n225474 , n47714 , 
     n47715 , n47716 , n47717 , n47718 , n47719 , n225481 , n225482 , n47722 , n47723 , n47724 , 
     n47725 , n225487 , n225488 , n47728 , n47729 , n47730 , n47731 , n47732 , n47733 , n225495 , 
     n225496 , n47736 , n47737 , n47738 , n47739 , n225501 , n225502 , n47742 , n47743 , n47744 , 
     n47745 , n47746 , n47747 , n225509 , n225510 , n47750 , n225512 , n47752 , n225514 , n225515 , 
     n47755 , n225517 , n225518 , n47758 , n47759 , n47760 , n47761 , n47762 , n47763 , n225525 , 
     n225526 , n47766 , n47767 , n47768 , n47769 , n47770 , n47771 , n47772 , n47773 , n225535 , 
     n225536 , n47776 , n47777 , n47778 , n47779 , n47780 , n47781 , n47782 , n47783 , n47784 , 
     n47785 , n225547 , n225548 , n47788 , n225550 , n225551 , n47791 , n47792 , n47793 , n47794 , 
     n47795 , n47796 , n47797 , n47798 , n225560 , n225561 , n47801 , n225563 , n225564 , n47804 , 
     n47805 , n47806 , n47807 , n47808 , n47809 , n47810 , n225572 , n225573 , n47813 , n47814 , 
     n47815 , n47816 , n47817 , n47818 , n225580 , n225581 , n47821 , n47822 , n47823 , n47824 , 
     n47825 , n47826 , n47827 , n47828 , n47829 , n47830 , n47831 , n225593 , n225594 , n47834 , 
     n225596 , n225597 , n47837 , n47838 , n47839 , n47840 , n47841 , n47842 , n225604 , n225605 , 
     n47845 , n225607 , n225608 , n47848 , n47849 , n47850 , n47851 , n47852 , n47853 , n47854 , 
     n47855 , n47856 , n47857 , n225619 , n225620 , n47860 , n225622 , n225623 , n47863 , n47864 , 
     n47865 , n47866 , n47867 , n47868 , n225630 , n225631 , n47871 , n47872 , n47873 , n47874 , 
     n47875 , n47876 , n225638 , n225639 , n47879 , n47880 , n47881 , n47882 , n225644 , n225645 , 
     n47885 , n47886 , n47887 , n47888 , n47889 , n47890 , n225652 , n225653 , n47893 , n47894 , 
     n225656 , n225657 , n47897 , n47898 , n47899 , n47900 , n47901 , n225663 , n225664 , n47904 , 
     n47905 , n47906 , n47907 , n47908 , n47909 , n47910 , n47911 , n225673 , n225674 , n47914 , 
     n225676 , n225677 , n47917 , n225679 , n225680 , n47920 , n225682 , n225683 , n47923 , n47924 , 
     n47925 , n47926 , n225688 , n225689 , n47929 , n225691 , n225692 , n47932 , n47933 , n225695 , 
     n225696 , n47936 , n47937 , n47938 , n47939 , n47940 , n47941 , n47942 , n47943 , n225705 , 
     n225706 , n47946 , n47947 , n47948 , n47949 , n47950 , n47951 , n225713 , n225714 , n47954 , 
     n225716 , n225717 , n47957 , n47958 , n47959 , n47960 , n47961 , n47962 , n47963 , n47964 , 
     n225726 , n225727 , n47967 , n47968 , n47969 , n47970 , n47971 , n47972 , n47973 , n47974 , 
     n225736 , n225737 , n225738 , n225739 , n47979 , n225741 , n225742 , n47982 , n47983 , n47984 , 
     n47985 , n47986 , n47987 , n47988 , n47989 , n47990 , n47991 , n225753 , n225754 , n47994 , 
     n225756 , n225757 , n47997 , n47998 , n47999 , n48000 , n225762 , n225763 , n48003 , n48004 , 
     n48005 , n48006 , n48007 , n48008 , n225770 , n225771 , n48011 , n48012 , n48013 , n48014 , 
     n48015 , n48016 , n225778 , n225779 , n48019 , n225781 , n225782 , n48022 , n48023 , n48024 , 
     n48025 , n48026 , n48027 , n48028 , n48029 , n48030 , n48031 , n225793 , n225794 , n48034 , 
     n225796 , n225797 , n48037 , n48038 , n48039 , n48040 , n48041 , n48042 , n225804 , n225805 , 
     n48045 , n48046 , n48047 , n48048 , n48049 , n48050 , n225812 , n225813 , n48053 , n48054 , 
     n48055 , n48056 , n48057 , n48058 , n225820 , n225821 , n48061 , n48062 , n48063 , n48064 , 
     n48065 , n225827 , n225828 , n225829 , n225830 , n48070 , n48071 , n48072 , n48073 , n225835 , 
     n225836 , n48076 , n48077 , n48078 , n48079 , n48080 , n225842 , n225843 , n48083 , n48084 , 
     n48085 , n48086 , n225848 , n225849 , n48089 , n48090 , n48091 , n48092 , n48093 , n48094 , 
     n48095 , n225857 , n225858 , n48098 , n48099 , n48100 , n48101 , n225863 , n225864 , n48104 , 
     n225866 , n225867 , n48107 , n225869 , n225870 , n48110 , n48111 , n48112 , n48113 , n48114 , 
     n48115 , n48116 , n48117 , n48118 , n48119 , n225881 , n225882 , n48122 , n48123 , n48124 , 
     n48125 , n225887 , n225888 , n48128 , n48129 , n48130 , n48131 , n48132 , n48133 , n225895 , 
     n225896 , n48136 , n48137 , n48138 , n48139 , n225901 , n225902 , n48142 , n48143 , n48144 , 
     n48145 , n225907 , n225908 , n48148 , n48149 , n48150 , n48151 , n225913 , n225914 , n48154 , 
     n48155 , n48156 , n48157 , n225919 , n225920 , n48160 , n48161 , n48162 , n48163 , n225925 , 
     n225926 , n48166 , n48167 , n48168 , n48169 , n48170 , n48171 , n48172 , n48173 , n48174 , 
     n48175 , n225937 , n225938 , n48178 , n48179 , n48180 , n48181 , n48182 , n48183 , n48184 , 
     n48185 , n225947 , n225948 , n48188 , n48189 , n48190 , n48191 , n225953 , n225954 , n48194 , 
     n225956 , n225957 , n48197 , n48198 , n48199 , n48200 , n48201 , n48202 , n48203 , n225965 , 
     n225966 , n48206 , n48207 , n48208 , n48209 , n48210 , n48211 , n48212 , n225974 , n225975 , 
     n48215 , n48216 , n48217 , n48218 , n225980 , n225981 , n48221 , n48222 , n48223 , n48224 , 
     n225986 , n225987 , n48227 , n225989 , n225990 , n48230 , n48231 , n48232 , n48233 , n48234 , 
     n48235 , n225997 , n225998 , n48238 , n226000 , n226001 , n48241 , n226003 , n226004 , n48244 , 
     n48245 , n48246 , n48247 , n48248 , n226010 , n226011 , n48251 , n48252 , n48253 , n48254 , 
     n48255 , n48256 , n48257 , n226019 , n226020 , n48260 , n48261 , n48262 , n48263 , n48264 , 
     n48265 , n48266 , n48267 , n48268 , n48269 , n226031 , n226032 , n48272 , n226034 , n226035 , 
     n48275 , n226037 , n226038 , n48278 , n226040 , n226041 , n48281 , n48282 , n48283 , n48284 , 
     n48285 , n48286 , n48287 , n48288 , n48289 , n48290 , n48291 , n226053 , n226054 , n48294 , 
     n48295 , n48296 , n48297 , n48298 , n48299 , n226061 , n226062 , n48302 , n48303 , n48304 , 
     n48305 , n48306 , n48307 , n48308 , n48309 , n48310 , n48311 , n48312 , n226074 , n226075 , 
     n48315 , n48316 , n48317 , n48318 , n48319 , n48320 , n48321 , n48322 , n226084 , n226085 , 
     n48325 , n226087 , n226088 , n48328 , n48329 , n48330 , n48331 , n226093 , n226094 , n48334 , 
     n226096 , n226097 , n48337 , n226099 , n226100 , n48340 , n48341 , n48342 , n48343 , n48344 , 
     n48345 , n48346 , n48347 , n226109 , n226110 , n48350 , n48351 , n48352 , n48353 , n48354 , 
     n48355 , n226117 , n226118 , n48358 , n48359 , n48360 , n48361 , n226123 , n226124 , n48364 , 
     n226126 , n226127 , n48367 , n48368 , n48369 , n48370 , n226132 , n226133 , n48373 , n48374 , 
     n48375 , n48376 , n48377 , n48378 , n48379 , n48380 , n48381 , n48382 , n226144 , n226145 , 
     n48385 , n226147 , n226148 , n48388 , n48389 , n48390 , n48391 , n48392 , n48393 , n226155 , 
     n226156 , n48396 , n48397 , n48398 , n48399 , n48400 , n48401 , n226163 , n226164 , n48404 , 
     n48405 , n48406 , n48407 , n226169 , n226170 , n48410 , n48411 , n48412 , n48413 , n48414 , 
     n48415 , n226177 , n226178 , n48418 , n48419 , n48420 , n48421 , n226183 , n226184 , n48424 , 
     n226186 , n226187 , n48427 , n48428 , n48429 , n48430 , n48431 , n48432 , n226194 , n226195 , 
     n48435 , n48436 , n48437 , n48438 , n226200 , n226201 , n48441 , n226203 , n226204 , n48444 , 
     n48445 , n48446 , n48447 , n48448 , n48449 , n48450 , n48451 , n48452 , n48453 , n226215 , 
     n226216 , n48456 , n226218 , n226219 , n48459 , n48460 , n48461 , n48462 , n226224 , n226225 , 
     n48465 , n48466 , n48467 , n48468 , n48469 , n48470 , n226232 , n226233 , n48473 , n226235 , 
     n226236 , n48476 , n226238 , n226239 , n48479 , n48480 , n48481 , n48482 , n48483 , n48484 , 
     n226246 , n226247 , n48487 , n48488 , n48489 , n48490 , n48491 , n48492 , n226254 , n226255 , 
     n48495 , n48496 , n48497 , n226259 , n226260 , n226261 , n226262 , n48502 , n48503 , n48504 , 
     n48505 , n48506 , n48507 , n226269 , n226270 , n48510 , n48511 , n48512 , n48513 , n226275 , 
     n226276 , n48516 , n226278 , n226279 , n48519 , n48520 , n48521 , n48522 , n226284 , n226285 , 
     n48525 , n48526 , n48527 , n48528 , n48529 , n48530 , n226292 , n226293 , n48533 , n48534 , 
     n48535 , n48536 , n48537 , n48538 , n226300 , n226301 , n48541 , n226303 , n226304 , n48544 , 
     n48545 , n48546 , n48547 , n48548 , n48549 , n48550 , n48551 , n226313 , n226314 , n48554 , 
     n48555 , n48556 , n48557 , n226319 , n226320 , n226321 , n226322 , n48562 , n48563 , n48564 , 
     n48565 , n226327 , n226328 , n48568 , n48569 , n48570 , n48571 , n226333 , n226334 , n48574 , 
     n48575 , n48576 , n48577 , n226339 , n226340 , n48580 , n48581 , n48582 , n48583 , n48584 , 
     n48585 , n48586 , n48587 , n226349 , n226350 , n48590 , n48591 , n48592 , n48593 , n48594 , 
     n48595 , n226357 , n226358 , n48598 , n226360 , n226361 , n48601 , n226363 , n226364 , n48604 , 
     n48605 , n48606 , n48607 , n226369 , n226370 , n48610 , n48611 , n48612 , n48613 , n48614 , 
     n48615 , n226377 , n226378 , n48618 , n48619 , n48620 , n48621 , n226383 , n226384 , n48624 , 
     n226386 , n48626 , n48627 , n48628 , n48629 , n48630 , n48631 , n48632 , n48633 , n48634 , 
     n48635 , n226397 , n226398 , n48638 , n48639 , n48640 , n48641 , n48642 , n48643 , n48644 , 
     n48645 , n226407 , n226408 , n48648 , n48649 , n226411 , n48651 , n48652 , n48653 , n48654 , 
     n226416 , n226417 , n48657 , n48658 , n48659 , n48660 , n48661 , n48662 , n226424 , n226425 , 
     n48665 , n48666 , n48667 , n48668 , n226430 , n226431 , n48671 , n226433 , n226434 , n48674 , 
     n48675 , n48676 , n48677 , n226439 , n226440 , n48680 , n226442 , n226443 , n48683 , n48684 , 
     n48685 , n48686 , n48687 , n48688 , n48689 , n48690 , n48691 , n48692 , n226454 , n226455 , 
     n48695 , n48696 , n48697 , n48698 , n226460 , n226461 , n48701 , n226463 , n226464 , n48704 , 
     n226466 , n226467 , n48707 , n48708 , n48709 , n48710 , n226472 , n226473 , n48713 , n226475 , 
     n226476 , n48716 , n48717 , n48718 , n48719 , n48720 , n48721 , n226483 , n226484 , n48724 , 
     n48725 , n48726 , n48727 , n226489 , n226490 , n48730 , n48731 , n48732 , n48733 , n48734 , 
     n48735 , n48736 , n48737 , n48738 , n48739 , n226501 , n226502 , n48742 , n48743 , n48744 , 
     n48745 , n48746 , n48747 , n48748 , n48749 , n48750 , n226512 , n226513 , n48753 , n48754 , 
     n48755 , n48756 , n48757 , n48758 , n48759 , n226521 , n226522 , n48762 , n226524 , n226525 , 
     n48765 , n226527 , n226528 , n48768 , n48769 , n48770 , n48771 , n48772 , n48773 , n226535 , 
     n226536 , n48776 , n48777 , n48778 , n48779 , n48780 , n48781 , n226543 , n226544 , n48784 , 
     n48785 , n48786 , n48787 , n48788 , n226550 , n226551 , n48791 , n48792 , n48793 , n48794 , 
     n226556 , n226557 , n48797 , n48798 , n48799 , n48800 , n48801 , n48802 , n48803 , n48804 , 
     n48805 , n48806 , n226568 , n226569 , n48809 , n48810 , n48811 , n48812 , n226574 , n226575 , 
     n48815 , n48816 , n48817 , n48818 , n48819 , n48820 , n226582 , n226583 , n48823 , n226585 , 
     n226586 , n48826 , n48827 , n48828 , n48829 , n48830 , n48831 , n48832 , n48833 , n226595 , 
     n226596 , n48836 , n48837 , n48838 , n48839 , n48840 , n48841 , n226603 , n226604 , n48844 , 
     n226606 , n226607 , n48847 , n226609 , n226610 , n48850 , n226612 , n226613 , n48853 , n226615 , 
     n226616 , n48856 , n226618 , n226619 , n48859 , n48860 , n48861 , n48862 , n226624 , n226625 , 
     n48865 , n48866 , n48867 , n48868 , n48869 , n48870 , n226632 , n226633 , n48873 , n48874 , 
     n48875 , n48876 , n48877 , n48878 , n226640 , n226641 , n48881 , n48882 , n48883 , n48884 , 
     n48885 , n48886 , n226648 , n226649 , n48889 , n48890 , n48891 , n48892 , n48893 , n48894 , 
     n48895 , n48896 , n48897 , n226659 , n226660 , n48900 , n48901 , n48902 , n48903 , n48904 , 
     n48905 , n226667 , n226668 , n48908 , n48909 , n48910 , n48911 , n48912 , n48913 , n48914 , 
     n48915 , n48916 , n48917 , n48918 , n226680 , n226681 , n48921 , n48922 , n48923 , n48924 , 
     n226686 , n226687 , n48927 , n226689 , n226690 , n48930 , n48931 , n48932 , n48933 , n48934 , 
     n48935 , n48936 , n48937 , n48938 , n48939 , n226701 , n226702 , n48942 , n48943 , n48944 , 
     n48945 , n226707 , n226708 , n48948 , n48949 , n48950 , n48951 , n48952 , n48953 , n48954 , 
     n48955 , n48956 , n48957 , n226719 , n226720 , n48960 , n48961 , n48962 , n48963 , n48964 , 
     n48965 , n48966 , n48967 , n226729 , n226730 , n48970 , n48971 , n48972 , n48973 , n48974 , 
     n48975 , n48976 , n48977 , n48978 , n48979 , n226741 , n226742 , n48982 , n48983 , n48984 , 
     n48985 , n48986 , n48987 , n48988 , n226750 , n226751 , n48991 , n48992 , n48993 , n48994 , 
     n226756 , n226757 , n48997 , n48998 , n48999 , n49000 , n226762 , n226763 , n49003 , n226765 , 
     n226766 , n49006 , n226768 , n226769 , n49009 , n226771 , n226772 , n49012 , n49013 , n49014 , 
     n49015 , n226777 , n226778 , n49018 , n49019 , n49020 , n49021 , n49022 , n49023 , n226785 , 
     n226786 , n49026 , n49027 , n49028 , n49029 , n49030 , n49031 , n226793 , n226794 , n49034 , 
     n49035 , n49036 , n49037 , n49038 , n49039 , n226801 , n226802 , n49042 , n49043 , n49044 , 
     n49045 , n226807 , n226808 , n49048 , n226810 , n226811 , n49051 , n49052 , n49053 , n49054 , 
     n49055 , n49056 , n226818 , n226819 , n49059 , n226821 , n226822 , n49062 , n49063 , n49064 , 
     n49065 , n49066 , n49067 , n49068 , n49069 , n49070 , n49071 , n49072 , n226834 , n226835 , 
     n49075 , n49076 , n49077 , n49078 , n49079 , n49080 , n49081 , n49082 , n49083 , n226845 , 
     n226846 , n49086 , n226848 , n226849 , n49089 , n226851 , n226852 , n49092 , n49093 , n49094 , 
     n49095 , n49096 , n49097 , n226859 , n226860 , n49100 , n49101 , n49102 , n49103 , n226865 , 
     n226866 , n49106 , n226868 , n226869 , n49109 , n226871 , n226872 , n49112 , n226874 , n226875 , 
     n49115 , n226877 , n226878 , n49118 , n49119 , n49120 , n49121 , n49122 , n49123 , n226885 , 
     n226886 , n49126 , n49127 , n49128 , n49129 , n226891 , n226892 , n49132 , n49133 , n49134 , 
     n49135 , n49136 , n49137 , n226899 , n226900 , n49140 , n226902 , n226903 , n49143 , n49144 , 
     n49145 , n49146 , n49147 , n49148 , n49149 , n49150 , n49151 , n49152 , n226914 , n226915 , 
     n49155 , n49156 , n226918 , n226919 , n49159 , n49160 , n49161 , n49162 , n49163 , n226925 , 
     n226926 , n226927 , n226928 , n49168 , n49169 , n49170 , n49171 , n226933 , n226934 , n49174 , 
     n226936 , n226937 , n49177 , n49178 , n49179 , n49180 , n49181 , n49182 , n49183 , n49184 , 
     n49185 , n226947 , n226948 , n49188 , n49189 , n49190 , n49191 , n49192 , n49193 , n226955 , 
     n226956 , n49196 , n226958 , n226959 , n49199 , n49200 , n49201 , n49202 , n49203 , n49204 , 
     n226966 , n226967 , n49207 , n49208 , n49209 , n49210 , n49211 , n49212 , n226974 , n226975 , 
     n49215 , n49216 , n49217 , n49218 , n49219 , n49220 , n226982 , n226983 , n49223 , n226985 , 
     n226986 , n49226 , n49227 , n49228 , n49229 , n226991 , n226992 , n49232 , n49233 , n49234 , 
     n49235 , n49236 , n49237 , n49238 , n49239 , n227001 , n227002 , n49242 , n227004 , n227005 , 
     n49245 , n227007 , n227008 , n49248 , n49249 , n227011 , n227012 , n49252 , n49253 , n49254 , 
     n49255 , n49256 , n227018 , n227019 , n49259 , n49260 , n49261 , n49262 , n227024 , n227025 , 
     n49265 , n49266 , n49267 , n49268 , n227030 , n227031 , n49271 , n49272 , n49273 , n49274 , 
     n49275 , n49276 , n227038 , n227039 , n49279 , n49280 , n49281 , n49282 , n227044 , n227045 , 
     n49285 , n49286 , n49287 , n227049 , n227050 , n49290 , n49291 , n49292 , n49293 , n49294 , 
     n49295 , n49296 , n49297 , n49298 , n49299 , n227061 , n227062 , n49302 , n49303 , n49304 , 
     n49305 , n49306 , n49307 , n49308 , n227070 , n227071 , n227072 , n227073 , n49313 , n227075 , 
     n227076 , n49316 , n49317 , n49318 , n49319 , n227081 , n227082 , n49322 , n49323 , n49324 , 
     n49325 , n227087 , n227088 , n49328 , n227090 , n227091 , n49331 , n49332 , n49333 , n49334 , 
     n227096 , n227097 , n49337 , n49338 , n49339 , n49340 , n49341 , n49342 , n49343 , n49344 , 
     n49345 , n49346 , n49347 , n49348 , n49349 , n227111 , n227112 , n49352 , n49353 , n49354 , 
     n49355 , n49356 , n227118 , n227119 , n49359 , n49360 , n49361 , n49362 , n49363 , n49364 , 
     n49365 , n49366 , n49367 , n227129 , n227130 , n49370 , n49371 , n49372 , n227134 , n227135 , 
     n49375 , n49376 , n49377 , n49378 , n49379 , n49380 , n227142 , n227143 , n49383 , n227145 , 
     n227146 , n49386 , n49387 , n49388 , n49389 , n227151 , n227152 , n49392 , n49393 , n49394 , 
     n49395 , n49396 , n49397 , n227159 , n227160 , n49400 , n227162 , n227163 , n49403 , n227165 , 
     n227166 , n49406 , n49407 , n49408 , n49409 , n49410 , n49411 , n227173 , n227174 , n49414 , 
     n49415 , n49416 , n49417 , n227179 , n227180 , n49420 , n49421 , n49422 , n49423 , n49424 , 
     n49425 , n49426 , n49427 , n49428 , n49429 , n227191 , n227192 , n49432 , n49433 , n49434 , 
     n49435 , n227197 , n227198 , n49438 , n49439 , n49440 , n49441 , n227203 , n227204 , n49444 , 
     n49445 , n49446 , n49447 , n49448 , n49449 , n227211 , n227212 , n49452 , n49453 , n49454 , 
     n49455 , n49456 , n49457 , n49458 , n49459 , n227221 , n227222 , n49462 , n49463 , n49464 , 
     n49465 , n49466 , n49467 , n227229 , n227230 , n49470 , n49471 , n49472 , n49473 , n49474 , 
     n49475 , n227237 , n227238 , n49478 , n227240 , n227241 , n49481 , n49482 , n49483 , n49484 , 
     n227246 , n227247 , n49487 , n227249 , n227250 , n49490 , n49491 , n49492 , n49493 , n49494 , 
     n49495 , n49496 , n49497 , n49498 , n49499 , n227261 , n227262 , n49502 , n49503 , n49504 , 
     n49505 , n49506 , n49507 , n227269 , n227270 , n49510 , n49511 , n49512 , n49513 , n49514 , 
     n49515 , n49516 , n49517 , n49518 , n49519 , n227281 , n227282 , n49522 , n49523 , n49524 , 
     n49525 , n49526 , n49527 , n49528 , n49529 , n227291 , n227292 , n49532 , n49533 , n49534 , 
     n49535 , n227297 , n227298 , n49538 , n227300 , n227301 , n49541 , n227303 , n227304 , n49544 , 
     n227306 , n227307 , n49547 , n49548 , n49549 , n49550 , n49551 , n49552 , n49553 , n49554 , 
     n49555 , n49556 , n227318 , n227319 , n49559 , n49560 , n49561 , n49562 , n49563 , n49564 , 
     n49565 , n49566 , n49567 , n49568 , n227330 , n227331 , n49571 , n49572 , n49573 , n49574 , 
     n49575 , n49576 , n49577 , n49578 , n49579 , n49580 , n227342 , n227343 , n49583 , n49584 , 
     n49585 , n49586 , n49587 , n49588 , n49589 , n49590 , n227352 , n227353 , n49593 , n49594 , 
     n49595 , n49596 , n49597 , n49598 , n227360 , n227361 , n49601 , n49602 , n49603 , n49604 , 
     n49605 , n49606 , n227368 , n227369 , n49609 , n227371 , n227372 , n49612 , n49613 , n227375 , 
     n227376 , n49616 , n49617 , n49618 , n49619 , n227381 , n227382 , n49622 , n227384 , n227385 , 
     n49625 , n49626 , n49627 , n49628 , n49629 , n49630 , n49631 , n49632 , n227394 , n227395 , 
     n49635 , n49636 , n49637 , n49638 , n49639 , n49640 , n49641 , n49642 , n227404 , n227405 , 
     n49645 , n49646 , n49647 , n49648 , n227410 , n227411 , n49651 , n49652 , n49653 , n49654 , 
     n227416 , n227417 , n49657 , n49658 , n49659 , n49660 , n227422 , n227423 , n49663 , n49664 , 
     n49665 , n49666 , n49667 , n49668 , n227430 , n227431 , n49671 , n49672 , n49673 , n49674 , 
     n227436 , n227437 , n49677 , n227439 , n227440 , n49680 , n49681 , n49682 , n227444 , n227445 , 
     n227446 , n227447 , n49687 , n49688 , n49689 , n49690 , n227452 , n227453 , n49693 , n49694 , 
     n49695 , n49696 , n49697 , n49698 , n227460 , n227461 , n49701 , n49702 , n49703 , n49704 , 
     n49705 , n49706 , n49707 , n49708 , n49709 , n49710 , n227472 , n227473 , n49713 , n49714 , 
     n49715 , n49716 , n49717 , n49718 , n227480 , n227481 , n49721 , n227483 , n227484 , n49724 , 
     n49725 , n49726 , n49727 , n227489 , n227490 , n49730 , n49731 , n49732 , n49733 , n227495 , 
     n227496 , n227497 , n227498 , n49738 , n49739 , n49740 , n49741 , n227503 , n227504 , n49744 , 
     n227506 , n227507 , n49747 , n49748 , n49749 , n49750 , n49751 , n49752 , n227514 , n227515 , 
     n49755 , n49756 , n49757 , n49758 , n227520 , n227521 , n49761 , n227523 , n227524 , n49764 , 
     n49765 , n49766 , n227528 , n49768 , n49769 , n49770 , n49771 , n49772 , n49773 , n49774 , 
     n49775 , n227537 , n227538 , n49778 , n227540 , n227541 , n49781 , n49782 , n49783 , n49784 , 
     n49785 , n49786 , n227548 , n227549 , n49789 , n49790 , n49791 , n49792 , n49793 , n49794 , 
     n227556 , n227557 , n49797 , n227559 , n227560 , n49800 , n49801 , n49802 , n49803 , n49804 , 
     n49805 , n227567 , n227568 , n49808 , n49809 , n49810 , n49811 , n227573 , n227574 , n49814 , 
     n227576 , n227577 , n49817 , n49818 , n49819 , n49820 , n49821 , n49822 , n49823 , n49824 , 
     n227586 , n227587 , n49827 , n227589 , n227590 , n49830 , n49831 , n49832 , n49833 , n227595 , 
     n227596 , n49836 , n227598 , n227599 , n49839 , n49840 , n49841 , n49842 , n227604 , n227605 , 
     n49845 , n227607 , n227608 , n49848 , n227610 , n227611 , n49851 , n49852 , n49853 , n49854 , 
     n49855 , n49856 , n227618 , n227619 , n49859 , n49860 , n49861 , n49862 , n227624 , n227625 , 
     n49865 , n49866 , n49867 , n49868 , n49869 , n227631 , n227632 , n49872 , n49873 , n49874 , 
     n49875 , n49876 , n49877 , n227639 , n227640 , n49880 , n49881 , n49882 , n49883 , n49884 , 
     n49885 , n227647 , n227648 , n49888 , n49889 , n49890 , n49891 , n49892 , n49893 , n227655 , 
     n227656 , n49896 , n49897 , n49898 , n49899 , n49900 , n49901 , n49902 , n49903 , n227665 , 
     n227666 , n49906 , n49907 , n49908 , n49909 , n49910 , n49911 , n227673 , n227674 , n49914 , 
     n49915 , n49916 , n49917 , n49918 , n49919 , n227681 , n227682 , n49922 , n227684 , n227685 , 
     n49925 , n227687 , n227688 , n49928 , n49929 , n49930 , n49931 , n227693 , n227694 , n49934 , 
     n49935 , n49936 , n227698 , n227699 , n49939 , n49940 , n49941 , n49942 , n49943 , n49944 , 
     n227706 , n227707 , n49947 , n49948 , n49949 , n49950 , n227712 , n227713 , n49953 , n49954 , 
     n49955 , n49956 , n227718 , n227719 , n49959 , n49960 , n49961 , n49962 , n49963 , n49964 , 
     n49965 , n49966 , n49967 , n49968 , n227730 , n227731 , n49971 , n49972 , n49973 , n49974 , 
     n49975 , n49976 , n227738 , n227739 , n49979 , n49980 , n49981 , n49982 , n227744 , n227745 , 
     n49985 , n49986 , n49987 , n49988 , n227750 , n227751 , n49991 , n49992 , n49993 , n49994 , 
     n227756 , n227757 , n49997 , n49998 , n49999 , n50000 , n227762 , n227763 , n50003 , n50004 , 
     n50005 , n50006 , n50007 , n50008 , n50009 , n50010 , n227772 , n227773 , n50013 , n227775 , 
     n227776 , n50016 , n50017 , n50018 , n50019 , n50020 , n50021 , n50022 , n50023 , n227785 , 
     n227786 , n50026 , n50027 , n50028 , n50029 , n50030 , n50031 , n50032 , n50033 , n227795 , 
     n227796 , n50036 , n50037 , n50038 , n50039 , n227801 , n227802 , n50042 , n50043 , n50044 , 
     n50045 , n50046 , n50047 , n227809 , n227810 , n50050 , n50051 , n50052 , n50053 , n50054 , 
     n50055 , n50056 , n50057 , n50058 , n50059 , n227821 , n227822 , n50062 , n50063 , n50064 , 
     n50065 , n50066 , n50067 , n227829 , n227830 , n50070 , n50071 , n50072 , n50073 , n50074 , 
     n50075 , n227837 , n227838 , n50078 , n50079 , n50080 , n50081 , n50082 , n50083 , n227845 , 
     n227846 , n50086 , n227848 , n227849 , n50089 , n227851 , n50091 , n50092 , n50093 , n50094 , 
     n227856 , n227857 , n50097 , n50098 , n50099 , n50100 , n227862 , n227863 , n50103 , n50104 , 
     n50105 , n50106 , n227868 , n227869 , n50109 , n50110 , n50111 , n50112 , n227874 , n227875 , 
     n50115 , n50116 , n50117 , n50118 , n227880 , n227881 , n50121 , n50122 , n50123 , n50124 , 
     n50125 , n50126 , n50127 , n50128 , n50129 , n50130 , n227892 , n227893 , n50133 , n50134 , 
     n50135 , n50136 , n50137 , n50138 , n50139 , n50140 , n227902 , n227903 , n50143 , n50144 , 
     n50145 , n50146 , n50147 , n50148 , n50149 , n227911 , n227912 , n50152 , n50153 , n50154 , 
     n50155 , n227917 , n227918 , n50158 , n227920 , n227921 , n50161 , n50162 , n50163 , n50164 , 
     n50165 , n50166 , n227928 , n227929 , n50169 , n50170 , n50171 , n50172 , n50173 , n50174 , 
     n227936 , n227937 , n50177 , n50178 , n50179 , n50180 , n50181 , n50182 , n227944 , n227945 , 
     n50185 , n50186 , n50187 , n50188 , n50189 , n50190 , n50191 , n50192 , n227954 , n227955 , 
     n50195 , n50196 , n50197 , n50198 , n227960 , n227961 , n50201 , n50202 , n50203 , n50204 , 
     n227966 , n227967 , n50207 , n50208 , n50209 , n50210 , n227972 , n227973 , n50213 , n50214 , 
     n50215 , n50216 , n50217 , n50218 , n227980 , n227981 , n50221 , n50222 , n50223 , n50224 , 
     n227986 , n227987 , n50227 , n50228 , n50229 , n50230 , n50231 , n50232 , n50233 , n50234 , 
     n227996 , n227997 , n50237 , n50238 , n50239 , n50240 , n50241 , n50242 , n228004 , n228005 , 
     n50245 , n228007 , n228008 , n50248 , n50249 , n50250 , n50251 , n50252 , n50253 , n228015 , 
     n228016 , n50256 , n50257 , n50258 , n50259 , n50260 , n50261 , n228023 , n228024 , n50264 , 
     n50265 , n228027 , n228028 , n50268 , n50269 , n50270 , n50271 , n228033 , n228034 , n50274 , 
     n50275 , n50276 , n50277 , n50278 , n50279 , n228041 , n228042 , n50282 , n50283 , n50284 , 
     n50285 , n228047 , n228048 , n50288 , n50289 , n50290 , n50291 , n228053 , n228054 , n50294 , 
     n50295 , n50296 , n50297 , n50298 , n50299 , n228061 , n228062 , n50302 , n50303 , n50304 , 
     n50305 , n50306 , n50307 , n228069 , n228070 , n50310 , n228072 , n228073 , n50313 , n50314 , 
     n50315 , n50316 , n228078 , n228079 , n50319 , n50320 , n50321 , n50322 , n228084 , n228085 , 
     n50325 , n50326 , n50327 , n50328 , n228090 , n228091 , n50331 , n228093 , n228094 , n50334 , 
     n50335 , n50336 , n50337 , n228099 , n228100 , n50340 , n50341 , n50342 , n50343 , n228105 , 
     n228106 , n50346 , n50347 , n50348 , n50349 , n228111 , n228112 , n50352 , n50353 , n50354 , 
     n50355 , n50356 , n50357 , n50358 , n228120 , n228121 , n50361 , n50362 , n50363 , n50364 , 
     n50365 , n50366 , n50367 , n228129 , n228130 , n50370 , n228132 , n228133 , n50373 , n50374 , 
     n50375 , n50376 , n228138 , n228139 , n50379 , n50380 , n50381 , n50382 , n228144 , n228145 , 
     n50385 , n50386 , n50387 , n50388 , n228150 , n228151 , n50391 , n50392 , n50393 , n50394 , 
     n228156 , n228157 , n50397 , n50398 , n50399 , n50400 , n50401 , n50402 , n50403 , n50404 , 
     n50405 , n50406 , n50407 , n228169 , n228170 , n50410 , n50411 , n50412 , n50413 , n228175 , 
     n228176 , n50416 , n50417 , n50418 , n50419 , n50420 , n228182 , n228183 , n50423 , n50424 , 
     n50425 , n50426 , n50427 , n50428 , n50429 , n50430 , n50431 , n50432 , n228194 , n228195 , 
     n50435 , n50436 , n50437 , n50438 , n228200 , n228201 , n50441 , n50442 , n50443 , n50444 , 
     n50445 , n50446 , n228208 , n228209 , n50449 , n228211 , n228212 , n50452 , n50453 , n50454 , 
     n50455 , n50456 , n50457 , n50458 , n50459 , n228221 , n228222 , n50462 , n50463 , n50464 , 
     n50465 , n50466 , n50467 , n50468 , n50469 , n228231 , n228232 , n50472 , n50473 , n50474 , 
     n50475 , n228237 , n228238 , n50478 , n50479 , n50480 , n50481 , n50482 , n50483 , n50484 , 
     n50485 , n50486 , n50487 , n228249 , n228250 , n50490 , n50491 , n50492 , n50493 , n228255 , 
     n228256 , n50496 , n228258 , n228259 , n50499 , n228261 , n228262 , n50502 , n228264 , n228265 , 
     n50505 , n50506 , n50507 , n50508 , n228270 , n228271 , n50511 , n50512 , n50513 , n50514 , 
     n228276 , n228277 , n50517 , n50518 , n228280 , n228281 , n50521 , n50522 , n50523 , n50524 , 
     n50525 , n228287 , n228288 , n50528 , n50529 , n50530 , n50531 , n50532 , n50533 , n50534 , 
     n50535 , n228297 , n228298 , n50538 , n50539 , n50540 , n50541 , n50542 , n50543 , n228305 , 
     n228306 , n50546 , n50547 , n50548 , n50549 , n228311 , n228312 , n50552 , n50553 , n50554 , 
     n50555 , n228317 , n228318 , n50558 , n50559 , n50560 , n50561 , n50562 , n50563 , n228325 , 
     n228326 , n50566 , n50567 , n50568 , n50569 , n228331 , n228332 , n50572 , n228334 , n228335 , 
     n50575 , n50576 , n50577 , n50578 , n50579 , n50580 , n50581 , n50582 , n50583 , n228345 , 
     n228346 , n50586 , n50587 , n50588 , n50589 , n228351 , n228352 , n50592 , n50593 , n50594 , 
     n50595 , n228357 , n228358 , n50598 , n50599 , n50600 , n50601 , n228363 , n228364 , n50604 , 
     n228366 , n228367 , n50607 , n50608 , n50609 , n50610 , n228372 , n228373 , n50613 , n50614 , 
     n50615 , n228377 , n228378 , n228379 , n228380 , n50620 , n228382 , n228383 , n50623 , n228385 , 
     n228386 , n50626 , n50627 , n50628 , n50629 , n228391 , n228392 , n50632 , n50633 , n50634 , 
     n50635 , n228397 , n228398 , n50638 , n50639 , n50640 , n50641 , n228403 , n228404 , n50644 , 
     n50645 , n50646 , n50647 , n50648 , n50649 , n50650 , n228412 , n228413 , n50653 , n50654 , 
     n50655 , n50656 , n50657 , n50658 , n228420 , n228421 , n50661 , n50662 , n50663 , n50664 , 
     n50665 , n228427 , n228428 , n50668 , n50669 , n50670 , n50671 , n228433 , n228434 , n50674 , 
     n50675 , n50676 , n50677 , n228439 , n228440 , n50680 , n50681 , n50682 , n50683 , n228445 , 
     n228446 , n50686 , n50687 , n50688 , n50689 , n50690 , n50691 , n50692 , n50693 , n50694 , 
     n228456 , n228457 , n50697 , n228459 , n228460 , n50700 , n50701 , n50702 , n50703 , n228465 , 
     n228466 , n50706 , n50707 , n228469 , n228470 , n228471 , n228472 , n50712 , n50713 , n50714 , 
     n50715 , n50716 , n50717 , n228479 , n228480 , n50720 , n50721 , n50722 , n50723 , n228485 , 
     n228486 , n50726 , n50727 , n50728 , n50729 , n50730 , n50731 , n228493 , n228494 , n50734 , 
     n50735 , n50736 , n50737 , n228499 , n228500 , n50740 , n50741 , n50742 , n50743 , n50744 , 
     n50745 , n228507 , n228508 , n50748 , n50749 , n50750 , n50751 , n228513 , n228514 , n50754 , 
     n50755 , n50756 , n50757 , n50758 , n50759 , n228521 , n228522 , n50762 , n50763 , n50764 , 
     n228526 , n228527 , n50767 , n50768 , n50769 , n50770 , n228532 , n228533 , n50773 , n50774 , 
     n50775 , n50776 , n228538 , n228539 , n50779 , n50780 , n50781 , n50782 , n50783 , n50784 , 
     n228546 , n228547 , n50787 , n50788 , n50789 , n50790 , n50791 , n50792 , n228554 , n228555 , 
     n50795 , n50796 , n50797 , n50798 , n228560 , n228561 , n50801 , n50802 , n50803 , n50804 , 
     n228566 , n228567 , n50807 , n228569 , n228570 , n50810 , n50811 , n50812 , n50813 , n50814 , 
     n50815 , n228577 , n228578 , n50818 , n50819 , n50820 , n50821 , n50822 , n50823 , n50824 , 
     n50825 , n228587 , n228588 , n50828 , n50829 , n50830 , n228592 , n228593 , n50833 , n50834 , 
     n50835 , n50836 , n50837 , n50838 , n50839 , n50840 , n228602 , n228603 , n50843 , n50844 , 
     n228606 , n228607 , n50847 , n50848 , n50849 , n228611 , n228612 , n50852 , n50853 , n50854 , 
     n50855 , n50856 , n50857 , n228619 , n228620 , n50860 , n50861 , n50862 , n50863 , n228625 , 
     n228626 , n50866 , n50867 , n50868 , n50869 , n228631 , n228632 , n50872 , n50873 , n50874 , 
     n50875 , n228637 , n228638 , n50878 , n50879 , n50880 , n50881 , n228643 , n228644 , n50884 , 
     n50885 , n228647 , n228648 , n50888 , n50889 , n50890 , n50891 , n228653 , n228654 , n50894 , 
     n50895 , n50896 , n50897 , n228659 , n228660 , n50900 , n50901 , n50902 , n50903 , n228665 , 
     n228666 , n50906 , n228668 , n228669 , n50909 , n50910 , n50911 , n50912 , n228674 , n228675 , 
     n50915 , n50916 , n50917 , n50918 , n228680 , n228681 , n50921 , n228683 , n228684 , n50924 , 
     n50925 , n50926 , n50927 , n228689 , n228690 , n50930 , n50931 , n50932 , n50933 , n228695 , 
     n228696 , n50936 , n50937 , n50938 , n50939 , n50940 , n50941 , n50942 , n50943 , n50944 , 
     n50945 , n228707 , n228708 , n50948 , n50949 , n50950 , n50951 , n50952 , n50953 , n228715 , 
     n228716 , n50956 , n50957 , n50958 , n50959 , n228721 , n228722 , n50962 , n228724 , n228725 , 
     n50965 , n50966 , n50967 , n50968 , n50969 , n50970 , n228732 , n228733 , n50973 , n50974 , 
     n50975 , n50976 , n228738 , n228739 , n50979 , n50980 , n50981 , n50982 , n50983 , n50984 , 
     n228746 , n228747 , n50987 , n228749 , n228750 , n50990 , n50991 , n50992 , n50993 , n50994 , 
     n50995 , n50996 , n228758 , n228759 , n228760 , n228761 , n51001 , n51002 , n51003 , n51004 , 
     n228766 , n228767 , n51007 , n51008 , n51009 , n51010 , n228772 , n228773 , n51013 , n228775 , 
     n228776 , n51016 , n51017 , n51018 , n51019 , n51020 , n51021 , n228783 , n228784 , n51024 , 
     n51025 , n51026 , n51027 , n228789 , n228790 , n51030 , n51031 , n51032 , n51033 , n228795 , 
     n228796 , n51036 , n51037 , n51038 , n51039 , n228801 , n228802 , n51042 , n51043 , n51044 , 
     n51045 , n228807 , n228808 , n51048 , n51049 , n51050 , n51051 , n51052 , n51053 , n51054 , 
     n51055 , n228817 , n228818 , n51058 , n228820 , n51060 , n51061 , n51062 , n51063 , n51064 , 
     n51065 , n228827 , n228828 , n51068 , n51069 , n51070 , n51071 , n228833 , n228834 , n51074 , 
     n51075 , n51076 , n51077 , n51078 , n51079 , n51080 , n51081 , n228843 , n228844 , n51084 , 
     n51085 , n51086 , n51087 , n51088 , n51089 , n228851 , n228852 , n51092 , n51093 , n51094 , 
     n51095 , n228857 , n228858 , n51098 , n51099 , n51100 , n51101 , n228863 , n228864 , n51104 , 
     n51105 , n51106 , n51107 , n228869 , n228870 , n51110 , n51111 , n51112 , n51113 , n51114 , 
     n51115 , n228877 , n228878 , n51118 , n51119 , n51120 , n51121 , n51122 , n51123 , n51124 , 
     n51125 , n51126 , n228888 , n228889 , n51129 , n51130 , n51131 , n51132 , n228894 , n228895 , 
     n51135 , n51136 , n51137 , n51138 , n228900 , n228901 , n51141 , n51142 , n51143 , n51144 , 
     n51145 , n51146 , n228908 , n228909 , n51149 , n51150 , n51151 , n51152 , n51153 , n51154 , 
     n51155 , n228917 , n228918 , n51158 , n51159 , n51160 , n51161 , n228923 , n228924 , n51164 , 
     n51165 , n51166 , n51167 , n228929 , n228930 , n51170 , n51171 , n51172 , n51173 , n228935 , 
     n228936 , n51176 , n51177 , n51178 , n51179 , n51180 , n51181 , n51182 , n228944 , n228945 , 
     n51185 , n51186 , n51187 , n51188 , n228950 , n228951 , n51191 , n51192 , n51193 , n51194 , 
     n228956 , n228957 , n51197 , n51198 , n51199 , n51200 , n51201 , n51202 , n228964 , n228965 , 
     n51205 , n51206 , n51207 , n51208 , n228970 , n228971 , n51211 , n228973 , n228974 , n51214 , 
     n51215 , n51216 , n51217 , n51218 , n51219 , n228981 , n228982 , n51222 , n51223 , n51224 , 
     n51225 , n228987 , n228988 , n51228 , n51229 , n51230 , n51231 , n51232 , n51233 , n228995 , 
     n228996 , n51236 , n51237 , n51238 , n51239 , n51240 , n51241 , n229003 , n229004 , n51244 , 
     n51245 , n51246 , n51247 , n51248 , n51249 , n229011 , n229012 , n51252 , n229014 , n229015 , 
     n51255 , n51256 , n51257 , n51258 , n229020 , n229021 , n51261 , n51262 , n51263 , n51264 , 
     n51265 , n51266 , n229028 , n229029 , n51269 , n51270 , n51271 , n51272 , n51273 , n51274 , 
     n229036 , n229037 , n51277 , n229039 , n229040 , n51280 , n51281 , n51282 , n51283 , n51284 , 
     n51285 , n51286 , n51287 , n229049 , n229050 , n51290 , n51291 , n51292 , n51293 , n51294 , 
     n51295 , n229057 , n229058 , n51298 , n229060 , n229061 , n51301 , n229063 , n229064 , n51304 , 
     n51305 , n51306 , n51307 , n229069 , n229070 , n51310 , n51311 , n51312 , n51313 , n51314 , 
     n51315 , n229077 , n229078 , n51318 , n229080 , n229081 , n51321 , n51322 , n51323 , n229085 , 
     n229086 , n229087 , n229088 , n51328 , n51329 , n51330 , n51331 , n229093 , n229094 , n51334 , 
     n51335 , n51336 , n229098 , n229099 , n51339 , n51340 , n51341 , n51342 , n51343 , n229105 , 
     n229106 , n51346 , n51347 , n51348 , n51349 , n229111 , n229112 , n51352 , n51353 , n51354 , 
     n51355 , n51356 , n51357 , n51358 , n51359 , n229121 , n229122 , n51362 , n51363 , n51364 , 
     n51365 , n229127 , n229128 , n51368 , n51369 , n51370 , n51371 , n229133 , n229134 , n51374 , 
     n51375 , n51376 , n51377 , n229139 , n229140 , n51380 , n51381 , n51382 , n51383 , n229145 , 
     n229146 , n51386 , n229148 , n229149 , n51389 , n51390 , n51391 , n51392 , n229154 , n229155 , 
     n51395 , n51396 , n51397 , n51398 , n51399 , n51400 , n51401 , n51402 , n51403 , n229165 , 
     n229166 , n51406 , n51407 , n51408 , n51409 , n51410 , n51411 , n51412 , n229174 , n229175 , 
     n51415 , n229177 , n229178 , n51418 , n51419 , n51420 , n51421 , n51422 , n51423 , n51424 , 
     n51425 , n229187 , n229188 , n51428 , n229190 , n229191 , n51431 , n229193 , n229194 , n51434 , 
     n51435 , n51436 , n51437 , n229199 , n229200 , n51440 , n51441 , n51442 , n51443 , n51444 , 
     n51445 , n51446 , n51447 , n229209 , n229210 , n51450 , n51451 , n51452 , n51453 , n51454 , 
     n51455 , n229217 , n229218 , n51458 , n51459 , n51460 , n51461 , n51462 , n51463 , n229225 , 
     n229226 , n51466 , n51467 , n51468 , n51469 , n229231 , n229232 , n51472 , n229234 , n229235 , 
     n51475 , n51476 , n51477 , n51478 , n229240 , n229241 , n51481 , n51482 , n51483 , n51484 , 
     n229246 , n229247 , n51487 , n229249 , n229250 , n51490 , n51491 , n51492 , n51493 , n229255 , 
     n229256 , n51496 , n229258 , n229259 , n51499 , n51500 , n51501 , n51502 , n51503 , n229265 , 
     n229266 , n229267 , n229268 , n51508 , n51509 , n51510 , n51511 , n51512 , n51513 , n229275 , 
     n229276 , n51516 , n51517 , n51518 , n51519 , n229281 , n229282 , n51522 , n51523 , n51524 , 
     n51525 , n229287 , n229288 , n51528 , n51529 , n51530 , n51531 , n229293 , n229294 , n51534 , 
     n51535 , n51536 , n51537 , n229299 , n229300 , n51540 , n51541 , n51542 , n51543 , n229305 , 
     n229306 , n51546 , n51547 , n51548 , n51549 , n229311 , n229312 , n51552 , n51553 , n51554 , 
     n229316 , n229317 , n229318 , n229319 , n51559 , n51560 , n51561 , n51562 , n51563 , n51564 , 
     n229326 , n229327 , n51567 , n51568 , n51569 , n51570 , n51571 , n51572 , n51573 , n51574 , 
     n51575 , n229337 , n229338 , n229339 , n229340 , n51580 , n51581 , n51582 , n51583 , n51584 , 
     n51585 , n229347 , n229348 , n51588 , n51589 , n51590 , n51591 , n51592 , n51593 , n229355 , 
     n229356 , n51596 , n51597 , n51598 , n51599 , n229361 , n229362 , n51602 , n229364 , n229365 , 
     n51605 , n51606 , n51607 , n51608 , n229370 , n229371 , n51611 , n51612 , n51613 , n51614 , 
     n229376 , n229377 , n51617 , n51618 , n51619 , n51620 , n51621 , n51622 , n229384 , n229385 , 
     n51625 , n229387 , n229388 , n51628 , n229390 , n229391 , n51631 , n229393 , n229394 , n51634 , 
     n51635 , n51636 , n51637 , n51638 , n51639 , n229401 , n229402 , n51642 , n229404 , n229405 , 
     n51645 , n51646 , n51647 , n51648 , n51649 , n229411 , n229412 , n51652 , n51653 , n51654 , 
     n51655 , n51656 , n229418 , n229419 , n51659 , n229421 , n229422 , n51662 , n51663 , n51664 , 
     n51665 , n51666 , n229428 , n229429 , n51669 , n51670 , n51671 , n51672 , n229434 , n229435 , 
     n51675 , n229437 , n229438 , n51678 , n51679 , n229441 , n229442 , n51682 , n51683 , n51684 , 
     n51685 , n51686 , n51687 , n51688 , n51689 , n229451 , n229452 , n51692 , n51693 , n51694 , 
     n51695 , n229457 , n229458 , n51698 , n51699 , n51700 , n51701 , n229463 , n229464 , n51704 , 
     n229466 , n229467 , n51707 , n51708 , n51709 , n51710 , n229472 , n229473 , n51713 , n51714 , 
     n51715 , n51716 , n229478 , n229479 , n51719 , n229481 , n229482 , n51722 , n51723 , n51724 , 
     n51725 , n229487 , n229488 , n51728 , n51729 , n51730 , n51731 , n229493 , n229494 , n51734 , 
     n51735 , n51736 , n51737 , n229499 , n229500 , n51740 , n51741 , n51742 , n51743 , n229505 , 
     n229506 , n51746 , n51747 , n51748 , n51749 , n51750 , n229512 , n229513 , n51753 , n51754 , 
     n51755 , n51756 , n229518 , n229519 , n51759 , n229521 , n229522 , n51762 , n229524 , n229525 , 
     n51765 , n51766 , n51767 , n51768 , n51769 , n229531 , n229532 , n51772 , n51773 , n51774 , 
     n51775 , n229537 , n229538 , n51778 , n229540 , n229541 , n51781 , n51782 , n51783 , n51784 , 
     n51785 , n229547 , n229548 , n51788 , n51789 , n229551 , n229552 , n51792 , n51793 , n51794 , 
     n51795 , n51796 , n51797 , n229559 , n229560 , n51800 , n51801 , n51802 , n51803 , n51804 , 
     n51805 , n51806 , n51807 , n229569 , n229570 , n51810 , n51811 , n51812 , n51813 , n51814 , 
     n51815 , n229577 , n229578 , n51818 , n51819 , n51820 , n51821 , n229583 , n229584 , n51824 , 
     n51825 , n51826 , n51827 , n229589 , n229590 , n51830 , n51831 , n51832 , n51833 , n229595 , 
     n229596 , n51836 , n229598 , n229599 , n51839 , n51840 , n51841 , n229603 , n229604 , n51844 , 
     n51845 , n51846 , n51847 , n229609 , n229610 , n51850 , n51851 , n51852 , n51853 , n51854 , 
     n51855 , n229617 , n229618 , n51858 , n51859 , n51860 , n51861 , n229623 , n229624 , n51864 , 
     n51865 , n51866 , n51867 , n229629 , n229630 , n51870 , n229632 , n229633 , n51873 , n51874 , 
     n51875 , n51876 , n229638 , n229639 , n51879 , n51880 , n51881 , n51882 , n51883 , n51884 , 
     n51885 , n51886 , n229648 , n229649 , n51889 , n51890 , n51891 , n51892 , n229654 , n229655 , 
     n51895 , n51896 , n51897 , n51898 , n229660 , n229661 , n51901 , n51902 , n51903 , n51904 , 
     n51905 , n51906 , n51907 , n51908 , n229670 , n229671 , n51911 , n229673 , n51913 , n51914 , 
     n51915 , n51916 , n229678 , n229679 , n51919 , n51920 , n51921 , n51922 , n229684 , n229685 , 
     n51925 , n51926 , n51927 , n51928 , n51929 , n51930 , n229692 , n229693 , n51933 , n51934 , 
     n51935 , n51936 , n229698 , n229699 , n51939 , n51940 , n51941 , n51942 , n229704 , n229705 , 
     n51945 , n51946 , n51947 , n51948 , n229710 , n229711 , n51951 , n229713 , n229714 , n51954 , 
     n51955 , n51956 , n51957 , n51958 , n229720 , n229721 , n51961 , n51962 , n51963 , n51964 , 
     n229726 , n229727 , n51967 , n51968 , n51969 , n51970 , n51971 , n51972 , n229734 , n229735 , 
     n51975 , n51976 , n51977 , n51978 , n229740 , n229741 , n51981 , n229743 , n229744 , n51984 , 
     n229746 , n229747 , n51987 , n229749 , n51989 , n51990 , n51991 , n51992 , n229754 , n229755 , 
     n51995 , n51996 , n51997 , n51998 , n51999 , n52000 , n229762 , n229763 , n52003 , n229765 , 
     n229766 , n52006 , n52007 , n52008 , n52009 , n229771 , n229772 , n52012 , n52013 , n52014 , 
     n52015 , n229777 , n229778 , n52018 , n52019 , n52020 , n52021 , n229783 , n229784 , n52024 , 
     n52025 , n52026 , n52027 , n52028 , n52029 , n229791 , n229792 , n52032 , n52033 , n52034 , 
     n52035 , n229797 , n229798 , n52038 , n52039 , n52040 , n52041 , n52042 , n52043 , n229805 , 
     n229806 , n52046 , n52047 , n52048 , n52049 , n52050 , n52051 , n52052 , n52053 , n52054 , 
     n229816 , n229817 , n52057 , n52058 , n52059 , n52060 , n229822 , n229823 , n52063 , n52064 , 
     n52065 , n52066 , n229828 , n229829 , n52069 , n52070 , n52071 , n52072 , n52073 , n52074 , 
     n229836 , n229837 , n52077 , n229839 , n229840 , n52080 , n52081 , n52082 , n52083 , n52084 , 
     n229846 , n229847 , n52087 , n52088 , n52089 , n52090 , n229852 , n229853 , n52093 , n52094 , 
     n52095 , n52096 , n52097 , n52098 , n229860 , n229861 , n52101 , n52102 , n52103 , n52104 , 
     n229866 , n229867 , n52107 , n229869 , n229870 , n52110 , n52111 , n52112 , n52113 , n52114 , 
     n52115 , n229877 , n229878 , n52118 , n52119 , n52120 , n52121 , n229883 , n229884 , n52124 , 
     n52125 , n52126 , n52127 , n52128 , n52129 , n229891 , n229892 , n52132 , n52133 , n52134 , 
     n52135 , n52136 , n52137 , n229899 , n229900 , n52140 , n52141 , n52142 , n52143 , n229905 , 
     n229906 , n52146 , n52147 , n52148 , n52149 , n229911 , n229912 , n52152 , n229914 , n229915 , 
     n52155 , n52156 , n52157 , n52158 , n229920 , n229921 , n52161 , n229923 , n229924 , n52164 , 
     n52165 , n52166 , n52167 , n229929 , n229930 , n52170 , n52171 , n52172 , n52173 , n229935 , 
     n229936 , n52176 , n229938 , n229939 , n52179 , n52180 , n52181 , n52182 , n52183 , n52184 , 
     n52185 , n52186 , n52187 , n52188 , n229950 , n229951 , n52191 , n52192 , n52193 , n52194 , 
     n229956 , n229957 , n52197 , n52198 , n52199 , n52200 , n52201 , n52202 , n229964 , n229965 , 
     n229966 , n229967 , n52207 , n52208 , n52209 , n52210 , n52211 , n52212 , n229974 , n229975 , 
     n52215 , n52216 , n52217 , n52218 , n229980 , n229981 , n52221 , n52222 , n52223 , n52224 , 
     n52225 , n52226 , n52227 , n52228 , n52229 , n229991 , n229992 , n52232 , n52233 , n52234 , 
     n52235 , n229997 , n229998 , n52238 , n52239 , n52240 , n52241 , n230003 , n230004 , n52244 , 
     n230006 , n230007 , n52247 , n52248 , n52249 , n52250 , n52251 , n52252 , n52253 , n52254 , 
     n52255 , n52256 , n230018 , n230019 , n52259 , n52260 , n52261 , n52262 , n230024 , n230025 , 
     n52265 , n52266 , n52267 , n52268 , n52269 , n230031 , n230032 , n52272 , n52273 , n52274 , 
     n52275 , n230037 , n230038 , n52278 , n52279 , n52280 , n52281 , n230043 , n230044 , n52284 , 
     n52285 , n52286 , n52287 , n52288 , n52289 , n230051 , n230052 , n52292 , n52293 , n52294 , 
     n52295 , n230057 , n230058 , n52298 , n52299 , n52300 , n52301 , n230063 , n230064 , n52304 , 
     n52305 , n52306 , n52307 , n230069 , n230070 , n52310 , n52311 , n230073 , n230074 , n52314 , 
     n52315 , n52316 , n52317 , n52318 , n52319 , n230081 , n230082 , n52322 , n52323 , n52324 , 
     n52325 , n52326 , n230088 , n230089 , n52329 , n52330 , n52331 , n52332 , n230094 , n230095 , 
     n52335 , n52336 , n52337 , n52338 , n52339 , n52340 , n230102 , n230103 , n52343 , n52344 , 
     n52345 , n52346 , n52347 , n52348 , n52349 , n52350 , n230112 , n230113 , n52353 , n52354 , 
     n52355 , n52356 , n230118 , n230119 , n52359 , n52360 , n52361 , n52362 , n230124 , n230125 , 
     n52365 , n52366 , n52367 , n52368 , n230130 , n230131 , n52371 , n52372 , n52373 , n52374 , 
     n52375 , n52376 , n52377 , n52378 , n52379 , n230141 , n230142 , n230143 , n230144 , n52384 , 
     n52385 , n52386 , n52387 , n230149 , n230150 , n52390 , n230152 , n230153 , n52393 , n230155 , 
     n230156 , n52396 , n52397 , n52398 , n52399 , n230161 , n230162 , n52402 , n52403 , n52404 , 
     n52405 , n230167 , n230168 , n52408 , n52409 , n52410 , n52411 , n52412 , n52413 , n230175 , 
     n230176 , n52416 , n230178 , n230179 , n52419 , n52420 , n52421 , n52422 , n230184 , n230185 , 
     n52425 , n52426 , n52427 , n52428 , n52429 , n52430 , n52431 , n52432 , n52433 , n230195 , 
     n230196 , n52436 , n230198 , n230199 , n52439 , n230201 , n230202 , n52442 , n230204 , n230205 , 
     n52445 , n230207 , n230208 , n230209 , n230210 , n52450 , n52451 , n52452 , n52453 , n230215 , 
     n230216 , n52456 , n52457 , n52458 , n52459 , n230221 , n230222 , n52462 , n52463 , n52464 , 
     n52465 , n230227 , n230228 , n52468 , n52469 , n52470 , n52471 , n230233 , n230234 , n52474 , 
     n230236 , n230237 , n52477 , n230239 , n230240 , n52480 , n230242 , n230243 , n52483 , n52484 , 
     n52485 , n52486 , n230248 , n230249 , n52489 , n52490 , n52491 , n52492 , n230254 , n230255 , 
     n52495 , n52496 , n52497 , n52498 , n230260 , n230261 , n52501 , n52502 , n52503 , n52504 , 
     n52505 , n52506 , n230268 , n230269 , n52509 , n230271 , n230272 , n52512 , n52513 , n52514 , 
     n52515 , n52516 , n52517 , n230279 , n230280 , n52520 , n52521 , n52522 , n52523 , n230285 , 
     n230286 , n52526 , n230288 , n230289 , n52529 , n52530 , n52531 , n52532 , n230294 , n230295 , 
     n52535 , n52536 , n52537 , n52538 , n230300 , n230301 , n52541 , n52542 , n52543 , n230305 , 
     n230306 , n230307 , n230308 , n52548 , n52549 , n52550 , n52551 , n230313 , n230314 , n52554 , 
     n52555 , n52556 , n52557 , n230319 , n230320 , n52560 , n52561 , n52562 , n52563 , n230325 , 
     n230326 , n52566 , n52567 , n52568 , n52569 , n52570 , n52571 , n230333 , n230334 , n52574 , 
     n52575 , n52576 , n52577 , n230339 , n230340 , n52580 , n52581 , n52582 , n52583 , n52584 , 
     n52585 , n230347 , n230348 , n52588 , n52589 , n52590 , n52591 , n230353 , n230354 , n52594 , 
     n52595 , n52596 , n52597 , n52598 , n52599 , n230361 , n230362 , n52602 , n52603 , n52604 , 
     n52605 , n230367 , n230368 , n52608 , n52609 , n52610 , n52611 , n230373 , n230374 , n52614 , 
     n52615 , n52616 , n52617 , n52618 , n230380 , n230381 , n52621 , n52622 , n52623 , n52624 , 
     n230386 , n230387 , n52627 , n52628 , n52629 , n52630 , n52631 , n52632 , n230394 , n230395 , 
     n52635 , n52636 , n52637 , n52638 , n52639 , n230401 , n230402 , n52642 , n52643 , n52644 , 
     n52645 , n230407 , n230408 , n52648 , n52649 , n52650 , n52651 , n230413 , n230414 , n52654 , 
     n230416 , n230417 , n52657 , n52658 , n52659 , n52660 , n230422 , n230423 , n52663 , n52664 , 
     n52665 , n52666 , n230428 , n230429 , n52669 , n52670 , n52671 , n52672 , n230434 , n230435 , 
     n52675 , n230437 , n230438 , n52678 , n52679 , n52680 , n52681 , n230443 , n230444 , n52684 , 
     n52685 , n52686 , n52687 , n230449 , n230450 , n52690 , n230452 , n230453 , n52693 , n230455 , 
     n230456 , n52696 , n230458 , n230459 , n52699 , n230461 , n230462 , n52702 , n52703 , n52704 , 
     n52705 , n52706 , n230468 , n230469 , n52709 , n52710 , n52711 , n52712 , n52713 , n52714 , 
     n52715 , n230477 , n230478 , n52718 , n230480 , n230481 , n52721 , n52722 , n52723 , n52724 , 
     n52725 , n230487 , n230488 , n52728 , n52729 , n52730 , n52731 , n230493 , n230494 , n52734 , 
     n52735 , n230497 , n230498 , n52738 , n52739 , n52740 , n52741 , n52742 , n230504 , n230505 , 
     n52745 , n52746 , n52747 , n52748 , n52749 , n230511 , n230512 , n52752 , n52753 , n52754 , 
     n52755 , n52756 , n52757 , n230519 , n230520 , n52760 , n52761 , n52762 , n52763 , n52764 , 
     n52765 , n52766 , n52767 , n52768 , n52769 , n52770 , n52771 , n230533 , n230534 , n52774 , 
     n230536 , n230537 , n52777 , n52778 , n52779 , n52780 , n230542 , n230543 , n52783 , n230545 , 
     n230546 , n52786 , n52787 , n52788 , n52789 , n230551 , n230552 , n52792 , n52793 , n52794 , 
     n52795 , n230557 , n230558 , n52798 , n52799 , n52800 , n52801 , n230563 , n230564 , n52804 , 
     n52805 , n52806 , n52807 , n52808 , n52809 , n230571 , n230572 , n52812 , n230574 , n230575 , 
     n52815 , n52816 , n52817 , n52818 , n52819 , n52820 , n230582 , n230583 , n52823 , n52824 , 
     n52825 , n52826 , n230588 , n230589 , n52829 , n230591 , n230592 , n52832 , n230594 , n230595 , 
     n52835 , n230597 , n52837 , n52838 , n52839 , n52840 , n230602 , n230603 , n52843 , n52844 , 
     n52845 , n52846 , n230608 , n230609 , n52849 , n52850 , n52851 , n52852 , n230614 , n230615 , 
     n52855 , n230617 , n230618 , n52858 , n52859 , n52860 , n52861 , n230623 , n230624 , n52864 , 
     n52865 , n52866 , n52867 , n230629 , n230630 , n52870 , n52871 , n52872 , n52873 , n230635 , 
     n230636 , n52876 , n52877 , n52878 , n52879 , n52880 , n52881 , n230643 , n230644 , n52884 , 
     n52885 , n52886 , n52887 , n230649 , n230650 , n52890 , n52891 , n52892 , n52893 , n52894 , 
     n52895 , n230657 , n230658 , n52898 , n52899 , n52900 , n52901 , n230663 , n230664 , n52904 , 
     n230666 , n230667 , n52907 , n230669 , n230670 , n52910 , n52911 , n52912 , n230674 , n230675 , 
     n52915 , n52916 , n52917 , n52918 , n230680 , n230681 , n52921 , n52922 , n52923 , n52924 , 
     n230686 , n230687 , n52927 , n230689 , n230690 , n52930 , n230692 , n230693 , n52933 , n52934 , 
     n52935 , n52936 , n52937 , n52938 , n230700 , n230701 , n52941 , n52942 , n52943 , n52944 , 
     n230706 , n230707 , n52947 , n52948 , n52949 , n52950 , n230712 , n230713 , n52953 , n52954 , 
     n52955 , n52956 , n230718 , n230719 , n52959 , n52960 , n52961 , n52962 , n52963 , n230725 , 
     n230726 , n52966 , n52967 , n52968 , n52969 , n230731 , n230732 , n52972 , n52973 , n52974 , 
     n52975 , n230737 , n230738 , n52978 , n230740 , n52980 , n52981 , n52982 , n52983 , n230745 , 
     n230746 , n52986 , n52987 , n52988 , n52989 , n52990 , n52991 , n230753 , n230754 , n52994 , 
     n52995 , n52996 , n52997 , n52998 , n52999 , n53000 , n53001 , n53002 , n230764 , n230765 , 
     n230766 , n230767 , n53007 , n53008 , n53009 , n53010 , n53011 , n53012 , n53013 , n53014 , 
     n53015 , n230777 , n230778 , n230779 , n230780 , n53020 , n230782 , n230783 , n53023 , n230785 , 
     n230786 , n53026 , n53027 , n53028 , n53029 , n230791 , n230792 , n53032 , n53033 , n53034 , 
     n53035 , n230797 , n230798 , n53038 , n53039 , n53040 , n53041 , n53042 , n53043 , n53044 , 
     n53045 , n230807 , n230808 , n230809 , n230810 , n53050 , n230812 , n230813 , n53053 , n53054 , 
     n53055 , n53056 , n230818 , n230819 , n53059 , n230821 , n230822 , n53062 , n53063 , n53064 , 
     n53065 , n230827 , n230828 , n53068 , n53069 , n53070 , n53071 , n230833 , n230834 , n53074 , 
     n53075 , n53076 , n53077 , n230839 , n230840 , n53080 , n53081 , n53082 , n53083 , n230845 , 
     n230846 , n53086 , n53087 , n53088 , n53089 , n230851 , n230852 , n53092 , n230854 , n230855 , 
     n53095 , n230857 , n230858 , n53098 , n53099 , n53100 , n53101 , n230863 , n230864 , n53104 , 
     n53105 , n53106 , n53107 , n230869 , n230870 , n53110 , n53111 , n53112 , n53113 , n230875 , 
     n230876 , n53116 , n53117 , n53118 , n53119 , n230881 , n230882 , n53122 , n53123 , n53124 , 
     n53125 , n230887 , n230888 , n53128 , n53129 , n53130 , n53131 , n230893 , n230894 , n53134 , 
     n53135 , n53136 , n53137 , n230899 , n230900 , n53140 , n230902 , n230903 , n53143 , n230905 , 
     n230906 , n53146 , n53147 , n53148 , n53149 , n230911 , n230912 , n53152 , n230914 , n230915 , 
     n53155 , n53156 , n53157 , n53158 , n230920 , n230921 , n53161 , n53162 , n53163 , n53164 , 
     n230926 , n230927 , n53167 , n53168 , n53169 , n53170 , n53171 , n230933 , n230934 , n53174 , 
     n53175 , n53176 , n53177 , n53178 , n230940 , n230941 , n53181 , n53182 , n53183 , n53184 , 
     n53185 , n53186 , n53187 , n53188 , n53189 , n53190 , n230952 , n230953 , n53193 , n53194 , 
     n230956 , n230957 , n53197 , n53198 , n53199 , n53200 , n53201 , n53202 , n53203 , n230965 , 
     n230966 , n53206 , n230968 , n230969 , n53209 , n53210 , n53211 , n53212 , n53213 , n53214 , 
     n53215 , n53216 , n53217 , n53218 , n230980 , n230981 , n53221 , n53222 , n53223 , n53224 , 
     n230986 , n230987 , n53227 , n53228 , n53229 , n53230 , n230992 , n230993 , n53233 , n230995 , 
     n230996 , n53236 , n230998 , n230999 , n53239 , n231001 , n231002 , n53242 , n53243 , n53244 , 
     n53245 , n231007 , n231008 , n53248 , n53249 , n53250 , n53251 , n231013 , n231014 , n53254 , 
     n53255 , n53256 , n53257 , n231019 , n231020 , n53260 , n53261 , n53262 , n53263 , n231025 , 
     n231026 , n53266 , n53267 , n53268 , n53269 , n231031 , n231032 , n53272 , n53273 , n53274 , 
     n53275 , n231037 , n231038 , n53278 , n231040 , n231041 , n53281 , n53282 , n53283 , n53284 , 
     n231046 , n231047 , n53287 , n53288 , n53289 , n53290 , n231052 , n231053 , n53293 , n53294 , 
     n53295 , n53296 , n53297 , n53298 , n231060 , n231061 , n53301 , n53302 , n53303 , n53304 , 
     n231066 , n231067 , n53307 , n53308 , n53309 , n53310 , n231072 , n231073 , n53313 , n53314 , 
     n53315 , n53316 , n231078 , n231079 , n53319 , n53320 , n53321 , n53322 , n53323 , n53324 , 
     n231086 , n231087 , n53327 , n53328 , n53329 , n53330 , n53331 , n53332 , n231094 , n231095 , 
     n231096 , n231097 , n53337 , n53338 , n53339 , n53340 , n231102 , n231103 , n53343 , n53344 , 
     n53345 , n53346 , n231108 , n231109 , n53349 , n53350 , n53351 , n53352 , n231114 , n231115 , 
     n53355 , n53356 , n53357 , n53358 , n231120 , n231121 , n53361 , n53362 , n53363 , n53364 , 
     n231126 , n231127 , n53367 , n53368 , n53369 , n53370 , n231132 , n231133 , n53373 , n231135 , 
     n231136 , n231137 , n231138 , n53378 , n53379 , n53380 , n231142 , n231143 , n231144 , n231145 , 
     n53385 , n53386 , n53387 , n53388 , n53389 , n53390 , n231152 , n231153 , n53393 , n231155 , 
     n231156 , n53396 , n231158 , n231159 , n53399 , n53400 , n53401 , n53402 , n231164 , n231165 , 
     n53405 , n53406 , n53407 , n53408 , n231170 , n231171 , n53411 , n53412 , n53413 , n53414 , 
     n231176 , n231177 , n53417 , n231179 , n231180 , n53420 , n231182 , n231183 , n53423 , n53424 , 
     n53425 , n53426 , n53427 , n53428 , n231190 , n231191 , n53431 , n53432 , n53433 , n53434 , 
     n53435 , n53436 , n231198 , n231199 , n53439 , n53440 , n53441 , n53442 , n231204 , n231205 , 
     n53445 , n231207 , n231208 , n53448 , n231210 , n231211 , n53451 , n53452 , n53453 , n53454 , 
     n231216 , n231217 , n53457 , n53458 , n53459 , n53460 , n231222 , n231223 , n53463 , n53464 , 
     n53465 , n53466 , n53467 , n53468 , n231230 , n231231 , n53471 , n53472 , n53473 , n53474 , 
     n231236 , n231237 , n53477 , n231239 , n53479 , n53480 , n53481 , n53482 , n231244 , n231245 , 
     n53485 , n53486 , n53487 , n53488 , n53489 , n53490 , n53491 , n53492 , n231254 , n231255 , 
     n53495 , n231257 , n231258 , n53498 , n53499 , n53500 , n53501 , n231263 , n231264 , n53504 , 
     n53505 , n53506 , n53507 , n231269 , n231270 , n53510 , n53511 , n53512 , n53513 , n231275 , 
     n231276 , n53516 , n53517 , n53518 , n53519 , n231281 , n231282 , n53522 , n53523 , n231285 , 
     n231286 , n53526 , n53527 , n53528 , n53529 , n231291 , n231292 , n53532 , n53533 , n53534 , 
     n53535 , n231297 , n231298 , n53538 , n53539 , n53540 , n53541 , n231303 , n231304 , n53544 , 
     n53545 , n53546 , n53547 , n231309 , n231310 , n53550 , n53551 , n53552 , n53553 , n231315 , 
     n231316 , n53556 , n53557 , n53558 , n53559 , n231321 , n231322 , n53562 , n231324 , n231325 , 
     n231326 , n231327 , n53567 , n231329 , n231330 , n53570 , n231332 , n53572 , n231334 , n231335 , 
     n53575 , n53576 , n53577 , n53578 , n231340 , n231341 , n53581 , n53582 , n53583 , n53584 , 
     n231346 , n231347 , n53587 , n53588 , n53589 , n53590 , n231352 , n231353 , n53593 , n53594 , 
     n53595 , n53596 , n231358 , n231359 , n53599 , n231361 , n231362 , n53602 , n53603 , n53604 , 
     n53605 , n231367 , n231368 , n53608 , n53609 , n53610 , n53611 , n231373 , n231374 , n53614 , 
     n53615 , n53616 , n53617 , n231379 , n231380 , n53620 , n53621 , n53622 , n53623 , n231385 , 
     n231386 , n53626 , n53627 , n53628 , n53629 , n231391 , n231392 , n53632 , n53633 , n53634 , 
     n53635 , n231397 , n231398 , n53638 , n53639 , n53640 , n53641 , n231403 , n231404 , n53644 , 
     n53645 , n53646 , n53647 , n53648 , n231410 , n231411 , n231412 , n231413 , n53653 , n53654 , 
     n53655 , n53656 , n53657 , n53658 , n53659 , n231421 , n231422 , n231423 , n231424 , n53664 , 
     n53665 , n53666 , n53667 , n53668 , n53669 , n53670 , n231432 , n231433 , n53673 , n53674 , 
     n53675 , n53676 , n231438 , n231439 , n53679 , n53680 , n53681 , n53682 , n231444 , n231445 , 
     n53685 , n53686 , n53687 , n53688 , n231450 , n231451 , n53691 , n53692 , n53693 , n53694 , 
     n53695 , n53696 , n53697 , n231459 , n231460 , n53700 , n53701 , n53702 , n53703 , n231465 , 
     n231466 , n53706 , n231468 , n231469 , n53709 , n53710 , n53711 , n53712 , n231474 , n231475 , 
     n53715 , n53716 , n53717 , n53718 , n231480 , n231481 , n53721 , n231483 , n231484 , n53724 , 
     n53725 , n53726 , n53727 , n231489 , n231490 , n53730 , n53731 , n53732 , n53733 , n53734 , 
     n53735 , n53736 , n53737 , n231499 , n231500 , n53740 , n231502 , n231503 , n53743 , n231505 , 
     n231506 , n53746 , n231508 , n231509 , n53749 , n53750 , n53751 , n53752 , n231514 , n231515 , 
     n53755 , n53756 , n53757 , n53758 , n231520 , n231521 , n53761 , n53762 , n53763 , n53764 , 
     n53765 , n53766 , n231528 , n231529 , n231530 , n231531 , n53771 , n53772 , n53773 , n53774 , 
     n231536 , n231537 , n53777 , n53778 , n53779 , n53780 , n231542 , n231543 , n53783 , n53784 , 
     n53785 , n53786 , n53787 , n53788 , n53789 , n231551 , n231552 , n231553 , n231554 , n53794 , 
     n53795 , n53796 , n53797 , n231559 , n231560 , n53800 , n53801 , n53802 , n53803 , n231565 , 
     n231566 , n53806 , n53807 , n53808 , n53809 , n53810 , n53811 , n231573 , n231574 , n53814 , 
     n53815 , n53816 , n53817 , n231579 , n231580 , n53820 , n53821 , n53822 , n53823 , n231585 , 
     n231586 , n53826 , n53827 , n231589 , n231590 , n231591 , n231592 , n53832 , n53833 , n53834 , 
     n53835 , n231597 , n231598 , n53838 , n53839 , n53840 , n53841 , n231603 , n231604 , n53844 , 
     n53845 , n53846 , n53847 , n231609 , n231610 , n53850 , n53851 , n53852 , n53853 , n231615 , 
     n231616 , n53856 , n53857 , n53858 , n53859 , n231621 , n231622 , n53862 , n53863 , n53864 , 
     n53865 , n231627 , n231628 , n53868 , n53869 , n53870 , n53871 , n231633 , n231634 , n53874 , 
     n53875 , n53876 , n53877 , n231639 , n231640 , n53880 , n53881 , n53882 , n53883 , n231645 , 
     n231646 , n53886 , n231648 , n231649 , n53889 , n53890 , n53891 , n53892 , n231654 , n231655 , 
     n53895 , n231657 , n231658 , n53898 , n53899 , n53900 , n53901 , n231663 , n231664 , n53904 , 
     n53905 , n53906 , n53907 , n231669 , n231670 , n53910 , n53911 , n53912 , n53913 , n231675 , 
     n231676 , n53916 , n53917 , n53918 , n53919 , n231681 , n231682 , n53922 , n53923 , n53924 , 
     n53925 , n231687 , n231688 , n53928 , n231690 , n231691 , n53931 , n231693 , n231694 , n53934 , 
     n53935 , n53936 , n53937 , n231699 , n231700 , n53940 , n231702 , n231703 , n53943 , n53944 , 
     n53945 , n53946 , n231708 , n231709 , n53949 , n53950 , n53951 , n53952 , n231714 , n231715 , 
     n53955 , n53956 , n53957 , n53958 , n53959 , n53960 , n231722 , n231723 , n53963 , n53964 , 
     n53965 , n53966 , n231728 , n231729 , n53969 , n53970 , n53971 , n53972 , n231734 , n231735 , 
     n53975 , n53976 , n53977 , n53978 , n231740 , n231741 , n53981 , n53982 , n53983 , n53984 , 
     n231746 , n231747 , n231748 , n231749 , n53989 , n53990 , n53991 , n53992 , n231754 , n231755 , 
     n53995 , n53996 , n53997 , n53998 , n231760 , n231761 , n54001 , n54002 , n54003 , n54004 , 
     n54005 , n54006 , n231768 , n231769 , n54009 , n54010 , n54011 , n54012 , n54013 , n231775 , 
     n231776 , n54016 , n54017 , n54018 , n54019 , n231781 , n231782 , n231783 , n231784 , n54024 , 
     n231786 , n231787 , n54027 , n231789 , n231790 , n54030 , n54031 , n54032 , n54033 , n231795 , 
     n231796 , n54036 , n54037 , n54038 , n54039 , n54040 , n231802 , n231803 , n54043 , n54044 , 
     n54045 , n54046 , n54047 , n231809 , n231810 , n54050 , n54051 , n54052 , n54053 , n231815 , 
     n231816 , n54056 , n54057 , n54058 , n54059 , n231821 , n231822 , n54062 , n231824 , n231825 , 
     n54065 , n231827 , n231828 , n54068 , n54069 , n54070 , n54071 , n231833 , n231834 , n54074 , 
     n54075 , n54076 , n54077 , n231839 , n231840 , n54080 , n54081 , n54082 , n54083 , n231845 , 
     n231846 , n54086 , n54087 , n54088 , n54089 , n231851 , n231852 , n54092 , n231854 , n231855 , 
     n54095 , n54096 , n54097 , n54098 , n231860 , n231861 , n54101 , n54102 , n54103 , n54104 , 
     n54105 , n54106 , n231868 , n231869 , n54109 , n54110 , n54111 , n54112 , n231874 , n231875 , 
     n54115 , n54116 , n54117 , n54118 , n231880 , n231881 , n54121 , n54122 , n54123 , n54124 , 
     n54125 , n54126 , n54127 , n54128 , n54129 , n231891 , n231892 , n231893 , n231894 , n54134 , 
     n231896 , n231897 , n54137 , n54138 , n54139 , n54140 , n231902 , n231903 , n54143 , n54144 , 
     n54145 , n54146 , n54147 , n54148 , n231910 , n231911 , n54151 , n54152 , n54153 , n54154 , 
     n54155 , n231917 , n231918 , n54158 , n231920 , n231921 , n54161 , n231923 , n231924 , n54164 , 
     n54165 , n54166 , n54167 , n231929 , n231930 , n54170 , n54171 , n54172 , n54173 , n54174 , 
     n54175 , n54176 , n54177 , n231939 , n231940 , n54180 , n54181 , n54182 , n54183 , n231945 , 
     n231946 , n54186 , n54187 , n54188 , n54189 , n231951 , n231952 , n54192 , n54193 , n54194 , 
     n54195 , n231957 , n231958 , n54198 , n54199 , n54200 , n54201 , n231963 , n231964 , n54204 , 
     n231966 , n54206 , n54207 , n54208 , n54209 , n54210 , n54211 , n231973 , n231974 , n54214 , 
     n231976 , n231977 , n54217 , n54218 , n54219 , n54220 , n54221 , n54222 , n231984 , n231985 , 
     n54225 , n54226 , n54227 , n54228 , n231990 , n231991 , n54231 , n54232 , n54233 , n54234 , 
     n231996 , n231997 , n54237 , n54238 , n54239 , n54240 , n232002 , n232003 , n54243 , n54244 , 
     n54245 , n54246 , n232008 , n232009 , n54249 , n232011 , n232012 , n54252 , n232014 , n54254 , 
     n54255 , n54256 , n54257 , n54258 , n232020 , n232021 , n54261 , n54262 , n54263 , n54264 , 
     n54265 , n54266 , n232028 , n232029 , n54269 , n54270 , n54271 , n54272 , n54273 , n232035 , 
     n232036 , n54276 , n54277 , n54278 , n54279 , n232041 , n232042 , n54282 , n54283 , n54284 , 
     n54285 , n232047 , n232048 , n54288 , n54289 , n54290 , n54291 , n232053 , n232054 , n54294 , 
     n54295 , n54296 , n54297 , n232059 , n232060 , n54300 , n54301 , n54302 , n54303 , n232065 , 
     n232066 , n54306 , n54307 , n54308 , n54309 , n232071 , n232072 , n54312 , n54313 , n54314 , 
     n54315 , n232077 , n232078 , n54318 , n54319 , n54320 , n54321 , n232083 , n232084 , n54324 , 
     n54325 , n54326 , n54327 , n232089 , n232090 , n54330 , n54331 , n54332 , n54333 , n232095 , 
     n232096 , n54336 , n54337 , n54338 , n54339 , n232101 , n232102 , n54342 , n54343 , n54344 , 
     n54345 , n54346 , n232108 , n232109 , n232110 , n232111 , n54351 , n232113 , n232114 , n54354 , 
     n54355 , n54356 , n54357 , n232119 , n232120 , n54360 , n232122 , n232123 , n54363 , n54364 , 
     n54365 , n54366 , n232128 , n232129 , n54369 , n54370 , n54371 , n54372 , n232134 , n232135 , 
     n54375 , n54376 , n54377 , n54378 , n232140 , n232141 , n54381 , n54382 , n54383 , n54384 , 
     n232146 , n232147 , n54387 , n232149 , n232150 , n54390 , n232152 , n232153 , n54393 , n232155 , 
     n232156 , n54396 , n54397 , n54398 , n54399 , n232161 , n232162 , n54402 , n54403 , n54404 , 
     n54405 , n232167 , n232168 , n54408 , n54409 , n54410 , n54411 , n232173 , n232174 , n54414 , 
     n54415 , n54416 , n54417 , n232179 , n232180 , n54420 , n54421 , n54422 , n54423 , n232185 , 
     n232186 , n54426 , n54427 , n54428 , n54429 , n232191 , n232192 , n54432 , n54433 , n54434 , 
     n54435 , n232197 , n232198 , n54438 , n54439 , n54440 , n54441 , n232203 , n232204 , n54444 , 
     n54445 , n54446 , n54447 , n232209 , n232210 , n54450 , n54451 , n54452 , n54453 , n232215 , 
     n232216 , n54456 , n54457 , n54458 , n54459 , n232221 , n232222 , n54462 , n232224 , n232225 , 
     n54465 , n232227 , n232228 , n54468 , n54469 , n54470 , n54471 , n232233 , n232234 , n54474 , 
     n54475 , n54476 , n54477 , n232239 , n232240 , n54480 , n232242 , n232243 , n54483 , n54484 , 
     n54485 , n54486 , n232248 , n232249 , n54489 , n54490 , n54491 , n54492 , n232254 , n232255 , 
     n54495 , n54496 , n54497 , n54498 , n232260 , n232261 , n54501 , n54502 , n54503 , n54504 , 
     n232266 , n232267 , n54507 , n54508 , n54509 , n54510 , n232272 , n232273 , n54513 , n54514 , 
     n54515 , n54516 , n232278 , n232279 , n54519 , n232281 , n232282 , n54522 , n232284 , n232285 , 
     n54525 , n54526 , n54527 , n54528 , n232290 , n232291 , n54531 , n232293 , n232294 , n54534 , 
     n54535 , n54536 , n54537 , n232299 , n232300 , n54540 , n54541 , n54542 , n54543 , n232305 , 
     n232306 , n54546 , n54547 , n54548 , n54549 , n232311 , n232312 , n54552 , n54553 , n54554 , 
     n54555 , n232317 , n232318 , n232319 , n232320 , n54560 , n54561 , n54562 , n54563 , n232325 , 
     n232326 , n54566 , n54567 , n54568 , n54569 , n232331 , n232332 , n54572 , n54573 , n54574 , 
     n54575 , n232337 , n232338 , n54578 , n54579 , n54580 , n54581 , n232343 , n232344 , n54584 , 
     n54585 , n54586 , n54587 , n232349 , n232350 , n54590 , n232352 , n232353 , n54593 , n54594 , 
     n54595 , n54596 , n54597 , n54598 , n54599 , n54600 , n54601 , n54602 , n54603 , n232365 , 
     n232366 , n232367 , n232368 , n54608 , n54609 , n54610 , n54611 , n232373 , n232374 , n54614 , 
     n54615 , n54616 , n54617 , n232379 , n232380 , n54620 , n54621 , n54622 , n54623 , n232385 , 
     n232386 , n54626 , n54627 , n54628 , n54629 , n232391 , n232392 , n54632 , n54633 , n54634 , 
     n54635 , n232397 , n232398 , n54638 , n54639 , n54640 , n54641 , n232403 , n232404 , n54644 , 
     n54645 , n54646 , n54647 , n232409 , n232410 , n54650 , n232412 , n232413 , n54653 , n54654 , 
     n54655 , n54656 , n232418 , n232419 , n54659 , n54660 , n54661 , n54662 , n54663 , n54664 , 
     n232426 , n232427 , n54667 , n54668 , n54669 , n54670 , n232432 , n232433 , n54673 , n232435 , 
     n232436 , n54676 , n54677 , n54678 , n54679 , n232441 , n232442 , n54682 , n232444 , n232445 , 
     n54685 , n232447 , n232448 , n54688 , n54689 , n54690 , n54691 , n54692 , n232454 , n232455 , 
     n54695 , n54696 , n54697 , n54698 , n54699 , n232461 , n232462 , n54702 , n54703 , n54704 , 
     n54705 , n54706 , n54707 , n54708 , n232470 , n232471 , n54711 , n54712 , n54713 , n54714 , 
     n232476 , n232477 , n54717 , n54718 , n54719 , n54720 , n232482 , n232483 , n54723 , n54724 , 
     n54725 , n54726 , n232488 , n232489 , n54729 , n54730 , n54731 , n54732 , n54733 , n54734 , 
     n232496 , n232497 , n54737 , n54738 , n54739 , n54740 , n232502 , n232503 , n54743 , n54744 , 
     n54745 , n54746 , n54747 , n54748 , n54749 , n54750 , n232512 , n232513 , n232514 , n232515 , 
     n54755 , n232517 , n232518 , n54758 , n232520 , n232521 , n54761 , n232523 , n232524 , n54764 , 
     n54765 , n232527 , n232528 , n54768 , n54769 , n54770 , n54771 , n54772 , n54773 , n54774 , 
     n54775 , n232537 , n232538 , n54778 , n54779 , n54780 , n54781 , n232543 , n232544 , n54784 , 
     n54785 , n54786 , n54787 , n232549 , n232550 , n54790 , n54791 , n54792 , n54793 , n232555 , 
     n232556 , n54796 , n232558 , n232559 , n54799 , n232561 , n232562 , n54802 , n54803 , n54804 , 
     n54805 , n232567 , n232568 , n54808 , n54809 , n54810 , n54811 , n232573 , n232574 , n54814 , 
     n54815 , n54816 , n54817 , n232579 , n232580 , n54820 , n232582 , n232583 , n54823 , n54824 , 
     n54825 , n54826 , n232588 , n232589 , n54829 , n54830 , n54831 , n54832 , n232594 , n232595 , 
     n54835 , n54836 , n54837 , n54838 , n232600 , n232601 , n54841 , n54842 , n54843 , n54844 , 
     n232606 , n232607 , n54847 , n54848 , n54849 , n54850 , n54851 , n54852 , n54853 , n54854 , 
     n54855 , n232617 , n232618 , n54858 , n54859 , n54860 , n54861 , n232623 , n232624 , n54864 , 
     n232626 , n232627 , n54867 , n54868 , n54869 , n54870 , n54871 , n232633 , n232634 , n54874 , 
     n54875 , n54876 , n54877 , n232639 , n232640 , n54880 , n54881 , n232643 , n232644 , n54884 , 
     n54885 , n54886 , n54887 , n232649 , n232650 , n54890 , n54891 , n54892 , n54893 , n232655 , 
     n232656 , n54896 , n232658 , n232659 , n54899 , n54900 , n54901 , n54902 , n232664 , n232665 , 
     n54905 , n54906 , n54907 , n54908 , n232670 , n232671 , n54911 , n54912 , n54913 , n54914 , 
     n232676 , n232677 , n54917 , n54918 , n54919 , n54920 , n232682 , n232683 , n54923 , n54924 , 
     n54925 , n54926 , n54927 , n232689 , n232690 , n232691 , n232692 , n54932 , n232694 , n232695 , 
     n54935 , n232697 , n232698 , n54938 , n54939 , n54940 , n54941 , n232703 , n232704 , n54944 , 
     n54945 , n232707 , n232708 , n54948 , n54949 , n54950 , n54951 , n232713 , n232714 , n54954 , 
     n54955 , n54956 , n54957 , n232719 , n232720 , n54960 , n54961 , n54962 , n54963 , n232725 , 
     n232726 , n54966 , n232728 , n232729 , n54969 , n54970 , n54971 , n54972 , n232734 , n232735 , 
     n54975 , n54976 , n54977 , n54978 , n232740 , n232741 , n54981 , n54982 , n54983 , n54984 , 
     n232746 , n232747 , n54987 , n232749 , n54989 , n54990 , n54991 , n54992 , n54993 , n54994 , 
     n232756 , n232757 , n54997 , n54998 , n54999 , n55000 , n232762 , n232763 , n55003 , n55004 , 
     n55005 , n55006 , n55007 , n55008 , n55009 , n55010 , n55011 , n232773 , n232774 , n232775 , 
     n232776 , n55016 , n232778 , n232779 , n55019 , n55020 , n55021 , n55022 , n232784 , n232785 , 
     n55025 , n55026 , n55027 , n55028 , n232790 , n232791 , n55031 , n55032 , n55033 , n55034 , 
     n232796 , n232797 , n55037 , n55038 , n55039 , n55040 , n232802 , n232803 , n55043 , n55044 , 
     n55045 , n55046 , n55047 , n55048 , n232810 , n232811 , n232812 , n232813 , n55053 , n232815 , 
     n232816 , n55056 , n232818 , n232819 , n55059 , n55060 , n55061 , n55062 , n55063 , n232825 , 
     n232826 , n55066 , n55067 , n55068 , n55069 , n55070 , n55071 , n232833 , n232834 , n55074 , 
     n55075 , n55076 , n55077 , n232839 , n232840 , n55080 , n55081 , n55082 , n55083 , n232845 , 
     n232846 , n55086 , n55087 , n55088 , n55089 , n232851 , n232852 , n55092 , n55093 , n55094 , 
     n55095 , n232857 , n232858 , n55098 , n55099 , n55100 , n55101 , n232863 , n232864 , n55104 , 
     n55105 , n55106 , n55107 , n55108 , n232870 , n232871 , n55111 , n55112 , n55113 , n55114 , 
     n232876 , n232877 , n55117 , n55118 , n55119 , n55120 , n55121 , n232883 , n232884 , n55124 , 
     n55125 , n232887 , n232888 , n55128 , n55129 , n55130 , n55131 , n232893 , n232894 , n55134 , 
     n55135 , n55136 , n55137 , n232899 , n232900 , n55140 , n55141 , n55142 , n55143 , n232905 , 
     n232906 , n55146 , n55147 , n55148 , n55149 , n232911 , n232912 , n55152 , n232914 , n232915 , 
     n55155 , n55156 , n55157 , n55158 , n55159 , n55160 , n232922 , n232923 , n55163 , n55164 , 
     n55165 , n55166 , n55167 , n232929 , n232930 , n55170 , n55171 , n55172 , n55173 , n232935 , 
     n232936 , n55176 , n55177 , n55178 , n55179 , n232941 , n232942 , n55182 , n55183 , n55184 , 
     n55185 , n232947 , n232948 , n55188 , n55189 , n55190 , n55191 , n232953 , n232954 , n55194 , 
     n232956 , n232957 , n55197 , n55198 , n55199 , n55200 , n232962 , n232963 , n55203 , n55204 , 
     n55205 , n55206 , n232968 , n232969 , n55209 , n232971 , n232972 , n55212 , n55213 , n55214 , 
     n55215 , n232977 , n232978 , n55218 , n55219 , n55220 , n55221 , n232983 , n232984 , n55224 , 
     n55225 , n55226 , n55227 , n232989 , n232990 , n55230 , n55231 , n55232 , n55233 , n232995 , 
     n232996 , n55236 , n232998 , n232999 , n55239 , n55240 , n55241 , n55242 , n55243 , n55244 , 
     n55245 , n55246 , n233008 , n233009 , n55249 , n55250 , n55251 , n55252 , n233014 , n233015 , 
     n55255 , n55256 , n55257 , n55258 , n233020 , n233021 , n55261 , n55262 , n55263 , n55264 , 
     n233026 , n233027 , n55267 , n55268 , n55269 , n55270 , n55271 , n55272 , n233034 , n233035 , 
     n55275 , n55276 , n55277 , n55278 , n233040 , n233041 , n55281 , n233043 , n233044 , n55284 , 
     n233046 , n233047 , n55287 , n55288 , n55289 , n55290 , n233052 , n233053 , n55293 , n55294 , 
     n55295 , n55296 , n233058 , n233059 , n55299 , n55300 , n55301 , n55302 , n55303 , n55304 , 
     n233066 , n233067 , n55307 , n55308 , n55309 , n55310 , n233072 , n233073 , n55313 , n55314 , 
     n55315 , n55316 , n233078 , n233079 , n55319 , n55320 , n55321 , n55322 , n233084 , n233085 , 
     n55325 , n55326 , n55327 , n55328 , n233090 , n233091 , n55331 , n55332 , n55333 , n55334 , 
     n233096 , n233097 , n55337 , n55338 , n55339 , n55340 , n233102 , n233103 , n55343 , n55344 , 
     n55345 , n55346 , n233108 , n233109 , n55349 , n55350 , n55351 , n55352 , n233114 , n233115 , 
     n55355 , n55356 , n55357 , n55358 , n233120 , n233121 , n55361 , n55362 , n55363 , n55364 , 
     n233126 , n233127 , n55367 , n55368 , n55369 , n55370 , n233132 , n233133 , n55373 , n55374 , 
     n55375 , n55376 , n233138 , n233139 , n55379 , n55380 , n55381 , n55382 , n233144 , n233145 , 
     n55385 , n55386 , n55387 , n55388 , n233150 , n233151 , n55391 , n55392 , n55393 , n55394 , 
     n233156 , n233157 , n55397 , n233159 , n233160 , n55400 , n55401 , n55402 , n55403 , n233165 , 
     n233166 , n55406 , n55407 , n55408 , n55409 , n55410 , n55411 , n55412 , n55413 , n55414 , 
     n55415 , n233177 , n233178 , n55418 , n55419 , n55420 , n55421 , n55422 , n55423 , n233185 , 
     n233186 , n55426 , n233188 , n233189 , n55429 , n233191 , n233192 , n55432 , n55433 , n55434 , 
     n55435 , n233197 , n233198 , n55438 , n55439 , n55440 , n55441 , n233203 , n233204 , n55444 , 
     n233206 , n233207 , n55447 , n55448 , n55449 , n55450 , n233212 , n233213 , n55453 , n55454 , 
     n55455 , n55456 , n233218 , n233219 , n55459 , n55460 , n55461 , n55462 , n233224 , n233225 , 
     n55465 , n55466 , n55467 , n55468 , n233230 , n233231 , n55471 , n233233 , n233234 , n55474 , 
     n55475 , n55476 , n55477 , n233239 , n233240 , n55480 , n55481 , n55482 , n55483 , n233245 , 
     n233246 , n55486 , n55487 , n55488 , n55489 , n233251 , n233252 , n55492 , n55493 , n55494 , 
     n55495 , n55496 , n233258 , n233259 , n55499 , n55500 , n55501 , n55502 , n233264 , n233265 , 
     n55505 , n55506 , n55507 , n55508 , n233270 , n233271 , n55511 , n55512 , n55513 , n55514 , 
     n233276 , n233277 , n55517 , n55518 , n55519 , n55520 , n233282 , n233283 , n55523 , n55524 , 
     n55525 , n55526 , n233288 , n233289 , n55529 , n55530 , n55531 , n55532 , n55533 , n55534 , 
     n233296 , n233297 , n55537 , n55538 , n233300 , n233301 , n55541 , n55542 , n55543 , n55544 , 
     n233306 , n233307 , n55547 , n55548 , n55549 , n55550 , n233312 , n233313 , n55553 , n233315 , 
     n233316 , n55556 , n233318 , n233319 , n55559 , n55560 , n55561 , n55562 , n233324 , n233325 , 
     n55565 , n55566 , n55567 , n55568 , n233330 , n233331 , n55571 , n55572 , n55573 , n55574 , 
     n233336 , n233337 , n55577 , n55578 , n55579 , n55580 , n233342 , n233343 , n55583 , n233345 , 
     n233346 , n55586 , n233348 , n233349 , n55589 , n55590 , n55591 , n55592 , n233354 , n233355 , 
     n55595 , n55596 , n55597 , n55598 , n233360 , n233361 , n55601 , n55602 , n55603 , n55604 , 
     n233366 , n233367 , n55607 , n233369 , n233370 , n55610 , n55611 , n55612 , n55613 , n233375 , 
     n233376 , n55616 , n233378 , n233379 , n55619 , n55620 , n55621 , n55622 , n55623 , n233385 , 
     n233386 , n55626 , n55627 , n55628 , n55629 , n55630 , n233392 , n233393 , n55633 , n55634 , 
     n55635 , n55636 , n233398 , n233399 , n55639 , n55640 , n55641 , n55642 , n233404 , n233405 , 
     n55645 , n55646 , n55647 , n55648 , n233410 , n233411 , n55651 , n55652 , n55653 , n55654 , 
     n233416 , n233417 , n55657 , n55658 , n55659 , n55660 , n233422 , n233423 , n55663 , n55664 , 
     n55665 , n55666 , n233428 , n233429 , n55669 , n233431 , n233432 , n55672 , n233434 , n233435 , 
     n55675 , n233437 , n55677 , n233439 , n233440 , n55680 , n55681 , n55682 , n55683 , n233445 , 
     n233446 , n55686 , n55687 , n55688 , n55689 , n233451 , n233452 , n55692 , n55693 , n55694 , 
     n55695 , n233457 , n233458 , n55698 , n55699 , n55700 , n55701 , n233463 , n233464 , n55704 , 
     n233466 , n233467 , n55707 , n233469 , n233470 , n55710 , n55711 , n55712 , n55713 , n55714 , 
     n233476 , n233477 , n55717 , n55718 , n55719 , n55720 , n55721 , n233483 , n233484 , n55724 , 
     n55725 , n55726 , n55727 , n233489 , n233490 , n55730 , n55731 , n55732 , n55733 , n233495 , 
     n233496 , n55736 , n55737 , n55738 , n55739 , n233501 , n233502 , n55742 , n55743 , n55744 , 
     n55745 , n233507 , n233508 , n55748 , n55749 , n55750 , n55751 , n233513 , n233514 , n233515 , 
     n233516 , n55756 , n233518 , n233519 , n55759 , n55760 , n55761 , n55762 , n55763 , n55764 , 
     n55765 , n55766 , n55767 , n55768 , n55769 , n55770 , n233532 , n233533 , n55773 , n55774 , 
     n55775 , n55776 , n233538 , n233539 , n55779 , n55780 , n55781 , n55782 , n55783 , n55784 , 
     n55785 , n55786 , n55787 , n233549 , n233550 , n233551 , n233552 , n55792 , n55793 , n55794 , 
     n55795 , n233557 , n233558 , n55798 , n55799 , n55800 , n55801 , n233563 , n233564 , n55804 , 
     n55805 , n55806 , n55807 , n233569 , n233570 , n55810 , n233572 , n233573 , n55813 , n55814 , 
     n55815 , n55816 , n233578 , n233579 , n55819 , n55820 , n55821 , n55822 , n233584 , n233585 , 
     n55825 , n55826 , n55827 , n55828 , n233590 , n233591 , n55831 , n55832 , n55833 , n55834 , 
     n55835 , n55836 , n55837 , n233599 , n233600 , n233601 , n233602 , n55842 , n55843 , n55844 , 
     n55845 , n233607 , n233608 , n55848 , n55849 , n55850 , n55851 , n233613 , n233614 , n55854 , 
     n55855 , n55856 , n55857 , n233619 , n233620 , n55860 , n55861 , n55862 , n55863 , n233625 , 
     n233626 , n55866 , n55867 , n55868 , n55869 , n233631 , n233632 , n55872 , n233634 , n233635 , 
     n233636 , n233637 , n55877 , n55878 , n233640 , n233641 , n55881 , n55882 , n55883 , n55884 , 
     n233646 , n233647 , n55887 , n55888 , n55889 , n55890 , n233652 , n233653 , n55893 , n55894 , 
     n55895 , n55896 , n55897 , n55898 , n233660 , n233661 , n233662 , n233663 , n55903 , n233665 , 
     n233666 , n55906 , n233668 , n233669 , n55909 , n55910 , n55911 , n55912 , n233674 , n233675 , 
     n55915 , n55916 , n55917 , n55918 , n233680 , n233681 , n55921 , n233683 , n55923 , n233685 , 
     n233686 , n55926 , n55927 , n55928 , n55929 , n233691 , n233692 , n55932 , n55933 , n55934 , 
     n55935 , n233697 , n233698 , n55938 , n55939 , n55940 , n55941 , n233703 , n233704 , n55944 , 
     n55945 , n55946 , n55947 , n233709 , n233710 , n55950 , n55951 , n55952 , n55953 , n233715 , 
     n233716 , n55956 , n55957 , n55958 , n55959 , n233721 , n233722 , n55962 , n55963 , n55964 , 
     n55965 , n233727 , n233728 , n55968 , n233730 , n233731 , n55971 , n55972 , n55973 , n55974 , 
     n233736 , n233737 , n55977 , n55978 , n55979 , n55980 , n233742 , n233743 , n55983 , n233745 , 
     n55985 , n55986 , n55987 , n55988 , n233750 , n233751 , n55991 , n55992 , n55993 , n55994 , 
     n233756 , n233757 , n55997 , n55998 , n55999 , n56000 , n233762 , n233763 , n56003 , n56004 , 
     n56005 , n56006 , n233768 , n233769 , n56009 , n56010 , n56011 , n56012 , n56013 , n56014 , 
     n233776 , n233777 , n56017 , n56018 , n56019 , n56020 , n56021 , n233783 , n233784 , n56024 , 
     n233786 , n233787 , n56027 , n56028 , n56029 , n56030 , n233792 , n233793 , n56033 , n56034 , 
     n56035 , n56036 , n233798 , n233799 , n56039 , n56040 , n56041 , n56042 , n233804 , n233805 , 
     n56045 , n56046 , n56047 , n56048 , n233810 , n233811 , n56051 , n233813 , n233814 , n56054 , 
     n233816 , n233817 , n56057 , n56058 , n56059 , n56060 , n233822 , n233823 , n56063 , n56064 , 
     n56065 , n56066 , n233828 , n233829 , n56069 , n56070 , n56071 , n56072 , n233834 , n233835 , 
     n56075 , n233837 , n233838 , n56078 , n233840 , n233841 , n233842 , n233843 , n233844 , n233845 , 
     n233846 , n233847 , n233848 , n233849 , n233850 , n233851 , n233852 , n233853 , n233854 , n233855 , 
     n233856 , n233857 , n233858 , n233859 , n233860 , n233861 , n233862 , n233863 , n233864 , n233865 , 
     n233866 , n233867 , n233868 , n233869 , n233870 , n233871 , n233872 , n233873 , n233874 , n233875 , 
     n233876 , n233877 , n233878 , n233879 , n233880 , n233881 , n233882 , n233883 , n233884 , n233885 , 
     n233886 , n233887 , n233888 , n233889 , n233890 , n233891 , n233892 , n233893 , n233894 , n233895 , 
     n233896 , n233897 , n233898 , n233899 , n233900 , n233901 , n233902 , n233903 , n233904 , n233905 , 
     n233906 , n233907 , n233908 , n233909 , n233910 , n233911 , n233912 , n233913 , n233914 , n233915 , 
     n233916 , n233917 , n233918 , n233919 , n233920 , n233921 , n233922 , n233923 , n233924 , n233925 , 
     n233926 , n233927 , n233928 , n233929 , n233930 , n233931 , n233932 , n233933 , n233934 , n233935 , 
     n233936 , n233937 , n233938 , n233939 , n233940 , n233941 , n233942 , n233943 , n233944 , n233945 , 
     n233946 , n233947 , n233948 , n233949 , n233950 , n233951 , n233952 , n233953 , n233954 , n233955 , 
     n233956 , n233957 , n233958 , n233959 , n233960 , n233961 , n233962 , n233963 , n233964 , n233965 , 
     n233966 , n233967 , n233968 , n233969 , n233970 , n233971 , n233972 , n233973 , n233974 , n233975 , 
     n233976 , n233977 , n233978 , n233979 , n233980 , n233981 , n233982 , n233983 , n233984 , n233985 , 
     n233986 , n233987 , n233988 , n233989 , n233990 , n233991 , n233992 , n233993 , n233994 , n233995 , 
     n233996 , n233997 , n233998 , n233999 , n234000 , n234001 , n234002 , n234003 , n234004 , n234005 , 
     n234006 , n234007 , n234008 , n234009 , n234010 , n234011 , n234012 , n234013 , n234014 , n234015 , 
     n234016 , n234017 , n234018 , n234019 , n234020 , n234021 , n234022 , n234023 , n234024 , n234025 , 
     n234026 , n234027 , n234028 , n234029 , n234030 , n234031 , n234032 , n234033 , n234034 , n234035 , 
     n234036 , n234037 , n234038 , n234039 , n234040 , n234041 , n234042 , n234043 , n234044 , n234045 , 
     n234046 , n234047 , n234048 , n234049 , n234050 , n234051 , n234052 , n234053 , n234054 , n234055 , 
     n234056 , n234057 , n234058 , n234059 , n234060 , n234061 , n234062 , n234063 , n234064 , n234065 , 
     n234066 , n234067 , n234068 , n234069 , n234070 , n234071 , n234072 , n234073 , n234074 , n234075 , 
     n234076 , n234077 , n234078 , n234079 , n234080 , n234081 , n234082 , n234083 , n234084 , n234085 , 
     n234086 , n234087 , n234088 , n234089 , n234090 , n234091 , n234092 , n234093 , n234094 , n234095 , 
     n234096 , n234097 , n234098 , n234099 , n234100 , n234101 , n234102 , n234103 , n234104 , n234105 , 
     n234106 , n234107 , n234108 , n234109 , n234110 , n234111 , n234112 , n234113 , n234114 , n234115 , 
     n234116 , n234117 , n234118 , n234119 , n234120 , n234121 , n234122 , n234123 , n234124 , n234125 , 
     n234126 , n234127 , n234128 , n234129 , n234130 , n234131 , n234132 , n234133 , n234134 , n234135 , 
     n234136 , n234137 , n234138 , n234139 , n234140 , n234141 , n234142 , n234143 , n234144 , n234145 , 
     n234146 , n234147 , n234148 , n234149 , n234150 , n234151 , n234152 , n234153 , n234154 , n234155 , 
     n234156 , n234157 , n234158 , n234159 , n234160 , n234161 , n234162 , n234163 , n234164 , n234165 , 
     n234166 , n234167 , n234168 , n234169 , n234170 , n234171 , n234172 , n234173 , n234174 , n234175 , 
     n234176 , n234177 , n234178 , n234179 , n234180 , n234181 , n234182 , n234183 , n234184 , n234185 , 
     n234186 , n234187 , n234188 , n234189 , n234190 , n234191 , n234192 , n234193 , n234194 , n234195 , 
     n234196 , n234197 , n234198 , n234199 , n234200 , n234201 , n234202 , n234203 , n234204 , n234205 , 
     n234206 , n234207 , n234208 , n234209 , n234210 , n234211 , n234212 , n234213 , n234214 , n234215 , 
     n234216 , n234217 , n234218 , n234219 , n234220 , n234221 , n234222 , n234223 , n234224 , n234225 , 
     n234226 , n234227 , n234228 , n234229 , n234230 , n234231 , n234232 , n234233 , n234234 , n234235 , 
     n234236 , n234237 , n234238 , n234239 , n234240 , n234241 , n234242 , n234243 , n234244 , n234245 , 
     n234246 , n234247 , n234248 , n234249 , n234250 , n234251 , n234252 , n234253 , n234254 , n234255 , 
     n234256 , n234257 , n234258 , n234259 , n234260 , n234261 , n234262 , n234263 , n234264 , n234265 , 
     n234266 , n234267 , n234268 , n234269 , n234270 , n234271 , n234272 , n234273 , n234274 , n234275 , 
     n234276 , n234277 , n234278 , n234279 , n234280 , n234281 , n234282 , n234283 , n234284 , n234285 , 
     n234286 , n234287 , n234288 , n234289 , n234290 , n234291 , n234292 , n234293 , n234294 , n234295 , 
     n234296 , n234297 , n234298 , n234299 , n234300 , n234301 , n234302 , n234303 , n234304 , n234305 , 
     n234306 , n234307 , n234308 , n234309 , n234310 , n234311 , n234312 , n234313 , n234314 , n234315 , 
     n234316 , n234317 , n234318 , n234319 , n234320 , n234321 , n234322 , n234323 , n234324 , n234325 , 
     n234326 , n234327 , n234328 , n234329 , n234330 , n234331 , n234332 , n234333 , n234334 , n234335 , 
     n234336 , n234337 , n234338 , n234339 , n234340 , n234341 , n234342 , n234343 , n234344 , n234345 , 
     n234346 , n234347 , n234348 , n234349 , n234350 , n234351 , n234352 , n234353 , n234354 , n234355 , 
     n234356 , n234357 , n234358 , n234359 , n234360 , n234361 , n234362 , n234363 , n234364 , n234365 , 
     n234366 , n234367 , n234368 , n234369 , n234370 , n234371 , n234372 , n234373 , n234374 , n234375 , 
     n234376 , n234377 , n234378 , n234379 , n234380 , n234381 , n234382 , n234383 , n234384 , n234385 , 
     n234386 , n234387 , n234388 , n234389 , n234390 , n234391 , n234392 , n234393 , n234394 , n234395 , 
     n234396 , n234397 , n234398 , n234399 , n234400 , n234401 , n234402 , n234403 , n234404 , n234405 , 
     n234406 , n234407 , n234408 , n234409 , n234410 , n234411 , n234412 , n234413 , n234414 , n234415 , 
     n234416 , n234417 , n234418 , n234419 , n234420 , n234421 , n234422 , n234423 , n234424 , n234425 , 
     n234426 , n234427 , n234428 , n234429 , n234430 , n234431 , n234432 , n234433 , n234434 , n234435 , 
     n234436 , n234437 , n234438 , n234439 , n234440 , n234441 , n234442 , n234443 , n234444 , n234445 , 
     n234446 , n234447 , n234448 , n234449 , n234450 , n234451 , n234452 , n234453 , n234454 , n234455 , 
     n234456 , n234457 , n234458 , n234459 , n234460 , n234461 , n234462 , n234463 , n234464 , n234465 , 
     n234466 , n234467 , n234468 , n234469 , n234470 , n234471 , n234472 , n234473 , n234474 , n234475 , 
     n234476 , n234477 , n234478 , n234479 , n234480 , n234481 , n234482 , n234483 , n234484 , n234485 , 
     n234486 , n234487 , n234488 , n234489 , n234490 , n234491 , n234492 , n234493 , n234494 , n234495 , 
     n234496 , n234497 , n234498 , n234499 , n234500 , n234501 , n234502 , n234503 , n234504 , n234505 , 
     n234506 , n234507 , n234508 , n234509 , n234510 , n234511 , n234512 , n234513 , n234514 , n234515 , 
     n234516 , n234517 , n234518 , n234519 , n234520 , n234521 , n234522 , n234523 , n234524 , n234525 , 
     n234526 , n234527 , n234528 , n234529 , n234530 , n234531 , n234532 , n234533 , n234534 , n234535 , 
     n234536 , n234537 , n234538 , n234539 , n234540 , n234541 , n234542 , n234543 , n234544 , n234545 , 
     n234546 , n234547 , n234548 , n234549 , n234550 , n234551 , n234552 , n234553 , n234554 , n234555 , 
     n234556 , n234557 , n234558 , n234559 , n234560 , n234561 , n234562 , n234563 , n234564 , n234565 , 
     n234566 , n234567 , n234568 , n234569 , n234570 , n234571 , n234572 , n234573 , n234574 , n234575 , 
     n234576 , n234577 , n234578 , n234579 , n234580 , n234581 , n234582 , n234583 , n234584 , n234585 , 
     n234586 , n234587 , n234588 , n234589 , n234590 , n234591 , n234592 , n234593 , n234594 , n234595 , 
     n234596 , n234597 , n234598 , n234599 , n234600 , n234601 , n234602 , n234603 , n234604 , n234605 , 
     n234606 , n234607 , n234608 , n234609 , n234610 , n234611 , n234612 , n234613 , n234614 , n234615 , 
     n234616 , n234617 , n234618 , n234619 , n234620 , n234621 , n234622 , n234623 , n234624 , n234625 , 
     n234626 , n234627 , n234628 , n234629 , n234630 , n234631 , n234632 , n234633 , n234634 , n234635 , 
     n234636 , n234637 , n234638 , n234639 , n234640 , n234641 , n234642 , n234643 , n234644 , n234645 , 
     n234646 , n234647 , n234648 , n234649 , n234650 , n234651 , n234652 , n234653 , n234654 , n234655 , 
     n234656 , n234657 , n234658 , n234659 , n234660 , n234661 , n234662 , n234663 , n234664 , n234665 , 
     n234666 , n234667 , n234668 , n234669 , n234670 , n234671 , n234672 , n234673 , n234674 , n234675 , 
     n234676 , n234677 , n234678 , n234679 , n234680 , n234681 , n234682 , n234683 , n234684 , n234685 , 
     n234686 , n234687 , n234688 , n234689 , n234690 , n234691 , n234692 , n234693 , n234694 , n234695 , 
     n234696 , n234697 , n234698 , n234699 , n234700 , n234701 , n234702 , n234703 , n234704 , n234705 , 
     n234706 , n234707 , n234708 , n234709 , n234710 , n234711 , n234712 , n234713 , n234714 , n234715 , 
     n234716 , n234717 , n234718 , n234719 , n234720 , n234721 , n234722 , n234723 , n234724 , n234725 , 
     n234726 , n234727 , n234728 , n234729 , n234730 , n234731 , n234732 , n234733 , n234734 , n234735 , 
     n234736 , n234737 , n234738 , n234739 , n234740 , n234741 , n234742 , n234743 , n234744 , n234745 , 
     n234746 , n234747 , n234748 , n234749 , n234750 , n234751 , n234752 , n234753 , n234754 , n234755 , 
     n234756 , n234757 , n234758 , n234759 , n234760 , n234761 , n234762 , n234763 , n234764 , n234765 , 
     n234766 , n234767 , n234768 , n234769 , n234770 , n234771 , n234772 , n234773 , n234774 , n234775 , 
     n234776 , n234777 , n234778 , n234779 , n234780 , n234781 , n234782 , n234783 , n234784 , n234785 , 
     n234786 , n234787 , n234788 , n234789 , n234790 , n234791 , n234792 , n234793 , n234794 , n234795 , 
     n234796 , n234797 , n234798 , n234799 , n234800 , n234801 , n234802 , n234803 , n234804 , n234805 , 
     n234806 , n234807 , n234808 , n234809 , n234810 , n234811 , n234812 , n234813 , n234814 , n234815 , 
     n234816 , n234817 , n234818 , n234819 , n234820 , n234821 , n234822 , n234823 , n234824 , n234825 , 
     n234826 , n234827 , n234828 , n234829 , n234830 , n234831 , n234832 , n234833 , n234834 , n234835 , 
     n234836 , n234837 , n234838 , n234839 , n234840 , n234841 , n234842 , n234843 , n234844 , n234845 , 
     n234846 , n234847 , n234848 , n234849 , n234850 , n234851 , n234852 , n234853 , n234854 , n234855 , 
     n234856 , n234857 , n234858 , n234859 , n234860 , n234861 , n234862 , n234863 , n234864 , n234865 , 
     n234866 , n234867 , n234868 , n234869 , n234870 , n234871 , n234872 , n234873 , n234874 , n234875 , 
     n234876 , n234877 , n234878 , n234879 , n234880 , n234881 , n234882 , n234883 , n234884 , n234885 , 
     n234886 , n234887 , n234888 , n234889 , n234890 , n234891 , n234892 , n234893 , n234894 , n234895 , 
     n234896 , n234897 , n234898 , n234899 , n234900 , n234901 , n234902 , n234903 , n234904 , n234905 , 
     n234906 , n234907 , n234908 , n234909 , n234910 , n234911 , n234912 , n234913 , n234914 , n234915 , 
     n234916 , n234917 , n234918 , n234919 , n234920 , n234921 , n234922 , n234923 , n234924 , n234925 , 
     n234926 , n234927 , n234928 , n234929 , n234930 , n234931 , n234932 , n234933 , n234934 , n234935 , 
     n234936 , n234937 , n234938 , n234939 , n234940 , n234941 , n234942 , n234943 , n234944 , n234945 , 
     n234946 , n234947 , n234948 , n234949 , n234950 , n234951 , n234952 , n234953 , n234954 , n234955 , 
     n234956 , n234957 , n234958 , n234959 , n234960 , n234961 , n234962 , n234963 , n234964 , n234965 , 
     n234966 , n234967 , n234968 , n234969 , n234970 , n234971 , n234972 , n234973 , n234974 , n234975 , 
     n234976 , n234977 , n234978 , n234979 , n234980 , n234981 , n234982 , n234983 , n234984 , n234985 , 
     n234986 , n234987 , n234988 , n234989 , n234990 , n234991 , n234992 , n234993 , n234994 , n234995 , 
     n234996 , n234997 , n234998 , n234999 , n235000 , n235001 , n235002 , n235003 , n235004 , n235005 , 
     n235006 , n235007 , n235008 , n235009 , n235010 , n235011 , n235012 , n235013 , n235014 , n235015 , 
     n235016 , n235017 , n235018 , n235019 , n235020 , n235021 , n235022 , n235023 , n235024 , n235025 , 
     n235026 , n235027 , n235028 , n235029 , n235030 , n235031 , n235032 , n235033 , n235034 , n235035 , 
     n235036 , n235037 , n235038 , n235039 , n235040 , n235041 , n235042 , n235043 , n235044 , n235045 , 
     n235046 , n235047 , n235048 , n235049 , n235050 , n235051 , n235052 , n235053 , n235054 , n235055 , 
     n235056 , n235057 , n235058 , n235059 , n235060 , n235061 , n235062 , n235063 , n235064 , n235065 , 
     n235066 , n235067 , n235068 , n235069 , n235070 , n235071 , n235072 , n235073 , n235074 , n235075 , 
     n235076 , n235077 , n235078 , n235079 , n235080 , n235081 , n235082 , n235083 , n235084 , n235085 , 
     n235086 , n235087 , n235088 , n235089 , n235090 , n235091 , n235092 , n235093 , n235094 , n235095 , 
     n235096 , n235097 , n235098 , n235099 , n235100 , n235101 , n235102 , n235103 , n235104 , n235105 , 
     n235106 , n235107 , n235108 , n235109 , n235110 , n235111 , n235112 , n235113 , n235114 , n235115 , 
     n235116 , n235117 , n235118 , n235119 , n235120 , n235121 , n235122 , n235123 , n235124 , n235125 , 
     n235126 , n235127 , n235128 , n235129 , n235130 , n235131 , n235132 , n235133 , n235134 , n235135 , 
     n235136 , n235137 , n235138 , n235139 , n235140 , n235141 , n235142 , n235143 , n235144 , n235145 , 
     n235146 , n235147 , n235148 , n235149 , n235150 , n235151 , n235152 , n235153 , n235154 , n235155 , 
     n235156 , n235157 , n235158 , n235159 , n235160 , n235161 , n235162 , n235163 , n235164 , n235165 , 
     n235166 , n235167 , n235168 , n235169 , n235170 , n235171 , n235172 , n235173 , n235174 , n235175 , 
     n235176 , n235177 , n235178 , n235179 , n235180 , n235181 , n235182 , n235183 , n235184 , n235185 , 
     n235186 , n235187 , n235188 , n235189 , n235190 , n235191 , n235192 , n235193 , n235194 , n235195 , 
     n235196 , n235197 , n235198 , n235199 , n235200 , n235201 , n235202 , n235203 , n235204 , n235205 , 
     n235206 , n235207 , n235208 , n235209 , n235210 , n235211 , n235212 , n235213 , n235214 , n235215 , 
     n235216 , n235217 , n235218 , n235219 , n235220 , n235221 , n235222 , n235223 , n235224 , n235225 , 
     n235226 , n235227 , n235228 , n235229 , n235230 , n235231 , n235232 , n235233 , n235234 , n235235 , 
     n235236 , n235237 , n235238 , n235239 , n235240 , n235241 , n235242 , n235243 , n235244 , n235245 , 
     n235246 , n235247 , n235248 , n235249 , n235250 , n235251 , n235252 , n235253 , n235254 , n235255 , 
     n235256 , n235257 , n235258 , n235259 , n235260 , n235261 , n235262 , n235263 , n235264 , n235265 , 
     n235266 , n235267 , n235268 , n235269 , n235270 , n235271 , n235272 , n235273 , n235274 , n235275 , 
     n235276 , n235277 , n235278 , n235279 , n235280 , n235281 , n235282 , n235283 , n235284 , n235285 , 
     n235286 , n235287 , n235288 , n235289 , n235290 , n235291 , n235292 , n235293 , n235294 , n235295 , 
     n235296 , n235297 , n235298 , n235299 , n235300 , n235301 , n235302 , n235303 , n235304 , n235305 , 
     n235306 , n235307 , n235308 , n235309 , n235310 , n235311 , n235312 , n235313 , n235314 , n235315 , 
     n235316 , n235317 , n235318 , n235319 , n235320 , n235321 , n235322 , n235323 , n235324 , n235325 , 
     n235326 , n235327 , n235328 , n235329 , n235330 , n235331 , n235332 , n235333 , n235334 , n235335 , 
     n235336 , n235337 , n235338 , n235339 , n235340 , n235341 , n235342 , n235343 , n235344 , n235345 , 
     n235346 , n235347 , n235348 , n235349 , n235350 , n235351 , n235352 , n235353 , n235354 , n235355 , 
     n235356 , n235357 , n235358 , n235359 , n235360 , n235361 , n235362 , n235363 , n235364 , n235365 , 
     n235366 , n235367 , n235368 , n235369 , n235370 , n235371 , n235372 , n235373 , n235374 , n235375 , 
     n235376 , n235377 , n235378 , n235379 , n235380 , n235381 , n235382 , n235383 , n235384 , n235385 , 
     n235386 , n235387 , n235388 , n235389 , n235390 , n235391 , n235392 , n235393 , n235394 , n235395 , 
     n235396 , n235397 , n235398 , n235399 , n235400 , n235401 , n235402 , n235403 , n235404 , n235405 , 
     n235406 , n235407 , n235408 , n235409 , n235410 , n235411 , n235412 , n235413 , n235414 , n235415 , 
     n235416 , n235417 , n235418 , n235419 , n235420 , n235421 , n235422 , n235423 , n235424 , n235425 , 
     n235426 , n235427 , n235428 , n235429 , n235430 , n235431 , n235432 , n235433 , n235434 , n235435 , 
     n235436 , n235437 , n235438 , n235439 , n235440 , n235441 , n235442 , n235443 , n235444 , n235445 , 
     n235446 , n235447 , n235448 , n235449 , n235450 , n235451 , n235452 , n235453 , n235454 , n235455 , 
     n235456 , n235457 , n235458 , n235459 , n235460 , n235461 , n235462 , n235463 , n235464 , n235465 , 
     n235466 , n235467 , n235468 , n235469 , n235470 , n235471 , n235472 , n235473 , n235474 , n235475 , 
     n235476 , n235477 , n235478 , n235479 , n235480 , n235481 , n235482 , n235483 , n235484 , n235485 , 
     n235486 , n235487 , n235488 , n235489 , n235490 , n235491 , n235492 , n235493 , n235494 , n235495 , 
     n235496 , n235497 , n235498 , n235499 , n235500 , n235501 , n235502 , n235503 , n235504 , n235505 , 
     n235506 , n235507 , n235508 , n235509 , n235510 , n235511 , n235512 , n235513 , n235514 , n235515 , 
     n235516 , n235517 , n235518 , n235519 , n235520 , n235521 , n235522 , n235523 , n235524 , n235525 , 
     n235526 , n235527 , n235528 , n235529 , n235530 , n235531 , n235532 , n235533 , n235534 , n235535 , 
     n235536 , n235537 , n235538 , n235539 , n235540 , n235541 , n235542 , n235543 , n235544 , n235545 , 
     n235546 , n235547 , n235548 , n235549 , n235550 , n235551 , n235552 , n235553 , n235554 , n235555 , 
     n235556 , n235557 , n235558 , n235559 , n235560 , n235561 , n235562 , n235563 , n235564 , n235565 , 
     n235566 , n235567 , n235568 , n235569 , n235570 , n235571 , n235572 , n235573 , n235574 , n235575 , 
     n235576 , n235577 , n235578 , n235579 , n235580 , n235581 , n235582 , n235583 , n235584 , n235585 , 
     n235586 , n235587 , n235588 , n235589 , n235590 , n235591 , n235592 , n235593 , n235594 , n235595 , 
     n235596 , n235597 , n235598 , n235599 , n235600 , n235601 , n235602 , n235603 , n235604 , n235605 , 
     n235606 , n235607 , n235608 , n235609 , n235610 , n235611 , n235612 , n235613 , n235614 , n235615 , 
     n235616 , n235617 , n235618 , n235619 , n235620 , n235621 , n235622 , n235623 , n235624 , n235625 , 
     n235626 , n235627 , n235628 , n235629 , n235630 , n235631 , n235632 , n235633 , n235634 , n235635 , 
     n235636 , n235637 , n235638 , n235639 , n235640 , n235641 , n235642 , n235643 , n235644 , n235645 , 
     n235646 , n235647 , n235648 , n235649 , n235650 , n235651 , n235652 , n235653 , n235654 , n235655 , 
     n235656 , n235657 , n235658 , n235659 , n235660 , n235661 , n235662 , n235663 , n235664 , n235665 , 
     n235666 , n235667 , n235668 , n235669 , n235670 , n235671 , n235672 , n235673 , n235674 , n235675 , 
     n235676 , n235677 , n235678 , n235679 , n235680 , n235681 , n235682 , n235683 , n235684 , n235685 , 
     n235686 , n235687 , n235688 , n235689 , n235690 , n235691 , n235692 , n235693 , n235694 , n235695 , 
     n235696 , n235697 , n235698 , n235699 , n235700 , n235701 , n235702 , n235703 , n235704 , n235705 , 
     n235706 , n235707 , n235708 , n235709 , n235710 , n235711 , n235712 , n235713 , n235714 , n235715 , 
     n235716 , n235717 , n235718 , n235719 , n235720 , n235721 , n235722 , n235723 , n235724 , n235725 , 
     n235726 , n235727 , n235728 , n235729 , n235730 , n235731 , n235732 , n235733 , n235734 , n235735 , 
     n235736 , n235737 , n235738 , n235739 , n235740 , n235741 , n235742 , n235743 , n235744 , n235745 , 
     n235746 , n235747 , n235748 , n235749 , n235750 , n235751 , n235752 , n235753 , n235754 , n235755 , 
     n235756 , n235757 , n235758 , n235759 , n235760 , n235761 , n235762 , n235763 , n235764 , n235765 , 
     n235766 , n235767 , n235768 , n235769 , n235770 , n235771 , n235772 , n235773 , n235774 , n235775 , 
     n235776 , n235777 , n235778 , n235779 , n235780 , n235781 , n235782 , n235783 , n235784 , n235785 , 
     n235786 , n235787 , n235788 , n235789 , n235790 , n235791 , n235792 , n235793 , n235794 , n235795 , 
     n235796 , n235797 , n235798 , n235799 , n235800 , n235801 , n235802 , n235803 , n235804 , n235805 , 
     n235806 , n235807 , n235808 , n235809 , n235810 , n235811 , n235812 , n235813 , n235814 , n235815 , 
     n235816 , n235817 , n235818 , n235819 , n235820 , n235821 , n235822 , n235823 , n235824 , n235825 , 
     n235826 , n235827 , n235828 , n235829 , n235830 , n235831 , n235832 , n235833 , n235834 , n235835 , 
     n235836 , n235837 , n235838 , n235839 , n235840 , n235841 , n235842 , n235843 , n235844 , n235845 , 
     n235846 , n235847 , n235848 , n235849 , n235850 , n235851 , n235852 , n235853 , n235854 , n235855 , 
     n235856 , n235857 , n235858 , n235859 , n235860 , n235861 , n235862 , n235863 , n235864 , n235865 , 
     n235866 , n235867 , n235868 , n235869 , n235870 , n235871 , n235872 , n235873 , n235874 , n235875 , 
     n235876 , n235877 , n235878 , n235879 , n235880 , n235881 , n235882 , n235883 , n235884 , n235885 , 
     n235886 , n235887 , n235888 , n235889 , n235890 , n235891 , n235892 , n235893 , n235894 , n235895 , 
     n235896 , n235897 , n235898 , n235899 , n235900 , n235901 , n235902 , n235903 , n235904 , n235905 , 
     n235906 , n235907 , n235908 , n235909 , n235910 , n235911 , n235912 , n235913 , n235914 , n235915 , 
     n235916 , n235917 , n235918 , n235919 , n235920 , n235921 , n235922 , n235923 , n235924 , n235925 , 
     n235926 , n235927 , n235928 , n235929 , n235930 , n235931 , n235932 , n235933 , n235934 , n235935 , 
     n235936 , n235937 , n235938 , n235939 , n235940 , n235941 , n235942 , n235943 , n235944 , n235945 , 
     n235946 , n235947 , n235948 , n235949 , n235950 , n235951 , n235952 , n235953 , n235954 , n235955 , 
     n235956 , n235957 , n235958 , n235959 , n235960 , n235961 , n235962 , n235963 , n235964 , n235965 , 
     n235966 , n235967 , n235968 , n235969 , n235970 , n235971 , n235972 , n235973 , n235974 , n235975 , 
     n235976 , n235977 , n235978 , n235979 , n235980 , n235981 , n235982 , n235983 , n235984 , n235985 , 
     n235986 , n235987 , n235988 , n235989 , n235990 , n235991 , n235992 , n235993 , n235994 , n235995 , 
     n235996 , n235997 , n235998 , n235999 , n236000 , n236001 , n236002 , n236003 , n236004 , n236005 , 
     n236006 , n236007 , n236008 , n236009 , n236010 , n236011 , n236012 , n236013 , n236014 , n236015 , 
     n236016 , n236017 , n236018 , n236019 , n236020 , n236021 , n236022 , n236023 , n236024 , n236025 , 
     n236026 , n236027 , n236028 , n236029 , n236030 , n236031 , n236032 , n236033 , n236034 , n236035 , 
     n236036 , n236037 , n236038 , n236039 , n236040 , n236041 , n236042 , n236043 , n236044 , n236045 , 
     n236046 , n236047 , n236048 , n236049 , n236050 , n236051 , n236052 , n236053 , n236054 , n236055 , 
     n236056 , n236057 , n236058 , n236059 , n236060 , n236061 , n236062 , n236063 , n236064 , n236065 , 
     n236066 , n236067 , n236068 , n236069 , n236070 , n236071 , n236072 , n236073 , n236074 , n236075 , 
     n236076 , n236077 , n236078 , n236079 , n236080 , n236081 , n236082 , n236083 , n236084 , n236085 , 
     n236086 , n236087 , n236088 , n236089 , n236090 , n236091 , n236092 , n236093 , n236094 , n236095 , 
     n236096 , n236097 , n236098 , n236099 , n236100 , n236101 , n236102 , n236103 , n236104 , n236105 , 
     n236106 , n236107 , n236108 , n236109 , n236110 , n236111 , n236112 , n236113 , n236114 , n236115 , 
     n236116 , n236117 , n236118 , n236119 , n236120 , n236121 , n236122 , n236123 , n236124 , n236125 , 
     n236126 , n236127 , n236128 , n236129 , n236130 , n236131 , n236132 , n236133 , n236134 , n236135 , 
     n236136 , n236137 , n236138 , n236139 , n236140 , n236141 , n236142 , n236143 , n236144 , n236145 , 
     n236146 , n236147 , n236148 , n236149 , n236150 , n236151 , n236152 , n236153 , n236154 , n236155 , 
     n236156 , n236157 , n236158 , n236159 , n236160 , n236161 , n236162 , n236163 , n236164 , n236165 , 
     n236166 , n236167 , n236168 , n236169 , n236170 , n236171 , n236172 , n236173 , n236174 , n236175 , 
     n236176 , n236177 , n236178 , n236179 , n236180 , n236181 , n236182 , n236183 , n236184 , n236185 , 
     n236186 , n236187 , n236188 , n236189 , n236190 , n236191 , n236192 , n236193 , n236194 , n236195 , 
     n236196 , n236197 , n236198 , n236199 , n236200 , n236201 , n236202 , n236203 , n236204 , n236205 , 
     n236206 , n236207 , n236208 , n236209 , n236210 , n236211 , n236212 , n236213 , n236214 , n236215 , 
     n236216 , n236217 , n236218 , n236219 , n236220 , n236221 , n236222 , n236223 , n236224 , n236225 , 
     n236226 , n236227 , n236228 , n236229 , n236230 , n236231 , n236232 , n236233 , n236234 , n236235 , 
     n236236 , n236237 , n236238 , n236239 , n236240 , n236241 , n236242 , n236243 , n236244 , n236245 , 
     n236246 , n236247 , n236248 , n236249 , n236250 , n236251 , n236252 , n236253 , n236254 , n236255 , 
     n236256 , n236257 , n236258 , n236259 , n236260 , n236261 , n236262 , n236263 , n236264 , n236265 , 
     n236266 , n236267 , n236268 , n236269 , n236270 , n236271 , n236272 , n236273 , n236274 , n236275 , 
     n236276 , n236277 , n236278 , n236279 , n236280 , n236281 , n236282 , n236283 , n236284 , n236285 , 
     n236286 , n236287 , n236288 , n236289 , n236290 , n236291 , n236292 , n236293 , n236294 , n236295 , 
     n236296 , n236297 , n236298 , n236299 , n236300 , n236301 , n236302 , n236303 , n236304 , n236305 , 
     n236306 , n236307 , n236308 , n236309 , n236310 , n236311 , n236312 , n236313 , n236314 , n236315 , 
     n236316 , n236317 , n236318 , n236319 , n236320 , n236321 , n236322 , n236323 , n236324 , n236325 , 
     n236326 , n236327 , n236328 , n236329 , n236330 , n236331 , n236332 , n236333 , n236334 , n236335 , 
     n236336 , n236337 , n236338 , n236339 , n236340 , n236341 , n236342 , n236343 , n236344 , n236345 , 
     n236346 , n236347 , n236348 , n236349 , n236350 , n236351 , n236352 , n236353 , n236354 , n236355 , 
     n236356 , n236357 , n236358 , n236359 , n236360 , n236361 , n236362 , n236363 , n236364 , n236365 , 
     n236366 , n236367 , n236368 , n236369 , n236370 , n236371 , n236372 , n236373 , n236374 , n236375 , 
     n236376 , n236377 , n236378 , n236379 , n236380 , n236381 , n236382 , n236383 , n236384 , n236385 , 
     n236386 , n236387 , n236388 , n236389 , n236390 , n236391 , n236392 , n236393 , n236394 , n236395 , 
     n236396 , n236397 , n236398 , n236399 , n236400 , n236401 , n236402 , n236403 , n236404 , n236405 , 
     n236406 , n236407 , n236408 , n236409 , n236410 , n236411 , n236412 , n236413 , n236414 , n236415 , 
     n236416 , n236417 , n236418 , n236419 , n236420 , n236421 , n236422 , n236423 , n236424 , n236425 , 
     n236426 , n236427 , n236428 , n236429 , n236430 , n236431 , n236432 , n236433 , n236434 , n236435 , 
     n236436 , n236437 , n236438 , n236439 , n236440 , n236441 , n236442 , n236443 , n236444 , n236445 , 
     n236446 , n236447 , n236448 , n236449 , n236450 , n236451 , n236452 , n236453 , n236454 , n236455 , 
     n236456 , n236457 , n236458 , n236459 , n236460 , n236461 , n236462 , n236463 , n236464 , n236465 , 
     n236466 , n236467 , n236468 , n236469 , n236470 , n236471 , n236472 , n236473 , n236474 , n236475 , 
     n236476 , n236477 , n236478 , n236479 , n236480 , n236481 , n236482 , n236483 , n236484 , n236485 , 
     n236486 , n236487 , n236488 , n236489 , n236490 , n236491 , n236492 , n236493 , n236494 , n236495 , 
     n236496 , n236497 , n236498 , n236499 , n236500 , n236501 , n236502 , n236503 , n236504 , n236505 , 
     n236506 , n236507 , n236508 , n236509 , n236510 , n236511 , n236512 , n236513 , n236514 , n236515 , 
     n236516 , n236517 , n236518 , n236519 , n236520 , n236521 , n236522 , n236523 , n236524 , n236525 , 
     n236526 , n236527 , n236528 , n236529 , n236530 , n236531 , n236532 , n236533 , n236534 , n236535 , 
     n236536 , n236537 , n236538 , n236539 , n236540 , n236541 , n236542 , n236543 , n236544 , n236545 , 
     n236546 , n236547 , n236548 , n236549 , n236550 , n236551 , n236552 , n236553 , n236554 , n236555 , 
     n236556 , n236557 , n236558 , n236559 , n236560 , n236561 , n236562 , n236563 , n236564 , n236565 , 
     n236566 , n236567 , n236568 , n236569 , n236570 , n236571 , n236572 , n236573 , n236574 , n236575 , 
     n236576 , n236577 , n236578 , n236579 , n236580 , n236581 , n236582 , n236583 , n236584 , n236585 , 
     n236586 , n236587 , n236588 , n236589 , n236590 , n236591 , n236592 , n236593 , n236594 , n236595 , 
     n236596 , n236597 , n236598 , n236599 , n236600 , n236601 , n236602 , n236603 , n236604 , n236605 , 
     n236606 , n236607 , n236608 , n236609 , n236610 , n236611 , n236612 , n236613 , n236614 , n236615 , 
     n236616 , n236617 , n236618 , n236619 , n236620 , n236621 , n236622 , n236623 , n236624 , n236625 , 
     n236626 , n236627 , n236628 , n236629 , n236630 , n236631 , n236632 , n236633 , n236634 , n236635 , 
     n236636 , n236637 , n236638 , n236639 , n236640 , n236641 , n236642 , n236643 , n236644 , n236645 , 
     n236646 , n236647 , n236648 , n236649 , n236650 , n236651 , n236652 , n236653 , n236654 , n236655 , 
     n236656 , n236657 , n236658 , n236659 , n236660 , n236661 , n236662 , n236663 , n236664 , n236665 , 
     n236666 , n236667 , n236668 , n236669 , n236670 , n236671 , n236672 , n236673 , n236674 , n236675 , 
     n236676 , n236677 , n236678 , n236679 , n236680 , n236681 , n236682 , n236683 , n236684 , n236685 , 
     n236686 , n236687 , n236688 , n236689 , n236690 , n236691 , n236692 , n236693 , n236694 , n236695 , 
     n236696 , n236697 , n236698 , n236699 , n236700 , n236701 , n236702 , n236703 , n236704 , n236705 , 
     n236706 , n236707 , n236708 , n236709 , n236710 , n236711 , n236712 , n236713 , n236714 , n236715 , 
     n236716 , n236717 , n236718 , n236719 , n236720 , n236721 , n236722 , n236723 , n236724 , n236725 , 
     n236726 , n236727 , n236728 , n236729 , n236730 , n236731 , n236732 , n236733 , n236734 , n236735 , 
     n236736 , n236737 , n236738 , n236739 , n236740 , n236741 , n236742 , n236743 , n236744 , n236745 , 
     n236746 , n236747 , n236748 , n236749 , n236750 , n236751 , n236752 , n236753 , n236754 , n236755 , 
     n236756 , n236757 , n236758 , n236759 , n236760 , n236761 , n236762 , n236763 , n236764 , n236765 , 
     n236766 , n236767 , n236768 , n236769 , n236770 , n236771 , n236772 , n236773 , n236774 , n236775 , 
     n236776 , n236777 , n236778 , n236779 , n236780 , n236781 , n236782 , n236783 , n236784 , n236785 , 
     n236786 , n236787 , n236788 , n236789 , n236790 , n236791 , n236792 , n236793 , n236794 , n236795 , 
     n236796 , n236797 , n236798 , n236799 , n236800 , n236801 , n236802 , n236803 , n236804 , n236805 , 
     n236806 , n236807 , n236808 , n236809 , n236810 , n236811 , n236812 , n236813 , n236814 , n236815 , 
     n236816 , n236817 , n236818 , n236819 , n236820 , n236821 , n236822 , n236823 , n236824 , n236825 , 
     n236826 , n236827 , n236828 , n236829 , n236830 , n236831 , n236832 , n236833 , n236834 , n236835 , 
     n236836 , n236837 , n236838 , n236839 , n236840 , n236841 , n236842 , n236843 , n236844 , n236845 , 
     n236846 , n236847 , n236848 , n236849 , n236850 , n236851 , n236852 , n236853 , n236854 , n236855 , 
     n236856 , n236857 , n236858 , n236859 , n236860 , n236861 , n236862 , n236863 , n236864 , n236865 , 
     n236866 , n236867 , n236868 , n236869 , n236870 , n236871 , n236872 , n236873 , n236874 , n236875 , 
     n236876 , n236877 , n236878 , n236879 , n236880 , n236881 , n236882 , n236883 , n236884 , n236885 , 
     n236886 , n236887 , n236888 , n236889 , n236890 , n236891 , n236892 , n236893 , n236894 , n236895 , 
     n236896 , n236897 , n236898 , n236899 , n236900 , n236901 , n236902 , n236903 , n236904 , n236905 , 
     n236906 , n236907 , n236908 , n236909 , n236910 , n236911 , n236912 , n236913 , n236914 , n236915 , 
     n236916 , n236917 , n236918 , n236919 , n236920 , n236921 , n236922 , n236923 , n236924 , n236925 , 
     n236926 , n236927 , n236928 , n236929 , n236930 , n236931 , n236932 , n236933 , n236934 , n236935 , 
     n236936 , n236937 , n236938 , n236939 , n236940 , n236941 , n236942 , n236943 , n236944 , n236945 , 
     n236946 , n236947 , n236948 , n236949 , n236950 , n236951 , n236952 , n236953 , n236954 , n236955 , 
     n236956 , n236957 , n236958 , n236959 , n236960 , n236961 , n236962 , n236963 , n236964 , n236965 , 
     n236966 , n236967 , n236968 , n236969 , n236970 , n236971 , n236972 , n236973 , n236974 , n236975 , 
     n236976 , n236977 , n236978 , n236979 , n236980 , n236981 , n236982 , n236983 , n236984 , n236985 , 
     n236986 , n236987 , n236988 , n236989 , n236990 , n236991 , n236992 , n236993 , n236994 , n236995 , 
     n236996 , n236997 , n236998 , n236999 , n237000 , n237001 , n237002 , n237003 , n237004 , n237005 , 
     n237006 , n237007 , n237008 , n237009 , n237010 , n237011 , n237012 , n237013 , n237014 , n237015 , 
     n237016 , n237017 , n237018 , n237019 , n237020 , n237021 , n237022 , n237023 , n237024 , n237025 , 
     n237026 , n237027 , n237028 , n237029 , n237030 , n237031 , n237032 , n237033 , n237034 , n237035 , 
     n237036 , n237037 , n237038 , n237039 , n237040 , n237041 , n237042 , n237043 , n237044 , n237045 , 
     n237046 , n237047 , n237048 , n237049 , n237050 , n237051 , n237052 , n237053 , n237054 , n237055 , 
     n237056 , n237057 , n237058 , n237059 , n237060 , n237061 , n237062 , n237063 , n237064 , n237065 , 
     n237066 , n237067 , n237068 , n237069 , n237070 , n237071 , n237072 , n237073 , n237074 , n237075 , 
     n237076 , n237077 , n237078 , n237079 , n237080 , n237081 , n237082 , n237083 , n237084 , n237085 , 
     n237086 , n237087 , n237088 , n237089 , n237090 , n237091 , n237092 , n237093 , n237094 , n237095 , 
     n237096 , n237097 , n237098 , n237099 , n237100 , n237101 , n237102 , n237103 , n237104 , n237105 , 
     n237106 , n237107 , n237108 , n237109 , n237110 , n237111 , n237112 , n237113 , n237114 , n237115 , 
     n237116 , n237117 , n237118 , n237119 , n237120 , n237121 , n237122 , n237123 , n237124 , n237125 , 
     n237126 , n237127 , n237128 , n237129 , n237130 , n237131 , n237132 , n237133 , n237134 , n237135 , 
     n237136 , n237137 , n237138 , n237139 , n237140 , n237141 , n237142 , n237143 , n237144 , n237145 , 
     n237146 , n237147 , n237148 , n237149 , n237150 , n237151 , n237152 , n237153 , n237154 , n237155 , 
     n237156 , n237157 , n237158 , n237159 , n237160 , n237161 , n237162 , n237163 , n237164 , n237165 , 
     n237166 , n237167 , n237168 , n237169 , n237170 , n237171 , n237172 , n237173 , n237174 , n237175 , 
     n237176 , n237177 , n237178 , n237179 , n237180 , n237181 , n237182 , n237183 , n237184 , n237185 , 
     n237186 , n237187 , n237188 , n237189 , n237190 , n237191 , n237192 , n237193 , n237194 , n237195 , 
     n237196 , n237197 , n237198 , n237199 , n237200 , n237201 , n237202 , n237203 , n237204 , n237205 , 
     n237206 , n237207 , n237208 , n237209 , n237210 , n237211 , n237212 , n237213 , n237214 , n237215 , 
     n237216 , n237217 , n237218 , n237219 , n237220 , n237221 , n237222 , n237223 , n237224 , n237225 , 
     n237226 , n237227 , n237228 , n237229 , n237230 , n237231 , n237232 , n237233 , n237234 , n237235 , 
     n237236 , n237237 , n237238 , n237239 , n237240 , n237241 , n237242 , n237243 , n237244 , n237245 , 
     n237246 , n237247 , n237248 , n237249 , n237250 , n237251 , n237252 , n237253 , n237254 , n237255 , 
     n237256 , n237257 , n237258 , n237259 , n237260 , n237261 , n237262 , n237263 , n237264 , n237265 , 
     n237266 , n237267 , n237268 , n237269 , n237270 , n237271 , n237272 , n237273 , n237274 , n237275 , 
     n237276 , n237277 , n237278 , n237279 , n237280 , n237281 , n237282 , n237283 , n237284 , n237285 , 
     n237286 , n237287 , n237288 , n237289 , n237290 , n237291 , n237292 , n237293 , n237294 , n237295 , 
     n237296 , n237297 , n237298 , n237299 , n237300 , n237301 , n237302 , n237303 , n237304 , n237305 , 
     n237306 , n237307 , n237308 , n237309 , n237310 , n237311 , n237312 , n237313 , n237314 , n237315 , 
     n237316 , n237317 , n237318 , n237319 , n237320 , n237321 , n237322 , n237323 , n237324 , n237325 , 
     n237326 , n237327 , n237328 , n237329 , n237330 , n237331 , n237332 , n237333 , n237334 , n237335 , 
     n237336 , n237337 , n237338 , n237339 , n237340 , n237341 , n237342 , n237343 , n237344 , n237345 , 
     n237346 , n237347 , n237348 , n237349 , n237350 , n237351 , n237352 , n237353 , n237354 , n237355 , 
     n237356 , n237357 , n237358 , n237359 , n237360 , n237361 , n237362 , n237363 , n237364 , n237365 , 
     n237366 , n237367 , n237368 , n237369 , n237370 , n237371 , n237372 , n237373 , n237374 , n237375 , 
     n237376 , n237377 , n237378 , n237379 , n237380 , n237381 , n237382 , n237383 , n237384 , n237385 , 
     n237386 , n237387 , n237388 , n237389 , n237390 , n237391 , n237392 , n237393 , n237394 , n237395 , 
     n237396 , n237397 , n237398 , n237399 , n237400 , n237401 , n237402 , n237403 , n237404 , n237405 , 
     n237406 , n237407 , n237408 , n237409 , n237410 , n237411 , n237412 , n237413 , n237414 , n237415 , 
     n237416 , n237417 , n237418 , n237419 , n237420 , n237421 , n237422 , n237423 , n237424 , n237425 , 
     n237426 , n237427 , n237428 , n237429 , n237430 , n237431 , n237432 , n237433 , n237434 , n237435 , 
     n237436 , n237437 , n237438 , n237439 , n237440 , n237441 , n237442 , n237443 , n237444 , n237445 , 
     n237446 , n237447 , n237448 , n237449 , n237450 , n237451 , n237452 , n237453 , n237454 , n237455 , 
     n237456 , n237457 , n237458 , n237459 , n237460 , n237461 , n237462 , n237463 , n237464 , n237465 , 
     n237466 , n237467 , n237468 , n237469 , n237470 , n237471 , n237472 , n237473 , n237474 , n237475 , 
     n237476 , n237477 , n237478 , n237479 , n237480 , n237481 , n237482 , n237483 , n237484 , n237485 , 
     n237486 , n237487 , n237488 , n237489 , n237490 , n237491 , n237492 , n237493 , n237494 , n237495 , 
     n237496 , n237497 , n237498 , n237499 , n237500 , n237501 , n237502 , n237503 , n237504 , n237505 , 
     n237506 , n237507 , n237508 , n237509 , n237510 , n237511 , n237512 , n237513 , n237514 , n237515 , 
     n237516 , n237517 , n237518 , n237519 , n237520 , n237521 , n237522 , n237523 , n237524 , n237525 , 
     n237526 , n237527 , n237528 , n237529 , n237530 , n237531 , n237532 , n237533 , n237534 , n237535 , 
     n237536 , n237537 , n237538 , n237539 , n237540 , n237541 , n237542 , n237543 , n237544 , n237545 , 
     n237546 , n237547 , n237548 , n237549 , n237550 , n237551 , n237552 , n237553 , n237554 , n237555 , 
     n237556 , n237557 , n237558 , n237559 , n237560 , n237561 , n237562 , n237563 , n237564 , n237565 , 
     n237566 , n237567 , n237568 , n237569 , n237570 , n237571 , n237572 , n237573 , n237574 , n237575 , 
     n237576 , n237577 , n237578 , n237579 , n237580 , n237581 , n237582 , n237583 , n237584 , n237585 , 
     n237586 , n237587 , n237588 , n237589 , n237590 , n237591 , n237592 , n237593 , n237594 , n237595 , 
     n237596 , n237597 , n237598 , n237599 , n237600 , n237601 , n237602 , n237603 , n237604 , n237605 , 
     n237606 , n237607 , n237608 , n237609 , n237610 , n237611 , n237612 , n237613 , n237614 , n237615 , 
     n237616 , n237617 , n237618 , n237619 , n237620 , n237621 , n237622 , n237623 , n237624 , n237625 , 
     n237626 , n237627 , n237628 , n237629 , n237630 , n237631 , n237632 , n237633 , n237634 , n237635 , 
     n237636 , n237637 , n237638 , n237639 , n237640 , n237641 , n237642 , n237643 , n237644 , n237645 , 
     n237646 , n237647 , n237648 , n237649 , n237650 , n237651 , n237652 , n237653 , n237654 , n237655 , 
     n237656 , n237657 , n237658 , n237659 , n237660 , n237661 , n237662 , n237663 , n237664 , n237665 , 
     n237666 , n237667 , n237668 , n237669 , n237670 , n237671 , n237672 , n237673 , n237674 , n237675 , 
     n237676 , n237677 , n237678 , n237679 , n237680 , n237681 , n237682 , n237683 , n237684 , n237685 , 
     n237686 , n237687 , n237688 , n237689 , n237690 , n237691 , n237692 , n237693 , n237694 , n237695 , 
     n237696 , n237697 , n237698 , n237699 , n237700 , n237701 , n237702 , n237703 , n237704 , n237705 , 
     n237706 , n237707 , n237708 , n237709 , n237710 , n237711 , n237712 , n237713 , n237714 , n237715 , 
     n237716 , n237717 , n237718 , n237719 , n237720 , n237721 , n237722 , n237723 , n237724 , n237725 , 
     n237726 , n237727 , n237728 , n237729 , n237730 , n237731 , n237732 , n237733 , n237734 , n237735 , 
     n237736 , n237737 , n237738 , n237739 , n237740 , n237741 , n237742 , n237743 , n237744 , n237745 , 
     n237746 , n237747 , n237748 , n237749 , n237750 , n237751 , n237752 , n237753 , n237754 , n237755 , 
     n237756 , n237757 , n237758 , n237759 , n237760 , n237761 , n237762 , n237763 , n237764 , n237765 , 
     n237766 , n237767 , n237768 , n237769 , n237770 , n237771 , n237772 , n237773 , n237774 , n237775 , 
     n237776 , n237777 , n237778 , n237779 , n237780 , n237781 , n237782 , n237783 , n237784 , n237785 , 
     n237786 , n237787 , n237788 , n237789 , n237790 , n237791 , n237792 , n237793 , n237794 , n237795 , 
     n237796 , n237797 , n237798 , n237799 , n237800 , n237801 , n237802 , n237803 , n237804 , n237805 , 
     n237806 , n237807 , n237808 , n237809 , n237810 , n237811 , n237812 , n237813 , n237814 , n237815 , 
     n237816 , n237817 , n237818 , n237819 , n237820 , n237821 , n237822 , n237823 , n237824 , n237825 , 
     n237826 , n237827 , n237828 , n237829 , n237830 , n237831 , n237832 , n237833 , n237834 , n237835 , 
     n237836 , n237837 , n237838 , n237839 , n237840 , n237841 , n237842 , n237843 , n237844 , n237845 , 
     n237846 , n237847 , n237848 , n237849 , n237850 , n237851 , n237852 , n237853 , n237854 , n237855 , 
     n237856 , n237857 , n237858 , n237859 , n237860 , n237861 , n237862 , n237863 , n237864 , n237865 , 
     n237866 , n237867 , n237868 , n237869 , n237870 , n237871 , n237872 , n237873 , n237874 , n237875 , 
     n237876 , n237877 , n237878 , n237879 , n237880 , n237881 , n237882 , n237883 , n237884 , n237885 , 
     n237886 , n237887 , n237888 , n237889 , n237890 , n237891 , n237892 , n237893 , n237894 , n237895 , 
     n237896 , n237897 , n237898 , n237899 , n237900 , n237901 , n237902 , n237903 , n237904 , n237905 , 
     n237906 , n237907 , n237908 , n237909 , n237910 , n237911 , n237912 , n237913 , n237914 , n237915 , 
     n237916 , n237917 , n237918 , n237919 , n237920 , n237921 , n237922 , n237923 , n237924 , n237925 , 
     n237926 , n237927 , n237928 , n237929 , n237930 , n237931 , n237932 , n237933 , n237934 , n237935 , 
     n237936 , n237937 , n237938 , n237939 , n237940 , n237941 , n237942 , n237943 , n237944 , n237945 , 
     n237946 , n237947 , n237948 , n237949 , n237950 , n237951 , n237952 , n237953 , n237954 , n237955 , 
     n237956 , n237957 , n237958 , n237959 , n237960 , n237961 , n237962 , n237963 , n237964 , n237965 , 
     n237966 , n237967 , n237968 , n237969 , n237970 , n237971 , n237972 , n237973 , n237974 , n237975 , 
     n237976 , n237977 , n237978 , n237979 , n237980 , n237981 , n237982 , n237983 , n237984 , n237985 , 
     n237986 , n237987 , n237988 , n237989 , n237990 , n237991 , n237992 , n237993 , n237994 , n237995 , 
     n237996 , n237997 , n237998 , n237999 , n238000 , n238001 , n238002 , n238003 , n238004 , n238005 , 
     n238006 , n238007 , n238008 , n238009 , n238010 , n238011 , n238012 , n238013 , n238014 , n238015 , 
     n238016 , n238017 , n238018 , n238019 , n238020 , n238021 , n238022 , n238023 , n238024 , n238025 , 
     n238026 , n238027 , n238028 , n238029 , n238030 , n238031 , n238032 , n238033 , n238034 , n238035 , 
     n238036 , n238037 , n238038 , n238039 , n238040 , n238041 , n238042 , n238043 , n238044 , n238045 , 
     n238046 , n238047 , n238048 , n238049 , n238050 , n238051 , n238052 , n238053 , n238054 , n238055 , 
     n238056 , n238057 , n238058 , n238059 , n238060 , n238061 , n238062 , n238063 , n238064 , n238065 , 
     n238066 , n238067 , n238068 , n238069 , n238070 , n238071 , n238072 , n238073 , n238074 , n238075 , 
     n238076 , n238077 , n238078 , n238079 , n238080 , n238081 , n238082 , n238083 , n238084 , n238085 , 
     n238086 , n238087 , n238088 , n238089 , n238090 , n238091 , n238092 , n238093 , n238094 , n238095 , 
     n238096 , n238097 , n238098 , n238099 , n238100 , n238101 , n238102 , n238103 , n238104 , n238105 , 
     n238106 , n238107 , n238108 , n238109 , n238110 , n238111 , n238112 , n238113 , n238114 , n238115 , 
     n238116 , n238117 , n238118 , n238119 , n238120 , n238121 , n238122 , n238123 , n238124 , n238125 , 
     n238126 , n238127 , n238128 , n238129 , n238130 , n238131 , n238132 , n238133 , n238134 , n238135 , 
     n238136 , n238137 , n238138 , n238139 , n238140 , n238141 , n238142 , n238143 , n238144 , n238145 , 
     n238146 , n238147 , n238148 , n238149 , n238150 , n238151 , n238152 , n238153 , n238154 , n238155 , 
     n238156 , n238157 , n238158 , n238159 , n238160 , n238161 , n238162 , n238163 , n238164 , n238165 , 
     n238166 , n238167 , n238168 , n238169 , n238170 , n238171 , n238172 , n238173 , n238174 , n238175 , 
     n238176 , n238177 , n238178 , n238179 , n238180 , n238181 , n238182 , n238183 , n238184 , n238185 , 
     n238186 , n238187 , n238188 , n238189 , n238190 , n238191 , n238192 , n238193 , n238194 , n238195 , 
     n238196 , n238197 , n238198 , n238199 , n238200 , n238201 , n238202 , n238203 , n238204 , n238205 , 
     n238206 , n238207 , n238208 , n238209 , n238210 , n238211 , n238212 , n238213 , n238214 , n238215 , 
     n238216 , n238217 , n238218 , n238219 , n238220 , n238221 , n238222 , n238223 , n238224 , n238225 , 
     n238226 , n238227 , n238228 , n238229 , n238230 , n238231 , n238232 , n238233 , n238234 , n238235 , 
     n238236 , n238237 , n238238 , n238239 , n238240 , n238241 , n238242 , n238243 , n238244 , n238245 , 
     n238246 , n238247 , n238248 , n238249 , n238250 , n238251 , n238252 , n238253 , n238254 , n238255 , 
     n238256 , n238257 , n238258 , n238259 , n238260 , n238261 , n238262 , n238263 , n238264 , n238265 , 
     n238266 , n238267 , n238268 , n238269 , n238270 , n238271 , n238272 , n238273 , n238274 , n238275 , 
     n238276 , n238277 , n238278 , n238279 , n238280 , n238281 , n238282 , n238283 , n238284 , n238285 , 
     n238286 , n238287 , n238288 , n238289 , n238290 , n238291 , n238292 , n238293 , n238294 , n238295 , 
     n238296 , n238297 , n238298 , n238299 , n238300 , n238301 , n238302 , n238303 , n238304 , n238305 , 
     n238306 , n238307 , n238308 , n238309 , n238310 , n238311 , n238312 , n238313 , n238314 , n238315 , 
     n238316 , n238317 , n238318 , n238319 , n238320 , n238321 , n238322 , n238323 , n238324 , n238325 , 
     n238326 , n238327 , n238328 , n238329 , n238330 , n238331 , n238332 , n238333 , n238334 , n238335 , 
     n238336 , n238337 , n238338 , n238339 , n238340 , n238341 , n238342 , n238343 , n238344 , n238345 , 
     n238346 , n238347 , n238348 , n238349 , n238350 , n238351 , n238352 , n238353 , n238354 , n238355 , 
     n238356 , n238357 , n238358 , n238359 , n238360 , n238361 , n238362 , n238363 , n238364 , n238365 , 
     n238366 , n238367 , n238368 , n238369 , n238370 , n238371 , n238372 , n238373 , n238374 , n238375 , 
     n238376 , n238377 , n238378 , n238379 , n238380 , n238381 , n238382 , n238383 , n238384 , n238385 , 
     n238386 , n238387 , n238388 , n238389 , n238390 , n238391 , n238392 , n238393 , n238394 , n238395 , 
     n238396 , n238397 , n238398 , n238399 , n238400 , n238401 , n238402 , n238403 , n238404 , n238405 , 
     n238406 , n238407 , n238408 , n238409 , n238410 , n238411 , n238412 , n238413 , n238414 , n238415 , 
     n238416 , n238417 , n238418 , n238419 , n238420 , n238421 , n238422 , n238423 , n238424 , n238425 , 
     n238426 , n238427 , n238428 , n238429 , n238430 , n238431 , n238432 , n238433 , n238434 , n238435 , 
     n238436 , n238437 , n238438 , n238439 , n238440 , n238441 , n238442 , n238443 , n238444 , n238445 , 
     n238446 , n238447 , n238448 , n238449 , n238450 , n238451 , n238452 , n238453 , n238454 , n238455 , 
     n238456 , n238457 , n238458 , n238459 , n238460 , n238461 , n238462 , n238463 , n238464 , n238465 , 
     n238466 , n238467 , n238468 , n238469 , n238470 , n238471 , n238472 , n238473 , n238474 , n238475 , 
     n238476 , n238477 , n238478 , n238479 , n238480 , n238481 , n238482 , n238483 , n238484 , n238485 , 
     n238486 , n238487 , n238488 , n238489 , n238490 , n238491 , n238492 , n238493 , n238494 , n238495 , 
     n238496 , n238497 , n238498 , n238499 , n238500 , n238501 , n238502 , n238503 , n238504 , n238505 , 
     n238506 , n238507 , n238508 , n238509 , n238510 , n238511 , n238512 , n238513 , n238514 , n238515 , 
     n238516 , n238517 , n238518 , n238519 , n238520 , n238521 , n238522 , n238523 , n238524 , n238525 , 
     n238526 , n238527 , n238528 , n238529 , n238530 , n238531 , n238532 , n238533 , n238534 , n238535 , 
     n238536 , n238537 , n238538 , n238539 , n238540 , n238541 , n238542 , n238543 , n238544 , n238545 , 
     n238546 , n238547 , n238548 , n238549 , n238550 , n238551 , n238552 , n238553 , n238554 , n238555 , 
     n238556 , n238557 , n238558 , n238559 , n238560 , n238561 , n238562 , n238563 , n238564 , n238565 , 
     n238566 , n238567 , n238568 , n238569 , n238570 , n238571 , n238572 , n238573 , n238574 , n238575 , 
     n238576 , n238577 , n238578 , n238579 , n238580 , n238581 , n238582 , n238583 , n238584 , n238585 , 
     n238586 , n238587 , n238588 , n238589 , n238590 , n238591 , n238592 , n238593 , n238594 , n238595 , 
     n238596 , n238597 , n238598 , n238599 , n238600 , n238601 , n238602 , n238603 , n238604 , n238605 , 
     n238606 , n238607 , n238608 , n238609 , n238610 , n238611 , n238612 , n238613 , n238614 , n238615 , 
     n238616 , n238617 , n238618 , n238619 , n238620 , n238621 , n238622 , n238623 , n238624 , n238625 , 
     n238626 , n238627 , n238628 , n238629 , n238630 , n238631 , n238632 , n238633 , n238634 , n238635 , 
     n238636 , n238637 , n238638 , n238639 , n238640 , n238641 , n238642 , n238643 , n238644 , n238645 , 
     n238646 , n238647 , n238648 , n238649 , n238650 , n238651 , n238652 , n238653 , n238654 , n238655 , 
     n238656 , n238657 , n238658 , n238659 , n238660 , n238661 , n238662 , n238663 , n238664 , n238665 , 
     n238666 , n238667 , n238668 , n238669 , n238670 , n238671 , n238672 , n238673 , n238674 , n238675 , 
     n238676 , n238677 , n238678 , n238679 , n238680 , n238681 , n238682 , n238683 , n238684 , n238685 , 
     n238686 , n238687 , n238688 , n238689 , n238690 , n238691 , n238692 , n238693 , n238694 , n238695 , 
     n238696 , n238697 , n238698 , n238699 , n238700 , n238701 , n238702 , n238703 , n238704 , n238705 , 
     n238706 , n238707 , n238708 , n238709 , n238710 , n238711 , n238712 , n238713 , n238714 , n238715 , 
     n238716 , n238717 , n238718 , n238719 , n238720 , n238721 , n238722 , n238723 , n238724 , n238725 , 
     n238726 , n238727 , n238728 , n238729 , n238730 , n238731 , n238732 , n238733 , n238734 , n238735 , 
     n238736 , n238737 , n238738 , n238739 , n238740 , n238741 , n238742 , n238743 , n238744 , n238745 , 
     n238746 , n238747 , n238748 , n238749 , n238750 , n238751 , n238752 , n238753 , n238754 , n238755 , 
     n238756 , n238757 , n238758 , n238759 , n238760 , n238761 , n238762 , n238763 , n238764 , n238765 , 
     n238766 , n238767 , n238768 , n238769 , n238770 , n238771 , n238772 , n238773 , n238774 , n238775 , 
     n238776 , n238777 , n238778 , n238779 , n238780 , n238781 , n238782 , n238783 , n238784 , n238785 , 
     n238786 , n238787 , n238788 , n238789 , n238790 , n238791 , n238792 , n238793 , n238794 , n238795 , 
     n238796 , n238797 , n238798 , n238799 , n238800 , n238801 , n238802 , n238803 , n238804 , n238805 , 
     n238806 , n238807 , n238808 , n238809 , n238810 , n238811 , n238812 , n238813 , n238814 , n238815 , 
     n238816 , n238817 , n238818 , n238819 , n238820 , n238821 , n238822 , n238823 , n238824 , n238825 , 
     n238826 , n238827 , n238828 , n238829 , n238830 , n238831 , n238832 , n238833 , n238834 , n238835 , 
     n238836 , n238837 , n238838 , n238839 , n238840 , n238841 , n238842 , n238843 , n238844 , n238845 , 
     n238846 , n238847 , n238848 , n238849 , n238850 , n238851 , n238852 , n238853 , n238854 , n238855 , 
     n238856 , n238857 , n238858 , n238859 , n238860 , n238861 , n238862 , n238863 , n238864 , n238865 , 
     n238866 , n238867 , n238868 , n238869 , n238870 , n238871 , n238872 , n238873 , n238874 , n238875 , 
     n238876 , n238877 , n238878 , n238879 , n238880 , n238881 , n238882 , n238883 , n238884 , n238885 , 
     n238886 , n238887 , n238888 , n238889 , n238890 , n238891 , n238892 , n238893 , n238894 , n238895 , 
     n238896 , n238897 , n238898 , n238899 , n238900 , n238901 , n238902 , n238903 , n238904 , n238905 , 
     n238906 , n238907 , n238908 , n238909 , n238910 , n238911 , n238912 , n238913 , n238914 , n238915 , 
     n238916 , n238917 , n238918 , n238919 , n238920 , n238921 , n238922 , n238923 , n238924 , n238925 , 
     n238926 , n238927 , n238928 , n238929 , n238930 , n238931 , n238932 , n238933 , n238934 , n238935 , 
     n238936 , n238937 , n238938 , n238939 , n238940 , n238941 , n238942 , n238943 , n238944 , n238945 , 
     n238946 , n238947 , n238948 , n238949 , n238950 , n238951 , n238952 , n238953 , n238954 , n238955 , 
     n238956 , n238957 , n238958 , n238959 , n238960 , n238961 , n238962 , n238963 , n238964 , n238965 , 
     n238966 , n238967 , n238968 , n238969 , n238970 , n238971 , n238972 , n238973 , n238974 , n238975 , 
     n238976 , n238977 , n238978 , n238979 , n238980 , n238981 , n238982 , n238983 , n238984 , n238985 , 
     n238986 , n238987 , n238988 , n238989 , n238990 , n238991 , n238992 , n238993 , n238994 , n238995 , 
     n238996 , n238997 , n238998 , n238999 , n239000 , n239001 , n239002 , n239003 , n239004 , n239005 , 
     n239006 , n239007 , n239008 , n239009 , n239010 , n239011 , n239012 , n239013 , n239014 , n239015 , 
     n239016 , n239017 , n239018 , n239019 , n239020 , n239021 , n239022 , n239023 , n239024 , n239025 , 
     n239026 , n239027 , n239028 , n239029 , n239030 , n239031 , n239032 , n239033 , n239034 , n239035 , 
     n239036 , n239037 , n239038 , n239039 , n239040 , n239041 , n239042 , n239043 , n239044 , n239045 , 
     n239046 , n239047 , n239048 , n239049 , n239050 , n239051 , n239052 , n239053 , n239054 , n239055 , 
     n239056 , n239057 , n239058 , n239059 , n239060 , n239061 , n239062 , n239063 , n239064 , n239065 , 
     n239066 , n239067 , n239068 , n239069 , n239070 , n239071 , n239072 , n239073 , n239074 , n239075 , 
     n239076 , n239077 , n239078 , n239079 , n239080 , n239081 , n239082 , n239083 , n239084 , n239085 , 
     n239086 , n239087 , n239088 , n239089 , n239090 , n239091 , n239092 , n239093 , n239094 , n239095 , 
     n239096 , n239097 , n239098 , n239099 , n239100 , n239101 , n239102 , n239103 , n239104 , n239105 , 
     n239106 , n239107 , n239108 , n239109 , n239110 , n239111 , n239112 , n239113 , n239114 , n239115 , 
     n239116 , n239117 , n239118 , n239119 , n239120 , n239121 , n239122 , n239123 , n239124 , n239125 , 
     n239126 , n239127 , n239128 , n239129 , n239130 , n239131 , n239132 , n239133 , n239134 , n239135 , 
     n239136 , n239137 , n239138 , n239139 , n239140 , n239141 , n239142 , n239143 , n239144 , n239145 , 
     n239146 , n239147 , n239148 , n239149 , n239150 , n239151 , n239152 , n239153 , n239154 , n239155 , 
     n239156 , n239157 , n239158 , n239159 , n239160 , n239161 , n239162 , n239163 , n239164 , n239165 , 
     n239166 , n239167 , n239168 , n239169 , n239170 , n239171 , n239172 , n239173 , n239174 , n239175 , 
     n239176 , n239177 , n239178 , n239179 , n239180 , n239181 , n239182 , n239183 , n239184 , n239185 , 
     n239186 , n239187 , n239188 , n239189 , n239190 , n239191 , n239192 , n239193 , n239194 , n239195 , 
     n239196 , n239197 , n239198 , n239199 , n239200 , n239201 , n239202 , n239203 , n239204 , n239205 , 
     n239206 , n239207 , n239208 , n239209 , n239210 , n239211 , n239212 , n239213 , n239214 , n239215 , 
     n239216 , n239217 , n239218 , n239219 , n239220 , n239221 , n239222 , n239223 , n239224 , n239225 , 
     n239226 , n239227 , n239228 , n239229 , n239230 , n239231 , n239232 , n239233 , n239234 , n239235 , 
     n239236 , n239237 , n239238 , n239239 , n239240 , n239241 , n239242 , n239243 , n239244 , n239245 , 
     n239246 , n239247 , n239248 , n239249 , n239250 , n239251 , n239252 , n239253 , n239254 , n239255 , 
     n239256 , n239257 , n239258 , n239259 , n239260 , n239261 , n239262 , n239263 , n239264 , n239265 , 
     n239266 , n239267 , n239268 , n239269 , n239270 , n239271 , n239272 , n239273 , n239274 , n239275 , 
     n239276 , n239277 , n239278 , n239279 , n239280 , n239281 , n239282 , n239283 , n239284 , n239285 , 
     n239286 , n239287 , n239288 , n239289 , n239290 , n239291 , n239292 , n239293 , n239294 , n239295 , 
     n239296 , n239297 , n239298 , n239299 , n239300 , n239301 , n239302 , n239303 , n239304 , n239305 , 
     n239306 , n239307 , n239308 , n239309 , n239310 , n239311 , n239312 , n239313 , n239314 , n239315 , 
     n239316 , n239317 , n239318 , n239319 , n239320 , n239321 , n239322 , n239323 , n239324 , n239325 , 
     n239326 , n239327 , n239328 , n239329 , n239330 , n239331 , n239332 , n239333 , n239334 , n239335 , 
     n239336 , n239337 , n239338 , n239339 , n239340 , n239341 , n239342 , n239343 , n239344 , n239345 , 
     n239346 , n239347 , n239348 , n239349 , n239350 , n239351 , n239352 , n239353 , n239354 , n239355 , 
     n239356 , n239357 , n239358 , n239359 , n239360 , n239361 , n239362 , n239363 , n239364 , n239365 , 
     n239366 , n239367 , n239368 , n239369 , n239370 , n239371 , n239372 , n239373 , n239374 , n239375 , 
     n239376 , n239377 , n239378 , n239379 , n239380 , n239381 , n239382 , n239383 , n239384 , n239385 , 
     n239386 , n239387 , n239388 , n239389 , n239390 , n239391 , n239392 , n239393 , n239394 , n239395 , 
     n239396 , n239397 , n239398 , n239399 , n239400 , n239401 , n239402 , n239403 , n239404 , n239405 , 
     n239406 , n239407 , n239408 , n239409 , n239410 , n239411 , n239412 , n239413 , n239414 , n239415 , 
     n239416 , n239417 , n239418 , n239419 , n239420 , n239421 , n239422 , n239423 , n239424 , n239425 , 
     n239426 , n239427 , n239428 , n239429 , n239430 , n239431 , n239432 , n239433 , n239434 , n239435 , 
     n239436 , n239437 , n239438 , n239439 , n239440 , n239441 , n239442 , n239443 , n239444 , n239445 , 
     n239446 , n239447 , n239448 , n239449 , n239450 , n239451 , n239452 , n239453 , n239454 , n239455 , 
     n239456 , n239457 , n239458 , n239459 , n239460 , n239461 , n239462 , n239463 , n239464 , n239465 , 
     n239466 , n239467 , n239468 , n239469 , n239470 , n239471 , n239472 , n239473 , n239474 , n239475 , 
     n239476 , n239477 , n239478 , n239479 , n239480 , n239481 , n239482 , n239483 , n239484 , n239485 , 
     n239486 , n239487 , n239488 , n239489 , n239490 , n239491 , n239492 , n239493 , n239494 , n239495 , 
     n239496 , n239497 , n239498 , n239499 , n239500 , n239501 , n239502 , n239503 , n239504 , n239505 , 
     n239506 , n239507 , n239508 , n239509 , n239510 , n239511 , n239512 , n239513 , n239514 , n239515 , 
     n239516 , n239517 , n239518 , n239519 , n239520 , n239521 , n239522 , n239523 , n239524 , n239525 , 
     n239526 , n239527 , n239528 , n239529 , n239530 , n239531 , n239532 , n239533 , n239534 , n239535 , 
     n239536 , n239537 , n239538 , n239539 , n239540 , n239541 , n239542 , n239543 , n239544 , n239545 , 
     n239546 , n239547 , n239548 , n239549 , n239550 , n239551 , n239552 , n239553 , n239554 , n239555 , 
     n239556 , n239557 , n239558 , n239559 , n239560 , n239561 , n239562 , n239563 , n239564 , n239565 , 
     n239566 , n239567 , n239568 , n239569 , n239570 , n239571 , n239572 , n239573 , n239574 , n239575 , 
     n239576 , n239577 , n239578 , n239579 , n239580 , n239581 , n239582 , n239583 , n239584 , n239585 , 
     n239586 , n239587 , n239588 , n239589 , n239590 , n239591 , n239592 , n239593 , n239594 , n239595 , 
     n239596 , n239597 , n239598 , n239599 , n239600 , n239601 , n239602 , n239603 , n239604 , n239605 , 
     n239606 , n239607 , n239608 , n239609 , n239610 , n239611 , n239612 , n239613 , n239614 , n239615 , 
     n239616 , n239617 , n239618 , n239619 , n239620 , n239621 , n239622 , n239623 , n239624 , n239625 , 
     n239626 , n239627 , n239628 , n239629 , n239630 , n239631 , n239632 , n239633 , n239634 , n239635 , 
     n239636 , n239637 , n239638 , n239639 , n239640 , n239641 , n239642 , n239643 , n239644 , n239645 , 
     n239646 , n239647 , n239648 , n239649 , n239650 , n239651 , n239652 , n239653 , n239654 , n239655 , 
     n239656 , n239657 , n239658 , n239659 , n239660 , n239661 , n239662 , n239663 , n239664 , n239665 , 
     n239666 , n239667 , n239668 , n239669 , n239670 , n239671 , n239672 , n239673 , n239674 , n239675 , 
     n239676 , n239677 , n239678 , n239679 , n239680 , n239681 , n239682 , n239683 , n239684 , n239685 , 
     n239686 , n239687 , n239688 , n239689 , n239690 , n239691 , n239692 , n239693 , n239694 , n239695 , 
     n239696 , n239697 , n239698 , n239699 , n239700 , n239701 , n239702 , n239703 , n239704 , n239705 , 
     n239706 , n239707 , n239708 , n239709 , n239710 , n239711 , n239712 , n239713 , n239714 , n239715 , 
     n239716 , n239717 , n239718 , n239719 , n239720 , n239721 , n239722 , n239723 , n239724 , n239725 , 
     n239726 , n239727 , n239728 , n239729 , n239730 , n239731 , n239732 , n239733 , n239734 , n239735 , 
     n239736 , n239737 , n239738 , n239739 , n239740 , n239741 , n239742 , n239743 , n239744 , n239745 , 
     n239746 , n239747 , n239748 , n239749 , n239750 , n239751 , n239752 , n239753 , n239754 , n239755 , 
     n239756 , n239757 , n239758 , n239759 , n239760 , n239761 , n239762 , n239763 , n239764 , n239765 , 
     n239766 , n239767 , n239768 , n239769 , n239770 , n239771 , n239772 , n239773 , n239774 , n239775 , 
     n239776 , n239777 , n239778 , n239779 , n239780 , n239781 , n239782 , n239783 , n239784 , n239785 , 
     n239786 , n239787 , n239788 , n239789 , n239790 , n239791 , n239792 , n239793 , n239794 , n239795 , 
     n239796 , n239797 , n239798 , n239799 , n239800 , n239801 , n239802 , n239803 , n239804 , n239805 , 
     n239806 , n239807 , n239808 , n239809 , n239810 , n239811 , n239812 , n239813 , n239814 , n239815 , 
     n239816 , n239817 , n239818 , n239819 , n239820 , n239821 , n239822 , n239823 , n239824 , n239825 , 
     n239826 , n239827 , n239828 , n239829 , n239830 , n239831 , n239832 , n239833 , n239834 , n239835 , 
     n239836 , n239837 , n239838 , n239839 , n239840 , n239841 , n239842 , n239843 , n239844 , n239845 , 
     n239846 , n239847 , n239848 , n239849 , n239850 , n239851 , n239852 , n239853 , n239854 , n239855 , 
     n239856 , n239857 , n239858 , n239859 , n239860 , n239861 , n239862 , n239863 , n239864 , n239865 , 
     n239866 , n239867 , n239868 , n239869 , n239870 , n239871 , n239872 , n239873 , n239874 , n239875 , 
     n239876 , n239877 , n239878 , n239879 , n239880 , n239881 , n239882 , n239883 , n239884 , n239885 , 
     n239886 , n239887 , n239888 , n239889 , n239890 , n239891 , n239892 , n239893 , n239894 , n239895 , 
     n239896 , n239897 , n239898 , n239899 , n239900 , n239901 , n239902 , n239903 , n239904 , n239905 , 
     n239906 , n239907 , n239908 , n239909 , n239910 , n239911 , n239912 , n239913 , n239914 , n239915 , 
     n239916 , n239917 , n239918 , n239919 , n239920 , n239921 , n239922 , n239923 , n239924 , n239925 , 
     n239926 , n239927 , n239928 , n239929 , n239930 , n239931 , n239932 , n239933 , n239934 , n239935 , 
     n239936 , n239937 , n239938 , n239939 , n239940 , n239941 , n239942 , n239943 , n239944 , n239945 , 
     n239946 , n239947 , n239948 , n239949 , n239950 , n239951 , n239952 , n239953 , n239954 , n239955 , 
     n239956 , n239957 , n239958 , n239959 , n239960 , n239961 , n239962 , n239963 , n239964 , n239965 , 
     n239966 , n239967 , n239968 , n239969 , n239970 , n239971 , n239972 , n239973 , n239974 , n239975 , 
     n239976 , n239977 , n239978 , n239979 , n239980 , n239981 , n239982 , n239983 , n239984 , n239985 , 
     n239986 , n239987 , n239988 , n239989 , n239990 , n239991 , n239992 , n239993 , n239994 , n239995 , 
     n239996 , n239997 , n239998 , n239999 , n240000 , n240001 , n240002 , n240003 , n240004 , n240005 , 
     n240006 , n240007 , n240008 , n240009 , n240010 , n240011 , n240012 , n240013 , n240014 , n240015 , 
     n240016 , n240017 , n240018 , n240019 , n240020 , n240021 , n240022 , n240023 , n240024 , n240025 , 
     n240026 , n240027 , n240028 , n240029 , n240030 , n240031 , n240032 , n240033 , n240034 , n240035 , 
     n240036 , n240037 , n240038 , n240039 , n240040 , n240041 , n240042 , n240043 , n240044 , n240045 , 
     n240046 , n240047 , n240048 , n240049 , n240050 , n240051 , n240052 , n240053 , n240054 , n240055 , 
     n240056 , n240057 , n240058 , n240059 , n240060 , n240061 , n240062 , n240063 , n240064 , n240065 , 
     n240066 , n240067 , n240068 , n240069 , n240070 , n240071 , n240072 , n240073 , n240074 , n240075 , 
     n240076 , n240077 , n240078 , n240079 , n240080 , n240081 , n240082 , n240083 , n240084 , n240085 , 
     n240086 , n240087 , n240088 , n240089 , n240090 , n240091 , n240092 , n240093 , n240094 , n240095 , 
     n240096 , n240097 , n240098 , n240099 , n240100 , n240101 , n240102 , n240103 , n240104 , n240105 , 
     n240106 , n240107 , n240108 , n240109 , n240110 , n240111 , n240112 , n240113 , n240114 , n240115 , 
     n240116 , n240117 , n240118 , n240119 , n240120 , n240121 , n240122 , n240123 , n240124 , n240125 , 
     n240126 , n240127 , n240128 , n240129 , n240130 , n240131 , n240132 , n240133 , n240134 , n240135 , 
     n240136 , n240137 , n240138 , n240139 , n240140 , n240141 , n240142 , n240143 , n240144 , n240145 , 
     n240146 , n240147 , n240148 , n240149 , n240150 , n240151 , n240152 , n240153 , n240154 , n240155 , 
     n240156 , n240157 , n240158 , n240159 , n240160 , n240161 , n240162 , n240163 , n240164 , n240165 , 
     n240166 , n240167 , n240168 , n240169 , n240170 , n240171 , n240172 , n240173 , n240174 , n240175 , 
     n240176 , n240177 , n240178 , n240179 , n240180 , n240181 , n240182 , n240183 , n240184 , n240185 , 
     n240186 , n240187 , n240188 , n240189 , n240190 , n240191 , n240192 , n240193 , n240194 , n240195 , 
     n240196 , n240197 , n240198 , n240199 , n240200 , n240201 , n240202 , n240203 , n240204 , n240205 , 
     n240206 , n240207 , n240208 , n240209 , n240210 , n240211 , n240212 , n240213 , n240214 , n240215 , 
     n240216 , n240217 , n240218 , n240219 , n240220 , n240221 , n240222 , n240223 , n240224 , n240225 , 
     n240226 , n240227 , n240228 , n240229 , n240230 , n240231 , n240232 , n240233 , n240234 , n240235 , 
     n240236 , n240237 , n240238 , n240239 , n240240 , n240241 , n240242 , n240243 , n240244 , n240245 , 
     n240246 , n240247 , n240248 , n240249 , n240250 , n240251 , n240252 , n240253 , n240254 , n240255 , 
     n240256 , n240257 , n240258 , n240259 , n240260 , n240261 , n240262 , n240263 , n240264 , n240265 , 
     n240266 , n240267 , n240268 , n240269 , n240270 , n240271 , n240272 , n240273 , n240274 , n240275 , 
     n240276 , n240277 , n240278 , n240279 , n240280 , n240281 , n240282 , n240283 , n240284 , n240285 , 
     n240286 , n240287 , n240288 , n240289 , n240290 , n240291 , n240292 , n240293 , n240294 , n240295 , 
     n240296 , n240297 , n240298 , n240299 , n240300 , n240301 , n240302 , n240303 , n240304 , n240305 , 
     n240306 , n240307 , n240308 , n240309 , n240310 , n240311 , n240312 , n240313 , n240314 , n240315 , 
     n240316 , n240317 , n240318 , n240319 , n240320 , n240321 , n240322 , n240323 , n240324 , n240325 , 
     n240326 , n240327 , n240328 , n240329 , n240330 , n240331 , n240332 , n240333 , n240334 , n240335 , 
     n240336 , n240337 , n240338 , n240339 , n240340 , n240341 , n240342 , n240343 , n240344 , n240345 , 
     n240346 , n240347 , n240348 , n240349 , n240350 , n240351 , n240352 , n240353 , n240354 , n240355 , 
     n240356 , n240357 , n240358 , n240359 , n240360 , n240361 , n240362 , n240363 , n240364 , n240365 , 
     n240366 , n240367 , n240368 , n240369 , n240370 , n240371 , n240372 , n240373 , n240374 , n240375 , 
     n240376 , n240377 , n240378 , n240379 , n240380 , n240381 , n240382 , n240383 , n240384 , n240385 , 
     n240386 , n240387 , n240388 , n240389 , n240390 , n240391 , n240392 , n240393 , n240394 , n240395 , 
     n240396 , n240397 , n240398 , n240399 , n240400 , n240401 , n240402 , n240403 , n240404 , n240405 , 
     n240406 , n240407 , n240408 , n240409 , n240410 , n240411 , n240412 , n240413 , n240414 , n240415 , 
     n240416 , n240417 , n240418 , n240419 , n240420 , n240421 , n240422 , n240423 , n240424 , n240425 , 
     n240426 , n240427 , n240428 , n240429 , n240430 , n240431 , n240432 , n240433 , n240434 , n240435 , 
     n240436 , n240437 , n240438 , n240439 , n240440 , n240441 , n240442 , n240443 , n240444 , n240445 , 
     n240446 , n240447 , n240448 , n240449 , n240450 , n240451 , n240452 , n240453 , n240454 , n240455 , 
     n240456 , n240457 , n240458 , n240459 , n240460 , n240461 , n240462 , n240463 , n240464 , n240465 , 
     n240466 , n240467 , n240468 , n240469 , n240470 , n240471 , n240472 , n240473 , n240474 , n240475 , 
     n240476 , n240477 , n240478 , n240479 , n240480 , n240481 , n240482 , n240483 , n240484 , n240485 , 
     n240486 , n240487 , n240488 , n240489 , n240490 , n240491 , n240492 , n240493 , n240494 , n240495 , 
     n240496 , n240497 , n240498 , n240499 , n240500 , n240501 , n240502 , n240503 , n240504 , n240505 , 
     n240506 , n240507 , n240508 , n240509 , n240510 , n240511 , n240512 , n240513 , n240514 , n240515 , 
     n240516 , n240517 , n240518 , n240519 , n240520 , n240521 , n240522 , n240523 , n240524 , n240525 , 
     n240526 , n240527 , n240528 , n240529 , n240530 , n240531 , n240532 , n240533 , n240534 , n240535 , 
     n240536 , n240537 , n240538 , n240539 , n240540 , n240541 , n240542 , n240543 , n240544 , n240545 , 
     n240546 , n240547 , n240548 , n240549 , n240550 , n240551 , n240552 , n240553 , n240554 , n240555 , 
     n240556 , n240557 , n240558 , n240559 , n240560 , n240561 , n240562 , n240563 , n240564 , n240565 , 
     n240566 , n240567 , n240568 , n240569 , n240570 , n240571 , n240572 , n240573 , n240574 , n240575 , 
     n240576 , n240577 , n240578 , n240579 , n240580 , n240581 , n240582 , n240583 , n240584 , n240585 , 
     n240586 , n240587 , n240588 , n240589 , n240590 , n240591 , n240592 , n240593 , n240594 , n240595 , 
     n240596 , n240597 , n240598 , n240599 , n240600 , n240601 , n240602 , n240603 , n240604 , n240605 , 
     n240606 , n240607 , n240608 , n240609 , n240610 , n240611 , n240612 , n240613 , n240614 , n240615 , 
     n240616 , n240617 , n240618 , n240619 , n240620 , n240621 , n240622 , n240623 , n240624 , n240625 , 
     n240626 , n240627 , n240628 , n240629 , n240630 , n240631 , n240632 , n240633 , n240634 , n240635 , 
     n240636 , n240637 , n240638 , n240639 , n240640 , n240641 , n240642 , n240643 , n240644 , n240645 , 
     n240646 , n240647 , n240648 , n240649 , n240650 , n240651 , n240652 , n240653 , n240654 , n240655 , 
     n240656 , n240657 , n240658 , n240659 , n240660 , n240661 , n240662 , n240663 , n240664 , n240665 , 
     n240666 , n240667 , n240668 , n240669 , n240670 , n240671 , n240672 , n240673 , n240674 , n240675 , 
     n240676 , n240677 , n240678 , n240679 , n240680 , n240681 , n240682 , n240683 , n240684 , n240685 , 
     n240686 , n240687 , n240688 , n240689 , n240690 , n240691 , n240692 , n240693 , n240694 , n240695 , 
     n240696 , n240697 , n240698 , n240699 , n240700 , n240701 , n240702 , n240703 , n240704 , n240705 , 
     n240706 , n240707 , n240708 , n240709 , n240710 , n240711 , n240712 , n240713 , n240714 , n240715 , 
     n240716 , n240717 , n240718 , n240719 , n240720 , n240721 , n240722 , n240723 , n240724 , n240725 , 
     n240726 , n240727 , n240728 , n240729 , n240730 , n240731 , n240732 , n240733 , n240734 , n240735 , 
     n240736 , n240737 , n240738 , n240739 , n240740 , n240741 , n240742 , n240743 , n240744 , n240745 , 
     n240746 , n240747 , n240748 , n240749 , n240750 , n240751 , n240752 , n240753 , n240754 , n240755 , 
     n240756 , n240757 , n240758 , n240759 , n240760 , n240761 , n240762 , n240763 , n240764 , n240765 , 
     n240766 , n240767 , n240768 , n240769 , n240770 , n240771 , n240772 , n240773 , n240774 , n240775 , 
     n240776 , n240777 , n240778 , n240779 , n240780 , n240781 , n240782 , n240783 , n240784 , n240785 , 
     n240786 , n240787 , n240788 , n240789 , n240790 , n240791 , n240792 , n240793 , n240794 , n240795 , 
     n240796 , n240797 , n240798 , n240799 , n240800 , n240801 , n240802 , n240803 , n240804 , n240805 , 
     n240806 , n240807 , n240808 , n240809 , n240810 , n240811 , n240812 , n240813 , n240814 , n240815 , 
     n240816 , n240817 , n240818 , n240819 , n240820 , n240821 , n240822 , n240823 , n240824 , n240825 , 
     n240826 , n240827 , n240828 , n240829 , n240830 , n240831 , n240832 , n240833 , n240834 , n240835 , 
     n240836 , n240837 , n240838 , n240839 , n240840 , n240841 , n240842 , n240843 , n240844 , n240845 , 
     n240846 , n240847 , n240848 , n240849 , n240850 , n240851 , n240852 , n240853 , n240854 , n240855 , 
     n240856 , n240857 , n240858 , n240859 , n240860 , n240861 , n240862 , n240863 , n240864 , n240865 , 
     n240866 , n240867 , n240868 , n240869 , n240870 , n240871 , n240872 , n240873 , n240874 , n240875 , 
     n240876 , n240877 , n240878 , n240879 , n240880 , n240881 , n240882 , n240883 , n240884 , n240885 , 
     n240886 , n240887 , n240888 , n240889 , n240890 , n240891 , n240892 , n240893 , n240894 , n240895 , 
     n240896 , n240897 , n240898 , n240899 , n240900 , n240901 , n240902 , n240903 , n240904 , n240905 , 
     n240906 , n240907 , n240908 , n240909 , n240910 , n240911 , n240912 , n240913 , n240914 , n240915 , 
     n240916 , n240917 , n240918 , n240919 , n240920 , n240921 , n240922 , n240923 , n240924 , n240925 , 
     n240926 , n240927 , n240928 , n240929 , n240930 , n240931 , n240932 , n240933 , n240934 , n240935 , 
     n240936 , n240937 , n240938 , n240939 , n240940 , n240941 , n240942 , n240943 , n240944 , n240945 , 
     n240946 , n240947 , n240948 , n240949 , n240950 , n240951 , n240952 , n240953 , n240954 , n240955 , 
     n240956 , n240957 , n240958 , n240959 , n240960 , n240961 , n240962 , n240963 , n240964 , n240965 , 
     n240966 , n240967 , n240968 , n240969 , n240970 , n240971 , n240972 , n240973 , n240974 , n240975 , 
     n240976 , n240977 , n240978 , n240979 , n240980 , n240981 , n240982 , n240983 , n240984 , n240985 , 
     n240986 , n240987 , n240988 , n240989 , n240990 , n240991 , n240992 , n240993 , n240994 , n240995 , 
     n240996 , n240997 , n240998 , n240999 , n241000 , n241001 , n241002 , n241003 , n241004 , n241005 , 
     n241006 , n241007 , n241008 , n241009 , n241010 , n241011 , n241012 , n241013 , n241014 , n241015 , 
     n241016 , n241017 , n241018 , n241019 , n241020 , n241021 , n241022 , n241023 , n241024 , n241025 , 
     n241026 , n241027 , n241028 , n241029 , n241030 , n241031 , n241032 , n241033 , n241034 , n241035 , 
     n241036 , n241037 , n241038 , n241039 , n241040 , n241041 , n241042 , n241043 , n241044 , n241045 , 
     n241046 , n241047 , n241048 , n241049 , n241050 , n241051 , n241052 , n241053 , n241054 , n241055 , 
     n241056 , n241057 , n241058 , n241059 , n241060 , n241061 , n241062 , n241063 , n241064 , n241065 , 
     n241066 , n241067 , n241068 , n241069 , n241070 , n241071 , n241072 , n241073 , n241074 , n241075 , 
     n241076 , n241077 , n241078 , n241079 , n241080 , n241081 , n241082 , n241083 , n241084 , n241085 , 
     n241086 , n241087 , n241088 , n241089 , n241090 , n241091 , n241092 , n241093 , n241094 , n241095 , 
     n241096 , n241097 , n241098 , n241099 , n241100 , n241101 , n241102 , n241103 , n241104 , n241105 , 
     n241106 , n241107 , n241108 , n241109 , n241110 , n241111 , n241112 , n241113 , n241114 , n241115 , 
     n241116 , n241117 , n241118 , n241119 , n241120 , n241121 , n241122 , n241123 , n241124 , n241125 , 
     n241126 , n241127 , n241128 , n241129 , n241130 , n241131 , n241132 , n241133 , n241134 , n241135 , 
     n241136 , n241137 , n241138 , n241139 , n241140 , n241141 , n241142 , n241143 , n241144 , n241145 , 
     n241146 , n241147 , n241148 , n241149 , n241150 , n241151 , n241152 , n241153 , n241154 , n241155 , 
     n241156 , n241157 , n241158 , n241159 , n241160 , n241161 , n241162 , n241163 , n241164 , n241165 , 
     n241166 , n241167 , n241168 , n241169 , n241170 , n241171 , n241172 , n241173 , n241174 , n241175 , 
     n241176 , n241177 , n241178 , n241179 , n241180 , n241181 , n241182 , n241183 , n241184 , n241185 , 
     n241186 , n241187 , n241188 , n241189 , n241190 , n241191 , n241192 , n241193 , n241194 , n241195 , 
     n241196 , n241197 , n241198 , n241199 , n241200 , n241201 , n241202 , n241203 , n241204 , n241205 , 
     n241206 , n241207 , n241208 , n241209 , n241210 , n241211 , n241212 , n241213 , n241214 , n241215 , 
     n241216 , n241217 , n241218 , n241219 , n241220 , n241221 , n241222 , n241223 , n241224 , n241225 , 
     n241226 , n241227 , n241228 , n241229 , n241230 , n241231 , n241232 , n241233 , n241234 , n241235 , 
     n241236 , n241237 , n241238 , n241239 , n241240 , n241241 , n241242 , n241243 , n241244 , n241245 , 
     n241246 , n241247 , n241248 , n241249 , n241250 , n241251 , n241252 , n241253 , n241254 , n241255 , 
     n241256 , n241257 , n241258 , n241259 , n241260 , n241261 , n241262 , n241263 , n241264 , n241265 , 
     n241266 , n241267 , n241268 , n241269 , n241270 , n241271 , n241272 , n241273 , n241274 , n241275 , 
     n241276 , n241277 , n241278 , n241279 , n241280 , n241281 , n241282 , n241283 , n241284 , n241285 , 
     n241286 , n241287 , n241288 , n241289 , n241290 , n241291 , n241292 , n241293 , n241294 , n241295 , 
     n241296 , n241297 , n241298 , n241299 , n241300 , n241301 , n241302 , n241303 , n241304 , n241305 , 
     n241306 , n241307 , n241308 , n241309 , n241310 , n241311 , n241312 , n241313 , n241314 , n241315 , 
     n241316 , n241317 , n241318 , n241319 , n241320 , n241321 , n241322 , n241323 , n241324 , n241325 , 
     n241326 , n241327 , n241328 , n241329 , n241330 , n241331 , n241332 , n241333 , n241334 , n241335 , 
     n241336 , n241337 , n241338 , n241339 , n241340 , n241341 , n241342 , n241343 , n241344 , n241345 , 
     n241346 , n241347 , n241348 , n241349 , n241350 , n241351 , n241352 , n241353 , n241354 , n241355 , 
     n241356 , n241357 , n241358 , n241359 , n241360 , n241361 , n241362 , n241363 , n241364 , n241365 , 
     n241366 , n241367 , n241368 , n241369 , n241370 , n241371 , n241372 , n241373 , n241374 , n241375 , 
     n241376 , n241377 , n241378 , n241379 , n241380 , n241381 , n241382 , n241383 , n241384 , n241385 , 
     n241386 , n241387 , n241388 , n241389 , n241390 , n241391 , n241392 , n241393 , n241394 , n241395 , 
     n241396 , n241397 , n241398 , n241399 , n241400 , n241401 , n241402 , n241403 , n241404 , n241405 , 
     n241406 , n241407 , n241408 , n241409 , n241410 , n241411 , n241412 , n241413 , n241414 , n241415 , 
     n241416 , n241417 , n241418 , n241419 , n241420 , n241421 , n241422 , n241423 , n241424 , n241425 , 
     n241426 , n241427 , n241428 , n241429 , n241430 , n241431 , n241432 , n241433 , n241434 , n241435 , 
     n241436 , n241437 , n241438 , n241439 , n241440 , n241441 , n241442 , n241443 , n241444 , n241445 , 
     n241446 , n241447 , n241448 , n241449 , n241450 , n241451 , n241452 , n241453 , n241454 , n241455 , 
     n241456 , n241457 , n241458 , n241459 , n241460 , n241461 , n241462 , n241463 , n241464 , n241465 , 
     n241466 , n241467 , n241468 , n241469 , n241470 , n241471 , n241472 , n241473 , n241474 , n241475 , 
     n241476 , n241477 , n241478 , n241479 , n241480 , n241481 , n241482 , n241483 , n241484 , n241485 , 
     n241486 , n241487 , n241488 , n241489 , n241490 , n241491 , n241492 , n241493 , n241494 , n241495 , 
     n241496 , n241497 , n241498 , n241499 , n241500 , n241501 , n241502 , n241503 , n241504 , n241505 , 
     n241506 , n241507 , n241508 , n241509 , n241510 , n241511 , n241512 , n241513 , n241514 , n241515 , 
     n241516 , n241517 , n241518 , n241519 , n241520 , n241521 , n241522 , n241523 , n241524 , n241525 , 
     n241526 , n241527 , n241528 , n241529 , n241530 , n241531 , n241532 , n241533 , n241534 , n241535 , 
     n241536 , n241537 , n241538 , n241539 , n241540 , n241541 , n241542 , n241543 , n241544 , n241545 , 
     n241546 , n241547 , n241548 , n241549 , n241550 , n241551 , n241552 , n241553 , n241554 , n241555 , 
     n241556 , n241557 , n241558 , n241559 , n241560 , n241561 , n241562 , n241563 , n241564 , n241565 , 
     n241566 , n241567 , n241568 , n241569 , n241570 , n241571 , n241572 , n241573 , n241574 , n241575 , 
     n241576 , n241577 , n241578 , n241579 , n241580 , n241581 , n241582 , n241583 , n241584 , n241585 , 
     n241586 , n241587 , n241588 , n241589 , n241590 , n241591 , n241592 , n241593 , n241594 , n241595 , 
     n241596 , n241597 , n241598 , n241599 , n241600 , n241601 , n241602 , n241603 , n241604 , n241605 , 
     n241606 , n241607 , n241608 , n241609 , n241610 , n241611 , n241612 , n241613 , n241614 , n241615 , 
     n241616 , n241617 , n241618 , n241619 , n241620 , n241621 , n241622 , n241623 , n241624 , n241625 , 
     n241626 , n241627 , n241628 , n241629 , n241630 , n241631 , n241632 , n241633 , n241634 , n241635 , 
     n241636 , n241637 , n241638 , n241639 , n241640 , n241641 , n241642 , n241643 , n241644 , n241645 , 
     n241646 , n241647 , n241648 , n241649 , n241650 , n241651 , n241652 , n241653 , n241654 , n241655 , 
     n241656 , n241657 , n241658 , n241659 , n241660 , n241661 , n241662 , n241663 , n241664 , n241665 , 
     n241666 , n241667 , n241668 , n241669 , n241670 , n241671 , n241672 , n241673 , n241674 , n241675 , 
     n241676 , n241677 , n241678 , n241679 , n241680 , n241681 , n241682 , n241683 , n241684 , n241685 , 
     n241686 , n241687 , n241688 , n241689 , n241690 , n241691 , n241692 , n241693 , n241694 , n241695 , 
     n241696 , n241697 , n241698 , n241699 , n241700 , n241701 , n241702 , n241703 , n241704 , n241705 , 
     n241706 , n241707 , n241708 , n241709 , n241710 , n241711 , n241712 , n241713 , n241714 , n241715 , 
     n241716 , n241717 , n241718 , n241719 , n241720 , n241721 , n241722 , n241723 , n241724 , n241725 , 
     n241726 , n241727 , n241728 , n241729 , n241730 , n241731 , n241732 , n241733 , n241734 , n241735 , 
     n241736 , n241737 , n241738 , n241739 , n241740 , n241741 , n241742 , n241743 , n241744 , n241745 , 
     n241746 , n241747 , n241748 , n241749 , n241750 , n241751 , n241752 , n241753 , n241754 , n241755 , 
     n241756 , n241757 , n241758 , n241759 , n241760 , n241761 , n241762 , n241763 , n241764 , n241765 , 
     n241766 , n241767 , n241768 , n241769 , n241770 , n241771 , n241772 , n241773 , n241774 , n241775 , 
     n241776 , n241777 , n241778 , n241779 , n241780 , n241781 , n241782 , n241783 , n241784 , n241785 , 
     n241786 , n241787 , n241788 , n241789 , n241790 , n241791 , n241792 , n241793 , n241794 , n241795 , 
     n241796 , n241797 , n241798 , n241799 , n241800 , n241801 , n241802 , n241803 , n241804 , n241805 , 
     n241806 , n241807 , n241808 , n241809 , n241810 , n241811 , n241812 , n241813 , n241814 , n241815 , 
     n241816 , n241817 , n241818 , n241819 , n241820 , n241821 , n241822 , n241823 , n241824 , n241825 , 
     n241826 , n241827 , n241828 , n241829 , n241830 , n241831 , n241832 , n241833 , n241834 , n241835 , 
     n241836 , n241837 , n241838 , n241839 , n241840 , n241841 , n241842 , n241843 , n241844 , n241845 , 
     n241846 , n241847 , n241848 , n241849 , n241850 , n241851 , n241852 , n241853 , n241854 , n241855 , 
     n241856 , n241857 , n241858 , n241859 , n241860 , n241861 , n241862 , n241863 , n241864 , n241865 , 
     n241866 , n241867 , n241868 , n241869 , n241870 , n241871 , n241872 , n241873 , n241874 , n241875 , 
     n241876 , n241877 , n241878 , n241879 , n241880 , n241881 , n241882 , n241883 , n241884 , n241885 , 
     n241886 , n241887 , n241888 , n241889 , n241890 , n241891 , n241892 , n241893 , n241894 , n241895 , 
     n241896 , n241897 , n241898 , n241899 , n241900 , n241901 , n241902 , n241903 , n241904 , n241905 , 
     n241906 , n241907 , n241908 , n241909 , n241910 , n241911 , n241912 , n241913 , n241914 , n241915 , 
     n241916 , n241917 , n241918 , n241919 , n241920 , n241921 , n241922 , n241923 , n241924 , n241925 , 
     n241926 , n241927 , n241928 , n241929 , n241930 , n241931 , n241932 , n241933 , n241934 , n241935 , 
     n241936 , n241937 , n241938 , n241939 , n241940 , n241941 , n241942 , n241943 , n241944 , n241945 , 
     n241946 , n241947 , n241948 , n241949 , n241950 , n241951 , n241952 , n241953 , n241954 , n241955 , 
     n241956 , n241957 , n241958 , n241959 , n241960 , n241961 , n241962 , n241963 , n241964 , n241965 , 
     n241966 , n241967 , n241968 , n241969 , n241970 , n241971 , n241972 , n241973 , n241974 , n241975 , 
     n241976 , n241977 , n241978 , n241979 , n241980 , n241981 , n241982 , n241983 , n241984 , n241985 , 
     n241986 , n241987 , n241988 , n241989 , n241990 , n241991 , n241992 , n241993 , n241994 , n241995 , 
     n241996 , n241997 , n241998 , n241999 , n242000 , n242001 , n242002 , n242003 , n242004 , n242005 , 
     n242006 , n242007 , n242008 , n242009 , n242010 , n242011 , n242012 , n242013 , n242014 , n242015 , 
     n242016 , n242017 , n242018 , n242019 , n242020 , n242021 , n242022 , n242023 , n242024 , n242025 , 
     n242026 , n242027 , n242028 , n242029 , n242030 , n242031 , n242032 , n242033 , n242034 , n242035 , 
     n242036 , n242037 , n242038 , n242039 , n242040 , n242041 , n242042 , n242043 , n242044 , n242045 , 
     n242046 , n242047 , n242048 , n242049 , n242050 , n242051 , n242052 , n242053 , n242054 , n242055 , 
     n242056 , n242057 , n242058 , n242059 , n242060 , n242061 , n242062 , n242063 , n242064 , n242065 , 
     n242066 , n242067 , n242068 , n242069 , n242070 , n242071 , n242072 , n242073 , n242074 , n242075 , 
     n242076 , n242077 , n242078 , n242079 , n242080 , n242081 , n242082 , n242083 , n242084 , n242085 , 
     n242086 , n242087 , n242088 , n242089 , n242090 , n242091 , n242092 , n242093 , n242094 , n242095 , 
     n242096 , n242097 , n242098 , n242099 , n242100 , n242101 , n242102 , n242103 , n242104 , n242105 , 
     n242106 , n242107 , n242108 , n242109 , n242110 , n242111 , n242112 , n242113 , n242114 , n242115 , 
     n242116 , n242117 , n242118 , n242119 , n242120 , n242121 , n242122 , n242123 , n242124 , n242125 , 
     n242126 , n242127 , n242128 , n242129 , n242130 , n242131 , n242132 , n242133 , n242134 , n242135 , 
     n242136 , n242137 , n242138 , n242139 , n242140 , n242141 , n242142 , n242143 , n242144 , n242145 , 
     n242146 , n242147 , n242148 , n242149 , n242150 , n242151 , n242152 , n242153 , n242154 , n242155 , 
     n242156 , n242157 , n242158 , n242159 , n242160 , n242161 , n242162 , n242163 , n242164 , n242165 , 
     n242166 , n242167 , n242168 , n242169 , n242170 , n242171 , n242172 , n242173 , n242174 , n242175 , 
     n242176 , n242177 , n242178 , n242179 , n242180 , n242181 , n242182 , n242183 , n242184 , n242185 , 
     n242186 , n242187 , n242188 , n242189 , n242190 , n242191 , n242192 , n242193 , n242194 , n242195 , 
     n242196 , n242197 , n242198 , n242199 , n242200 , n242201 , n242202 , n242203 , n242204 , n242205 , 
     n242206 , n242207 , n242208 , n242209 , n242210 , n242211 , n242212 , n242213 , n242214 , n242215 , 
     n242216 , n242217 , n242218 , n242219 , n242220 , n242221 , n242222 , n242223 , n242224 , n242225 , 
     n242226 , n242227 , n242228 , n242229 , n242230 , n242231 , n242232 , n242233 , n242234 , n242235 , 
     n242236 , n242237 , n242238 , n242239 , n242240 , n242241 , n242242 , n242243 , n242244 , n242245 , 
     n242246 , n242247 , n242248 , n242249 , n242250 , n242251 , n242252 , n242253 , n242254 , n242255 , 
     n242256 , n242257 , n242258 , n242259 , n242260 , n242261 , n242262 , n242263 , n242264 , n242265 , 
     n242266 , n242267 , n242268 , n242269 , n242270 , n242271 , n242272 , n242273 , n242274 , n242275 , 
     n242276 , n242277 , n242278 , n242279 , n242280 , n242281 , n242282 , n242283 , n242284 , n242285 , 
     n242286 , n242287 , n242288 , n242289 , n242290 , n242291 , n242292 , n242293 , n242294 , n242295 , 
     n242296 , n242297 , n242298 , n242299 , n242300 , n242301 , n242302 , n242303 , n242304 , n242305 , 
     n242306 , n242307 , n242308 , n242309 , n242310 , n242311 , n242312 , n242313 , n242314 , n242315 , 
     n242316 , n242317 , n242318 , n242319 , n242320 , n242321 , n242322 , n242323 , n242324 , n242325 , 
     n242326 , n242327 , n242328 , n242329 , n242330 , n242331 , n242332 , n242333 , n242334 , n242335 , 
     n242336 , n242337 , n242338 , n242339 , n242340 , n242341 , n242342 , n242343 , n242344 , n242345 , 
     n242346 , n242347 , n242348 , n242349 , n242350 , n242351 , n242352 , n242353 , n242354 , n242355 , 
     n242356 , n242357 , n242358 , n242359 , n242360 , n242361 , n242362 , n242363 , n242364 , n242365 , 
     n242366 , n242367 , n242368 , n242369 , n242370 , n242371 , n242372 , n242373 , n242374 , n242375 , 
     n242376 , n242377 , n242378 , n242379 , n242380 , n242381 , n242382 , n242383 , n242384 , n242385 , 
     n242386 , n242387 , n242388 , n242389 , n242390 , n242391 , n242392 , n242393 , n242394 , n242395 , 
     n242396 , n242397 , n242398 , n242399 , n242400 , n242401 , n242402 , n242403 , n242404 , n242405 , 
     n242406 , n242407 , n242408 , n242409 , n242410 , n242411 , n242412 , n242413 , n242414 , n242415 , 
     n242416 , n242417 , n242418 , n242419 , n242420 , n242421 , n242422 , n242423 , n242424 , n242425 , 
     n242426 , n242427 , n242428 , n242429 , n242430 , n242431 , n242432 , n242433 , n242434 , n242435 , 
     n242436 , n242437 , n242438 , n242439 , n242440 , n242441 , n242442 , n242443 , n242444 , n242445 , 
     n242446 , n242447 , n242448 , n242449 , n242450 , n242451 , n242452 , n242453 , n242454 , n242455 , 
     n242456 , n242457 , n242458 , n242459 , n242460 , n242461 , n242462 , n242463 , n242464 , n242465 , 
     n242466 , n242467 , n242468 , n242469 , n242470 , n242471 , n242472 , n242473 , n242474 , n242475 , 
     n242476 , n242477 , n242478 , n242479 , n242480 , n242481 , n242482 , n242483 , n242484 , n242485 , 
     n242486 , n242487 , n242488 , n242489 , n242490 , n242491 , n242492 , n242493 , n242494 , n242495 , 
     n242496 , n242497 , n242498 , n242499 , n242500 , n242501 , n242502 , n242503 , n242504 , n242505 , 
     n242506 , n242507 , n242508 , n242509 , n242510 , n242511 , n242512 , n242513 , n242514 , n242515 , 
     n242516 , n242517 , n242518 , n242519 , n242520 , n242521 , n242522 , n242523 , n242524 , n242525 , 
     n242526 , n242527 , n242528 , n242529 , n242530 , n242531 , n242532 , n242533 , n242534 , n242535 , 
     n242536 , n242537 , n242538 , n242539 , n242540 , n242541 , n242542 , n242543 , n242544 , n242545 , 
     n242546 , n242547 , n242548 , n242549 , n242550 , n242551 , n242552 , n242553 , n242554 , n242555 , 
     n242556 , n242557 , n242558 , n242559 , n242560 , n242561 , n242562 , n242563 , n242564 , n242565 , 
     n242566 , n242567 , n242568 , n242569 , n242570 , n242571 , n242572 , n242573 , n242574 , n242575 , 
     n242576 , n242577 , n242578 , n242579 , n242580 , n242581 , n242582 , n242583 , n242584 , n242585 , 
     n242586 , n242587 , n242588 , n242589 , n242590 , n242591 , n242592 , n242593 , n242594 , n242595 , 
     n242596 , n242597 , n242598 , n242599 , n242600 , n242601 , n242602 , n242603 , n242604 , n242605 , 
     n242606 , n242607 , n242608 , n242609 , n242610 , n242611 , n242612 , n242613 , n242614 , n242615 , 
     n242616 , n242617 , n242618 , n242619 , n242620 , n242621 , n242622 , n242623 , n242624 , n242625 , 
     n242626 , n242627 , n242628 , n242629 , n242630 , n242631 , n242632 , n242633 , n242634 , n242635 , 
     n242636 , n242637 , n242638 , n242639 , n242640 , n242641 , n242642 , n242643 , n242644 , n242645 , 
     n242646 , n242647 , n242648 , n242649 , n242650 , n242651 , n242652 , n242653 , n242654 , n242655 , 
     n242656 , n242657 , n242658 , n242659 , n242660 , n242661 , n242662 , n242663 , n242664 , n242665 , 
     n242666 , n242667 , n242668 , n242669 , n242670 , n242671 , n242672 , n242673 , n242674 , n242675 , 
     n242676 , n242677 , n242678 , n242679 , n242680 , n242681 , n242682 , n242683 , n242684 , n242685 , 
     n242686 , n242687 , n242688 , n242689 , n242690 , n242691 , n242692 , n242693 , n242694 , n242695 , 
     n242696 , n242697 , n242698 , n242699 , n242700 , n242701 , n242702 , n242703 , n242704 , n242705 , 
     n242706 , n242707 , n242708 , n242709 , n242710 , n242711 , n242712 , n242713 , n242714 , n242715 , 
     n242716 , n242717 , n242718 , n242719 , n242720 , n242721 , n242722 , n242723 , n242724 , n242725 , 
     n242726 , n242727 , n242728 , n242729 , n242730 , n242731 , n242732 , n242733 , n242734 , n242735 , 
     n242736 , n242737 , n242738 , n242739 , n242740 , n242741 , n242742 , n242743 , n242744 , n242745 , 
     n242746 , n242747 , n242748 , n242749 , n242750 , n242751 , n242752 , n242753 , n242754 , n242755 , 
     n242756 , n242757 , n242758 , n242759 , n242760 , n242761 , n242762 , n242763 , n242764 , n242765 , 
     n242766 , n242767 , n242768 , n242769 , n242770 , n242771 , n242772 , n242773 , n242774 , n242775 , 
     n242776 , n242777 , n242778 , n242779 , n242780 , n242781 , n242782 , n242783 , n242784 , n242785 , 
     n242786 , n242787 , n242788 , n242789 , n242790 , n242791 , n242792 , n242793 , n242794 , n242795 , 
     n242796 , n242797 , n242798 , n242799 , n242800 , n242801 , n242802 , n242803 , n242804 , n242805 , 
     n242806 , n242807 , n242808 , n242809 , n242810 , n242811 , n242812 , n242813 , n242814 , n242815 , 
     n242816 , n242817 , n242818 , n242819 , n242820 , n242821 , n242822 , n242823 , n242824 , n242825 , 
     n242826 , n242827 , n242828 , n242829 , n242830 , n242831 , n242832 , n242833 , n242834 , n242835 , 
     n242836 , n242837 , n242838 , n242839 , n242840 , n242841 , n242842 , n242843 , n242844 , n242845 , 
     n242846 , n242847 , n242848 , n242849 , n242850 , n242851 , n242852 , n242853 , n242854 , n242855 , 
     n242856 , n242857 , n242858 , n242859 , n242860 , n242861 , n242862 , n242863 , n242864 , n242865 , 
     n242866 , n242867 , n242868 , n242869 , n242870 , n242871 , n242872 , n242873 , n242874 , n242875 , 
     n242876 , n242877 , n242878 , n242879 , n242880 , n242881 , n242882 , n242883 , n242884 , n242885 , 
     n242886 , n242887 , n242888 , n242889 , n242890 , n242891 , n242892 , n242893 , n242894 , n242895 , 
     n242896 , n242897 , n242898 , n242899 , n242900 , n242901 , n242902 , n242903 , n242904 , n242905 , 
     n242906 , n242907 , n242908 , n242909 , n242910 , n242911 , n242912 , n242913 , n242914 , n242915 , 
     n242916 , n242917 , n242918 , n242919 , n242920 , n242921 , n242922 , n242923 , n242924 , n242925 , 
     n242926 , n242927 , n242928 , n242929 , n242930 , n242931 , n242932 , n242933 , n242934 , n242935 , 
     n242936 , n242937 , n242938 , n242939 , n242940 , n242941 , n242942 , n242943 , n242944 , n242945 , 
     n242946 , n242947 , n242948 , n242949 , n242950 , n242951 , n242952 , n242953 , n242954 , n242955 , 
     n242956 , n242957 , n242958 , n242959 , n242960 , n242961 , n242962 , n242963 , n242964 , n242965 , 
     n242966 , n242967 , n242968 , n242969 , n242970 , n242971 , n242972 , n242973 , n242974 , n242975 , 
     n242976 , n242977 , n242978 , n242979 , n242980 , n242981 , n242982 , n242983 , n242984 , n242985 , 
     n242986 , n242987 , n242988 , n242989 , n242990 , n242991 , n242992 , n242993 , n242994 , n242995 , 
     n242996 , n242997 , n242998 , n242999 , n243000 , n243001 , n243002 , n243003 , n243004 , n243005 , 
     n243006 , n243007 , n243008 , n243009 , n243010 , n243011 , n243012 , n243013 , n243014 , n243015 , 
     n243016 , n243017 , n243018 , n243019 , n243020 , n243021 , n243022 , n243023 , n243024 , n243025 , 
     n243026 , n243027 , n243028 , n243029 , n243030 , n243031 , n243032 , n243033 , n243034 , n243035 , 
     n243036 , n243037 , n243038 , n243039 , n243040 , n243041 , n243042 , n243043 , n243044 , n243045 , 
     n243046 , n243047 , n243048 , n243049 , n243050 , n243051 , n243052 , n243053 , n243054 , n243055 , 
     n243056 , n243057 , n243058 , n243059 , n243060 , n243061 , n243062 , n243063 , n243064 , n243065 , 
     n243066 , n243067 , n243068 , n243069 , n243070 , n243071 , n243072 , n243073 , n243074 , n243075 , 
     n243076 , n243077 , n243078 , n243079 , n243080 , n243081 , n243082 , n243083 , n243084 , n243085 , 
     n243086 , n243087 , n243088 , n243089 , n243090 , n243091 , n243092 , n243093 , n243094 , n243095 , 
     n243096 , n243097 , n243098 , n243099 , n243100 , n243101 , n243102 , n243103 , n243104 , n243105 , 
     n243106 , n243107 , n243108 , n243109 , n243110 , n243111 , n243112 , n243113 , n243114 , n243115 , 
     n243116 , n243117 , n243118 , n243119 , n243120 , n243121 , n243122 , n243123 , n243124 , n243125 , 
     n243126 , n243127 , n243128 , n243129 , n243130 , n243131 , n243132 , n243133 , n243134 , n243135 , 
     n243136 , n243137 , n243138 , n243139 , n243140 , n243141 , n243142 , n243143 , n243144 , n243145 , 
     n243146 , n243147 , n243148 , n243149 , n243150 , n243151 , n243152 , n243153 , n243154 , n243155 , 
     n243156 , n243157 , n243158 , n243159 , n243160 , n243161 , n243162 , n243163 , n243164 , n243165 , 
     n243166 , n243167 , n243168 , n243169 , n243170 , n243171 , n243172 , n243173 , n243174 , n243175 , 
     n243176 , n243177 , n243178 , n243179 , n243180 , n243181 , n243182 , n243183 , n243184 , n243185 , 
     n243186 , n243187 , n243188 , n243189 , n243190 , n243191 , n243192 , n243193 , n243194 , n243195 , 
     n243196 , n243197 , n243198 , n243199 , n243200 , n243201 , n243202 , n243203 , n243204 , n243205 , 
     n243206 , n243207 , n243208 , n243209 , n243210 , n243211 , n243212 , n243213 , n243214 , n243215 , 
     n243216 , n243217 , n243218 , n243219 , n243220 , n243221 , n243222 , n243223 , n243224 , n243225 , 
     n243226 , n243227 , n243228 , n243229 , n243230 , n243231 , n243232 , n243233 , n243234 , n243235 , 
     n243236 , n243237 , n243238 , n243239 , n243240 , n243241 , n243242 , n243243 , n243244 , n243245 , 
     n243246 , n243247 , n243248 , n243249 , n243250 , n243251 , n243252 , n243253 , n243254 , n243255 , 
     n243256 , n243257 , n243258 , n243259 , n243260 , n243261 , n243262 , n243263 , n243264 , n243265 , 
     n243266 , n243267 , n243268 , n243269 , n243270 , n243271 , n243272 , n243273 , n243274 , n243275 , 
     n243276 , n243277 , n243278 , n243279 , n243280 , n243281 , n243282 , n243283 , n243284 , n243285 , 
     n243286 , n243287 , n243288 , n243289 , n243290 , n243291 , n243292 , n243293 , n243294 , n243295 , 
     n243296 , n243297 , n243298 , n243299 , n243300 , n243301 , n243302 , n243303 , n243304 , n243305 , 
     n243306 , n243307 , n243308 , n243309 , n243310 , n243311 , n243312 , n243313 , n243314 , n243315 , 
     n243316 , n243317 , n243318 , n243319 , n243320 , n243321 , n243322 , n243323 , n243324 , n243325 , 
     n243326 , n243327 , n243328 , n243329 , n243330 , n243331 , n243332 , n243333 , n243334 , n243335 , 
     n243336 , n243337 , n243338 , n243339 , n243340 , n243341 , n243342 , n243343 , n243344 , n243345 , 
     n243346 , n243347 , n243348 , n243349 , n243350 , n243351 , n243352 , n243353 , n243354 , n243355 , 
     n243356 , n243357 , n243358 , n243359 , n243360 , n243361 , n243362 , n243363 , n243364 , n243365 , 
     n243366 , n243367 , n243368 , n243369 , n243370 , n243371 , n243372 , n243373 , n243374 , n243375 , 
     n243376 , n243377 , n243378 , n243379 , n243380 , n243381 , n243382 , n243383 , n243384 , n243385 , 
     n243386 , n243387 , n243388 , n243389 , n243390 , n243391 , n243392 , n243393 , n243394 , n243395 , 
     n243396 , n243397 , n243398 , n243399 , n243400 , n243401 , n243402 , n243403 , n243404 , n243405 , 
     n243406 , n243407 , n243408 , n243409 , n243410 , n243411 , n243412 , n243413 , n243414 , n243415 , 
     n243416 , n243417 , n243418 , n243419 , n243420 , n243421 , n243422 , n243423 , n243424 , n243425 , 
     n243426 , n243427 , n243428 , n243429 , n243430 , n243431 , n243432 , n243433 , n243434 , n243435 , 
     n243436 , n243437 , n243438 , n243439 , n243440 , n243441 , n243442 , n243443 , n243444 , n243445 , 
     n243446 , n243447 , n243448 , n243449 , n243450 , n243451 , n243452 , n243453 , n243454 , n243455 , 
     n243456 , n243457 , n243458 , n243459 , n243460 , n243461 , n243462 , n243463 , n243464 , n243465 , 
     n243466 , n243467 , n243468 , n243469 , n243470 , n243471 , n243472 , n243473 , n243474 , n243475 , 
     n243476 , n243477 , n243478 , n243479 , n243480 , n243481 , n243482 , n243483 , n243484 , n243485 , 
     n243486 , n243487 , n243488 , n243489 , n243490 , n243491 , n243492 , n243493 , n243494 , n243495 , 
     n243496 , n243497 , n243498 , n243499 , n243500 , n243501 , n243502 , n243503 , n243504 , n243505 , 
     n243506 , n243507 , n243508 , n243509 , n243510 , n243511 , n243512 , n243513 , n243514 , n243515 , 
     n243516 , n243517 , n243518 , n243519 , n243520 , n243521 , n243522 , n243523 , n243524 , n243525 , 
     n243526 , n243527 , n243528 , n243529 , n243530 , n243531 , n243532 , n243533 , n243534 , n243535 , 
     n243536 , n243537 , n243538 , n243539 , n243540 , n243541 , n243542 , n243543 , n243544 , n243545 , 
     n243546 , n243547 , n243548 , n243549 , n243550 , n243551 , n243552 , n243553 , n243554 , n243555 , 
     n243556 , n243557 , n243558 , n243559 , n243560 , n243561 , n243562 , n243563 , n243564 , n243565 , 
     n243566 , n243567 , n243568 , n243569 , n243570 , n243571 , n243572 , n243573 , n243574 , n243575 , 
     n243576 , n243577 , n243578 , n243579 , n243580 , n243581 , n243582 , n243583 , n243584 , n243585 , 
     n243586 , n243587 , n243588 , n243589 , n243590 , n243591 , n243592 , n243593 , n243594 , n243595 , 
     n243596 , n243597 , n243598 , n243599 , n243600 , n243601 , n243602 , n243603 , n243604 , n243605 , 
     n243606 , n243607 , n243608 , n243609 , n243610 , n243611 , n243612 , n243613 , n243614 , n243615 , 
     n243616 , n243617 , n243618 , n243619 , n243620 , n243621 , n243622 , n243623 , n243624 , n243625 , 
     n243626 , n243627 , n243628 , n243629 , n243630 , n243631 , n243632 , n243633 , n243634 , n243635 , 
     n243636 , n243637 , n243638 , n243639 , n243640 , n243641 , n243642 , n243643 , n243644 , n243645 , 
     n243646 , n243647 , n243648 , n243649 , n243650 , n243651 , n243652 , n243653 , n243654 , n243655 , 
     n243656 , n243657 , n243658 , n243659 , n243660 , n243661 , n243662 , n243663 , n243664 , n243665 , 
     n243666 , n243667 , n243668 , n243669 , n243670 , n243671 , n243672 , n243673 , n243674 , n243675 , 
     n243676 , n243677 , n243678 , n243679 , n243680 , n243681 , n243682 , n243683 , n243684 , n243685 , 
     n243686 , n243687 , n243688 , n243689 , n243690 , n243691 , n243692 , n243693 , n243694 , n243695 , 
     n243696 , n243697 , n243698 , n243699 , n243700 , n243701 , n243702 , n243703 , n243704 , n243705 , 
     n243706 , n243707 , n243708 , n243709 , n243710 , n243711 , n243712 , n243713 , n243714 , n243715 , 
     n243716 , n243717 , n243718 , n243719 , n243720 , n243721 , n243722 , n243723 , n243724 , n243725 , 
     n243726 , n243727 , n243728 , n243729 , n243730 , n243731 , n243732 , n243733 , n243734 , n243735 , 
     n243736 , n243737 , n243738 , n243739 , n243740 , n243741 , n243742 , n243743 , n243744 , n243745 , 
     n243746 , n243747 , n243748 , n243749 , n243750 , n243751 , n243752 , n243753 , n243754 , n243755 , 
     n243756 , n243757 , n243758 , n243759 , n243760 , n243761 , n243762 , n243763 , n243764 , n243765 , 
     n243766 , n243767 , n243768 , n243769 , n243770 , n243771 , n243772 , n243773 , n243774 , n243775 , 
     n243776 , n243777 , n243778 , n243779 , n243780 , n243781 , n243782 , n243783 , n243784 , n243785 , 
     n243786 , n243787 , n243788 , n243789 , n243790 , n243791 , n243792 , n243793 , n243794 , n243795 , 
     n243796 , n243797 , n243798 , n243799 , n243800 , n243801 , n243802 , n243803 , n243804 , n243805 , 
     n243806 , n243807 , n243808 , n243809 , n243810 , n243811 , n243812 , n243813 , n243814 , n243815 , 
     n243816 , n243817 , n243818 , n243819 , n243820 , n243821 , n243822 , n243823 , n243824 , n243825 , 
     n243826 , n243827 , n243828 , n243829 , n243830 , n243831 , n243832 , n243833 , n243834 , n243835 , 
     n243836 , n243837 , n243838 , n243839 , n243840 , n243841 , n243842 , n243843 , n243844 , n243845 , 
     n243846 , n243847 , n243848 , n243849 , n243850 , n243851 , n243852 , n243853 , n243854 , n243855 , 
     n243856 , n243857 , n243858 , n243859 , n243860 , n243861 , n243862 , n243863 , n243864 , n243865 , 
     n243866 , n243867 , n243868 , n243869 , n243870 , n243871 , n243872 , n243873 , n243874 , n243875 , 
     n243876 , n243877 , n243878 , n243879 , n243880 , n243881 , n243882 , n243883 , n243884 , n243885 , 
     n243886 , n243887 , n243888 , n243889 , n243890 , n243891 , n243892 , n243893 , n243894 , n243895 , 
     n243896 , n243897 , n243898 , n243899 , n243900 , n243901 , n243902 , n243903 , n243904 , n243905 , 
     n243906 , n243907 , n243908 , n243909 , n243910 , n243911 , n243912 , n243913 , n243914 , n243915 , 
     n243916 , n243917 , n243918 , n243919 , n243920 , n243921 , n243922 , n243923 , n243924 , n243925 , 
     n243926 , n243927 , n243928 , n243929 , n243930 , n243931 , n243932 , n243933 , n243934 , n243935 , 
     n243936 , n243937 , n243938 , n243939 , n243940 , n243941 , n243942 , n243943 , n243944 , n243945 , 
     n243946 , n243947 , n243948 , n243949 , n243950 , n243951 , n243952 , n243953 , n243954 , n243955 , 
     n243956 , n243957 , n243958 , n243959 , n243960 , n243961 , n243962 , n243963 , n243964 , n243965 , 
     n243966 , n243967 , n243968 , n243969 , n243970 , n243971 , n243972 , n243973 , n243974 , n243975 , 
     n243976 , n243977 , n243978 , n243979 , n243980 , n243981 , n243982 , n243983 , n243984 , n243985 , 
     n243986 , n243987 , n243988 , n243989 , n243990 , n243991 , n243992 , n243993 , n243994 , n243995 , 
     n243996 , n243997 , n243998 , n243999 , n244000 , n244001 , n244002 , n244003 , n244004 , n244005 , 
     n244006 , n244007 , n244008 , n244009 , n244010 , n244011 , n244012 , n244013 , n244014 , n244015 , 
     n244016 , n244017 , n244018 , n244019 , n244020 , n244021 , n244022 , n244023 , n244024 , n244025 , 
     n244026 , n244027 , n244028 , n244029 , n244030 , n244031 , n244032 , n244033 , n244034 , n244035 , 
     n244036 , n244037 , n244038 , n244039 , n244040 , n244041 , n244042 , n244043 , n244044 , n244045 , 
     n244046 , n244047 , n244048 , n244049 , n244050 , n244051 , n244052 , n244053 , n244054 , n244055 , 
     n244056 , n244057 , n244058 , n244059 , n244060 , n244061 , n244062 , n244063 , n244064 , n244065 , 
     n244066 , n244067 , n244068 , n244069 , n244070 , n244071 , n244072 , n244073 , n244074 , n244075 , 
     n244076 , n244077 , n244078 , n244079 , n244080 , n244081 , n244082 , n244083 , n244084 , n244085 , 
     n244086 , n244087 , n244088 , n244089 , n244090 , n244091 , n244092 , n244093 , n244094 , n244095 , 
     n244096 , n244097 , n244098 , n244099 , n244100 , n244101 , n244102 , n244103 , n244104 , n244105 , 
     n244106 , n244107 , n244108 , n244109 , n244110 , n244111 , n244112 , n244113 , n244114 , n244115 , 
     n244116 , n244117 , n244118 , n244119 , n244120 , n244121 , n244122 , n244123 , n244124 , n244125 , 
     n244126 , n244127 , n244128 , n244129 , n244130 , n244131 , n244132 , n244133 , n244134 , n244135 , 
     n244136 , n244137 , n244138 , n244139 , n244140 , n244141 , n244142 , n244143 , n244144 , n244145 , 
     n244146 , n244147 , n244148 , n244149 , n244150 , n244151 , n244152 , n244153 , n244154 , n244155 , 
     n244156 , n244157 , n244158 , n244159 , n244160 , n244161 , n244162 , n244163 , n244164 , n244165 , 
     n244166 , n244167 , n244168 , n244169 , n244170 , n244171 , n244172 , n244173 , n244174 , n244175 , 
     n244176 , n244177 , n244178 , n244179 , n244180 , n244181 , n244182 , n244183 , n244184 , n244185 , 
     n244186 , n244187 , n244188 , n244189 , n244190 , n244191 , n244192 , n244193 , n244194 , n244195 , 
     n244196 , n244197 , n244198 , n244199 , n244200 , n244201 , n244202 , n244203 , n244204 , n244205 , 
     n244206 , n244207 , n244208 , n244209 , n244210 , n244211 , n244212 , n244213 , n244214 , n244215 , 
     n244216 , n244217 , n244218 , n244219 , n244220 , n244221 , n244222 , n244223 , n244224 , n244225 , 
     n244226 , n244227 , n244228 , n244229 , n244230 , n244231 , n244232 , n244233 , n244234 , n244235 , 
     n244236 , n244237 , n244238 , n244239 , n244240 , n244241 , n244242 , n244243 , n244244 , n244245 , 
     n244246 , n244247 , n244248 , n244249 , n244250 , n244251 , n244252 , n244253 , n244254 , n244255 , 
     n244256 , n244257 , n244258 , n244259 , n244260 , n244261 , n244262 , n244263 , n244264 , n244265 , 
     n244266 , n244267 , n244268 , n244269 , n244270 , n244271 , n244272 , n244273 , n244274 , n244275 , 
     n244276 , n244277 , n244278 , n244279 , n244280 , n244281 , n244282 , n244283 , n244284 , n244285 , 
     n244286 , n244287 , n244288 , n244289 , n244290 , n244291 , n244292 , n244293 , n244294 , n244295 , 
     n244296 , n244297 , n244298 , n244299 , n244300 , n244301 , n244302 , n244303 , n244304 , n244305 , 
     n244306 , n244307 , n244308 , n244309 , n244310 , n244311 , n244312 , n244313 , n244314 , n244315 , 
     n244316 , n244317 , n244318 , n244319 , n244320 , n244321 , n244322 , n244323 , n244324 , n244325 , 
     n244326 , n244327 , n244328 , n244329 , n244330 , n244331 , n244332 , n244333 , n244334 , n244335 , 
     n244336 , n244337 , n244338 , n244339 , n244340 , n244341 , n244342 , n244343 , n244344 , n244345 , 
     n244346 , n244347 , n244348 , n244349 , n244350 , n244351 , n244352 , n244353 , n244354 , n244355 , 
     n244356 , n244357 , n244358 , n244359 , n244360 , n244361 , n244362 , n244363 , n244364 , n244365 , 
     n244366 , n244367 , n244368 , n244369 , n244370 , n244371 , n244372 , n244373 , n244374 , n244375 , 
     n244376 , n244377 , n244378 , n244379 , n244380 , n244381 , n244382 , n244383 , n244384 , n244385 , 
     n244386 , n244387 , n244388 , n244389 , n244390 , n244391 , n244392 , n244393 , n244394 , n244395 , 
     n244396 , n244397 , n244398 , n244399 , n244400 , n244401 , n244402 , n244403 , n244404 , n244405 , 
     n244406 , n244407 , n244408 , n244409 , n244410 , n244411 , n244412 , n244413 , n244414 , n244415 , 
     n244416 , n244417 , n244418 , n244419 , n244420 , n244421 , n244422 , n244423 , n244424 , n244425 , 
     n244426 , n244427 , n244428 , n244429 , n244430 , n244431 , n244432 , n244433 , n244434 , n244435 , 
     n244436 , n244437 , n244438 , n244439 , n244440 , n244441 , n244442 , n244443 , n244444 , n244445 , 
     n244446 , n244447 , n244448 , n244449 , n244450 , n244451 , n244452 , n244453 , n244454 , n244455 , 
     n244456 , n244457 , n244458 , n244459 , n244460 , n244461 , n244462 , n244463 , n244464 , n244465 , 
     n244466 , n244467 , n244468 , n244469 , n244470 , n244471 , n244472 , n244473 , n244474 , n244475 , 
     n244476 , n244477 , n244478 , n244479 , n244480 , n244481 , n244482 , n244483 , n244484 , n244485 , 
     n244486 , n244487 , n244488 , n244489 , n244490 , n244491 , n244492 , n244493 , n244494 , n244495 , 
     n244496 , n244497 , n244498 , n244499 , n244500 , n244501 , n244502 , n244503 , n244504 , n244505 , 
     n244506 , n244507 , n244508 , n244509 , n244510 , n244511 , n244512 , n244513 , n244514 , n244515 , 
     n244516 , n244517 , n244518 , n244519 , n244520 , n244521 , n244522 , n244523 , n244524 , n244525 , 
     n244526 , n244527 , n244528 , n244529 , n244530 , n244531 , n244532 , n244533 , n244534 , n244535 , 
     n244536 , n244537 , n244538 , n244539 , n244540 , n244541 , n244542 , n244543 , n244544 , n244545 , 
     n244546 , n244547 , n244548 , n244549 , n244550 , n244551 , n244552 , n244553 , n244554 , n244555 , 
     n244556 , n244557 , n244558 , n244559 , n244560 , n244561 , n244562 , n244563 , n244564 , n244565 , 
     n244566 , n244567 , n244568 , n244569 , n244570 , n244571 , n244572 , n244573 , n244574 , n244575 , 
     n244576 , n244577 , n244578 , n244579 , n244580 , n244581 , n244582 , n244583 , n244584 , n244585 , 
     n244586 , n244587 , n244588 , n244589 , n244590 , n244591 , n244592 , n244593 , n244594 , n244595 , 
     n244596 , n244597 , n244598 , n244599 , n244600 , n244601 , n244602 , n244603 , n244604 , n244605 , 
     n244606 , n244607 , n244608 , n244609 , n244610 , n244611 , n244612 , n244613 , n244614 , n244615 , 
     n244616 , n244617 , n244618 , n244619 , n244620 , n244621 , n244622 , n244623 , n244624 , n244625 , 
     n244626 , n244627 , n244628 , n244629 , n244630 , n244631 , n244632 , n244633 , n244634 , n244635 , 
     n244636 , n244637 , n244638 , n244639 , n244640 , n244641 , n244642 , n244643 , n244644 , n244645 , 
     n244646 , n244647 , n244648 , n244649 , n244650 , n244651 , n244652 , n244653 , n244654 , n244655 , 
     n244656 , n244657 , n244658 , n244659 , n244660 , n244661 , n244662 , n244663 , n244664 , n244665 , 
     n244666 , n244667 , n244668 , n244669 , n244670 , n244671 , n244672 , n244673 , n244674 , n244675 , 
     n244676 , n244677 , n244678 , n244679 , n244680 , n244681 , n244682 , n244683 , n244684 , n244685 , 
     n244686 , n244687 , n244688 , n244689 , n244690 , n244691 , n244692 , n244693 , n244694 , n244695 , 
     n244696 , n244697 , n244698 , n244699 , n244700 , n244701 , n244702 , n244703 , n244704 , n244705 , 
     n244706 , n244707 , n244708 , n244709 , n244710 , n244711 , n244712 , n244713 , n244714 , n244715 , 
     n244716 , n244717 , n244718 , n244719 , n244720 , n244721 , n244722 , n244723 , n244724 , n244725 , 
     n244726 , n244727 , n244728 , n244729 , n244730 , n244731 , n244732 , n244733 , n244734 , n244735 , 
     n244736 , n244737 , n244738 , n244739 , n244740 , n244741 , n244742 , n244743 , n244744 , n244745 , 
     n244746 , n244747 , n244748 , n244749 , n244750 , n244751 , n244752 , n244753 , n244754 , n244755 , 
     n244756 , n244757 , n244758 , n244759 , n244760 , n244761 , n244762 , n244763 , n244764 , n244765 , 
     n244766 , n244767 , n244768 , n244769 , n244770 , n244771 , n244772 , n244773 , n244774 , n244775 , 
     n244776 , n244777 , n244778 , n244779 , n244780 , n244781 , n244782 , n244783 , n244784 , n244785 , 
     n244786 , n244787 , n244788 , n244789 , n244790 , n244791 , n244792 , n244793 , n244794 , n244795 , 
     n244796 , n244797 , n244798 , n244799 , n244800 , n244801 , n244802 , n244803 , n244804 , n244805 , 
     n244806 , n244807 , n244808 , n244809 , n244810 , n244811 , n244812 , n244813 , n244814 , n244815 , 
     n244816 , n244817 , n244818 , n244819 , n244820 , n244821 , n244822 , n244823 , n244824 , n244825 , 
     n244826 , n244827 , n244828 , n244829 , n244830 , n244831 , n244832 , n244833 , n244834 , n244835 , 
     n244836 , n244837 , n244838 , n244839 , n244840 , n244841 , n244842 , n244843 , n244844 , n244845 , 
     n244846 , n244847 , n244848 , n244849 , n244850 , n244851 , n244852 , n244853 , n244854 , n244855 , 
     n244856 , n244857 , n244858 , n244859 , n244860 , n244861 , n244862 , n244863 , n244864 , n244865 , 
     n244866 , n244867 , n244868 , n244869 , n244870 , n244871 , n244872 , n244873 , n244874 , n244875 , 
     n244876 , n244877 , n244878 , n244879 , n244880 , n244881 , n244882 , n244883 , n244884 , n244885 , 
     n244886 , n244887 , n244888 , n244889 , n244890 , n244891 , n244892 , n244893 , n244894 , n244895 , 
     n244896 , n244897 , n244898 , n244899 , n244900 , n244901 , n244902 , n244903 , n244904 , n244905 , 
     n244906 , n244907 , n244908 , n244909 , n244910 , n244911 , n244912 , n244913 , n244914 , n244915 , 
     n244916 , n244917 , n244918 , n244919 , n244920 , n244921 , n244922 , n244923 , n244924 , n244925 , 
     n244926 , n244927 , n244928 , n244929 , n244930 , n244931 , n244932 , n244933 , n244934 , n244935 , 
     n244936 , n244937 , n244938 , n244939 , n244940 , n244941 , n244942 , n244943 , n244944 , n244945 , 
     n244946 , n244947 , n244948 , n244949 , n244950 , n244951 , n244952 , n244953 , n244954 , n244955 , 
     n244956 , n244957 , n244958 , n244959 , n244960 , n244961 , n244962 , n244963 , n244964 , n244965 , 
     n244966 , n244967 , n244968 , n244969 , n244970 , n244971 , n244972 , n244973 , n244974 , n244975 , 
     n244976 , n244977 , n244978 , n244979 , n244980 , n244981 , n244982 , n244983 , n244984 , n244985 , 
     n244986 , n244987 , n244988 , n244989 , n244990 , n244991 , n244992 , n244993 , n244994 , n244995 , 
     n244996 , n244997 , n244998 , n244999 , n245000 , n245001 , n245002 , n245003 , n245004 , n245005 , 
     n245006 , n245007 , n245008 , n245009 , n245010 , n245011 , n245012 , n245013 , n245014 , n245015 , 
     n245016 , n245017 , n245018 , n245019 , n245020 , n245021 , n245022 , n245023 , n245024 , n245025 , 
     n245026 , n245027 , n245028 , n245029 , n245030 , n245031 , n245032 , n245033 , n245034 , n245035 , 
     n245036 , n245037 , n245038 , n245039 , n245040 , n245041 , n245042 , n245043 , n245044 , n245045 , 
     n245046 , n245047 , n245048 , n245049 , n245050 , n245051 , n245052 , n245053 , n245054 , n245055 , 
     n245056 , n245057 , n245058 , n245059 , n245060 , n245061 , n245062 , n245063 , n245064 , n245065 , 
     n245066 , n245067 , n245068 , n245069 , n245070 , n245071 , n245072 , n245073 , n245074 , n245075 , 
     n245076 , n245077 , n245078 , n245079 , n245080 , n245081 , n245082 , n245083 , n245084 , n245085 , 
     n245086 , n245087 , n245088 , n245089 , n245090 , n245091 , n245092 , n245093 , n245094 , n245095 , 
     n245096 , n245097 , n245098 , n245099 , n245100 , n245101 , n245102 , n245103 , n245104 , n245105 , 
     n245106 , n245107 , n245108 , n245109 , n245110 , n245111 , n245112 , n245113 , n245114 , n245115 , 
     n245116 , n245117 , n245118 , n245119 , n245120 , n245121 , n245122 , n245123 , n245124 , n245125 , 
     n245126 , n245127 , n245128 , n245129 , n245130 , n245131 , n245132 , n245133 , n245134 , n245135 , 
     n245136 , n245137 , n245138 , n245139 , n245140 , n245141 , n245142 , n245143 , n245144 , n245145 , 
     n245146 , n245147 , n245148 , n245149 , n245150 , n245151 , n245152 , n245153 , n245154 , n245155 , 
     n245156 , n245157 , n245158 , n245159 , n245160 , n245161 , n245162 , n245163 , n245164 , n245165 , 
     n245166 , n245167 , n245168 , n245169 , n245170 , n245171 , n245172 , n245173 , n245174 , n245175 , 
     n245176 , n245177 , n245178 , n245179 , n245180 , n245181 , n245182 , n245183 , n245184 , n245185 , 
     n245186 , n245187 , n245188 , n245189 , n245190 , n245191 , n245192 , n245193 , n245194 , n245195 , 
     n245196 , n245197 , n245198 , n245199 , n245200 , n245201 , n245202 , n245203 , n245204 , n245205 , 
     n245206 , n245207 , n245208 , n245209 , n245210 , n245211 , n245212 , n245213 , n245214 , n245215 , 
     n245216 , n245217 , n245218 , n245219 , n245220 , n245221 , n245222 , n245223 , n245224 , n245225 , 
     n245226 , n245227 , n245228 , n245229 , n245230 , n245231 , n245232 , n245233 , n245234 , n245235 , 
     n245236 , n245237 , n245238 , n245239 , n245240 , n245241 , n245242 , n245243 , n245244 , n245245 , 
     n245246 , n245247 , n245248 , n245249 , n245250 , n245251 , n245252 , n245253 , n245254 , n245255 , 
     n245256 , n245257 , n245258 , n245259 , n245260 , n245261 , n245262 , n245263 , n245264 , n245265 , 
     n245266 , n245267 , n245268 , n245269 , n245270 , n245271 , n245272 , n245273 , n245274 , n245275 , 
     n245276 , n245277 , n245278 , n245279 , n245280 , n245281 , n245282 , n245283 , n245284 , n245285 , 
     n245286 , n245287 , n245288 , n245289 , n245290 , n245291 , n245292 , n245293 , n245294 , n245295 , 
     n245296 , n245297 , n245298 , n245299 , n245300 , n245301 , n245302 , n245303 , n245304 , n245305 , 
     n245306 , n245307 , n245308 , n245309 , n245310 , n245311 , n245312 , n245313 , n245314 , n245315 , 
     n245316 , n245317 , n245318 , n245319 , n245320 , n245321 , n245322 , n245323 , n245324 , n245325 , 
     n245326 , n245327 , n245328 , n245329 , n245330 , n245331 , n245332 , n245333 , n245334 , n245335 , 
     n245336 , n245337 , n245338 , n245339 , n245340 , n245341 , n245342 , n245343 , n245344 , n245345 , 
     n245346 , n245347 , n245348 , n245349 , n245350 , n245351 , n245352 , n245353 , n245354 , n245355 , 
     n245356 , n245357 , n245358 , n245359 , n245360 , n245361 , n245362 , n245363 , n245364 , n245365 , 
     n245366 , n245367 , n245368 , n245369 , n245370 , n245371 , n245372 , n245373 , n245374 , n245375 , 
     n245376 , n245377 , n245378 , n245379 , n245380 , n245381 , n245382 , n245383 , n245384 , n245385 , 
     n245386 , n245387 , n245388 , n245389 , n245390 , n245391 , n245392 , n245393 , n245394 , n245395 , 
     n245396 , n245397 , n245398 , n245399 , n245400 , n245401 , n245402 , n245403 , n245404 , n245405 , 
     n245406 , n245407 , n245408 , n245409 , n245410 , n245411 , n245412 , n245413 , n245414 , n245415 , 
     n245416 , n245417 , n245418 , n245419 , n245420 , n245421 , n245422 , n245423 , n245424 , n245425 , 
     n245426 , n245427 , n245428 , n245429 , n245430 , n245431 , n245432 , n245433 , n245434 , n245435 , 
     n245436 , n245437 , n245438 , n245439 , n245440 , n245441 , n245442 , n245443 , n245444 , n245445 , 
     n245446 , n245447 , n245448 , n245449 , n245450 , n245451 , n245452 , n245453 , n245454 , n245455 , 
     n245456 , n245457 , n245458 , n245459 , n245460 , n245461 , n245462 , n245463 , n245464 , n245465 , 
     n245466 , n245467 , n245468 , n245469 , n245470 , n245471 , n245472 , n245473 , n245474 , n245475 , 
     n245476 , n245477 , n245478 , n245479 , n245480 , n245481 , n245482 , n245483 , n245484 , n245485 , 
     n245486 , n245487 , n245488 , n245489 , n245490 , n245491 , n245492 , n245493 , n245494 , n245495 , 
     n245496 , n245497 , n245498 , n245499 , n245500 , n245501 , n245502 , n245503 , n245504 , n245505 , 
     n245506 , n245507 , n245508 , n245509 , n245510 , n245511 , n245512 , n245513 , n245514 , n245515 , 
     n245516 , n245517 , n245518 , n245519 , n245520 , n245521 , n245522 , n245523 , n245524 , n245525 , 
     n245526 , n245527 , n245528 , n245529 , n245530 , n245531 , n245532 , n245533 , n245534 , n245535 , 
     n245536 , n245537 , n245538 , n245539 , n245540 , n245541 , n245542 , n245543 , n245544 , n245545 , 
     n245546 , n245547 , n245548 , n245549 , n245550 , n245551 , n245552 , n245553 , n245554 , n245555 , 
     n245556 , n245557 , n245558 , n245559 , n245560 , n245561 , n245562 , n245563 , n245564 , n245565 , 
     n245566 , n245567 , n245568 , n245569 , n245570 , n245571 , n245572 , n245573 , n245574 , n245575 , 
     n245576 , n245577 , n245578 , n245579 , n245580 , n245581 , n245582 , n245583 , n245584 , n245585 , 
     n245586 , n245587 , n245588 , n245589 , n245590 , n245591 , n245592 , n245593 , n245594 , n245595 , 
     n245596 , n245597 , n245598 , n245599 , n245600 , n245601 , n245602 , n245603 , n245604 , n245605 , 
     n245606 , n245607 , n245608 , n245609 , n245610 , n245611 , n245612 , n245613 , n245614 , n245615 , 
     n245616 , n245617 , n245618 , n245619 , n245620 , n245621 , n245622 , n245623 , n245624 , n245625 , 
     n245626 , n245627 , n245628 , n245629 , n245630 , n245631 , n245632 , n245633 , n245634 , n245635 , 
     n245636 , n245637 , n245638 , n245639 , n245640 , n245641 , n245642 , n245643 , n245644 , n245645 , 
     n245646 , n245647 , n245648 , n245649 , n245650 , n245651 , n245652 , n245653 , n245654 , n245655 , 
     n245656 , n245657 , n245658 , n245659 , n245660 , n245661 , n245662 , n245663 , n245664 , n245665 , 
     n245666 , n245667 , n245668 , n245669 , n245670 , n245671 , n245672 , n245673 , n245674 , n245675 , 
     n245676 , n245677 , n245678 , n245679 , n245680 , n245681 , n245682 , n245683 , n245684 , n245685 , 
     n245686 , n245687 , n245688 , n245689 , n245690 , n245691 , n245692 , n245693 , n245694 , n245695 , 
     n245696 , n245697 , n245698 , n245699 , n245700 , n245701 , n245702 , n245703 , n245704 , n245705 , 
     n245706 , n245707 , n245708 , n245709 , n245710 , n245711 , n245712 , n245713 , n245714 , n245715 , 
     n245716 , n245717 , n245718 , n245719 , n245720 , n245721 , n245722 , n245723 , n245724 , n245725 , 
     n245726 , n245727 , n245728 , n245729 , n245730 , n245731 , n245732 , n245733 , n245734 , n245735 , 
     n245736 , n245737 , n245738 , n245739 , n245740 , n245741 , n245742 , n245743 , n245744 , n245745 , 
     n245746 , n245747 , n245748 , n245749 , n245750 , n245751 , n245752 , n245753 , n245754 , n245755 , 
     n245756 , n245757 , n245758 , n245759 , n245760 , n245761 , n245762 , n245763 , n245764 , n245765 , 
     n245766 , n245767 , n245768 , n245769 , n245770 , n245771 , n245772 , n245773 , n245774 , n245775 , 
     n245776 , n245777 , n245778 , n245779 , n245780 , n245781 , n245782 , n245783 , n245784 , n245785 , 
     n245786 , n245787 , n245788 , n245789 , n245790 , n245791 , n245792 , n245793 , n245794 , n245795 , 
     n245796 , n245797 , n245798 , n245799 , n245800 , n245801 , n245802 , n245803 , n245804 , n245805 , 
     n245806 , n245807 , n245808 , n245809 , n245810 , n245811 , n245812 , n245813 , n245814 , n245815 , 
     n245816 , n245817 , n245818 , n245819 , n245820 , n245821 , n245822 , n245823 , n245824 , n245825 , 
     n245826 , n245827 , n245828 , n245829 , n245830 , n245831 , n245832 , n245833 , n245834 , n245835 , 
     n245836 , n245837 , n245838 , n245839 , n245840 , n245841 , n245842 , n245843 , n245844 , n245845 , 
     n245846 , n245847 , n245848 , n245849 , n245850 , n245851 , n245852 , n245853 , n245854 , n245855 , 
     n245856 , n245857 , n245858 , n245859 , n245860 , n245861 , n245862 , n245863 , n245864 , n245865 , 
     n245866 , n245867 , n245868 , n245869 , n245870 , n245871 , n245872 , n245873 , n245874 , n245875 , 
     n245876 , n245877 , n245878 , n245879 , n245880 , n245881 , n245882 , n245883 , n245884 , n245885 , 
     n245886 , n245887 , n245888 , n245889 , n245890 , n245891 , n245892 , n245893 , n245894 , n245895 , 
     n245896 , n245897 , n245898 , n245899 , n245900 , n245901 , n245902 , n245903 , n245904 , n245905 , 
     n245906 , n245907 , n245908 , n245909 , n245910 , n245911 , n245912 , n245913 , n245914 , n245915 , 
     n245916 , n245917 , n245918 , n245919 , n245920 , n245921 , n245922 , n245923 , n245924 , n245925 , 
     n245926 , n245927 , n245928 , n245929 , n245930 , n245931 , n245932 , n245933 , n245934 , n245935 , 
     n245936 , n245937 , n245938 , n245939 , n245940 , n245941 , n245942 , n245943 , n245944 , n245945 , 
     n245946 , n245947 , n245948 , n245949 , n245950 , n245951 , n245952 , n245953 , n245954 , n245955 , 
     n245956 , n245957 , n245958 , n245959 , n245960 , n245961 , n245962 , n245963 , n245964 , n245965 , 
     n245966 , n245967 , n245968 , n245969 , n245970 , n245971 , n245972 , n245973 , n245974 , n245975 , 
     n245976 , n245977 , n245978 , n245979 , n245980 , n245981 , n245982 , n245983 , n245984 , n245985 , 
     n245986 , n245987 , n245988 , n245989 , n245990 , n245991 , n245992 , n245993 , n245994 , n245995 , 
     n245996 , n245997 , n245998 , n245999 , n246000 , n246001 , n246002 , n246003 , n246004 , n246005 , 
     n246006 , n246007 , n246008 , n246009 , n246010 , n246011 , n246012 , n246013 , n246014 , n246015 , 
     n246016 , n246017 , n246018 , n246019 , n246020 , n246021 , n246022 , n246023 , n246024 , n246025 , 
     n246026 , n246027 , n246028 , n246029 , n246030 , n246031 , n246032 , n246033 , n246034 , n246035 , 
     n246036 , n246037 , n246038 , n246039 , n246040 , n246041 , n246042 , n246043 , n246044 , n246045 , 
     n246046 , n246047 , n246048 , n246049 , n246050 , n246051 , n246052 , n246053 , n246054 , n246055 , 
     n246056 , n246057 , n246058 , n246059 , n246060 , n246061 , n246062 , n246063 , n246064 , n246065 , 
     n246066 , n246067 , n246068 , n246069 , n246070 , n246071 , n246072 , n246073 , n246074 , n246075 , 
     n246076 , n246077 , n246078 , n246079 , n246080 , n246081 , n246082 , n246083 , n246084 , n246085 , 
     n246086 , n246087 , n246088 , n246089 , n246090 , n246091 , n246092 , n246093 , n246094 , n246095 , 
     n246096 , n246097 , n246098 , n246099 , n246100 , n246101 , n246102 , n246103 , n246104 , n246105 , 
     n246106 , n246107 , n246108 , n246109 , n246110 , n246111 , n246112 , n246113 , n246114 , n246115 , 
     n246116 , n246117 , n246118 , n246119 , n246120 , n246121 , n246122 , n246123 , n246124 , n246125 , 
     n246126 , n246127 , n246128 , n246129 , n246130 , n246131 , n246132 , n246133 , n246134 , n246135 , 
     n246136 , n246137 , n246138 , n246139 , n246140 , n246141 , n246142 , n246143 , n246144 , n246145 , 
     n246146 , n246147 , n246148 , n246149 , n246150 , n246151 , n246152 , n246153 , n246154 , n246155 , 
     n246156 , n246157 , n246158 , n246159 , n246160 , n246161 , n246162 , n246163 , n246164 , n246165 , 
     n246166 , n246167 , n246168 , n246169 , n246170 , n246171 , n246172 , n246173 , n246174 , n246175 , 
     n246176 , n246177 , n246178 , n246179 , n246180 , n246181 , n246182 , n246183 , n246184 , n246185 , 
     n246186 , n246187 , n246188 , n246189 , n246190 , n246191 , n246192 , n246193 , n246194 , n246195 , 
     n246196 , n246197 , n246198 , n246199 , n246200 , n246201 , n246202 , n246203 , n246204 , n246205 , 
     n246206 , n246207 , n246208 , n246209 , n246210 , n246211 , n246212 , n246213 , n246214 , n246215 , 
     n246216 , n246217 , n246218 , n246219 , n246220 , n246221 , n246222 , n246223 , n246224 , n246225 , 
     n246226 , n246227 , n246228 , n246229 , n246230 , n246231 , n246232 , n246233 , n246234 , n246235 , 
     n246236 , n246237 , n246238 , n246239 , n246240 , n246241 , n246242 , n246243 , n246244 , n246245 , 
     n246246 , n246247 , n246248 , n246249 , n246250 , n246251 , n246252 , n246253 , n246254 , n246255 , 
     n246256 , n246257 , n246258 , n246259 , n246260 , n246261 , n246262 , n246263 , n246264 , n246265 , 
     n246266 , n246267 , n246268 , n246269 , n246270 , n246271 , n246272 , n246273 , n246274 , n246275 , 
     n246276 , n246277 , n246278 , n246279 , n246280 , n246281 , n246282 , n246283 , n246284 , n246285 , 
     n246286 , n246287 , n246288 , n246289 , n246290 , n246291 , n246292 , n246293 , n246294 , n246295 , 
     n246296 , n246297 , n246298 , n246299 , n246300 , n246301 , n246302 , n246303 , n246304 , n246305 , 
     n246306 , n246307 , n246308 , n246309 , n246310 , n246311 , n246312 , n246313 , n246314 , n246315 , 
     n246316 , n246317 , n246318 , n246319 , n246320 , n246321 , n246322 , n246323 , n246324 , n246325 , 
     n246326 , n246327 , n246328 , n246329 , n246330 , n246331 , n246332 , n246333 , n246334 , n246335 , 
     n246336 , n246337 , n246338 , n246339 , n246340 , n246341 , n246342 , n246343 , n246344 , n246345 , 
     n246346 , n246347 , n246348 , n246349 , n246350 , n246351 , n246352 , n246353 , n246354 , n246355 , 
     n246356 , n246357 , n246358 , n246359 , n246360 , n246361 , n246362 , n246363 , n246364 , n246365 , 
     n246366 , n246367 , n246368 , n246369 , n246370 , n246371 , n246372 , n246373 , n246374 , n246375 , 
     n246376 , n246377 , n246378 , n246379 , n246380 , n246381 , n246382 , n246383 , n246384 , n246385 , 
     n246386 , n246387 , n246388 , n246389 , n246390 , n246391 , n246392 , n246393 , n246394 , n246395 , 
     n246396 , n246397 , n246398 , n246399 , n246400 , n246401 , n246402 , n246403 , n246404 , n246405 , 
     n246406 , n246407 , n246408 , n246409 , n246410 , n246411 , n246412 , n246413 , n246414 , n246415 , 
     n246416 , n246417 , n246418 , n246419 , n246420 , n246421 , n246422 , n246423 , n246424 , n246425 , 
     n246426 , n246427 , n246428 , n246429 , n246430 , n246431 , n246432 , n246433 , n246434 , n246435 , 
     n246436 , n246437 , n246438 , n246439 , n246440 , n246441 , n246442 , n246443 , n246444 , n246445 , 
     n246446 , n246447 , n246448 , n246449 , n246450 , n246451 , n246452 , n246453 , n246454 , n246455 , 
     n246456 , n246457 , n246458 , n246459 , n246460 , n246461 , n246462 , n246463 , n246464 , n246465 , 
     n246466 , n246467 , n246468 , n246469 , n246470 , n246471 , n246472 , n246473 , n246474 , n246475 , 
     n246476 , n246477 , n246478 , n246479 , n246480 , n246481 , n246482 , n246483 , n246484 , n246485 , 
     n246486 , n246487 , n246488 , n246489 , n246490 , n246491 , n246492 , n246493 , n246494 , n246495 , 
     n246496 , n246497 , n246498 , n246499 , n246500 , n246501 , n246502 , n246503 , n246504 , n246505 , 
     n246506 , n246507 , n246508 , n246509 , n246510 , n246511 , n246512 , n246513 , n246514 , n246515 , 
     n246516 , n246517 , n246518 , n246519 , n246520 , n246521 , n246522 , n246523 , n246524 , n246525 , 
     n246526 , n246527 , n246528 , n246529 , n246530 , n246531 , n246532 , n246533 , n246534 , n246535 , 
     n246536 , n246537 , n246538 , n246539 , n246540 , n246541 , n246542 , n246543 , n246544 , n246545 , 
     n246546 , n246547 , n246548 , n246549 , n246550 , n246551 , n246552 , n246553 , n246554 , n246555 , 
     n246556 , n246557 , n246558 , n246559 , n246560 , n246561 , n246562 , n246563 , n246564 , n246565 , 
     n246566 , n246567 , n246568 , n246569 , n246570 , n246571 , n246572 , n246573 , n246574 , n246575 , 
     n246576 , n246577 , n246578 , n246579 , n246580 , n246581 , n246582 , n246583 , n246584 , n246585 , 
     n246586 , n246587 , n246588 , n246589 , n246590 , n246591 , n246592 , n246593 , n246594 , n246595 , 
     n246596 , n246597 , n246598 , n246599 , n246600 , n246601 , n246602 , n246603 , n246604 , n246605 , 
     n246606 , n246607 , n246608 , n246609 , n246610 , n246611 , n246612 , n246613 , n246614 , n246615 , 
     n246616 , n246617 , n246618 , n246619 , n246620 , n246621 , n246622 , n246623 , n246624 , n246625 , 
     n246626 , n246627 , n246628 , n246629 , n246630 , n246631 , n246632 , n246633 , n246634 , n246635 , 
     n246636 , n246637 , n246638 , n246639 , n246640 , n246641 , n246642 , n246643 , n246644 , n246645 , 
     n246646 , n246647 , n246648 , n246649 , n246650 , n246651 , n246652 , n246653 , n246654 , n246655 , 
     n246656 , n246657 , n246658 , n246659 , n246660 , n246661 , n246662 , n246663 , n246664 , n246665 , 
     n246666 , n246667 , n246668 , n246669 , n246670 , n246671 , n246672 , n246673 , n246674 , n246675 , 
     n246676 , n246677 , n246678 , n246679 , n246680 , n246681 , n246682 , n246683 , n246684 , n246685 , 
     n246686 , n246687 , n246688 , n246689 , n246690 , n246691 , n246692 , n246693 , n246694 , n246695 , 
     n246696 , n246697 , n246698 , n246699 , n246700 , n246701 , n246702 , n246703 , n246704 , n246705 , 
     n246706 , n246707 , n246708 , n246709 , n246710 , n246711 , n246712 , n246713 , n246714 , n246715 , 
     n246716 , n246717 , n246718 , n246719 , n246720 , n246721 , n246722 , n246723 , n246724 , n246725 , 
     n246726 , n246727 , n246728 , n246729 , n246730 , n246731 , n246732 , n246733 , n246734 , n246735 , 
     n246736 , n246737 , n246738 , n246739 , n246740 , n246741 , n246742 , n246743 , n246744 , n246745 , 
     n246746 , n246747 , n246748 , n246749 , n246750 , n246751 , n246752 , n246753 , n246754 , n246755 , 
     n246756 , n246757 , n246758 , n246759 , n246760 , n246761 , n246762 , n246763 , n246764 , n246765 , 
     n246766 , n246767 , n246768 , n246769 , n246770 , n246771 , n246772 , n246773 , n246774 , n246775 , 
     n246776 , n246777 , n246778 , n246779 , n246780 , n246781 , n246782 , n246783 , n246784 , n246785 , 
     n246786 , n246787 , n246788 , n246789 , n246790 , n246791 , n246792 , n246793 , n246794 , n246795 , 
     n246796 , n246797 , n246798 , n246799 , n246800 , n246801 , n246802 , n246803 , n246804 , n246805 , 
     n246806 , n246807 , n246808 , n246809 , n246810 , n246811 , n246812 , n246813 , n246814 , n246815 , 
     n246816 , n246817 , n246818 , n246819 , n246820 , n246821 , n246822 , n246823 , n246824 , n246825 , 
     n246826 , n246827 , n246828 , n246829 , n246830 , n246831 , n246832 , n246833 , n246834 , n246835 , 
     n246836 , n246837 , n246838 , n246839 , n246840 , n246841 , n246842 , n246843 , n246844 , n246845 , 
     n246846 , n246847 , n246848 , n246849 , n246850 , n246851 , n246852 , n246853 , n246854 , n246855 , 
     n246856 , n246857 , n246858 , n246859 , n246860 , n246861 , n246862 , n246863 , n246864 , n246865 , 
     n246866 , n246867 , n246868 , n246869 , n246870 , n246871 , n246872 , n246873 , n246874 , n246875 , 
     n246876 , n246877 , n246878 , n246879 , n246880 , n246881 , n246882 , n246883 , n246884 , n246885 , 
     n246886 , n246887 , n246888 , n246889 , n246890 , n246891 , n246892 , n246893 , n246894 , n246895 , 
     n246896 , n246897 , n246898 , n246899 , n246900 , n246901 , n246902 , n246903 , n246904 , n246905 , 
     n246906 , n246907 , n246908 , n246909 , n246910 , n246911 , n246912 , n246913 , n246914 , n246915 , 
     n246916 , n246917 , n246918 , n246919 , n246920 , n246921 , n246922 , n246923 , n246924 , n246925 , 
     n246926 , n246927 , n246928 , n246929 , n246930 , n246931 , n246932 , n246933 , n246934 , n246935 , 
     n246936 , n246937 , n246938 , n246939 , n246940 , n246941 , n246942 , n246943 , n246944 , n246945 , 
     n246946 , n246947 , n246948 , n246949 , n246950 , n246951 , n246952 , n246953 , n246954 , n246955 , 
     n246956 , n246957 , n246958 , n246959 , n246960 , n246961 , n246962 , n246963 , n246964 , n246965 , 
     n246966 , n246967 , n246968 , n246969 , n246970 , n246971 , n246972 , n246973 , n246974 , n246975 , 
     n246976 , n246977 , n246978 , n246979 , n246980 , n246981 , n246982 , n246983 , n246984 , n246985 , 
     n246986 , n246987 , n246988 , n246989 , n246990 , n246991 , n246992 , n246993 , n246994 , n246995 , 
     n246996 , n246997 , n246998 , n246999 , n247000 , n247001 , n247002 , n247003 , n247004 , n247005 , 
     n247006 , n247007 , n247008 , n247009 , n247010 , n247011 , n247012 , n247013 , n247014 , n247015 , 
     n247016 , n247017 , n247018 , n247019 , n247020 , n247021 , n247022 , n247023 , n247024 , n247025 , 
     n247026 , n247027 , n247028 , n247029 , n247030 , n247031 , n247032 , n247033 , n247034 , n247035 , 
     n247036 , n247037 , n247038 , n247039 , n247040 , n247041 , n247042 , n247043 , n247044 , n247045 , 
     n247046 , n247047 , n247048 , n247049 , n247050 , n247051 , n247052 , n247053 , n247054 , n247055 , 
     n247056 , n247057 , n247058 , n247059 , n247060 , n247061 , n247062 , n247063 , n247064 , n247065 , 
     n247066 , n247067 , n247068 , n247069 , n247070 , n247071 , n247072 , n247073 , n247074 , n247075 , 
     n247076 , n247077 , n247078 , n247079 , n247080 , n247081 , n247082 , n247083 , n247084 , n247085 , 
     n247086 , n247087 , n247088 , n247089 , n247090 , n247091 , n247092 , n247093 , n247094 , n247095 , 
     n247096 , n247097 , n247098 , n247099 , n247100 , n247101 , n247102 , n247103 , n247104 , n247105 , 
     n247106 , n247107 , n247108 , n247109 , n247110 , n247111 , n247112 , n247113 , n247114 , n247115 , 
     n247116 , n247117 , n247118 , n247119 , n247120 , n247121 , n247122 , n247123 , n247124 , n247125 , 
     n247126 , n247127 , n247128 , n247129 , n247130 , n247131 , n247132 , n247133 , n247134 , n247135 , 
     n247136 , n247137 , n247138 , n247139 , n247140 , n247141 , n247142 , n247143 , n247144 , n247145 , 
     n247146 , n247147 , n247148 , n247149 , n247150 , n247151 , n247152 , n247153 , n247154 , n247155 , 
     n247156 , n247157 , n247158 , n247159 , n247160 , n247161 , n247162 , n247163 , n247164 , n247165 , 
     n247166 , n247167 , n247168 , n247169 , n247170 , n247171 , n247172 , n247173 , n247174 , n247175 , 
     n247176 , n247177 , n247178 , n247179 , n247180 , n247181 , n247182 , n247183 , n247184 , n247185 , 
     n247186 , n247187 , n247188 , n247189 , n247190 , n247191 , n247192 , n247193 , n247194 , n247195 , 
     n247196 , n247197 , n247198 , n247199 , n247200 , n247201 , n247202 , n247203 , n247204 , n247205 , 
     n247206 , n247207 , n247208 , n247209 , n247210 , n247211 , n247212 , n247213 , n247214 , n247215 , 
     n247216 , n247217 , n247218 , n247219 , n247220 , n247221 , n247222 , n247223 , n247224 , n247225 , 
     n247226 , n247227 , n247228 , n247229 , n247230 , n247231 , n247232 , n247233 , n247234 , n247235 , 
     n247236 , n247237 , n247238 , n247239 , n247240 , n247241 , n247242 , n247243 , n247244 , n247245 , 
     n247246 , n247247 , n247248 , n247249 , n247250 , n247251 , n247252 , n247253 , n247254 , n247255 , 
     n247256 , n247257 , n247258 , n247259 , n247260 , n247261 , n247262 , n247263 , n247264 , n247265 , 
     n247266 , n247267 , n247268 , n247269 , n247270 , n247271 , n247272 , n247273 , n247274 , n247275 , 
     n247276 , n247277 , n247278 , n247279 , n247280 , n247281 , n247282 , n247283 , n247284 , n247285 , 
     n247286 , n247287 , n247288 , n247289 , n247290 , n247291 , n247292 , n247293 , n247294 , n247295 , 
     n247296 , n247297 , n247298 , n247299 , n247300 , n247301 , n247302 , n247303 , n247304 , n247305 , 
     n247306 , n247307 , n247308 , n247309 , n247310 , n247311 , n247312 , n247313 , n247314 , n247315 , 
     n247316 , n247317 , n247318 , n247319 , n247320 , n247321 , n247322 , n247323 , n247324 , n247325 , 
     n247326 , n247327 , n247328 , n247329 , n247330 , n247331 , n247332 , n247333 , n247334 , n247335 , 
     n247336 , n247337 , n247338 , n247339 , n247340 , n247341 , n247342 , n247343 , n247344 , n247345 , 
     n247346 , n247347 , n247348 , n247349 , n247350 , n247351 , n247352 , n247353 , n247354 , n247355 , 
     n247356 , n247357 , n247358 , n247359 , n247360 , n247361 , n247362 , n247363 , n247364 , n247365 , 
     n247366 , n247367 , n247368 , n247369 , n247370 , n247371 , n247372 , n247373 , n247374 , n247375 , 
     n247376 , n247377 , n247378 , n247379 , n247380 , n247381 , n247382 , n247383 , n247384 , n247385 , 
     n247386 , n247387 , n247388 , n247389 , n247390 , n247391 , n247392 , n247393 , n247394 , n247395 , 
     n247396 , n247397 , n247398 , n247399 , n247400 , n247401 , n247402 , n247403 , n247404 , n247405 , 
     n247406 , n247407 , n247408 , n247409 , n247410 , n247411 , n247412 , n247413 , n247414 , n247415 , 
     n247416 , n247417 , n247418 , n247419 , n247420 , n247421 , n247422 , n247423 , n247424 , n247425 , 
     n247426 , n247427 , n247428 , n247429 , n247430 , n247431 , n247432 , n247433 , n247434 , n247435 , 
     n247436 , n247437 , n247438 , n247439 , n247440 , n247441 , n247442 , n247443 , n247444 , n247445 , 
     n247446 , n247447 , n247448 , n247449 , n247450 , n247451 , n247452 , n247453 , n247454 , n247455 , 
     n247456 , n247457 , n247458 , n247459 , n247460 , n247461 , n247462 , n247463 , n247464 , n247465 , 
     n247466 , n247467 , n247468 , n247469 , n247470 , n247471 , n247472 , n247473 , n247474 , n247475 , 
     n247476 , n247477 , n247478 , n247479 , n247480 , n247481 , n247482 , n247483 , n247484 , n247485 , 
     n247486 , n247487 , n247488 , n247489 , n247490 , n247491 , n247492 , n247493 , n247494 , n247495 , 
     n247496 , n247497 , n247498 , n247499 , n247500 , n247501 , n247502 , n247503 , n247504 , n247505 , 
     n247506 , n247507 , n247508 , n247509 , n247510 , n247511 , n247512 , n247513 , n247514 , n247515 , 
     n247516 , n247517 , n247518 , n247519 , n247520 , n247521 , n247522 , n247523 , n247524 , n247525 , 
     n247526 , n247527 , n247528 , n247529 , n247530 , n247531 , n247532 , n247533 , n247534 , n247535 , 
     n247536 , n247537 , n247538 , n247539 , n247540 , n247541 , n247542 , n247543 , n247544 , n247545 , 
     n247546 , n247547 , n247548 , n247549 , n247550 , n247551 , n247552 , n247553 , n247554 , n247555 , 
     n247556 , n247557 , n247558 , n247559 , n247560 , n247561 , n247562 , n247563 , n247564 , n247565 , 
     n247566 , n247567 , n247568 , n247569 , n247570 , n247571 , n247572 , n247573 , n247574 , n247575 , 
     n247576 , n247577 , n247578 , n247579 , n247580 , n247581 , n247582 , n247583 , n247584 , n247585 , 
     n247586 , n247587 , n247588 , n247589 , n247590 , n247591 , n247592 , n247593 , n247594 , n247595 , 
     n247596 , n247597 , n247598 , n247599 , n247600 , n247601 , n247602 , n247603 , n247604 , n247605 , 
     n247606 , n247607 , n247608 , n247609 , n247610 , n247611 , n247612 , n247613 , n247614 , n247615 , 
     n247616 , n247617 , n247618 , n247619 , n247620 , n247621 , n247622 , n247623 , n247624 , n247625 , 
     n247626 , n247627 , n247628 , n247629 , n247630 , n247631 , n247632 , n247633 , n247634 , n247635 , 
     n247636 , n247637 , n247638 , n247639 , n247640 , n247641 , n247642 , n247643 , n247644 , n247645 , 
     n247646 , n247647 , n247648 , n247649 , n247650 , n247651 , n247652 , n247653 , n247654 , n247655 , 
     n247656 , n247657 , n247658 , n247659 , n247660 , n247661 , n247662 , n247663 , n247664 , n247665 , 
     n247666 , n247667 , n247668 , n247669 , n247670 , n247671 , n247672 , n247673 , n247674 , n247675 , 
     n247676 , n247677 , n247678 , n247679 , n247680 , n247681 , n247682 , n247683 , n247684 , n247685 , 
     n247686 , n247687 , n247688 , n247689 , n247690 , n247691 , n247692 , n247693 , n247694 , n247695 , 
     n247696 , n247697 , n247698 , n247699 , n247700 , n247701 , n247702 , n247703 , n247704 , n247705 , 
     n247706 , n247707 , n247708 , n247709 , n247710 , n247711 , n247712 , n247713 , n247714 , n247715 , 
     n247716 , n247717 , n247718 , n247719 , n247720 , n247721 , n247722 , n247723 , n247724 , n247725 , 
     n247726 , n247727 , n247728 , n247729 , n247730 , n247731 , n247732 , n247733 , n247734 , n247735 , 
     n247736 , n247737 , n247738 , n247739 , n247740 , n247741 , n247742 , n247743 , n247744 , n247745 , 
     n247746 , n247747 , n247748 , n247749 , n247750 , n247751 , n247752 , n247753 , n247754 , n247755 , 
     n247756 , n247757 , n247758 , n247759 , n247760 , n247761 , n247762 , n247763 , n247764 , n247765 , 
     n247766 , n247767 , n247768 , n247769 , n247770 , n247771 , n247772 , n247773 , n247774 , n247775 , 
     n247776 , n247777 , n247778 , n247779 , n247780 , n247781 , n247782 , n247783 , n247784 , n247785 , 
     n247786 , n247787 , n247788 , n247789 , n247790 , n247791 , n247792 , n247793 , n247794 , n247795 , 
     n247796 , n247797 , n247798 , n247799 , n247800 , n247801 , n247802 , n247803 , n247804 , n247805 , 
     n247806 , n247807 , n247808 , n247809 , n247810 , n247811 , n247812 , n247813 , n247814 , n247815 , 
     n247816 , n247817 , n247818 , n247819 , n247820 , n247821 , n247822 , n247823 , n247824 , n247825 , 
     n247826 , n247827 , n247828 , n247829 , n247830 , n247831 , n247832 , n247833 , n247834 , n247835 , 
     n247836 , n247837 , n247838 , n247839 , n247840 , n247841 , n247842 , n247843 , n247844 , n247845 , 
     n247846 , n247847 , n247848 , n247849 , n247850 , n247851 , n247852 , n247853 , n247854 , n247855 , 
     n247856 , n247857 , n247858 , n247859 , n247860 , n247861 , n247862 , n247863 , n247864 , n247865 , 
     n247866 , n247867 , n247868 , n247869 , n247870 , n247871 , n247872 , n247873 , n247874 , n247875 , 
     n247876 , n247877 , n247878 , n247879 , n247880 , n247881 , n247882 , n247883 , n247884 , n247885 , 
     n247886 , n247887 , n247888 , n247889 , n247890 , n247891 , n247892 , n247893 , n247894 , n247895 , 
     n247896 , n247897 , n247898 , n247899 , n247900 , n247901 , n247902 , n247903 , n247904 , n247905 , 
     n247906 , n247907 , n247908 , n247909 , n247910 , n247911 , n247912 , n247913 , n247914 , n247915 , 
     n247916 , n247917 , n247918 , n247919 , n247920 , n247921 , n247922 , n247923 , n247924 , n247925 , 
     n247926 , n247927 , n247928 , n247929 , n247930 , n247931 , n247932 , n247933 , n247934 , n247935 , 
     n247936 , n247937 , n247938 , n247939 , n247940 , n247941 , n247942 , n247943 , n247944 , n247945 , 
     n247946 , n247947 , n247948 , n247949 , n247950 , n247951 , n247952 , n247953 , n247954 , n247955 , 
     n247956 , n247957 , n247958 , n247959 , n247960 , n247961 , n247962 , n247963 , n247964 , n247965 , 
     n247966 , n247967 , n247968 , n247969 , n247970 , n247971 , n247972 , n247973 , n247974 , n247975 , 
     n247976 , n247977 , n247978 , n247979 , n247980 , n247981 , n247982 , n247983 , n247984 , n247985 , 
     n247986 , n247987 , n247988 , n247989 , n247990 , n247991 , n247992 , n247993 , n247994 , n247995 , 
     n247996 , n247997 , n247998 , n247999 , n248000 , n248001 , n248002 , n248003 , n248004 , n248005 , 
     n248006 , n248007 , n248008 , n248009 , n248010 , n248011 , n248012 , n248013 , n248014 , n248015 , 
     n248016 , n248017 , n248018 , n248019 , n248020 , n248021 , n248022 , n248023 , n248024 , n248025 , 
     n248026 , n248027 , n248028 , n248029 , n248030 , n248031 , n248032 , n248033 , n248034 , n248035 , 
     n248036 , n248037 , n248038 , n248039 , n248040 , n248041 , n248042 , n248043 , n248044 , n248045 , 
     n248046 , n248047 , n248048 , n248049 , n248050 , n248051 , n248052 , n248053 , n248054 , n248055 , 
     n248056 , n248057 , n248058 , n248059 , n248060 , n248061 , n248062 , n248063 , n248064 , n248065 , 
     n248066 , n248067 , n248068 , n248069 , n248070 , n248071 , n248072 , n248073 , n248074 , n248075 , 
     n248076 , n248077 , n248078 , n248079 , n248080 , n248081 , n248082 , n248083 , n248084 , n248085 , 
     n248086 , n248087 , n248088 , n248089 , n248090 , n248091 , n248092 , n248093 , n248094 , n248095 , 
     n248096 , n248097 , n248098 , n248099 , n248100 , n248101 , n248102 , n248103 , n248104 , n248105 , 
     n248106 , n248107 , n248108 , n248109 , n248110 , n248111 , n248112 , n248113 , n248114 , n248115 , 
     n248116 , n248117 , n248118 , n248119 , n248120 , n248121 , n248122 , n248123 , n248124 , n248125 , 
     n248126 , n248127 , n248128 , n248129 , n248130 , n248131 , n248132 , n248133 , n248134 , n248135 , 
     n248136 , n248137 , n248138 , n248139 , n248140 , n248141 , n248142 , n248143 , n248144 , n248145 , 
     n248146 , n248147 , n248148 , n248149 , n248150 , n248151 , n248152 , n248153 , n248154 , n248155 , 
     n248156 , n248157 , n248158 , n248159 , n248160 , n248161 , n248162 , n248163 , n248164 , n248165 , 
     n248166 , n248167 , n248168 , n248169 , n248170 , n248171 , n248172 , n248173 , n248174 , n248175 , 
     n248176 , n248177 , n248178 , n248179 , n248180 , n248181 , n248182 , n248183 , n248184 , n248185 , 
     n248186 , n248187 , n248188 , n248189 , n248190 , n248191 , n248192 , n248193 , n248194 , n248195 , 
     n248196 , n248197 , n248198 , n248199 , n248200 , n248201 , n248202 , n248203 , n248204 , n248205 , 
     n248206 , n248207 , n248208 , n248209 , n248210 , n248211 , n248212 , n248213 , n248214 , n248215 , 
     n248216 , n248217 , n248218 , n248219 , n248220 , n248221 , n248222 , n248223 , n248224 , n248225 , 
     n248226 , n248227 , n248228 , n248229 , n248230 , n248231 , n248232 , n248233 , n248234 , n248235 , 
     n248236 , n248237 , n248238 , n248239 , n248240 , n248241 , n248242 , n248243 , n248244 , n248245 , 
     n248246 , n248247 , n248248 , n248249 , n248250 , n248251 , n248252 , n248253 , n248254 , n248255 , 
     n248256 , n248257 , n248258 , n248259 , n248260 , n248261 , n248262 , n248263 , n248264 , n248265 , 
     n248266 , n248267 , n248268 , n248269 , n248270 , n248271 , n248272 , n248273 , n248274 , n248275 , 
     n248276 , n248277 , n248278 , n248279 , n248280 , n248281 , n248282 , n248283 , n248284 , n248285 , 
     n248286 , n248287 , n248288 , n248289 , n248290 , n248291 , n248292 , n248293 , n248294 , n248295 , 
     n248296 , n248297 , n248298 , n248299 , n248300 , n248301 , n248302 , n248303 , n248304 , n248305 , 
     n248306 , n248307 , n248308 , n248309 , n248310 , n248311 , n248312 , n248313 , n248314 , n248315 , 
     n248316 , n248317 , n248318 , n248319 , n248320 , n248321 , n248322 , n248323 , n248324 , n248325 , 
     n248326 , n248327 , n248328 , n248329 , n248330 , n248331 , n248332 , n248333 , n248334 , n248335 , 
     n248336 , n248337 , n248338 , n248339 , n248340 , n248341 , n248342 , n248343 , n248344 , n248345 , 
     n248346 , n248347 , n248348 , n248349 , n248350 , n248351 , n248352 , n248353 , n248354 , n248355 , 
     n248356 , n248357 , n248358 , n248359 , n248360 , n248361 , n248362 , n248363 , n248364 , n248365 , 
     n248366 , n248367 , n248368 , n248369 , n248370 , n248371 , n248372 , n248373 , n248374 , n248375 , 
     n248376 , n248377 , n248378 , n248379 , n248380 , n248381 , n248382 , n248383 , n248384 , n248385 , 
     n248386 , n248387 , n248388 , n248389 , n248390 , n248391 , n248392 , n248393 , n248394 , n248395 , 
     n248396 , n248397 , n248398 , n248399 , n248400 , n248401 , n248402 , n248403 , n248404 , n248405 , 
     n248406 , n248407 , n248408 , n248409 , n248410 , n248411 , n248412 , n248413 , n248414 , n248415 , 
     n248416 , n248417 , n248418 , n248419 , n248420 , n248421 , n248422 , n248423 , n248424 , n248425 , 
     n248426 , n248427 , n248428 , n248429 , n248430 , n248431 , n248432 , n248433 , n248434 , n248435 , 
     n248436 , n248437 , n248438 , n248439 , n248440 , n248441 , n248442 , n248443 , n248444 , n248445 , 
     n248446 , n248447 , n248448 , n248449 , n248450 , n248451 , n248452 , n248453 , n248454 , n248455 , 
     n248456 , n248457 , n248458 , n248459 , n248460 , n248461 , n248462 , n248463 , n248464 , n248465 , 
     n248466 , n248467 , n248468 , n248469 , n248470 , n248471 , n248472 , n248473 , n248474 , n248475 , 
     n248476 , n248477 , n248478 , n248479 , n248480 , n248481 , n248482 , n248483 , n248484 , n248485 , 
     n248486 , n248487 , n248488 , n248489 , n248490 , n248491 , n248492 , n248493 , n248494 , n248495 , 
     n248496 , n248497 , n248498 , n248499 , n248500 , n248501 , n248502 , n248503 , n248504 , n248505 , 
     n248506 , n248507 , n248508 , n248509 , n248510 , n248511 , n248512 , n248513 , n248514 , n248515 , 
     n248516 , n248517 , n248518 , n248519 , n248520 , n248521 , n248522 , n248523 , n248524 , n248525 , 
     n248526 , n248527 , n248528 , n248529 , n248530 , n248531 , n248532 , n248533 , n248534 , n248535 , 
     n248536 , n248537 , n248538 , n248539 , n248540 , n248541 , n248542 , n248543 , n248544 , n248545 , 
     n248546 , n248547 , n248548 , n248549 , n248550 , n248551 , n248552 , n248553 , n248554 , n248555 , 
     n248556 , n248557 , n248558 , n248559 , n248560 , n248561 , n248562 , n248563 , n248564 , n248565 , 
     n248566 , n248567 , n248568 , n248569 , n248570 , n248571 , n248572 , n248573 , n248574 , n248575 , 
     n248576 , n248577 , n248578 , n248579 , n248580 , n248581 , n248582 , n248583 , n248584 , n248585 , 
     n248586 , n248587 , n248588 , n248589 , n248590 , n248591 , n248592 , n248593 , n248594 , n248595 , 
     n248596 , n248597 , n248598 , n248599 , n248600 , n248601 , n248602 , n248603 , n248604 , n248605 , 
     n248606 , n248607 , n248608 , n248609 , n248610 , n248611 , n248612 , n248613 , n248614 , n248615 , 
     n248616 , n248617 , n248618 , n248619 , n248620 , n248621 , n248622 , n248623 , n248624 , n248625 , 
     n248626 , n248627 , n248628 , n248629 , n248630 , n248631 , n248632 , n248633 , n248634 , n248635 , 
     n248636 , n248637 , n248638 , n248639 , n248640 , n248641 , n248642 , n248643 , n248644 , n248645 , 
     n248646 , n248647 , n248648 , n248649 , n248650 , n248651 , n248652 , n248653 , n248654 , n248655 , 
     n248656 , n248657 , n248658 , n248659 , n248660 , n248661 , n248662 , n248663 , n248664 , n248665 , 
     n248666 , n248667 , n248668 , n248669 , n248670 , n248671 , n248672 , n248673 , n248674 , n248675 , 
     n248676 , n248677 , n248678 , n248679 , n248680 , n248681 , n248682 , n248683 , n248684 , n248685 , 
     n248686 , n248687 , n248688 , n248689 , n248690 , n248691 , n248692 , n248693 , n248694 , n248695 , 
     n248696 , n248697 , n248698 , n248699 , n248700 , n248701 , n248702 , n248703 , n248704 , n248705 , 
     n248706 , n248707 , n248708 , n248709 , n248710 , n248711 , n248712 , n248713 , n248714 , n248715 , 
     n248716 , n248717 , n248718 , n248719 , n248720 , n248721 , n248722 , n248723 , n248724 , n248725 , 
     n248726 , n248727 , n248728 , n248729 , n248730 , n248731 , n248732 , n248733 , n248734 , n248735 , 
     n248736 , n248737 , n248738 , n248739 , n248740 , n248741 , n248742 , n248743 , n248744 , n248745 , 
     n248746 , n248747 , n248748 , n248749 , n248750 , n248751 , n248752 , n248753 , n248754 , n248755 , 
     n248756 , n248757 , n248758 , n248759 , n248760 , n248761 , n248762 , n248763 , n248764 , n248765 , 
     n248766 , n248767 , n248768 , n248769 , n248770 , n248771 , n248772 , n248773 , n248774 , n248775 , 
     n248776 , n248777 , n248778 , n248779 , n248780 , n248781 , n248782 , n248783 , n248784 , n248785 , 
     n248786 , n248787 , n248788 , n248789 , n248790 , n248791 , n248792 , n248793 , n248794 , n248795 , 
     n248796 , n248797 , n248798 , n248799 , n248800 , n248801 , n248802 , n248803 , n248804 , n248805 , 
     n248806 , n248807 , n248808 , n248809 , n248810 , n248811 , n248812 , n248813 , n248814 , n248815 , 
     n248816 , n248817 , n248818 , n248819 , n248820 , n248821 , n248822 , n248823 , n248824 , n248825 , 
     n248826 , n248827 , n248828 , n248829 , n248830 , n248831 , n248832 , n248833 , n248834 , n248835 , 
     n248836 , n248837 , n248838 , n248839 , n248840 , n248841 , n248842 , n248843 , n248844 , n248845 , 
     n248846 , n248847 , n248848 , n248849 , n248850 , n248851 , n248852 , n248853 , n248854 , n248855 , 
     n248856 , n248857 , n248858 , n248859 , n248860 , n248861 , n248862 , n248863 , n248864 , n248865 , 
     n248866 , n248867 , n248868 , n248869 , n248870 , n248871 , n248872 , n248873 , n248874 , n248875 , 
     n248876 , n248877 , n248878 , n248879 , n248880 , n248881 , n248882 , n248883 , n248884 , n248885 , 
     n248886 , n248887 , n248888 , n248889 , n248890 , n248891 , n248892 , n248893 , n248894 , n248895 , 
     n248896 , n248897 , n248898 , n248899 , n248900 , n248901 , n248902 , n248903 , n248904 , n248905 , 
     n248906 , n248907 , n248908 , n248909 , n248910 , n248911 , n248912 , n248913 , n248914 , n248915 , 
     n248916 , n248917 , n248918 , n248919 , n248920 , n248921 , n248922 , n248923 , n248924 , n248925 , 
     n248926 , n248927 , n248928 , n248929 , n248930 , n248931 , n248932 , n248933 , n248934 , n248935 , 
     n248936 , n248937 , n248938 , n248939 , n248940 , n248941 , n248942 , n248943 , n248944 , n248945 , 
     n248946 , n248947 , n248948 , n248949 , n248950 , n248951 , n248952 , n248953 , n248954 , n248955 , 
     n248956 , n248957 , n248958 , n248959 , n248960 , n248961 , n248962 , n248963 , n248964 , n248965 , 
     n248966 , n248967 , n248968 , n248969 , n248970 , n248971 , n248972 , n248973 , n248974 , n248975 , 
     n248976 , n248977 , n248978 , n248979 , n248980 , n248981 , n248982 , n248983 , n248984 , n248985 , 
     n248986 , n248987 , n248988 , n248989 , n248990 , n248991 , n248992 , n248993 , n248994 , n248995 , 
     n248996 , n248997 , n248998 , n248999 , n249000 , n249001 , n249002 , n249003 , n249004 , n249005 , 
     n249006 , n249007 , n249008 , n249009 , n249010 , n249011 , n249012 , n249013 , n249014 , n249015 , 
     n249016 , n249017 , n249018 , n249019 , n249020 , n249021 , n249022 , n249023 , n249024 , n249025 , 
     n249026 , n249027 , n249028 , n249029 , n249030 , n249031 , n249032 , n249033 , n249034 , n249035 , 
     n249036 , n249037 , n249038 , n249039 , n249040 , n249041 , n249042 , n249043 , n249044 , n249045 , 
     n249046 , n249047 , n249048 , n249049 , n249050 , n249051 , n249052 , n249053 , n249054 , n249055 , 
     n249056 , n249057 , n249058 , n249059 , n249060 , n249061 , n249062 , n249063 , n249064 , n249065 , 
     n249066 , n249067 , n249068 , n249069 , n249070 , n249071 , n249072 , n249073 , n249074 , n249075 , 
     n249076 , n249077 , n249078 , n249079 , n249080 , n249081 , n249082 , n249083 , n249084 , n249085 , 
     n249086 , n249087 , n249088 , n249089 , n249090 , n249091 , n249092 , n249093 , n249094 , n249095 , 
     n249096 , n249097 , n249098 , n249099 , n249100 , n249101 , n249102 , n249103 , n249104 , n249105 , 
     n249106 , n249107 , n249108 , n249109 , n249110 , n249111 , n249112 , n249113 , n249114 , n249115 , 
     n249116 , n249117 , n249118 , n249119 , n249120 , n249121 , n249122 , n249123 , n249124 , n249125 , 
     n249126 , n249127 , n249128 , n249129 , n249130 , n249131 , n249132 , n249133 , n249134 , n249135 , 
     n249136 , n249137 , n249138 , n249139 , n249140 , n249141 , n249142 , n249143 , n249144 , n249145 , 
     n249146 , n249147 , n249148 , n249149 , n249150 , n249151 , n249152 , n249153 , n249154 , n249155 , 
     n249156 , n249157 , n249158 , n249159 , n249160 , n249161 , n249162 , n249163 , n249164 , n249165 , 
     n249166 , n249167 , n249168 , n249169 , n249170 , n249171 , n249172 , n249173 , n249174 , n249175 , 
     n249176 , n249177 , n249178 , n249179 , n249180 , n249181 , n249182 , n249183 , n249184 , n249185 , 
     n249186 , n249187 , n249188 , n249189 , n249190 , n249191 , n249192 , n249193 , n249194 , n249195 , 
     n249196 , n249197 , n249198 , n249199 , n249200 , n249201 , n249202 , n249203 , n249204 , n249205 , 
     n249206 , n249207 , n249208 , n249209 , n249210 , n249211 , n249212 , n249213 , n249214 , n249215 , 
     n249216 , n249217 , n249218 , n249219 , n249220 , n249221 , n249222 , n249223 , n249224 , n249225 , 
     n249226 , n249227 , n249228 , n249229 , n249230 , n249231 , n249232 , n249233 , n249234 , n249235 , 
     n249236 , n249237 , n249238 , n249239 , n249240 , n249241 , n249242 , n249243 , n249244 , n249245 , 
     n249246 , n249247 , n249248 , n249249 , n249250 , n249251 , n249252 , n249253 , n249254 , n249255 , 
     n249256 , n249257 , n249258 , n249259 , n249260 , n249261 , n249262 , n249263 , n249264 , n249265 , 
     n249266 , n249267 , n249268 , n249269 , n249270 , n249271 , n249272 , n249273 , n249274 , n249275 , 
     n249276 , n249277 , n249278 , n249279 , n249280 , n249281 , n249282 , n249283 , n249284 , n249285 , 
     n249286 , n249287 , n249288 , n249289 , n249290 , n249291 , n249292 , n249293 , n249294 , n249295 , 
     n249296 , n249297 , n249298 , n249299 , n249300 , n249301 , n249302 , n249303 , n249304 , n249305 , 
     n249306 , n249307 , n249308 , n249309 , n249310 , n249311 , n249312 , n249313 , n249314 , n249315 , 
     n249316 , n249317 , n249318 , n249319 , n249320 , n249321 , n249322 , n249323 , n249324 , n249325 , 
     n249326 , n249327 , n249328 , n249329 , n249330 , n249331 , n249332 , n249333 , n249334 , n249335 , 
     n249336 , n249337 , n249338 , n249339 , n249340 , n249341 , n249342 , n249343 , n249344 , n249345 , 
     n249346 , n249347 , n249348 , n249349 , n249350 , n249351 , n249352 , n249353 , n249354 , n249355 , 
     n249356 , n249357 , n249358 , n249359 , n249360 , n249361 , n249362 , n249363 , n249364 , n249365 , 
     n249366 , n249367 , n249368 , n249369 , n249370 , n249371 , n249372 , n249373 , n249374 , n249375 , 
     n249376 , n249377 , n249378 , n249379 , n249380 , n249381 , n249382 , n249383 , n249384 , n249385 , 
     n249386 , n249387 , n249388 , n249389 , n249390 , n249391 , n249392 , n249393 , n249394 , n249395 , 
     n249396 , n249397 , n249398 , n249399 , n249400 , n249401 , n249402 , n249403 , n249404 , n249405 , 
     n249406 , n249407 , n249408 , n249409 , n249410 , n249411 , n249412 , n249413 , n249414 , n249415 , 
     n249416 , n249417 , n249418 , n249419 , n249420 , n249421 , n249422 , n249423 , n249424 , n249425 , 
     n249426 , n249427 , n249428 , n249429 , n249430 , n249431 , n249432 , n249433 , n249434 , n249435 , 
     n249436 , n249437 , n249438 , n249439 , n249440 , n249441 , n249442 , n249443 , n249444 , n249445 , 
     n249446 , n249447 , n249448 , n249449 , n249450 , n249451 , n249452 , n249453 , n249454 , n249455 , 
     n249456 , n249457 , n249458 , n249459 , n249460 , n249461 , n249462 , n249463 , n249464 , n249465 , 
     n249466 , n249467 , n249468 , n249469 , n249470 , n249471 , n249472 , n249473 , n249474 , n249475 , 
     n249476 , n249477 , n249478 , n249479 , n249480 , n249481 , n249482 , n249483 , n249484 , n249485 , 
     n249486 , n249487 , n249488 , n249489 , n249490 , n249491 , n249492 , n249493 , n249494 , n249495 , 
     n249496 , n249497 , n249498 , n249499 , n249500 , n249501 , n249502 , n249503 , n249504 , n249505 , 
     n249506 , n249507 , n249508 , n249509 , n249510 , n249511 , n249512 , n249513 , n249514 , n249515 , 
     n249516 , n249517 , n249518 , n249519 , n249520 , n249521 , n249522 , n249523 , n249524 , n249525 , 
     n249526 , n249527 , n249528 , n249529 , n249530 , n249531 , n249532 , n249533 , n249534 , n249535 , 
     n249536 , n249537 , n249538 , n249539 , n249540 , n249541 , n249542 , n249543 , n249544 , n249545 , 
     n249546 , n249547 , n249548 , n249549 , n249550 , n249551 , n249552 , n249553 , n249554 , n249555 , 
     n249556 , n249557 , n249558 , n249559 , n249560 , n249561 , n249562 , n249563 , n249564 , n249565 , 
     n249566 , n249567 , n249568 , n249569 , n249570 , n249571 , n249572 , n249573 , n249574 , n249575 , 
     n249576 , n249577 , n249578 , n249579 , n249580 , n249581 , n249582 , n249583 , n249584 , n249585 , 
     n249586 , n249587 , n249588 , n249589 , n249590 , n249591 , n249592 , n249593 , n249594 , n249595 , 
     n249596 , n249597 , n249598 , n249599 , n249600 , n249601 , n249602 , n249603 , n249604 , n249605 , 
     n249606 , n249607 , n249608 , n249609 , n249610 , n249611 , n249612 , n249613 , n249614 , n249615 , 
     n249616 , n249617 , n249618 , n249619 , n249620 , n249621 , n249622 , n249623 , n249624 , n249625 , 
     n249626 , n249627 , n249628 , n249629 , n249630 , n249631 , n249632 , n249633 , n249634 , n249635 , 
     n249636 , n249637 , n249638 , n249639 , n249640 , n249641 , n249642 , n249643 , n249644 , n249645 , 
     n249646 , n249647 , n249648 , n249649 , n249650 , n249651 , n249652 , n249653 , n249654 , n249655 , 
     n249656 , n249657 , n249658 , n249659 , n249660 , n249661 , n249662 , n249663 , n249664 , n249665 , 
     n249666 , n249667 , n249668 , n249669 , n249670 , n249671 , n249672 , n249673 , n249674 , n249675 , 
     n249676 , n249677 , n249678 , n249679 , n249680 , n249681 , n249682 , n249683 , n249684 , n249685 , 
     n249686 , n249687 , n249688 , n249689 , n249690 , n249691 , n249692 , n249693 , n249694 , n249695 , 
     n249696 , n249697 , n249698 , n249699 , n249700 , n249701 , n249702 , n249703 , n249704 , n249705 , 
     n249706 , n249707 , n249708 , n249709 , n249710 , n249711 , n249712 , n249713 , n249714 , n249715 , 
     n249716 , n249717 , n249718 , n249719 , n249720 , n249721 , n249722 , n249723 , n249724 , n249725 , 
     n249726 , n249727 , n249728 , n249729 , n249730 , n249731 , n249732 , n249733 , n249734 , n249735 , 
     n249736 , n249737 , n249738 , n249739 , n249740 , n249741 , n249742 , n249743 , n249744 , n249745 , 
     n249746 , n249747 , n249748 , n249749 , n249750 , n249751 , n249752 , n249753 , n249754 , n249755 , 
     n249756 , n249757 , n249758 , n249759 , n249760 , n249761 , n249762 , n249763 , n249764 , n249765 , 
     n249766 , n249767 , n249768 , n249769 , n249770 , n249771 , n249772 , n249773 , n249774 , n249775 , 
     n249776 , n249777 , n249778 , n249779 , n249780 , n249781 , n249782 , n249783 , n249784 , n249785 , 
     n249786 , n249787 , n249788 , n249789 , n249790 , n249791 , n249792 , n249793 , n249794 , n249795 , 
     n249796 , n249797 , n249798 , n249799 , n249800 , n249801 , n249802 , n249803 , n249804 , n249805 , 
     n249806 , n249807 , n249808 , n249809 , n249810 , n249811 , n249812 , n249813 , n249814 , n249815 , 
     n249816 , n249817 , n249818 , n249819 , n249820 , n249821 , n249822 , n249823 , n249824 , n249825 , 
     n249826 , n249827 , n249828 , n249829 , n249830 , n249831 , n249832 , n249833 , n249834 , n249835 , 
     n249836 , n249837 , n249838 , n249839 , n249840 , n249841 , n249842 , n249843 , n249844 , n249845 , 
     n249846 , n249847 , n249848 , n249849 , n249850 , n249851 , n249852 , n249853 , n249854 , n249855 , 
     n249856 , n249857 , n249858 , n249859 , n249860 , n249861 , n249862 , n249863 , n249864 , n249865 , 
     n249866 , n249867 , n249868 , n249869 , n249870 , n249871 , n249872 , n249873 , n249874 , n249875 , 
     n249876 , n249877 , n249878 , n249879 , n249880 , n249881 , n249882 , n249883 , n249884 , n249885 , 
     n249886 , n249887 , n249888 , n249889 , n249890 , n249891 , n249892 , n249893 , n249894 , n249895 , 
     n249896 , n249897 , n249898 , n249899 , n249900 , n249901 , n249902 , n249903 , n249904 , n249905 , 
     n249906 , n249907 , n249908 , n249909 , n249910 , n249911 , n249912 , n249913 , n249914 , n249915 , 
     n249916 , n249917 , n249918 , n249919 , n249920 , n249921 , n249922 , n249923 , n249924 , n249925 , 
     n249926 , n249927 , n249928 , n249929 , n249930 , n249931 , n249932 , n249933 , n249934 , n249935 , 
     n249936 , n249937 , n249938 , n249939 , n249940 , n249941 , n249942 , n249943 , n249944 , n249945 , 
     n249946 , n249947 , n249948 , n249949 , n249950 , n249951 , n249952 , n249953 , n249954 , n249955 , 
     n249956 , n249957 , n249958 , n249959 , n249960 , n249961 , n249962 , n249963 , n249964 , n249965 , 
     n249966 , n249967 , n249968 , n249969 , n249970 , n249971 , n249972 , n249973 , n249974 , n249975 , 
     n249976 , n249977 , n249978 , n249979 , n249980 , n249981 , n249982 , n249983 , n249984 , n249985 , 
     n249986 , n249987 , n249988 , n249989 , n249990 , n249991 , n249992 , n249993 , n249994 , n249995 , 
     n249996 , n249997 , n249998 , n249999 , n250000 , n250001 , n250002 , n250003 , n250004 , n250005 , 
     n250006 , n250007 , n250008 , n250009 , n250010 , n250011 , n250012 , n250013 , n250014 , n250015 , 
     n250016 , n250017 , n250018 , n250019 , n250020 , n250021 , n250022 , n250023 , n250024 , n250025 , 
     n250026 , n250027 , n250028 , n250029 , n250030 , n250031 , n250032 , n250033 , n250034 , n250035 , 
     n250036 , n250037 , n250038 , n250039 , n250040 , n250041 , n250042 , n250043 , n250044 , n250045 , 
     n250046 , n250047 , n250048 , n250049 , n250050 , n250051 , n250052 , n250053 , n250054 , n250055 , 
     n250056 , n250057 , n250058 , n250059 , n250060 , n250061 , n250062 , n250063 , n250064 , n250065 , 
     n250066 , n250067 , n250068 , n250069 , n250070 , n250071 , n250072 , n250073 , n250074 , n250075 , 
     n250076 , n250077 , n250078 , n250079 , n250080 , n250081 , n250082 , n250083 , n250084 , n250085 , 
     n250086 , n250087 , n250088 , n250089 , n250090 , n250091 , n250092 , n250093 , n250094 , n250095 , 
     n250096 , n250097 , n250098 , n250099 , n250100 , n250101 , n250102 , n250103 , n250104 , n250105 , 
     n250106 , n250107 , n250108 , n250109 , n250110 , n250111 , n250112 , n250113 , n250114 , n250115 , 
     n250116 , n250117 , n250118 , n250119 , n250120 , n250121 , n250122 , n250123 , n250124 , n250125 , 
     n250126 , n250127 , n250128 , n250129 , n250130 , n250131 , n250132 , n250133 , n250134 , n250135 , 
     n250136 , n250137 , n250138 , n250139 , n250140 , n250141 , n250142 , n250143 , n250144 , n250145 , 
     n250146 , n250147 , n250148 , n250149 , n250150 , n250151 , n250152 , n250153 , n250154 , n250155 , 
     n250156 , n250157 , n250158 , n250159 , n250160 , n250161 , n250162 , n250163 , n250164 , n250165 , 
     n250166 , n250167 , n250168 , n250169 , n250170 , n250171 , n250172 , n250173 , n250174 , n250175 , 
     n250176 , n250177 , n250178 , n250179 , n250180 , n250181 , n250182 , n250183 , n250184 , n250185 , 
     n250186 , n250187 , n250188 , n250189 , n250190 , n250191 , n250192 , n250193 , n250194 , n250195 , 
     n250196 , n250197 , n250198 , n250199 , n250200 , n250201 , n250202 , n250203 , n250204 , n250205 , 
     n250206 , n250207 , n250208 , n250209 , n250210 , n250211 , n250212 , n250213 , n250214 , n250215 , 
     n250216 , n250217 , n250218 , n250219 , n250220 , n250221 , n250222 , n250223 , n250224 , n250225 , 
     n250226 , n250227 , n250228 , n250229 , n250230 , n250231 , n250232 , n250233 , n250234 , n250235 , 
     n250236 , n250237 , n250238 , n250239 , n250240 , n250241 , n250242 , n250243 , n250244 , n250245 , 
     n250246 , n250247 , n250248 , n250249 , n250250 , n250251 , n250252 , n250253 , n250254 , n250255 , 
     n250256 , n250257 , n250258 , n250259 , n250260 , n250261 , n250262 , n250263 , n250264 , n250265 , 
     n250266 , n250267 , n250268 , n250269 , n250270 , n250271 , n250272 , n250273 , n250274 , n250275 , 
     n250276 , n250277 , n250278 , n250279 , n250280 , n250281 , n250282 , n250283 , n250284 , n250285 , 
     n250286 , n250287 , n250288 , n250289 , n250290 , n250291 , n250292 , n250293 , n250294 , n250295 , 
     n250296 , n250297 , n250298 , n250299 , n250300 , n250301 , n250302 , n250303 , n250304 , n250305 , 
     n250306 , n250307 , n250308 , n250309 , n250310 , n250311 , n250312 , n250313 , n250314 , n250315 , 
     n250316 , n250317 , n250318 , n250319 , n250320 , n250321 , n250322 , n250323 , n250324 , n250325 , 
     n250326 , n250327 , n250328 , n250329 , n250330 , n250331 , n250332 , n250333 , n250334 , n250335 , 
     n250336 , n250337 , n250338 , n250339 , n250340 , n250341 , n250342 , n250343 , n250344 , n250345 , 
     n250346 , n250347 , n250348 , n250349 , n250350 , n250351 , n250352 , n250353 , n250354 , n250355 , 
     n250356 , n250357 , n250358 , n250359 , n250360 , n250361 , n250362 , n250363 , n250364 , n250365 , 
     n250366 , n250367 , n250368 , n250369 , n250370 , n250371 , n250372 , n250373 , n250374 , n250375 , 
     n250376 , n250377 , n250378 , n250379 , n250380 , n250381 , n250382 , n250383 , n250384 , n250385 , 
     n250386 , n250387 , n250388 , n250389 , n250390 , n250391 , n250392 , n250393 , n250394 , n250395 , 
     n250396 , n250397 , n250398 , n250399 , n250400 , n250401 , n250402 , n250403 , n250404 , n250405 , 
     n250406 , n250407 , n250408 , n250409 , n250410 , n250411 , n250412 , n250413 , n250414 , n250415 , 
     n250416 , n250417 , n250418 , n250419 , n250420 , n250421 , n250422 , n250423 , n250424 , n250425 , 
     n250426 , n250427 , n250428 , n250429 , n250430 , n250431 , n250432 , n250433 , n250434 , n250435 , 
     n250436 , n250437 , n250438 , n250439 , n250440 , n250441 , n250442 , n250443 , n250444 , n250445 , 
     n250446 , n250447 , n250448 , n250449 , n250450 , n250451 , n250452 , n250453 , n250454 , n250455 , 
     n250456 , n250457 , n250458 , n250459 , n250460 , n250461 , n250462 , n250463 , n250464 , n250465 , 
     n250466 , n250467 , n250468 , n250469 , n250470 , n250471 , n250472 , n250473 , n250474 , n250475 , 
     n250476 , n250477 , n250478 , n250479 , n250480 , n250481 , n250482 , n250483 , n250484 , n250485 , 
     n250486 , n250487 , n250488 , n250489 , n250490 , n250491 , n250492 , n250493 , n250494 , n250495 , 
     n250496 , n250497 , n250498 , n250499 , n250500 , n250501 , n250502 , n250503 , n250504 , n250505 , 
     n250506 , n250507 , n250508 , n250509 , n250510 , n250511 , n250512 , n250513 , n250514 , n250515 , 
     n250516 , n250517 , n250518 , n250519 , n250520 , n250521 , n250522 , n250523 , n250524 , n250525 , 
     n250526 , n250527 , n250528 , n250529 , n250530 , n250531 , n250532 , n250533 , n250534 , n250535 , 
     n250536 , n250537 , n250538 , n250539 , n250540 , n250541 , n250542 , n250543 , n250544 , n250545 , 
     n250546 , n250547 , n250548 , n250549 , n250550 , n250551 , n250552 , n250553 , n250554 , n250555 , 
     n250556 , n250557 , n250558 , n250559 , n250560 , n250561 , n250562 , n250563 , n250564 , n250565 , 
     n250566 , n250567 , n250568 , n250569 , n250570 , n250571 , n250572 , n250573 , n250574 , n250575 , 
     n250576 , n250577 , n250578 , n250579 , n250580 , n250581 , n250582 , n250583 , n250584 , n250585 , 
     n250586 , n250587 , n250588 , n250589 , n250590 , n250591 , n250592 , n250593 , n250594 , n250595 , 
     n250596 , n250597 , n250598 , n250599 , n250600 , n250601 , n250602 , n250603 , n250604 , n250605 , 
     n250606 , n250607 , n250608 , n250609 , n250610 , n250611 , n250612 , n250613 , n250614 , n250615 , 
     n250616 , n250617 , n250618 , n250619 , n250620 , n250621 , n250622 , n250623 , n250624 , n250625 , 
     n250626 , n250627 , n250628 , n250629 , n250630 , n250631 , n250632 , n250633 , n250634 , n250635 , 
     n250636 , n250637 , n250638 , n250639 , n250640 , n250641 , n250642 , n250643 , n250644 , n250645 , 
     n250646 , n250647 , n250648 , n250649 , n250650 , n250651 , n250652 , n250653 , n250654 , n250655 , 
     n250656 , n250657 , n250658 , n250659 , n250660 , n250661 , n250662 , n250663 , n250664 , n250665 , 
     n250666 , n250667 , n250668 , n250669 , n250670 , n250671 , n250672 , n250673 , n250674 , n250675 , 
     n250676 , n250677 , n250678 , n250679 , n250680 , n250681 , n250682 , n250683 , n250684 , n250685 , 
     n250686 , n250687 , n250688 , n250689 , n250690 , n250691 , n250692 , n250693 , n250694 , n250695 , 
     n250696 , n250697 , n250698 , n250699 , n250700 , n250701 , n250702 , n250703 , n250704 , n250705 , 
     n250706 , n250707 , n250708 , n250709 , n250710 , n250711 , n250712 , n250713 , n250714 , n250715 , 
     n250716 , n250717 , n250718 , n250719 , n250720 , n250721 , n250722 , n250723 , n250724 , n250725 , 
     n250726 , n250727 , n250728 , n250729 , n250730 , n250731 , n250732 , n250733 , n250734 , n250735 , 
     n250736 , n250737 , n250738 , n250739 , n250740 , n250741 , n250742 , n250743 , n250744 , n250745 , 
     n250746 , n250747 , n250748 , n250749 , n250750 , n250751 , n250752 , n250753 , n250754 , n250755 , 
     n250756 , n250757 , n250758 , n250759 , n250760 , n250761 , n250762 , n250763 , n250764 , n250765 , 
     n250766 , n250767 , n250768 , n250769 , n250770 , n250771 , n250772 , n250773 , n250774 , n250775 , 
     n250776 , n250777 , n250778 , n250779 , n250780 , n250781 , n250782 , n250783 , n250784 , n250785 , 
     n250786 , n250787 , n250788 , n250789 , n250790 , n250791 , n250792 , n250793 , n250794 , n250795 , 
     n250796 , n250797 , n250798 , n250799 , n250800 , n250801 , n250802 , n250803 , n250804 , n250805 , 
     n250806 , n250807 , n250808 , n250809 , n250810 , n250811 , n250812 , n250813 , n250814 , n250815 , 
     n250816 , n250817 , n250818 , n250819 , n250820 , n250821 , n250822 , n250823 , n250824 , n250825 , 
     n250826 , n250827 , n250828 , n250829 , n250830 , n250831 , n250832 , n250833 , n250834 , n250835 , 
     n250836 , n250837 , n250838 , n250839 , n250840 , n250841 , n250842 , n250843 , n250844 , n250845 , 
     n250846 , n250847 , n250848 , n250849 , n250850 , n250851 , n250852 , n250853 , n250854 , n250855 , 
     n250856 , n250857 , n250858 , n250859 , n250860 , n250861 , n250862 , n250863 , n250864 , n250865 , 
     n250866 , n250867 , n250868 , n250869 , n250870 , n250871 , n250872 , n250873 , n250874 , n250875 , 
     n250876 , n250877 , n250878 , n250879 , n250880 , n250881 , n250882 , n250883 , n250884 , n250885 , 
     n250886 , n250887 , n250888 , n250889 , n250890 , n250891 , n250892 , n250893 , n250894 , n250895 , 
     n250896 , n250897 , n250898 , n250899 , n250900 , n250901 , n250902 , n250903 , n250904 , n250905 , 
     n250906 , n250907 , n250908 , n250909 , n250910 , n250911 , n250912 , n250913 , n250914 , n250915 , 
     n250916 , n250917 , n250918 , n250919 , n250920 , n250921 , n250922 , n250923 , n250924 , n250925 , 
     n250926 , n250927 , n250928 , n250929 , n250930 , n250931 , n250932 , n250933 , n250934 , n250935 , 
     n250936 , n250937 , n250938 , n250939 , n250940 , n250941 , n250942 , n250943 , n250944 , n250945 , 
     n250946 , n250947 , n250948 , n250949 , n250950 , n250951 , n250952 , n250953 , n250954 , n250955 , 
     n250956 , n250957 , n250958 , n250959 , n250960 , n250961 , n250962 , n250963 , n250964 , n250965 , 
     n250966 , n250967 , n250968 , n250969 , n250970 , n250971 , n250972 , n250973 , n250974 , n250975 , 
     n250976 , n250977 , n250978 , n250979 , n250980 , n250981 , n250982 , n250983 , n250984 , n250985 , 
     n250986 , n250987 , n250988 , n250989 , n250990 , n250991 , n250992 , n250993 , n250994 , n250995 , 
     n250996 , n250997 , n250998 , n250999 , n251000 , n251001 , n251002 , n251003 , n251004 , n251005 , 
     n251006 , n251007 , n251008 , n251009 , n251010 , n251011 , n251012 , n251013 , n251014 , n251015 , 
     n251016 , n251017 , n251018 , n251019 , n251020 , n251021 , n251022 , n251023 , n251024 , n251025 , 
     n251026 , n251027 , n251028 , n251029 , n251030 , n251031 , n251032 , n251033 , n251034 , n251035 , 
     n251036 , n251037 , n251038 , n251039 , n251040 , n251041 , n251042 , n251043 , n251044 , n251045 , 
     n251046 , n251047 , n251048 , n251049 , n251050 , n251051 , n251052 , n251053 , n251054 , n251055 , 
     n251056 , n251057 , n251058 , n251059 , n251060 , n251061 , n251062 , n251063 , n251064 , n251065 , 
     n251066 , n251067 , n251068 , n251069 , n251070 , n251071 , n251072 , n251073 , n251074 , n251075 , 
     n251076 , n251077 , n251078 , n251079 , n251080 , n251081 , n251082 , n251083 , n251084 , n251085 , 
     n251086 , n251087 , n251088 , n251089 , n251090 , n251091 , n251092 , n251093 , n251094 , n251095 , 
     n251096 , n251097 , n251098 , n251099 , n251100 , n251101 , n251102 , n251103 , n251104 , n251105 , 
     n251106 , n251107 , n251108 , n251109 , n251110 , n251111 , n251112 , n251113 , n251114 , n251115 , 
     n251116 , n251117 , n251118 , n251119 , n251120 , n251121 , n251122 , n251123 , n251124 , n251125 , 
     n251126 , n251127 , n251128 , n251129 , n251130 , n251131 , n251132 , n251133 , n251134 , n251135 , 
     n251136 , n251137 , n251138 , n251139 , n251140 , n251141 , n251142 , n251143 , n251144 , n251145 , 
     n251146 , n251147 , n251148 , n251149 , n251150 , n251151 , n251152 , n251153 , n251154 , n251155 , 
     n251156 , n251157 , n251158 , n251159 , n251160 , n251161 , n251162 , n251163 , n251164 , n251165 , 
     n251166 , n251167 , n251168 , n251169 , n251170 , n251171 , n251172 , n251173 , n251174 , n251175 , 
     n251176 , n251177 , n251178 , n251179 , n251180 , n251181 , n251182 , n251183 , n251184 , n251185 , 
     n251186 , n251187 , n251188 , n251189 , n251190 , n251191 , n251192 , n251193 , n251194 , n251195 , 
     n251196 , n251197 , n251198 , n251199 , n251200 , n251201 , n251202 , n251203 , n251204 , n251205 , 
     n251206 , n251207 , n251208 , n251209 , n251210 , n251211 , n251212 , n251213 , n251214 , n251215 , 
     n251216 , n251217 , n251218 , n251219 , n251220 , n251221 , n251222 , n251223 , n251224 , n251225 , 
     n251226 , n251227 , n251228 , n251229 , n251230 , n251231 , n251232 , n251233 , n251234 , n251235 , 
     n251236 , n251237 , n251238 , n251239 , n251240 , n251241 , n251242 , n251243 , n251244 , n251245 , 
     n251246 , n251247 , n251248 , n251249 , n251250 , n251251 , n251252 , n251253 , n251254 , n251255 , 
     n251256 , n251257 , n251258 , n251259 , n251260 , n251261 , n251262 , n251263 , n251264 , n251265 , 
     n251266 , n251267 , n251268 , n251269 , n251270 , n251271 , n251272 , n251273 , n251274 , n251275 , 
     n251276 , n251277 , n251278 , n251279 , n251280 , n251281 , n251282 , n251283 , n251284 , n251285 , 
     n251286 , n251287 , n251288 , n251289 , n251290 , n251291 , n251292 , n251293 , n251294 , n251295 , 
     n251296 , n251297 , n251298 , n251299 , n251300 , n251301 , n251302 , n251303 , n251304 , n251305 , 
     n251306 , n251307 , n251308 , n251309 , n251310 , n251311 , n251312 , n251313 , n251314 , n251315 , 
     n251316 , n251317 , n251318 , n251319 , n251320 , n251321 , n251322 , n251323 , n251324 , n251325 , 
     n251326 , n251327 , n251328 , n251329 , n251330 , n251331 , n251332 , n251333 , n251334 , n251335 , 
     n251336 , n251337 , n251338 , n251339 , n251340 , n251341 , n251342 , n251343 , n251344 , n251345 , 
     n251346 , n251347 , n251348 , n251349 , n251350 , n251351 , n251352 , n251353 , n251354 , n251355 , 
     n251356 , n251357 , n251358 , n251359 , n251360 , n251361 , n251362 , n251363 , n251364 , n251365 , 
     n251366 , n251367 , n251368 , n251369 , n251370 , n251371 , n251372 , n251373 , n251374 , n251375 , 
     n251376 , n251377 , n251378 , n251379 , n251380 , n251381 , n251382 , n251383 , n251384 , n251385 , 
     n251386 , n251387 , n251388 , n251389 , n251390 , n251391 , n251392 , n251393 , n251394 , n251395 , 
     n251396 , n251397 , n251398 , n251399 , n251400 , n251401 , n251402 , n251403 , n251404 , n251405 , 
     n251406 , n251407 , n251408 , n251409 , n251410 , n251411 , n251412 , n251413 , n251414 , n251415 , 
     n251416 , n251417 , n251418 , n251419 , n251420 , n251421 , n251422 , n251423 , n251424 , n251425 , 
     n251426 , n251427 , n251428 , n251429 , n251430 , n251431 , n251432 , n251433 , n251434 , n251435 , 
     n251436 , n251437 , n251438 , n251439 , n251440 , n251441 , n251442 , n251443 , n251444 , n251445 , 
     n251446 , n251447 , n251448 , n251449 , n251450 , n251451 , n251452 , n251453 , n251454 , n251455 , 
     n251456 , n251457 , n251458 , n251459 , n251460 , n251461 , n251462 , n251463 , n251464 , n251465 , 
     n251466 , n251467 , n251468 , n251469 , n251470 , n251471 , n251472 , n251473 , n251474 , n251475 , 
     n251476 , n251477 , n251478 , n251479 , n251480 , n251481 , n251482 , n251483 , n251484 , n251485 , 
     n251486 , n251487 , n251488 , n251489 , n251490 , n251491 , n251492 , n251493 , n251494 , n251495 , 
     n251496 , n251497 , n251498 , n251499 , n251500 , n251501 , n251502 , n251503 , n251504 , n251505 , 
     n251506 , n251507 , n251508 , n251509 , n251510 , n251511 , n251512 , n251513 , n251514 , n251515 , 
     n251516 , n251517 , n251518 , n251519 , n251520 , n251521 , n251522 , n251523 , n251524 , n251525 , 
     n251526 , n251527 , n251528 , n251529 , n251530 , n251531 , n251532 , n251533 , n251534 , n251535 , 
     n251536 , n251537 , n251538 , n251539 , n251540 , n251541 , n251542 , n251543 , n251544 , n251545 , 
     n251546 , n251547 , n251548 , n251549 , n251550 , n251551 , n251552 , n251553 , n251554 , n251555 , 
     n251556 , n251557 , n251558 , n251559 , n251560 , n251561 , n251562 , n251563 , n251564 , n251565 , 
     n251566 , n251567 , n251568 , n251569 , n251570 , n251571 , n251572 , n251573 , n251574 , n251575 , 
     n251576 , n251577 , n251578 , n251579 , n251580 , n251581 , n251582 , n251583 , n251584 , n251585 , 
     n251586 , n251587 , n251588 , n251589 , n251590 , n251591 , n251592 , n251593 , n251594 , n251595 , 
     n251596 , n251597 , n251598 , n251599 , n251600 , n251601 , n251602 , n251603 , n251604 , n251605 , 
     n251606 , n251607 , n251608 , n251609 , n251610 , n251611 , n251612 , n251613 , n251614 , n251615 , 
     n251616 , n251617 , n251618 , n251619 , n251620 , n251621 , n251622 , n251623 , n251624 , n251625 , 
     n251626 , n251627 , n251628 , n251629 , n251630 , n251631 , n251632 , n251633 , n251634 , n251635 , 
     n251636 , n251637 , n251638 , n251639 , n251640 , n251641 , n251642 , n251643 , n251644 , n251645 , 
     n251646 , n251647 , n251648 , n251649 , n251650 , n251651 , n251652 , n251653 , n251654 , n251655 , 
     n251656 , n251657 , n251658 , n251659 , n251660 , n251661 , n251662 , n251663 , n251664 , n251665 , 
     n251666 , n251667 , n251668 , n251669 , n251670 , n251671 , n251672 , n251673 , n251674 , n251675 , 
     n251676 , n251677 , n251678 , n251679 , n251680 , n251681 , n251682 , n251683 , n251684 , n251685 , 
     n251686 , n251687 , n251688 , n251689 , n251690 , n251691 , n251692 , n251693 , n251694 , n251695 , 
     n251696 , n251697 , n251698 , n251699 , n251700 , n251701 , n251702 , n251703 , n251704 , n251705 , 
     n251706 , n251707 , n251708 , n251709 , n251710 , n251711 , n251712 , n251713 , n251714 , n251715 , 
     n251716 , n251717 , n251718 , n251719 , n251720 , n251721 , n251722 , n251723 , n251724 , n251725 , 
     n251726 , n251727 , n251728 , n251729 , n251730 , n251731 , n251732 , n251733 , n251734 , n251735 , 
     n251736 , n251737 , n251738 , n251739 , n251740 , n251741 , n251742 , n251743 , n251744 , n251745 , 
     n251746 , n251747 , n251748 , n251749 , n251750 , n251751 , n251752 , n251753 , n251754 , n251755 , 
     n251756 , n251757 , n251758 , n251759 , n251760 , n251761 , n251762 , n251763 , n251764 , n251765 , 
     n251766 , n251767 , n251768 , n251769 , n251770 , n251771 , n251772 , n251773 , n251774 , n251775 , 
     n251776 , n251777 , n251778 , n251779 , n251780 , n251781 , n251782 , n251783 , n251784 , n251785 , 
     n251786 , n251787 , n251788 , n251789 , n251790 , n251791 , n251792 , n251793 , n251794 , n251795 , 
     n251796 , n251797 , n251798 , n251799 , n251800 , n251801 , n251802 , n251803 , n251804 , n251805 , 
     n251806 , n251807 , n251808 , n251809 , n251810 , n251811 , n251812 , n251813 , n251814 , n251815 , 
     n251816 , n251817 , n251818 , n251819 , n251820 , n251821 , n251822 , n251823 , n251824 , n251825 , 
     n251826 , n251827 , n251828 , n251829 , n251830 , n251831 , n251832 , n251833 , n251834 , n251835 , 
     n251836 , n251837 , n251838 , n251839 , n251840 , n251841 , n251842 , n251843 , n251844 , n251845 , 
     n251846 , n251847 , n251848 , n251849 , n251850 , n251851 , n251852 , n251853 , n251854 , n251855 , 
     n251856 , n251857 , n251858 , n251859 , n251860 , n251861 , n251862 , n251863 , n251864 , n251865 , 
     n251866 , n251867 , n251868 , n251869 , n251870 , n251871 , n251872 , n251873 , n251874 , n251875 , 
     n251876 , n251877 , n251878 , n251879 , n251880 , n251881 , n251882 , n251883 , n251884 , n251885 , 
     n251886 , n251887 , n251888 , n251889 , n251890 , n251891 , n251892 , n251893 , n251894 , n251895 , 
     n251896 , n251897 , n251898 , n251899 , n251900 , n251901 , n251902 , n251903 , n251904 , n251905 , 
     n251906 , n251907 , n251908 , n251909 , n251910 , n251911 , n251912 , n251913 , n251914 , n251915 , 
     n251916 , n251917 , n251918 , n251919 , n251920 , n251921 , n251922 , n251923 , n251924 , n251925 , 
     n251926 , n251927 , n251928 , n251929 , n251930 , n251931 , n251932 , n251933 , n251934 , n251935 , 
     n251936 , n251937 , n251938 , n251939 , n251940 , n251941 , n251942 , n251943 , n251944 , n251945 , 
     n251946 , n251947 , n251948 , n251949 , n251950 , n251951 , n251952 , n251953 , n251954 , n251955 , 
     n251956 , n251957 , n251958 , n251959 , n251960 , n251961 , n251962 , n251963 , n251964 , n251965 , 
     n251966 , n251967 , n251968 , n251969 , n251970 , n251971 , n251972 , n251973 , n251974 , n251975 , 
     n251976 , n251977 , n251978 , n251979 , n251980 , n251981 , n251982 , n251983 , n251984 , n251985 , 
     n251986 , n251987 , n251988 , n251989 , n251990 , n251991 , n251992 , n251993 , n251994 , n251995 , 
     n251996 , n251997 , n251998 , n251999 , n252000 , n252001 , n252002 , n252003 , n252004 , n252005 , 
     n252006 , n252007 , n252008 , n252009 , n252010 , n252011 , n252012 , n252013 , n252014 , n252015 , 
     n252016 , n252017 , n252018 , n252019 , n252020 , n252021 , n252022 , n252023 , n252024 , n252025 , 
     n252026 , n252027 , n252028 , n252029 , n252030 , n252031 , n252032 , n252033 , n252034 , n252035 , 
     n252036 , n252037 , n252038 , n252039 , n252040 , n252041 , n252042 , n252043 , n252044 , n252045 , 
     n252046 , n252047 , n252048 , n252049 , n252050 , n252051 , n252052 , n252053 , n252054 , n252055 , 
     n252056 , n252057 , n252058 , n252059 , n252060 , n252061 , n252062 , n252063 , n252064 , n252065 , 
     n252066 , n252067 , n252068 , n252069 , n252070 , n252071 , n252072 , n252073 , n252074 , n252075 , 
     n252076 , n252077 , n252078 , n252079 , n252080 , n252081 , n252082 , n252083 , n252084 , n252085 , 
     n252086 , n252087 , n252088 , n252089 , n252090 , n252091 , n252092 , n252093 , n252094 , n252095 , 
     n252096 , n252097 , n252098 , n252099 , n252100 , n252101 , n252102 , n252103 , n252104 , n252105 , 
     n252106 , n252107 , n252108 , n252109 , n252110 , n252111 , n252112 , n252113 , n252114 , n252115 , 
     n252116 , n252117 , n252118 , n252119 , n252120 , n252121 , n252122 , n252123 , n252124 , n252125 , 
     n252126 , n252127 , n252128 , n252129 , n252130 , n252131 , n252132 , n252133 , n252134 , n252135 , 
     n252136 , n252137 , n252138 , n252139 , n252140 , n252141 , n252142 , n252143 , n252144 , n252145 , 
     n252146 , n252147 , n252148 , n252149 , n252150 , n252151 , n252152 , n252153 , n252154 , n252155 , 
     n252156 , n252157 , n252158 , n252159 , n252160 , n252161 , n252162 , n252163 , n252164 , n252165 , 
     n252166 , n252167 , n252168 , n252169 , n252170 , n252171 , n252172 , n252173 , n252174 , n252175 , 
     n252176 , n252177 , n252178 , n252179 , n252180 , n252181 , n252182 , n252183 , n252184 , n252185 , 
     n252186 , n252187 , n252188 , n252189 , n252190 , n252191 , n252192 , n252193 , n252194 , n252195 , 
     n252196 , n252197 , n252198 , n252199 , n252200 , n252201 , n252202 , n252203 , n252204 , n252205 , 
     n252206 , n252207 , n252208 , n252209 , n252210 , n252211 , n252212 , n252213 , n252214 , n252215 , 
     n252216 , n252217 , n252218 , n252219 , n252220 , n252221 , n252222 , n252223 , n252224 , n252225 , 
     n252226 , n252227 , n252228 , n252229 , n252230 , n252231 , n252232 , n252233 , n252234 , n252235 , 
     n252236 , n252237 , n252238 , n252239 , n252240 , n252241 , n252242 , n252243 , n252244 , n252245 , 
     n252246 , n252247 , n252248 , n252249 , n252250 , n252251 , n252252 , n252253 , n252254 , n252255 , 
     n252256 , n252257 , n252258 , n252259 , n252260 , n252261 , n252262 , n252263 , n252264 , n252265 , 
     n252266 , n252267 , n252268 , n252269 , n252270 , n252271 , n252272 , n252273 , n252274 , n252275 , 
     n252276 , n252277 , n252278 , n252279 , n252280 , n252281 , n252282 , n252283 , n252284 , n252285 , 
     n252286 , n252287 , n252288 , n252289 , n252290 , n252291 , n252292 , n252293 , n252294 , n252295 , 
     n252296 , n252297 , n252298 , n252299 , n252300 , n252301 , n252302 , n252303 , n252304 , n252305 , 
     n252306 , n252307 , n252308 , n252309 , n252310 , n252311 , n252312 , n252313 , n252314 , n252315 , 
     n252316 , n252317 , n252318 , n252319 , n252320 , n252321 , n252322 , n252323 , n252324 , n252325 , 
     n252326 , n252327 , n252328 , n252329 , n252330 , n252331 , n252332 , n252333 , n252334 , n252335 , 
     n252336 , n252337 , n252338 , n252339 , n252340 , n252341 , n252342 , n252343 , n252344 , n252345 , 
     n252346 , n252347 , n252348 , n252349 , n252350 , n252351 , n252352 , n252353 , n252354 , n252355 , 
     n252356 , n252357 , n252358 , n252359 , n252360 , n252361 , n252362 , n252363 , n252364 , n252365 , 
     n252366 , n252367 , n252368 , n252369 , n252370 , n252371 , n252372 , n252373 , n252374 , n252375 , 
     n252376 , n252377 , n252378 , n252379 , n252380 , n252381 , n252382 , n252383 , n252384 , n252385 , 
     n252386 , n252387 , n252388 , n252389 , n252390 , n252391 , n252392 , n252393 , n252394 , n252395 , 
     n252396 , n252397 , n252398 , n252399 , n252400 , n252401 , n252402 , n252403 , n252404 , n252405 , 
     n252406 , n252407 , n252408 , n252409 , n252410 , n252411 , n252412 , n252413 , n252414 , n252415 , 
     n252416 , n252417 , n252418 , n252419 , n252420 , n252421 , n252422 , n252423 , n252424 , n252425 , 
     n252426 , n252427 , n252428 , n252429 , n252430 , n252431 , n252432 , n252433 , n252434 , n252435 , 
     n252436 , n252437 , n252438 , n252439 , n252440 , n252441 , n252442 , n252443 , n252444 , n252445 , 
     n252446 , n252447 , n252448 , n252449 , n252450 , n252451 , n252452 , n252453 , n252454 , n252455 , 
     n252456 , n252457 , n252458 , n252459 , n252460 , n252461 , n252462 , n252463 , n252464 , n252465 , 
     n252466 , n252467 , n252468 , n252469 , n252470 , n252471 , n252472 , n252473 , n252474 , n252475 , 
     n252476 , n252477 , n252478 , n252479 , n252480 , n252481 , n252482 , n252483 , n252484 , n252485 , 
     n252486 , n252487 , n252488 , n252489 , n252490 , n252491 , n252492 , n252493 , n252494 , n252495 , 
     n252496 , n252497 , n252498 , n252499 , n252500 , n252501 , n252502 , n252503 , n252504 , n252505 , 
     n252506 , n252507 , n252508 , n252509 , n252510 , n252511 , n252512 , n252513 , n252514 , n252515 , 
     n252516 , n252517 , n252518 , n252519 , n252520 , n252521 , n252522 , n252523 , n252524 , n252525 , 
     n252526 , n252527 , n252528 , n252529 , n252530 , n252531 , n252532 , n252533 , n252534 , n252535 , 
     n252536 , n252537 , n252538 , n252539 , n252540 , n252541 , n252542 , n252543 , n252544 , n252545 , 
     n252546 , n252547 , n252548 , n252549 , n252550 , n252551 , n252552 , n252553 , n252554 , n252555 , 
     n252556 , n252557 , n252558 , n252559 , n252560 , n252561 , n252562 , n252563 , n252564 , n252565 , 
     n252566 , n252567 , n252568 , n252569 , n252570 , n252571 , n252572 , n252573 , n252574 , n252575 , 
     n252576 , n252577 , n252578 , n252579 , n252580 , n252581 , n252582 , n252583 , n252584 , n252585 , 
     n252586 , n252587 , n252588 , n252589 , n252590 , n252591 , n252592 , n252593 , n252594 , n252595 , 
     n252596 , n252597 , n252598 , n252599 , n252600 , n252601 , n252602 , n252603 , n252604 , n252605 , 
     n252606 , n252607 , n252608 , n252609 , n252610 , n252611 , n252612 , n252613 , n252614 , n252615 , 
     n252616 , n252617 , n252618 , n252619 , n252620 , n252621 , n252622 , n252623 , n252624 , n252625 , 
     n252626 , n252627 , n252628 , n252629 , n252630 , n252631 , n252632 , n252633 , n252634 , n252635 , 
     n252636 , n252637 , n252638 , n252639 , n252640 , n252641 , n252642 , n252643 , n252644 , n252645 , 
     n252646 , n252647 , n252648 , n252649 , n252650 , n252651 , n252652 , n252653 , n252654 , n252655 , 
     n252656 , n252657 , n252658 , n252659 , n252660 , n252661 , n252662 , n252663 , n252664 , n252665 , 
     n252666 , n252667 , n252668 , n252669 , n252670 , n252671 , n252672 , n252673 , n252674 , n252675 , 
     n252676 , n252677 , n252678 , n252679 , n252680 , n252681 , n252682 , n252683 , n252684 , n252685 , 
     n252686 , n252687 , n252688 , n252689 , n252690 , n252691 , n252692 , n252693 , n252694 , n252695 , 
     n252696 , n252697 , n252698 , n252699 , n252700 , n252701 , n252702 , n252703 , n252704 , n252705 , 
     n252706 , n252707 , n252708 , n252709 , n252710 , n252711 , n252712 , n252713 , n252714 , n252715 , 
     n252716 , n252717 , n252718 , n252719 , n252720 , n252721 , n252722 , n252723 , n252724 , n252725 , 
     n252726 , n252727 , n252728 , n252729 , n252730 , n252731 , n252732 , n252733 , n252734 , n252735 , 
     n252736 , n252737 , n252738 , n252739 , n252740 , n252741 , n252742 , n252743 , n252744 , n252745 , 
     n252746 , n252747 , n252748 , n252749 , n252750 , n252751 , n252752 , n252753 , n252754 , n252755 , 
     n252756 , n252757 , n252758 , n252759 , n252760 , n252761 , n252762 , n252763 , n252764 , n252765 , 
     n252766 , n252767 , n252768 , n252769 , n252770 , n252771 , n252772 , n252773 , n252774 , n252775 , 
     n252776 , n252777 , n252778 , n252779 , n252780 , n252781 , n252782 , n252783 , n252784 , n252785 , 
     n252786 , n252787 , n252788 , n252789 , n252790 , n252791 , n252792 , n252793 , n252794 , n252795 , 
     n252796 , n252797 , n252798 , n252799 , n252800 , n252801 , n252802 , n252803 , n252804 , n252805 , 
     n252806 , n252807 , n252808 , n252809 , n252810 , n252811 , n252812 , n252813 , n252814 , n252815 , 
     n252816 , n252817 , n252818 , n252819 , n252820 , n252821 , n252822 , n252823 , n252824 , n252825 , 
     n252826 , n252827 , n252828 , n252829 , n252830 , n252831 , n252832 , n252833 , n252834 , n252835 , 
     n252836 , n252837 , n252838 , n252839 , n252840 , n252841 , n252842 , n252843 , n252844 , n252845 , 
     n252846 , n252847 , n252848 , n252849 , n252850 , n252851 , n252852 , n252853 , n252854 , n252855 , 
     n252856 , n252857 , n252858 , n252859 , n252860 , n252861 , n252862 , n252863 , n252864 , n252865 , 
     n252866 , n252867 , n252868 , n252869 , n252870 , n252871 , n252872 , n252873 , n252874 , n252875 , 
     n252876 , n252877 , n252878 , n252879 , n252880 , n252881 , n252882 , n252883 , n252884 , n252885 , 
     n252886 , n252887 , n252888 , n252889 , n252890 , n252891 , n252892 , n252893 , n252894 , n252895 , 
     n252896 , n252897 , n252898 , n252899 , n252900 , n252901 , n252902 , n252903 , n252904 , n252905 , 
     n252906 , n252907 , n252908 , n252909 , n252910 , n252911 , n252912 , n252913 , n252914 , n252915 , 
     n252916 , n252917 , n252918 , n252919 , n252920 , n252921 , n252922 , n252923 , n252924 , n252925 , 
     n252926 , n252927 , n252928 , n252929 , n252930 , n252931 , n252932 , n252933 , n252934 , n252935 , 
     n252936 , n252937 , n252938 , n252939 , n252940 , n252941 , n252942 , n252943 , n252944 , n252945 , 
     n252946 , n252947 , n252948 , n252949 , n252950 , n252951 , n252952 , n252953 , n252954 , n252955 , 
     n252956 , n252957 , n252958 , n252959 , n252960 , n252961 , n252962 , n252963 , n252964 , n252965 , 
     n252966 , n252967 , n252968 , n252969 , n252970 , n252971 , n252972 , n252973 , n252974 , n252975 , 
     n252976 , n252977 , n252978 , n252979 , n252980 , n252981 , n252982 , n252983 , n252984 , n252985 , 
     n252986 , n252987 , n252988 , n252989 , n252990 , n252991 , n252992 , n252993 , n252994 , n252995 , 
     n252996 , n252997 , n252998 , n252999 , n253000 , n253001 , n253002 , n253003 , n253004 , n253005 , 
     n253006 , n253007 , n253008 , n253009 , n253010 , n253011 , n253012 , n253013 , n253014 , n253015 , 
     n253016 , n253017 , n253018 , n253019 , n253020 , n253021 , n253022 , n253023 , n253024 , n253025 , 
     n253026 , n253027 , n253028 , n253029 , n253030 , n253031 , n253032 , n253033 , n253034 , n253035 , 
     n253036 , n253037 , n253038 , n253039 , n253040 , n253041 , n253042 , n253043 , n253044 , n253045 , 
     n253046 , n253047 , n253048 , n253049 , n253050 , n253051 , n253052 , n253053 , n253054 , n253055 , 
     n253056 , n253057 , n253058 , n253059 , n253060 , n253061 , n253062 , n253063 , n253064 , n253065 , 
     n253066 , n253067 , n253068 , n253069 , n253070 , n253071 , n253072 , n253073 , n253074 , n253075 , 
     n253076 , n253077 , n253078 , n253079 , n253080 , n253081 , n253082 , n253083 , n253084 , n253085 , 
     n253086 , n253087 , n253088 , n253089 , n253090 , n253091 , n253092 , n253093 , n253094 , n253095 , 
     n253096 , n253097 , n253098 , n253099 , n253100 , n253101 , n253102 , n253103 , n253104 , n253105 , 
     n253106 , n253107 , n253108 , n253109 , n253110 , n253111 , n253112 , n253113 , n253114 , n253115 , 
     n253116 , n253117 , n253118 , n253119 , n253120 , n253121 , n253122 , n253123 , n253124 , n253125 , 
     n253126 , n253127 , n253128 , n253129 , n253130 , n253131 , n253132 , n253133 , n253134 , n253135 , 
     n253136 , n253137 , n253138 , n253139 , n253140 , n253141 , n253142 , n253143 , n253144 , n253145 , 
     n253146 , n253147 , n253148 , n253149 , n253150 , n253151 , n253152 , n253153 , n253154 , n253155 , 
     n253156 , n253157 , n253158 , n253159 , n253160 , n253161 , n253162 , n253163 , n253164 , n253165 , 
     n253166 , n253167 , n253168 , n253169 , n253170 , n253171 , n253172 , n253173 , n253174 , n253175 , 
     n253176 , n253177 , n253178 , n253179 , n253180 , n253181 , n253182 , n253183 , n253184 , n253185 , 
     n253186 , n253187 , n253188 , n253189 , n253190 , n253191 , n253192 , n253193 , n253194 , n253195 , 
     n253196 , n253197 , n253198 , n253199 , n253200 , n253201 , n253202 , n253203 , n253204 , n253205 , 
     n253206 , n253207 , n253208 , n253209 , n253210 , n253211 , n253212 , n253213 , n253214 , n253215 , 
     n253216 , n253217 , n253218 , n253219 , n253220 , n253221 , n253222 , n253223 , n253224 , n253225 , 
     n253226 , n253227 , n253228 , n253229 , n253230 , n253231 , n253232 , n253233 , n253234 , n253235 , 
     n253236 , n253237 , n253238 , n253239 , n253240 , n253241 , n253242 , n253243 , n253244 , n253245 , 
     n253246 , n253247 , n253248 , n253249 , n253250 , n253251 , n253252 , n253253 , n253254 , n253255 , 
     n253256 , n253257 , n253258 , n253259 , n253260 , n253261 , n253262 , n253263 , n253264 , n253265 , 
     n253266 , n253267 , n253268 , n253269 , n253270 , n253271 , n253272 , n253273 , n253274 , n253275 , 
     n253276 , n253277 , n253278 , n253279 , n253280 , n253281 , n253282 , n253283 , n253284 , n253285 , 
     n253286 , n253287 , n253288 , n253289 , n253290 , n253291 , n253292 , n253293 , n253294 , n253295 , 
     n253296 , n253297 , n253298 , n253299 , n253300 , n253301 , n253302 , n253303 , n253304 , n253305 , 
     n253306 , n253307 , n253308 , n253309 , n253310 , n253311 , n253312 , n253313 , n253314 , n253315 , 
     n253316 , n253317 , n253318 , n253319 , n253320 , n253321 , n253322 , n253323 , n253324 , n253325 , 
     n253326 , n253327 , n253328 , n253329 , n253330 , n253331 , n253332 , n253333 , n253334 , n253335 , 
     n253336 , n253337 , n253338 , n253339 , n253340 , n253341 , n253342 , n253343 , n253344 , n253345 , 
     n253346 , n253347 , n253348 , n253349 , n253350 , n253351 , n253352 , n253353 , n253354 , n253355 , 
     n253356 , n253357 , n253358 , n253359 , n253360 , n253361 , n253362 , n253363 , n253364 , n253365 , 
     n253366 , n253367 , n253368 , n253369 , n253370 , n253371 , n253372 , n253373 , n253374 , n253375 , 
     n253376 , n253377 , n253378 , n253379 , n253380 , n253381 , n253382 , n253383 , n253384 , n253385 , 
     n253386 , n253387 , n253388 , n253389 , n253390 , n253391 , n253392 , n253393 , n253394 , n253395 , 
     n253396 , n253397 , n253398 , n253399 , n253400 , n253401 , n253402 , n253403 , n253404 , n253405 , 
     n253406 , n253407 , n253408 , n253409 , n253410 , n253411 , n253412 , n253413 , n253414 , n253415 , 
     n253416 , n253417 , n253418 , n253419 , n253420 , n253421 , n253422 , n253423 , n253424 , n253425 , 
     n253426 , n253427 , n253428 , n253429 , n253430 , n253431 , n253432 , n253433 , n253434 , n253435 , 
     n253436 , n253437 , n253438 , n253439 , n253440 , n253441 , n253442 , n253443 , n253444 , n253445 , 
     n253446 , n253447 , n253448 , n253449 , n253450 , n253451 , n253452 , n253453 , n253454 , n253455 , 
     n253456 , n253457 , n253458 , n253459 , n253460 , n253461 , n253462 , n253463 , n253464 , n253465 , 
     n253466 , n253467 , n253468 , n253469 , n253470 , n253471 , n253472 , n253473 , n253474 , n253475 , 
     n253476 , n253477 , n253478 , n253479 , n253480 , n253481 , n253482 , n253483 , n253484 , n253485 , 
     n253486 , n253487 , n253488 , n253489 , n253490 , n253491 , n253492 , n253493 , n253494 , n253495 , 
     n253496 , n253497 , n253498 , n253499 , n253500 , n253501 , n253502 , n253503 , n253504 , n253505 , 
     n253506 , n253507 , n253508 , n253509 , n253510 , n253511 , n253512 , n253513 , n253514 , n253515 , 
     n253516 , n253517 , n253518 , n253519 , n253520 , n253521 , n253522 , n253523 , n253524 , n253525 , 
     n253526 , n253527 , n253528 , n253529 , n253530 , n253531 , n253532 , n253533 , n253534 , n253535 , 
     n253536 , n253537 , n253538 , n253539 , n253540 , n253541 , n253542 , n253543 , n253544 , n253545 , 
     n253546 , n253547 , n253548 , n253549 , n253550 , n253551 , n253552 , n253553 , n253554 , n253555 , 
     n253556 , n253557 , n253558 , n253559 , n253560 , n253561 , n253562 , n253563 , n253564 , n253565 , 
     n253566 , n253567 , n253568 , n253569 , n253570 , n253571 , n253572 , n253573 , n253574 , n253575 , 
     n253576 , n253577 , n253578 , n253579 , n253580 , n253581 , n253582 , n253583 , n253584 , n253585 , 
     n253586 , n253587 , n253588 , n253589 , n253590 , n253591 , n253592 , n253593 , n253594 , n253595 , 
     n253596 , n253597 , n253598 , n253599 , n253600 , n253601 , n253602 , n253603 , n253604 , n253605 , 
     n253606 , n253607 , n253608 , n253609 , n253610 , n253611 , n253612 , n253613 , n253614 , n253615 , 
     n253616 , n253617 , n253618 , n253619 , n253620 , n253621 , n253622 , n253623 , n253624 , n253625 , 
     n253626 , n253627 , n253628 , n253629 , n253630 , n253631 , n253632 , n253633 , n253634 , n253635 , 
     n253636 , n253637 , n253638 , n253639 , n253640 , n253641 , n253642 , n253643 , n253644 , n253645 , 
     n253646 , n253647 , n253648 , n253649 , n253650 , n253651 , n253652 , n253653 , n253654 , n253655 , 
     n253656 , n253657 , n253658 , n253659 , n253660 , n253661 , n253662 , n253663 , n253664 , n253665 , 
     n253666 , n253667 , n253668 , n253669 , n253670 , n253671 , n253672 , n253673 , n253674 , n253675 , 
     n253676 , n253677 , n253678 , n253679 , n253680 , n253681 , n253682 , n253683 , n253684 , n253685 , 
     n253686 , n253687 , n253688 , n253689 , n253690 , n253691 , n253692 , n253693 , n253694 , n253695 , 
     n253696 , n253697 , n253698 , n253699 , n253700 , n253701 , n253702 , n253703 , n253704 , n253705 , 
     n253706 , n253707 , n253708 , n253709 , n253710 , n253711 , n253712 , n253713 , n253714 , n253715 , 
     n253716 , n253717 , n253718 , n253719 , n253720 , n253721 , n253722 , n253723 , n253724 , n253725 , 
     n253726 , n253727 , n253728 , n253729 , n253730 , n253731 , n253732 , n253733 , n253734 , n253735 , 
     n253736 , n253737 , n253738 , n253739 , n253740 , n253741 , n253742 , n253743 , n253744 , n253745 , 
     n253746 , n253747 , n253748 , n253749 , n253750 , n253751 , n253752 , n253753 , n253754 , n253755 , 
     n253756 , n253757 , n253758 , n253759 , n253760 , n253761 , n253762 , n253763 , n253764 , n253765 , 
     n253766 , n253767 , n253768 , n253769 , n253770 , n253771 , n253772 , n253773 , n253774 , n253775 , 
     n253776 , n253777 , n253778 , n253779 , n253780 , n253781 , n253782 , n253783 , n253784 , n253785 , 
     n253786 , n253787 , n253788 , n253789 , n253790 , n253791 , n253792 , n253793 , n253794 , n253795 , 
     n253796 , n253797 , n253798 , n253799 , n253800 , n253801 , n253802 , n253803 , n253804 , n253805 , 
     n253806 , n253807 , n253808 , n253809 , n253810 , n253811 , n253812 , n253813 , n253814 , n253815 , 
     n253816 , n253817 , n253818 , n253819 , n253820 , n253821 , n253822 , n253823 , n253824 , n253825 , 
     n253826 , n253827 , n253828 , n253829 , n253830 , n253831 , n253832 , n253833 , n253834 , n253835 , 
     n253836 , n253837 , n253838 , n253839 , n253840 , n253841 , n253842 , n253843 , n253844 , n253845 , 
     n253846 , n253847 , n253848 , n253849 , n253850 , n253851 , n253852 , n253853 , n253854 , n253855 , 
     n253856 , n253857 , n253858 , n253859 , n253860 , n253861 , n253862 , n253863 , n253864 , n253865 , 
     n253866 , n253867 , n253868 , n253869 , n253870 , n253871 , n253872 , n253873 , n253874 , n253875 , 
     n253876 , n253877 , n253878 , n253879 , n253880 , n253881 , n253882 , n253883 , n253884 , n253885 , 
     n253886 , n253887 , n253888 , n253889 , n253890 , n253891 , n253892 , n253893 , n253894 , n253895 , 
     n253896 , n253897 , n253898 , n253899 , n253900 , n253901 , n253902 , n253903 , n253904 , n253905 , 
     n253906 , n253907 , n253908 , n253909 , n253910 , n253911 , n253912 , n253913 , n253914 , n253915 , 
     n253916 , n253917 , n253918 , n253919 , n253920 , n253921 , n253922 , n253923 , n253924 , n253925 , 
     n253926 , n253927 , n253928 , n253929 , n253930 , n253931 , n253932 , n253933 , n253934 , n253935 , 
     n253936 , n253937 , n253938 , n253939 , n253940 , n253941 , n253942 , n253943 , n253944 , n253945 , 
     n253946 , n253947 , n253948 , n253949 , n253950 , n253951 , n253952 , n253953 , n253954 , n253955 , 
     n253956 , n253957 , n253958 , n253959 , n253960 , n253961 , n253962 , n253963 , n253964 , n253965 , 
     n253966 , n253967 , n253968 , n253969 , n253970 , n253971 , n253972 , n253973 , n253974 , n253975 , 
     n253976 , n253977 , n253978 , n253979 , n253980 , n253981 , n253982 , n253983 , n253984 , n253985 , 
     n253986 , n253987 , n253988 , n253989 , n253990 , n253991 , n253992 , n253993 , n253994 , n253995 , 
     n253996 , n253997 , n253998 , n253999 , n254000 , n254001 , n254002 , n254003 , n254004 , n254005 , 
     n254006 , n254007 , n254008 , n254009 , n254010 , n254011 , n254012 , n254013 , n254014 , n254015 , 
     n254016 , n254017 , n254018 , n254019 , n254020 , n254021 , n254022 , n254023 , n254024 , n254025 , 
     n254026 , n254027 , n254028 , n254029 , n254030 , n254031 , n254032 , n254033 , n254034 , n254035 , 
     n254036 , n254037 , n254038 , n254039 , n254040 , n254041 , n254042 , n254043 , n254044 , n254045 , 
     n254046 , n254047 , n254048 , n254049 , n254050 , n254051 , n254052 , n254053 , n254054 , n254055 , 
     n254056 , n254057 , n254058 , n254059 , n254060 , n254061 , n254062 , n254063 , n254064 , n254065 , 
     n254066 , n254067 , n254068 , n254069 , n254070 , n254071 , n254072 , n254073 , n254074 , n254075 , 
     n254076 , n254077 , n254078 , n254079 , n254080 , n254081 , n254082 , n254083 , n254084 , n254085 , 
     n254086 , n254087 , n254088 , n254089 , n254090 , n254091 , n254092 , n254093 , n254094 , n254095 , 
     n254096 , n254097 , n254098 , n254099 , n254100 , n254101 , n254102 , n254103 , n254104 , n254105 , 
     n254106 , n254107 , n254108 , n254109 , n254110 , n254111 , n254112 , n254113 , n254114 , n254115 , 
     n254116 , n254117 , n254118 , n254119 , n254120 , n254121 , n254122 , n254123 , n254124 , n254125 , 
     n254126 , n254127 , n254128 , n254129 , n254130 , n254131 , n254132 , n254133 , n254134 , n254135 , 
     n254136 , n254137 , n254138 , n254139 , n254140 , n254141 , n254142 , n254143 , n254144 , n254145 , 
     n254146 , n254147 , n254148 , n254149 , n254150 , n254151 , n254152 , n254153 , n254154 , n254155 , 
     n254156 , n254157 , n254158 , n254159 , n254160 , n254161 , n254162 , n254163 , n254164 , n254165 , 
     n254166 , n254167 , n254168 , n254169 , n254170 , n254171 , n254172 , n254173 , n254174 , n254175 , 
     n254176 , n254177 , n254178 , n254179 , n254180 , n254181 , n254182 , n254183 , n254184 , n254185 , 
     n254186 , n254187 , n254188 , n254189 , n254190 , n254191 , n254192 , n254193 , n254194 , n254195 , 
     n254196 , n254197 , n254198 , n254199 , n254200 , n254201 , n254202 , n254203 , n254204 , n254205 , 
     n254206 , n254207 , n254208 , n254209 , n254210 , n254211 , n254212 , n254213 , n254214 , n254215 , 
     n254216 , n254217 , n254218 , n254219 , n254220 , n254221 , n254222 , n254223 , n254224 , n254225 , 
     n254226 , n254227 , n254228 , n254229 , n254230 , n254231 , n254232 , n254233 , n254234 , n254235 , 
     n254236 , n254237 , n254238 , n254239 , n254240 , n254241 , n254242 , n254243 , n254244 , n254245 , 
     n254246 , n254247 , n254248 , n254249 , n254250 , n254251 , n254252 , n254253 , n254254 , n254255 , 
     n254256 , n254257 , n254258 , n254259 , n254260 , n254261 , n254262 , n254263 , n254264 , n254265 , 
     n254266 , n254267 , n254268 , n254269 , n254270 , n254271 , n254272 , n254273 , n254274 , n254275 , 
     n254276 , n254277 , n254278 , n254279 , n254280 , n254281 , n254282 , n254283 , n254284 , n254285 , 
     n254286 , n254287 , n254288 , n254289 , n254290 , n254291 , n254292 , n254293 , n254294 , n254295 , 
     n254296 , n254297 , n254298 , n254299 , n254300 , n254301 , n254302 , n254303 , n254304 , n254305 , 
     n254306 , n254307 , n254308 , n254309 , n254310 , n254311 , n254312 , n254313 , n254314 , n254315 , 
     n254316 , n254317 , n254318 , n254319 , n254320 , n254321 , n254322 , n254323 , n254324 , n254325 , 
     n254326 , n254327 , n254328 , n254329 , n254330 , n254331 , n254332 , n254333 , n254334 , n254335 , 
     n254336 , n254337 , n254338 , n254339 , n254340 , n254341 , n254342 , n254343 , n254344 , n254345 , 
     n254346 , n254347 , n254348 , n254349 , n254350 , n254351 , n254352 , n254353 , n254354 , n254355 , 
     n254356 , n254357 , n254358 , n254359 , n254360 , n254361 , n254362 , n254363 , n254364 , n254365 , 
     n254366 , n254367 , n254368 , n254369 , n254370 , n254371 , n254372 , n254373 , n254374 , n254375 , 
     n254376 , n254377 , n254378 , n254379 , n254380 , n254381 , n254382 , n254383 , n254384 , n254385 , 
     n254386 , n254387 , n254388 , n254389 , n254390 , n254391 , n254392 , n254393 , n254394 , n254395 , 
     n254396 , n254397 , n254398 , n254399 , n254400 , n254401 , n254402 , n254403 , n254404 , n254405 , 
     n254406 , n254407 , n254408 , n254409 , n254410 , n254411 , n254412 , n254413 , n254414 , n254415 , 
     n254416 , n254417 , n254418 , n254419 , n254420 , n254421 , n254422 , n254423 , n254424 , n254425 , 
     n254426 , n254427 , n254428 , n254429 , n254430 , n254431 , n254432 , n254433 , n254434 , n254435 , 
     n254436 , n254437 , n254438 , n254439 , n254440 , n254441 , n254442 , n254443 , n254444 , n254445 , 
     n254446 , n254447 , n254448 , n254449 , n254450 , n254451 , n254452 , n254453 , n254454 , n254455 , 
     n254456 , n254457 , n254458 , n254459 , n254460 , n254461 , n254462 , n254463 , n254464 , n254465 , 
     n254466 , n254467 , n254468 , n254469 , n254470 , n254471 , n254472 , n254473 , n254474 , n254475 , 
     n254476 , n254477 , n254478 , n254479 , n254480 , n254481 , n254482 , n254483 , n254484 , n254485 , 
     n254486 , n254487 , n254488 , n254489 , n254490 , n254491 , n254492 , n254493 , n254494 , n254495 , 
     n254496 , n254497 , n254498 , n254499 , n254500 , n254501 , n254502 , n254503 , n254504 , n254505 , 
     n254506 , n254507 , n254508 , n254509 , n254510 , n254511 , n254512 , n254513 , n254514 , n254515 , 
     n254516 , n254517 , n254518 , n254519 , n254520 , n254521 , n254522 , n254523 , n254524 , n254525 , 
     n254526 , n254527 , n254528 , n254529 , n254530 , n254531 , n254532 , n254533 , n254534 , n254535 , 
     n254536 , n254537 , n254538 , n254539 , n254540 , n254541 , n254542 , n254543 , n254544 , n254545 , 
     n254546 , n254547 , n254548 , n254549 , n254550 , n254551 , n254552 , n254553 , n254554 , n254555 , 
     n254556 , n254557 , n254558 , n254559 , n254560 , n254561 , n254562 , n254563 , n254564 , n254565 , 
     n254566 , n254567 , n254568 , n254569 , n254570 , n254571 , n254572 , n254573 , n254574 , n254575 , 
     n254576 , n254577 , n254578 , n254579 , n254580 , n254581 , n254582 , n254583 , n254584 , n254585 , 
     n254586 , n254587 , n254588 , n254589 , n254590 , n254591 , n254592 , n254593 , n254594 , n254595 , 
     n254596 , n254597 , n254598 , n254599 , n254600 , n254601 , n254602 , n254603 , n254604 , n254605 , 
     n254606 , n254607 , n254608 , n254609 , n254610 , n254611 , n254612 , n254613 , n254614 , n254615 , 
     n254616 , n254617 , n254618 , n254619 , n254620 , n254621 , n254622 , n254623 , n254624 , n254625 , 
     n254626 , n254627 , n254628 , n254629 , n254630 , n254631 , n254632 , n254633 , n254634 , n254635 , 
     n254636 , n254637 , n254638 , n254639 , n254640 , n254641 , n254642 , n254643 , n254644 , n254645 , 
     n254646 , n254647 , n254648 , n254649 , n254650 , n254651 , n254652 , n254653 , n254654 , n254655 , 
     n254656 , n254657 , n254658 , n254659 , n254660 , n254661 , n254662 , n254663 , n254664 , n254665 , 
     n254666 , n254667 , n254668 , n254669 , n254670 , n254671 , n254672 , n254673 , n254674 , n254675 , 
     n254676 , n254677 , n254678 , n254679 , n254680 , n254681 , n254682 , n254683 , n254684 , n254685 , 
     n254686 , n254687 , n254688 , n254689 , n254690 , n254691 , n254692 , n254693 , n254694 , n254695 , 
     n254696 , n254697 , n254698 , n254699 , n254700 , n254701 , n254702 , n254703 , n254704 , n254705 , 
     n254706 , n254707 , n254708 , n254709 , n254710 , n254711 , n254712 , n254713 , n254714 , n254715 , 
     n254716 , n254717 , n254718 , n254719 , n254720 , n254721 , n254722 , n254723 , n254724 , n254725 , 
     n254726 , n254727 , n254728 , n254729 , n254730 , n254731 , n254732 , n254733 , n254734 , n254735 , 
     n254736 , n254737 , n254738 , n254739 , n254740 , n254741 , n254742 , n254743 , n254744 , n254745 , 
     n254746 , n254747 , n254748 , n254749 , n254750 , n254751 , n254752 , n254753 , n254754 , n254755 , 
     n254756 , n254757 , n254758 , n254759 , n254760 , n254761 , n254762 , n254763 , n254764 , n254765 , 
     n254766 , n254767 , n254768 , n254769 , n254770 , n254771 , n254772 , n254773 , n254774 , n254775 , 
     n254776 , n254777 , n254778 , n254779 , n254780 , n254781 , n254782 , n254783 , n254784 , n254785 , 
     n254786 , n254787 , n254788 , n254789 , n254790 , n254791 , n254792 , n254793 , n254794 , n254795 , 
     n254796 , n254797 , n254798 , n254799 , n254800 , n254801 , n254802 , n254803 , n254804 , n254805 , 
     n254806 , n254807 , n254808 , n254809 , n254810 , n254811 , n254812 , n254813 , n254814 , n254815 , 
     n254816 , n254817 , n254818 , n254819 , n254820 , n254821 , n254822 , n254823 , n254824 , n254825 , 
     n254826 , n254827 , n254828 , n254829 , n254830 , n254831 , n254832 , n254833 , n254834 , n254835 , 
     n254836 , n254837 , n254838 , n254839 , n254840 , n254841 , n254842 , n254843 , n254844 , n254845 , 
     n254846 , n254847 , n254848 , n254849 , n254850 , n254851 , n254852 , n254853 , n254854 , n254855 , 
     n254856 , n254857 , n254858 , n254859 , n254860 , n254861 , n254862 , n254863 , n254864 , n254865 , 
     n254866 , n254867 , n254868 , n254869 , n254870 , n254871 , n254872 , n254873 , n254874 , n254875 , 
     n254876 , n254877 , n254878 , n254879 , n254880 , n254881 , n254882 , n254883 , n254884 , n254885 , 
     n254886 , n254887 , n254888 , n254889 , n254890 , n254891 , n254892 , n254893 , n254894 , n254895 , 
     n254896 , n254897 , n254898 , n254899 , n254900 , n254901 , n254902 , n254903 , n254904 , n254905 , 
     n254906 , n254907 , n254908 , n254909 , n254910 , n254911 , n254912 , n254913 , n254914 , n254915 , 
     n254916 , n254917 , n254918 , n254919 , n254920 , n254921 , n254922 , n254923 , n254924 , n254925 , 
     n254926 , n254927 , n254928 , n254929 , n254930 , n254931 , n254932 , n254933 , n254934 , n254935 , 
     n254936 , n254937 , n254938 , n254939 , n254940 , n254941 , n254942 , n254943 , n254944 , n254945 , 
     n254946 , n254947 , n254948 , n254949 , n254950 , n254951 , n254952 , n254953 , n254954 , n254955 , 
     n254956 , n254957 , n254958 , n254959 , n254960 , n254961 , n254962 , n254963 , n254964 , n254965 , 
     n254966 , n254967 , n254968 , n254969 , n254970 , n254971 , n254972 , n254973 , n254974 , n254975 , 
     n254976 , n254977 , n254978 , n254979 , n254980 , n254981 , n254982 , n254983 , n254984 , n254985 , 
     n254986 , n254987 , n254988 , n254989 , n254990 , n254991 , n254992 , n254993 , n254994 , n254995 , 
     n254996 , n254997 , n254998 , n254999 , n255000 , n255001 , n255002 , n255003 , n255004 , n255005 , 
     n255006 , n255007 , n255008 , n255009 , n255010 , n255011 , n255012 , n255013 , n255014 , n255015 , 
     n255016 , n255017 , n255018 , n255019 , n255020 , n255021 , n255022 , n255023 , n255024 , n255025 , 
     n255026 , n255027 , n255028 , n255029 , n255030 , n255031 , n255032 , n255033 , n255034 , n255035 , 
     n255036 , n255037 , n255038 , n255039 , n255040 , n255041 , n255042 , n255043 , n255044 , n255045 , 
     n255046 , n255047 , n255048 , n255049 , n255050 , n255051 , n255052 , n255053 , n255054 , n255055 , 
     n255056 , n255057 , n255058 , n255059 , n255060 , n255061 , n255062 , n255063 , n255064 , n255065 , 
     n255066 , n255067 , n255068 , n255069 , n255070 , n255071 , n255072 , n255073 , n255074 , n255075 , 
     n255076 , n255077 , n255078 , n255079 , n255080 , n255081 , n255082 , n255083 , n255084 , n255085 , 
     n255086 , n255087 , n255088 , n255089 , n255090 , n255091 , n255092 , n255093 , n255094 , n255095 , 
     n255096 , n255097 , n255098 , n255099 , n255100 , n255101 , n255102 , n255103 , n255104 , n255105 , 
     n255106 , n255107 , n255108 , n255109 , n255110 , n255111 , n255112 , n255113 , n255114 , n255115 , 
     n255116 , n255117 , n255118 , n255119 , n255120 , n255121 , n255122 , n255123 , n255124 , n255125 , 
     n255126 , n255127 , n255128 , n255129 , n255130 , n255131 , n255132 , n255133 , n255134 , n255135 , 
     n255136 , n255137 , n255138 , n255139 , n255140 , n255141 , n255142 , n255143 , n255144 , n255145 , 
     n255146 , n255147 , n255148 , n255149 , n255150 , n255151 , n255152 , n255153 , n255154 , n255155 , 
     n255156 , n255157 , n255158 , n255159 , n255160 , n255161 , n255162 , n255163 , n255164 , n255165 , 
     n255166 , n255167 , n255168 , n255169 , n255170 , n255171 , n255172 , n255173 , n255174 , n255175 , 
     n255176 , n255177 , n255178 , n255179 , n255180 , n255181 , n255182 , n255183 , n255184 , n255185 , 
     n255186 , n255187 , n255188 , n255189 , n255190 , n255191 , n255192 , n255193 , n255194 , n255195 , 
     n255196 , n255197 , n255198 , n255199 , n255200 , n255201 , n255202 , n255203 , n255204 , n255205 , 
     n255206 , n255207 , n255208 , n255209 , n255210 , n255211 , n255212 , n255213 , n255214 , n255215 , 
     n255216 , n255217 , n255218 , n255219 , n255220 , n255221 , n255222 , n255223 , n255224 , n255225 , 
     n255226 , n255227 , n255228 , n255229 , n255230 , n255231 , n255232 , n255233 , n255234 , n255235 , 
     n255236 , n255237 , n255238 , n255239 , n255240 , n255241 , n255242 , n255243 , n255244 , n255245 , 
     n255246 , n255247 , n255248 , n255249 , n255250 , n255251 , n255252 , n255253 , n255254 , n255255 , 
     n255256 , n255257 , n255258 , n255259 , n255260 , n255261 , n255262 , n255263 , n255264 , n255265 , 
     n255266 , n255267 , n255268 , n255269 , n255270 , n255271 , n255272 , n255273 , n255274 , n255275 , 
     n255276 , n255277 , n255278 , n255279 , n255280 , n255281 , n255282 , n255283 , n255284 , n255285 , 
     n255286 , n255287 , n255288 , n255289 , n255290 , n255291 , n255292 , n255293 , n255294 , n255295 , 
     n255296 , n255297 , n255298 , n255299 , n255300 , n255301 , n255302 , n255303 , n255304 , n255305 , 
     n255306 , n255307 , n255308 , n255309 , n255310 , n255311 , n255312 , n255313 , n255314 , n255315 , 
     n255316 , n255317 , n255318 , n255319 , n255320 , n255321 , n255322 , n255323 , n255324 , n255325 , 
     n255326 , n255327 , n255328 , n255329 , n255330 , n255331 , n255332 , n255333 , n255334 , n255335 , 
     n255336 , n255337 , n255338 , n255339 , n255340 , n255341 , n255342 , n255343 , n255344 , n255345 , 
     n255346 , n255347 , n255348 , n255349 , n255350 , n255351 , n255352 , n255353 , n255354 , n255355 , 
     n255356 , n255357 , n255358 , n255359 , n255360 , n255361 , n255362 , n255363 , n255364 , n255365 , 
     n255366 , n255367 , n255368 , n255369 , n255370 , n255371 , n255372 , n255373 , n255374 , n255375 , 
     n255376 , n255377 , n255378 , n255379 , n255380 , n255381 , n255382 , n255383 , n255384 , n255385 , 
     n255386 , n255387 , n255388 , n255389 , n255390 , n255391 , n255392 , n255393 , n255394 , n255395 , 
     n255396 , n255397 , n255398 , n255399 , n255400 , n255401 , n255402 , n255403 , n255404 , n255405 , 
     n255406 , n255407 , n255408 , n255409 , n255410 , n255411 , n255412 , n255413 , n255414 , n255415 , 
     n255416 , n255417 , n255418 , n255419 , n255420 , n255421 , n255422 , n255423 , n255424 , n255425 , 
     n255426 , n255427 , n255428 , n255429 , n255430 , n255431 , n255432 , n255433 , n255434 , n255435 , 
     n255436 , n255437 , n255438 , n255439 , n255440 , n255441 , n255442 , n255443 , n255444 , n255445 , 
     n255446 , n255447 , n255448 , n255449 , n255450 , n255451 , n255452 , n255453 , n255454 , n255455 , 
     n255456 , n255457 , n255458 , n255459 , n255460 , n255461 , n255462 , n255463 , n255464 , n255465 , 
     n255466 , n255467 , n255468 , n255469 , n255470 , n255471 , n255472 , n255473 , n255474 , n255475 , 
     n255476 , n255477 , n255478 , n255479 , n255480 , n255481 , n255482 , n255483 , n255484 , n255485 , 
     n255486 , n255487 , n255488 , n255489 , n255490 , n255491 , n255492 , n255493 , n255494 , n255495 , 
     n255496 , n255497 , n255498 , n255499 , n255500 , n255501 , n255502 , n255503 , n255504 , n255505 , 
     n255506 , n255507 , n255508 , n255509 , n255510 , n255511 , n255512 , n255513 , n255514 , n255515 , 
     n255516 , n255517 , n255518 , n255519 , n255520 , n255521 , n255522 , n255523 , n255524 , n255525 , 
     n255526 , n255527 , n255528 , n255529 , n255530 , n255531 , n255532 , n255533 , n255534 , n255535 , 
     n255536 , n255537 , n255538 , n255539 , n255540 , n255541 , n255542 , n255543 , n255544 , n255545 , 
     n255546 , n255547 , n255548 , n255549 , n255550 , n255551 , n255552 , n255553 , n255554 , n255555 , 
     n255556 , n255557 , n255558 , n255559 , n255560 , n255561 , n255562 , n255563 , n255564 , n255565 , 
     n255566 , n255567 , n255568 , n255569 , n255570 , n255571 , n255572 , n255573 , n255574 , n255575 , 
     n255576 , n255577 , n255578 , n255579 , n255580 , n255581 , n255582 , n255583 , n255584 , n255585 , 
     n255586 , n255587 , n255588 , n255589 , n255590 , n255591 , n255592 , n255593 , n255594 , n255595 , 
     n255596 , n255597 , n255598 , n255599 , n255600 , n255601 , n255602 , n255603 , n255604 , n255605 , 
     n255606 , n255607 , n255608 , n255609 , n255610 , n255611 , n255612 , n255613 , n255614 , n255615 , 
     n255616 , n255617 , n255618 , n255619 , n255620 , n255621 , n255622 , n255623 , n255624 , n255625 , 
     n255626 , n255627 , n255628 , n255629 , n255630 , n255631 , n255632 , n255633 , n255634 , n255635 , 
     n255636 , n255637 , n255638 , n255639 , n255640 , n255641 , n255642 , n255643 , n255644 , n255645 , 
     n255646 , n255647 , n255648 , n255649 , n255650 , n255651 , n255652 , n255653 , n255654 , n255655 , 
     n255656 , n255657 , n255658 , n255659 , n255660 , n255661 , n255662 , n255663 , n255664 , n255665 , 
     n255666 , n255667 , n255668 , n255669 , n255670 , n255671 , n255672 , n255673 , n255674 , n255675 , 
     n255676 , n255677 , n255678 , n255679 , n255680 , n255681 , n255682 , n255683 , n255684 , n255685 , 
     n255686 , n255687 , n255688 , n255689 , n255690 , n255691 , n255692 , n255693 , n255694 , n255695 , 
     n255696 , n255697 , n255698 , n255699 , n255700 , n255701 , n255702 , n255703 , n255704 , n255705 , 
     n255706 , n255707 , n255708 , n255709 , n255710 , n255711 , n255712 , n255713 , n255714 , n255715 , 
     n255716 , n255717 , n255718 , n255719 , n255720 , n255721 , n255722 , n255723 , n255724 , n255725 , 
     n255726 , n255727 , n255728 , n255729 , n255730 , n255731 , n255732 , n255733 , n255734 , n255735 , 
     n255736 , n255737 , n255738 , n255739 , n255740 , n255741 , n255742 , n255743 , n255744 , n255745 , 
     n255746 , n255747 , n255748 , n255749 , n255750 , n255751 , n255752 , n255753 , n255754 , n255755 , 
     n255756 , n255757 , n255758 , n255759 , n255760 , n255761 , n255762 , n255763 , n255764 , n255765 , 
     n255766 , n255767 , n255768 , n255769 , n255770 , n255771 , n255772 , n255773 , n255774 , n255775 , 
     n255776 , n255777 , n255778 , n255779 , n255780 , n255781 , n255782 , n255783 , n255784 , n255785 , 
     n255786 , n255787 , n255788 , n255789 , n255790 , n255791 , n255792 , n255793 , n255794 , n255795 , 
     n255796 , n255797 , n255798 , n255799 , n255800 , n255801 , n255802 , n255803 , n255804 , n255805 , 
     n255806 , n255807 , n255808 , n255809 , n255810 , n255811 , n255812 , n255813 , n255814 , n255815 , 
     n255816 , n255817 , n255818 , n255819 , n255820 , n255821 , n255822 , n255823 , n255824 , n255825 , 
     n255826 , n255827 , n255828 , n255829 , n255830 , n255831 , n255832 , n255833 , n255834 , n255835 , 
     n255836 , n255837 , n255838 , n255839 , n255840 , n255841 , n255842 , n255843 , n255844 , n255845 , 
     n255846 , n255847 , n255848 , n255849 , n255850 , n255851 , n255852 , n255853 , n255854 , n255855 , 
     n255856 , n255857 , n255858 , n255859 , n255860 , n255861 , n255862 , n255863 , n255864 , n255865 , 
     n255866 , n255867 , n255868 , n255869 , n255870 , n255871 , n255872 , n255873 , n255874 , n255875 , 
     n255876 , n255877 , n255878 , n255879 , n255880 , n255881 , n255882 , n255883 , n255884 , n255885 , 
     n255886 , n255887 , n255888 , n255889 , n255890 , n255891 , n255892 , n255893 , n255894 , n255895 , 
     n255896 , n255897 , n255898 , n255899 , n255900 , n255901 , n255902 , n255903 , n255904 , n255905 , 
     n255906 , n255907 , n255908 , n255909 , n255910 , n255911 , n255912 , n255913 , n255914 , n255915 , 
     n255916 , n255917 , n255918 , n255919 , n255920 , n255921 , n255922 , n255923 , n255924 , n255925 , 
     n255926 , n255927 , n255928 , n255929 , n255930 , n255931 , n255932 , n255933 , n255934 , n255935 , 
     n255936 , n255937 , n255938 , n255939 , n255940 , n255941 , n255942 , n255943 , n255944 , n255945 , 
     n255946 , n255947 , n255948 , n255949 , n255950 , n255951 , n255952 , n255953 , n255954 , n255955 , 
     n255956 , n255957 , n255958 , n255959 , n255960 , n255961 , n255962 , n255963 , n255964 , n255965 , 
     n255966 , n255967 , n255968 , n255969 , n255970 , n255971 , n255972 , n255973 , n255974 , n255975 , 
     n255976 , n255977 , n255978 , n255979 , n255980 , n255981 , n255982 , n255983 , n255984 , n255985 , 
     n255986 , n255987 , n255988 , n255989 , n255990 , n255991 , n255992 , n255993 , n255994 , n255995 , 
     n255996 , n255997 , n255998 , n255999 , n256000 , n256001 , n256002 , n256003 , n256004 , n256005 , 
     n256006 , n256007 , n256008 , n256009 , n256010 , n256011 , n256012 , n256013 , n256014 , n256015 , 
     n256016 , n256017 , n256018 , n256019 , n256020 , n256021 , n256022 , n256023 , n256024 , n256025 , 
     n256026 , n256027 , n256028 , n256029 , n256030 , n256031 , n256032 , n256033 , n256034 , n256035 , 
     n256036 , n256037 , n256038 , n256039 , n256040 , n256041 , n256042 , n256043 , n256044 , n256045 , 
     n256046 , n256047 , n256048 , n256049 , n256050 , n256051 , n256052 , n256053 , n256054 , n256055 , 
     n256056 , n256057 , n256058 , n256059 , n256060 , n256061 , n256062 , n256063 , n256064 , n256065 , 
     n256066 , n256067 , n256068 , n256069 , n256070 , n256071 , n256072 , n256073 , n256074 , n256075 , 
     n256076 , n256077 , n256078 , n256079 , n256080 , n256081 , n256082 , n256083 , n256084 , n256085 , 
     n256086 , n256087 , n256088 , n256089 , n256090 , n256091 , n256092 , n256093 , n256094 , n256095 , 
     n256096 , n256097 , n256098 , n256099 , n256100 , n256101 , n256102 , n256103 , n256104 , n256105 , 
     n256106 , n256107 , n256108 , n256109 , n256110 , n256111 , n256112 , n256113 , n256114 , n256115 , 
     n256116 , n256117 , n256118 , n256119 , n256120 , n256121 , n256122 , n256123 , n256124 , n256125 , 
     n256126 , n256127 , n256128 , n256129 , n256130 , n256131 , n256132 , n256133 , n256134 , n256135 , 
     n256136 , n256137 , n256138 , n256139 , n256140 , n256141 , n256142 , n256143 , n256144 , n256145 , 
     n256146 , n256147 , n256148 , n256149 , n256150 , n256151 , n256152 , n256153 , n256154 , n256155 , 
     n256156 , n256157 , n256158 , n256159 , n256160 , n256161 , n256162 , n256163 , n256164 , n256165 , 
     n256166 , n256167 , n256168 , n256169 , n256170 , n256171 , n256172 , n256173 , n256174 , n256175 , 
     n256176 , n256177 , n256178 , n256179 , n256180 , n256181 , n256182 , n256183 , n256184 , n256185 , 
     n256186 , n256187 , n256188 , n256189 , n256190 , n256191 , n256192 , n256193 , n256194 , n256195 , 
     n256196 , n256197 , n256198 , n256199 , n256200 , n256201 , n256202 , n256203 , n256204 , n256205 , 
     n256206 , n256207 , n256208 , n256209 , n256210 , n256211 , n256212 , n256213 , n256214 , n256215 , 
     n256216 , n256217 , n256218 , n256219 , n256220 , n256221 , n256222 , n256223 , n256224 , n256225 , 
     n256226 , n256227 , n256228 , n256229 , n256230 , n256231 , n256232 , n256233 , n256234 , n256235 , 
     n256236 , n256237 , n256238 , n256239 , n256240 , n256241 , n256242 , n256243 , n256244 , n256245 , 
     n256246 , n256247 , n256248 , n256249 , n256250 , n256251 , n256252 , n256253 , n256254 , n256255 , 
     n256256 , n256257 , n256258 , n256259 , n256260 , n256261 , n256262 , n256263 , n256264 , n256265 , 
     n256266 , n256267 , n256268 , n256269 , n256270 , n256271 , n256272 , n256273 , n256274 , n256275 , 
     n256276 , n256277 , n256278 , n256279 , n256280 , n256281 , n256282 , n256283 , n256284 , n256285 , 
     n256286 , n256287 , n256288 , n256289 , n256290 , n256291 , n256292 , n256293 , n256294 , n256295 , 
     n256296 , n256297 , n256298 , n256299 , n256300 , n256301 , n256302 , n256303 , n256304 , n256305 , 
     n256306 , n256307 , n256308 , n256309 , n256310 , n256311 , n256312 , n256313 , n256314 , n256315 , 
     n256316 , n256317 , n256318 , n256319 , n256320 , n256321 , n256322 , n256323 , n256324 , n256325 , 
     n256326 , n256327 , n256328 , n256329 , n256330 , n256331 , n256332 , n256333 , n256334 , n256335 , 
     n256336 , n256337 , n256338 , n256339 , n256340 , n256341 , n256342 , n256343 , n256344 , n256345 , 
     n256346 , n256347 , n256348 , n256349 , n256350 , n256351 , n256352 , n256353 , n256354 , n256355 , 
     n256356 , n256357 , n256358 , n256359 , n256360 , n256361 , n256362 , n256363 , n256364 , n256365 , 
     n256366 , n256367 , n256368 , n256369 , n256370 , n256371 , n256372 , n256373 , n256374 , n256375 , 
     n256376 , n256377 , n256378 , n256379 , n256380 , n256381 , n256382 , n256383 , n256384 , n256385 , 
     n256386 , n256387 , n256388 , n256389 , n256390 , n256391 , n256392 , n256393 , n256394 , n256395 , 
     n256396 , n256397 , n256398 , n256399 , n256400 , n256401 , n256402 , n256403 , n256404 , n256405 , 
     n256406 , n256407 , n256408 , n256409 , n256410 , n256411 , n256412 , n256413 , n256414 , n256415 , 
     n256416 , n256417 , n256418 , n256419 , n256420 , n256421 , n256422 , n256423 , n256424 , n256425 , 
     n256426 , n256427 , n256428 , n256429 , n256430 , n256431 , n256432 , n256433 , n256434 , n256435 , 
     n256436 , n256437 , n256438 , n256439 , n256440 , n256441 , n256442 , n256443 , n256444 , n256445 , 
     n256446 , n256447 , n256448 , n256449 , n256450 , n256451 , n256452 , n256453 , n256454 , n256455 , 
     n256456 , n256457 , n256458 , n256459 , n256460 , n256461 , n256462 , n256463 , n256464 , n256465 , 
     n256466 , n256467 , n256468 , n256469 , n256470 , n256471 , n256472 , n256473 , n256474 , n256475 , 
     n256476 , n256477 , n256478 , n256479 , n256480 , n256481 , n256482 , n256483 , n256484 , n256485 , 
     n256486 , n256487 , n256488 , n256489 , n256490 , n256491 , n256492 , n256493 , n256494 , n256495 , 
     n256496 , n256497 , n256498 , n256499 , n256500 , n256501 , n256502 , n256503 , n256504 , n256505 , 
     n256506 , n256507 , n256508 , n256509 , n256510 , n256511 , n256512 , n256513 , n256514 , n256515 , 
     n256516 , n256517 , n256518 , n256519 , n256520 , n256521 , n256522 , n256523 , n256524 , n256525 , 
     n256526 , n256527 , n256528 , n256529 , n256530 , n256531 , n256532 , n256533 , n256534 , n256535 , 
     n256536 , n256537 , n256538 , n256539 , n256540 , n256541 , n256542 , n256543 , n256544 , n256545 , 
     n256546 , n256547 , n256548 , n256549 , n256550 , n256551 , n256552 , n256553 , n256554 , n256555 , 
     n256556 , n256557 , n256558 , n256559 , n256560 , n256561 , n256562 , n256563 , n256564 , n256565 , 
     n256566 , n256567 , n256568 , n256569 , n256570 , n256571 , n256572 , n256573 , n256574 , n256575 , 
     n256576 , n256577 , n256578 , n256579 , n256580 , n256581 , n256582 , n256583 , n256584 , n256585 , 
     n256586 , n256587 , n256588 , n256589 , n256590 , n256591 , n256592 , n256593 , n256594 , n256595 , 
     n256596 , n256597 , n256598 , n256599 , n256600 , n256601 , n256602 , n256603 , n256604 , n256605 , 
     n256606 , n256607 , n256608 , n256609 , n256610 , n256611 , n256612 , n256613 , n256614 , n256615 , 
     n256616 , n256617 , n256618 , n256619 , n256620 , n256621 , n256622 , n256623 , n256624 , n256625 , 
     n256626 , n256627 , n256628 , n256629 , n256630 , n256631 , n256632 , n256633 , n256634 , n256635 , 
     n256636 , n256637 , n256638 , n256639 , n256640 , n256641 , n256642 , n256643 , n256644 , n256645 , 
     n256646 , n256647 , n256648 , n256649 , n256650 , n256651 , n256652 , n256653 , n256654 , n256655 , 
     n256656 , n256657 , n256658 , n256659 , n256660 , n256661 , n256662 , n256663 , n256664 , n256665 , 
     n256666 , n256667 , n256668 , n256669 , n256670 , n256671 , n256672 , n256673 , n256674 , n256675 , 
     n256676 , n256677 , n256678 , n256679 , n256680 , n256681 , n256682 , n256683 , n256684 , n256685 , 
     n256686 , n256687 , n256688 , n256689 , n256690 , n256691 , n256692 , n256693 , n256694 , n256695 , 
     n256696 , n256697 , n256698 , n256699 , n256700 , n256701 , n256702 , n256703 , n256704 , n256705 , 
     n256706 , n256707 , n256708 , n256709 , n256710 , n256711 , n256712 , n256713 , n256714 , n256715 , 
     n256716 , n256717 , n256718 , n256719 , n256720 , n256721 , n256722 , n256723 , n256724 , n256725 , 
     n256726 , n256727 , n256728 , n256729 , n256730 , n256731 , n256732 , n256733 , n256734 , n256735 , 
     n256736 , n256737 , n256738 , n256739 , n256740 , n256741 , n256742 , n256743 , n256744 , n256745 , 
     n256746 , n256747 , n256748 , n256749 , n256750 , n256751 , n256752 , n256753 , n256754 , n256755 , 
     n256756 , n256757 , n256758 , n256759 , n256760 , n256761 , n256762 , n256763 , n256764 , n256765 , 
     n256766 , n256767 , n256768 , n256769 , n256770 , n256771 , n256772 , n256773 , n256774 , n256775 , 
     n256776 , n256777 , n256778 , n256779 , n256780 , n256781 , n256782 , n256783 , n256784 , n256785 , 
     n256786 , n256787 , n256788 , n256789 , n256790 , n256791 , n256792 , n256793 , n256794 , n256795 , 
     n256796 , n256797 , n256798 , n256799 , n256800 , n256801 , n256802 , n256803 , n256804 , n256805 , 
     n256806 , n256807 , n256808 , n256809 , n256810 , n256811 , n256812 , n256813 , n256814 , n256815 , 
     n256816 , n256817 , n256818 , n256819 , n256820 , n256821 , n256822 , n256823 , n256824 , n256825 , 
     n256826 , n256827 , n256828 , n256829 , n256830 , n256831 , n256832 , n256833 , n256834 , n256835 , 
     n256836 , n256837 , n256838 , n256839 , n256840 , n256841 , n256842 , n256843 , n256844 , n256845 , 
     n256846 , n256847 , n256848 , n256849 , n256850 , n256851 , n256852 , n256853 , n256854 , n256855 , 
     n256856 , n256857 , n256858 , n256859 , n256860 , n256861 , n256862 , n256863 , n256864 , n256865 , 
     n256866 , n256867 , n256868 , n256869 , n256870 , n256871 , n256872 , n256873 , n256874 , n256875 , 
     n256876 , n256877 , n256878 , n256879 , n256880 , n256881 , n256882 , n256883 , n256884 , n256885 , 
     n256886 , n256887 , n256888 , n256889 , n256890 , n256891 , n256892 , n256893 , n256894 , n256895 , 
     n256896 , n256897 , n256898 , n256899 , n256900 , n256901 , n256902 , n256903 , n256904 , n256905 , 
     n256906 , n256907 , n256908 , n256909 , n256910 , n256911 , n256912 , n256913 , n256914 , n256915 , 
     n256916 , n256917 , n256918 , n256919 , n256920 , n256921 , n256922 , n256923 , n256924 , n256925 , 
     n256926 , n256927 , n256928 , n256929 , n256930 , n256931 , n256932 , n256933 , n256934 , n256935 , 
     n256936 , n256937 , n256938 , n256939 , n256940 , n256941 , n256942 , n256943 , n256944 , n256945 , 
     n256946 , n256947 , n256948 , n256949 , n256950 , n256951 , n256952 , n256953 , n256954 , n256955 , 
     n256956 , n256957 , n256958 , n256959 , n256960 , n256961 , n256962 , n256963 , n256964 , n256965 , 
     n256966 , n256967 , n256968 , n256969 , n256970 , n256971 , n256972 , n256973 , n256974 , n256975 , 
     n256976 , n256977 , n256978 , n256979 , n256980 , n256981 , n256982 , n256983 , n256984 , n256985 , 
     n256986 , n256987 , n256988 , n256989 , n256990 , n256991 , n256992 , n256993 , n256994 , n256995 , 
     n256996 , n256997 , n256998 , n256999 , n257000 , n257001 , n257002 , n257003 , n257004 , n257005 , 
     n257006 , n257007 , n257008 , n257009 , n257010 , n257011 , n257012 , n257013 , n257014 , n257015 , 
     n257016 , n257017 , n257018 , n257019 , n257020 , n257021 , n257022 , n257023 , n257024 , n257025 , 
     n257026 , n257027 , n257028 , n257029 , n257030 , n257031 , n257032 , n257033 , n257034 , n257035 , 
     n257036 , n257037 , n257038 , n257039 , n257040 , n257041 , n257042 , n257043 , n257044 , n257045 , 
     n257046 , n257047 , n257048 , n257049 , n257050 , n257051 , n257052 , n257053 , n257054 , n257055 , 
     n257056 , n257057 , n257058 , n257059 , n257060 , n257061 , n257062 , n257063 , n257064 , n257065 , 
     n257066 , n257067 , n257068 , n257069 , n257070 , n257071 , n257072 , n257073 , n257074 , n257075 , 
     n257076 , n257077 , n257078 , n257079 , n257080 , n257081 , n257082 , n257083 , n257084 , n257085 , 
     n257086 , n257087 , n257088 , n257089 , n257090 , n257091 , n257092 , n257093 , n257094 , n257095 , 
     n257096 , n257097 , n257098 , n257099 , n257100 , n257101 , n257102 , n257103 , n257104 , n257105 , 
     n257106 , n257107 , n257108 , n257109 , n257110 , n257111 , n257112 , n257113 , n257114 , n257115 , 
     n257116 , n257117 , n257118 , n257119 , n257120 , n257121 , n257122 , n257123 , n257124 , n257125 , 
     n257126 , n257127 , n257128 , n257129 , n257130 , n257131 , n257132 , n257133 , n257134 , n257135 , 
     n257136 , n257137 , n257138 , n257139 , n257140 , n257141 , n257142 , n257143 , n257144 , n257145 , 
     n257146 , n257147 , n257148 , n257149 , n257150 , n257151 , n257152 , n257153 , n257154 , n257155 , 
     n257156 , n257157 , n257158 , n257159 , n257160 , n257161 , n257162 , n257163 , n257164 , n257165 , 
     n257166 , n257167 , n257168 , n257169 , n257170 , n257171 , n257172 , n257173 , n257174 , n257175 , 
     n257176 , n257177 , n257178 , n257179 , n257180 , n257181 , n257182 , n257183 , n257184 , n257185 , 
     n257186 , n257187 , n257188 , n257189 , n257190 , n257191 , n257192 , n257193 , n257194 , n257195 , 
     n257196 , n257197 , n257198 , n257199 , n257200 , n257201 , n257202 , n257203 , n257204 , n257205 , 
     n257206 , n257207 , n257208 , n257209 , n257210 , n257211 , n257212 , n257213 , n257214 , n257215 , 
     n257216 , n257217 , n257218 , n257219 , n257220 , n257221 , n257222 , n257223 , n257224 , n257225 , 
     n257226 , n257227 , n257228 , n257229 , n257230 , n257231 , n257232 , n257233 , n257234 , n257235 , 
     n257236 , n257237 , n257238 , n257239 , n257240 , n257241 , n257242 , n257243 , n257244 , n257245 , 
     n257246 , n257247 , n257248 , n257249 , n257250 , n257251 , n257252 , n257253 , n257254 , n257255 , 
     n257256 , n257257 , n257258 , n257259 , n257260 , n257261 , n257262 , n257263 , n257264 , n257265 , 
     n257266 , n257267 , n257268 , n257269 , n257270 , n257271 , n257272 , n257273 , n257274 , n257275 , 
     n257276 , n257277 , n257278 , n257279 , n257280 , n257281 , n257282 , n257283 , n257284 , n257285 , 
     n257286 , n257287 , n257288 , n257289 , n257290 , n257291 , n257292 , n257293 , n257294 , n257295 , 
     n257296 , n257297 , n257298 , n257299 , n257300 , n257301 , n257302 , n257303 , n257304 , n257305 , 
     n257306 , n257307 , n257308 , n257309 , n257310 , n257311 , n257312 , n257313 , n257314 , n257315 , 
     n257316 , n257317 , n257318 , n257319 , n257320 , n257321 , n257322 , n257323 , n257324 , n257325 , 
     n257326 , n257327 , n257328 , n257329 , n257330 , n257331 , n257332 , n257333 , n257334 , n257335 , 
     n257336 , n257337 , n257338 , n257339 , n257340 , n257341 , n257342 , n257343 , n257344 , n257345 , 
     n257346 , n257347 , n257348 , n257349 , n257350 , n257351 , n257352 , n257353 , n257354 , n257355 , 
     n257356 , n257357 , n257358 , n257359 , n257360 , n257361 , n257362 , n257363 , n257364 , n257365 , 
     n257366 , n257367 , n257368 , n257369 , n257370 , n257371 , n257372 , n257373 , n257374 , n257375 , 
     n257376 , n257377 , n257378 , n257379 , n257380 , n257381 , n257382 , n257383 , n257384 , n257385 , 
     n257386 , n257387 , n257388 , n257389 , n257390 , n257391 , n257392 , n257393 , n257394 , n257395 , 
     n257396 , n257397 , n257398 , n257399 , n257400 , n257401 , n257402 , n257403 , n257404 , n257405 , 
     n257406 , n257407 , n257408 , n257409 , n257410 , n257411 , n257412 , n257413 , n257414 , n257415 , 
     n257416 , n257417 , n257418 , n257419 , n257420 , n257421 , n257422 , n257423 , n257424 , n257425 , 
     n257426 , n257427 , n257428 , n257429 , n257430 , n257431 , n257432 , n257433 , n257434 , n257435 , 
     n257436 , n257437 , n257438 , n257439 , n257440 , n257441 , n257442 , n257443 , n257444 , n257445 , 
     n257446 , n257447 , n257448 , n257449 , n257450 , n257451 , n257452 , n257453 , n257454 , n257455 , 
     n257456 , n257457 , n257458 , n257459 , n257460 , n257461 , n257462 , n257463 , n257464 , n257465 , 
     n257466 , n257467 , n257468 , n257469 , n257470 , n257471 , n257472 , n257473 , n257474 , n257475 , 
     n257476 , n257477 , n257478 , n257479 , n257480 , n257481 , n257482 , n257483 , n257484 , n257485 , 
     n257486 , n257487 , n257488 , n257489 , n257490 , n257491 , n257492 , n257493 , n257494 , n257495 , 
     n257496 , n257497 , n257498 , n257499 , n257500 , n257501 , n257502 , n257503 , n257504 , n257505 , 
     n257506 , n257507 , n257508 , n257509 , n257510 , n257511 , n257512 , n257513 , n257514 , n257515 , 
     n257516 , n257517 , n257518 , n257519 , n257520 , n257521 , n257522 , n257523 , n257524 , n257525 , 
     n257526 , n257527 , n257528 , n257529 , n257530 , n257531 , n257532 , n257533 , n257534 , n257535 , 
     n257536 , n257537 , n257538 , n257539 , n257540 , n257541 , n257542 , n257543 , n257544 , n257545 , 
     n257546 , n257547 , n257548 , n257549 , n257550 , n257551 , n257552 , n257553 , n257554 , n257555 , 
     n257556 , n257557 , n257558 , n257559 , n257560 , n257561 , n257562 , n257563 , n257564 , n257565 , 
     n257566 , n257567 , n257568 , n257569 , n257570 , n257571 , n257572 , n257573 , n257574 , n257575 , 
     n257576 , n257577 , n257578 , n257579 , n257580 , n257581 , n257582 , n257583 , n257584 , n257585 , 
     n257586 , n257587 , n257588 , n257589 , n257590 , n257591 , n257592 , n257593 , n257594 , n257595 , 
     n257596 , n257597 , n257598 , n257599 , n257600 , n257601 , n257602 , n257603 , n257604 , n257605 , 
     n257606 , n257607 , n257608 , n257609 , n257610 , n257611 , n257612 , n257613 , n257614 , n257615 , 
     n257616 , n257617 , n257618 , n257619 , n257620 , n257621 , n257622 , n257623 , n257624 , n257625 , 
     n257626 , n257627 , n257628 , n257629 , n257630 , n257631 , n257632 , n257633 , n257634 , n257635 , 
     n257636 , n257637 , n257638 , n257639 , n257640 , n257641 , n257642 , n257643 , n257644 , n257645 , 
     n257646 , n257647 , n257648 , n257649 , n257650 , n257651 , n257652 , n257653 , n257654 , n257655 , 
     n257656 , n257657 , n257658 , n257659 , n257660 , n257661 , n257662 , n257663 , n257664 , n257665 , 
     n257666 , n257667 , n257668 , n257669 , n257670 , n257671 , n257672 , n257673 , n257674 , n257675 , 
     n257676 , n257677 , n257678 , n257679 , n257680 , n257681 , n257682 , n257683 , n257684 , n257685 , 
     n257686 , n257687 , n257688 , n257689 , n257690 , n257691 , n257692 , n257693 , n257694 , n257695 , 
     n257696 , n257697 , n257698 , n257699 , n257700 , n257701 , n257702 , n257703 , n257704 , n257705 , 
     n257706 , n257707 , n257708 , n257709 , n257710 , n257711 , n257712 , n257713 , n257714 , n257715 , 
     n257716 , n257717 , n257718 , n257719 , n257720 , n257721 , n257722 , n257723 , n257724 , n257725 , 
     n257726 , n257727 , n257728 , n257729 , n257730 , n257731 , n257732 , n257733 , n257734 , n257735 , 
     n257736 , n257737 , n257738 , n257739 , n257740 , n257741 , n257742 , n257743 , n257744 , n257745 , 
     n257746 , n257747 , n257748 , n257749 , n257750 , n257751 , n257752 , n257753 , n257754 , n257755 , 
     n257756 , n257757 , n257758 , n257759 , n257760 , n257761 , n257762 , n257763 , n257764 , n257765 , 
     n257766 , n257767 , n257768 , n257769 , n257770 , n257771 , n257772 , n257773 , n257774 , n257775 , 
     n257776 , n257777 , n257778 , n257779 , n257780 , n257781 , n257782 , n257783 , n257784 , n257785 , 
     n257786 , n257787 , n257788 , n257789 , n257790 , n257791 , n257792 , n257793 , n257794 , n257795 , 
     n257796 , n257797 , n257798 , n257799 , n257800 , n257801 , n257802 , n257803 , n257804 , n257805 , 
     n257806 , n257807 , n257808 , n257809 , n257810 , n257811 , n257812 , n257813 , n257814 , n257815 , 
     n257816 , n257817 , n257818 , n257819 , n257820 , n257821 , n257822 , n257823 , n257824 , n257825 , 
     n257826 , n257827 , n257828 , n257829 , n257830 , n257831 , n257832 , n257833 , n257834 , n257835 , 
     n257836 , n257837 , n257838 , n257839 , n257840 , n257841 , n257842 , n257843 , n257844 , n257845 , 
     n257846 , n257847 , n257848 , n257849 , n257850 , n257851 , n257852 , n257853 , n257854 , n257855 , 
     n257856 , n257857 , n257858 , n257859 , n257860 , n257861 , n257862 , n257863 , n257864 , n257865 , 
     n257866 , n257867 , n257868 , n257869 , n257870 , n257871 , n257872 , n257873 , n257874 , n257875 , 
     n257876 , n257877 , n257878 , n257879 , n257880 , n257881 , n257882 , n257883 , n257884 , n257885 , 
     n257886 , n257887 , n257888 , n257889 , n257890 , n257891 , n257892 , n257893 , n257894 , n257895 , 
     n257896 , n257897 , n257898 , n257899 , n257900 , n257901 , n257902 , n257903 , n257904 , n257905 , 
     n257906 , n257907 , n257908 , n257909 , n257910 , n257911 , n257912 , n257913 , n257914 , n257915 , 
     n257916 , n257917 , n257918 , n257919 , n257920 , n257921 , n257922 , n257923 , n257924 , n257925 , 
     n257926 , n257927 , n257928 , n257929 , n257930 , n257931 , n257932 , n257933 , n257934 , n257935 , 
     n257936 , n257937 , n257938 , n257939 , n257940 , n257941 , n257942 , n257943 , n257944 , n257945 , 
     n257946 , n257947 , n257948 , n257949 , n257950 , n257951 , n257952 , n257953 , n257954 , n257955 , 
     n257956 , n257957 , n257958 , n257959 , n257960 , n257961 , n257962 , n257963 , n257964 , n257965 , 
     n257966 , n257967 , n257968 , n257969 , n257970 , n257971 , n257972 , n257973 , n257974 , n257975 , 
     n257976 , n257977 , n257978 , n257979 , n257980 , n257981 , n257982 , n257983 , n257984 , n257985 , 
     n257986 , n257987 , n257988 , n257989 , n257990 , n257991 , n257992 , n257993 , n257994 , n257995 , 
     n257996 , n257997 , n257998 , n257999 , n258000 , n258001 , n258002 , n258003 , n258004 , n258005 , 
     n258006 , n258007 , n258008 , n258009 , n258010 , n258011 , n258012 , n258013 , n258014 , n258015 , 
     n258016 , n258017 , n258018 , n258019 , n258020 , n258021 , n258022 , n258023 , n258024 , n258025 , 
     n258026 , n258027 , n258028 , n258029 , n258030 , n258031 , n258032 , n258033 , n258034 , n258035 , 
     n258036 , n258037 , n258038 , n258039 , n258040 , n258041 , n258042 , n258043 , n258044 , n258045 , 
     n258046 , n258047 , n258048 , n258049 , n258050 , n258051 , n258052 , n258053 , n258054 , n258055 , 
     n258056 , n258057 , n258058 , n258059 , n258060 , n258061 , n258062 , n258063 , n258064 , n258065 , 
     n258066 , n258067 , n258068 , n258069 , n258070 , n258071 , n258072 , n258073 , n258074 , n258075 , 
     n258076 , n258077 , n258078 , n258079 , n258080 , n258081 , n258082 , n258083 , n258084 , n258085 , 
     n258086 , n258087 , n258088 , n258089 , n258090 , n258091 , n258092 , n258093 , n258094 , n258095 , 
     n258096 , n258097 , n258098 , n258099 , n258100 , n258101 , n258102 , n258103 , n258104 , n258105 , 
     n258106 , n258107 , n258108 , n258109 , n258110 , n258111 , n258112 , n258113 , n258114 , n258115 , 
     n258116 , n258117 , n258118 , n258119 , n258120 , n258121 , n258122 , n258123 , n258124 , n258125 , 
     n258126 , n258127 , n258128 , n258129 , n258130 , n258131 , n258132 , n258133 , n258134 , n258135 , 
     n258136 , n258137 , n258138 , n258139 , n258140 , n258141 , n258142 , n258143 , n258144 , n258145 , 
     n258146 , n258147 , n258148 , n258149 , n258150 , n258151 , n258152 , n258153 , n258154 , n258155 , 
     n258156 , n258157 , n258158 , n258159 , n258160 , n258161 , n258162 , n258163 , n258164 , n258165 , 
     n258166 , n258167 , n258168 , n258169 , n258170 , n258171 , n258172 , n258173 , n258174 , n258175 , 
     n258176 , n258177 , n258178 , n258179 , n258180 , n258181 , n258182 , n258183 , n258184 , n258185 , 
     n258186 , n258187 , n258188 , n258189 , n258190 , n258191 , n258192 , n258193 , n258194 , n258195 , 
     n258196 , n258197 , n258198 , n258199 , n258200 , n258201 , n258202 , n258203 , n258204 , n258205 , 
     n258206 , n258207 , n258208 , n258209 , n258210 , n258211 , n258212 , n258213 , n258214 , n258215 , 
     n258216 , n258217 , n258218 , n258219 , n258220 , n258221 , n258222 , n258223 , n258224 , n258225 , 
     n258226 , n258227 , n258228 , n258229 , n258230 , n258231 , n258232 , n258233 , n258234 , n258235 , 
     n258236 , n258237 , n258238 , n258239 , n258240 , n258241 , n258242 , n258243 , n258244 , n258245 , 
     n258246 , n258247 , n258248 , n258249 , n258250 , n258251 , n258252 , n258253 , n258254 , n258255 , 
     n258256 , n258257 , n258258 , n258259 , n258260 , n258261 , n258262 , n258263 , n258264 , n258265 , 
     n258266 , n258267 , n258268 , n258269 , n258270 , n258271 , n258272 , n258273 , n258274 , n258275 , 
     n258276 , n258277 , n258278 , n258279 , n258280 , n258281 , n258282 , n258283 , n258284 , n258285 , 
     n258286 , n258287 , n258288 , n258289 , n258290 , n258291 , n258292 , n258293 , n258294 , n258295 , 
     n258296 , n258297 , n258298 , n258299 , n258300 , n258301 , n258302 , n258303 , n258304 , n258305 , 
     n258306 , n258307 , n258308 , n258309 , n258310 , n258311 , n258312 , n258313 , n258314 , n258315 , 
     n258316 , n258317 , n258318 , n258319 , n258320 , n258321 , n258322 , n258323 , n258324 , n258325 , 
     n258326 , n258327 , n258328 , n258329 , n258330 , n258331 , n258332 , n258333 , n258334 , n258335 , 
     n258336 , n258337 , n258338 , n258339 , n258340 , n258341 , n258342 , n258343 , n258344 , n258345 , 
     n258346 , n258347 , n258348 , n258349 , n258350 , n258351 , n258352 , n258353 , n258354 , n258355 , 
     n258356 , n258357 , n258358 , n258359 , n258360 , n258361 , n258362 , n258363 , n258364 , n258365 , 
     n258366 , n258367 , n258368 , n258369 , n258370 , n258371 , n258372 , n258373 , n258374 , n258375 , 
     n258376 , n258377 , n258378 , n258379 , n258380 , n258381 , n258382 , n258383 , n258384 , n258385 , 
     n258386 , n258387 , n258388 , n258389 , n258390 , n258391 , n258392 , n258393 , n258394 , n258395 , 
     n258396 , n258397 , n258398 , n258399 , n258400 , n258401 , n258402 , n258403 , n258404 , n258405 , 
     n258406 , n258407 , n258408 , n258409 , n258410 , n258411 , n258412 , n258413 , n258414 , n258415 , 
     n258416 , n258417 , n258418 , n258419 , n258420 , n258421 , n258422 , n258423 , n258424 , n258425 , 
     n258426 , n258427 , n258428 , n258429 , n258430 , n258431 , n258432 , n258433 , n258434 , n258435 , 
     n258436 , n258437 , n258438 , n258439 , n258440 , n258441 , n258442 , n258443 , n258444 , n258445 , 
     n258446 , n258447 , n258448 , n258449 , n258450 , n258451 , n258452 , n258453 , n258454 , n258455 , 
     n258456 , n258457 , n258458 , n258459 , n258460 , n258461 , n258462 , n258463 , n258464 , n258465 , 
     n258466 , n258467 , n258468 , n258469 , n258470 , n258471 , n258472 , n258473 , n258474 , n258475 , 
     n258476 , n258477 , n258478 , n258479 , n258480 , n258481 , n258482 , n258483 , n258484 , n258485 , 
     n258486 , n258487 , n258488 , n258489 , n258490 , n258491 , n258492 , n258493 , n258494 , n258495 , 
     n258496 , n258497 , n258498 , n258499 , n258500 , n258501 , n258502 , n258503 , n258504 , n258505 , 
     n258506 , n258507 , n258508 , n258509 , n258510 , n258511 , n258512 , n258513 , n258514 , n258515 , 
     n258516 , n258517 , n258518 , n258519 , n258520 , n258521 , n258522 , n258523 , n258524 , n258525 , 
     n258526 , n258527 , n258528 , n258529 , n258530 , n258531 , n258532 , n258533 , n258534 , n258535 , 
     n258536 , n258537 , n258538 , n258539 , n258540 , n258541 , n258542 , n258543 , n258544 , n258545 , 
     n258546 , n258547 , n258548 , n258549 , n258550 , n258551 , n258552 , n258553 , n258554 , n258555 , 
     n258556 , n258557 , n258558 , n258559 , n258560 , n258561 , n258562 , n258563 , n258564 , n258565 , 
     n258566 , n258567 , n258568 , n258569 , n258570 , n258571 , n258572 , n258573 , n258574 , n258575 , 
     n258576 , n258577 , n258578 , n258579 , n258580 , n258581 , n258582 , n258583 , n258584 , n258585 , 
     n258586 , n258587 , n258588 , n258589 , n258590 , n258591 , n258592 , n258593 , n258594 , n258595 , 
     n258596 , n258597 , n258598 , n258599 , n258600 , n258601 , n258602 , n258603 , n258604 , n258605 , 
     n258606 , n258607 , n258608 , n258609 , n258610 , n258611 , n258612 , n258613 , n258614 , n258615 , 
     n258616 , n258617 , n258618 , n258619 , n258620 , n258621 , n258622 , n258623 , n258624 , n258625 , 
     n258626 , n258627 , n258628 , n258629 , n258630 , n258631 , n258632 , n258633 , n258634 , n258635 , 
     n258636 , n258637 , n258638 , n258639 , n258640 , n258641 , n258642 , n258643 , n258644 , n258645 , 
     n258646 , n258647 , n258648 , n258649 , n258650 , n258651 , n258652 , n258653 , n258654 , n258655 , 
     n258656 , n258657 , n258658 , n258659 , n258660 , n258661 , n258662 , n258663 , n258664 , n258665 , 
     n258666 , n258667 , n258668 , n258669 , n258670 , n258671 , n258672 , n258673 , n258674 , n258675 , 
     n258676 , n258677 , n258678 , n258679 , n258680 , n258681 , n258682 , n258683 , n258684 , n258685 , 
     n258686 , n258687 , n258688 , n258689 , n258690 , n258691 , n258692 , n258693 , n258694 , n258695 , 
     n258696 , n258697 , n258698 , n258699 , n258700 , n258701 , n258702 , n258703 , n258704 , n258705 , 
     n258706 , n258707 , n258708 , n258709 , n258710 , n258711 , n258712 , n258713 , n258714 , n258715 , 
     n258716 , n258717 , n258718 , n258719 , n258720 , n258721 , n258722 , n258723 , n258724 , n258725 , 
     n258726 , n258727 , n258728 , n258729 , n258730 , n258731 , n258732 , n258733 , n258734 , n258735 , 
     n258736 , n258737 , n258738 , n258739 , n258740 , n258741 , n258742 , n258743 , n258744 , n258745 , 
     n258746 , n258747 , n258748 , n258749 , n258750 , n258751 , n258752 , n258753 , n258754 , n258755 , 
     n258756 , n258757 , n258758 , n258759 , n258760 , n258761 , n258762 , n258763 , n258764 , n258765 , 
     n258766 , n258767 , n258768 , n258769 , n258770 , n258771 , n258772 , n258773 , n258774 , n258775 , 
     n258776 , n258777 , n258778 , n258779 , n258780 , n258781 , n258782 , n258783 , n258784 , n258785 , 
     n258786 , n258787 , n258788 , n258789 , n258790 , n258791 , n258792 , n258793 , n258794 , n258795 , 
     n258796 , n258797 , n258798 , n258799 , n258800 , n258801 , n258802 , n258803 , n258804 , n258805 , 
     n258806 , n258807 , n258808 , n258809 , n258810 , n258811 , n258812 , n258813 , n258814 , n258815 , 
     n258816 , n258817 , n258818 , n258819 , n258820 , n258821 , n258822 , n258823 , n258824 , n258825 , 
     n258826 , n258827 , n258828 , n258829 , n258830 , n258831 , n258832 , n258833 , n258834 , n258835 , 
     n258836 , n258837 , n258838 , n258839 , n258840 , n258841 , n258842 , n258843 , n258844 , n258845 , 
     n258846 , n258847 , n258848 , n258849 , n258850 , n258851 , n258852 , n258853 , n258854 , n258855 , 
     n258856 , n258857 , n258858 , n258859 , n258860 , n258861 , n258862 , n258863 , n258864 , n258865 , 
     n258866 , n258867 , n258868 , n258869 , n258870 , n258871 , n258872 , n258873 , n258874 , n258875 , 
     n258876 , n258877 , n258878 , n258879 , n258880 , n258881 , n258882 , n258883 , n258884 , n258885 , 
     n258886 , n258887 , n258888 , n258889 , n258890 , n258891 , n258892 , n258893 , n258894 , n258895 , 
     n258896 , n258897 , n258898 , n258899 , n258900 , n258901 , n258902 , n258903 , n258904 , n258905 , 
     n258906 , n258907 , n258908 , n258909 , n258910 , n258911 , n258912 , n258913 , n258914 , n258915 , 
     n258916 , n258917 , n258918 , n258919 , n258920 , n258921 , n258922 , n258923 , n258924 , n258925 , 
     n258926 , n258927 , n258928 , n258929 , n258930 , n258931 , n258932 , n258933 , n258934 , n258935 , 
     n258936 , n258937 , n258938 , n258939 , n258940 , n258941 , n258942 , n258943 , n258944 , n258945 , 
     n258946 , n258947 , n258948 , n258949 , n258950 , n258951 , n258952 , n258953 , n258954 , n258955 , 
     n258956 , n258957 , n258958 , n258959 , n258960 , n258961 , n258962 , n258963 , n258964 , n258965 , 
     n258966 , n258967 , n258968 , n258969 , n258970 , n258971 , n258972 , n258973 , n258974 , n258975 , 
     n258976 , n258977 , n258978 , n258979 , n258980 , n258981 , n258982 , n258983 , n258984 , n258985 , 
     n258986 , n258987 , n258988 , n258989 , n258990 , n258991 , n258992 , n258993 , n258994 , n258995 , 
     n258996 , n258997 , n258998 , n258999 , n259000 , n259001 , n259002 , n259003 , n259004 , n259005 , 
     n259006 , n259007 , n259008 , n259009 , n259010 , n259011 , n259012 , n259013 , n259014 , n259015 , 
     n259016 , n259017 , n259018 , n259019 , n259020 , n259021 , n259022 , n259023 , n259024 , n259025 , 
     n259026 , n259027 , n259028 , n259029 , n259030 , n259031 , n259032 , n259033 , n259034 , n259035 , 
     n259036 , n259037 , n259038 , n259039 , n259040 , n259041 , n259042 , n259043 , n259044 , n259045 , 
     n259046 , n259047 , n259048 , n259049 , n259050 , n259051 , n259052 , n259053 , n259054 , n259055 , 
     n259056 , n259057 , n259058 , n259059 , n259060 , n259061 , n259062 , n259063 , n259064 , n259065 , 
     n259066 , n259067 , n259068 , n259069 , n259070 , n259071 , n259072 , n259073 , n259074 , n259075 , 
     n259076 , n259077 , n259078 , n259079 , n259080 , n259081 , n259082 , n259083 , n259084 , n259085 , 
     n259086 , n259087 , n259088 , n259089 , n259090 , n259091 , n259092 , n259093 , n259094 , n259095 , 
     n259096 , n259097 , n259098 , n259099 , n259100 , n259101 , n259102 , n259103 , n259104 , n259105 , 
     n259106 , n259107 , n259108 , n259109 , n259110 , n259111 , n259112 , n259113 , n259114 , n259115 , 
     n259116 , n259117 , n259118 , n259119 , n259120 , n259121 , n259122 , n259123 , n259124 , n259125 , 
     n259126 , n259127 , n259128 , n259129 , n259130 , n259131 , n259132 , n259133 , n259134 , n259135 , 
     n259136 , n259137 , n259138 , n259139 , n259140 , n259141 , n259142 , n259143 , n259144 , n259145 , 
     n259146 , n259147 , n259148 , n259149 , n259150 , n259151 , n259152 , n259153 , n259154 , n259155 , 
     n259156 , n259157 , n259158 , n259159 , n259160 , n259161 , n259162 , n259163 , n259164 , n259165 , 
     n259166 , n259167 , n259168 , n259169 , n259170 , n259171 , n259172 , n259173 , n259174 , n259175 , 
     n259176 , n259177 , n259178 , n259179 , n259180 , n259181 , n259182 , n259183 , n259184 , n259185 , 
     n259186 , n259187 , n259188 , n259189 , n259190 , n259191 , n259192 , n259193 , n259194 , n259195 , 
     n259196 , n259197 , n259198 , n259199 , n259200 , n259201 , n259202 , n259203 , n259204 , n259205 , 
     n259206 , n259207 , n259208 , n259209 , n259210 , n259211 , n259212 , n259213 , n259214 , n259215 , 
     n259216 , n259217 , n259218 , n259219 , n259220 , n259221 , n259222 , n259223 , n259224 , n259225 , 
     n259226 , n259227 , n259228 , n259229 , n259230 , n259231 , n259232 , n259233 , n259234 , n259235 , 
     n259236 , n259237 , n259238 , n259239 , n259240 , n259241 , n259242 , n259243 , n259244 , n259245 , 
     n259246 , n259247 , n259248 , n259249 , n259250 , n259251 , n259252 , n259253 , n259254 , n259255 , 
     n259256 , n259257 , n259258 , n259259 , n259260 , n259261 , n259262 , n259263 , n259264 , n259265 , 
     n259266 , n259267 , n259268 , n259269 , n259270 , n259271 , n259272 , n259273 , n259274 , n259275 , 
     n259276 , n259277 , n259278 , n259279 , n259280 , n259281 , n259282 , n259283 , n259284 , n259285 , 
     n259286 , n259287 , n259288 , n259289 , n259290 , n259291 , n259292 , n259293 , n259294 , n259295 , 
     n259296 , n259297 , n259298 , n259299 , n259300 , n259301 , n259302 , n259303 , n259304 , n259305 , 
     n259306 , n259307 , n259308 , n259309 , n259310 , n259311 , n259312 , n259313 , n259314 , n259315 , 
     n259316 , n259317 , n259318 , n259319 , n259320 , n259321 , n259322 , n259323 , n259324 , n259325 , 
     n259326 , n259327 , n259328 , n259329 , n259330 , n259331 , n259332 , n259333 , n259334 , n259335 , 
     n259336 , n259337 , n259338 , n259339 , n259340 , n259341 , n259342 , n259343 , n259344 , n259345 , 
     n259346 , n259347 , n259348 , n259349 , n259350 , n259351 , n259352 , n259353 , n259354 , n259355 , 
     n259356 , n259357 , n259358 , n259359 , n259360 , n259361 , n259362 , n259363 , n259364 , n259365 , 
     n259366 , n259367 , n259368 , n259369 , n259370 , n259371 , n259372 , n259373 , n259374 , n259375 , 
     n259376 , n259377 , n259378 , n259379 , n259380 , n259381 , n259382 , n259383 , n259384 , n259385 , 
     n259386 , n259387 , n259388 , n259389 , n259390 , n259391 , n259392 , n259393 , n259394 , n259395 , 
     n259396 , n259397 , n259398 , n259399 , n259400 , n259401 , n259402 , n259403 , n259404 , n259405 , 
     n259406 , n259407 , n259408 , n259409 , n259410 , n259411 , n259412 , n259413 , n259414 , n259415 , 
     n259416 , n259417 , n259418 , n259419 , n259420 , n259421 , n259422 , n259423 , n259424 , n259425 , 
     n259426 , n259427 , n259428 , n259429 , n259430 , n259431 , n259432 , n259433 , n259434 , n259435 , 
     n259436 , n259437 , n259438 , n259439 , n259440 , n259441 , n259442 , n259443 , n259444 , n259445 , 
     n259446 , n259447 , n259448 , n259449 , n259450 , n259451 , n259452 , n259453 , n259454 , n259455 , 
     n259456 , n259457 , n259458 , n259459 , n259460 , n259461 , n259462 , n259463 , n259464 , n259465 , 
     n259466 , n259467 , n259468 , n259469 , n259470 , n259471 , n259472 , n259473 , n259474 , n259475 , 
     n259476 , n259477 , n259478 , n259479 , n259480 , n259481 , n259482 , n259483 , n259484 , n259485 , 
     n259486 , n259487 , n259488 , n259489 , n259490 , n259491 , n259492 , n259493 , n259494 , n259495 , 
     n259496 , n259497 , n259498 , n259499 , n259500 , n259501 , n259502 , n259503 , n259504 , n259505 , 
     n259506 , n259507 , n259508 , n259509 , n259510 , n259511 , n259512 , n259513 , n259514 , n259515 , 
     n259516 , n259517 , n259518 , n259519 , n259520 , n259521 , n259522 , n259523 , n259524 , n259525 , 
     n259526 , n259527 , n259528 , n259529 , n259530 , n259531 , n259532 , n259533 , n259534 , n259535 , 
     n259536 , n259537 , n259538 , n259539 , n259540 , n259541 , n259542 , n259543 , n259544 , n259545 , 
     n259546 , n259547 , n259548 , n259549 , n259550 , n259551 , n259552 , n259553 , n259554 , n259555 , 
     n259556 , n259557 , n259558 , n259559 , n259560 , n259561 , n259562 , n259563 , n259564 , n259565 , 
     n259566 , n259567 , n259568 , n259569 , n259570 , n259571 , n259572 , n259573 , n259574 , n259575 , 
     n259576 , n259577 , n259578 , n259579 , n259580 , n259581 , n259582 , n259583 , n259584 , n259585 , 
     n259586 , n259587 , n259588 , n259589 , n259590 , n259591 , n259592 , n259593 , n259594 , n259595 , 
     n259596 , n259597 , n259598 , n259599 , n259600 , n259601 , n259602 , n259603 , n259604 , n259605 , 
     n259606 , n259607 , n259608 , n259609 , n259610 , n259611 , n259612 , n259613 , n259614 , n259615 , 
     n259616 , n259617 , n259618 , n259619 , n259620 , n259621 , n259622 , n259623 , n259624 , n259625 , 
     n259626 , n259627 , n259628 , n259629 , n259630 , n259631 , n259632 , n259633 , n259634 , n259635 , 
     n259636 , n259637 , n259638 , n259639 , n259640 , n259641 , n259642 , n259643 , n259644 , n259645 , 
     n259646 , n259647 , n259648 , n259649 , n259650 , n259651 , n259652 , n259653 , n259654 , n259655 , 
     n259656 , n259657 , n259658 , n259659 , n259660 , n259661 , n259662 , n259663 , n259664 , n259665 , 
     n259666 , n259667 , n259668 , n259669 , n259670 , n259671 , n259672 , n259673 , n259674 , n259675 , 
     n259676 , n259677 , n259678 , n259679 , n259680 , n259681 , n259682 , n259683 , n259684 , n259685 , 
     n259686 , n259687 , n259688 , n259689 , n259690 , n259691 , n259692 , n259693 , n259694 , n259695 , 
     n259696 , n259697 , n259698 , n259699 , n259700 , n259701 , n259702 , n259703 , n259704 , n259705 , 
     n259706 , n259707 , n259708 , n259709 , n259710 , n259711 , n259712 , n259713 , n259714 , n259715 , 
     n259716 , n259717 , n259718 , n259719 , n259720 , n259721 , n259722 , n259723 , n259724 , n259725 , 
     n259726 , n259727 , n259728 , n259729 , n259730 , n259731 , n259732 , n259733 , n259734 , n259735 , 
     n259736 , n259737 , n259738 , n259739 , n259740 , n259741 , n259742 , n259743 , n259744 , n259745 , 
     n259746 , n259747 , n259748 , n259749 , n259750 , n259751 , n259752 , n259753 , n259754 , n259755 , 
     n259756 , n259757 , n259758 , n259759 , n259760 , n259761 , n259762 , n259763 , n259764 , n259765 , 
     n259766 , n259767 , n259768 , n259769 , n259770 , n259771 , n259772 , n259773 , n259774 , n259775 , 
     n259776 , n259777 , n259778 , n259779 , n259780 , n259781 , n259782 , n259783 , n259784 , n259785 , 
     n259786 , n259787 , n259788 , n259789 , n259790 , n259791 , n259792 , n259793 , n259794 , n259795 , 
     n259796 , n259797 , n259798 , n259799 , n259800 , n259801 , n259802 , n259803 , n259804 , n259805 , 
     n259806 , n259807 , n259808 , n259809 , n259810 , n259811 , n259812 , n259813 , n259814 , n259815 , 
     n259816 , n259817 , n259818 , n259819 , n259820 , n259821 , n259822 , n259823 , n259824 , n259825 , 
     n259826 , n259827 , n259828 , n259829 , n259830 , n259831 , n259832 , n259833 , n259834 , n259835 , 
     n259836 , n259837 , n259838 , n259839 , n259840 , n259841 , n259842 , n259843 , n259844 , n259845 , 
     n259846 , n259847 , n259848 , n259849 , n259850 , n259851 , n259852 , n259853 , n259854 , n259855 , 
     n259856 , n259857 , n259858 , n259859 , n259860 , n259861 , n259862 , n259863 , n259864 , n259865 , 
     n259866 , n259867 , n259868 , n259869 , n259870 , n259871 , n259872 , n259873 , n259874 , n259875 , 
     n259876 , n259877 , n259878 , n259879 , n259880 , n259881 , n259882 , n259883 , n259884 , n259885 , 
     n259886 , n259887 , n259888 , n259889 , n259890 , n259891 , n259892 , n259893 , n259894 , n259895 , 
     n259896 , n259897 , n259898 , n259899 , n259900 , n259901 , n259902 , n259903 , n259904 , n259905 , 
     n259906 , n259907 , n259908 , n259909 , n259910 , n259911 , n259912 , n259913 , n259914 , n259915 , 
     n259916 , n259917 , n259918 , n259919 , n259920 , n259921 , n259922 , n259923 , n259924 , n259925 , 
     n259926 , n259927 , n259928 , n259929 , n259930 , n259931 , n259932 , n259933 , n259934 , n259935 , 
     n259936 , n259937 , n259938 , n259939 , n259940 , n259941 , n259942 , n259943 , n259944 , n259945 , 
     n259946 , n259947 , n259948 , n259949 , n259950 , n259951 , n259952 , n259953 , n259954 , n259955 , 
     n259956 , n259957 , n259958 , n259959 , n259960 , n259961 , n259962 , n259963 , n259964 , n259965 , 
     n259966 , n259967 , n259968 , n259969 , n259970 , n259971 , n259972 , n259973 , n259974 , n259975 , 
     n259976 , n259977 , n259978 , n259979 , n259980 , n259981 , n259982 , n259983 , n259984 , n259985 , 
     n259986 , n259987 , n259988 , n259989 , n259990 , n259991 , n259992 , n259993 , n259994 , n259995 , 
     n259996 , n259997 , n259998 , n259999 , n260000 , n260001 , n260002 , n260003 , n260004 , n260005 , 
     n260006 , n260007 , n260008 , n260009 , n260010 , n260011 , n260012 , n260013 , n260014 , n260015 , 
     n260016 , n260017 , n260018 , n260019 , n260020 , n260021 , n260022 , n260023 , n260024 , n260025 , 
     n260026 , n260027 , n260028 , n260029 , n260030 , n260031 , n260032 , n260033 , n260034 , n260035 , 
     n260036 , n260037 , n260038 , n260039 , n260040 , n260041 , n260042 , n260043 , n260044 , n260045 , 
     n260046 , n260047 , n260048 , n260049 , n260050 , n260051 , n260052 , n260053 , n260054 , n260055 , 
     n260056 , n260057 , n260058 , n260059 , n260060 , n260061 , n260062 , n260063 , n260064 , n260065 , 
     n260066 , n260067 , n260068 , n260069 , n260070 , n260071 , n260072 , n260073 , n260074 , n260075 , 
     n260076 , n260077 , n260078 , n260079 , n260080 , n260081 , n260082 , n260083 , n260084 , n260085 , 
     n260086 , n260087 , n260088 , n260089 , n260090 , n260091 , n260092 , n260093 , n260094 , n260095 , 
     n260096 , n260097 , n260098 , n260099 , n260100 , n260101 , n260102 , n260103 , n260104 , n260105 , 
     n260106 , n260107 , n260108 , n260109 , n260110 , n260111 , n260112 , n260113 , n260114 , n260115 , 
     n260116 , n260117 , n260118 , n260119 , n260120 , n260121 , n260122 , n260123 , n260124 , n260125 , 
     n260126 , n260127 , n260128 , n260129 , n260130 , n260131 , n260132 , n260133 , n260134 , n260135 , 
     n260136 , n260137 , n260138 , n260139 , n260140 , n260141 , n260142 , n260143 , n260144 , n260145 , 
     n260146 , n260147 , n260148 , n260149 , n260150 , n260151 , n260152 , n260153 , n260154 , n260155 , 
     n260156 , n260157 , n260158 , n260159 , n260160 , n260161 , n260162 , n260163 , n260164 , n260165 , 
     n260166 , n260167 , n260168 , n260169 , n260170 , n260171 , n260172 , n260173 , n260174 , n260175 , 
     n260176 , n260177 , n260178 , n260179 , n260180 , n260181 , n260182 , n260183 , n260184 , n260185 , 
     n260186 , n260187 , n260188 , n260189 , n260190 , n260191 , n260192 , n260193 , n260194 , n260195 , 
     n260196 , n260197 , n260198 , n260199 , n260200 , n260201 , n260202 , n260203 , n260204 , n260205 , 
     n260206 , n260207 , n260208 , n260209 , n260210 , n260211 , n260212 , n260213 , n260214 , n260215 , 
     n260216 , n260217 , n260218 , n260219 , n260220 , n260221 , n260222 , n260223 , n260224 , n260225 , 
     n260226 , n260227 , n260228 , n260229 , n260230 , n260231 , n260232 , n260233 , n260234 , n260235 , 
     n260236 , n260237 , n260238 , n260239 , n260240 , n260241 , n260242 , n260243 , n260244 , n260245 , 
     n260246 , n260247 , n260248 , n260249 , n260250 , n260251 , n260252 , n260253 , n260254 , n260255 , 
     n260256 , n260257 , n260258 , n260259 , n260260 , n260261 , n260262 , n260263 , n260264 , n260265 , 
     n260266 , n260267 , n260268 , n260269 , n260270 , n260271 , n260272 , n260273 , n260274 , n260275 , 
     n260276 , n260277 , n260278 , n260279 , n260280 , n260281 , n260282 , n260283 , n260284 , n260285 , 
     n260286 , n260287 , n260288 , n260289 , n260290 , n260291 , n260292 , n260293 , n260294 , n260295 , 
     n260296 , n260297 , n260298 , n260299 , n260300 , n260301 , n260302 , n260303 , n260304 , n260305 , 
     n260306 , n260307 , n260308 , n260309 , n260310 , n260311 , n260312 , n260313 , n260314 , n260315 , 
     n260316 , n260317 , n260318 , n260319 , n260320 , n260321 , n260322 , n260323 , n260324 , n260325 , 
     n260326 , n260327 , n260328 , n260329 , n260330 , n260331 , n260332 , n260333 , n260334 , n260335 , 
     n260336 , n260337 , n260338 , n260339 , n260340 , n260341 , n260342 , n260343 , n260344 , n260345 , 
     n260346 , n260347 , n260348 , n260349 , n260350 , n260351 , n260352 , n260353 , n260354 , n260355 , 
     n260356 , n260357 , n260358 , n260359 , n260360 , n260361 , n260362 , n260363 , n260364 , n260365 , 
     n260366 , n260367 , n260368 , n260369 , n260370 , n260371 , n260372 , n260373 , n260374 , n260375 , 
     n260376 , n260377 , n260378 , n260379 , n260380 , n260381 , n260382 , n260383 , n260384 , n260385 , 
     n260386 , n260387 , n260388 , n260389 , n260390 , n260391 , n260392 , n260393 , n260394 , n260395 , 
     n260396 , n260397 , n260398 , n260399 , n260400 , n260401 , n260402 , n260403 , n260404 , n260405 , 
     n260406 , n260407 , n260408 , n260409 , n260410 , n260411 , n260412 , n260413 , n260414 , n260415 , 
     n260416 , n260417 , n260418 , n260419 , n260420 , n260421 , n260422 , n260423 , n260424 , n260425 , 
     n260426 , n260427 , n260428 , n260429 , n260430 , n260431 , n260432 , n260433 , n260434 , n260435 , 
     n260436 , n260437 , n260438 , n260439 , n260440 , n260441 , n260442 , n260443 , n260444 , n260445 , 
     n260446 , n260447 , n260448 , n260449 , n260450 , n260451 , n260452 , n260453 , n260454 , n260455 , 
     n260456 , n260457 , n260458 , n260459 , n260460 , n260461 , n260462 , n260463 , n260464 , n260465 , 
     n260466 , n260467 , n260468 , n260469 , n260470 , n260471 , n260472 , n260473 , n260474 , n260475 , 
     n260476 , n260477 , n260478 , n260479 , n260480 , n260481 , n260482 , n260483 , n260484 , n260485 , 
     n260486 , n260487 , n260488 , n260489 , n260490 , n260491 , n260492 , n260493 , n260494 , n260495 , 
     n260496 , n260497 , n260498 , n260499 , n260500 , n260501 , n260502 , n260503 , n260504 , n260505 , 
     n260506 , n260507 , n260508 , n260509 , n260510 , n260511 , n260512 , n260513 , n260514 , n260515 , 
     n260516 , n260517 , n260518 , n260519 , n260520 , n260521 , n260522 , n260523 , n260524 , n260525 , 
     n260526 , n260527 , n260528 , n260529 , n260530 , n260531 , n260532 , n260533 , n260534 , n260535 , 
     n260536 , n260537 , n260538 , n260539 , n260540 , n260541 , n260542 , n260543 , n260544 , n260545 , 
     n260546 , n260547 , n260548 , n260549 , n260550 , n260551 , n260552 , n260553 , n260554 , n260555 , 
     n260556 , n260557 , n260558 , n260559 , n260560 , n260561 , n260562 , n260563 , n260564 , n260565 , 
     n260566 , n260567 , n260568 , n260569 , n260570 , n260571 , n260572 , n260573 , n260574 , n260575 , 
     n260576 , n260577 , n260578 , n260579 , n260580 , n260581 , n260582 , n260583 , n260584 , n260585 , 
     n260586 , n260587 , n260588 , n260589 , n260590 , n260591 , n260592 , n260593 , n260594 , n260595 , 
     n260596 , n260597 , n260598 , n260599 , n260600 , n260601 , n260602 , n260603 , n260604 , n260605 , 
     n260606 , n260607 , n260608 , n260609 , n260610 , n260611 , n260612 , n260613 , n260614 , n260615 , 
     n260616 , n260617 , n260618 , n260619 , n260620 , n260621 , n260622 , n260623 , n260624 , n260625 , 
     n260626 , n260627 , n260628 , n260629 , n260630 , n260631 , n260632 , n260633 , n260634 , n260635 , 
     n260636 , n260637 , n260638 , n260639 , n260640 , n260641 , n260642 , n260643 , n260644 , n260645 , 
     n260646 , n260647 , n260648 , n260649 , n260650 , n260651 , n260652 , n260653 , n260654 , n260655 , 
     n260656 , n260657 , n260658 , n260659 , n260660 , n260661 , n260662 , n260663 , n260664 , n260665 , 
     n260666 , n260667 , n260668 , n260669 , n260670 , n260671 , n260672 , n260673 , n260674 , n260675 , 
     n260676 , n260677 , n260678 , n260679 , n260680 , n260681 , n260682 , n260683 , n260684 , n260685 , 
     n260686 , n260687 , n260688 , n260689 , n260690 , n260691 , n260692 , n260693 , n260694 , n260695 , 
     n260696 , n260697 , n260698 , n260699 , n260700 , n260701 , n260702 , n260703 , n260704 , n260705 , 
     n260706 , n260707 , n260708 , n260709 , n260710 , n260711 , n260712 , n260713 , n260714 , n260715 , 
     n260716 , n260717 , n260718 , n260719 , n260720 , n260721 , n260722 , n260723 , n260724 , n260725 , 
     n260726 , n260727 , n260728 , n260729 , n260730 , n260731 , n260732 , n260733 , n260734 , n260735 , 
     n260736 , n260737 , n260738 , n260739 , n260740 , n260741 , n260742 , n260743 , n260744 , n260745 , 
     n260746 , n260747 , n260748 , n260749 , n260750 , n260751 , n260752 , n260753 , n260754 , n260755 , 
     n260756 , n260757 , n260758 , n260759 , n260760 , n260761 , n260762 , n260763 , n260764 , n260765 , 
     n260766 , n260767 , n260768 , n260769 , n260770 , n260771 , n260772 , n260773 , n260774 , n260775 , 
     n260776 , n260777 , n260778 , n260779 , n260780 , n260781 , n260782 , n260783 , n260784 , n260785 , 
     n260786 , n260787 , n260788 , n260789 , n260790 , n260791 , n260792 , n260793 , n260794 , n260795 , 
     n260796 , n260797 , n260798 , n260799 , n260800 , n260801 , n260802 , n260803 , n260804 , n260805 , 
     n260806 , n260807 , n260808 , n260809 , n260810 , n260811 , n260812 , n260813 , n260814 , n260815 , 
     n260816 , n260817 , n260818 , n260819 , n260820 , n260821 , n260822 , n260823 , n260824 , n260825 , 
     n260826 , n260827 , n260828 , n260829 , n260830 , n260831 , n260832 , n260833 , n260834 , n260835 , 
     n260836 , n260837 , n260838 , n260839 , n260840 , n260841 , n260842 , n260843 , n260844 , n260845 , 
     n260846 , n260847 , n260848 , n260849 , n260850 , n260851 , n260852 , n260853 , n260854 , n260855 , 
     n260856 , n260857 , n260858 , n260859 , n260860 , n260861 , n260862 , n260863 , n260864 , n260865 , 
     n260866 , n260867 , n260868 , n260869 , n260870 , n260871 , n260872 , n260873 , n260874 , n260875 , 
     n260876 , n260877 , n260878 , n260879 , n260880 , n260881 , n260882 , n260883 , n260884 , n260885 , 
     n260886 , n260887 , n260888 , n260889 , n260890 , n260891 , n260892 , n260893 , n260894 , n260895 , 
     n260896 , n260897 , n260898 , n260899 , n260900 , n260901 , n260902 , n260903 , n260904 , n260905 , 
     n260906 , n260907 , n260908 , n260909 , n260910 , n260911 , n260912 , n260913 , n260914 , n260915 , 
     n260916 , n260917 , n260918 , n260919 , n260920 , n260921 , n260922 , n260923 , n260924 , n260925 , 
     n260926 , n260927 , n260928 , n260929 , n260930 , n260931 , n260932 , n260933 , n260934 , n260935 , 
     n260936 , n260937 , n260938 , n260939 , n260940 , n260941 , n260942 , n260943 , n260944 , n260945 , 
     n260946 , n260947 , n260948 , n260949 , n260950 , n260951 , n260952 , n260953 , n260954 , n260955 , 
     n260956 , n260957 , n260958 , n260959 , n260960 , n260961 , n260962 , n260963 , n260964 , n260965 , 
     n260966 , n260967 , n260968 , n260969 , n260970 , n260971 , n260972 , n260973 , n260974 , n260975 , 
     n260976 , n260977 , n260978 , n260979 , n260980 , n260981 , n260982 , n260983 , n260984 , n260985 , 
     n260986 , n260987 , n260988 , n260989 , n260990 , n260991 , n260992 , n260993 , n260994 , n260995 , 
     n260996 , n260997 , n260998 , n260999 , n261000 , n261001 , n261002 , n261003 , n261004 , n261005 , 
     n261006 , n261007 , n261008 , n261009 , n261010 , n261011 , n261012 , n261013 , n261014 , n261015 , 
     n261016 , n261017 , n261018 , n261019 , n261020 , n261021 , n261022 , n261023 , n261024 , n261025 , 
     n261026 , n261027 , n261028 , n261029 , n261030 , n261031 , n261032 , n261033 , n261034 , n261035 , 
     n261036 , n261037 , n261038 , n261039 , n261040 , n261041 , n261042 , n261043 , n261044 , n261045 , 
     n261046 , n261047 , n261048 , n261049 , n261050 , n261051 , n261052 , n261053 , n261054 , n261055 , 
     n261056 , n261057 , n261058 , n261059 , n261060 , n261061 , n261062 , n261063 , n261064 , n261065 , 
     n261066 , n261067 , n261068 , n261069 , n261070 , n261071 , n261072 , n261073 , n261074 , n261075 , 
     n261076 , n261077 , n261078 , n261079 , n261080 , n261081 , n261082 , n261083 , n261084 , n261085 , 
     n261086 , n261087 , n261088 , n261089 , n261090 , n261091 , n261092 , n261093 , n261094 , n261095 , 
     n261096 , n261097 , n261098 , n261099 , n261100 , n261101 , n261102 , n261103 , n261104 , n261105 , 
     n261106 , n261107 , n261108 , n261109 , n261110 , n261111 , n261112 , n261113 , n261114 , n261115 , 
     n261116 , n261117 , n261118 , n261119 , n261120 , n261121 , n261122 , n261123 , n261124 , n261125 , 
     n261126 , n261127 , n261128 , n261129 , n261130 , n261131 , n261132 , n261133 , n261134 , n261135 , 
     n261136 , n261137 , n261138 , n261139 , n261140 , n261141 , n261142 , n261143 , n261144 , n261145 , 
     n261146 , n261147 , n261148 , n261149 , n261150 , n261151 , n261152 , n261153 , n261154 , n261155 , 
     n261156 , n261157 , n261158 , n261159 , n261160 , n261161 , n261162 , n261163 , n261164 , n261165 , 
     n261166 , n261167 , n261168 , n261169 , n261170 , n261171 , n261172 , n261173 , n261174 , n261175 , 
     n261176 , n261177 , n261178 , n261179 , n261180 , n261181 , n261182 , n261183 , n261184 , n261185 , 
     n261186 , n261187 , n261188 , n261189 , n261190 , n261191 , n261192 , n261193 , n261194 , n261195 , 
     n261196 , n261197 , n261198 , n261199 , n261200 , n261201 , n261202 , n261203 , n261204 , n261205 , 
     n261206 , n261207 , n261208 , n261209 , n261210 , n261211 , n261212 , n261213 , n261214 , n261215 , 
     n261216 , n261217 , n261218 , n261219 , n261220 , n261221 , n261222 , n261223 , n261224 , n261225 , 
     n261226 , n261227 , n261228 , n261229 , n261230 , n261231 , n261232 , n261233 , n261234 , n261235 , 
     n261236 , n261237 , n261238 , n261239 , n261240 , n261241 , n261242 , n261243 , n261244 , n261245 , 
     n261246 , n261247 , n261248 , n261249 , n261250 , n261251 , n261252 , n261253 , n261254 , n261255 , 
     n261256 , n261257 , n261258 , n261259 , n261260 , n261261 , n261262 , n261263 , n261264 , n261265 , 
     n261266 , n261267 , n261268 , n261269 , n261270 , n261271 , n261272 , n261273 , n261274 , n261275 , 
     n261276 , n261277 , n261278 , n261279 , n261280 , n261281 , n261282 , n261283 , n261284 , n261285 , 
     n261286 , n261287 , n261288 , n261289 , n261290 , n261291 , n261292 , n261293 , n261294 , n261295 , 
     n261296 , n261297 , n261298 , n261299 , n261300 , n261301 , n261302 , n261303 , n261304 , n261305 , 
     n261306 , n261307 , n261308 , n261309 , n261310 , n261311 , n261312 , n261313 , n261314 , n261315 , 
     n261316 , n261317 , n261318 , n261319 , n261320 , n261321 , n261322 , n261323 , n261324 , n261325 , 
     n261326 , n261327 , n261328 , n261329 , n261330 , n261331 , n261332 , n261333 , n261334 , n261335 , 
     n261336 , n261337 , n261338 , n261339 , n261340 , n261341 , n261342 , n261343 , n261344 , n261345 , 
     n261346 , n261347 , n261348 , n261349 , n261350 , n261351 , n261352 , n261353 , n261354 , n261355 , 
     n261356 , n261357 , n261358 , n261359 , n261360 , n261361 , n261362 , n261363 , n261364 , n261365 , 
     n261366 , n261367 , n261368 , n261369 , n261370 , n261371 , n261372 , n261373 , n261374 , n261375 , 
     n261376 , n261377 , n261378 , n261379 , n261380 , n261381 , n261382 , n261383 , n261384 , n261385 , 
     n261386 , n261387 , n261388 , n261389 , n261390 , n261391 , n261392 , n261393 , n261394 , n261395 , 
     n261396 , n261397 , n261398 , n261399 , n261400 , n261401 , n261402 , n261403 , n261404 , n261405 , 
     n261406 , n261407 , n261408 , n261409 , n261410 , n261411 , n261412 , n261413 , n261414 , n261415 , 
     n261416 , n261417 , n261418 , n261419 , n261420 , n261421 , n261422 , n261423 , n261424 , n261425 , 
     n261426 , n261427 , n261428 , n261429 , n261430 , n261431 , n261432 , n261433 , n261434 , n261435 , 
     n261436 , n261437 , n261438 , n261439 , n261440 , n261441 , n261442 , n261443 , n261444 , n261445 , 
     n261446 , n261447 , n261448 , n261449 , n261450 , n261451 , n261452 , n261453 , n261454 , n261455 , 
     n261456 , n261457 , n261458 , n261459 , n261460 , n261461 , n261462 , n261463 , n261464 , n261465 , 
     n261466 , n261467 , n261468 , n261469 , n261470 , n261471 , n261472 , n261473 , n261474 , n261475 , 
     n261476 , n261477 , n261478 , n261479 , n261480 , n261481 , n261482 , n261483 , n261484 , n261485 , 
     n261486 , n261487 , n261488 , n261489 , n261490 , n261491 , n261492 , n261493 , n261494 , n261495 , 
     n261496 , n261497 , n261498 , n261499 , n261500 , n261501 , n261502 , n261503 , n261504 , n261505 , 
     n261506 , n261507 , n261508 , n261509 , n261510 , n261511 , n261512 , n261513 , n261514 , n261515 , 
     n261516 , n261517 , n261518 , n261519 , n261520 , n261521 , n261522 , n261523 , n261524 , n261525 , 
     n261526 , n261527 , n261528 , n261529 , n261530 , n261531 , n261532 , n261533 , n261534 , n261535 , 
     n261536 , n261537 , n261538 , n261539 , n261540 , n261541 , n261542 , n261543 , n261544 , n261545 , 
     n261546 , n261547 , n261548 , n261549 , n261550 , n261551 , n261552 , n261553 , n261554 , n261555 , 
     n261556 , n261557 , n261558 , n261559 , n261560 , n261561 , n261562 , n261563 , n261564 , n261565 , 
     n261566 , n261567 , n261568 , n261569 , n261570 , n261571 , n261572 , n261573 , n261574 , n261575 , 
     n261576 , n261577 , n261578 , n261579 , n261580 , n261581 , n261582 , n261583 , n261584 , n261585 , 
     n261586 , n261587 , n261588 , n261589 , n261590 , n261591 , n261592 , n261593 , n261594 , n261595 , 
     n261596 , n261597 , n261598 , n261599 , n261600 , n261601 , n261602 , n261603 , n261604 , n261605 , 
     n261606 , n261607 , n261608 , n261609 , n261610 , n261611 , n261612 , n261613 , n261614 , n261615 , 
     n261616 , n261617 , n261618 , n261619 , n261620 , n261621 , n261622 , n261623 , n261624 , n261625 , 
     n261626 , n261627 , n261628 , n261629 , n261630 , n261631 , n261632 , n261633 , n261634 , n261635 , 
     n261636 , n261637 , n261638 , n261639 , n261640 , n261641 , n261642 , n261643 , n261644 , n261645 , 
     n261646 , n261647 , n261648 , n261649 , n261650 , n261651 , n261652 , n261653 , n261654 , n261655 , 
     n261656 , n261657 , n261658 , n261659 , n261660 , n261661 , n261662 , n261663 , n261664 , n261665 , 
     n261666 , n261667 , n261668 , n261669 , n261670 , n261671 , n261672 , n261673 , n261674 , n261675 , 
     n261676 , n261677 , n261678 , n261679 , n261680 , n261681 , n261682 , n261683 , n261684 , n261685 , 
     n261686 , n261687 , n261688 , n261689 , n261690 , n261691 , n261692 , n261693 , n261694 , n261695 , 
     n261696 , n261697 , n261698 , n261699 , n261700 , n261701 , n261702 , n261703 , n261704 , n261705 , 
     n261706 , n261707 , n261708 , n261709 , n261710 , n261711 , n261712 , n261713 , n261714 , n261715 , 
     n261716 , n261717 , n261718 , n261719 , n261720 , n261721 , n261722 , n261723 , n261724 , n261725 , 
     n261726 , n261727 , n261728 , n261729 , n261730 , n261731 , n261732 , n261733 , n261734 , n261735 , 
     n261736 , n261737 , n261738 , n261739 , n261740 , n261741 , n261742 , n261743 , n261744 , n261745 , 
     n261746 , n261747 , n261748 , n261749 , n261750 , n261751 , n261752 , n261753 , n261754 , n261755 , 
     n261756 , n261757 , n261758 , n261759 , n261760 , n261761 , n261762 , n261763 , n261764 , n261765 , 
     n261766 , n261767 , n261768 , n261769 , n261770 , n261771 , n261772 , n261773 , n261774 , n261775 , 
     n261776 , n261777 , n261778 , n261779 , n261780 , n261781 , n261782 , n261783 , n261784 , n261785 , 
     n261786 , n261787 , n261788 , n261789 , n261790 , n261791 , n261792 , n261793 , n261794 , n261795 , 
     n261796 , n261797 , n261798 , n261799 , n261800 , n261801 , n261802 , n261803 , n261804 , n261805 , 
     n261806 , n261807 , n261808 , n261809 , n261810 , n261811 , n261812 , n261813 , n261814 , n261815 , 
     n261816 , n261817 , n261818 , n261819 , n261820 , n261821 , n261822 , n261823 , n261824 , n261825 , 
     n261826 , n261827 , n261828 , n261829 , n261830 , n261831 , n261832 , n261833 , n261834 , n261835 , 
     n261836 , n261837 , n261838 , n261839 , n261840 , n261841 , n261842 , n261843 , n261844 , n261845 , 
     n261846 , n261847 , n261848 , n261849 , n261850 , n261851 , n261852 , n261853 , n261854 , n261855 , 
     n261856 , n261857 , n261858 , n261859 , n261860 , n261861 , n261862 , n261863 , n261864 , n261865 , 
     n261866 , n261867 , n261868 , n261869 , n261870 , n261871 , n261872 , n261873 , n261874 , n261875 , 
     n261876 , n261877 , n261878 , n261879 , n261880 , n261881 , n261882 , n261883 , n261884 , n261885 , 
     n261886 , n261887 , n261888 , n261889 , n261890 , n261891 , n261892 , n261893 , n261894 , n261895 , 
     n261896 , n261897 , n261898 , n261899 , n261900 , n261901 , n261902 , n261903 , n261904 , n261905 , 
     n261906 , n261907 , n261908 , n261909 , n261910 , n261911 , n261912 , n261913 , n261914 , n261915 , 
     n261916 , n261917 , n261918 , n261919 , n261920 , n261921 , n261922 , n261923 , n261924 , n261925 , 
     n261926 , n261927 , n261928 , n261929 , n261930 , n261931 , n261932 , n261933 , n261934 , n261935 , 
     n261936 , n261937 , n261938 , n261939 , n261940 , n261941 , n261942 , n261943 , n261944 , n261945 , 
     n261946 , n261947 , n261948 , n261949 , n261950 , n261951 , n261952 , n261953 , n261954 , n261955 , 
     n261956 , n261957 , n261958 , n261959 , n261960 , n261961 , n261962 , n261963 , n261964 , n261965 , 
     n261966 , n261967 , n261968 , n261969 , n261970 , n261971 , n261972 , n261973 , n261974 , n261975 , 
     n261976 , n261977 , n261978 , n261979 , n261980 , n261981 , n261982 , n261983 , n261984 , n261985 , 
     n261986 , n261987 , n261988 , n261989 , n261990 , n261991 , n261992 , n261993 , n261994 , n261995 , 
     n261996 , n261997 , n261998 , n261999 , n262000 , n262001 , n262002 , n262003 , n262004 , n262005 , 
     n262006 , n262007 , n262008 , n262009 , n262010 , n262011 , n262012 , n262013 , n262014 , n262015 , 
     n262016 , n262017 , n262018 , n262019 , n262020 , n262021 , n262022 , n262023 , n262024 , n262025 , 
     n262026 , n262027 , n262028 , n262029 , n262030 , n262031 , n262032 , n262033 , n262034 , n262035 , 
     n262036 , n262037 , n262038 , n262039 , n262040 , n262041 , n262042 , n262043 , n262044 , n262045 , 
     n262046 , n262047 , n262048 , n262049 , n262050 , n262051 , n262052 , n262053 , n262054 , n262055 , 
     n262056 , n262057 , n262058 , n262059 , n262060 , n262061 , n262062 , n262063 , n262064 , n262065 , 
     n262066 , n262067 , n262068 , n262069 , n262070 , n262071 , n262072 , n262073 , n262074 , n262075 , 
     n262076 , n262077 , n262078 , n262079 , n262080 , n262081 , n262082 , n262083 , n262084 , n262085 , 
     n262086 , n262087 , n262088 , n262089 , n262090 , n262091 , n262092 , n262093 , n262094 , n262095 , 
     n262096 , n262097 , n262098 , n262099 , n262100 , n262101 , n262102 , n262103 , n262104 , n262105 , 
     n262106 , n262107 , n262108 , n262109 , n262110 , n262111 , n262112 , n262113 , n262114 , n262115 , 
     n262116 , n262117 , n262118 , n262119 , n262120 , n262121 , n262122 , n262123 , n262124 , n262125 , 
     n262126 , n262127 , n262128 , n262129 , n262130 , n262131 , n262132 , n262133 , n262134 , n262135 , 
     n262136 , n262137 , n262138 , n262139 , n262140 , n262141 , n262142 , n262143 , n262144 , n262145 , 
     n262146 , n262147 , n262148 , n262149 , n262150 , n262151 , n262152 , n262153 , n262154 , n262155 , 
     n262156 , n262157 , n262158 , n262159 , n262160 , n262161 , n262162 , n262163 , n262164 , n262165 , 
     n262166 , n262167 , n262168 , n262169 , n262170 , n262171 , n262172 , n262173 , n262174 , n262175 , 
     n262176 , n262177 , n262178 , n262179 , n262180 , n262181 , n262182 , n262183 , n262184 , n262185 , 
     n262186 , n262187 , n262188 , n262189 , n262190 , n262191 , n262192 , n262193 , n262194 , n262195 , 
     n262196 , n262197 , n262198 , n262199 , n262200 , n262201 , n262202 , n262203 , n262204 , n262205 , 
     n262206 , n262207 , n262208 , n262209 , n262210 , n262211 , n262212 , n262213 , n262214 , n262215 , 
     n262216 , n262217 , n262218 , n262219 , n262220 , n262221 , n262222 , n262223 , n262224 , n262225 , 
     n262226 , n262227 , n262228 , n262229 , n262230 , n262231 , n262232 , n262233 , n262234 , n262235 , 
     n262236 , n262237 , n262238 , n262239 , n262240 , n262241 , n262242 , n262243 , n262244 , n262245 , 
     n262246 , n262247 , n262248 , n262249 , n262250 , n262251 , n262252 , n262253 , n262254 , n262255 , 
     n262256 , n262257 , n262258 , n262259 , n262260 , n262261 , n262262 , n262263 , n262264 , n262265 , 
     n262266 , n262267 , n262268 , n262269 , n262270 , n262271 , n262272 , n262273 , n262274 , n262275 , 
     n262276 , n262277 , n262278 , n262279 , n262280 , n262281 , n262282 , n262283 , n262284 , n262285 , 
     n262286 , n262287 , n262288 , n262289 , n262290 , n262291 , n262292 , n262293 , n262294 , n262295 , 
     n262296 , n262297 , n262298 , n262299 , n262300 , n262301 , n262302 , n262303 , n262304 , n262305 , 
     n262306 , n262307 , n262308 , n262309 , n262310 , n262311 , n262312 , n262313 , n262314 , n262315 , 
     n262316 , n262317 , n262318 , n262319 , n262320 , n262321 , n262322 , n262323 , n262324 , n262325 , 
     n262326 , n262327 , n262328 , n262329 , n262330 , n262331 , n262332 , n262333 , n262334 , n262335 , 
     n262336 , n262337 , n262338 , n262339 , n262340 , n262341 , n262342 , n262343 , n262344 , n262345 , 
     n262346 , n262347 , n262348 , n262349 , n262350 , n262351 , n262352 , n262353 , n262354 , n262355 , 
     n262356 , n262357 , n262358 , n262359 , n262360 , n262361 , n262362 , n262363 , n262364 , n262365 , 
     n262366 , n262367 , n262368 , n262369 , n262370 , n262371 , n262372 , n262373 , n262374 , n262375 , 
     n262376 , n262377 , n262378 , n262379 , n262380 , n262381 , n262382 , n262383 , n262384 , n262385 , 
     n262386 , n262387 , n262388 , n262389 , n262390 , n262391 , n262392 , n262393 , n262394 , n262395 , 
     n262396 , n262397 , n262398 , n262399 , n262400 , n262401 , n262402 , n262403 , n262404 , n262405 , 
     n262406 , n262407 , n262408 , n262409 , n262410 , n262411 , n262412 , n262413 , n262414 , n262415 , 
     n262416 , n262417 , n262418 , n262419 , n262420 , n262421 , n262422 , n262423 , n262424 , n262425 , 
     n262426 , n262427 , n262428 , n262429 , n262430 , n262431 , n262432 , n262433 , n262434 , n262435 , 
     n262436 , n262437 , n262438 , n262439 , n262440 , n262441 , n262442 , n262443 , n262444 , n262445 , 
     n262446 , n262447 , n262448 , n262449 , n262450 , n262451 , n262452 , n262453 , n262454 , n262455 , 
     n262456 , n262457 , n262458 , n262459 , n262460 , n262461 , n262462 , n262463 , n262464 , n262465 , 
     n262466 , n262467 , n262468 , n262469 , n262470 , n262471 , n262472 , n262473 , n262474 , n262475 , 
     n262476 , n262477 , n262478 , n262479 , n262480 , n262481 , n262482 , n262483 , n262484 , n262485 , 
     n262486 , n262487 , n262488 , n262489 , n262490 , n262491 , n262492 , n262493 , n262494 , n262495 , 
     n262496 , n262497 , n262498 , n262499 , n262500 , n262501 , n262502 , n262503 , n262504 , n262505 , 
     n262506 , n262507 , n262508 , n262509 , n262510 , n262511 , n262512 , n262513 , n262514 , n262515 , 
     n262516 , n262517 , n262518 , n262519 , n262520 , n262521 , n262522 , n262523 , n262524 , n262525 , 
     n262526 , n262527 , n262528 , n262529 , n262530 , n262531 , n262532 , n262533 , n262534 , n262535 , 
     n262536 , n262537 , n262538 , n262539 , n262540 , n262541 , n262542 , n262543 , n262544 , n262545 , 
     n262546 , n262547 , n262548 , n262549 , n262550 , n262551 , n262552 , n262553 , n262554 , n262555 , 
     n262556 , n262557 , n262558 , n262559 , n262560 , n262561 , n262562 , n262563 , n262564 , n262565 , 
     n262566 , n262567 , n262568 , n262569 , n262570 , n262571 , n262572 , n262573 , n262574 , n262575 , 
     n262576 , n262577 , n262578 , n262579 , n262580 , n262581 , n262582 , n262583 , n262584 , n262585 , 
     n262586 , n262587 , n262588 , n262589 , n262590 , n262591 , n262592 , n262593 , n262594 , n262595 , 
     n262596 , n262597 , n262598 , n262599 , n262600 , n262601 , n262602 , n262603 , n262604 , n262605 , 
     n262606 , n262607 , n262608 , n262609 , n262610 , n262611 , n262612 , n262613 , n262614 , n262615 , 
     n262616 , n262617 , n262618 , n262619 , n262620 , n262621 , n262622 , n262623 , n262624 , n262625 , 
     n262626 , n262627 , n262628 , n262629 , n262630 , n262631 , n262632 , n262633 , n262634 , n262635 , 
     n262636 , n262637 , n262638 , n262639 , n262640 , n262641 , n262642 , n262643 , n262644 , n262645 , 
     n262646 , n262647 , n262648 , n262649 , n262650 , n262651 , n262652 , n262653 , n262654 , n262655 , 
     n262656 , n262657 , n262658 , n262659 , n262660 , n262661 , n262662 , n262663 , n262664 , n262665 , 
     n262666 , n262667 , n262668 , n262669 , n262670 , n262671 , n262672 , n262673 , n262674 , n262675 , 
     n262676 , n262677 , n262678 , n262679 , n262680 , n262681 , n262682 , n262683 , n262684 , n262685 , 
     n262686 , n262687 , n262688 , n262689 , n262690 , n262691 , n262692 , n262693 , n262694 , n262695 , 
     n262696 , n262697 , n262698 , n262699 , n262700 , n262701 , n262702 , n262703 , n262704 , n262705 , 
     n262706 , n262707 , n262708 , n262709 , n262710 , n262711 , n262712 , n262713 , n262714 , n262715 , 
     n262716 , n262717 , n262718 , n262719 , n262720 , n262721 , n262722 , n262723 , n262724 , n262725 , 
     n262726 , n262727 , n262728 , n262729 , n262730 , n262731 , n262732 , n262733 , n262734 , n262735 , 
     n262736 , n262737 , n262738 , n262739 , n262740 , n262741 , n262742 , n262743 , n262744 , n262745 , 
     n262746 , n262747 , n262748 , n262749 , n262750 , n262751 , n262752 , n262753 , n262754 , n262755 , 
     n262756 , n262757 , n262758 , n262759 , n262760 , n262761 , n262762 , n262763 , n262764 , n262765 , 
     n262766 , n262767 , n262768 , n262769 , n262770 , n262771 , n262772 , n262773 , n262774 , n262775 , 
     n262776 , n262777 , n262778 , n262779 , n262780 , n262781 , n262782 , n262783 , n262784 , n262785 , 
     n262786 , n262787 , n262788 , n262789 , n262790 , n262791 , n262792 , n262793 , n262794 , n262795 , 
     n262796 , n262797 , n262798 , n262799 , n262800 , n262801 , n262802 , n262803 , n262804 , n262805 , 
     n262806 , n262807 , n262808 , n262809 , n262810 , n262811 , n262812 , n262813 , n262814 , n262815 , 
     n262816 , n262817 , n262818 , n262819 , n262820 , n262821 , n262822 , n262823 , n262824 , n262825 , 
     n262826 , n262827 , n262828 , n262829 , n262830 , n262831 , n262832 , n262833 , n262834 , n262835 , 
     n262836 , n262837 , n262838 , n262839 , n262840 , n262841 , n262842 , n262843 , n262844 , n262845 , 
     n262846 , n262847 , n262848 , n262849 , n262850 , n262851 , n262852 , n262853 , n262854 , n262855 , 
     n262856 , n262857 , n262858 , n262859 , n262860 , n262861 , n262862 , n262863 , n262864 , n262865 , 
     n262866 , n262867 , n262868 , n262869 , n262870 , n262871 , n262872 , n262873 , n262874 , n262875 , 
     n262876 , n262877 , n262878 , n262879 , n262880 , n262881 , n262882 , n262883 , n262884 , n262885 , 
     n262886 , n262887 , n262888 , n262889 , n262890 , n262891 , n262892 , n262893 , n262894 , n262895 , 
     n262896 , n262897 , n262898 , n262899 , n262900 , n262901 , n262902 , n262903 , n262904 , n262905 , 
     n262906 , n262907 , n262908 , n262909 , n262910 , n262911 , n262912 , n262913 , n262914 , n262915 , 
     n262916 , n262917 , n262918 , n262919 , n262920 , n262921 , n262922 , n262923 , n262924 , n262925 , 
     n262926 , n262927 , n262928 , n262929 , n262930 , n262931 , n262932 , n262933 , n262934 , n262935 , 
     n262936 , n262937 , n262938 , n262939 , n262940 , n262941 , n262942 , n262943 , n262944 , n262945 , 
     n262946 , n262947 , n262948 , n262949 , n262950 , n262951 , n262952 , n262953 , n262954 , n262955 , 
     n262956 , n262957 , n262958 , n262959 , n262960 , n262961 , n262962 , n262963 , n262964 , n262965 , 
     n262966 , n262967 , n262968 , n262969 , n262970 , n262971 , n262972 , n262973 , n262974 , n262975 , 
     n262976 , n262977 , n262978 , n262979 , n262980 , n262981 , n262982 , n262983 , n262984 , n262985 , 
     n262986 , n262987 , n262988 , n262989 , n262990 , n262991 , n262992 , n262993 , n262994 , n262995 , 
     n262996 , n262997 , n262998 , n262999 , n263000 , n263001 , n263002 , n263003 , n263004 , n263005 , 
     n263006 , n263007 , n263008 , n263009 , n263010 , n263011 , n263012 , n263013 , n263014 , n263015 , 
     n263016 , n263017 , n263018 , n263019 , n263020 , n263021 , n263022 , n263023 , n263024 , n263025 , 
     n263026 , n263027 , n263028 , n263029 , n263030 , n263031 , n263032 , n263033 , n263034 , n263035 , 
     n263036 , n263037 , n263038 , n263039 , n263040 , n263041 , n263042 , n263043 , n263044 , n263045 , 
     n263046 , n263047 , n263048 , n263049 , n263050 , n263051 , n263052 , n263053 , n263054 , n263055 , 
     n263056 , n263057 , n263058 , n263059 , n263060 , n263061 , n263062 , n263063 , n263064 , n263065 , 
     n263066 , n263067 , n263068 , n263069 , n263070 , n263071 , n263072 , n263073 , n263074 , n263075 , 
     n263076 , n263077 , n263078 , n263079 , n263080 , n263081 , n263082 , n263083 , n263084 , n263085 , 
     n263086 , n263087 , n263088 , n263089 , n263090 , n263091 , n263092 , n263093 , n263094 , n263095 , 
     n263096 , n263097 , n263098 , n263099 , n263100 , n263101 , n263102 , n263103 , n263104 , n263105 , 
     n263106 , n263107 , n263108 , n263109 , n263110 , n263111 , n263112 , n263113 , n263114 , n263115 , 
     n263116 , n263117 , n263118 , n263119 , n263120 , n263121 , n263122 , n263123 , n263124 , n263125 , 
     n263126 , n263127 , n263128 , n263129 , n263130 , n263131 , n263132 , n263133 , n263134 , n263135 , 
     n263136 , n263137 , n263138 , n263139 , n263140 , n263141 , n263142 , n263143 , n263144 , n263145 , 
     n263146 , n263147 , n263148 , n263149 , n263150 , n263151 , n263152 , n263153 , n263154 , n263155 , 
     n263156 , n263157 , n263158 , n263159 , n263160 , n263161 , n263162 , n263163 , n263164 , n263165 , 
     n263166 , n263167 , n263168 , n263169 , n263170 , n263171 , n263172 , n263173 , n263174 , n263175 , 
     n263176 , n263177 , n263178 , n263179 , n263180 , n263181 , n263182 , n263183 , n263184 , n263185 , 
     n263186 , n263187 , n263188 , n263189 , n263190 , n263191 , n263192 , n263193 , n263194 , n263195 , 
     n263196 , n263197 , n263198 , n263199 , n263200 , n263201 , n263202 , n263203 , n263204 , n263205 , 
     n263206 , n263207 , n263208 , n263209 , n263210 , n263211 , n263212 , n263213 , n263214 , n263215 , 
     n263216 , n263217 , n263218 , n263219 , n263220 , n263221 , n263222 , n263223 , n263224 , n263225 , 
     n263226 , n263227 , n263228 , n263229 , n263230 , n263231 , n263232 , n263233 , n263234 , n263235 , 
     n263236 , n263237 , n263238 , n263239 , n263240 , n263241 , n263242 , n263243 , n263244 , n263245 , 
     n263246 , n263247 , n263248 , n263249 , n263250 , n263251 , n263252 , n263253 , n263254 , n263255 , 
     n263256 , n263257 , n263258 , n263259 , n263260 , n263261 , n263262 , n263263 , n263264 , n263265 , 
     n263266 , n263267 , n263268 , n263269 , n263270 , n263271 , n263272 , n263273 , n263274 , n263275 , 
     n263276 , n263277 , n263278 , n263279 , n263280 , n263281 , n263282 , n263283 , n263284 , n263285 , 
     n263286 , n263287 , n263288 , n263289 , n263290 , n263291 , n263292 , n263293 , n263294 , n263295 , 
     n263296 , n263297 , n263298 , n263299 , n263300 , n263301 , n263302 , n263303 , n263304 , n263305 , 
     n263306 , n263307 , n263308 , n263309 , n263310 , n263311 , n263312 , n263313 , n263314 , n263315 , 
     n263316 , n263317 , n263318 , n263319 , n263320 , n263321 , n263322 , n263323 , n263324 , n263325 , 
     n263326 , n263327 , n263328 , n263329 , n263330 , n263331 , n263332 , n263333 , n263334 , n263335 , 
     n263336 , n263337 , n263338 , n263339 , n263340 , n263341 , n263342 , n263343 , n263344 , n263345 , 
     n263346 , n263347 , n263348 , n263349 , n263350 , n263351 , n263352 , n263353 , n263354 , n263355 , 
     n263356 , n263357 , n263358 , n263359 , n263360 , n263361 , n263362 , n263363 , n263364 , n263365 , 
     n263366 , n263367 , n263368 , n263369 , n263370 , n263371 , n263372 , n263373 , n263374 , n263375 , 
     n263376 , n263377 , n263378 , n263379 , n263380 , n263381 , n263382 , n263383 , n263384 , n263385 , 
     n263386 , n263387 , n263388 , n263389 , n263390 , n263391 , n263392 , n263393 , n263394 , n263395 , 
     n263396 , n263397 , n263398 , n263399 , n263400 , n263401 , n263402 , n263403 , n263404 , n263405 , 
     n263406 , n263407 , n263408 , n263409 , n263410 , n263411 , n263412 , n263413 , n263414 , n263415 , 
     n263416 , n263417 , n263418 , n263419 , n263420 , n263421 , n263422 , n263423 , n263424 , n263425 , 
     n263426 , n263427 , n263428 , n263429 , n263430 , n263431 , n263432 , n263433 , n263434 , n263435 , 
     n263436 , n263437 , n263438 , n263439 , n263440 , n263441 , n263442 , n263443 , n263444 , n263445 , 
     n263446 , n263447 , n263448 , n263449 , n263450 , n263451 , n263452 , n263453 , n263454 , n263455 , 
     n263456 , n263457 , n263458 , n263459 , n263460 , n263461 , n263462 , n263463 , n263464 , n263465 , 
     n263466 , n263467 , n263468 , n263469 , n263470 , n263471 , n263472 , n263473 , n263474 , n263475 , 
     n263476 , n263477 , n263478 , n263479 , n263480 , n263481 , n263482 , n263483 , n263484 , n263485 , 
     n263486 , n263487 , n263488 , n263489 , n263490 , n263491 , n263492 , n263493 , n263494 , n263495 , 
     n263496 , n263497 , n263498 , n263499 , n263500 , n263501 , n263502 , n263503 , n263504 , n263505 , 
     n263506 , n263507 , n263508 , n263509 , n263510 , n263511 , n263512 , n263513 , n263514 , n263515 , 
     n263516 , n263517 , n263518 , n263519 , n263520 , n263521 , n263522 , n263523 , n263524 , n263525 , 
     n263526 , n263527 , n263528 , n263529 , n263530 , n263531 , n263532 , n263533 , n263534 , n263535 , 
     n263536 , n263537 , n263538 , n263539 , n263540 , n263541 , n263542 , n263543 , n263544 , n263545 , 
     n263546 , n263547 , n263548 , n263549 , n263550 , n263551 , n263552 , n263553 , n263554 , n263555 , 
     n263556 , n263557 , n263558 , n263559 , n263560 , n263561 , n263562 , n263563 , n263564 , n263565 , 
     n263566 , n263567 , n263568 , n263569 , n263570 , n263571 , n263572 , n263573 , n263574 , n263575 , 
     n263576 , n263577 , n263578 , n263579 , n263580 , n263581 , n263582 , n263583 , n263584 , n263585 , 
     n263586 , n263587 , n263588 , n263589 , n263590 , n263591 , n263592 , n263593 , n263594 , n263595 , 
     n263596 , n263597 , n263598 , n263599 , n263600 , n263601 , n263602 , n263603 , n263604 , n263605 , 
     n263606 , n263607 , n263608 , n263609 , n263610 , n263611 , n263612 , n263613 , n263614 , n263615 , 
     n263616 , n263617 , n263618 , n263619 , n263620 , n263621 , n263622 , n263623 , n263624 , n263625 , 
     n263626 , n263627 , n263628 , n263629 , n263630 , n263631 , n263632 , n263633 , n263634 , n263635 , 
     n263636 , n263637 , n263638 , n263639 , n263640 , n263641 , n263642 , n263643 , n263644 , n263645 , 
     n263646 , n263647 , n263648 , n263649 , n263650 , n263651 , n263652 , n263653 , n263654 , n263655 , 
     n263656 , n263657 , n263658 , n263659 , n263660 , n263661 , n263662 , n263663 , n263664 , n263665 , 
     n263666 , n263667 , n263668 , n263669 , n263670 , n263671 , n263672 , n263673 , n263674 , n263675 , 
     n263676 , n263677 , n263678 , n263679 , n263680 , n263681 , n263682 , n263683 , n263684 , n263685 , 
     n263686 , n263687 , n263688 , n263689 , n263690 , n263691 , n263692 , n263693 , n263694 , n263695 , 
     n263696 , n263697 , n263698 , n263699 , n263700 , n263701 , n263702 , n263703 , n263704 , n263705 , 
     n263706 , n263707 , n263708 , n263709 , n263710 , n263711 , n263712 , n263713 , n263714 , n263715 , 
     n263716 , n263717 , n263718 , n263719 , n263720 , n263721 , n263722 , n263723 , n263724 , n263725 , 
     n263726 , n263727 , n263728 , n263729 , n263730 , n263731 , n263732 , n263733 , n263734 , n263735 , 
     n263736 , n263737 , n263738 , n263739 , n263740 , n263741 , n263742 , n263743 , n263744 , n263745 , 
     n263746 , n263747 , n263748 , n263749 , n263750 , n263751 , n263752 , n263753 , n263754 , n263755 , 
     n263756 , n263757 , n263758 , n263759 , n263760 , n263761 , n263762 , n263763 , n263764 , n263765 , 
     n263766 , n263767 , n263768 , n263769 , n263770 , n263771 , n263772 , n263773 , n263774 , n263775 , 
     n263776 , n263777 , n263778 , n263779 , n263780 , n263781 , n263782 , n263783 , n263784 , n263785 , 
     n263786 , n263787 , n263788 , n263789 , n263790 , n263791 , n263792 , n263793 , n263794 , n263795 , 
     n263796 , n263797 , n263798 , n263799 , n263800 , n263801 , n263802 , n263803 , n263804 , n263805 , 
     n263806 , n263807 , n263808 , n263809 , n263810 , n263811 , n263812 , n263813 , n263814 , n263815 , 
     n263816 , n263817 , n263818 , n263819 , n263820 , n263821 , n263822 , n263823 , n263824 , n263825 , 
     n263826 , n263827 , n263828 , n263829 , n263830 , n263831 , n263832 , n263833 , n263834 , n263835 , 
     n263836 , n263837 , n263838 , n263839 , n263840 , n263841 , n263842 , n263843 , n263844 , n263845 , 
     n263846 , n263847 , n263848 , n263849 , n263850 , n263851 , n263852 , n263853 , n263854 , n263855 , 
     n263856 , n263857 , n263858 , n263859 , n263860 , n263861 , n263862 , n263863 , n263864 , n263865 , 
     n263866 , n263867 , n263868 , n263869 , n263870 , n263871 , n263872 , n263873 , n263874 , n263875 , 
     n263876 , n263877 , n263878 , n263879 , n263880 , n263881 , n263882 , n263883 , n263884 , n263885 , 
     n263886 , n263887 , n263888 , n263889 , n263890 , n263891 , n263892 , n263893 , n263894 , n263895 , 
     n263896 , n263897 , n263898 , n263899 , n263900 , n263901 , n263902 , n263903 , n263904 , n263905 , 
     n263906 , n263907 , n263908 , n263909 , n263910 , n263911 , n263912 , n263913 , n263914 , n263915 , 
     n263916 , n263917 , n263918 , n263919 , n263920 , n263921 , n263922 , n263923 , n263924 , n263925 , 
     n263926 , n263927 , n263928 , n263929 , n263930 , n263931 , n263932 , n263933 , n263934 , n263935 , 
     n263936 , n263937 , n263938 , n263939 , n263940 , n263941 , n263942 , n263943 , n263944 , n263945 , 
     n263946 , n263947 , n263948 , n263949 , n263950 , n263951 , n263952 , n263953 , n263954 , n263955 , 
     n263956 , n263957 , n263958 , n263959 , n263960 , n263961 , n263962 , n263963 , n263964 , n263965 , 
     n263966 , n263967 , n263968 , n263969 , n263970 , n263971 , n263972 , n263973 , n263974 , n263975 , 
     n263976 , n263977 , n263978 , n263979 , n263980 , n263981 , n263982 , n263983 , n263984 , n263985 , 
     n263986 , n263987 , n263988 , n263989 , n263990 , n263991 , n263992 , n263993 , n263994 , n263995 , 
     n263996 , n263997 , n263998 , n263999 , n264000 , n264001 , n264002 , n264003 , n264004 , n264005 , 
     n264006 , n264007 , n264008 , n264009 , n264010 , n264011 , n264012 , n264013 , n264014 , n264015 , 
     n264016 , n264017 , n264018 , n264019 , n264020 , n264021 , n264022 , n264023 , n264024 , n264025 , 
     n264026 , n264027 , n264028 , n264029 , n264030 , n264031 , n264032 , n264033 , n264034 , n264035 , 
     n264036 , n264037 , n264038 , n264039 , n264040 , n264041 , n264042 , n264043 , n264044 , n264045 , 
     n264046 , n264047 , n264048 , n264049 , n264050 , n264051 , n264052 , n264053 , n264054 , n264055 , 
     n264056 , n264057 , n264058 , n264059 , n264060 , n264061 , n264062 , n264063 , n264064 , n264065 , 
     n264066 , n264067 , n264068 , n264069 , n264070 , n264071 , n264072 , n264073 , n264074 , n264075 , 
     n264076 , n264077 , n264078 , n264079 , n264080 , n264081 , n264082 , n264083 , n264084 , n264085 , 
     n264086 , n264087 , n264088 , n264089 , n264090 , n264091 , n264092 , n264093 , n264094 , n264095 , 
     n264096 , n264097 , n264098 , n264099 , n264100 , n264101 , n264102 , n264103 , n264104 , n264105 , 
     n264106 , n264107 , n264108 , n264109 , n264110 , n264111 , n264112 , n264113 , n264114 , n264115 , 
     n264116 , n264117 , n264118 , n264119 , n264120 , n264121 , n264122 , n264123 , n264124 , n264125 , 
     n264126 , n264127 , n264128 , n264129 , n264130 , n264131 , n264132 , n264133 , n264134 , n264135 , 
     n264136 , n264137 , n264138 , n264139 , n264140 , n264141 , n264142 , n264143 , n264144 , n264145 , 
     n264146 , n264147 , n264148 , n264149 , n264150 , n264151 , n264152 , n264153 , n264154 , n264155 , 
     n264156 , n264157 , n264158 , n264159 , n264160 , n264161 , n264162 , n264163 , n264164 , n264165 , 
     n264166 , n264167 , n264168 , n264169 , n264170 , n264171 , n264172 , n264173 , n264174 , n264175 , 
     n264176 , n264177 , n264178 , n264179 , n264180 , n264181 , n264182 , n264183 , n264184 , n264185 , 
     n264186 , n264187 , n264188 , n264189 , n264190 , n264191 , n264192 , n264193 , n264194 , n264195 , 
     n264196 , n264197 , n264198 , n264199 , n264200 , n264201 , n264202 , n264203 , n264204 , n264205 , 
     n264206 , n264207 , n264208 , n264209 , n264210 , n264211 , n264212 , n264213 , n264214 , n264215 , 
     n264216 , n264217 , n264218 , n264219 , n264220 , n264221 , n264222 , n264223 , n264224 , n264225 , 
     n264226 , n264227 , n264228 , n264229 , n264230 , n264231 , n264232 , n264233 , n264234 , n264235 , 
     n264236 , n264237 , n264238 , n264239 , n264240 , n264241 , n264242 , n264243 , n264244 , n264245 , 
     n264246 , n264247 , n264248 , n264249 , n264250 , n264251 , n264252 , n264253 , n264254 , n264255 , 
     n264256 , n264257 , n264258 , n264259 , n264260 , n264261 , n264262 , n264263 , n264264 , n264265 , 
     n264266 , n264267 , n264268 , n264269 , n264270 , n264271 , n264272 , n264273 , n264274 , n264275 , 
     n264276 , n264277 , n264278 , n264279 , n264280 , n264281 , n264282 , n264283 , n264284 , n264285 , 
     n264286 , n264287 , n264288 , n264289 , n264290 , n264291 , n264292 , n264293 , n264294 , n264295 , 
     n264296 , n264297 , n264298 , n264299 , n264300 , n264301 , n264302 , n264303 , n264304 , n264305 , 
     n264306 , n264307 , n264308 , n264309 , n264310 , n264311 , n264312 , n264313 , n264314 , n264315 , 
     n264316 , n264317 , n264318 , n264319 , n264320 , n264321 , n264322 , n264323 , n264324 , n264325 , 
     n264326 , n264327 , n264328 , n264329 , n264330 , n264331 , n264332 , n264333 , n264334 , n264335 , 
     n264336 , n264337 , n264338 , n264339 , n264340 , n264341 , n264342 , n264343 , n264344 , n264345 , 
     n264346 , n264347 , n264348 , n264349 , n264350 , n264351 , n264352 , n264353 , n264354 , n264355 , 
     n264356 , n264357 , n264358 , n264359 , n264360 , n264361 , n264362 , n264363 , n264364 , n264365 , 
     n264366 , n264367 , n264368 , n264369 , n264370 , n264371 , n264372 , n264373 , n264374 , n264375 , 
     n264376 , n264377 , n264378 , n264379 , n264380 , n264381 , n264382 , n264383 , n264384 , n264385 , 
     n264386 , n264387 , n264388 , n264389 , n264390 , n264391 , n264392 , n264393 , n264394 , n264395 , 
     n264396 , n264397 , n264398 , n264399 , n264400 , n264401 , n264402 , n264403 , n264404 , n264405 , 
     n264406 , n264407 , n264408 , n264409 , n264410 , n264411 , n264412 , n264413 , n264414 , n264415 , 
     n264416 , n264417 , n264418 , n264419 , n264420 , n264421 , n264422 , n264423 , n264424 , n264425 , 
     n264426 , n264427 , n264428 , n264429 , n264430 , n264431 , n264432 , n264433 , n264434 , n264435 , 
     n264436 , n264437 , n264438 , n264439 , n264440 , n264441 , n264442 , n264443 , n264444 , n264445 , 
     n264446 , n264447 , n264448 , n264449 , n264450 , n264451 , n264452 , n264453 , n264454 , n264455 , 
     n264456 , n264457 , n264458 , n264459 , n264460 , n264461 , n264462 , n264463 , n264464 , n264465 , 
     n264466 , n264467 , n264468 , n264469 , n264470 , n264471 , n264472 , n264473 , n264474 , n264475 , 
     n264476 , n264477 , n264478 , n264479 , n264480 , n264481 , n264482 , n264483 , n264484 , n264485 , 
     n264486 , n264487 , n264488 , n264489 , n264490 , n264491 , n264492 , n264493 , n264494 , n264495 , 
     n264496 , n264497 , n264498 , n264499 , n264500 , n264501 , n264502 , n264503 , n264504 , n264505 , 
     n264506 , n264507 , n264508 , n264509 , n264510 , n264511 , n264512 , n264513 , n264514 , n264515 , 
     n264516 , n264517 , n264518 , n264519 , n264520 , n264521 , n264522 , n264523 , n264524 , n264525 , 
     n264526 , n264527 , n264528 , n264529 , n264530 , n264531 , n264532 , n264533 , n264534 , n264535 , 
     n264536 , n264537 , n264538 , n264539 , n264540 , n264541 , n264542 , n264543 , n264544 , n264545 , 
     n264546 , n264547 , n264548 , n264549 , n264550 , n264551 , n264552 , n264553 , n264554 , n264555 , 
     n264556 , n264557 , n264558 , n264559 , n264560 , n264561 , n264562 , n264563 , n264564 , n264565 , 
     n264566 , n264567 , n264568 , n264569 , n264570 , n264571 , n264572 , n264573 , n264574 , n264575 , 
     n264576 , n264577 , n264578 , n264579 , n264580 , n264581 , n264582 , n264583 , n264584 , n264585 , 
     n264586 , n264587 , n264588 , n264589 , n264590 , n264591 , n264592 , n264593 , n264594 , n264595 , 
     n264596 , n264597 , n264598 , n264599 , n264600 , n264601 , n264602 , n264603 , n264604 , n264605 , 
     n264606 , n264607 , n264608 , n264609 , n264610 , n264611 , n264612 , n264613 , n264614 , n264615 , 
     n264616 , n264617 , n264618 , n264619 , n264620 , n264621 , n264622 , n264623 , n264624 , n264625 , 
     n264626 , n264627 , n264628 , n264629 , n264630 , n264631 , n264632 , n264633 , n264634 , n264635 , 
     n264636 , n264637 , n264638 , n264639 , n264640 , n264641 , n264642 , n264643 , n264644 , n264645 , 
     n264646 , n264647 , n264648 , n264649 , n264650 , n264651 , n264652 , n264653 , n264654 , n264655 , 
     n264656 , n264657 , n264658 , n264659 , n264660 , n264661 , n264662 , n264663 , n264664 , n264665 , 
     n264666 , n264667 , n264668 , n264669 , n264670 , n264671 , n264672 , n264673 , n264674 , n264675 , 
     n264676 , n264677 , n264678 , n264679 , n264680 , n264681 , n264682 , n264683 , n264684 , n264685 , 
     n264686 , n264687 , n264688 , n264689 , n264690 , n264691 , n264692 , n264693 , n264694 , n264695 , 
     n264696 , n264697 , n264698 , n264699 , n264700 , n264701 , n264702 , n264703 , n264704 , n264705 , 
     n264706 , n264707 , n264708 , n264709 , n264710 , n264711 , n264712 , n264713 , n264714 , n264715 , 
     n264716 , n264717 , n264718 , n264719 , n264720 , n264721 , n264722 , n264723 , n264724 , n264725 , 
     n264726 , n264727 , n264728 , n264729 , n264730 , n264731 , n264732 , n264733 , n264734 , n264735 , 
     n264736 , n264737 , n264738 , n264739 , n264740 , n264741 , n264742 , n264743 , n264744 , n264745 , 
     n264746 , n264747 , n264748 , n264749 , n264750 , n264751 , n264752 , n264753 , n264754 , n264755 , 
     n264756 , n264757 , n264758 , n264759 , n264760 , n264761 , n264762 , n264763 , n264764 , n264765 , 
     n264766 , n264767 , n264768 , n264769 , n264770 , n264771 , n264772 , n264773 , n264774 , n264775 , 
     n264776 , n264777 , n264778 , n264779 , n264780 , n264781 , n264782 , n264783 , n264784 , n264785 , 
     n264786 , n264787 , n264788 , n264789 , n264790 , n264791 , n264792 , n264793 , n264794 , n264795 , 
     n264796 , n264797 , n264798 , n264799 , n264800 , n264801 , n264802 , n264803 , n264804 , n264805 , 
     n264806 , n264807 , n264808 , n264809 , n264810 , n264811 , n264812 , n264813 , n264814 , n264815 , 
     n264816 , n264817 , n264818 , n264819 , n264820 , n264821 , n264822 , n264823 , n264824 , n264825 , 
     n264826 , n264827 , n264828 , n264829 , n264830 , n264831 , n264832 , n264833 , n264834 , n264835 , 
     n264836 , n264837 , n264838 , n264839 , n264840 , n264841 , n264842 , n264843 , n264844 , n264845 , 
     n264846 , n264847 , n264848 , n264849 , n264850 , n264851 , n264852 , n264853 , n264854 , n264855 , 
     n264856 , n264857 , n264858 , n264859 , n264860 , n264861 , n264862 , n264863 , n264864 , n264865 , 
     n264866 , n264867 , n264868 , n264869 , n264870 , n264871 , n264872 , n264873 , n264874 , n264875 , 
     n264876 , n264877 , n264878 , n264879 , n264880 , n264881 , n264882 , n264883 , n264884 , n264885 , 
     n264886 , n264887 , n264888 , n264889 , n264890 , n264891 , n264892 , n264893 , n264894 , n264895 , 
     n264896 , n264897 , n264898 , n264899 , n264900 , n264901 , n264902 , n264903 , n264904 , n264905 , 
     n264906 , n264907 , n264908 , n264909 , n264910 , n264911 , n264912 , n264913 , n264914 , n264915 , 
     n264916 , n264917 , n264918 , n264919 , n264920 , n264921 , n264922 , n264923 , n264924 , n264925 , 
     n264926 , n264927 , n264928 , n264929 , n264930 , n264931 , n264932 , n264933 , n264934 , n264935 , 
     n264936 , n264937 , n264938 , n264939 , n264940 , n264941 , n264942 , n264943 , n264944 , n264945 , 
     n264946 , n264947 , n264948 , n264949 , n264950 , n264951 , n264952 , n264953 , n264954 , n264955 , 
     n264956 , n264957 , n264958 , n264959 , n264960 , n264961 , n264962 , n264963 , n264964 , n264965 , 
     n264966 , n264967 , n264968 , n264969 , n264970 , n264971 , n264972 , n264973 , n264974 , n264975 , 
     n264976 , n264977 , n264978 , n264979 , n264980 , n264981 , n264982 , n264983 , n264984 , n264985 , 
     n264986 , n264987 , n264988 , n264989 , n264990 , n264991 , n264992 , n264993 , n264994 , n264995 , 
     n264996 , n264997 , n264998 , n264999 , n265000 , n265001 , n265002 , n265003 , n265004 , n265005 , 
     n265006 , n265007 , n265008 , n265009 , n265010 , n265011 , n265012 , n265013 , n265014 , n265015 , 
     n265016 , n265017 , n265018 , n265019 , n265020 , n265021 , n265022 , n265023 , n265024 , n265025 , 
     n265026 , n265027 , n265028 , n265029 , n265030 , n265031 , n265032 , n265033 , n265034 , n265035 , 
     n265036 , n265037 , n265038 , n265039 , n265040 , n265041 , n265042 , n265043 , n265044 , n265045 , 
     n265046 , n265047 , n265048 , n265049 , n265050 , n265051 , n265052 , n265053 , n265054 , n265055 , 
     n265056 , n265057 , n265058 , n265059 , n265060 , n265061 , n265062 , n265063 , n265064 , n265065 , 
     n265066 , n265067 , n265068 , n265069 , n265070 , n265071 , n265072 , n265073 , n265074 , n265075 , 
     n265076 , n265077 , n265078 , n265079 , n265080 , n265081 , n265082 , n265083 , n265084 , n265085 , 
     n265086 , n265087 , n265088 , n265089 , n265090 , n265091 , n265092 , n265093 , n265094 , n265095 , 
     n265096 , n265097 , n265098 , n265099 , n265100 , n265101 , n265102 , n265103 , n265104 , n265105 , 
     n265106 , n265107 , n265108 , n265109 , n265110 , n265111 , n265112 , n265113 , n265114 , n265115 , 
     n265116 , n265117 , n265118 , n265119 , n265120 , n265121 , n265122 , n265123 , n265124 , n265125 , 
     n265126 , n265127 , n265128 , n265129 , n265130 , n265131 , n265132 , n265133 , n265134 , n265135 , 
     n265136 , n265137 , n265138 , n265139 , n265140 , n265141 , n265142 , n265143 , n265144 , n265145 , 
     n265146 , n265147 , n265148 , n265149 , n265150 , n265151 , n265152 , n265153 , n265154 , n265155 , 
     n265156 , n265157 , n265158 , n265159 , n265160 , n265161 , n265162 , n265163 , n265164 , n265165 , 
     n265166 , n265167 , n265168 , n265169 , n265170 , n265171 , n265172 , n265173 , n265174 , n265175 , 
     n265176 , n265177 , n265178 , n265179 , n265180 , n265181 , n265182 , n265183 , n265184 , n265185 , 
     n265186 , n265187 , n265188 , n265189 , n265190 , n265191 , n265192 , n265193 , n265194 , n265195 , 
     n265196 , n265197 , n265198 , n265199 , n265200 , n265201 , n265202 , n265203 , n265204 , n265205 , 
     n265206 , n265207 , n265208 , n265209 , n265210 , n265211 , n265212 , n265213 , n265214 , n265215 , 
     n265216 , n265217 , n265218 , n265219 , n265220 , n265221 , n265222 , n265223 , n265224 , n265225 , 
     n265226 , n265227 , n265228 , n265229 , n265230 , n265231 , n265232 , n265233 , n265234 , n265235 , 
     n265236 , n265237 , n265238 , n265239 , n265240 , n265241 , n265242 , n265243 , n265244 , n265245 , 
     n265246 , n265247 , n265248 , n265249 , n265250 , n265251 , n265252 , n265253 , n265254 , n265255 , 
     n265256 , n265257 , n265258 , n265259 , n265260 , n265261 , n265262 , n265263 , n265264 , n265265 , 
     n265266 , n265267 , n265268 , n265269 , n265270 , n265271 , n265272 , n265273 , n265274 , n265275 , 
     n265276 , n265277 , n265278 , n265279 , n265280 , n265281 , n265282 , n265283 , n265284 , n265285 , 
     n265286 , n265287 , n265288 , n265289 , n265290 , n265291 , n265292 , n265293 , n265294 , n265295 , 
     n265296 , n265297 , n265298 , n265299 , n265300 , n265301 , n265302 , n265303 , n265304 , n265305 , 
     n265306 , n265307 , n265308 , n265309 , n265310 , n265311 , n265312 , n265313 , n265314 , n265315 , 
     n265316 , n265317 , n265318 , n265319 , n265320 , n265321 , n265322 , n265323 , n265324 , n265325 , 
     n265326 , n265327 , n265328 , n265329 , n265330 , n265331 , n265332 , n265333 , n265334 , n265335 , 
     n265336 , n265337 , n265338 , n265339 , n265340 , n265341 , n265342 , n265343 , n265344 , n265345 , 
     n265346 , n265347 , n265348 , n265349 , n265350 , n265351 , n265352 , n265353 , n265354 , n265355 , 
     n265356 , n265357 , n265358 , n265359 , n265360 , n265361 , n265362 , n265363 , n265364 , n265365 , 
     n265366 , n265367 , n265368 , n265369 , n265370 , n265371 , n265372 , n265373 , n265374 , n265375 , 
     n265376 , n265377 , n265378 , n265379 , n265380 , n265381 , n265382 , n265383 , n265384 , n265385 , 
     n265386 , n265387 , n265388 , n265389 , n265390 , n265391 , n265392 , n265393 , n265394 , n265395 , 
     n265396 , n265397 , n265398 , n265399 , n265400 , n265401 , n265402 , n265403 , n265404 , n265405 , 
     n265406 , n265407 , n265408 , n265409 , n265410 , n265411 , n265412 , n265413 , n265414 , n265415 , 
     n265416 , n265417 , n265418 , n265419 , n265420 , n265421 , n265422 , n265423 , n265424 , n265425 , 
     n265426 , n265427 , n265428 , n265429 , n265430 , n265431 , n265432 , n265433 , n265434 , n265435 , 
     n265436 , n265437 , n265438 , n265439 , n265440 , n265441 , n265442 , n265443 , n265444 , n265445 , 
     n265446 , n265447 , n265448 , n265449 , n265450 , n265451 , n265452 , n265453 , n265454 , n265455 , 
     n265456 , n265457 , n265458 , n265459 , n265460 , n265461 , n265462 , n265463 , n265464 , n265465 , 
     n265466 , n265467 , n265468 , n265469 , n265470 , n265471 , n265472 , n265473 , n265474 , n265475 , 
     n265476 , n265477 , n265478 , n265479 , n265480 , n265481 , n265482 , n265483 , n265484 , n265485 , 
     n265486 , n265487 , n265488 , n265489 , n265490 , n265491 , n265492 , n265493 , n265494 , n265495 , 
     n265496 , n265497 , n265498 , n265499 , n265500 , n265501 , n265502 , n265503 , n265504 , n265505 , 
     n265506 , n265507 , n265508 , n265509 , n265510 , n265511 , n265512 , n265513 , n265514 , n265515 , 
     n265516 , n265517 , n265518 , n265519 , n265520 , n265521 , n265522 , n265523 , n265524 , n265525 , 
     n265526 , n265527 , n265528 , n265529 , n265530 , n265531 , n265532 , n265533 , n265534 , n265535 , 
     n265536 , n265537 , n265538 , n265539 , n265540 , n265541 , n265542 , n265543 , n265544 , n265545 , 
     n265546 , n265547 , n265548 , n265549 , n265550 , n265551 , n265552 , n265553 , n265554 , n265555 , 
     n265556 , n265557 , n265558 , n265559 , n265560 , n265561 , n265562 , n265563 , n265564 , n265565 , 
     n265566 , n265567 , n265568 , n265569 , n265570 , n265571 , n265572 , n265573 , n265574 , n265575 , 
     n265576 , n265577 , n265578 , n265579 , n265580 , n265581 , n265582 , n265583 , n265584 , n265585 , 
     n265586 , n265587 , n265588 , n265589 , n265590 , n265591 , n265592 , n265593 , n265594 , n265595 , 
     n265596 , n265597 , n265598 , n265599 , n265600 , n265601 , n265602 , n265603 , n265604 , n265605 , 
     n265606 , n265607 , n265608 , n265609 , n265610 , n265611 , n265612 , n265613 , n265614 , n265615 , 
     n265616 , n265617 , n265618 , n265619 , n265620 , n265621 , n265622 , n265623 , n265624 , n265625 , 
     n265626 , n265627 , n265628 , n265629 , n265630 , n265631 , n265632 , n265633 , n265634 , n265635 , 
     n265636 , n265637 , n265638 , n265639 , n265640 , n265641 , n265642 , n265643 , n265644 , n265645 , 
     n265646 , n265647 , n265648 , n265649 , n265650 , n265651 , n265652 , n265653 , n265654 , n265655 , 
     n265656 , n265657 , n265658 , n265659 , n265660 , n265661 , n265662 , n265663 , n265664 , n265665 , 
     n265666 , n265667 , n265668 , n265669 , n265670 , n265671 , n265672 , n265673 , n265674 , n265675 , 
     n265676 , n265677 , n265678 , n265679 , n265680 , n265681 , n265682 , n265683 , n265684 , n265685 , 
     n265686 , n265687 , n265688 , n265689 , n265690 , n265691 , n265692 , n265693 , n265694 , n265695 , 
     n265696 , n265697 , n265698 , n265699 , n265700 , n265701 , n265702 , n265703 , n265704 , n265705 , 
     n265706 , n265707 , n265708 , n265709 , n265710 , n265711 , n265712 , n265713 , n265714 , n265715 , 
     n265716 , n265717 , n265718 , n265719 , n265720 , n265721 , n265722 , n265723 , n265724 , n265725 , 
     n265726 , n265727 , n265728 , n265729 , n265730 , n265731 , n265732 , n265733 , n265734 , n265735 , 
     n265736 , n265737 , n265738 , n265739 , n265740 , n265741 , n265742 , n265743 , n265744 , n265745 , 
     n265746 , n265747 , n265748 , n265749 , n265750 , n265751 , n265752 , n265753 , n265754 , n265755 , 
     n265756 , n265757 , n265758 , n265759 , n265760 , n265761 , n265762 , n265763 , n265764 , n265765 , 
     n265766 , n265767 , n265768 , n265769 , n265770 , n265771 , n265772 , n265773 , n265774 , n265775 , 
     n265776 , n265777 , n265778 , n265779 , n265780 , n265781 , n265782 , n265783 , n265784 , n265785 , 
     n265786 , n265787 , n265788 , n265789 , n265790 , n265791 , n265792 , n265793 , n265794 , n265795 , 
     n265796 , n265797 , n265798 , n265799 , n265800 , n265801 , n265802 , n265803 , n265804 , n265805 , 
     n265806 , n265807 , n265808 , n265809 , n265810 , n265811 , n265812 , n265813 , n265814 , n265815 , 
     n265816 , n265817 , n265818 , n265819 , n265820 , n265821 , n265822 , n265823 , n265824 , n265825 , 
     n265826 , n265827 , n265828 , n265829 , n265830 , n265831 , n265832 , n265833 , n265834 , n265835 , 
     n265836 , n265837 , n265838 , n265839 , n265840 , n265841 , n265842 , n265843 , n265844 , n265845 , 
     n265846 , n265847 , n265848 , n265849 , n265850 , n265851 , n265852 , n265853 , n265854 , n265855 , 
     n265856 , n265857 , n265858 , n265859 , n265860 , n265861 , n265862 , n265863 , n265864 , n265865 , 
     n265866 , n265867 , n265868 , n265869 , n265870 , n265871 , n265872 , n265873 , n265874 , n265875 , 
     n265876 , n265877 , n265878 , n265879 , n265880 , n265881 , n265882 , n265883 , n265884 , n265885 , 
     n265886 , n265887 , n265888 , n265889 , n265890 , n265891 , n265892 , n265893 , n265894 , n265895 , 
     n265896 , n265897 , n265898 , n265899 , n265900 , n265901 , n265902 , n265903 , n265904 , n265905 , 
     n265906 , n265907 , n265908 , n265909 , n265910 , n265911 , n265912 , n265913 , n265914 , n265915 , 
     n265916 , n265917 , n265918 , n265919 , n265920 , n265921 , n265922 , n265923 , n265924 , n265925 , 
     n265926 , n265927 , n265928 , n265929 , n265930 , n265931 , n265932 , n265933 , n265934 , n265935 , 
     n265936 , n265937 , n265938 , n265939 , n265940 , n265941 , n265942 , n265943 , n265944 , n265945 , 
     n265946 , n265947 , n265948 , n265949 , n265950 , n265951 , n265952 , n265953 , n265954 , n265955 , 
     n265956 , n265957 , n265958 , n265959 , n265960 , n265961 , n265962 , n265963 , n265964 , n265965 , 
     n265966 , n265967 , n265968 , n265969 , n265970 , n265971 , n265972 , n265973 , n265974 , n265975 , 
     n265976 , n265977 , n265978 , n265979 , n265980 , n265981 , n265982 , n265983 , n265984 , n265985 , 
     n265986 , n265987 , n265988 , n265989 , n265990 , n265991 , n265992 , n265993 , n265994 , n265995 , 
     n265996 , n265997 , n265998 , n265999 , n266000 , n266001 , n266002 , n266003 , n266004 , n266005 , 
     n266006 , n266007 , n266008 , n266009 , n266010 , n266011 , n266012 , n266013 , n266014 , n266015 , 
     n266016 , n266017 , n266018 , n266019 , n266020 , n266021 , n266022 , n266023 , n266024 , n266025 , 
     n266026 , n266027 , n266028 , n266029 , n266030 , n266031 , n266032 , n266033 , n266034 , n266035 , 
     n266036 , n266037 , n266038 , n266039 , n266040 , n266041 , n266042 , n266043 , n266044 , n266045 , 
     n266046 , n266047 , n266048 , n266049 , n266050 , n266051 , n266052 , n266053 , n266054 , n266055 , 
     n266056 , n266057 , n266058 , n266059 , n266060 , n266061 , n266062 , n266063 , n266064 , n266065 , 
     n266066 , n266067 , n266068 , n266069 , n266070 , n266071 , n266072 , n266073 , n266074 , n266075 , 
     n266076 , n266077 , n266078 , n266079 , n266080 , n266081 , n266082 , n266083 , n266084 , n266085 , 
     n266086 , n266087 , n266088 , n266089 , n266090 , n266091 , n266092 , n266093 , n266094 , n266095 , 
     n266096 , n266097 , n266098 , n266099 , n266100 , n266101 , n266102 , n266103 , n266104 , n266105 , 
     n266106 , n266107 , n266108 , n266109 , n266110 , n266111 , n266112 , n266113 , n266114 , n266115 , 
     n266116 , n266117 , n266118 , n266119 , n266120 , n266121 , n266122 , n266123 , n266124 , n266125 , 
     n266126 , n266127 , n266128 , n266129 , n266130 , n266131 , n266132 , n266133 , n266134 , n266135 , 
     n266136 , n266137 , n266138 , n266139 , n266140 , n266141 , n266142 , n266143 , n266144 , n266145 , 
     n266146 , n266147 , n266148 , n266149 , n266150 , n266151 , n266152 , n266153 , n266154 , n266155 , 
     n266156 , n266157 , n266158 , n266159 , n266160 , n266161 , n266162 , n266163 , n266164 , n266165 , 
     n266166 , n266167 , n266168 , n266169 , n266170 , n266171 , n266172 , n266173 , n266174 , n266175 , 
     n266176 , n266177 , n266178 , n266179 , n266180 , n266181 , n266182 , n266183 , n266184 , n266185 , 
     n266186 , n266187 , n266188 , n266189 , n266190 , n266191 , n266192 , n266193 , n266194 , n266195 , 
     n266196 , n266197 , n266198 , n266199 , n266200 , n266201 , n266202 , n266203 , n266204 , n266205 , 
     n266206 , n266207 , n266208 , n266209 , n266210 , n266211 , n266212 , n266213 , n266214 , n266215 , 
     n266216 , n266217 , n266218 , n266219 , n266220 , n266221 , n266222 , n266223 , n266224 , n266225 , 
     n266226 , n266227 , n266228 , n266229 , n266230 , n266231 , n266232 , n266233 , n266234 , n266235 , 
     n266236 , n266237 , n266238 , n266239 , n266240 , n266241 , n266242 , n266243 , n266244 , n266245 , 
     n266246 , n266247 , n266248 , n266249 , n266250 , n266251 , n266252 , n266253 , n266254 , n266255 , 
     n266256 , n266257 , n266258 , n266259 , n266260 , n266261 , n266262 , n266263 , n266264 , n266265 , 
     n266266 , n266267 , n266268 , n266269 , n266270 , n266271 , n266272 , n266273 , n266274 , n266275 , 
     n266276 , n266277 , n266278 , n266279 , n266280 , n266281 , n266282 , n266283 , n266284 , n266285 , 
     n266286 , n266287 , n266288 , n266289 , n266290 , n266291 , n266292 , n266293 , n266294 , n266295 , 
     n266296 , n266297 , n266298 , n266299 , n266300 , n266301 , n266302 , n266303 , n266304 , n266305 , 
     n266306 , n266307 , n266308 , n266309 , n266310 , n266311 , n266312 , n266313 , n266314 , n266315 , 
     n266316 , n266317 , n266318 , n266319 , n266320 , n266321 , n266322 , n266323 , n266324 , n266325 , 
     n266326 , n266327 , n266328 , n266329 , n266330 , n266331 , n266332 , n266333 , n266334 , n266335 , 
     n266336 , n266337 , n266338 , n266339 , n266340 , n266341 , n266342 , n266343 , n266344 , n266345 , 
     n266346 , n266347 , n266348 , n266349 , n266350 , n266351 , n266352 , n266353 , n266354 , n266355 , 
     n266356 , n266357 , n266358 , n266359 , n266360 , n266361 , n266362 , n266363 , n266364 , n266365 , 
     n266366 , n266367 , n266368 , n266369 , n266370 , n266371 , n266372 , n266373 , n266374 , n266375 , 
     n266376 , n266377 , n266378 , n266379 , n266380 , n266381 , n266382 , n266383 , n266384 , n266385 , 
     n266386 , n266387 , n266388 , n266389 , n266390 , n266391 , n266392 , n266393 , n266394 , n266395 , 
     n266396 , n266397 , n266398 , n266399 , n266400 , n266401 , n266402 , n266403 , n266404 , n266405 , 
     n266406 , n266407 , n266408 , n266409 , n266410 , n266411 , n266412 , n266413 , n266414 , n266415 , 
     n266416 , n266417 , n266418 , n266419 , n266420 , n266421 , n266422 , n266423 , n266424 , n266425 , 
     n266426 , n266427 , n266428 , n266429 , n266430 , n266431 , n266432 , n266433 , n266434 , n266435 , 
     n266436 , n266437 , n266438 , n266439 , n266440 , n266441 , n266442 , n266443 , n266444 , n266445 , 
     n266446 , n266447 , n266448 , n266449 , n266450 , n266451 , n266452 , n266453 , n266454 , n266455 , 
     n266456 , n266457 , n266458 , n266459 , n266460 , n266461 , n266462 , n266463 , n266464 , n266465 , 
     n266466 , n266467 , n266468 , n266469 , n266470 , n266471 , n266472 , n266473 , n266474 , n266475 , 
     n266476 , n266477 , n266478 , n266479 , n266480 , n266481 , n266482 , n266483 , n266484 , n266485 , 
     n266486 , n266487 , n266488 , n266489 , n266490 , n266491 , n266492 , n266493 , n266494 , n266495 , 
     n266496 , n266497 , n266498 , n266499 , n266500 , n266501 , n266502 , n266503 , n266504 , n266505 , 
     n266506 , n266507 , n266508 , n266509 , n266510 , n266511 , n266512 , n266513 , n266514 , n266515 , 
     n266516 , n266517 , n266518 , n266519 , n266520 , n266521 , n266522 , n266523 , n266524 , n266525 , 
     n266526 , n266527 , n266528 , n266529 , n266530 , n266531 , n266532 , n266533 , n266534 , n266535 , 
     n266536 , n266537 , n266538 , n266539 , n266540 , n266541 , n266542 , n266543 , n266544 , n266545 , 
     n266546 , n266547 , n266548 , n266549 , n266550 , n266551 , n266552 , n266553 , n266554 , n266555 , 
     n266556 , n266557 , n266558 , n266559 , n266560 , n266561 , n266562 , n266563 , n266564 , n266565 , 
     n266566 , n266567 , n266568 , n266569 , n266570 , n266571 , n266572 , n266573 , n266574 , n266575 , 
     n266576 , n266577 , n266578 , n266579 , n266580 , n266581 , n266582 , n266583 , n266584 , n266585 , 
     n266586 , n266587 , n266588 , n266589 , n266590 , n266591 , n266592 , n266593 , n266594 , n266595 , 
     n266596 , n266597 , n266598 , n266599 , n266600 , n266601 , n266602 , n266603 , n266604 , n266605 , 
     n266606 , n266607 , n266608 , n266609 , n266610 , n266611 , n266612 , n266613 , n266614 , n266615 , 
     n266616 , n266617 , n266618 , n266619 , n266620 , n266621 , n266622 , n266623 , n266624 , n266625 , 
     n266626 , n266627 , n266628 , n266629 , n266630 , n266631 , n266632 , n266633 , n266634 , n266635 , 
     n266636 , n266637 , n266638 , n266639 , n266640 , n266641 , n266642 , n266643 , n266644 , n266645 , 
     n266646 , n266647 , n266648 , n266649 , n266650 , n266651 , n266652 , n266653 , n266654 , n266655 , 
     n266656 , n266657 , n266658 , n266659 , n266660 , n266661 , n266662 , n266663 , n266664 , n266665 , 
     n266666 , n266667 , n266668 , n266669 , n266670 , n266671 , n266672 , n266673 , n266674 , n266675 , 
     n266676 , n266677 , n266678 , n266679 , n266680 , n266681 , n266682 , n266683 , n266684 , n266685 , 
     n266686 , n266687 , n266688 , n266689 , n266690 , n266691 , n266692 , n266693 , n266694 , n266695 , 
     n266696 , n266697 , n266698 , n266699 , n266700 , n266701 , n266702 , n266703 , n266704 , n266705 , 
     n266706 , n266707 , n266708 , n266709 , n266710 , n266711 , n266712 , n266713 , n266714 , n266715 , 
     n266716 , n266717 , n266718 , n266719 , n266720 , n266721 , n266722 , n266723 , n266724 , n266725 , 
     n266726 , n266727 , n266728 , n266729 , n266730 , n266731 , n266732 , n266733 , n266734 , n266735 , 
     n266736 , n266737 , n266738 , n266739 , n266740 , n266741 , n266742 , n266743 , n266744 , n266745 , 
     n266746 , n266747 , n266748 , n266749 , n266750 , n266751 , n266752 , n266753 , n266754 , n266755 , 
     n266756 , n266757 , n266758 , n266759 , n266760 , n266761 , n266762 , n266763 , n266764 , n266765 , 
     n266766 , n266767 , n266768 , n266769 , n266770 , n266771 , n266772 , n266773 , n266774 , n266775 , 
     n266776 , n266777 , n266778 , n266779 , n266780 , n266781 , n266782 , n266783 , n266784 , n266785 , 
     n266786 , n266787 , n266788 , n266789 , n266790 , n266791 , n266792 , n266793 , n266794 , n266795 , 
     n266796 , n266797 , n266798 , n266799 , n266800 , n266801 , n266802 , n266803 , n266804 , n266805 , 
     n266806 , n266807 , n266808 , n266809 , n266810 , n266811 , n266812 , n266813 , n266814 , n266815 , 
     n266816 , n266817 , n266818 , n266819 , n266820 , n266821 , n266822 , n266823 , n266824 , n266825 , 
     n266826 , n266827 , n266828 , n266829 , n266830 , n266831 , n266832 , n266833 , n266834 , n266835 , 
     n266836 , n266837 , n266838 , n266839 , n266840 , n266841 , n266842 , n266843 , n266844 , n266845 , 
     n266846 , n266847 , n266848 , n266849 , n266850 , n266851 , n266852 , n266853 , n266854 , n266855 , 
     n266856 , n266857 , n266858 , n266859 , n266860 , n266861 , n266862 , n266863 , n266864 , n266865 , 
     n266866 , n266867 , n266868 , n266869 , n266870 , n266871 , n266872 , n266873 , n266874 , n266875 , 
     n266876 , n266877 , n266878 , n266879 , n266880 , n266881 , n266882 , n266883 , n266884 , n266885 , 
     n266886 , n266887 , n266888 , n266889 , n266890 , n266891 , n266892 , n266893 , n266894 , n266895 , 
     n266896 , n266897 , n266898 , n266899 , n266900 , n266901 , n266902 , n266903 , n266904 , n266905 , 
     n266906 , n266907 , n266908 , n266909 , n266910 , n266911 , n266912 , n266913 , n266914 , n266915 , 
     n266916 , n266917 , n266918 , n266919 , n266920 , n266921 , n266922 , n266923 , n266924 , n266925 , 
     n266926 , n266927 , n266928 , n266929 , n266930 , n266931 , n266932 , n266933 , n266934 , n266935 , 
     n266936 , n266937 , n266938 , n266939 , n266940 , n266941 , n266942 , n266943 , n266944 , n266945 , 
     n266946 , n266947 , n266948 , n266949 , n266950 , n266951 , n266952 , n266953 , n266954 , n266955 , 
     n266956 , n266957 , n266958 , n266959 , n266960 , n266961 , n266962 , n266963 , n266964 , n266965 , 
     n266966 , n266967 , n266968 , n266969 , n266970 , n266971 , n266972 , n266973 , n266974 , n266975 , 
     n266976 , n266977 , n266978 , n266979 , n266980 , n266981 , n266982 , n266983 , n266984 , n266985 , 
     n266986 , n266987 , n266988 , n266989 , n266990 , n266991 , n266992 , n266993 , n266994 , n266995 , 
     n266996 , n266997 , n266998 , n266999 , n267000 , n267001 , n267002 , n267003 , n267004 , n267005 , 
     n267006 , n267007 , n267008 , n267009 , n267010 , n267011 , n267012 , n267013 , n267014 , n267015 , 
     n267016 , n267017 , n267018 , n267019 , n267020 , n267021 , n267022 , n267023 , n267024 , n267025 , 
     n267026 , n267027 , n267028 , n267029 , n267030 , n267031 , n267032 , n267033 , n267034 , n267035 , 
     n267036 , n267037 , n267038 , n267039 , n267040 , n267041 , n267042 , n267043 , n267044 , n267045 , 
     n267046 , n267047 , n267048 , n267049 , n267050 , n267051 , n267052 , n267053 , n267054 , n267055 , 
     n267056 , n267057 , n267058 , n267059 , n267060 , n267061 , n267062 , n267063 , n267064 , n267065 , 
     n267066 , n267067 , n267068 , n267069 , n267070 , n267071 , n267072 , n267073 , n267074 , n267075 , 
     n267076 , n267077 , n267078 , n267079 , n267080 , n267081 , n267082 , n267083 , n267084 , n267085 , 
     n267086 , n267087 , n267088 , n267089 , n267090 , n267091 , n267092 , n267093 , n267094 , n267095 , 
     n267096 , n267097 , n267098 , n267099 , n267100 , n267101 , n267102 , n267103 , n267104 , n267105 , 
     n267106 , n267107 , n267108 , n267109 , n267110 , n267111 , n267112 , n267113 , n267114 , n267115 , 
     n267116 , n267117 , n267118 , n267119 , n267120 , n267121 , n267122 , n267123 , n267124 , n267125 , 
     n267126 , n267127 , n267128 , n267129 , n267130 , n267131 , n267132 , n267133 , n267134 , n267135 , 
     n267136 , n267137 , n267138 , n267139 , n267140 , n267141 , n267142 , n267143 , n267144 , n267145 , 
     n267146 , n267147 , n267148 , n267149 , n267150 , n267151 , n267152 , n267153 , n267154 , n267155 , 
     n267156 , n267157 , n267158 , n267159 , n267160 , n267161 , n267162 , n267163 , n267164 , n267165 , 
     n267166 , n267167 , n267168 , n267169 , n267170 , n267171 , n267172 , n267173 , n267174 , n267175 , 
     n267176 , n267177 , n267178 , n267179 , n267180 , n267181 , n267182 , n267183 , n267184 , n267185 , 
     n267186 , n267187 , n267188 , n267189 , n267190 , n267191 , n267192 , n267193 , n267194 , n267195 , 
     n267196 , n267197 , n267198 , n267199 , n267200 , n267201 , n267202 , n267203 , n267204 , n267205 , 
     n267206 , n267207 , n267208 , n267209 , n267210 , n267211 , n267212 , n267213 , n267214 , n267215 , 
     n267216 , n267217 , n267218 , n267219 , n267220 , n267221 , n267222 , n267223 , n267224 , n267225 , 
     n267226 , n267227 , n267228 , n267229 , n267230 , n267231 , n267232 , n267233 , n267234 , n267235 , 
     n267236 , n267237 , n267238 , n267239 , n267240 , n267241 , n267242 , n267243 , n267244 , n267245 , 
     n267246 , n267247 , n267248 , n267249 , n267250 , n267251 , n267252 , n267253 , n267254 , n267255 , 
     n267256 , n267257 , n267258 , n267259 , n267260 , n267261 , n267262 , n267263 , n267264 , n267265 , 
     n267266 , n267267 , n267268 , n267269 , n267270 , n267271 , n267272 , n267273 , n267274 , n267275 , 
     n267276 , n267277 , n267278 , n267279 , n267280 , n267281 , n267282 , n267283 , n267284 , n267285 , 
     n267286 , n267287 , n267288 , n267289 , n267290 , n267291 , n267292 , n267293 , n267294 , n267295 , 
     n267296 , n267297 , n267298 , n267299 , n267300 , n267301 , n267302 , n267303 , n267304 , n267305 , 
     n267306 , n267307 , n267308 , n267309 , n267310 , n267311 , n267312 , n267313 , n267314 , n267315 , 
     n267316 , n267317 , n267318 , n267319 , n267320 , n267321 , n267322 , n267323 , n267324 , n267325 , 
     n267326 , n267327 , n267328 , n267329 , n267330 , n267331 , n267332 , n267333 , n267334 , n267335 , 
     n267336 , n267337 , n267338 , n267339 , n267340 , n267341 , n267342 , n267343 , n267344 , n267345 , 
     n267346 , n267347 , n267348 , n267349 , n267350 , n267351 , n267352 , n267353 , n267354 , n267355 , 
     n267356 , n267357 , n267358 , n267359 , n267360 , n267361 , n267362 , n267363 , n267364 , n267365 , 
     n267366 , n267367 , n267368 , n267369 , n267370 , n267371 , n267372 , n267373 , n267374 , n267375 , 
     n267376 , n267377 , n267378 , n267379 , n267380 , n267381 , n267382 , n267383 , n267384 , n267385 , 
     n267386 , n267387 , n267388 , n267389 , n267390 , n267391 , n267392 , n267393 , n267394 , n267395 , 
     n267396 , n267397 , n267398 , n267399 , n267400 , n267401 , n267402 , n267403 , n267404 , n267405 , 
     n267406 , n267407 , n267408 , n267409 , n267410 , n267411 , n267412 , n267413 , n267414 , n267415 , 
     n267416 , n267417 , n267418 , n267419 , n267420 , n267421 , n267422 , n267423 , n267424 , n267425 , 
     n267426 , n267427 , n267428 , n267429 , n267430 , n267431 , n267432 , n267433 , n267434 , n267435 , 
     n267436 , n267437 , n267438 , n267439 , n267440 , n267441 , n267442 , n267443 , n267444 , n267445 , 
     n267446 , n267447 , n267448 , n267449 , n267450 , n267451 , n267452 , n267453 , n267454 , n267455 , 
     n267456 , n267457 , n267458 , n267459 , n267460 , n267461 , n267462 , n267463 , n267464 , n267465 , 
     n267466 , n267467 , n267468 , n267469 , n267470 , n267471 , n267472 , n267473 , n267474 , n267475 , 
     n267476 , n267477 , n267478 , n267479 , n267480 , n267481 , n267482 , n267483 , n267484 , n267485 , 
     n267486 , n267487 , n267488 , n267489 , n267490 , n267491 , n267492 , n267493 , n267494 , n267495 , 
     n267496 , n267497 , n267498 , n267499 , n267500 , n267501 , n267502 , n267503 , n267504 , n267505 , 
     n267506 , n267507 , n267508 , n267509 , n267510 , n267511 , n267512 , n267513 , n267514 , n267515 , 
     n267516 , n267517 , n267518 , n267519 , n267520 , n267521 , n267522 , n267523 , n267524 , n267525 , 
     n267526 , n267527 , n267528 , n267529 , n267530 , n267531 , n267532 , n267533 , n267534 , n267535 , 
     n267536 , n267537 , n267538 , n267539 , n267540 , n267541 , n267542 , n267543 , n267544 , n267545 , 
     n267546 , n267547 , n267548 , n267549 , n267550 , n267551 , n267552 , n267553 , n267554 , n267555 , 
     n267556 , n267557 , n267558 , n267559 , n267560 , n267561 , n267562 , n267563 , n267564 , n267565 , 
     n267566 , n267567 , n267568 , n267569 , n267570 , n267571 , n267572 , n267573 , n267574 , n267575 , 
     n267576 , n267577 , n267578 , n267579 , n267580 , n267581 , n267582 , n267583 , n267584 , n267585 , 
     n267586 , n267587 , n267588 , n267589 , n267590 , n267591 , n267592 , n267593 , n267594 , n267595 , 
     n267596 , n267597 , n267598 , n267599 , n267600 , n267601 , n267602 , n267603 , n267604 , n267605 , 
     n267606 , n267607 , n267608 , n267609 , n267610 , n267611 , n267612 , n267613 , n267614 , n267615 , 
     n267616 , n267617 , n267618 , n267619 , n267620 , n267621 , n267622 , n267623 , n267624 , n267625 , 
     n267626 , n267627 , n267628 , n267629 , n267630 , n267631 , n267632 , n267633 , n267634 , n267635 , 
     n267636 , n267637 , n267638 , n267639 , n267640 , n267641 , n267642 , n267643 , n267644 , n267645 , 
     n267646 , n267647 , n267648 , n267649 , n267650 , n267651 , n267652 , n267653 , n267654 , n267655 , 
     n267656 , n267657 , n267658 , n267659 , n267660 , n267661 , n267662 , n267663 , n267664 , n267665 , 
     n267666 , n267667 , n267668 , n267669 , n267670 , n267671 , n267672 , n267673 , n267674 , n267675 , 
     n267676 , n267677 , n267678 , n267679 , n267680 , n267681 , n267682 , n267683 , n267684 , n267685 , 
     n267686 , n267687 , n267688 , n267689 , n267690 , n267691 , n267692 , n267693 , n267694 , n267695 , 
     n267696 , n267697 , n267698 , n267699 , n267700 , n267701 , n267702 , n267703 , n267704 , n267705 , 
     n267706 , n267707 , n267708 , n267709 , n267710 , n267711 , n267712 , n267713 , n267714 , n267715 , 
     n267716 , n267717 , n267718 , n267719 , n267720 , n267721 , n267722 , n267723 , n267724 , n267725 , 
     n267726 , n267727 , n267728 , n267729 , n267730 , n267731 , n267732 , n267733 , n267734 , n267735 , 
     n267736 , n267737 , n267738 , n267739 , n267740 , n267741 , n267742 , n267743 , n267744 , n267745 , 
     n267746 , n267747 , n267748 , n267749 , n267750 , n267751 , n267752 , n267753 , n267754 , n267755 , 
     n267756 , n267757 , n267758 , n267759 , n267760 , n267761 , n267762 , n267763 , n267764 , n267765 , 
     n267766 , n267767 , n267768 , n267769 , n267770 , n267771 , n267772 , n267773 , n267774 , n267775 , 
     n267776 , n267777 , n267778 , n267779 , n267780 , n267781 , n267782 , n267783 , n267784 , n267785 , 
     n267786 , n267787 , n267788 , n267789 , n267790 , n267791 , n267792 , n267793 , n267794 , n267795 , 
     n267796 , n267797 , n267798 , n267799 , n267800 , n267801 , n267802 , n267803 , n267804 , n267805 , 
     n267806 , n267807 , n267808 , n267809 , n267810 , n267811 , n267812 , n267813 , n267814 , n267815 , 
     n267816 , n267817 , n267818 , n267819 , n267820 , n267821 , n267822 , n267823 , n267824 , n267825 , 
     n267826 , n267827 , n267828 , n267829 , n267830 , n267831 , n267832 , n267833 , n267834 , n267835 , 
     n267836 , n267837 , n267838 , n267839 , n267840 , n267841 , n267842 , n267843 , n267844 , n267845 , 
     n267846 , n267847 , n267848 , n267849 , n267850 , n267851 , n267852 , n267853 , n267854 , n267855 , 
     n267856 , n267857 , n267858 , n267859 , n267860 , n267861 , n267862 , n267863 , n267864 , n267865 , 
     n267866 , n267867 , n267868 , n267869 , n267870 , n267871 , n267872 , n267873 , n267874 , n267875 , 
     n267876 , n267877 , n267878 , n267879 , n267880 , n267881 , n267882 , n267883 , n267884 , n267885 , 
     n267886 , n267887 , n267888 , n267889 , n267890 , n267891 , n267892 , n267893 , n267894 , n267895 , 
     n267896 , n267897 , n267898 , n267899 , n267900 , n267901 , n267902 , n267903 , n267904 , n267905 , 
     n267906 , n267907 , n267908 , n267909 , n267910 , n267911 , n267912 , n267913 , n267914 , n267915 , 
     n267916 , n267917 , n267918 , n267919 , n267920 , n267921 , n267922 , n267923 , n267924 , n267925 , 
     n267926 , n267927 , n267928 , n267929 , n267930 , n267931 , n267932 , n267933 , n267934 , n267935 , 
     n267936 , n267937 , n267938 , n267939 , n267940 , n267941 , n267942 , n267943 , n267944 , n267945 , 
     n267946 , n267947 , n267948 , n267949 , n267950 , n267951 , n267952 , n267953 , n267954 , n267955 , 
     n267956 , n267957 , n267958 , n267959 , n267960 , n267961 , n267962 , n267963 , n267964 , n267965 , 
     n267966 , n267967 , n267968 , n267969 , n267970 , n267971 , n267972 , n267973 , n267974 , n267975 , 
     n267976 , n267977 , n267978 , n267979 , n267980 , n267981 , n267982 , n267983 , n267984 , n267985 , 
     n267986 , n267987 , n267988 , n267989 , n267990 , n267991 , n267992 , n267993 , n267994 , n267995 , 
     n267996 , n267997 , n267998 , n267999 , n268000 , n268001 , n268002 , n268003 , n268004 , n268005 , 
     n268006 , n268007 , n268008 , n268009 , n268010 , n268011 , n268012 , n268013 , n268014 , n268015 , 
     n268016 , n268017 , n268018 , n268019 , n268020 , n268021 , n268022 , n268023 , n268024 , n268025 , 
     n268026 , n268027 , n268028 , n268029 , n268030 , n268031 , n268032 , n268033 , n268034 , n268035 , 
     n268036 , n268037 , n268038 , n268039 , n268040 , n268041 , n268042 , n268043 , n268044 , n268045 , 
     n268046 , n268047 , n268048 , n268049 , n268050 , n268051 , n268052 , n268053 , n268054 , n268055 , 
     n268056 , n268057 , n268058 , n268059 , n268060 , n268061 , n268062 , n268063 , n268064 , n268065 , 
     n268066 , n268067 , n268068 , n268069 , n268070 , n268071 , n268072 , n268073 , n268074 , n268075 , 
     n268076 , n268077 , n268078 , n268079 , n268080 , n268081 , n268082 , n268083 , n268084 , n268085 , 
     n268086 , n268087 , n268088 , n268089 , n268090 , n268091 , n268092 , n268093 , n268094 , n268095 , 
     n268096 , n268097 , n268098 , n268099 , n268100 , n268101 , n268102 , n268103 , n268104 , n268105 , 
     n268106 , n268107 , n268108 , n268109 , n268110 , n268111 , n268112 , n268113 , n268114 , n268115 , 
     n268116 , n268117 , n268118 , n268119 , n268120 , n268121 , n268122 , n268123 , n268124 , n268125 , 
     n268126 , n268127 , n268128 , n268129 , n268130 , n268131 , n268132 , n268133 , n268134 , n268135 , 
     n268136 , n268137 , n268138 , n268139 , n268140 , n268141 , n268142 , n268143 , n268144 , n268145 , 
     n268146 , n268147 , n268148 , n268149 , n268150 , n268151 , n268152 , n268153 , n268154 , n268155 , 
     n268156 , n268157 , n268158 , n268159 , n268160 , n268161 , n268162 , n268163 , n268164 , n268165 , 
     n268166 , n268167 , n268168 , n268169 , n268170 , n268171 , n268172 , n268173 , n268174 , n268175 , 
     n268176 , n268177 , n268178 , n268179 , n268180 , n268181 , n268182 , n268183 , n268184 , n268185 , 
     n268186 , n268187 , n268188 , n268189 , n268190 , n268191 , n268192 , n268193 , n268194 , n268195 , 
     n268196 , n268197 , n268198 , n268199 , n268200 , n268201 , n268202 , n268203 , n268204 , n268205 , 
     n268206 , n268207 , n268208 , n268209 , n268210 , n268211 , n268212 , n268213 , n268214 , n268215 , 
     n268216 , n268217 , n268218 , n268219 , n268220 , n268221 , n268222 , n268223 , n268224 , n268225 , 
     n268226 , n268227 , n268228 , n268229 , n268230 , n268231 , n268232 , n268233 , n268234 , n268235 , 
     n268236 , n268237 , n268238 , n268239 , n268240 , n268241 , n268242 , n268243 , n268244 , n268245 , 
     n268246 , n268247 , n268248 , n268249 , n268250 , n268251 , n268252 , n268253 , n268254 , n268255 , 
     n268256 , n268257 , n268258 , n268259 , n268260 , n268261 , n268262 , n268263 , n268264 , n268265 , 
     n268266 , n268267 , n268268 , n268269 , n268270 , n268271 , n268272 , n268273 , n268274 , n268275 , 
     n268276 , n268277 , n268278 , n268279 , n268280 , n268281 , n268282 , n268283 , n268284 , n268285 , 
     n268286 , n268287 , n268288 , n268289 , n268290 , n268291 , n268292 , n268293 , n268294 , n268295 , 
     n268296 , n268297 , n268298 , n268299 , n268300 , n268301 , n268302 , n268303 , n268304 , n268305 , 
     n268306 , n268307 , n268308 , n268309 , n268310 , n268311 , n268312 , n268313 , n268314 , n268315 , 
     n268316 , n268317 , n268318 , n268319 , n268320 , n268321 , n268322 , n268323 , n268324 , n268325 , 
     n268326 , n268327 , n268328 , n268329 , n268330 , n268331 , n268332 , n268333 , n268334 , n268335 , 
     n268336 , n268337 , n268338 , n268339 , n268340 , n268341 , n268342 , n268343 , n268344 , n268345 , 
     n268346 , n268347 , n268348 , n268349 , n268350 , n268351 , n268352 , n268353 , n268354 , n268355 , 
     n268356 , n268357 , n268358 , n268359 , n268360 , n268361 , n268362 , n268363 , n268364 , n268365 , 
     n268366 , n268367 , n268368 , n268369 , n268370 , n268371 , n268372 , n268373 , n268374 , n268375 , 
     n268376 , n268377 , n268378 , n268379 , n268380 , n268381 , n268382 , n268383 , n268384 , n268385 , 
     n268386 , n268387 , n268388 , n268389 , n268390 , n268391 , n268392 , n268393 , n268394 , n268395 , 
     n268396 , n268397 , n268398 , n268399 , n268400 , n268401 , n268402 , n268403 , n268404 , n268405 , 
     n268406 , n268407 , n268408 , n268409 , n268410 , n268411 , n268412 , n268413 , n268414 , n268415 , 
     n268416 , n268417 , n268418 , n268419 , n268420 , n268421 , n268422 , n268423 , n268424 , n268425 , 
     n268426 , n268427 , n268428 , n268429 , n268430 , n268431 , n268432 , n268433 , n268434 , n268435 , 
     n268436 , n268437 , n268438 , n268439 , n268440 , n268441 , n268442 , n268443 , n268444 , n268445 , 
     n268446 , n268447 , n268448 , n268449 , n268450 , n268451 , n268452 , n268453 , n268454 , n268455 , 
     n268456 , n268457 , n268458 , n268459 , n268460 , n268461 , n268462 , n268463 , n268464 , n268465 , 
     n268466 , n268467 , n268468 , n268469 , n268470 , n268471 , n268472 , n268473 , n268474 , n268475 , 
     n268476 , n268477 , n268478 , n268479 , n268480 , n268481 , n268482 , n268483 , n268484 , n268485 , 
     n268486 , n268487 , n268488 , n268489 , n268490 , n268491 , n268492 , n268493 , n268494 , n268495 , 
     n268496 , n268497 , n268498 , n268499 , n268500 , n268501 , n268502 , n268503 , n268504 , n268505 , 
     n268506 , n268507 , n268508 , n268509 , n268510 , n268511 , n268512 , n268513 , n268514 , n268515 , 
     n268516 , n268517 , n268518 , n268519 , n268520 , n268521 , n268522 , n268523 , n268524 , n268525 , 
     n268526 , n268527 , n268528 , n268529 , n268530 , n268531 , n268532 , n268533 , n268534 , n268535 , 
     n268536 , n268537 , n268538 , n268539 , n268540 , n268541 , n268542 , n268543 , n268544 , n268545 , 
     n268546 , n268547 , n268548 , n268549 , n268550 , n268551 , n268552 , n268553 , n268554 , n268555 , 
     n268556 , n268557 , n268558 , n268559 , n268560 , n268561 , n268562 , n268563 , n268564 , n268565 , 
     n268566 , n268567 , n268568 , n268569 , n268570 , n268571 , n268572 , n268573 , n268574 , n268575 , 
     n268576 , n268577 , n268578 , n268579 , n268580 , n268581 , n268582 , n268583 , n268584 , n268585 , 
     n268586 , n268587 , n268588 , n268589 , n268590 , n268591 , n268592 , n268593 , n268594 , n268595 , 
     n268596 , n268597 , n268598 , n268599 , n268600 , n268601 , n268602 , n268603 , n268604 , n268605 , 
     n268606 , n268607 , n268608 , n268609 , n268610 , n268611 , n268612 , n268613 , n268614 , n268615 , 
     n268616 , n268617 , n268618 , n268619 , n268620 , n268621 , n268622 , n268623 , n268624 , n268625 , 
     n268626 , n268627 , n268628 , n268629 , n268630 , n268631 , n268632 , n268633 , n268634 , n268635 , 
     n268636 , n268637 , n268638 , n268639 , n268640 , n268641 , n268642 , n268643 , n268644 , n268645 , 
     n268646 , n268647 , n268648 , n268649 , n268650 , n268651 , n268652 , n268653 , n268654 , n268655 , 
     n268656 , n268657 , n268658 , n268659 , n268660 , n268661 , n268662 , n268663 , n268664 , n268665 , 
     n268666 , n268667 , n268668 , n268669 , n268670 , n268671 , n268672 , n268673 , n268674 , n268675 , 
     n268676 , n268677 , n268678 , n268679 , n268680 , n268681 , n268682 , n268683 , n268684 , n268685 , 
     n268686 , n268687 , n268688 , n268689 , n268690 , n268691 , n268692 , n268693 , n268694 , n268695 , 
     n268696 , n268697 , n268698 , n268699 , n268700 , n268701 , n268702 , n268703 , n268704 , n268705 , 
     n268706 , n268707 , n268708 , n268709 , n268710 , n268711 , n268712 , n268713 , n268714 , n268715 , 
     n268716 , n268717 , n268718 , n268719 , n268720 , n268721 , n268722 , n268723 , n268724 , n268725 , 
     n268726 , n268727 , n268728 , n268729 , n268730 , n268731 , n268732 , n268733 , n268734 , n268735 , 
     n268736 , n268737 , n268738 , n268739 , n268740 , n268741 , n268742 , n268743 , n268744 , n268745 , 
     n268746 , n268747 , n268748 , n268749 , n268750 , n268751 , n268752 , n268753 , n268754 , n268755 , 
     n268756 , n268757 , n268758 , n268759 , n268760 , n268761 , n268762 , n268763 , n268764 , n268765 , 
     n268766 , n268767 , n268768 , n268769 , n268770 , n268771 , n268772 , n268773 , n268774 , n268775 , 
     n268776 , n268777 , n268778 , n268779 , n268780 , n268781 , n268782 , n268783 , n268784 , n268785 , 
     n268786 , n268787 , n268788 , n268789 , n268790 , n268791 , n268792 , n268793 , n268794 , n268795 , 
     n268796 , n268797 , n268798 , n268799 , n268800 , n268801 , n268802 , n268803 , n268804 , n268805 , 
     n268806 , n268807 , n268808 , n268809 , n268810 , n268811 , n268812 , n268813 , n268814 , n268815 , 
     n268816 , n268817 , n268818 , n268819 , n268820 , n268821 , n268822 , n268823 , n268824 , n268825 , 
     n268826 , n268827 , n268828 , n268829 , n268830 , n268831 , n268832 , n268833 , n268834 , n268835 , 
     n268836 , n268837 , n268838 , n268839 , n268840 , n268841 , n268842 , n268843 , n268844 , n268845 , 
     n268846 , n268847 , n268848 , n268849 , n268850 , n268851 , n268852 , n268853 , n268854 , n268855 , 
     n268856 , n268857 , n268858 , n268859 , n268860 , n268861 , n268862 , n268863 , n268864 , n268865 , 
     n268866 , n268867 , n268868 , n268869 , n268870 , n268871 , n268872 , n268873 , n268874 , n268875 , 
     n268876 , n268877 , n268878 , n268879 , n268880 , n268881 , n268882 , n268883 , n268884 , n268885 , 
     n268886 , n268887 , n268888 , n268889 , n268890 , n268891 , n268892 , n268893 , n268894 , n268895 , 
     n268896 , n268897 , n268898 , n268899 , n268900 , n268901 , n268902 , n268903 , n268904 , n268905 , 
     n268906 , n268907 , n268908 , n268909 , n268910 , n268911 , n268912 , n268913 , n268914 , n268915 , 
     n268916 , n268917 , n268918 , n268919 , n268920 , n268921 , n268922 , n268923 , n268924 , n268925 , 
     n268926 , n268927 , n268928 , n268929 , n268930 , n268931 , n268932 , n268933 , n268934 , n268935 , 
     n268936 , n268937 , n268938 , n268939 , n268940 , n268941 , n268942 , n268943 , n268944 , n268945 , 
     n268946 , n268947 , n268948 , n268949 , n268950 , n268951 , n268952 , n268953 , n268954 , n268955 , 
     n268956 , n268957 , n268958 , n268959 , n268960 , n268961 , n268962 , n268963 , n268964 , n268965 , 
     n268966 , n268967 , n268968 , n268969 , n268970 , n268971 , n268972 , n268973 , n268974 , n268975 , 
     n268976 , n268977 , n268978 , n268979 , n268980 , n268981 , n268982 , n268983 , n268984 , n268985 , 
     n268986 , n268987 , n268988 , n268989 , n268990 , n268991 , n268992 , n268993 , n268994 , n268995 , 
     n268996 , n268997 , n268998 , n268999 , n269000 , n269001 , n269002 , n269003 , n269004 , n269005 , 
     n269006 , n269007 , n269008 , n269009 , n269010 , n269011 , n269012 , n269013 , n269014 , n269015 , 
     n269016 , n269017 , n269018 , n269019 , n269020 , n269021 , n269022 , n269023 , n269024 , n269025 , 
     n269026 , n269027 , n269028 , n269029 , n269030 , n269031 , n269032 , n269033 , n269034 , n269035 , 
     n269036 , n269037 , n269038 , n269039 , n269040 , n269041 , n269042 , n269043 , n269044 , n269045 , 
     n269046 , n269047 , n269048 , n269049 , n269050 , n269051 , n269052 , n269053 , n269054 , n269055 , 
     n269056 , n269057 , n269058 , n269059 , n269060 , n269061 , n269062 , n269063 , n269064 , n269065 , 
     n269066 , n269067 , n269068 , n269069 , n269070 , n269071 , n269072 , n269073 , n269074 , n269075 , 
     n269076 , n269077 , n269078 , n269079 , n269080 , n269081 , n269082 , n269083 , n269084 , n269085 , 
     n269086 , n269087 , n269088 , n269089 , n269090 , n269091 , n269092 , n269093 , n269094 , n269095 , 
     n269096 , n269097 , n269098 , n269099 , n269100 , n269101 , n269102 , n269103 , n269104 , n269105 , 
     n269106 , n269107 , n269108 , n269109 , n269110 , n269111 , n269112 , n269113 , n269114 , n269115 , 
     n269116 , n269117 , n269118 , n269119 , n269120 , n269121 , n269122 , n269123 , n269124 , n269125 , 
     n269126 , n269127 , n269128 , n269129 , n269130 , n269131 , n269132 , n269133 , n269134 , n269135 , 
     n269136 , n269137 , n269138 , n269139 , n269140 , n269141 , n269142 , n269143 , n269144 , n269145 , 
     n269146 , n269147 , n269148 , n269149 , n269150 , n269151 , n269152 , n269153 , n269154 , n269155 , 
     n269156 , n269157 , n269158 , n269159 , n269160 , n269161 , n269162 , n269163 , n269164 , n269165 , 
     n269166 , n269167 , n269168 , n269169 , n269170 , n269171 , n269172 , n269173 , n269174 , n269175 , 
     n269176 , n269177 , n269178 , n269179 , n269180 , n269181 , n269182 , n269183 , n269184 , n269185 , 
     n269186 , n269187 , n269188 , n269189 , n269190 , n269191 , n269192 , n269193 , n269194 , n269195 , 
     n269196 , n269197 , n269198 , n269199 , n269200 , n269201 , n269202 , n269203 , n269204 , n269205 , 
     n269206 , n269207 , n269208 , n269209 , n269210 , n269211 , n269212 , n269213 , n269214 , n269215 , 
     n269216 , n269217 , n269218 , n269219 , n269220 , n269221 , n269222 , n269223 , n269224 , n269225 , 
     n269226 , n269227 , n269228 , n269229 , n269230 , n269231 , n269232 , n269233 , n269234 , n269235 , 
     n269236 , n269237 , n269238 , n269239 , n269240 , n269241 , n269242 , n269243 , n269244 , n269245 , 
     n269246 , n269247 , n269248 , n269249 , n269250 , n269251 , n269252 , n269253 , n269254 , n269255 , 
     n269256 , n269257 , n269258 , n269259 , n269260 , n269261 , n269262 , n269263 , n269264 , n269265 , 
     n269266 , n269267 , n269268 , n269269 , n269270 , n269271 , n269272 , n269273 , n269274 , n269275 , 
     n269276 , n269277 , n269278 , n269279 , n269280 , n269281 , n269282 , n269283 , n269284 , n269285 , 
     n269286 , n269287 , n269288 , n269289 , n269290 , n269291 , n269292 , n269293 , n269294 , n269295 , 
     n269296 , n269297 , n269298 , n269299 , n269300 , n269301 , n269302 , n269303 , n269304 , n269305 , 
     n269306 , n269307 , n269308 , n269309 , n269310 , n269311 , n269312 , n269313 , n269314 , n269315 , 
     n269316 , n269317 , n269318 , n269319 , n269320 , n269321 , n269322 , n269323 , n269324 , n269325 , 
     n269326 , n269327 , n269328 , n269329 , n269330 , n269331 , n269332 , n269333 , n269334 , n269335 , 
     n269336 , n269337 , n269338 , n269339 , n269340 , n269341 , n269342 , n269343 , n269344 , n269345 , 
     n269346 , n269347 , n269348 , n269349 , n269350 , n269351 , n269352 , n269353 , n269354 , n269355 , 
     n269356 , n269357 , n269358 , n269359 , n269360 , n269361 , n269362 , n269363 , n269364 , n269365 , 
     n269366 , n269367 , n269368 , n269369 , n269370 , n269371 , n269372 , n269373 , n269374 , n269375 , 
     n269376 , n269377 , n269378 , n269379 , n269380 , n269381 , n269382 , n269383 , n269384 , n269385 , 
     n269386 , n269387 , n269388 , n269389 , n269390 , n269391 , n269392 , n269393 , n269394 , n269395 , 
     n269396 , n269397 , n269398 , n269399 , n269400 , n269401 , n269402 , n269403 , n269404 , n269405 , 
     n269406 , n269407 , n269408 , n269409 , n269410 , n269411 , n269412 , n269413 , n269414 , n269415 , 
     n269416 , n269417 , n269418 , n269419 , n269420 , n269421 , n269422 , n269423 , n269424 , n269425 , 
     n269426 , n269427 , n269428 , n269429 , n269430 , n269431 , n269432 , n269433 , n269434 , n269435 , 
     n269436 , n269437 , n269438 , n269439 , n269440 , n269441 , n269442 , n269443 , n269444 , n269445 , 
     n269446 , n269447 , n269448 , n269449 , n269450 , n269451 , n269452 , n269453 , n269454 , n269455 , 
     n269456 , n269457 , n269458 , n269459 , n269460 , n269461 , n269462 , n269463 , n269464 , n269465 , 
     n269466 , n269467 , n269468 , n269469 , n269470 , n269471 , n269472 , n269473 , n269474 , n269475 , 
     n269476 , n269477 , n269478 , n269479 , n269480 , n269481 , n269482 , n269483 , n269484 , n269485 , 
     n269486 , n269487 , n269488 , n269489 , n269490 , n269491 , n269492 , n269493 , n269494 , n269495 , 
     n269496 , n269497 , n269498 , n269499 , n269500 , n269501 , n269502 , n269503 , n269504 , n269505 , 
     n269506 , n269507 , n269508 , n269509 , n269510 , n269511 , n269512 , n269513 , n269514 , n269515 , 
     n269516 , n269517 , n269518 , n269519 , n269520 , n269521 , n269522 , n269523 , n269524 , n269525 , 
     n269526 , n269527 , n269528 , n269529 , n269530 , n269531 , n269532 , n269533 , n269534 , n269535 , 
     n269536 , n269537 , n269538 , n269539 , n269540 , n269541 , n269542 , n269543 , n269544 , n269545 , 
     n269546 , n269547 , n269548 , n269549 , n269550 , n269551 , n269552 , n269553 , n269554 , n269555 , 
     n269556 , n269557 , n269558 , n269559 , n269560 , n269561 , n269562 , n269563 , n269564 , n269565 , 
     n269566 , n269567 , n269568 , n269569 , n269570 , n269571 , n269572 , n269573 , n269574 , n269575 , 
     n269576 , n269577 , n269578 , n269579 , n269580 , n269581 , n269582 , n269583 , n269584 , n269585 , 
     n269586 , n269587 , n269588 , n269589 , n269590 , n269591 , n269592 , n269593 , n269594 , n269595 , 
     n269596 , n269597 , n269598 , n269599 , n269600 , n269601 , n269602 , n269603 , n269604 , n269605 , 
     n269606 , n269607 , n269608 , n269609 , n269610 , n269611 , n269612 , n269613 , n269614 , n269615 , 
     n269616 , n269617 , n269618 , n269619 , n269620 , n269621 , n269622 , n269623 , n269624 , n269625 , 
     n269626 , n269627 , n269628 , n269629 , n269630 , n269631 , n269632 , n269633 , n269634 , n269635 , 
     n269636 , n269637 , n269638 , n269639 , n269640 , n269641 , n269642 , n269643 , n269644 , n269645 , 
     n269646 , n269647 , n269648 , n269649 , n269650 , n269651 , n269652 , n269653 , n269654 , n269655 , 
     n269656 , n269657 , n269658 , n269659 , n269660 , n269661 , n269662 , n269663 , n269664 , n269665 , 
     n269666 , n269667 , n269668 , n269669 , n269670 , n269671 , n269672 , n269673 , n269674 , n269675 , 
     n269676 , n269677 , n269678 , n269679 , n269680 , n269681 , n269682 , n269683 , n269684 , n269685 , 
     n269686 , n269687 , n269688 , n269689 , n269690 , n269691 , n269692 , n269693 , n269694 , n269695 , 
     n269696 , n269697 , n269698 , n269699 , n269700 , n269701 , n269702 , n269703 , n269704 , n269705 , 
     n269706 , n269707 , n269708 , n269709 , n269710 , n269711 , n269712 , n269713 , n269714 , n269715 , 
     n269716 , n269717 , n269718 , n269719 , n269720 , n269721 , n269722 , n269723 , n269724 , n269725 , 
     n269726 , n269727 , n269728 , n269729 , n269730 , n269731 , n269732 , n269733 , n269734 , n269735 , 
     n269736 , n269737 , n269738 , n269739 , n269740 , n269741 , n269742 , n269743 , n269744 , n269745 , 
     n269746 , n269747 , n269748 , n269749 , n269750 , n269751 , n269752 , n269753 , n269754 , n269755 , 
     n269756 , n269757 , n269758 , n269759 , n269760 , n269761 , n269762 , n269763 , n269764 , n269765 , 
     n269766 , n269767 , n269768 , n269769 , n269770 , n269771 , n269772 , n269773 , n269774 , n269775 , 
     n269776 , n269777 , n269778 , n269779 , n269780 , n269781 , n269782 , n269783 , n269784 , n269785 , 
     n269786 , n269787 , n269788 , n269789 , n269790 , n269791 , n269792 , n269793 , n269794 , n269795 , 
     n269796 , n269797 , n269798 , n269799 , n269800 , n269801 , n269802 , n269803 , n269804 , n269805 , 
     n269806 , n269807 , n269808 , n269809 , n269810 , n269811 , n269812 , n269813 , n269814 , n269815 , 
     n269816 , n269817 , n269818 , n269819 , n269820 , n269821 , n269822 , n269823 , n269824 , n269825 , 
     n269826 , n269827 , n269828 , n269829 , n269830 , n269831 , n269832 , n269833 , n269834 , n269835 , 
     n269836 , n269837 , n269838 , n269839 , n269840 , n269841 , n269842 , n269843 , n269844 , n269845 , 
     n269846 , n269847 , n269848 , n269849 , n269850 , n269851 , n269852 , n269853 , n269854 , n269855 , 
     n269856 , n269857 , n269858 , n269859 , n269860 , n269861 , n269862 , n269863 , n269864 , n269865 , 
     n269866 , n269867 , n269868 , n269869 , n269870 , n269871 , n269872 , n269873 , n269874 , n269875 , 
     n269876 , n269877 , n269878 , n269879 , n269880 , n269881 , n269882 , n269883 , n269884 , n269885 , 
     n269886 , n269887 , n269888 , n269889 , n269890 , n269891 , n269892 , n269893 , n269894 , n269895 , 
     n269896 , n269897 , n269898 , n269899 , n269900 , n269901 , n269902 , n269903 , n269904 , n269905 , 
     n269906 , n269907 , n269908 , n269909 , n269910 , n269911 , n269912 , n269913 , n269914 , n269915 , 
     n269916 , n269917 , n269918 , n269919 , n269920 , n269921 , n269922 , n269923 , n269924 , n269925 , 
     n269926 , n269927 , n269928 , n269929 , n269930 , n269931 , n269932 , n269933 , n269934 , n269935 , 
     n269936 , n269937 , n269938 , n269939 , n269940 , n269941 , n269942 , n269943 , n269944 , n269945 , 
     n269946 , n269947 , n269948 , n269949 , n269950 , n269951 , n269952 , n269953 , n269954 , n269955 , 
     n269956 , n269957 , n269958 , n269959 , n269960 , n269961 , n269962 , n269963 , n269964 , n269965 , 
     n269966 , n269967 , n269968 , n269969 , n269970 , n269971 , n269972 , n269973 , n269974 , n269975 , 
     n269976 , n269977 , n269978 , n269979 , n269980 , n269981 , n269982 , n269983 , n269984 , n269985 , 
     n269986 , n269987 , n269988 , n269989 , n269990 , n269991 , n269992 , n269993 , n269994 , n269995 , 
     n269996 , n269997 , n269998 , n269999 , n270000 , n270001 , n270002 , n270003 , n270004 , n270005 , 
     n270006 , n270007 , n270008 , n270009 , n270010 , n270011 , n270012 , n270013 , n270014 , n270015 , 
     n270016 , n270017 , n270018 , n270019 , n270020 , n270021 , n270022 , n270023 , n270024 , n270025 , 
     n270026 , n270027 , n270028 , n270029 , n270030 , n270031 , n270032 , n270033 , n270034 , n270035 , 
     n270036 , n270037 , n270038 , n270039 , n270040 , n270041 , n270042 , n270043 , n270044 , n270045 , 
     n270046 , n270047 , n270048 , n270049 , n270050 , n270051 , n270052 , n270053 , n270054 , n270055 , 
     n270056 , n270057 , n270058 , n270059 , n270060 , n270061 , n270062 , n270063 , n270064 , n270065 , 
     n270066 , n270067 , n270068 , n270069 , n270070 , n270071 , n270072 , n270073 , n270074 , n270075 , 
     n270076 , n270077 , n270078 , n270079 , n270080 , n270081 , n270082 , n270083 , n270084 , n270085 , 
     n270086 , n270087 , n270088 , n270089 , n270090 , n270091 , n270092 , n270093 , n270094 , n270095 , 
     n270096 , n270097 , n270098 , n270099 , n270100 , n270101 , n270102 , n270103 , n270104 , n270105 , 
     n270106 , n270107 , n270108 , n270109 , n270110 , n270111 , n270112 , n270113 , n270114 , n270115 , 
     n270116 , n270117 , n270118 , n270119 , n270120 , n270121 , n270122 , n270123 , n270124 , n270125 , 
     n270126 , n270127 , n270128 , n270129 , n270130 , n270131 , n270132 , n270133 , n270134 , n270135 , 
     n270136 , n270137 , n270138 , n270139 , n270140 , n270141 , n270142 , n270143 , n270144 , n270145 , 
     n270146 , n270147 , n270148 , n270149 , n270150 , n270151 , n270152 , n270153 , n270154 , n270155 , 
     n270156 , n270157 , n270158 , n270159 , n270160 , n270161 , n270162 , n270163 , n270164 , n270165 , 
     n270166 , n270167 , n270168 , n270169 , n270170 , n270171 , n270172 , n270173 , n270174 , n270175 , 
     n270176 , n270177 , n270178 , n270179 , n270180 , n270181 , n270182 , n270183 , n270184 , n270185 , 
     n270186 , n270187 , n270188 , n270189 , n270190 , n270191 , n270192 , n270193 , n270194 , n270195 , 
     n270196 , n270197 , n270198 , n270199 , n270200 , n270201 , n270202 , n270203 , n270204 , n270205 , 
     n270206 , n270207 , n270208 , n270209 , n270210 , n270211 , n270212 , n270213 , n270214 , n270215 , 
     n270216 , n270217 , n270218 , n270219 , n270220 , n270221 , n270222 , n270223 , n270224 , n270225 , 
     n270226 , n270227 , n270228 , n270229 , n270230 , n270231 , n270232 , n270233 , n270234 , n270235 , 
     n270236 , n270237 , n270238 , n270239 , n270240 , n270241 , n270242 , n270243 , n270244 , n270245 , 
     n270246 , n270247 , n270248 , n270249 , n270250 , n270251 , n270252 , n270253 , n270254 , n270255 , 
     n270256 , n270257 , n270258 , n270259 , n270260 , n270261 , n270262 , n270263 , n270264 , n270265 , 
     n270266 , n270267 , n270268 , n270269 , n270270 , n270271 , n270272 , n270273 , n270274 , n270275 , 
     n270276 , n270277 , n270278 , n270279 , n270280 , n270281 , n270282 , n270283 , n270284 , n270285 , 
     n270286 , n270287 , n270288 , n270289 , n270290 , n270291 , n270292 , n270293 , n270294 , n270295 , 
     n270296 , n270297 , n270298 , n270299 , n270300 , n270301 , n270302 , n270303 , n270304 , n270305 , 
     n270306 , n270307 , n270308 , n270309 , n270310 , n270311 , n270312 , n270313 , n270314 , n270315 , 
     n270316 , n270317 , n270318 , n270319 , n270320 , n270321 , n270322 , n270323 , n270324 , n270325 , 
     n270326 , n270327 , n270328 , n270329 , n270330 , n270331 , n270332 , n270333 , n270334 , n270335 , 
     n270336 , n270337 , n270338 , n270339 , n270340 , n270341 , n270342 , n270343 , n270344 , n270345 , 
     n270346 , n270347 , n270348 , n270349 , n270350 , n270351 , n270352 , n270353 , n270354 , n270355 , 
     n270356 , n270357 , n270358 , n270359 , n270360 , n270361 , n270362 , n270363 , n270364 , n270365 , 
     n270366 , n270367 , n270368 , n270369 , n270370 , n270371 , n270372 , n270373 , n270374 , n270375 , 
     n270376 , n270377 , n270378 , n270379 , n270380 , n270381 , n270382 , n270383 , n270384 , n270385 , 
     n270386 , n270387 , n270388 , n270389 , n270390 , n270391 , n270392 , n270393 , n270394 , n270395 , 
     n270396 , n270397 , n270398 , n270399 , n270400 , n270401 , n270402 , n270403 , n270404 , n270405 , 
     n270406 , n270407 , n270408 , n270409 , n270410 , n270411 , n270412 , n270413 , n270414 , n270415 , 
     n270416 , n270417 , n270418 , n270419 , n270420 , n270421 , n270422 , n270423 , n270424 , n270425 , 
     n270426 , n270427 , n270428 , n270429 , n270430 , n270431 , n270432 , n270433 , n270434 , n270435 , 
     n270436 , n270437 , n270438 , n270439 , n270440 , n270441 , n270442 , n270443 , n270444 , n270445 , 
     n270446 , n270447 , n270448 , n270449 , n270450 , n270451 , n270452 , n270453 , n270454 , n270455 , 
     n270456 , n270457 , n270458 , n270459 , n270460 , n270461 , n270462 , n270463 , n270464 , n270465 , 
     n270466 , n270467 , n270468 , n270469 , n270470 , n270471 , n270472 , n270473 , n270474 , n270475 , 
     n270476 , n270477 , n270478 , n270479 , n270480 , n270481 , n270482 , n270483 , n270484 , n270485 , 
     n270486 , n270487 , n270488 , n270489 , n270490 , n270491 , n270492 , n270493 , n270494 , n270495 , 
     n270496 , n270497 , n270498 , n270499 , n270500 , n270501 , n270502 , n270503 , n270504 , n270505 , 
     n270506 , n270507 , n270508 , n270509 , n270510 , n270511 , n270512 , n270513 , n270514 , n270515 , 
     n270516 , n270517 , n270518 , n270519 , n270520 , n270521 , n270522 , n270523 , n270524 , n270525 , 
     n270526 , n270527 , n270528 , n270529 , n270530 , n270531 , n270532 , n270533 , n270534 , n270535 , 
     n270536 , n270537 , n270538 , n270539 , n270540 , n270541 , n270542 , n270543 , n270544 , n270545 , 
     n270546 , n270547 , n270548 , n270549 , n270550 , n270551 , n270552 , n270553 , n270554 , n270555 , 
     n270556 , n270557 , n270558 , n270559 , n270560 , n270561 , n270562 , n270563 , n270564 , n270565 , 
     n270566 , n270567 , n270568 , n270569 , n270570 , n270571 , n270572 , n270573 , n270574 , n270575 , 
     n270576 , n270577 , n270578 , n270579 , n270580 , n270581 , n270582 , n270583 , n270584 , n270585 , 
     n270586 , n270587 , n270588 , n270589 , n270590 , n270591 , n270592 , n270593 , n270594 , n270595 , 
     n270596 , n270597 , n270598 , n270599 , n270600 , n270601 , n270602 , n270603 , n270604 , n270605 , 
     n270606 , n270607 , n270608 , n270609 , n270610 , n270611 , n270612 , n270613 , n270614 , n270615 , 
     n270616 , n270617 , n270618 , n270619 , n270620 , n270621 , n270622 , n270623 , n270624 , n270625 , 
     n270626 , n270627 , n270628 , n270629 , n270630 , n270631 , n270632 , n270633 , n270634 , n270635 , 
     n270636 , n270637 , n270638 , n270639 , n270640 , n270641 , n270642 , n270643 , n270644 , n270645 , 
     n270646 , n270647 , n270648 , n270649 , n270650 , n270651 , n270652 , n270653 , n270654 , n270655 , 
     n270656 , n270657 , n270658 , n270659 , n270660 , n270661 , n270662 , n270663 , n270664 , n270665 , 
     n270666 , n270667 , n270668 , n270669 , n270670 , n270671 , n270672 , n270673 , n270674 , n270675 , 
     n270676 , n270677 , n270678 , n270679 , n270680 , n270681 , n270682 , n270683 , n270684 , n270685 , 
     n270686 , n270687 , n270688 , n270689 , n270690 , n270691 , n270692 , n270693 , n270694 , n270695 , 
     n270696 , n270697 , n270698 , n270699 , n270700 , n270701 , n270702 , n270703 , n270704 , n270705 , 
     n270706 , n270707 , n270708 , n270709 , n270710 , n270711 , n270712 , n270713 , n270714 , n270715 , 
     n270716 , n270717 , n270718 , n270719 , n270720 , n270721 , n270722 , n270723 , n270724 , n270725 , 
     n270726 , n270727 , n270728 , n270729 , n270730 , n270731 , n270732 , n270733 , n270734 , n270735 , 
     n270736 , n270737 , n270738 , n270739 , n270740 , n270741 , n270742 , n270743 , n270744 , n270745 , 
     n270746 , n270747 , n270748 , n270749 , n270750 , n270751 , n270752 , n270753 , n270754 , n270755 , 
     n270756 , n270757 , n270758 , n270759 , n270760 , n270761 , n270762 , n270763 , n270764 , n270765 , 
     n270766 , n270767 , n270768 , n270769 , n270770 , n270771 , n270772 , n270773 , n270774 , n270775 , 
     n270776 , n270777 , n270778 , n270779 , n270780 , n270781 , n270782 , n270783 , n270784 , n270785 , 
     n270786 , n270787 , n270788 , n270789 , n270790 , n270791 , n270792 , n270793 , n270794 , n270795 , 
     n270796 , n270797 , n270798 , n270799 , n270800 , n270801 , n270802 , n270803 , n270804 , n270805 , 
     n270806 , n270807 , n270808 , n270809 , n270810 , n270811 , n270812 , n270813 , n270814 , n270815 , 
     n270816 , n270817 , n270818 , n270819 , n270820 , n270821 , n270822 , n270823 , n270824 , n270825 , 
     n270826 , n270827 , n270828 , n270829 , n270830 , n270831 , n270832 , n270833 , n270834 , n270835 , 
     n270836 , n270837 , n270838 , n270839 , n270840 , n270841 , n270842 , n270843 , n270844 , n270845 , 
     n270846 , n270847 , n270848 , n270849 , n270850 , n270851 , n270852 , n270853 , n270854 , n270855 , 
     n270856 , n270857 , n270858 , n270859 , n270860 , n270861 , n270862 , n270863 , n270864 , n270865 , 
     n270866 , n270867 , n270868 , n270869 , n270870 , n270871 , n270872 , n270873 , n270874 , n270875 , 
     n270876 , n270877 , n270878 , n270879 , n270880 , n270881 , n270882 , n270883 , n270884 , n270885 , 
     n270886 , n270887 , n270888 , n270889 , n270890 , n270891 , n270892 , n270893 , n270894 , n270895 , 
     n270896 , n270897 , n270898 , n270899 , n270900 , n270901 , n270902 , n270903 , n270904 , n270905 , 
     n270906 , n270907 , n270908 , n270909 , n270910 , n270911 , n270912 , n270913 , n270914 , n270915 , 
     n270916 , n270917 , n270918 , n270919 , n270920 , n270921 , n270922 , n270923 , n270924 , n270925 , 
     n270926 , n270927 , n270928 , n270929 , n270930 , n270931 , n270932 , n270933 , n270934 , n270935 , 
     n270936 , n270937 , n270938 , n270939 , n270940 , n270941 , n270942 , n270943 , n270944 , n270945 , 
     n270946 , n270947 , n270948 , n270949 , n270950 , n270951 , n270952 , n270953 , n270954 , n270955 , 
     n270956 , n270957 , n270958 , n270959 , n270960 , n270961 , n270962 , n270963 , n270964 , n270965 , 
     n270966 , n270967 , n270968 , n270969 , n270970 , n270971 , n270972 , n270973 , n270974 , n270975 , 
     n270976 , n270977 , n270978 , n270979 , n270980 , n270981 , n270982 , n270983 , n270984 , n270985 , 
     n270986 , n270987 , n270988 , n270989 , n270990 , n270991 , n270992 , n270993 , n270994 , n270995 , 
     n270996 , n270997 , n270998 , n270999 , n271000 , n271001 , n271002 , n271003 , n271004 , n271005 , 
     n271006 , n271007 , n271008 , n271009 , n271010 , n271011 , n271012 , n271013 , n271014 , n271015 , 
     n271016 , n271017 , n271018 , n271019 , n271020 , n271021 , n271022 , n271023 , n271024 , n271025 , 
     n271026 , n271027 , n271028 , n271029 , n271030 , n271031 , n271032 , n271033 , n271034 , n271035 , 
     n271036 , n271037 , n271038 , n271039 , n271040 , n271041 , n271042 , n271043 , n271044 , n271045 , 
     n271046 , n271047 , n271048 , n271049 , n271050 , n271051 , n271052 , n271053 , n271054 , n271055 , 
     n271056 , n271057 , n271058 , n271059 , n271060 , n271061 , n271062 , n271063 , n271064 , n271065 , 
     n271066 , n271067 , n271068 , n271069 , n271070 , n271071 , n271072 , n271073 , n271074 , n271075 , 
     n271076 , n271077 , n271078 , n271079 , n271080 , n271081 , n271082 , n271083 , n271084 , n271085 , 
     n271086 , n271087 , n271088 , n271089 , n271090 , n271091 , n271092 , n271093 , n271094 , n271095 , 
     n271096 , n271097 , n271098 , n271099 , n271100 , n271101 , n271102 , n271103 , n271104 , n271105 , 
     n271106 , n271107 , n271108 , n271109 , n271110 , n271111 , n271112 , n271113 , n271114 , n271115 , 
     n271116 , n271117 , n271118 , n271119 , n271120 , n271121 , n271122 , n271123 , n271124 , n271125 , 
     n271126 , n271127 , n271128 , n271129 , n271130 , n271131 , n271132 , n271133 , n271134 , n271135 , 
     n271136 , n271137 , n271138 , n271139 , n271140 , n271141 , n271142 , n271143 , n271144 , n271145 , 
     n271146 , n271147 , n271148 , n271149 , n271150 , n271151 , n271152 , n271153 , n271154 , n271155 , 
     n271156 , n271157 , n271158 , n271159 , n271160 , n271161 , n271162 , n271163 , n271164 , n271165 , 
     n271166 , n271167 , n271168 , n271169 , n271170 , n271171 , n271172 , n271173 , n271174 , n271175 , 
     n271176 , n271177 , n271178 , n271179 , n271180 , n271181 , n271182 , n271183 , n271184 , n271185 , 
     n271186 , n271187 , n271188 , n271189 , n271190 , n271191 , n271192 , n271193 , n271194 , n271195 , 
     n271196 , n271197 , n271198 , n271199 , n271200 , n271201 , n271202 , n271203 , n271204 , n271205 , 
     n271206 , n271207 , n271208 , n271209 , n271210 , n271211 , n271212 , n271213 , n271214 , n271215 , 
     n271216 , n271217 , n271218 , n271219 , n271220 , n271221 , n271222 , n271223 , n271224 , n271225 , 
     n271226 , n271227 , n271228 , n271229 , n271230 , n271231 , n271232 , n271233 , n271234 , n271235 , 
     n271236 , n271237 , n271238 , n271239 , n271240 , n271241 , n271242 , n271243 , n271244 , n271245 , 
     n271246 , n271247 , n271248 , n271249 , n271250 , n271251 , n271252 , n271253 , n271254 , n271255 , 
     n271256 , n271257 , n271258 , n271259 , n271260 , n271261 , n271262 , n271263 , n271264 , n271265 , 
     n271266 , n271267 , n271268 , n271269 , n271270 , n271271 , n271272 , n271273 , n271274 , n271275 , 
     n271276 , n271277 , n271278 , n271279 , n271280 , n271281 , n271282 , n271283 , n271284 , n271285 , 
     n271286 , n271287 , n271288 , n271289 , n271290 , n271291 , n271292 , n271293 , n271294 , n271295 , 
     n271296 , n271297 , n271298 , n271299 , n271300 , n271301 , n271302 , n271303 , n271304 , n271305 , 
     n271306 , n271307 , n271308 , n271309 , n271310 , n271311 , n271312 , n271313 , n271314 , n271315 , 
     n271316 , n271317 , n271318 , n271319 , n271320 , n271321 , n271322 , n271323 , n271324 , n271325 , 
     n271326 , n271327 , n271328 , n271329 , n271330 , n271331 , n271332 , n271333 , n271334 , n271335 , 
     n271336 , n271337 , n271338 , n271339 , n271340 , n271341 , n271342 , n271343 , n271344 , n271345 , 
     n271346 , n271347 , n271348 , n271349 , n271350 , n271351 , n271352 , n271353 , n271354 , n271355 , 
     n271356 , n271357 , n271358 , n271359 , n271360 , n271361 , n271362 , n271363 , n271364 , n271365 , 
     n271366 , n271367 , n271368 , n271369 , n271370 , n271371 , n271372 , n271373 , n271374 , n271375 , 
     n271376 , n271377 , n271378 , n271379 , n271380 , n271381 , n271382 , n271383 , n271384 , n271385 , 
     n271386 , n271387 , n271388 , n271389 , n271390 , n271391 , n271392 , n271393 , n271394 , n271395 , 
     n271396 , n271397 , n271398 , n271399 , n271400 , n271401 , n271402 , n271403 , n271404 , n271405 , 
     n271406 , n271407 , n271408 , n271409 , n271410 , n271411 , n271412 , n271413 , n271414 , n271415 , 
     n271416 , n271417 , n271418 , n271419 , n271420 , n271421 , n271422 , n271423 , n271424 , n271425 , 
     n271426 , n271427 , n271428 , n271429 , n271430 , n271431 , n271432 , n271433 , n271434 , n271435 , 
     n271436 , n271437 , n271438 , n271439 , n271440 , n271441 , n271442 , n271443 , n271444 , n271445 , 
     n271446 , n271447 , n271448 , n271449 , n271450 , n271451 , n271452 , n271453 , n271454 , n271455 , 
     n271456 , n271457 , n271458 , n271459 , n271460 , n271461 , n271462 , n271463 , n271464 , n271465 , 
     n271466 , n271467 , n271468 , n271469 , n271470 , n271471 , n271472 , n271473 , n271474 , n271475 , 
     n271476 , n271477 , n271478 , n271479 , n271480 , n271481 , n271482 , n271483 , n271484 , n271485 , 
     n271486 , n271487 , n271488 , n271489 , n271490 , n271491 , n271492 , n271493 , n271494 , n271495 , 
     n271496 , n271497 , n271498 , n271499 , n271500 , n271501 , n271502 , n271503 , n271504 , n271505 , 
     n271506 , n271507 , n271508 , n271509 , n271510 , n271511 , n271512 , n271513 , n271514 , n271515 , 
     n271516 , n271517 , n271518 , n271519 , n271520 , n271521 , n271522 , n271523 , n271524 , n271525 , 
     n271526 , n271527 , n271528 , n271529 , n271530 , n271531 , n271532 , n271533 , n271534 , n271535 , 
     n271536 , n271537 , n271538 , n271539 , n271540 , n271541 , n271542 , n271543 , n271544 , n271545 , 
     n271546 , n271547 , n271548 , n271549 , n271550 , n271551 , n271552 , n271553 , n271554 , n271555 , 
     n271556 , n271557 , n271558 , n271559 , n271560 , n271561 , n271562 , n271563 , n271564 , n271565 , 
     n271566 , n271567 , n271568 , n271569 , n271570 , n271571 , n271572 , n271573 , n271574 , n271575 , 
     n271576 , n271577 , n271578 , n271579 , n271580 , n271581 , n271582 , n271583 , n271584 , n271585 , 
     n271586 , n271587 , n271588 , n271589 , n271590 , n271591 , n271592 , n271593 , n271594 , n271595 , 
     n271596 , n271597 , n271598 , n271599 , n271600 , n271601 , n271602 , n271603 , n271604 , n271605 , 
     n271606 , n271607 , n271608 , n271609 , n271610 , n271611 , n271612 , n271613 , n271614 , n271615 , 
     n271616 , n271617 , n271618 , n271619 , n271620 , n271621 , n271622 , n271623 , n271624 , n271625 , 
     n271626 , n271627 , n271628 , n271629 , n271630 , n271631 , n271632 , n271633 , n271634 , n271635 , 
     n271636 , n271637 , n271638 , n271639 , n271640 , n271641 , n271642 , n271643 , n271644 , n271645 , 
     n271646 , n271647 , n271648 , n271649 , n271650 , n271651 , n271652 , n271653 , n271654 , n271655 , 
     n271656 , n271657 , n271658 , n271659 , n271660 , n271661 , n271662 , n271663 , n271664 , n271665 , 
     n271666 , n271667 , n271668 , n271669 , n271670 , n271671 , n271672 , n271673 , n271674 , n271675 , 
     n271676 , n271677 , n271678 , n271679 , n271680 , n271681 , n271682 , n271683 , n271684 , n271685 , 
     n271686 , n271687 , n271688 , n271689 , n271690 , n271691 , n271692 , n271693 , n271694 , n271695 , 
     n271696 , n271697 , n271698 , n271699 , n271700 , n271701 , n271702 , n271703 , n271704 , n271705 , 
     n271706 , n271707 , n271708 , n271709 , n271710 , n271711 , n271712 , n271713 , n271714 , n271715 , 
     n271716 , n271717 , n271718 , n271719 , n271720 , n271721 , n271722 , n271723 , n271724 , n271725 , 
     n271726 , n271727 , n271728 , n271729 , n271730 , n271731 , n271732 , n271733 , n271734 , n271735 , 
     n271736 , n271737 , n271738 , n271739 , n271740 , n271741 , n271742 , n271743 , n271744 , n271745 , 
     n271746 , n271747 , n271748 , n271749 , n271750 , n271751 , n271752 , n271753 , n271754 , n271755 , 
     n271756 , n271757 , n271758 , n271759 , n271760 , n271761 , n271762 , n271763 , n271764 , n271765 , 
     n271766 , n271767 , n271768 , n271769 , n271770 , n271771 , n271772 , n271773 , n271774 , n271775 , 
     n271776 , n271777 , n271778 , n271779 , n271780 , n271781 , n271782 , n271783 , n271784 , n271785 , 
     n271786 , n271787 , n271788 , n271789 , n271790 , n271791 , n271792 , n271793 , n271794 , n271795 , 
     n271796 , n271797 , n271798 , n271799 , n271800 , n271801 , n271802 , n271803 , n271804 , n271805 , 
     n271806 , n271807 , n271808 , n271809 , n271810 , n271811 , n271812 , n271813 , n271814 , n271815 , 
     n271816 , n271817 , n271818 , n271819 , n271820 , n271821 , n271822 , n271823 , n271824 , n271825 , 
     n271826 , n271827 , n271828 , n271829 , n271830 , n271831 , n271832 , n271833 , n271834 , n271835 , 
     n271836 , n271837 , n271838 , n271839 , n271840 , n271841 , n271842 , n271843 , n271844 , n271845 , 
     n271846 , n271847 , n271848 , n271849 , n271850 , n271851 , n271852 , n271853 , n271854 , n271855 , 
     n271856 , n271857 , n271858 , n271859 , n271860 , n271861 , n271862 , n271863 , n271864 , n271865 , 
     n271866 , n271867 , n271868 , n271869 , n271870 , n271871 , n271872 , n271873 , n271874 , n271875 , 
     n271876 , n271877 , n271878 , n271879 , n271880 , n271881 , n271882 , n271883 , n271884 , n271885 , 
     n271886 , n271887 , n271888 , n271889 , n271890 , n271891 , n271892 , n271893 , n271894 , n271895 , 
     n271896 , n271897 , n271898 , n271899 , n271900 , n271901 , n271902 , n271903 , n271904 , n271905 , 
     n271906 , n271907 , n271908 , n271909 , n271910 , n271911 , n271912 , n271913 , n271914 , n271915 , 
     n271916 , n271917 , n271918 , n271919 , n271920 , n271921 , n271922 , n271923 , n271924 , n271925 , 
     n271926 , n271927 , n271928 , n271929 , n271930 , n271931 , n271932 , n271933 , n271934 , n271935 , 
     n271936 , n271937 , n271938 , n271939 , n271940 , n271941 , n271942 , n271943 , n271944 , n271945 , 
     n271946 , n271947 , n271948 , n271949 , n271950 , n271951 , n271952 , n271953 , n271954 , n271955 , 
     n271956 , n271957 , n271958 , n271959 , n271960 , n271961 , n271962 , n271963 , n271964 , n271965 , 
     n271966 , n271967 , n271968 , n271969 , n271970 , n271971 , n271972 , n271973 , n271974 , n271975 , 
     n271976 , n271977 , n271978 , n271979 , n271980 , n271981 , n271982 , n271983 , n271984 , n271985 , 
     n271986 , n271987 , n271988 , n271989 , n271990 , n271991 , n271992 , n271993 , n271994 , n271995 , 
     n271996 , n271997 , n271998 , n271999 , n272000 , n272001 , n272002 , n272003 , n272004 , n272005 , 
     n272006 , n272007 , n272008 , n272009 , n272010 , n272011 , n272012 , n272013 , n272014 , n272015 , 
     n272016 , n272017 , n272018 , n272019 , n272020 , n272021 , n272022 , n272023 , n272024 , n272025 , 
     n272026 , n272027 , n272028 , n272029 , n272030 , n272031 , n272032 , n272033 , n272034 , n272035 , 
     n272036 , n272037 , n272038 , n272039 , n272040 , n272041 , n272042 , n272043 , n272044 , n272045 , 
     n272046 , n272047 , n272048 , n272049 , n272050 , n272051 , n272052 , n272053 , n272054 , n272055 , 
     n272056 , n272057 , n272058 , n272059 , n272060 , n272061 , n272062 , n272063 , n272064 , n272065 , 
     n272066 , n272067 , n272068 , n272069 , n272070 , n272071 , n272072 , n272073 , n272074 , n272075 , 
     n272076 , n272077 , n272078 , n272079 , n272080 , n272081 , n272082 , n272083 , n272084 , n272085 , 
     n272086 , n272087 , n272088 , n272089 , n272090 , n272091 , n272092 , n272093 , n272094 , n272095 , 
     n272096 , n272097 , n272098 , n272099 , n272100 , n272101 , n272102 , n272103 , n272104 , n272105 , 
     n272106 , n272107 , n272108 , n272109 , n272110 , n272111 , n272112 , n272113 , n272114 , n272115 , 
     n272116 , n272117 , n272118 , n272119 , n272120 , n272121 , n272122 , n272123 , n272124 , n272125 , 
     n272126 , n272127 , n272128 , n272129 , n272130 , n272131 , n272132 , n272133 , n272134 , n272135 , 
     n272136 , n272137 , n272138 , n272139 , n272140 , n272141 , n272142 , n272143 , n272144 , n272145 , 
     n272146 , n272147 , n272148 , n272149 , n272150 , n272151 , n272152 , n272153 , n272154 , n272155 , 
     n272156 , n272157 , n272158 , n272159 , n272160 , n272161 , n272162 , n272163 , n272164 , n272165 , 
     n272166 , n272167 , n272168 , n272169 , n272170 , n272171 , n272172 , n272173 , n272174 , n272175 , 
     n272176 , n272177 , n272178 , n272179 , n272180 , n272181 , n272182 , n272183 , n272184 , n272185 , 
     n272186 , n272187 , n272188 , n272189 , n272190 , n272191 , n272192 , n272193 , n272194 , n272195 , 
     n272196 , n272197 , n272198 , n272199 , n272200 , n272201 , n272202 , n272203 , n272204 , n272205 , 
     n272206 , n272207 , n272208 , n272209 , n272210 , n272211 , n272212 , n272213 , n272214 , n272215 , 
     n272216 , n272217 , n272218 , n272219 , n272220 , n272221 , n272222 , n272223 , n272224 , n272225 , 
     n272226 , n272227 , n272228 , n272229 , n272230 , n272231 , n272232 , n272233 , n272234 , n272235 , 
     n272236 , n272237 , n272238 , n272239 , n272240 , n272241 , n272242 , n272243 , n272244 , n272245 , 
     n272246 , n272247 , n272248 , n272249 , n272250 , n272251 , n272252 , n272253 , n272254 , n272255 , 
     n272256 , n272257 , n272258 , n272259 , n272260 , n272261 , n272262 , n272263 , n272264 , n272265 , 
     n272266 , n272267 , n272268 , n272269 , n272270 , n272271 , n272272 , n272273 , n272274 , n272275 , 
     n272276 , n272277 , n272278 , n272279 , n272280 , n272281 , n272282 , n272283 , n272284 , n272285 , 
     n272286 , n272287 , n272288 , n272289 , n272290 , n272291 , n272292 , n272293 , n272294 , n272295 , 
     n272296 , n272297 , n272298 , n272299 , n272300 , n272301 , n272302 , n272303 , n272304 , n272305 , 
     n272306 , n272307 , n272308 , n272309 , n272310 , n272311 , n272312 , n272313 , n272314 , n272315 , 
     n272316 , n272317 , n272318 , n272319 , n272320 , n272321 , n272322 , n272323 , n272324 , n272325 , 
     n272326 , n272327 , n272328 , n272329 , n272330 , n272331 , n272332 , n272333 , n272334 , n272335 , 
     n272336 , n272337 , n272338 , n272339 , n272340 , n272341 , n272342 , n272343 , n272344 , n272345 , 
     n272346 , n272347 , n272348 , n272349 , n272350 , n272351 , n272352 , n272353 , n272354 , n272355 , 
     n272356 , n272357 , n272358 , n272359 , n272360 , n272361 , n272362 , n272363 , n272364 , n272365 , 
     n272366 , n272367 , n272368 , n272369 , n272370 , n272371 , n272372 , n272373 , n272374 , n272375 , 
     n272376 , n272377 , n272378 , n272379 , n272380 , n272381 , n272382 , n272383 , n272384 , n272385 , 
     n272386 , n272387 , n272388 , n272389 , n272390 , n272391 , n272392 , n272393 , n272394 , n272395 , 
     n272396 , n272397 , n272398 , n272399 , n272400 , n272401 , n272402 , n272403 , n272404 , n272405 , 
     n272406 , n272407 , n272408 , n272409 , n272410 , n272411 , n272412 , n272413 , n272414 , n272415 , 
     n272416 , n272417 , n272418 , n272419 , n272420 , n272421 , n272422 , n272423 , n272424 , n272425 , 
     n272426 , n272427 , n272428 , n272429 , n272430 , n272431 , n272432 , n272433 , n272434 , n272435 , 
     n272436 , n272437 , n272438 , n272439 , n272440 , n272441 , n272442 , n272443 , n272444 , n272445 , 
     n272446 , n272447 , n272448 , n272449 , n272450 , n272451 , n272452 , n272453 , n272454 , n272455 , 
     n272456 , n272457 , n272458 , n272459 , n272460 , n272461 , n272462 , n272463 , n272464 , n272465 , 
     n272466 , n272467 , n272468 , n272469 , n272470 , n272471 , n272472 , n272473 , n272474 , n272475 , 
     n272476 , n272477 , n272478 , n272479 , n272480 , n272481 , n272482 , n272483 , n272484 , n272485 , 
     n272486 , n272487 , n272488 , n272489 , n272490 , n272491 , n272492 , n272493 , n272494 , n272495 , 
     n272496 , n272497 , n272498 , n272499 , n272500 , n272501 , n272502 , n272503 , n272504 , n272505 , 
     n272506 , n272507 , n272508 , n272509 , n272510 , n272511 , n272512 , n272513 , n272514 , n272515 , 
     n272516 , n272517 , n272518 , n272519 , n272520 , n272521 , n272522 , n272523 , n272524 , n272525 , 
     n272526 , n272527 , n272528 , n272529 , n272530 , n272531 , n272532 , n272533 , n272534 , n272535 , 
     n272536 , n272537 , n272538 , n272539 , n272540 , n272541 , n272542 , n272543 , n272544 , n272545 , 
     n272546 , n272547 , n272548 , n272549 , n272550 , n272551 , n272552 , n272553 , n272554 , n272555 , 
     n272556 , n272557 , n272558 , n272559 , n272560 , n272561 , n272562 , n272563 , n272564 , n272565 , 
     n272566 , n272567 , n272568 , n272569 , n272570 , n272571 , n272572 , n272573 , n272574 , n272575 , 
     n272576 , n272577 , n272578 , n272579 , n272580 , n272581 , n272582 , n272583 , n272584 , n272585 , 
     n272586 , n272587 , n272588 , n272589 , n272590 , n272591 , n272592 , n272593 , n272594 , n272595 , 
     n272596 , n272597 , n272598 , n272599 , n272600 , n272601 , n272602 , n272603 , n272604 , n272605 , 
     n272606 , n272607 , n272608 , n272609 , n272610 , n272611 , n272612 , n272613 , n272614 , n272615 , 
     n272616 , n272617 , n272618 , n272619 , n272620 , n272621 , n272622 , n272623 , n272624 , n272625 , 
     n272626 , n272627 , n272628 , n272629 , n272630 , n272631 , n272632 , n272633 , n272634 , n272635 , 
     n272636 , n272637 , n272638 , n272639 , n272640 , n272641 , n272642 , n272643 , n272644 , n272645 , 
     n272646 , n272647 , n272648 , n272649 , n272650 , n272651 , n272652 , n272653 , n272654 , n272655 , 
     n272656 , n272657 , n272658 , n272659 , n272660 , n272661 , n272662 , n272663 , n272664 , n272665 , 
     n272666 , n272667 , n272668 , n272669 , n272670 , n272671 , n272672 , n272673 , n272674 , n272675 , 
     n272676 , n272677 , n272678 , n272679 , n272680 , n272681 , n272682 , n272683 , n272684 , n272685 , 
     n272686 , n272687 , n272688 , n272689 , n272690 , n272691 , n272692 , n272693 , n272694 , n272695 , 
     n272696 , n272697 , n272698 , n272699 , n272700 , n272701 , n272702 , n272703 , n272704 , n272705 , 
     n272706 , n272707 , n272708 , n272709 , n272710 , n272711 , n272712 , n272713 , n272714 , n272715 , 
     n272716 , n272717 , n272718 , n272719 , n272720 , n272721 , n272722 , n272723 , n272724 , n272725 , 
     n272726 , n272727 , n272728 , n272729 , n272730 , n272731 , n272732 , n272733 , n272734 , n272735 , 
     n272736 , n272737 , n272738 , n272739 , n272740 , n272741 , n272742 , n272743 , n272744 , n272745 , 
     n272746 , n272747 , n272748 , n272749 , n272750 , n272751 , n272752 , n272753 , n272754 , n272755 , 
     n272756 , n272757 , n272758 , n272759 , n272760 , n272761 , n272762 , n272763 , n272764 , n272765 , 
     n272766 , n272767 , n272768 , n272769 , n272770 , n272771 , n272772 , n272773 , n272774 , n272775 , 
     n272776 , n272777 , n272778 , n272779 , n272780 , n272781 , n272782 , n272783 , n272784 , n272785 , 
     n272786 , n272787 , n272788 , n272789 , n272790 , n272791 , n272792 , n272793 , n272794 , n272795 , 
     n272796 , n272797 , n272798 , n272799 , n272800 , n272801 , n272802 , n272803 , n272804 , n272805 , 
     n272806 , n272807 , n272808 , n272809 , n272810 , n272811 , n272812 , n272813 , n272814 , n272815 , 
     n272816 , n272817 , n272818 , n272819 , n272820 , n272821 , n272822 , n272823 , n272824 , n272825 , 
     n272826 , n272827 , n272828 , n272829 , n272830 , n272831 , n272832 , n272833 , n272834 , n272835 , 
     n272836 , n272837 , n272838 , n272839 , n272840 , n272841 , n272842 , n272843 , n272844 , n272845 , 
     n272846 , n272847 , n272848 , n272849 , n272850 , n272851 , n272852 , n272853 , n272854 , n272855 , 
     n272856 , n272857 , n272858 , n272859 , n272860 , n272861 , n272862 , n272863 , n272864 , n272865 , 
     n272866 , n272867 , n272868 , n272869 , n272870 , n272871 , n272872 , n272873 , n272874 , n272875 , 
     n272876 , n272877 , n272878 , n272879 , n272880 , n272881 , n272882 , n272883 , n272884 , n272885 , 
     n272886 , n272887 , n272888 , n272889 , n272890 , n272891 , n272892 , n272893 , n272894 , n272895 , 
     n272896 , n272897 , n272898 , n272899 , n272900 , n272901 , n272902 , n272903 , n272904 , n272905 , 
     n272906 , n272907 , n272908 , n272909 , n272910 , n272911 , n272912 , n272913 , n272914 , n272915 , 
     n272916 , n272917 , n272918 , n272919 , n272920 , n272921 , n272922 , n272923 , n272924 , n272925 , 
     n272926 , n272927 , n272928 , n272929 , n272930 , n272931 , n272932 , n272933 , n272934 , n272935 , 
     n272936 , n272937 , n272938 , n272939 , n272940 , n272941 , n272942 , n272943 , n272944 , n272945 , 
     n272946 , n272947 , n272948 , n272949 , n272950 , n272951 , n272952 , n272953 , n272954 , n272955 , 
     n272956 , n272957 , n272958 , n272959 , n272960 , n272961 , n272962 , n272963 , n272964 , n272965 , 
     n272966 , n272967 , n272968 , n272969 , n272970 , n272971 , n272972 , n272973 , n272974 , n272975 , 
     n272976 , n272977 , n272978 , n272979 , n272980 , n272981 , n272982 , n272983 , n272984 , n272985 , 
     n272986 , n272987 , n272988 , n272989 , n272990 , n272991 , n272992 , n272993 , n272994 , n272995 , 
     n272996 , n272997 , n272998 , n272999 , n273000 , n273001 , n273002 , n273003 , n273004 , n273005 , 
     n273006 , n273007 , n273008 , n273009 , n273010 , n273011 , n273012 , n273013 , n273014 , n273015 , 
     n273016 , n273017 , n273018 , n273019 , n273020 , n273021 , n273022 , n273023 , n273024 , n273025 , 
     n273026 , n273027 , n273028 , n273029 , n273030 , n273031 , n273032 , n273033 , n273034 , n273035 , 
     n273036 , n273037 , n273038 , n273039 , n273040 , n273041 , n273042 , n273043 , n273044 , n273045 , 
     n273046 , n273047 , n273048 , n273049 , n273050 , n273051 , n273052 , n273053 , n273054 , n273055 , 
     n273056 , n273057 , n273058 , n273059 , n273060 , n273061 , n273062 , n273063 , n273064 , n273065 , 
     n273066 , n273067 , n273068 , n273069 , n273070 , n273071 , n273072 , n273073 , n273074 , n273075 , 
     n273076 , n273077 , n273078 , n273079 , n273080 , n273081 , n273082 , n273083 , n273084 , n273085 , 
     n273086 , n273087 , n273088 , n273089 , n273090 , n273091 , n273092 , n273093 , n273094 , n273095 , 
     n273096 , n273097 , n273098 , n273099 , n273100 , n273101 , n273102 , n273103 , n273104 , n273105 , 
     n273106 , n273107 , n273108 , n273109 , n273110 , n273111 , n273112 , n273113 , n273114 , n273115 , 
     n273116 , n273117 , n273118 , n273119 , n273120 , n273121 , n273122 , n273123 , n273124 , n273125 , 
     n273126 , n273127 , n273128 , n273129 , n273130 , n273131 , n273132 , n273133 , n273134 , n273135 , 
     n273136 , n273137 , n273138 , n273139 , n273140 , n273141 , n273142 , n273143 , n273144 , n273145 , 
     n273146 , n273147 , n273148 , n273149 , n273150 , n273151 , n273152 , n273153 , n273154 , n273155 , 
     n273156 , n273157 , n273158 , n273159 , n273160 , n273161 , n273162 , n273163 , n273164 , n273165 , 
     n273166 , n273167 , n273168 , n273169 , n273170 , n273171 , n273172 , n273173 , n273174 , n273175 , 
     n273176 , n273177 , n273178 , n273179 , n273180 , n273181 , n273182 , n273183 , n273184 , n273185 , 
     n273186 , n273187 , n273188 , n273189 , n273190 , n273191 , n273192 , n273193 , n273194 , n273195 , 
     n273196 , n273197 , n273198 , n273199 , n273200 , n273201 , n273202 , n273203 , n273204 , n273205 , 
     n273206 , n273207 , n273208 , n273209 , n273210 , n273211 , n273212 , n273213 , n273214 , n273215 , 
     n273216 , n273217 , n273218 , n273219 , n273220 , n273221 , n273222 , n273223 , n273224 , n273225 , 
     n273226 , n273227 , n273228 , n273229 , n273230 , n273231 , n273232 , n273233 , n273234 , n273235 , 
     n273236 , n273237 , n273238 , n273239 , n273240 , n273241 , n273242 , n273243 , n273244 , n273245 , 
     n273246 , n273247 , n273248 , n273249 , n273250 , n273251 , n273252 , n273253 , n273254 , n273255 , 
     n273256 , n273257 , n273258 , n273259 , n273260 , n273261 , n273262 , n273263 , n273264 , n273265 , 
     n273266 , n273267 , n273268 , n273269 , n273270 , n273271 , n273272 , n273273 , n273274 , n273275 , 
     n273276 , n273277 , n273278 , n273279 , n273280 , n273281 , n273282 , n273283 , n273284 , n273285 , 
     n273286 , n273287 , n273288 , n273289 , n273290 , n273291 , n273292 , n273293 , n273294 , n273295 , 
     n273296 , n273297 , n273298 , n273299 , n273300 , n273301 , n273302 , n273303 , n273304 , n273305 , 
     n273306 , n273307 , n273308 , n273309 , n273310 , n273311 , n273312 , n273313 , n273314 , n273315 , 
     n273316 , n273317 , n273318 , n273319 , n273320 , n273321 , n273322 , n273323 , n273324 , n273325 , 
     n273326 , n273327 , n273328 , n273329 , n273330 , n273331 , n273332 , n273333 , n273334 , n273335 , 
     n273336 , n273337 , n273338 , n273339 , n273340 , n273341 , n273342 , n273343 , n273344 , n273345 , 
     n273346 , n273347 , n273348 , n273349 , n273350 , n273351 , n273352 , n273353 , n273354 , n273355 , 
     n273356 , n273357 , n273358 , n273359 , n273360 , n273361 , n273362 , n273363 , n273364 , n273365 , 
     n273366 , n273367 , n273368 , n273369 , n273370 , n273371 , n273372 , n273373 , n273374 , n273375 , 
     n273376 , n273377 , n273378 , n273379 , n273380 , n273381 , n273382 , n273383 , n273384 , n273385 , 
     n273386 , n273387 , n273388 , n273389 , n273390 , n273391 , n273392 , n273393 , n273394 , n273395 , 
     n273396 , n273397 , n273398 , n273399 , n273400 , n273401 , n273402 , n273403 , n273404 , n273405 , 
     n273406 , n273407 , n273408 , n273409 , n273410 , n273411 , n273412 , n273413 , n273414 , n273415 , 
     n273416 , n273417 , n273418 , n273419 , n273420 , n273421 , n273422 , n273423 , n273424 , n273425 , 
     n273426 , n273427 , n273428 , n273429 , n273430 , n273431 , n273432 , n273433 , n273434 , n273435 , 
     n273436 , n273437 , n273438 , n273439 , n273440 , n273441 , n273442 , n273443 , n273444 , n273445 , 
     n273446 , n273447 , n273448 , n273449 , n273450 , n273451 , n273452 , n273453 , n273454 , n273455 , 
     n273456 , n273457 , n273458 , n273459 , n273460 , n273461 , n273462 , n273463 , n273464 , n273465 , 
     n273466 , n273467 , n273468 , n273469 , n273470 , n273471 , n273472 , n273473 , n273474 , n273475 , 
     n273476 , n273477 , n273478 , n273479 , n273480 , n273481 , n273482 , n273483 , n273484 , n273485 , 
     n273486 , n273487 , n273488 , n273489 , n273490 , n273491 , n273492 , n273493 , n273494 , n273495 , 
     n273496 , n273497 , n273498 , n273499 , n273500 , n273501 , n273502 , n273503 , n273504 , n273505 , 
     n273506 , n273507 , n273508 , n273509 , n273510 , n273511 , n273512 , n273513 , n273514 , n273515 , 
     n273516 , n273517 , n273518 , n273519 , n273520 , n273521 , n273522 , n273523 , n273524 , n273525 , 
     n273526 , n273527 , n273528 , n273529 , n273530 , n273531 , n273532 , n273533 , n273534 , n273535 , 
     n273536 , n273537 , n273538 , n273539 , n273540 , n273541 , n273542 , n273543 , n273544 , n273545 , 
     n273546 , n273547 , n273548 , n273549 , n273550 , n273551 , n273552 , n273553 , n273554 , n273555 , 
     n273556 , n273557 , n273558 , n273559 , n273560 , n273561 , n273562 , n273563 , n273564 , n273565 , 
     n273566 , n273567 , n273568 , n273569 , n273570 , n273571 , n273572 , n273573 , n273574 , n273575 , 
     n273576 , n273577 , n273578 , n273579 , n273580 , n273581 , n273582 , n273583 , n273584 , n273585 , 
     n273586 , n273587 , n273588 , n273589 , n273590 , n273591 , n273592 , n273593 , n273594 , n273595 , 
     n273596 , n273597 , n273598 , n273599 , n273600 , n273601 , n273602 , n273603 , n273604 , n273605 , 
     n273606 , n273607 , n273608 , n273609 , n273610 , n273611 , n273612 , n273613 , n273614 , n273615 , 
     n273616 , n273617 , n273618 , n273619 , n273620 , n273621 , n273622 , n273623 , n273624 , n273625 , 
     n273626 , n273627 , n273628 , n273629 , n273630 , n273631 , n273632 , n273633 , n273634 , n273635 , 
     n273636 , n273637 , n273638 , n273639 , n273640 , n273641 , n273642 , n273643 , n273644 , n273645 , 
     n273646 , n273647 , n273648 , n273649 , n273650 , n273651 , n273652 , n273653 , n273654 , n273655 , 
     n273656 , n273657 , n273658 , n273659 , n273660 , n273661 , n273662 , n273663 , n273664 , n273665 , 
     n273666 , n273667 , n273668 , n273669 , n273670 , n273671 , n273672 , n273673 , n273674 , n273675 , 
     n273676 , n273677 , n273678 , n273679 , n273680 , n273681 , n273682 , n273683 , n273684 , n273685 , 
     n273686 , n273687 , n273688 , n273689 , n273690 , n273691 , n273692 , n273693 , n273694 , n273695 , 
     n273696 , n273697 , n273698 , n273699 , n273700 , n273701 , n273702 , n273703 , n273704 , n273705 , 
     n273706 , n273707 , n273708 , n273709 , n273710 , n273711 , n273712 , n273713 , n273714 , n273715 , 
     n273716 , n273717 , n273718 , n273719 , n273720 , n273721 , n273722 , n273723 , n273724 , n273725 , 
     n273726 , n273727 , n273728 , n273729 , n273730 , n273731 , n273732 , n273733 , n273734 , n273735 , 
     n273736 , n273737 , n273738 , n273739 , n273740 , n273741 , n273742 , n273743 , n273744 , n273745 , 
     n273746 , n273747 , n273748 , n273749 , n273750 , n273751 , n273752 , n273753 , n273754 , n273755 , 
     n273756 , n273757 , n273758 , n273759 , n273760 , n273761 , n273762 , n273763 , n273764 , n273765 , 
     n273766 , n273767 , n273768 , n273769 , n273770 , n273771 , n273772 , n273773 , n273774 , n273775 , 
     n273776 , n273777 , n273778 , n273779 , n273780 , n273781 , n273782 , n273783 , n273784 , n273785 , 
     n273786 , n273787 , n273788 , n273789 , n273790 , n273791 , n273792 , n273793 , n273794 , n273795 , 
     n273796 , n273797 , n273798 , n273799 , n273800 , n273801 , n273802 , n273803 , n273804 , n273805 , 
     n273806 , n273807 , n273808 , n273809 , n273810 , n273811 , n273812 , n273813 , n273814 , n273815 , 
     n273816 , n273817 , n273818 , n273819 , n273820 , n273821 , n273822 , n273823 , n273824 , n273825 , 
     n273826 , n273827 , n273828 , n273829 , n273830 , n273831 , n273832 , n273833 , n273834 , n273835 , 
     n273836 , n273837 , n273838 , n273839 , n273840 , n273841 , n273842 , n273843 , n273844 , n273845 , 
     n273846 , n273847 , n273848 , n273849 , n273850 , n273851 , n273852 , n273853 , n273854 , n273855 , 
     n273856 , n273857 , n273858 , n273859 , n273860 , n273861 , n273862 , n273863 , n273864 , n273865 , 
     n273866 , n273867 , n273868 , n273869 , n273870 , n273871 , n273872 , n273873 , n273874 , n273875 , 
     n273876 , n273877 , n273878 , n273879 , n273880 , n273881 , n273882 , n273883 , n273884 , n273885 , 
     n273886 , n273887 , n273888 , n273889 , n273890 , n273891 , n273892 , n273893 , n273894 , n273895 , 
     n273896 , n273897 , n273898 , n273899 , n273900 , n273901 , n273902 , n273903 , n273904 , n273905 , 
     n273906 , n273907 , n273908 , n273909 , n273910 , n273911 , n273912 , n273913 , n273914 , n273915 , 
     n273916 , n273917 , n273918 , n273919 , n273920 , n273921 , n273922 , n273923 , n273924 , n273925 , 
     n273926 , n273927 , n273928 , n273929 , n273930 , n273931 , n273932 , n273933 , n273934 , n273935 , 
     n273936 , n273937 , n273938 , n273939 , n273940 , n273941 , n273942 , n273943 , n273944 , n273945 , 
     n273946 , n273947 , n273948 , n273949 , n273950 , n273951 , n273952 , n273953 , n273954 , n273955 , 
     n273956 , n273957 , n273958 , n273959 , n273960 , n273961 , n273962 , n273963 , n273964 , n273965 , 
     n273966 , n273967 , n273968 , n273969 , n273970 , n273971 , n273972 , n273973 , n273974 , n273975 , 
     n273976 , n273977 , n273978 , n273979 , n273980 , n273981 , n273982 , n273983 , n273984 , n273985 , 
     n273986 , n273987 , n273988 , n273989 , n273990 , n273991 , n273992 , n273993 , n273994 , n273995 , 
     n273996 , n273997 , n273998 , n273999 , n274000 , n274001 , n274002 , n274003 , n274004 , n274005 , 
     n274006 , n274007 , n274008 , n274009 , n274010 , n274011 , n274012 , n274013 , n274014 , n274015 , 
     n274016 , n274017 , n274018 , n274019 , n274020 , n274021 , n274022 , n274023 , n274024 , n274025 , 
     n274026 , n274027 , n274028 , n274029 , n274030 , n274031 , n274032 , n274033 , n274034 , n274035 , 
     n274036 , n274037 , n274038 , n274039 , n274040 , n274041 , n274042 , n274043 , n274044 , n274045 , 
     n274046 , n274047 , n274048 , n274049 , n274050 , n274051 , n274052 , n274053 , n274054 , n274055 , 
     n274056 , n274057 , n274058 , n274059 , n274060 , n274061 , n274062 , n274063 , n274064 , n274065 , 
     n274066 , n274067 , n274068 , n274069 , n274070 , n274071 , n274072 , n274073 , n274074 , n274075 , 
     n274076 , n274077 , n274078 , n274079 , n274080 , n274081 , n274082 , n274083 , n274084 , n274085 , 
     n274086 , n274087 , n274088 , n274089 , n274090 , n274091 , n274092 , n274093 , n274094 , n274095 , 
     n274096 , n274097 , n274098 , n274099 , n274100 , n274101 , n274102 , n274103 , n274104 , n274105 , 
     n274106 , n274107 , n274108 , n274109 , n274110 , n274111 , n274112 , n274113 , n274114 , n274115 , 
     n274116 , n274117 , n274118 , n274119 , n274120 , n274121 , n274122 , n274123 , n274124 , n274125 , 
     n274126 , n274127 , n274128 , n274129 , n274130 , n274131 , n274132 , n274133 , n274134 , n274135 , 
     n274136 , n274137 , n274138 , n274139 , n274140 , n274141 , n274142 , n274143 , n274144 , n274145 , 
     n274146 , n274147 , n274148 , n274149 , n274150 , n274151 , n274152 , n274153 , n274154 , n274155 , 
     n274156 , n274157 , n274158 , n274159 , n274160 , n274161 , n274162 , n274163 , n274164 , n274165 , 
     n274166 , n274167 , n274168 , n274169 , n274170 , n274171 , n274172 , n274173 , n274174 , n274175 , 
     n274176 , n274177 , n274178 , n274179 , n274180 , n274181 , n274182 , n274183 , n274184 , n274185 , 
     n274186 , n274187 , n274188 , n274189 , n274190 , n274191 , n274192 , n274193 , n274194 , n274195 , 
     n274196 , n274197 , n274198 , n274199 , n274200 , n274201 , n274202 , n274203 , n274204 , n274205 , 
     n274206 , n274207 , n274208 , n274209 , n274210 , n274211 , n274212 , n274213 , n274214 , n274215 , 
     n274216 , n274217 , n274218 , n274219 , n274220 , n274221 , n274222 , n274223 , n274224 , n274225 , 
     n274226 , n274227 , n274228 , n274229 , n274230 , n274231 , n274232 , n274233 , n274234 , n274235 , 
     n274236 , n274237 , n274238 , n274239 , n274240 , n274241 , n274242 , n274243 , n274244 , n274245 , 
     n274246 , n274247 , n274248 , n274249 , n274250 , n274251 , n274252 , n274253 , n274254 , n274255 , 
     n274256 , n274257 , n274258 , n274259 , n274260 , n274261 , n274262 , n274263 , n274264 , n274265 , 
     n274266 , n274267 , n274268 , n274269 , n274270 , n274271 , n274272 , n274273 , n274274 , n274275 , 
     n274276 , n274277 , n274278 , n274279 , n274280 , n274281 , n274282 , n274283 , n274284 , n274285 , 
     n274286 , n274287 , n274288 , n274289 , n274290 , n274291 , n274292 , n274293 , n274294 , n274295 , 
     n274296 , n274297 , n274298 , n274299 , n274300 , n274301 , n274302 , n274303 , n274304 , n274305 , 
     n274306 , n274307 , n274308 , n274309 , n274310 , n274311 , n274312 , n274313 , n274314 , n274315 , 
     n274316 , n274317 , n274318 , n274319 , n274320 , n274321 , n274322 , n274323 , n274324 , n274325 , 
     n274326 , n274327 , n274328 , n274329 , n274330 , n274331 , n274332 , n274333 , n274334 , n274335 , 
     n274336 , n274337 , n274338 , n274339 , n274340 , n274341 , n274342 , n274343 , n274344 , n274345 , 
     n274346 , n274347 , n274348 , n274349 , n274350 , n274351 , n274352 , n274353 , n274354 , n274355 , 
     n274356 , n274357 , n274358 , n274359 , n274360 , n274361 , n274362 , n274363 , n274364 , n274365 , 
     n274366 , n274367 , n274368 , n274369 , n274370 , n274371 , n274372 , n274373 , n274374 , n274375 , 
     n274376 , n274377 , n274378 , n274379 , n274380 , n274381 , n274382 , n274383 , n274384 , n274385 , 
     n274386 , n274387 , n274388 , n274389 , n274390 , n274391 , n274392 , n274393 , n274394 , n274395 , 
     n274396 , n274397 , n274398 , n274399 , n274400 , n274401 , n274402 , n274403 , n274404 , n274405 , 
     n274406 , n274407 , n274408 , n274409 , n274410 , n274411 , n274412 , n274413 , n274414 , n274415 , 
     n274416 , n274417 , n274418 , n274419 , n274420 , n274421 , n274422 , n274423 , n274424 , n274425 , 
     n274426 , n274427 , n274428 , n274429 , n274430 , n274431 , n274432 , n274433 , n274434 , n274435 , 
     n274436 , n274437 , n274438 , n274439 , n274440 , n274441 , n274442 , n274443 , n274444 , n274445 , 
     n274446 , n274447 , n274448 , n274449 , n274450 , n274451 , n274452 , n274453 , n274454 , n274455 , 
     n274456 , n274457 , n274458 , n274459 , n274460 , n274461 , n274462 , n274463 , n274464 , n274465 , 
     n274466 , n274467 , n274468 , n274469 , n274470 , n274471 , n274472 , n274473 , n274474 , n274475 , 
     n274476 , n274477 , n274478 , n274479 , n274480 , n274481 , n274482 , n274483 , n274484 , n274485 , 
     n274486 , n274487 , n274488 , n274489 , n274490 , n274491 , n274492 , n274493 , n274494 , n274495 , 
     n274496 , n274497 , n274498 , n274499 , n274500 , n274501 , n274502 , n274503 , n274504 , n274505 , 
     n274506 , n274507 , n274508 , n274509 , n274510 , n274511 , n274512 , n274513 , n274514 , n274515 , 
     n274516 , n274517 , n274518 , n274519 , n274520 , n274521 , n274522 , n274523 , n274524 , n274525 , 
     n274526 , n274527 , n274528 , n274529 , n274530 , n274531 , n274532 , n274533 , n274534 , n274535 , 
     n274536 , n274537 , n274538 , n274539 , n274540 , n274541 , n274542 , n274543 , n274544 , n274545 , 
     n274546 , n274547 , n274548 , n274549 , n274550 , n274551 , n274552 , n274553 , n274554 , n274555 , 
     n274556 , n274557 , n274558 , n274559 , n274560 , n274561 , n274562 , n274563 , n274564 , n274565 , 
     n274566 , n274567 , n274568 , n274569 , n274570 , n274571 , n274572 , n274573 , n274574 , n274575 , 
     n274576 , n274577 , n274578 , n274579 , n274580 , n274581 , n274582 , n274583 , n274584 , n274585 , 
     n274586 , n274587 , n274588 , n274589 , n274590 , n274591 , n274592 , n274593 , n274594 , n274595 , 
     n274596 , n274597 , n274598 , n274599 , n274600 , n274601 , n274602 , n274603 , n274604 , n274605 , 
     n274606 , n274607 , n274608 , n274609 , n274610 , n274611 , n274612 , n274613 , n274614 , n274615 , 
     n274616 , n274617 , n274618 , n274619 , n274620 , n274621 , n274622 , n274623 , n274624 , n274625 , 
     n274626 , n274627 , n274628 , n274629 , n274630 , n274631 , n274632 , n274633 , n274634 , n274635 , 
     n274636 , n274637 , n274638 , n274639 , n274640 , n274641 , n274642 , n274643 , n274644 , n274645 , 
     n274646 , n274647 , n274648 , n274649 , n274650 , n274651 , n274652 , n274653 , n274654 , n274655 , 
     n274656 , n274657 , n274658 , n274659 , n274660 , n274661 , n274662 , n274663 , n274664 , n274665 , 
     n274666 , n274667 , n274668 , n274669 , n274670 , n274671 , n274672 , n274673 , n274674 , n274675 , 
     n274676 , n274677 , n274678 , n274679 , n274680 , n274681 , n274682 , n274683 , n274684 , n274685 , 
     n274686 , n274687 , n274688 , n274689 , n274690 , n274691 , n274692 , n274693 , n274694 , n274695 , 
     n274696 , n274697 , n274698 , n274699 , n274700 , n274701 , n274702 , n274703 , n274704 , n274705 , 
     n274706 , n274707 , n274708 , n274709 , n274710 , n274711 , n274712 , n274713 , n274714 , n274715 , 
     n274716 , n274717 , n274718 , n274719 , n274720 , n274721 , n274722 , n274723 , n274724 , n274725 , 
     n274726 , n274727 , n274728 , n274729 , n274730 , n274731 , n274732 , n274733 , n274734 , n274735 , 
     n274736 , n274737 , n274738 , n274739 , n274740 , n274741 , n274742 , n274743 , n274744 , n274745 , 
     n274746 , n274747 , n274748 , n274749 , n274750 , n274751 , n274752 , n274753 , n274754 , n274755 , 
     n274756 , n274757 , n274758 , n274759 , n274760 , n274761 , n274762 , n274763 , n274764 , n274765 , 
     n274766 , n274767 , n274768 , n274769 , n274770 , n274771 , n274772 , n274773 , n274774 , n274775 , 
     n274776 , n274777 , n274778 , n274779 , n274780 , n274781 , n274782 , n274783 , n274784 , n274785 , 
     n274786 , n274787 , n274788 , n274789 , n274790 , n274791 , n274792 , n274793 , n274794 , n274795 , 
     n274796 , n274797 , n274798 , n274799 , n274800 , n274801 , n274802 , n274803 , n274804 , n274805 , 
     n274806 , n274807 , n274808 , n274809 , n274810 , n274811 , n274812 , n274813 , n274814 , n274815 , 
     n274816 , n274817 , n274818 , n274819 , n274820 , n274821 , n274822 , n274823 , n274824 , n274825 , 
     n274826 , n274827 , n274828 , n274829 , n274830 , n274831 , n274832 , n274833 , n274834 , n274835 , 
     n274836 , n274837 , n274838 , n274839 , n274840 , n274841 , n274842 , n274843 , n274844 , n274845 , 
     n274846 , n274847 , n274848 , n274849 , n274850 , n274851 , n274852 , n274853 , n274854 , n274855 , 
     n274856 , n274857 , n274858 , n274859 , n274860 , n274861 , n274862 , n274863 , n274864 , n274865 , 
     n274866 , n274867 , n274868 , n274869 , n274870 , n274871 , n274872 , n274873 , n274874 , n274875 , 
     n274876 , n274877 , n274878 , n274879 , n274880 , n274881 , n274882 , n274883 , n274884 , n274885 , 
     n274886 , n274887 , n274888 , n274889 , n274890 , n274891 , n274892 , n274893 , n274894 , n274895 , 
     n274896 , n274897 , n274898 , n274899 , n274900 , n274901 , n274902 , n274903 , n274904 , n274905 , 
     n274906 , n274907 , n274908 , n274909 , n274910 , n274911 , n274912 , n274913 , n274914 , n274915 , 
     n274916 , n274917 , n274918 , n274919 , n274920 , n274921 , n274922 , n274923 , n274924 , n274925 , 
     n274926 , n274927 , n274928 , n274929 , n274930 , n274931 , n274932 , n274933 , n274934 , n274935 , 
     n274936 , n274937 , n274938 , n274939 , n274940 , n274941 , n274942 , n274943 , n274944 , n274945 , 
     n274946 , n274947 , n274948 , n274949 , n274950 , n274951 , n274952 , n274953 , n274954 , n274955 , 
     n274956 , n274957 , n274958 , n274959 , n274960 , n274961 , n274962 , n274963 , n274964 , n274965 , 
     n274966 , n274967 , n274968 , n274969 , n274970 , n274971 , n274972 , n274973 , n274974 , n274975 , 
     n274976 , n274977 , n274978 , n274979 , n274980 , n274981 , n274982 , n274983 , n274984 , n274985 , 
     n274986 , n274987 , n274988 , n274989 , n274990 , n274991 , n274992 , n274993 , n274994 , n274995 , 
     n274996 , n274997 , n274998 , n274999 , n275000 , n275001 , n275002 , n275003 , n275004 , n275005 , 
     n275006 , n275007 , n275008 , n275009 , n275010 , n275011 , n275012 , n275013 , n275014 , n275015 , 
     n275016 , n275017 , n275018 , n275019 , n275020 , n275021 , n275022 , n275023 , n275024 , n275025 , 
     n275026 , n275027 , n275028 , n275029 , n275030 , n275031 , n275032 , n275033 , n275034 , n275035 , 
     n275036 , n275037 , n275038 , n275039 , n275040 , n275041 , n275042 , n275043 , n275044 , n275045 , 
     n275046 , n275047 , n275048 , n275049 , n275050 , n275051 , n275052 , n275053 , n275054 , n275055 , 
     n275056 , n275057 , n275058 , n275059 , n275060 , n275061 , n275062 , n275063 , n275064 , n275065 , 
     n275066 , n275067 , n275068 , n275069 , n275070 , n275071 , n275072 , n275073 , n275074 , n275075 , 
     n275076 , n275077 , n275078 , n275079 , n275080 , n275081 , n275082 , n275083 , n275084 , n275085 , 
     n275086 , n275087 , n275088 , n275089 , n275090 , n275091 , n275092 , n275093 , n275094 , n275095 , 
     n275096 , n275097 , n275098 , n275099 , n275100 , n275101 , n275102 , n275103 , n275104 , n275105 , 
     n275106 , n275107 , n275108 , n275109 , n275110 , n275111 , n275112 , n275113 , n275114 , n275115 , 
     n275116 , n275117 , n275118 , n275119 , n275120 , n275121 , n275122 , n275123 , n275124 , n275125 , 
     n275126 , n275127 , n275128 , n275129 , n275130 , n275131 , n275132 , n275133 , n275134 , n275135 , 
     n275136 , n275137 , n275138 , n275139 , n275140 , n275141 , n275142 , n275143 , n275144 , n275145 , 
     n275146 , n275147 , n275148 , n275149 , n275150 , n275151 , n275152 , n275153 , n275154 , n275155 , 
     n275156 , n275157 , n275158 , n275159 , n275160 , n275161 , n275162 , n275163 , n275164 , n275165 , 
     n275166 , n275167 , n275168 , n275169 , n275170 , n275171 , n275172 , n275173 , n275174 , n275175 , 
     n275176 , n275177 , n275178 , n275179 , n275180 , n275181 , n275182 , n275183 , n275184 , n275185 , 
     n275186 , n275187 , n275188 , n275189 , n275190 , n275191 , n275192 , n275193 , n275194 , n275195 , 
     n275196 , n275197 , n275198 , n275199 , n275200 , n275201 , n275202 , n275203 , n275204 , n275205 , 
     n275206 , n275207 , n275208 , n275209 , n275210 , n275211 , n275212 , n275213 , n275214 , n275215 , 
     n275216 , n275217 , n275218 , n275219 , n275220 , n275221 , n275222 , n275223 , n275224 , n275225 , 
     n275226 , n275227 , n275228 , n275229 , n275230 , n275231 , n275232 , n275233 , n275234 , n275235 , 
     n275236 , n275237 , n275238 , n275239 , n275240 , n275241 , n275242 , n275243 , n275244 , n275245 , 
     n275246 , n275247 , n275248 , n275249 , n275250 , n275251 , n275252 , n275253 , n275254 , n275255 , 
     n275256 , n275257 , n275258 , n275259 , n275260 , n275261 , n275262 , n275263 , n275264 , n275265 , 
     n275266 , n275267 , n275268 , n275269 , n275270 , n275271 , n275272 , n275273 , n275274 , n275275 , 
     n275276 , n275277 , n275278 , n275279 , n275280 , n275281 , n275282 , n275283 , n275284 , n275285 , 
     n275286 , n275287 , n275288 , n275289 , n275290 , n275291 , n275292 , n275293 , n275294 , n275295 , 
     n275296 , n275297 , n275298 , n275299 , n275300 , n275301 , n275302 , n275303 , n275304 , n275305 , 
     n275306 , n275307 , n275308 , n275309 , n275310 , n275311 , n275312 , n275313 , n275314 , n275315 , 
     n275316 , n275317 , n275318 , n275319 , n275320 , n275321 , n275322 , n275323 , n275324 , n275325 , 
     n275326 , n275327 , n275328 , n275329 , n275330 , n275331 , n275332 , n275333 , n275334 , n275335 , 
     n275336 , n275337 , n275338 , n275339 , n275340 , n275341 , n275342 , n275343 , n275344 , n275345 , 
     n275346 , n275347 , n275348 , n275349 , n275350 , n275351 , n275352 , n275353 , n275354 , n275355 , 
     n275356 , n275357 , n275358 , n275359 , n275360 , n275361 , n275362 , n275363 , n275364 , n275365 , 
     n275366 , n275367 , n275368 , n275369 , n275370 , n275371 , n275372 , n275373 , n275374 , n275375 , 
     n275376 , n275377 , n275378 , n275379 , n275380 , n275381 , n275382 , n275383 , n275384 , n275385 , 
     n275386 , n275387 , n275388 , n275389 , n275390 , n275391 , n275392 , n275393 , n275394 , n275395 , 
     n275396 , n275397 , n275398 , n275399 , n275400 , n275401 , n275402 , n275403 , n275404 , n275405 , 
     n275406 , n275407 , n275408 , n275409 , n275410 , n275411 , n275412 , n275413 , n275414 , n275415 , 
     n275416 , n275417 , n275418 , n275419 , n275420 , n275421 , n275422 , n275423 , n275424 , n275425 , 
     n275426 , n275427 , n275428 , n275429 , n275430 , n275431 , n275432 , n275433 , n275434 , n275435 , 
     n275436 , n275437 , n275438 , n275439 , n275440 , n275441 , n275442 , n275443 , n275444 , n275445 , 
     n275446 , n275447 , n275448 , n275449 , n275450 , n275451 , n275452 , n275453 , n275454 , n275455 , 
     n275456 , n275457 , n275458 , n275459 , n275460 , n275461 , n275462 , n275463 , n275464 , n275465 , 
     n275466 , n275467 , n275468 , n275469 , n275470 , n275471 , n275472 , n275473 , n275474 , n275475 , 
     n275476 , n275477 , n275478 , n275479 , n275480 , n275481 , n275482 , n275483 , n275484 , n275485 , 
     n275486 , n275487 , n275488 , n275489 , n275490 , n275491 , n275492 , n275493 , n275494 , n275495 , 
     n275496 , n275497 , n275498 , n275499 , n275500 , n275501 , n275502 , n275503 , n275504 , n275505 , 
     n275506 , n275507 , n275508 , n275509 , n275510 , n275511 , n275512 , n275513 , n275514 , n275515 , 
     n275516 , n275517 , n275518 , n275519 , n275520 , n275521 , n275522 , n275523 , n275524 , n275525 , 
     n275526 , n275527 , n275528 , n275529 , n275530 , n275531 , n275532 , n275533 , n275534 , n275535 , 
     n275536 , n275537 , n275538 , n275539 , n275540 , n275541 , n275542 , n275543 , n275544 , n275545 , 
     n275546 , n275547 , n275548 , n275549 , n275550 , n275551 , n275552 , n275553 , n275554 , n275555 , 
     n275556 , n275557 , n275558 , n275559 , n275560 , n275561 , n275562 , n275563 , n275564 , n275565 , 
     n275566 , n275567 , n275568 , n275569 , n275570 , n275571 , n275572 , n275573 , n275574 , n275575 , 
     n275576 , n275577 , n275578 , n275579 , n275580 , n275581 , n275582 , n275583 , n275584 , n275585 , 
     n275586 , n275587 , n275588 , n275589 , n275590 , n275591 , n275592 , n275593 , n275594 , n275595 , 
     n275596 , n275597 , n275598 , n275599 , n275600 , n275601 , n275602 , n275603 , n275604 , n275605 , 
     n275606 , n275607 , n275608 , n275609 , n275610 , n275611 , n275612 , n275613 , n275614 , n275615 , 
     n275616 , n275617 , n275618 , n275619 , n275620 , n275621 , n275622 , n275623 , n275624 , n275625 , 
     n275626 , n275627 , n275628 , n275629 , n275630 , n275631 , n275632 , n275633 , n275634 , n275635 , 
     n275636 , n275637 , n275638 , n275639 , n275640 , n275641 , n275642 , n275643 , n275644 , n275645 , 
     n275646 , n275647 , n275648 , n275649 , n275650 , n275651 , n275652 , n275653 , n275654 , n275655 , 
     n275656 , n275657 , n275658 , n275659 , n275660 , n275661 , n275662 , n275663 , n275664 , n275665 , 
     n275666 , n275667 , n275668 , n275669 , n275670 , n275671 , n275672 , n275673 , n275674 , n275675 , 
     n275676 , n275677 , n275678 , n275679 , n275680 , n275681 , n275682 , n275683 , n275684 , n275685 , 
     n275686 , n275687 , n275688 , n275689 , n275690 , n275691 , n275692 , n275693 , n275694 , n275695 , 
     n275696 , n275697 , n275698 , n275699 , n275700 , n275701 , n275702 , n275703 , n275704 , n275705 , 
     n275706 , n275707 , n275708 , n275709 , n275710 , n275711 , n275712 , n275713 , n275714 , n275715 , 
     n275716 , n275717 , n275718 , n275719 , n275720 , n275721 , n275722 , n275723 , n275724 , n275725 , 
     n275726 , n275727 , n275728 , n275729 , n275730 , n275731 , n275732 , n275733 , n275734 , n275735 , 
     n275736 , n275737 , n275738 , n275739 , n275740 , n275741 , n275742 , n275743 , n275744 , n275745 , 
     n275746 , n275747 , n275748 , n275749 , n275750 , n275751 , n275752 , n275753 , n275754 , n275755 , 
     n275756 , n275757 , n275758 , n275759 , n275760 , n275761 , n275762 , n275763 , n275764 , n275765 , 
     n275766 , n275767 , n275768 , n275769 , n275770 , n275771 , n275772 , n275773 , n275774 , n275775 , 
     n275776 , n275777 , n275778 , n275779 , n275780 , n275781 , n275782 , n275783 , n275784 , n275785 , 
     n275786 , n275787 , n275788 , n275789 , n275790 , n275791 , n275792 , n275793 , n275794 , n275795 , 
     n275796 , n275797 , n275798 , n275799 , n275800 , n275801 , n275802 , n275803 , n275804 , n275805 , 
     n275806 , n275807 , n275808 , n275809 , n275810 , n275811 , n275812 , n275813 , n275814 , n275815 , 
     n275816 , n275817 , n275818 , n275819 , n275820 , n275821 , n275822 , n275823 , n275824 , n275825 , 
     n275826 , n275827 , n275828 , n275829 , n275830 , n275831 , n275832 , n275833 , n275834 , n275835 , 
     n275836 , n275837 , n275838 , n275839 , n275840 , n275841 , n275842 , n275843 , n275844 , n275845 , 
     n275846 , n275847 , n275848 , n275849 , n275850 , n275851 , n275852 , n275853 , n275854 , n275855 , 
     n275856 , n275857 , n275858 , n275859 , n275860 , n275861 , n275862 , n275863 , n275864 , n275865 , 
     n275866 , n275867 , n275868 , n275869 , n275870 , n275871 , n275872 , n275873 , n275874 , n275875 , 
     n275876 , n275877 , n275878 , n275879 , n275880 , n275881 , n275882 , n275883 , n275884 , n275885 , 
     n275886 , n275887 , n275888 , n275889 , n275890 , n275891 , n275892 , n275893 , n275894 , n275895 , 
     n275896 , n275897 , n275898 , n275899 , n275900 , n275901 , n275902 , n275903 , n275904 , n275905 , 
     n275906 , n275907 , n275908 , n275909 , n275910 , n275911 , n275912 , n275913 , n275914 , n275915 , 
     n275916 , n275917 , n275918 , n275919 , n275920 , n275921 , n275922 , n275923 , n275924 , n275925 , 
     n275926 , n275927 , n275928 , n275929 , n275930 , n275931 , n275932 , n275933 , n275934 , n275935 , 
     n275936 , n275937 , n275938 , n275939 , n275940 , n275941 , n275942 , n275943 , n275944 , n275945 , 
     n275946 , n275947 , n275948 , n275949 , n275950 , n275951 , n275952 , n275953 , n275954 , n275955 , 
     n275956 , n275957 , n275958 , n275959 , n275960 , n275961 , n275962 , n275963 , n275964 , n275965 , 
     n275966 , n275967 , n275968 , n275969 , n275970 , n275971 , n275972 , n275973 , n275974 , n275975 , 
     n275976 , n275977 , n275978 , n275979 , n275980 , n275981 , n275982 , n275983 , n275984 , n275985 , 
     n275986 , n275987 , n275988 , n275989 , n275990 , n275991 , n275992 , n275993 , n275994 , n275995 , 
     n275996 , n275997 , n275998 , n275999 , n276000 , n276001 , n276002 , n276003 , n276004 , n276005 , 
     n276006 , n276007 , n276008 , n276009 , n276010 , n276011 , n276012 , n276013 , n276014 , n276015 , 
     n276016 , n276017 , n276018 , n276019 , n276020 , n276021 , n276022 , n276023 , n276024 , n276025 , 
     n276026 , n276027 , n276028 , n276029 , n276030 , n276031 , n276032 , n276033 , n276034 , n276035 , 
     n276036 , n276037 , n276038 , n276039 , n276040 , n276041 , n276042 , n276043 , n276044 , n276045 , 
     n276046 , n276047 , n276048 , n276049 , n276050 , n276051 , n276052 , n276053 , n276054 , n276055 , 
     n276056 , n276057 , n276058 , n276059 , n276060 , n276061 , n276062 , n276063 , n276064 , n276065 , 
     n276066 , n276067 , n276068 , n276069 , n276070 , n276071 , n276072 , n276073 , n276074 , n276075 , 
     n276076 , n276077 , n276078 , n276079 , n276080 , n276081 , n276082 , n276083 , n276084 , n276085 , 
     n276086 , n276087 , n276088 , n276089 , n276090 , n276091 , n276092 , n276093 , n276094 , n276095 , 
     n276096 , n276097 , n276098 , n276099 , n276100 , n276101 , n276102 , n276103 , n276104 , n276105 , 
     n276106 , n276107 , n276108 , n276109 , n276110 , n276111 , n276112 , n276113 , n276114 , n276115 , 
     n276116 , n276117 , n276118 , n276119 , n276120 , n276121 , n276122 , n276123 , n276124 , n276125 , 
     n276126 , n276127 , n276128 , n276129 , n276130 , n276131 , n276132 , n276133 , n276134 , n276135 , 
     n276136 , n276137 , n276138 , n276139 , n276140 , n276141 , n276142 , n276143 , n276144 , n276145 , 
     n276146 , n276147 , n276148 , n276149 , n276150 , n276151 , n276152 , n276153 , n276154 , n276155 , 
     n276156 , n276157 , n276158 , n276159 , n276160 , n276161 , n276162 , n276163 , n276164 , n276165 , 
     n276166 , n276167 , n276168 , n276169 , n276170 , n276171 , n276172 , n276173 , n276174 , n276175 , 
     n276176 , n276177 , n276178 , n276179 , n276180 , n276181 , n276182 , n276183 , n276184 , n276185 , 
     n276186 , n276187 , n276188 , n276189 , n276190 , n276191 , n276192 , n276193 , n276194 , n276195 , 
     n276196 , n276197 , n276198 , n276199 , n276200 , n276201 , n276202 , n276203 , n276204 , n276205 , 
     n276206 , n276207 , n276208 , n276209 , n276210 , n276211 , n276212 , n276213 , n276214 , n276215 , 
     n276216 , n276217 , n276218 , n276219 , n276220 , n276221 , n276222 , n276223 , n276224 , n276225 , 
     n276226 , n276227 , n276228 , n276229 , n276230 , n276231 , n276232 , n276233 , n276234 , n276235 , 
     n276236 , n276237 , n276238 , n276239 , n276240 , n276241 , n276242 , n276243 , n276244 , n276245 , 
     n276246 , n276247 , n276248 , n276249 , n276250 , n276251 , n276252 , n276253 , n276254 , n276255 , 
     n276256 , n276257 , n276258 , n276259 , n276260 , n276261 , n276262 , n276263 , n276264 , n276265 , 
     n276266 , n276267 , n276268 , n276269 , n276270 , n276271 , n276272 , n276273 , n276274 , n276275 , 
     n276276 , n276277 , n276278 , n276279 , n276280 , n276281 , n276282 , n276283 , n276284 , n276285 , 
     n276286 , n276287 , n276288 , n276289 , n276290 , n276291 , n276292 , n276293 , n276294 , n276295 , 
     n276296 , n276297 , n276298 , n276299 , n276300 , n276301 , n276302 , n276303 , n276304 , n276305 , 
     n276306 , n276307 , n276308 , n276309 , n276310 , n276311 , n276312 , n276313 , n276314 , n276315 , 
     n276316 , n276317 , n276318 , n276319 , n276320 , n276321 , n276322 , n276323 , n276324 , n276325 , 
     n276326 , n276327 , n276328 , n276329 , n276330 , n276331 , n276332 , n276333 , n276334 , n276335 , 
     n276336 , n276337 , n276338 , n276339 , n276340 , n276341 , n276342 , n276343 , n276344 , n276345 , 
     n276346 , n276347 , n276348 , n276349 , n276350 , n276351 , n276352 , n276353 , n276354 , n276355 , 
     n276356 , n276357 , n276358 , n276359 , n276360 , n276361 , n276362 , n276363 , n276364 , n276365 , 
     n276366 , n276367 , n276368 , n276369 , n276370 , n276371 , n276372 , n276373 , n276374 , n276375 , 
     n276376 , n276377 , n276378 , n276379 , n276380 , n276381 , n276382 , n276383 , n276384 , n276385 , 
     n276386 , n276387 , n276388 , n276389 , n276390 , n276391 , n276392 , n276393 , n276394 , n276395 , 
     n276396 , n276397 , n276398 , n276399 , n276400 , n276401 , n276402 , n276403 , n276404 , n276405 , 
     n276406 , n276407 , n276408 , n276409 , n276410 , n276411 , n276412 , n276413 , n276414 , n276415 , 
     n276416 , n276417 , n276418 , n276419 , n276420 , n276421 , n276422 , n276423 , n276424 , n276425 , 
     n276426 , n276427 , n276428 , n276429 , n276430 , n276431 , n276432 , n276433 , n276434 , n276435 , 
     n276436 , n276437 , n276438 , n276439 , n276440 , n276441 , n276442 , n276443 , n276444 , n276445 , 
     n276446 , n276447 , n276448 , n276449 , n276450 , n276451 , n276452 , n276453 , n276454 , n276455 , 
     n276456 , n276457 , n276458 , n276459 , n276460 , n276461 , n276462 , n276463 , n276464 , n276465 , 
     n276466 , n276467 , n276468 , n276469 , n276470 , n276471 , n276472 , n276473 , n276474 , n276475 , 
     n276476 , n276477 , n276478 , n276479 , n276480 , n276481 , n276482 , n276483 , n276484 , n276485 , 
     n276486 , n276487 , n276488 , n276489 , n276490 , n276491 , n276492 , n276493 , n276494 , n276495 , 
     n276496 , n276497 , n276498 , n276499 , n276500 , n276501 , n276502 , n276503 , n276504 , n276505 , 
     n276506 , n276507 , n276508 , n276509 , n276510 , n276511 , n276512 , n276513 , n276514 , n276515 , 
     n276516 , n276517 , n276518 , n276519 , n276520 , n276521 , n276522 , n276523 , n276524 , n276525 , 
     n276526 , n276527 , n276528 , n276529 , n276530 , n276531 , n276532 , n276533 , n276534 , n276535 , 
     n276536 , n276537 , n276538 , n276539 , n276540 , n276541 , n276542 , n276543 , n276544 , n276545 , 
     n276546 , n276547 , n276548 , n276549 , n276550 , n276551 , n276552 , n276553 , n276554 , n276555 , 
     n276556 , n276557 , n276558 , n276559 , n276560 , n276561 , n276562 , n276563 , n276564 , n276565 , 
     n276566 , n276567 , n276568 , n276569 , n276570 , n276571 , n276572 , n276573 , n276574 , n276575 , 
     n276576 , n276577 , n276578 , n276579 , n276580 , n276581 , n276582 , n276583 , n276584 , n276585 , 
     n276586 , n276587 , n276588 , n276589 , n276590 , n276591 , n276592 , n276593 , n276594 , n276595 , 
     n276596 , n276597 , n276598 , n276599 , n276600 , n276601 , n276602 , n276603 , n276604 , n276605 , 
     n276606 , n276607 , n276608 , n276609 , n276610 , n276611 , n276612 , n276613 , n276614 , n276615 , 
     n276616 , n276617 , n276618 , n276619 , n276620 , n276621 , n276622 , n276623 , n276624 , n276625 , 
     n276626 , n276627 , n276628 , n276629 , n276630 , n276631 , n276632 , n276633 , n276634 , n276635 , 
     n276636 , n276637 , n276638 , n276639 , n276640 , n276641 , n276642 , n276643 , n276644 , n276645 , 
     n276646 , n276647 , n276648 , n276649 , n276650 , n276651 , n276652 , n276653 , n276654 , n276655 , 
     n276656 , n276657 , n276658 , n276659 , n276660 , n276661 , n276662 , n276663 , n276664 , n276665 , 
     n276666 , n276667 , n276668 , n276669 , n276670 , n276671 , n276672 , n276673 , n276674 , n276675 , 
     n276676 , n276677 , n276678 , n276679 , n276680 , n276681 , n276682 , n276683 , n276684 , n276685 , 
     n276686 , n276687 , n276688 , n276689 , n276690 , n276691 , n276692 , n276693 , n276694 , n276695 , 
     n276696 , n276697 , n276698 , n276699 , n276700 , n276701 , n276702 , n276703 , n276704 , n276705 , 
     n276706 , n276707 , n276708 , n276709 , n276710 , n276711 , n276712 , n276713 , n276714 , n276715 , 
     n276716 , n276717 , n276718 , n276719 , n276720 , n276721 , n276722 , n276723 , n276724 , n276725 , 
     n276726 , n276727 , n276728 , n276729 , n276730 , n276731 , n276732 , n276733 , n276734 , n276735 , 
     n276736 , n276737 , n276738 , n276739 , n276740 , n276741 , n276742 , n276743 , n276744 , n276745 , 
     n276746 , n276747 , n276748 , n276749 , n276750 , n276751 , n276752 , n276753 , n276754 , n276755 , 
     n276756 , n276757 , n276758 , n276759 , n276760 , n276761 , n276762 , n276763 , n276764 , n276765 , 
     n276766 , n276767 , n276768 , n276769 , n276770 , n276771 , n276772 , n276773 , n276774 , n276775 , 
     n276776 , n276777 , n276778 , n276779 , n276780 , n276781 , n276782 , n276783 , n276784 , n276785 , 
     n276786 , n276787 , n276788 , n276789 , n276790 , n276791 , n276792 , n276793 , n276794 , n276795 , 
     n276796 , n276797 , n276798 , n276799 , n276800 , n276801 , n276802 , n276803 , n276804 , n276805 , 
     n276806 , n276807 , n276808 , n276809 , n276810 , n276811 , n276812 , n276813 , n276814 , n276815 , 
     n276816 , n276817 , n276818 , n276819 , n276820 , n276821 , n276822 , n276823 , n276824 , n276825 , 
     n276826 , n276827 , n276828 , n276829 , n276830 , n276831 , n276832 , n276833 , n276834 , n276835 , 
     n276836 , n276837 , n276838 , n276839 , n276840 , n276841 , n276842 , n276843 , n276844 , n276845 , 
     n276846 , n276847 , n276848 , n276849 , n276850 , n276851 , n276852 , n276853 , n276854 , n276855 , 
     n276856 , n276857 , n276858 , n276859 , n276860 , n276861 , n276862 , n276863 , n276864 , n276865 , 
     n276866 , n276867 , n276868 , n276869 , n276870 , n276871 , n276872 , n276873 , n276874 , n276875 , 
     n276876 , n276877 , n276878 , n276879 , n276880 , n276881 , n276882 , n276883 , n276884 , n276885 , 
     n276886 , n276887 , n276888 , n276889 , n276890 , n276891 , n276892 , n276893 , n276894 , n276895 , 
     n276896 , n276897 , n276898 , n276899 , n276900 , n276901 , n276902 , n276903 , n276904 , n276905 , 
     n276906 , n276907 , n276908 , n276909 , n276910 , n276911 , n276912 , n276913 , n276914 , n276915 , 
     n276916 , n276917 , n276918 , n276919 , n276920 , n276921 , n276922 , n276923 , n276924 , n276925 , 
     n276926 , n276927 , n276928 , n276929 , n276930 , n276931 , n276932 , n276933 , n276934 , n276935 , 
     n276936 , n276937 , n276938 , n276939 , n276940 , n276941 , n276942 , n276943 , n276944 , n276945 , 
     n276946 , n276947 , n276948 , n276949 , n276950 , n276951 , n276952 , n276953 , n276954 , n276955 , 
     n276956 , n276957 , n276958 , n276959 , n276960 , n276961 , n276962 , n276963 , n276964 , n276965 , 
     n276966 , n276967 , n276968 , n276969 , n276970 , n276971 , n276972 , n276973 , n276974 , n276975 , 
     n276976 , n276977 , n276978 , n276979 , n276980 , n276981 , n276982 , n276983 , n276984 , n276985 , 
     n276986 , n276987 , n276988 , n276989 , n276990 , n276991 , n276992 , n276993 , n276994 , n276995 , 
     n276996 , n276997 , n276998 , n276999 , n277000 , n277001 , n277002 , n277003 , n277004 , n277005 , 
     n277006 , n277007 , n277008 , n277009 , n277010 , n277011 , n277012 , n277013 , n277014 , n277015 , 
     n277016 , n277017 , n277018 , n277019 , n277020 , n277021 , n277022 , n277023 , n277024 , n277025 , 
     n277026 , n277027 , n277028 , n277029 , n277030 , n277031 , n277032 , n277033 , n277034 , n277035 , 
     n277036 , n277037 , n277038 , n277039 , n277040 , n277041 , n277042 , n277043 , n277044 , n277045 , 
     n277046 , n277047 , n277048 , n277049 , n277050 , n277051 , n277052 , n277053 , n277054 , n277055 , 
     n277056 , n277057 , n277058 , n277059 , n277060 , n277061 , n277062 , n277063 , n277064 , n277065 , 
     n277066 , n277067 , n277068 , n277069 , n277070 , n277071 , n277072 , n277073 , n277074 , n277075 , 
     n277076 , n277077 , n277078 , n277079 , n277080 , n277081 , n277082 , n277083 , n277084 , n277085 , 
     n277086 , n277087 , n277088 , n277089 , n277090 , n277091 , n277092 , n277093 , n277094 , n277095 , 
     n277096 , n277097 , n277098 , n277099 , n277100 , n277101 , n277102 , n277103 , n277104 , n277105 , 
     n277106 , n277107 , n277108 , n277109 , n277110 , n277111 , n277112 , n277113 , n277114 , n277115 , 
     n277116 , n277117 , n277118 , n277119 , n277120 , n277121 , n277122 , n277123 , n277124 , n277125 , 
     n277126 , n277127 , n277128 , n277129 , n277130 , n277131 , n277132 , n277133 , n277134 , n277135 , 
     n277136 , n277137 , n277138 , n277139 , n277140 , n277141 , n277142 , n277143 , n277144 , n277145 , 
     n277146 , n277147 , n277148 , n277149 , n277150 , n277151 , n277152 , n277153 , n277154 , n277155 , 
     n277156 , n277157 , n277158 , n277159 , n277160 , n277161 , n277162 , n277163 , n277164 , n277165 , 
     n277166 , n277167 , n277168 , n277169 , n277170 , n277171 , n277172 , n277173 , n277174 , n277175 , 
     n277176 , n277177 , n277178 , n277179 , n277180 , n277181 , n277182 , n277183 , n277184 , n277185 , 
     n277186 , n277187 , n277188 , n277189 , n277190 , n277191 , n277192 , n277193 , n277194 , n277195 , 
     n277196 , n277197 , n277198 , n277199 , n277200 , n277201 , n277202 , n277203 , n277204 , n277205 , 
     n277206 , n277207 , n277208 , n277209 , n277210 , n277211 , n277212 , n277213 , n277214 , n277215 , 
     n277216 , n277217 , n277218 , n277219 , n277220 , n277221 , n277222 , n277223 , n277224 , n277225 , 
     n277226 , n277227 , n277228 , n277229 , n277230 , n277231 , n277232 , n277233 , n277234 , n277235 , 
     n277236 , n277237 , n277238 , n277239 , n277240 , n277241 , n277242 , n277243 , n277244 , n277245 , 
     n277246 , n277247 , n277248 , n277249 , n277250 , n277251 , n277252 , n277253 , n277254 , n277255 , 
     n277256 , n277257 , n277258 , n277259 , n277260 , n277261 , n277262 , n277263 , n277264 , n277265 , 
     n277266 , n277267 , n277268 , n277269 , n277270 , n277271 , n277272 , n277273 , n277274 , n277275 , 
     n277276 , n277277 , n277278 , n277279 , n277280 , n277281 , n277282 , n277283 , n277284 , n277285 , 
     n277286 , n277287 , n277288 , n277289 , n277290 , n277291 , n277292 , n277293 , n277294 , n277295 , 
     n277296 , n277297 , n277298 , n277299 , n277300 , n277301 , n277302 , n277303 , n277304 , n277305 , 
     n277306 , n277307 , n277308 , n277309 , n277310 , n277311 , n277312 , n277313 , n277314 , n277315 , 
     n277316 , n277317 , n277318 , n277319 , n277320 , n277321 , n277322 , n277323 , n277324 , n277325 , 
     n277326 , n277327 , n277328 , n277329 , n277330 , n277331 , n277332 , n277333 , n277334 , n277335 , 
     n277336 , n277337 , n277338 , n277339 , n277340 , n277341 , n277342 , n277343 , n277344 , n277345 , 
     n277346 , n277347 , n277348 , n277349 , n277350 , n277351 , n277352 , n277353 , n277354 , n277355 , 
     n277356 , n277357 , n277358 , n277359 , n277360 , n277361 , n277362 , n277363 , n277364 , n277365 , 
     n277366 , n277367 , n277368 , n277369 , n277370 , n277371 , n277372 , n277373 , n277374 , n277375 , 
     n277376 , n277377 , n277378 , n277379 , n277380 , n277381 , n277382 , n277383 , n277384 , n277385 , 
     n277386 , n277387 , n277388 , n277389 , n277390 , n277391 , n277392 , n277393 , n277394 , n277395 , 
     n277396 , n277397 , n277398 , n277399 , n277400 , n277401 , n277402 , n277403 , n277404 , n277405 , 
     n277406 , n277407 , n277408 , n277409 , n277410 , n277411 , n277412 , n277413 , n277414 , n277415 , 
     n277416 , n277417 , n277418 , n277419 , n277420 , n277421 , n277422 , n277423 , n277424 , n277425 , 
     n277426 , n277427 , n277428 , n277429 , n277430 , n277431 , n277432 , n277433 , n277434 , n277435 , 
     n277436 , n277437 , n277438 , n277439 , n277440 , n277441 , n277442 , n277443 , n277444 , n277445 , 
     n277446 , n277447 , n277448 , n277449 , n277450 , n277451 , n277452 , n277453 , n277454 , n277455 , 
     n277456 , n277457 , n277458 , n277459 , n277460 , n277461 , n277462 , n277463 , n277464 , n277465 , 
     n277466 , n277467 , n277468 , n277469 , n277470 , n277471 , n277472 , n277473 , n277474 , n277475 , 
     n277476 , n277477 , n277478 , n277479 , n277480 , n277481 , n277482 , n277483 , n277484 , n277485 , 
     n277486 , n277487 , n277488 , n277489 , n277490 , n277491 , n277492 , n277493 , n277494 , n277495 , 
     n277496 , n277497 , n277498 , n277499 , n277500 , n277501 , n277502 , n277503 , n277504 , n277505 , 
     n277506 , n277507 , n277508 , n277509 , n277510 , n277511 , n277512 , n277513 , n277514 , n277515 , 
     n277516 , n277517 , n277518 , n277519 , n277520 , n277521 , n277522 , n277523 , n277524 , n277525 , 
     n277526 , n277527 , n277528 , n277529 , n277530 , n277531 , n277532 , n277533 , n277534 , n277535 , 
     n277536 , n277537 , n277538 , n277539 , n277540 , n277541 , n277542 , n277543 , n277544 , n277545 , 
     n277546 , n277547 , n277548 , n277549 , n277550 , n277551 , n277552 , n277553 , n277554 , n277555 , 
     n277556 , n277557 , n277558 , n277559 , n277560 , n277561 , n277562 , n277563 , n277564 , n277565 , 
     n277566 , n277567 , n277568 , n277569 , n277570 , n277571 , n277572 , n277573 , n277574 , n277575 , 
     n277576 , n277577 , n277578 , n277579 , n277580 , n277581 , n277582 , n277583 , n277584 , n277585 , 
     n277586 , n277587 , n277588 , n277589 , n277590 , n277591 , n277592 , n277593 , n277594 , n277595 , 
     n277596 , n277597 , n277598 , n277599 , n277600 , n277601 , n277602 , n277603 , n277604 , n277605 , 
     n277606 , n277607 , n277608 , n277609 , n277610 , n277611 , n277612 , n277613 , n277614 , n277615 , 
     n277616 , n277617 , n277618 , n277619 , n277620 , n277621 , n277622 , n277623 , n277624 , n277625 , 
     n277626 , n277627 , n277628 , n277629 , n277630 , n277631 , n277632 , n277633 , n277634 , n277635 , 
     n277636 , n277637 , n277638 , n277639 , n277640 , n277641 , n277642 , n277643 , n277644 , n277645 , 
     n277646 , n277647 , n277648 , n277649 , n277650 , n277651 , n277652 , n277653 , n277654 , n277655 , 
     n277656 , n277657 , n277658 , n277659 , n277660 , n277661 , n277662 , n277663 , n277664 , n277665 , 
     n277666 , n277667 , n277668 , n277669 , n277670 , n277671 , n277672 , n277673 , n277674 , n277675 , 
     n277676 , n277677 , n277678 , n277679 , n277680 , n277681 , n277682 , n277683 , n277684 , n277685 , 
     n277686 , n277687 , n277688 , n277689 , n277690 , n277691 , n277692 , n277693 , n277694 , n277695 , 
     n277696 , n277697 , n277698 , n277699 , n277700 , n277701 , n277702 , n277703 , n277704 , n277705 , 
     n277706 , n277707 , n277708 , n277709 , n277710 , n277711 , n277712 , n277713 , n277714 , n277715 , 
     n277716 , n277717 , n277718 , n277719 , n277720 , n277721 , n277722 , n277723 , n277724 , n277725 , 
     n277726 , n277727 , n277728 , n277729 , n277730 , n277731 , n277732 , n277733 , n277734 , n277735 , 
     n277736 , n277737 , n277738 , n277739 , n277740 , n277741 , n277742 , n277743 , n277744 , n277745 , 
     n277746 , n277747 , n277748 , n277749 , n277750 , n277751 , n277752 , n277753 , n277754 , n277755 , 
     n277756 , n277757 , n277758 , n277759 , n277760 , n277761 , n277762 , n277763 , n277764 , n277765 , 
     n277766 , n277767 , n277768 , n277769 , n277770 , n277771 , n277772 , n277773 , n277774 , n277775 , 
     n277776 , n277777 , n277778 , n277779 , n277780 , n277781 , n277782 , n277783 , n277784 , n277785 , 
     n277786 , n277787 , n277788 , n277789 , n277790 , n277791 , n277792 , n277793 , n277794 , n277795 , 
     n277796 , n277797 , n277798 , n277799 , n277800 , n277801 , n277802 , n277803 , n277804 , n277805 , 
     n277806 , n277807 , n277808 , n277809 , n277810 , n277811 , n277812 , n277813 , n277814 , n277815 , 
     n277816 , n277817 , n277818 , n277819 , n277820 , n277821 , n277822 , n277823 , n277824 , n277825 , 
     n277826 , n277827 , n277828 , n277829 , n277830 , n277831 , n277832 , n277833 , n277834 , n277835 , 
     n277836 , n277837 , n277838 , n277839 , n277840 , n277841 , n277842 , n277843 , n277844 , n277845 , 
     n277846 , n277847 , n277848 , n277849 , n277850 , n277851 , n277852 , n277853 , n277854 , n277855 , 
     n277856 , n277857 , n277858 , n277859 , n277860 , n277861 , n277862 , n277863 , n277864 , n277865 , 
     n277866 , n277867 , n277868 , n277869 , n277870 , n277871 , n277872 , n277873 , n277874 , n277875 , 
     n277876 , n277877 , n277878 , n277879 , n277880 , n277881 , n277882 , n277883 , n277884 , n277885 , 
     n277886 , n277887 , n277888 , n277889 , n277890 , n277891 , n277892 , n277893 , n277894 , n277895 , 
     n277896 , n277897 , n277898 , n277899 , n277900 , n277901 , n277902 , n277903 , n277904 , n277905 , 
     n277906 , n277907 , n277908 , n277909 , n277910 , n277911 , n277912 , n277913 , n277914 , n277915 , 
     n277916 , n277917 , n277918 , n277919 , n277920 , n277921 , n277922 , n277923 , n277924 , n277925 , 
     n277926 , n277927 , n277928 , n277929 , n277930 , n277931 , n277932 , n277933 , n277934 , n277935 , 
     n277936 , n277937 , n277938 , n277939 , n277940 , n277941 , n277942 , n277943 , n277944 , n277945 , 
     n277946 , n277947 , n277948 , n277949 , n277950 , n277951 , n277952 , n277953 , n277954 , n277955 , 
     n277956 , n277957 , n277958 , n277959 , n277960 , n277961 , n277962 , n277963 , n277964 , n277965 , 
     n277966 , n277967 , n277968 , n277969 , n277970 , n277971 , n277972 , n277973 , n277974 , n277975 , 
     n277976 , n277977 , n277978 , n277979 , n277980 , n277981 , n277982 , n277983 , n277984 , n277985 , 
     n277986 , n277987 , n277988 , n277989 , n277990 , n277991 , n277992 , n277993 , n277994 , n277995 , 
     n277996 , n277997 , n277998 , n277999 , n278000 , n278001 , n278002 , n278003 , n278004 , n278005 , 
     n278006 , n278007 , n278008 , n278009 , n278010 , n278011 , n278012 , n278013 , n278014 , n278015 , 
     n278016 , n278017 , n278018 , n278019 , n278020 , n278021 , n278022 , n278023 , n278024 , n278025 , 
     n278026 , n278027 , n278028 , n278029 , n278030 , n278031 , n278032 , n278033 , n278034 , n278035 , 
     n278036 , n278037 , n278038 , n278039 , n278040 , n278041 , n278042 , n278043 , n278044 , n278045 , 
     n278046 , n278047 , n278048 , n278049 , n278050 , n278051 , n278052 , n278053 , n278054 , n278055 , 
     n278056 , n278057 , n278058 , n278059 , n278060 , n278061 , n278062 , n278063 , n278064 , n278065 , 
     n278066 , n278067 , n278068 , n278069 , n278070 , n278071 , n278072 , n278073 , n278074 , n278075 , 
     n278076 , n278077 , n278078 , n278079 , n278080 , n278081 , n278082 , n278083 , n278084 , n278085 , 
     n278086 , n278087 , n278088 , n278089 , n278090 , n278091 , n278092 , n278093 , n278094 , n278095 , 
     n278096 , n278097 , n278098 , n278099 , n278100 , n278101 , n278102 , n278103 , n278104 , n278105 , 
     n278106 , n278107 , n278108 , n278109 , n278110 , n278111 , n278112 , n278113 , n278114 , n278115 , 
     n278116 , n278117 , n278118 , n278119 , n278120 , n278121 , n278122 , n278123 , n278124 , n278125 , 
     n278126 , n278127 , n278128 , n278129 , n278130 , n278131 , n278132 , n278133 , n278134 , n278135 , 
     n278136 , n278137 , n278138 , n278139 , n278140 , n278141 , n278142 , n278143 , n278144 , n278145 , 
     n278146 , n278147 , n278148 , n278149 , n278150 , n278151 , n278152 , n278153 , n278154 , n278155 , 
     n278156 , n278157 , n278158 , n278159 , n278160 , n278161 , n278162 , n278163 , n278164 , n278165 , 
     n278166 , n278167 , n278168 , n278169 , n278170 , n278171 , n278172 , n278173 , n278174 , n278175 , 
     n278176 , n278177 , n278178 , n278179 , n278180 , n278181 , n278182 , n278183 , n278184 , n278185 , 
     n278186 , n278187 , n278188 , n278189 , n278190 , n278191 , n278192 , n278193 , n278194 , n278195 , 
     n278196 , n278197 , n278198 , n278199 , n278200 , n278201 , n278202 , n278203 , n278204 , n278205 , 
     n278206 , n278207 , n278208 , n278209 , n278210 , n278211 , n278212 , n278213 , n278214 , n278215 , 
     n278216 , n278217 , n278218 , n278219 , n278220 , n278221 , n278222 , n278223 , n278224 , n278225 , 
     n278226 , n278227 , n278228 , n278229 , n278230 , n278231 , n278232 , n278233 , n278234 , n278235 , 
     n278236 , n278237 , n278238 , n278239 , n278240 , n278241 , n278242 , n278243 , n278244 , n278245 , 
     n278246 , n278247 , n278248 , n278249 , n278250 , n278251 , n278252 , n278253 , n278254 , n278255 , 
     n278256 , n278257 , n278258 , n278259 , n278260 , n278261 , n278262 , n278263 , n278264 , n278265 , 
     n278266 , n278267 , n278268 , n278269 , n278270 , n278271 , n278272 , n278273 , n278274 , n278275 , 
     n278276 , n278277 , n278278 , n278279 , n278280 , n278281 , n278282 , n278283 , n278284 , n278285 , 
     n278286 , n278287 , n278288 , n278289 , n278290 , n278291 , n278292 , n278293 , n278294 , n278295 , 
     n278296 , n278297 , n278298 , n278299 , n278300 , n278301 , n278302 , n278303 , n278304 , n278305 , 
     n278306 , n278307 , n278308 , n278309 , n278310 , n278311 , n278312 , n278313 , n278314 , n278315 , 
     n278316 , n278317 , n278318 , n278319 , n278320 , n278321 , n278322 , n278323 , n278324 , n278325 , 
     n278326 , n278327 , n278328 , n278329 , n278330 , n278331 , n278332 , n278333 , n278334 , n278335 , 
     n278336 , n278337 , n278338 , n278339 , n278340 , n278341 , n278342 , n278343 , n278344 , n278345 , 
     n278346 , n278347 , n278348 , n278349 , n278350 , n278351 , n278352 , n278353 , n278354 , n278355 , 
     n278356 , n278357 , n278358 , n278359 , n278360 , n278361 , n278362 , n278363 , n278364 , n278365 , 
     n278366 , n278367 , n278368 , n278369 , n278370 , n278371 , n278372 , n278373 , n278374 , n278375 , 
     n278376 , n278377 , n278378 , n278379 , n278380 , n278381 , n278382 , n278383 , n278384 , n278385 , 
     n278386 , n278387 , n278388 , n278389 , n278390 , n278391 , n278392 , n278393 , n278394 , n278395 , 
     n278396 , n278397 , n278398 , n278399 , n278400 , n278401 , n278402 , n278403 , n278404 , n278405 , 
     n278406 , n278407 , n278408 , n278409 , n278410 , n278411 , n278412 , n278413 , n278414 , n278415 , 
     n278416 , n278417 , n278418 , n278419 , n278420 , n278421 , n278422 , n278423 , n278424 , n278425 , 
     n278426 , n278427 , n278428 , n278429 , n278430 , n278431 , n278432 , n278433 , n278434 , n278435 , 
     n278436 , n278437 , n278438 , n278439 , n278440 , n278441 , n278442 , n278443 , n278444 , n278445 , 
     n278446 , n278447 , n278448 , n278449 , n278450 , n278451 , n278452 , n278453 , n278454 , n278455 , 
     n278456 , n278457 , n278458 , n278459 , n278460 , n278461 , n278462 , n278463 , n278464 , n278465 , 
     n278466 , n278467 , n278468 , n278469 , n278470 , n278471 , n278472 , n278473 , n278474 , n278475 , 
     n278476 , n278477 , n278478 , n278479 , n278480 , n278481 , n278482 , n278483 , n278484 , n278485 , 
     n278486 , n278487 , n278488 , n278489 , n278490 , n278491 , n278492 , n278493 , n278494 , n278495 , 
     n278496 , n278497 , n278498 , n278499 , n278500 , n278501 , n278502 , n278503 , n278504 , n278505 , 
     n278506 , n278507 , n278508 , n278509 , n278510 , n278511 , n278512 , n278513 , n278514 , n278515 , 
     n278516 , n278517 , n278518 , n278519 , n278520 , n278521 , n278522 , n278523 , n278524 , n278525 , 
     n278526 , n278527 , n278528 , n278529 , n278530 , n278531 , n278532 , n278533 , n278534 , n278535 , 
     n278536 , n278537 , n278538 , n278539 , n278540 , n278541 , n278542 , n278543 , n278544 , n278545 , 
     n278546 , n278547 , n278548 , n278549 , n278550 , n278551 , n278552 , n278553 , n278554 , n278555 , 
     n278556 , n278557 , n278558 , n278559 , n278560 , n278561 , n278562 , n278563 , n278564 , n278565 , 
     n278566 , n278567 , n278568 , n278569 , n278570 , n278571 , n278572 , n278573 , n278574 , n278575 , 
     n278576 , n278577 , n278578 , n278579 , n278580 , n278581 , n278582 , n278583 , n278584 , n278585 , 
     n278586 , n278587 , n278588 , n278589 , n278590 , n278591 , n278592 , n278593 , n278594 , n278595 , 
     n278596 , n278597 , n278598 , n278599 , n278600 , n278601 , n278602 , n278603 , n278604 , n278605 , 
     n278606 , n278607 , n278608 , n278609 , n278610 , n278611 , n278612 , n278613 , n278614 , n278615 , 
     n278616 , n278617 , n278618 , n278619 , n278620 , n278621 , n278622 , n278623 , n278624 , n278625 , 
     n278626 , n278627 , n278628 , n278629 , n278630 , n278631 , n278632 , n278633 , n278634 , n278635 , 
     n278636 , n278637 , n278638 , n278639 , n278640 , n278641 , n278642 , n278643 , n278644 , n278645 , 
     n278646 , n278647 , n278648 , n278649 , n278650 , n278651 , n278652 , n278653 , n278654 , n278655 , 
     n278656 , n278657 , n278658 , n278659 , n278660 , n278661 , n278662 , n278663 , n278664 , n278665 , 
     n278666 , n278667 , n278668 , n278669 , n278670 , n278671 , n278672 , n278673 , n278674 , n278675 , 
     n278676 , n278677 , n278678 , n278679 , n278680 , n278681 , n278682 , n278683 , n278684 , n278685 , 
     n278686 , n278687 , n278688 , n278689 , n278690 , n278691 , n278692 , n278693 , n278694 , n278695 , 
     n278696 , n278697 , n278698 , n278699 , n278700 , n278701 , n278702 , n278703 , n278704 , n278705 , 
     n278706 , n278707 , n278708 , n278709 , n278710 , n278711 , n278712 , n278713 , n278714 , n278715 , 
     n278716 , n278717 , n278718 , n278719 , n278720 , n278721 , n278722 , n278723 , n278724 , n278725 , 
     n278726 , n278727 , n278728 , n278729 , n278730 , n278731 , n278732 , n278733 , n278734 , n278735 , 
     n278736 , n278737 , n278738 , n278739 , n278740 , n278741 , n278742 , n278743 , n278744 , n278745 , 
     n278746 , n278747 , n278748 , n278749 , n278750 , n278751 , n278752 , n278753 , n278754 , n278755 , 
     n278756 , n278757 , n278758 , n278759 , n278760 , n278761 , n278762 , n278763 , n278764 , n278765 , 
     n278766 , n278767 , n278768 , n278769 , n278770 , n278771 , n278772 , n278773 , n278774 , n278775 , 
     n278776 , n278777 , n278778 , n278779 , n278780 , n278781 , n278782 , n278783 , n278784 , n278785 , 
     n278786 , n278787 , n278788 , n278789 , n278790 , n278791 , n278792 , n278793 , n278794 , n278795 , 
     n278796 , n278797 , n278798 , n278799 , n278800 , n278801 , n278802 , n278803 , n278804 , n278805 , 
     n278806 , n278807 , n278808 , n278809 , n278810 , n278811 , n278812 , n278813 , n278814 , n278815 , 
     n278816 , n278817 , n278818 , n278819 , n278820 , n278821 , n278822 , n278823 , n278824 , n278825 , 
     n278826 , n278827 , n278828 , n278829 , n278830 , n278831 , n278832 , n278833 , n278834 , n278835 , 
     n278836 , n278837 , n278838 , n278839 , n278840 , n278841 , n278842 , n278843 , n278844 , n278845 , 
     n278846 , n278847 , n278848 , n278849 , n278850 , n278851 , n278852 , n278853 , n278854 , n278855 , 
     n278856 , n278857 , n278858 , n278859 , n278860 , n278861 , n278862 , n278863 , n278864 , n278865 , 
     n278866 , n278867 , n278868 , n278869 , n278870 , n278871 , n278872 , n278873 , n278874 , n278875 , 
     n278876 , n278877 , n278878 , n278879 , n278880 , n278881 , n278882 , n278883 , n278884 , n278885 , 
     n278886 , n278887 , n278888 , n278889 , n278890 , n278891 , n278892 , n278893 , n278894 , n278895 , 
     n278896 , n278897 , n278898 , n278899 , n278900 , n278901 , n278902 , n278903 , n278904 , n278905 , 
     n278906 , n278907 , n278908 , n278909 , n278910 , n278911 , n278912 , n278913 , n278914 , n278915 , 
     n278916 , n278917 , n278918 , n278919 , n278920 , n278921 , n278922 , n278923 , n278924 , n278925 , 
     n278926 , n278927 , n278928 , n278929 , n278930 , n278931 , n278932 , n278933 , n278934 , n278935 , 
     n278936 , n278937 , n278938 , n278939 , n278940 , n278941 , n278942 , n278943 , n278944 , n278945 , 
     n278946 , n278947 , n278948 , n278949 , n278950 , n278951 , n278952 , n278953 , n278954 , n278955 , 
     n278956 , n278957 , n278958 , n278959 , n278960 , n278961 , n278962 , n278963 , n278964 , n278965 , 
     n278966 , n278967 , n278968 , n278969 , n278970 , n278971 , n278972 , n278973 , n278974 , n278975 , 
     n278976 , n278977 , n278978 , n278979 , n278980 , n278981 , n278982 , n278983 , n278984 , n278985 , 
     n278986 , n278987 , n278988 , n278989 , n278990 , n278991 , n278992 , n278993 , n278994 , n278995 , 
     n278996 , n278997 , n278998 , n278999 , n279000 , n279001 , n279002 , n279003 , n279004 , n279005 , 
     n279006 , n279007 , n279008 , n279009 , n279010 , n279011 , n279012 , n279013 , n279014 , n279015 , 
     n279016 , n279017 , n279018 , n279019 , n279020 , n279021 , n279022 , n279023 , n279024 , n279025 , 
     n279026 , n279027 , n279028 , n279029 , n279030 , n279031 , n279032 , n279033 , n279034 , n279035 , 
     n279036 , n279037 , n279038 , n279039 , n279040 , n279041 , n279042 , n279043 , n279044 , n279045 , 
     n279046 , n279047 , n279048 , n279049 , n279050 , n279051 , n279052 , n279053 , n279054 , n279055 , 
     n279056 , n279057 , n279058 , n279059 , n279060 , n279061 , n279062 , n279063 , n279064 , n279065 , 
     n279066 , n279067 , n279068 , n279069 , n279070 , n279071 , n279072 , n279073 , n279074 , n279075 , 
     n279076 , n279077 , n279078 , n279079 , n279080 , n279081 , n279082 , n279083 , n279084 , n279085 , 
     n279086 , n279087 , n279088 , n279089 , n279090 , n279091 , n279092 , n279093 , n279094 , n279095 , 
     n279096 , n279097 , n279098 , n279099 , n279100 , n279101 , n279102 , n279103 , n279104 , n279105 , 
     n279106 , n279107 , n279108 , n279109 , n279110 , n279111 , n279112 , n279113 , n279114 , n279115 , 
     n279116 , n279117 , n279118 , n279119 , n279120 , n279121 , n279122 , n279123 , n279124 , n279125 , 
     n279126 , n279127 , n279128 , n279129 , n279130 , n279131 , n279132 , n279133 , n279134 , n279135 , 
     n279136 , n279137 , n279138 , n279139 , n279140 , n279141 , n279142 , n279143 , n279144 , n279145 , 
     n279146 , n279147 , n279148 , n279149 , n279150 , n279151 , n279152 , n279153 , n279154 , n279155 , 
     n279156 , n279157 , n279158 , n279159 , n279160 , n279161 , n279162 , n279163 , n279164 , n279165 , 
     n279166 , n279167 , n279168 , n279169 , n279170 , n279171 , n279172 , n279173 , n279174 , n279175 , 
     n279176 , n279177 , n279178 , n279179 , n279180 , n279181 , n279182 , n279183 , n279184 , n279185 , 
     n279186 , n279187 , n279188 , n279189 , n279190 , n279191 , n279192 , n279193 , n279194 , n279195 , 
     n279196 , n279197 , n279198 , n279199 , n279200 , n279201 , n279202 , n279203 , n279204 , n279205 , 
     n279206 , n279207 , n279208 , n279209 , n279210 , n279211 , n279212 , n279213 , n279214 , n279215 , 
     n279216 , n279217 , n279218 , n279219 , n279220 , n279221 , n279222 , n279223 , n279224 , n279225 , 
     n279226 , n279227 , n279228 , n279229 , n279230 , n279231 , n279232 , n279233 , n279234 , n279235 , 
     n279236 , n279237 , n279238 , n279239 , n279240 , n279241 , n279242 , n279243 , n279244 , n279245 , 
     n279246 , n279247 , n279248 , n279249 , n279250 , n279251 , n279252 , n279253 , n279254 , n279255 , 
     n279256 , n279257 , n279258 , n279259 , n279260 , n279261 , n279262 , n279263 , n279264 , n279265 , 
     n279266 , n279267 , n279268 , n279269 , n279270 , n279271 , n279272 , n279273 , n279274 , n279275 , 
     n279276 , n279277 , n279278 , n279279 , n279280 , n279281 , n279282 , n279283 , n279284 , n279285 , 
     n279286 , n279287 , n279288 , n279289 , n279290 , n279291 , n279292 , n279293 , n279294 , n279295 , 
     n279296 , n279297 , n279298 , n279299 , n279300 , n279301 , n279302 , n279303 , n279304 , n279305 , 
     n279306 , n279307 , n279308 , n279309 , n279310 , n279311 , n279312 , n279313 , n279314 , n279315 , 
     n279316 , n279317 , n279318 , n279319 , n279320 , n279321 , n279322 , n279323 , n279324 , n279325 , 
     n279326 , n279327 , n279328 , n279329 , n279330 , n279331 , n279332 , n279333 , n279334 , n279335 , 
     n279336 , n279337 , n279338 , n279339 , n279340 , n279341 , n279342 , n279343 , n279344 , n279345 , 
     n279346 , n279347 , n279348 , n279349 , n279350 , n279351 , n279352 , n279353 , n279354 , n279355 , 
     n279356 , n279357 , n279358 , n279359 , n279360 , n279361 , n279362 , n279363 , n279364 , n279365 , 
     n279366 , n279367 , n279368 , n279369 , n279370 , n279371 , n279372 , n279373 , n279374 , n279375 , 
     n279376 , n279377 , n279378 , n279379 , n279380 , n279381 , n279382 , n279383 , n279384 , n279385 , 
     n279386 , n279387 , n279388 , n279389 , n279390 , n279391 , n279392 , n279393 , n279394 , n279395 , 
     n279396 , n279397 , n279398 , n279399 , n279400 , n279401 , n279402 , n279403 , n279404 , n279405 , 
     n279406 , n279407 , n279408 , n279409 , n279410 , n279411 , n279412 , n279413 , n279414 , n279415 , 
     n279416 , n279417 , n279418 , n279419 , n279420 , n279421 , n279422 , n279423 , n279424 , n279425 , 
     n279426 , n279427 , n279428 , n279429 , n279430 , n279431 , n279432 , n279433 , n279434 , n279435 , 
     n279436 , n279437 , n279438 , n279439 , n279440 , n279441 , n279442 , n279443 , n279444 , n279445 , 
     n279446 , n279447 , n279448 , n279449 , n279450 , n279451 , n279452 , n279453 , n279454 , n279455 , 
     n279456 , n279457 , n279458 , n279459 , n279460 , n279461 , n279462 , n279463 , n279464 , n279465 , 
     n279466 , n279467 , n279468 , n279469 , n279470 , n279471 , n279472 , n279473 , n279474 , n279475 , 
     n279476 , n279477 , n279478 , n279479 , n279480 , n279481 , n279482 , n279483 , n279484 , n279485 , 
     n279486 , n279487 , n279488 , n279489 , n279490 , n279491 , n279492 , n279493 , n279494 , n279495 , 
     n279496 , n279497 , n279498 , n279499 , n279500 , n279501 , n279502 , n279503 , n279504 , n279505 , 
     n279506 , n279507 , n279508 , n279509 , n279510 , n279511 , n279512 , n279513 , n279514 , n279515 , 
     n279516 , n279517 , n279518 , n279519 , n279520 , n279521 , n279522 , n279523 , n279524 , n279525 , 
     n279526 , n279527 , n279528 , n279529 , n279530 , n279531 , n279532 , n279533 , n279534 , n279535 , 
     n279536 , n279537 , n279538 , n279539 , n279540 , n279541 , n279542 , n279543 , n279544 , n279545 , 
     n279546 , n279547 , n279548 , n279549 , n279550 , n279551 , n279552 , n279553 , n279554 , n279555 , 
     n279556 , n279557 , n279558 , n279559 , n279560 , n279561 , n279562 , n279563 , n279564 , n279565 , 
     n279566 , n279567 , n279568 , n279569 , n279570 , n279571 , n279572 , n279573 , n279574 , n279575 , 
     n279576 , n279577 , n279578 , n279579 , n279580 , n279581 , n279582 , n279583 , n279584 , n279585 , 
     n279586 , n279587 , n279588 , n279589 , n279590 , n279591 , n279592 , n279593 , n279594 , n279595 , 
     n279596 , n279597 , n279598 , n279599 , n279600 , n279601 , n279602 , n279603 , n279604 , n279605 , 
     n279606 , n279607 , n279608 , n279609 , n279610 , n279611 , n279612 , n279613 , n279614 , n279615 , 
     n279616 , n279617 , n279618 , n279619 , n279620 , n279621 , n279622 , n279623 , n279624 , n279625 , 
     n279626 , n279627 , n279628 , n279629 , n279630 , n279631 , n279632 , n279633 , n279634 , n279635 , 
     n279636 , n279637 , n279638 , n279639 , n279640 , n279641 , n279642 , n279643 , n279644 , n279645 , 
     n279646 , n279647 , n279648 , n279649 , n279650 , n279651 , n279652 , n279653 , n279654 , n279655 , 
     n279656 , n279657 , n279658 , n279659 , n279660 , n279661 , n279662 , n279663 , n279664 , n279665 , 
     n279666 , n279667 , n279668 , n279669 , n279670 , n279671 , n279672 , n279673 , n279674 , n279675 , 
     n279676 , n279677 , n279678 , n279679 , n279680 , n279681 , n279682 , n279683 , n279684 , n279685 , 
     n279686 , n279687 , n279688 , n279689 , n279690 , n279691 , n279692 , n279693 , n279694 , n279695 , 
     n279696 , n279697 , n279698 , n279699 , n279700 , n279701 , n279702 , n279703 , n279704 , n279705 , 
     n279706 , n279707 , n279708 , n279709 , n279710 , n279711 , n279712 , n279713 , n279714 , n279715 , 
     n279716 , n279717 , n279718 , n279719 , n279720 , n279721 , n279722 , n279723 , n279724 , n279725 , 
     n279726 , n279727 , n279728 , n279729 , n279730 , n279731 , n279732 , n279733 , n279734 , n279735 , 
     n279736 , n279737 , n279738 , n279739 , n279740 , n279741 , n279742 , n279743 , n279744 , n279745 , 
     n279746 , n279747 , n279748 , n279749 , n279750 , n279751 , n279752 , n279753 , n279754 , n279755 , 
     n279756 , n279757 , n279758 , n279759 , n279760 , n279761 , n279762 , n279763 , n279764 , n279765 , 
     n279766 , n279767 , n279768 , n279769 , n279770 , n279771 , n279772 , n279773 , n279774 , n279775 , 
     n279776 , n279777 , n279778 , n279779 , n279780 , n279781 , n279782 , n279783 , n279784 , n279785 , 
     n279786 , n279787 , n279788 , n279789 , n279790 , n279791 , n279792 , n279793 , n279794 , n279795 , 
     n279796 , n279797 , n279798 , n279799 , n279800 , n279801 , n279802 , n279803 , n279804 , n279805 , 
     n279806 , n279807 , n279808 , n279809 , n279810 , n279811 , n279812 , n279813 , n279814 , n279815 , 
     n279816 , n279817 , n279818 , n279819 , n279820 , n279821 , n279822 , n279823 , n279824 , n279825 , 
     n279826 , n279827 , n279828 , n279829 , n279830 , n279831 , n279832 , n279833 , n279834 , n279835 , 
     n279836 , n279837 , n279838 , n279839 , n279840 , n279841 , n279842 , n279843 , n279844 , n279845 , 
     n279846 , n279847 , n279848 , n279849 , n279850 , n279851 , n279852 , n279853 , n279854 , n279855 , 
     n279856 , n279857 , n279858 , n279859 , n279860 , n279861 , n279862 , n279863 , n279864 , n279865 , 
     n279866 , n279867 , n279868 , n279869 , n279870 , n279871 , n279872 , n279873 , n279874 , n279875 , 
     n279876 , n279877 , n279878 , n279879 , n279880 , n279881 , n279882 , n279883 , n279884 , n279885 , 
     n279886 , n279887 , n279888 , n279889 , n279890 , n279891 , n279892 , n279893 , n279894 , n279895 , 
     n279896 , n279897 , n279898 , n279899 , n279900 , n279901 , n279902 , n279903 , n279904 , n279905 , 
     n279906 , n279907 , n279908 , n279909 , n279910 , n279911 , n279912 , n279913 , n279914 , n279915 , 
     n279916 , n279917 , n279918 , n279919 , n279920 , n279921 , n279922 , n279923 , n279924 , n279925 , 
     n279926 , n279927 , n279928 , n279929 , n279930 , n279931 , n279932 , n279933 , n279934 , n279935 , 
     n279936 , n279937 , n279938 , n279939 , n279940 , n279941 , n279942 , n279943 , n279944 , n279945 , 
     n279946 , n279947 , n279948 , n279949 , n279950 , n279951 , n279952 , n279953 , n279954 , n279955 , 
     n279956 , n279957 , n279958 , n279959 , n279960 , n279961 , n279962 , n279963 , n279964 , n279965 , 
     n279966 , n279967 , n279968 , n279969 , n279970 , n279971 , n279972 , n279973 , n279974 , n279975 , 
     n279976 , n279977 , n279978 , n279979 , n279980 , n279981 , n279982 , n279983 , n279984 , n279985 , 
     n279986 , n279987 , n279988 , n279989 , n279990 , n279991 , n279992 , n279993 , n279994 , n279995 , 
     n279996 , n279997 , n279998 , n279999 , n280000 , n280001 , n280002 , n280003 , n280004 , n280005 , 
     n280006 , n280007 , n280008 , n280009 , n280010 , n280011 , n280012 , n280013 , n280014 , n280015 , 
     n280016 , n280017 , n280018 , n280019 , n280020 , n280021 , n280022 , n280023 , n280024 , n280025 , 
     n280026 , n280027 , n280028 , n280029 , n280030 , n280031 , n280032 , n280033 , n280034 , n280035 , 
     n280036 , n280037 , n280038 , n280039 , n280040 , n280041 , n280042 , n280043 , n280044 , n280045 , 
     n280046 , n280047 , n280048 , n280049 , n280050 , n280051 , n280052 , n280053 , n280054 , n280055 , 
     n280056 , n280057 , n280058 , n280059 , n280060 , n280061 , n280062 , n280063 , n280064 , n280065 , 
     n280066 , n280067 , n280068 , n280069 , n280070 , n280071 , n280072 , n280073 , n280074 , n280075 , 
     n280076 , n280077 , n280078 , n280079 , n280080 , n280081 , n280082 , n280083 , n280084 , n280085 , 
     n280086 , n280087 , n280088 , n280089 , n280090 , n280091 , n280092 , n280093 , n280094 , n280095 , 
     n280096 , n280097 , n280098 , n280099 , n280100 , n280101 , n280102 , n280103 , n280104 , n280105 , 
     n280106 , n280107 , n280108 , n280109 , n280110 , n280111 , n280112 , n280113 , n280114 , n280115 , 
     n280116 , n280117 , n280118 , n280119 , n280120 , n280121 , n280122 , n280123 , n280124 , n280125 , 
     n280126 , n280127 , n280128 , n280129 , n280130 , n280131 , n280132 , n280133 , n280134 , n280135 , 
     n280136 , n280137 , n280138 , n280139 , n280140 , n280141 , n280142 , n280143 , n280144 , n280145 , 
     n280146 , n280147 , n280148 , n280149 , n280150 , n280151 , n280152 , n280153 , n280154 , n280155 , 
     n280156 , n280157 , n280158 , n280159 , n280160 , n280161 , n280162 , n280163 , n280164 , n280165 , 
     n280166 , n280167 , n280168 , n280169 , n280170 , n280171 , n280172 , n280173 , n280174 , n280175 , 
     n280176 , n280177 , n280178 , n280179 , n280180 , n280181 , n280182 , n280183 , n280184 , n280185 , 
     n280186 , n280187 , n280188 , n280189 , n280190 , n280191 , n280192 , n280193 , n280194 , n280195 , 
     n280196 , n280197 , n280198 , n280199 , n280200 , n280201 , n280202 , n280203 , n280204 , n280205 , 
     n280206 , n280207 , n280208 , n280209 , n280210 , n280211 , n280212 , n280213 , n280214 , n280215 , 
     n280216 , n280217 , n280218 , n280219 , n280220 , n280221 , n280222 , n280223 , n280224 , n280225 , 
     n280226 , n280227 , n280228 , n280229 , n280230 , n280231 , n280232 , n280233 , n280234 , n280235 , 
     n280236 , n280237 , n280238 , n280239 , n280240 , n280241 , n280242 , n280243 , n280244 , n280245 , 
     n280246 , n280247 , n280248 , n280249 , n280250 , n280251 , n280252 , n280253 , n280254 , n280255 , 
     n280256 , n280257 , n280258 , n280259 , n280260 , n280261 , n280262 , n280263 , n280264 , n280265 , 
     n280266 , n280267 , n280268 , n280269 , n280270 , n280271 , n280272 , n280273 , n280274 , n280275 , 
     n280276 , n280277 , n280278 , n280279 , n280280 , n280281 , n280282 , n280283 , n280284 , n280285 , 
     n280286 , n280287 , n280288 , n280289 , n280290 , n280291 , n280292 , n280293 , n280294 , n280295 , 
     n280296 , n280297 , n280298 , n280299 , n280300 , n280301 , n280302 , n280303 , n280304 , n280305 , 
     n280306 , n280307 , n280308 , n280309 , n280310 , n280311 , n280312 , n280313 , n280314 , n280315 , 
     n280316 , n280317 , n280318 , n280319 , n280320 , n280321 , n280322 , n280323 , n280324 , n280325 , 
     n280326 , n280327 , n280328 , n280329 , n280330 , n280331 , n280332 , n280333 , n280334 , n280335 , 
     n280336 , n280337 , n280338 , n280339 , n280340 , n280341 , n280342 , n280343 , n280344 , n280345 , 
     n280346 , n280347 , n280348 , n280349 , n280350 , n280351 , n280352 , n280353 , n280354 , n280355 , 
     n280356 , n280357 , n280358 , n280359 , n280360 , n280361 , n280362 , n280363 , n280364 , n280365 , 
     n280366 , n280367 , n280368 , n280369 , n280370 , n280371 , n280372 , n280373 , n280374 , n280375 , 
     n280376 , n280377 , n280378 , n280379 , n280380 , n280381 , n280382 , n280383 , n280384 , n280385 , 
     n280386 , n280387 , n280388 , n280389 , n280390 , n280391 , n280392 , n280393 , n280394 , n280395 , 
     n280396 , n280397 , n280398 , n280399 , n280400 , n280401 , n280402 , n280403 , n280404 , n280405 , 
     n280406 , n280407 , n280408 , n280409 , n280410 , n280411 , n280412 , n280413 , n280414 , n280415 , 
     n280416 , n280417 , n280418 , n280419 , n280420 , n280421 , n280422 , n280423 , n280424 , n280425 , 
     n280426 , n280427 , n280428 , n280429 , n280430 , n280431 , n280432 , n280433 , n280434 , n280435 , 
     n280436 , n280437 , n280438 , n280439 , n280440 , n280441 , n280442 , n280443 , n280444 , n280445 , 
     n280446 , n280447 , n280448 , n280449 , n280450 , n280451 , n280452 , n280453 , n280454 , n280455 , 
     n280456 , n280457 , n280458 , n280459 , n280460 , n280461 , n280462 , n280463 , n280464 , n280465 , 
     n280466 , n280467 , n280468 , n280469 , n280470 , n280471 , n280472 , n280473 , n280474 , n280475 , 
     n280476 , n280477 , n280478 , n280479 , n280480 , n280481 , n280482 , n280483 , n280484 , n280485 , 
     n280486 , n280487 , n280488 , n280489 , n280490 , n280491 , n280492 , n280493 , n280494 , n280495 , 
     n280496 , n280497 , n280498 , n280499 , n280500 , n280501 , n280502 , n280503 , n280504 , n280505 , 
     n280506 , n280507 , n280508 , n280509 , n280510 , n280511 , n280512 , n280513 , n280514 , n280515 , 
     n280516 , n280517 , n280518 , n280519 , n280520 , n280521 , n280522 , n280523 , n280524 , n280525 , 
     n280526 , n280527 , n280528 , n280529 , n280530 , n280531 , n280532 , n280533 , n280534 , n280535 , 
     n280536 , n280537 , n280538 , n280539 , n280540 , n280541 , n280542 , n280543 , n280544 , n280545 , 
     n280546 , n280547 , n280548 , n280549 , n280550 , n280551 , n280552 , n280553 , n280554 , n280555 , 
     n280556 , n280557 , n280558 , n280559 , n280560 , n280561 , n280562 , n280563 , n280564 , n280565 , 
     n280566 , n280567 , n280568 , n280569 , n280570 , n280571 , n280572 , n280573 , n280574 , n280575 , 
     n280576 , n280577 , n280578 , n280579 , n280580 , n280581 , n280582 , n280583 , n280584 , n280585 , 
     n280586 , n280587 , n280588 , n280589 , n280590 , n280591 , n280592 , n280593 , n280594 , n280595 , 
     n280596 , n280597 , n280598 , n280599 , n280600 , n280601 , n280602 , n280603 , n280604 , n280605 , 
     n280606 , n280607 , n280608 , n280609 , n280610 , n280611 , n280612 , n280613 , n280614 , n280615 , 
     n280616 , n280617 , n280618 , n280619 , n280620 , n280621 , n280622 , n280623 , n280624 , n280625 , 
     n280626 , n280627 , n280628 , n280629 , n280630 , n280631 , n280632 , n280633 , n280634 , n280635 , 
     n280636 , n280637 , n280638 , n280639 , n280640 , n280641 , n280642 , n280643 , n280644 , n280645 , 
     n280646 , n280647 , n280648 , n280649 , n280650 , n280651 , n280652 , n280653 , n280654 , n280655 , 
     n280656 , n280657 , n280658 , n280659 , n280660 , n280661 , n280662 , n280663 , n280664 , n280665 , 
     n280666 , n280667 , n280668 , n280669 , n280670 , n280671 , n280672 , n280673 , n280674 , n280675 , 
     n280676 , n280677 , n280678 , n280679 , n280680 , n280681 , n280682 , n280683 , n280684 , n280685 , 
     n280686 , n280687 , n280688 , n280689 , n280690 , n280691 , n280692 , n280693 , n280694 , n280695 , 
     n280696 , n280697 , n280698 , n280699 , n280700 , n280701 , n280702 , n280703 , n280704 , n280705 , 
     n280706 , n280707 , n280708 , n280709 , n280710 , n280711 , n280712 , n280713 , n280714 , n280715 , 
     n280716 , n280717 , n280718 , n280719 , n280720 , n280721 , n280722 , n280723 , n280724 , n280725 , 
     n280726 , n280727 , n280728 , n280729 , n280730 , n280731 , n280732 , n280733 , n280734 , n280735 , 
     n280736 , n280737 , n280738 , n280739 , n280740 , n280741 , n280742 , n280743 , n280744 , n280745 , 
     n280746 , n280747 , n280748 , n280749 , n280750 , n280751 , n280752 , n280753 , n280754 , n280755 , 
     n280756 , n280757 , n280758 , n280759 , n280760 , n280761 , n280762 , n280763 , n280764 , n280765 , 
     n280766 , n280767 , n280768 , n280769 , n280770 , n280771 , n280772 , n280773 , n280774 , n280775 , 
     n280776 , n280777 , n280778 , n280779 , n280780 , n280781 , n280782 , n280783 , n280784 , n280785 , 
     n280786 , n280787 , n280788 , n280789 , n280790 , n280791 , n280792 , n280793 , n280794 , n280795 , 
     n280796 , n280797 , n280798 , n280799 , n280800 , n280801 , n280802 , n280803 , n280804 , n280805 , 
     n280806 , n280807 , n280808 , n280809 , n280810 , n280811 , n280812 , n280813 , n280814 , n280815 , 
     n280816 , n280817 , n280818 , n280819 , n280820 , n280821 , n280822 , n280823 , n280824 , n280825 , 
     n280826 , n280827 , n280828 , n280829 , n280830 , n280831 , n280832 , n280833 , n280834 , n280835 , 
     n280836 , n280837 , n280838 , n280839 , n280840 , n280841 , n280842 , n280843 , n280844 , n280845 , 
     n280846 , n280847 , n280848 , n280849 , n280850 , n280851 , n280852 , n280853 , n280854 , n280855 , 
     n280856 , n280857 , n280858 , n280859 , n280860 , n280861 , n280862 , n280863 , n280864 , n280865 , 
     n280866 , n280867 , n280868 , n280869 , n280870 , n280871 , n280872 , n280873 , n280874 , n280875 , 
     n280876 , n280877 , n280878 , n280879 , n280880 , n280881 , n280882 , n280883 , n280884 , n280885 , 
     n280886 , n280887 , n280888 , n280889 , n280890 , n280891 , n280892 , n280893 , n280894 , n280895 , 
     n280896 , n280897 , n280898 , n280899 , n280900 , n280901 , n280902 , n280903 , n280904 , n280905 , 
     n280906 , n280907 , n280908 , n280909 , n280910 , n280911 , n280912 , n280913 , n280914 , n280915 , 
     n280916 , n280917 , n280918 , n280919 , n280920 , n280921 , n280922 , n280923 , n280924 , n280925 , 
     n280926 , n280927 , n280928 , n280929 , n280930 , n280931 , n280932 , n280933 , n280934 , n280935 , 
     n280936 , n280937 , n280938 , n280939 , n280940 , n280941 , n280942 , n280943 , n280944 , n280945 , 
     n280946 , n280947 , n280948 , n280949 , n280950 , n280951 , n280952 , n280953 , n280954 , n280955 , 
     n280956 , n280957 , n280958 , n280959 , n280960 , n280961 , n280962 , n280963 , n280964 , n280965 , 
     n280966 , n280967 , n280968 , n280969 , n280970 , n280971 , n280972 , n280973 , n280974 , n280975 , 
     n280976 , n280977 , n280978 , n280979 , n280980 , n280981 , n280982 , n280983 , n280984 , n280985 , 
     n280986 , n280987 , n280988 , n280989 , n280990 , n280991 , n280992 , n280993 , n280994 , n280995 , 
     n280996 , n280997 , n280998 , n280999 , n281000 , n281001 , n281002 , n281003 , n281004 , n281005 , 
     n281006 , n281007 , n281008 , n281009 , n281010 , n281011 , n281012 , n281013 , n281014 , n281015 , 
     n281016 , n281017 , n281018 , n281019 , n281020 , n281021 , n281022 , n281023 , n281024 , n281025 , 
     n281026 , n281027 , n281028 , n281029 , n281030 , n281031 , n281032 , n281033 , n281034 , n281035 , 
     n281036 , n281037 , n281038 , n281039 , n281040 , n281041 , n281042 , n281043 , n281044 , n281045 , 
     n281046 , n281047 , n281048 , n281049 , n281050 , n281051 , n281052 , n281053 , n281054 , n281055 , 
     n281056 , n281057 , n281058 , n281059 , n281060 , n281061 , n281062 , n281063 , n281064 , n281065 , 
     n281066 , n281067 , n281068 , n281069 , n281070 , n281071 , n281072 , n281073 , n281074 , n281075 , 
     n281076 , n281077 , n281078 , n281079 , n281080 , n281081 , n281082 , n281083 , n281084 , n281085 , 
     n281086 , n281087 , n281088 , n281089 , n281090 , n281091 , n281092 , n281093 , n281094 , n281095 , 
     n281096 , n281097 , n281098 , n281099 , n281100 , n281101 , n281102 , n281103 , n281104 , n281105 , 
     n281106 , n281107 , n281108 , n281109 , n281110 , n281111 , n281112 , n281113 , n281114 , n281115 , 
     n281116 , n281117 , n281118 , n281119 , n281120 , n281121 , n281122 , n281123 , n281124 , n281125 , 
     n281126 , n281127 , n281128 , n281129 , n281130 , n281131 , n281132 , n281133 , n281134 , n281135 , 
     n281136 , n281137 , n281138 , n281139 , n281140 , n281141 , n281142 , n281143 , n281144 , n281145 , 
     n281146 , n281147 , n281148 , n281149 , n281150 , n281151 , n281152 , n281153 , n281154 , n281155 , 
     n281156 , n281157 , n281158 , n281159 , n281160 , n281161 , n281162 , n281163 , n281164 , n281165 , 
     n281166 , n281167 , n281168 , n281169 , n281170 , n281171 , n281172 , n281173 , n281174 , n281175 , 
     n281176 , n281177 , n281178 , n281179 , n281180 , n281181 , n281182 , n281183 , n281184 , n281185 , 
     n281186 , n281187 , n281188 , n281189 , n281190 , n281191 , n281192 , n281193 , n281194 , n281195 , 
     n281196 , n281197 , n281198 , n281199 , n281200 , n281201 , n281202 , n281203 , n281204 , n281205 , 
     n281206 , n281207 , n281208 , n281209 , n281210 , n281211 , n281212 , n281213 , n281214 , n281215 , 
     n281216 , n281217 , n281218 , n281219 , n281220 , n281221 , n281222 , n281223 , n281224 , n281225 , 
     n281226 , n281227 , n281228 , n281229 , n281230 , n281231 , n281232 , n281233 , n281234 , n281235 , 
     n281236 , n281237 , n281238 , n281239 , n281240 , n281241 , n281242 , n281243 , n281244 , n281245 , 
     n281246 , n281247 , n281248 , n281249 , n281250 , n281251 , n281252 , n281253 , n281254 , n281255 , 
     n281256 , n281257 , n281258 , n281259 , n281260 , n281261 , n281262 , n281263 , n281264 , n281265 , 
     n281266 , n281267 , n281268 , n281269 , n281270 , n281271 , n281272 , n281273 , n281274 , n281275 , 
     n281276 , n281277 , n281278 , n281279 , n281280 , n281281 , n281282 , n281283 , n281284 , n281285 , 
     n281286 , n281287 , n281288 , n281289 , n281290 , n281291 , n281292 , n281293 , n281294 , n281295 , 
     n281296 , n281297 , n281298 , n281299 , n281300 , n281301 , n281302 , n281303 , n281304 , n281305 , 
     n281306 , n281307 , n281308 , n281309 , n281310 , n281311 , n281312 , n281313 , n281314 , n281315 , 
     n281316 , n281317 , n281318 , n281319 , n281320 , n281321 , n281322 , n281323 , n281324 , n281325 , 
     n281326 , n281327 , n281328 , n281329 , n281330 , n281331 , n281332 , n281333 , n281334 , n281335 , 
     n281336 , n281337 , n281338 , n281339 , n281340 , n281341 , n281342 , n281343 , n281344 , n281345 , 
     n281346 , n281347 , n281348 , n281349 , n281350 , n281351 , n281352 , n281353 , n281354 , n281355 , 
     n281356 , n281357 , n281358 , n281359 , n281360 , n281361 , n281362 , n281363 , n281364 , n281365 , 
     n281366 , n281367 , n281368 , n281369 , n281370 , n281371 , n281372 , n281373 , n281374 , n281375 , 
     n281376 , n281377 , n281378 , n281379 , n281380 , n281381 , n281382 , n281383 , n281384 , n281385 , 
     n281386 , n281387 , n281388 , n281389 , n281390 , n281391 , n281392 , n281393 , n281394 , n281395 , 
     n281396 , n281397 , n281398 , n281399 , n281400 , n281401 , n281402 , n281403 , n281404 , n281405 , 
     n281406 , n281407 , n281408 , n281409 , n281410 , n281411 , n281412 , n281413 , n281414 , n281415 , 
     n281416 , n281417 , n281418 , n281419 , n281420 , n281421 , n281422 , n281423 , n281424 , n281425 , 
     n281426 , n281427 , n281428 , n281429 , n281430 , n281431 , n281432 , n281433 , n281434 , n281435 , 
     n281436 , n281437 , n281438 , n281439 , n281440 , n281441 , n281442 , n281443 , n281444 , n281445 , 
     n281446 , n281447 , n281448 , n281449 , n281450 , n281451 , n281452 , n281453 , n281454 , n281455 , 
     n281456 , n281457 , n281458 , n281459 , n281460 , n281461 , n281462 , n281463 , n281464 , n281465 , 
     n281466 , n281467 , n281468 , n281469 , n281470 , n281471 , n281472 , n281473 , n281474 , n281475 , 
     n281476 , n281477 , n281478 , n281479 , n281480 , n281481 , n281482 , n281483 , n281484 , n281485 , 
     n281486 , n281487 , n281488 , n281489 , n281490 , n281491 , n281492 , n281493 , n281494 , n281495 , 
     n281496 , n281497 , n281498 , n281499 , n281500 , n281501 , n281502 , n281503 , n281504 , n281505 , 
     n281506 , n281507 , n281508 , n281509 , n281510 , n281511 , n281512 , n281513 , n281514 , n281515 , 
     n281516 , n281517 , n281518 , n281519 , n281520 , n281521 , n281522 , n281523 , n281524 , n281525 , 
     n281526 , n281527 , n281528 , n281529 , n281530 , n281531 , n281532 , n281533 , n281534 , n281535 , 
     n281536 , n281537 , n281538 , n281539 , n281540 , n281541 , n281542 , n281543 , n281544 , n281545 , 
     n281546 , n281547 , n281548 , n281549 , n281550 , n281551 , n281552 , n281553 , n281554 , n281555 , 
     n281556 , n281557 , n281558 , n281559 , n281560 , n281561 , n281562 , n281563 , n281564 , n281565 , 
     n281566 , n281567 , n281568 , n281569 , n281570 , n281571 , n281572 , n281573 , n281574 , n281575 , 
     n281576 , n281577 , n281578 , n281579 , n281580 , n281581 , n281582 , n281583 , n281584 , n281585 , 
     n281586 , n281587 , n281588 , n281589 , n281590 , n281591 , n281592 , n281593 , n281594 , n281595 , 
     n281596 , n281597 , n281598 , n281599 , n281600 , n281601 , n281602 , n281603 , n281604 , n281605 , 
     n281606 , n281607 , n281608 , n281609 , n281610 , n281611 , n281612 , n281613 , n281614 , n281615 , 
     n281616 , n281617 , n281618 , n281619 , n281620 , n281621 , n281622 , n281623 , n281624 , n281625 , 
     n281626 , n281627 , n281628 , n281629 , n281630 , n281631 , n281632 , n281633 , n281634 , n281635 , 
     n281636 , n281637 , n281638 , n281639 , n281640 , n281641 , n281642 , n281643 , n281644 , n281645 , 
     n281646 , n281647 , n281648 , n281649 , n281650 , n281651 , n281652 , n281653 , n281654 , n281655 , 
     n281656 , n281657 , n281658 , n281659 , n281660 , n281661 , n281662 , n281663 , n281664 , n281665 , 
     n281666 , n281667 , n281668 , n281669 , n281670 , n281671 , n281672 , n281673 , n281674 , n281675 , 
     n281676 , n281677 , n281678 , n281679 , n281680 , n281681 , n281682 , n281683 , n281684 , n281685 , 
     n281686 , n281687 , n281688 , n281689 , n281690 , n281691 , n281692 , n281693 , n281694 , n281695 , 
     n281696 , n281697 , n281698 , n281699 , n281700 , n281701 , n281702 , n281703 , n281704 , n281705 , 
     n281706 , n281707 , n281708 , n281709 , n281710 , n281711 , n281712 , n281713 , n281714 , n281715 , 
     n281716 , n281717 , n281718 , n281719 , n281720 , n281721 , n281722 , n281723 , n281724 , n281725 , 
     n281726 , n281727 , n281728 , n281729 , n281730 , n281731 , n281732 , n281733 , n281734 , n281735 , 
     n281736 , n281737 , n281738 , n281739 , n281740 , n281741 , n281742 , n281743 , n281744 , n281745 , 
     n281746 , n281747 , n281748 , n281749 , n281750 , n281751 , n281752 , n281753 , n281754 , n281755 , 
     n281756 , n281757 , n281758 , n281759 , n281760 , n281761 , n281762 , n281763 , n281764 , n281765 , 
     n281766 , n281767 , n281768 , n281769 , n281770 , n281771 , n281772 , n281773 , n281774 , n281775 , 
     n281776 , n281777 , n281778 , n281779 , n281780 , n281781 , n281782 , n281783 , n281784 , n281785 , 
     n281786 , n281787 , n281788 , n281789 , n281790 , n281791 , n281792 , n281793 , n281794 , n281795 , 
     n281796 , n281797 , n281798 , n281799 , n281800 , n281801 , n281802 , n281803 , n281804 , n281805 , 
     n281806 , n281807 , n281808 , n281809 , n281810 , n281811 , n281812 , n281813 , n281814 , n281815 , 
     n281816 , n281817 , n281818 , n281819 , n281820 , n281821 , n281822 , n281823 , n281824 , n281825 , 
     n281826 , n281827 , n281828 , n281829 , n281830 , n281831 , n281832 , n281833 , n281834 , n281835 , 
     n281836 , n281837 , n281838 , n281839 , n281840 , n281841 , n281842 , n281843 , n281844 , n281845 , 
     n281846 , n281847 , n281848 , n281849 , n281850 , n281851 , n281852 , n281853 , n281854 , n281855 , 
     n281856 , n281857 , n281858 , n281859 , n281860 , n281861 , n281862 , n281863 , n281864 , n281865 , 
     n281866 , n281867 , n281868 , n281869 , n281870 , n281871 , n281872 , n281873 , n281874 , n281875 , 
     n281876 , n281877 , n281878 , n281879 , n281880 , n281881 , n281882 , n281883 , n281884 , n281885 , 
     n281886 , n281887 , n281888 , n281889 , n281890 , n281891 , n281892 , n281893 , n281894 , n281895 , 
     n281896 , n281897 , n281898 , n281899 , n281900 , n281901 , n281902 , n281903 , n281904 , n281905 , 
     n281906 , n281907 , n281908 , n281909 , n281910 , n281911 , n281912 , n281913 , n281914 , n281915 , 
     n281916 , n281917 , n281918 , n281919 , n281920 , n281921 , n281922 , n281923 , n281924 , n281925 , 
     n281926 , n281927 , n281928 , n281929 , n281930 , n281931 , n281932 , n281933 , n281934 , n281935 , 
     n281936 , n281937 , n281938 , n281939 , n281940 , n281941 , n281942 , n281943 , n281944 , n281945 , 
     n281946 , n281947 , n281948 , n281949 , n281950 , n281951 , n281952 , n281953 , n281954 , n281955 , 
     n281956 , n281957 , n281958 , n281959 , n281960 , n281961 , n281962 , n281963 , n281964 , n281965 , 
     n281966 , n281967 , n281968 , n281969 , n281970 , n281971 , n281972 , n281973 , n281974 , n281975 , 
     n281976 , n281977 , n281978 , n281979 , n281980 , n281981 , n281982 , n281983 , n281984 , n281985 , 
     n281986 , n281987 , n281988 , n281989 , n281990 , n281991 , n281992 , n281993 , n281994 , n281995 , 
     n281996 , n281997 , n281998 , n281999 , n282000 , n282001 , n282002 , n282003 , n282004 , n282005 , 
     n282006 , n282007 , n282008 , n282009 , n282010 , n282011 , n282012 , n282013 , n282014 , n282015 , 
     n282016 , n282017 , n282018 , n282019 , n282020 , n282021 , n282022 , n282023 , n282024 , n282025 , 
     n282026 , n282027 , n282028 , n282029 , n282030 , n282031 , n282032 , n282033 , n282034 , n282035 , 
     n282036 , n282037 , n282038 , n282039 , n282040 , n282041 , n282042 , n282043 , n282044 , n282045 , 
     n282046 , n282047 , n282048 , n282049 , n282050 , n282051 , n282052 , n282053 , n282054 , n282055 , 
     n282056 , n282057 , n282058 , n282059 , n282060 , n282061 , n282062 , n282063 , n282064 , n282065 , 
     n282066 , n282067 , n282068 , n282069 , n282070 , n282071 , n282072 , n282073 , n282074 , n282075 , 
     n282076 , n282077 , n282078 , n282079 , n282080 , n282081 , n282082 , n282083 , n282084 , n282085 , 
     n282086 , n282087 , n282088 , n282089 , n282090 , n282091 , n282092 , n282093 , n282094 , n282095 , 
     n282096 , n282097 , n282098 , n282099 , n282100 , n282101 , n282102 , n282103 , n282104 , n282105 , 
     n282106 , n282107 , n282108 , n282109 , n282110 , n282111 , n282112 , n282113 , n282114 , n282115 , 
     n282116 , n282117 , n282118 , n282119 , n282120 , n282121 , n282122 , n282123 , n282124 , n282125 , 
     n282126 , n282127 , n282128 , n282129 , n282130 , n282131 , n282132 , n282133 , n282134 , n282135 , 
     n282136 , n282137 , n282138 , n282139 , n282140 , n282141 , n282142 , n282143 , n282144 , n282145 , 
     n282146 , n282147 , n282148 , n282149 , n282150 , n282151 , n282152 , n282153 , n282154 , n282155 , 
     n282156 , n282157 , n282158 , n282159 , n282160 , n282161 , n282162 , n282163 , n282164 , n282165 , 
     n282166 , n282167 , n282168 , n282169 , n282170 , n282171 , n282172 , n282173 , n282174 , n282175 , 
     n282176 , n282177 , n282178 , n282179 , n282180 , n282181 , n282182 , n282183 , n282184 , n282185 , 
     n282186 , n282187 , n282188 , n282189 , n282190 , n282191 , n282192 , n282193 , n282194 , n282195 , 
     n282196 , n282197 , n282198 , n282199 , n282200 , n282201 , n282202 , n282203 , n282204 , n282205 , 
     n282206 , n282207 , n282208 , n282209 , n282210 , n282211 , n282212 , n282213 , n282214 , n282215 , 
     n282216 , n282217 , n282218 , n282219 , n282220 , n282221 , n282222 , n282223 , n282224 , n282225 , 
     n282226 , n282227 , n282228 , n282229 , n282230 , n282231 , n282232 , n282233 , n282234 , n282235 , 
     n282236 , n282237 , n282238 , n282239 , n282240 , n282241 , n282242 , n282243 , n282244 , n282245 , 
     n282246 , n282247 , n282248 , n282249 , n282250 , n282251 , n282252 , n282253 , n282254 , n282255 , 
     n282256 , n282257 , n282258 , n282259 , n282260 , n282261 , n282262 , n282263 , n282264 , n282265 , 
     n282266 , n282267 , n282268 , n282269 , n282270 , n282271 , n282272 , n282273 , n282274 , n282275 , 
     n282276 , n282277 , n282278 , n282279 , n282280 , n282281 , n282282 , n282283 , n282284 , n282285 , 
     n282286 , n282287 , n282288 , n282289 , n282290 , n282291 , n282292 , n282293 , n282294 , n282295 , 
     n282296 , n282297 , n282298 , n282299 , n282300 , n282301 , n282302 , n282303 , n282304 , n282305 , 
     n282306 , n282307 , n282308 , n282309 , n282310 , n282311 , n282312 , n282313 , n282314 , n282315 , 
     n282316 , n282317 , n282318 , n282319 , n282320 , n282321 , n282322 , n282323 , n282324 , n282325 , 
     n282326 , n282327 , n282328 , n282329 , n282330 , n282331 , n282332 , n282333 , n282334 , n282335 , 
     n282336 , n282337 , n282338 , n282339 , n282340 , n282341 , n282342 , n282343 , n282344 , n282345 , 
     n282346 , n282347 , n282348 , n282349 , n282350 , n282351 , n282352 , n282353 , n282354 , n282355 , 
     n282356 , n282357 , n282358 , n282359 , n282360 , n282361 , n282362 , n282363 , n282364 , n282365 , 
     n282366 , n282367 , n282368 , n282369 , n282370 , n282371 , n282372 , n282373 , n282374 , n282375 , 
     n282376 , n282377 , n282378 , n282379 , n282380 , n282381 , n282382 , n282383 , n282384 , n282385 , 
     n282386 , n282387 , n282388 , n282389 , n282390 , n282391 , n282392 , n282393 , n282394 , n282395 , 
     n282396 , n282397 , n282398 , n282399 , n282400 , n282401 , n282402 , n282403 , n282404 , n282405 , 
     n282406 , n282407 , n282408 , n282409 , n282410 , n282411 , n282412 , n282413 , n282414 , n282415 , 
     n282416 , n282417 , n282418 , n282419 , n282420 , n282421 , n282422 , n282423 , n282424 , n282425 , 
     n282426 , n282427 , n282428 , n282429 , n282430 , n282431 , n282432 , n282433 , n282434 , n282435 , 
     n282436 , n282437 , n282438 , n282439 , n282440 , n282441 , n282442 , n282443 , n282444 , n282445 , 
     n282446 , n282447 , n282448 , n282449 , n282450 , n282451 , n282452 , n282453 , n282454 , n282455 , 
     n282456 , n282457 , n282458 , n282459 , n282460 , n282461 , n282462 , n282463 , n282464 , n282465 , 
     n282466 , n282467 , n282468 , n282469 , n282470 , n282471 , n282472 , n282473 , n282474 , n282475 , 
     n282476 , n282477 , n282478 , n282479 , n282480 , n282481 , n282482 , n282483 , n282484 , n282485 , 
     n282486 , n282487 , n282488 , n282489 , n282490 , n282491 , n282492 , n282493 , n282494 , n282495 , 
     n282496 , n282497 , n282498 , n282499 , n282500 , n282501 , n282502 , n282503 , n282504 , n282505 , 
     n282506 , n282507 , n282508 , n282509 , n282510 , n282511 , n282512 , n282513 , n282514 , n282515 , 
     n282516 , n282517 , n282518 , n282519 , n282520 , n282521 , n282522 , n282523 , n282524 , n282525 , 
     n282526 , n282527 , n282528 , n282529 , n282530 , n282531 , n282532 , n282533 , n282534 , n282535 , 
     n282536 , n282537 , n282538 , n282539 , n282540 , n282541 , n282542 , n282543 , n282544 , n282545 , 
     n282546 , n282547 , n282548 , n282549 , n282550 , n282551 , n282552 , n282553 , n282554 , n282555 , 
     n282556 , n282557 , n282558 , n282559 , n282560 , n282561 , n282562 , n282563 , n282564 , n282565 , 
     n282566 , n282567 , n282568 , n282569 , n282570 , n282571 , n282572 , n282573 , n282574 , n282575 , 
     n282576 , n282577 , n282578 , n282579 , n282580 , n282581 , n282582 , n282583 , n282584 , n282585 , 
     n282586 , n282587 , n282588 , n282589 , n282590 , n282591 , n282592 , n282593 , n282594 , n282595 , 
     n282596 , n282597 , n282598 , n282599 , n282600 , n282601 , n282602 , n282603 , n282604 , n282605 , 
     n282606 , n282607 , n282608 , n282609 , n282610 , n282611 , n282612 , n282613 , n282614 , n282615 , 
     n282616 , n282617 , n282618 , n282619 , n282620 , n282621 , n282622 , n282623 , n282624 , n282625 , 
     n282626 , n282627 , n282628 , n282629 , n282630 , n282631 , n282632 , n282633 , n282634 , n282635 , 
     n282636 , n282637 , n282638 , n282639 , n282640 , n282641 , n282642 , n282643 , n282644 , n282645 , 
     n282646 , n282647 , n282648 , n282649 , n282650 , n282651 , n282652 , n282653 , n282654 , n282655 , 
     n282656 , n282657 , n282658 , n282659 , n282660 , n282661 , n282662 , n282663 , n282664 , n282665 , 
     n282666 , n282667 , n282668 , n282669 , n282670 , n282671 , n282672 , n282673 , n282674 , n282675 , 
     n282676 , n282677 , n282678 , n282679 , n282680 , n282681 , n282682 , n282683 , n282684 , n282685 , 
     n282686 , n282687 , n282688 , n282689 , n282690 , n282691 , n282692 , n282693 , n282694 , n282695 , 
     n282696 , n282697 , n282698 , n282699 , n282700 , n282701 , n282702 , n282703 , n282704 , n282705 , 
     n282706 , n282707 , n282708 , n282709 , n282710 , n282711 , n282712 , n282713 , n282714 , n282715 , 
     n282716 , n282717 , n282718 , n282719 , n282720 , n282721 , n282722 , n282723 , n282724 , n282725 , 
     n282726 , n282727 , n282728 , n282729 , n282730 , n282731 , n282732 , n282733 , n282734 , n282735 , 
     n282736 , n282737 , n282738 , n282739 , n282740 , n282741 , n282742 , n282743 , n282744 , n282745 , 
     n282746 , n282747 , n282748 , n282749 , n282750 , n282751 , n282752 , n282753 , n282754 , n282755 , 
     n282756 , n282757 , n282758 , n282759 , n282760 , n282761 , n282762 , n282763 , n282764 , n282765 , 
     n282766 , n282767 , n282768 , n282769 , n282770 , n282771 , n282772 , n282773 , n282774 , n282775 , 
     n282776 , n282777 , n282778 , n282779 , n282780 , n282781 , n282782 , n282783 , n282784 , n282785 , 
     n282786 , n282787 , n282788 , n282789 , n282790 , n282791 , n282792 , n282793 , n282794 , n282795 , 
     n282796 , n282797 , n282798 , n282799 , n282800 , n282801 , n282802 , n282803 , n282804 , n282805 , 
     n282806 , n282807 , n282808 , n282809 , n282810 , n282811 , n282812 , n282813 , n282814 , n282815 , 
     n282816 , n282817 , n282818 , n282819 , n282820 , n282821 , n282822 , n282823 , n282824 , n282825 , 
     n282826 , n282827 , n282828 , n282829 , n282830 , n282831 , n282832 , n282833 , n282834 , n282835 , 
     n282836 , n282837 , n282838 , n282839 , n282840 , n282841 , n282842 , n282843 , n282844 , n282845 , 
     n282846 , n282847 , n282848 , n282849 , n282850 , n282851 , n282852 , n282853 , n282854 , n282855 , 
     n282856 , n282857 , n282858 , n282859 , n282860 , n282861 , n282862 , n282863 , n282864 , n282865 , 
     n282866 , n282867 , n282868 , n282869 , n282870 , n282871 , n282872 , n282873 , n282874 , n282875 , 
     n282876 , n282877 , n282878 , n282879 , n282880 , n282881 , n282882 , n282883 , n282884 , n282885 , 
     n282886 , n282887 , n282888 , n282889 , n282890 , n282891 , n282892 , n282893 , n282894 , n282895 , 
     n282896 , n282897 , n282898 , n282899 , n282900 , n282901 , n282902 , n282903 , n282904 , n282905 , 
     n282906 , n282907 , n282908 , n282909 , n282910 , n282911 , n282912 , n282913 , n282914 , n282915 , 
     n282916 , n282917 , n282918 , n282919 , n282920 , n282921 , n282922 , n282923 , n282924 , n282925 , 
     n282926 , n282927 , n282928 , n282929 , n282930 , n282931 , n282932 , n282933 , n282934 , n282935 , 
     n282936 , n282937 , n282938 , n282939 , n282940 , n282941 , n282942 , n282943 , n282944 , n282945 , 
     n282946 , n282947 , n282948 , n282949 , n282950 , n282951 , n282952 , n282953 , n282954 , n282955 , 
     n282956 , n282957 , n282958 , n282959 , n282960 , n282961 , n282962 , n282963 , n282964 , n282965 , 
     n282966 , n282967 , n282968 , n282969 , n282970 , n282971 , n282972 , n282973 , n282974 , n282975 , 
     n282976 , n282977 , n282978 , n282979 , n282980 , n282981 , n282982 , n282983 , n282984 , n282985 , 
     n282986 , n282987 , n282988 , n282989 , n282990 , n282991 , n282992 , n282993 , n282994 , n282995 , 
     n282996 , n282997 , n282998 , n282999 , n283000 , n283001 , n283002 , n283003 , n283004 , n283005 , 
     n283006 , n283007 , n283008 , n283009 , n283010 , n283011 , n283012 , n283013 , n283014 , n283015 , 
     n283016 , n283017 , n283018 , n283019 , n283020 , n283021 , n283022 , n283023 , n283024 , n283025 , 
     n283026 , n283027 , n283028 , n283029 , n283030 , n283031 , n283032 , n283033 , n283034 , n283035 , 
     n283036 , n283037 , n283038 , n283039 , n283040 , n283041 , n283042 , n283043 , n283044 , n283045 , 
     n283046 , n283047 , n283048 , n283049 , n283050 , n283051 , n283052 , n283053 , n283054 , n283055 , 
     n283056 , n283057 , n283058 , n283059 , n283060 , n283061 , n283062 , n283063 , n283064 , n283065 , 
     n283066 , n283067 , n283068 , n283069 , n283070 , n283071 , n283072 , n283073 , n283074 , n283075 , 
     n283076 , n283077 , n283078 , n283079 , n283080 , n283081 , n283082 , n283083 , n283084 , n283085 , 
     n283086 , n283087 , n283088 , n283089 , n283090 , n283091 , n283092 , n283093 , n283094 , n283095 , 
     n283096 , n283097 , n283098 , n283099 , n283100 , n283101 , n283102 , n283103 , n283104 , n283105 , 
     n283106 , n283107 , n283108 , n283109 , n283110 , n283111 , n283112 , n283113 , n283114 , n283115 , 
     n283116 , n283117 , n283118 , n283119 , n283120 , n283121 , n283122 , n283123 , n283124 , n283125 , 
     n283126 , n283127 , n283128 , n283129 , n283130 , n283131 , n283132 , n283133 , n283134 , n283135 , 
     n283136 , n283137 , n283138 , n283139 , n283140 , n283141 , n283142 , n283143 , n283144 , n283145 , 
     n283146 , n283147 , n283148 , n283149 , n283150 , n283151 , n283152 , n283153 , n283154 , n283155 , 
     n283156 , n283157 , n283158 , n283159 , n283160 , n283161 , n283162 , n283163 , n283164 , n283165 , 
     n283166 , n283167 , n283168 , n283169 , n283170 , n283171 , n283172 , n283173 , n283174 , n283175 , 
     n283176 , n283177 , n283178 , n283179 , n283180 , n283181 , n283182 , n283183 , n283184 , n283185 , 
     n283186 , n283187 , n283188 , n283189 , n283190 , n283191 , n283192 , n283193 , n283194 , n283195 , 
     n283196 , n283197 , n283198 , n283199 , n283200 , n283201 , n283202 , n283203 , n283204 , n283205 , 
     n283206 , n283207 , n283208 , n283209 , n283210 , n283211 , n283212 , n283213 , n283214 , n283215 , 
     n283216 , n283217 , n283218 , n283219 , n283220 , n283221 , n283222 , n283223 , n283224 , n283225 , 
     n283226 , n283227 , n283228 , n283229 , n283230 , n283231 , n283232 , n283233 , n283234 , n283235 , 
     n283236 , n283237 , n283238 , n283239 , n283240 , n283241 , n283242 , n283243 , n283244 , n283245 , 
     n283246 , n283247 , n283248 , n283249 , n283250 , n283251 , n283252 , n283253 , n283254 , n283255 , 
     n283256 , n283257 , n283258 , n283259 , n283260 , n283261 , n283262 , n283263 , n283264 , n283265 , 
     n283266 , n283267 , n283268 , n283269 , n283270 , n283271 , n283272 , n283273 , n283274 , n283275 , 
     n283276 , n283277 , n283278 , n283279 , n283280 , n283281 , n283282 , n283283 , n283284 , n283285 , 
     n283286 , n283287 , n283288 , n283289 , n283290 , n283291 , n283292 , n283293 , n283294 , n283295 , 
     n283296 , n283297 , n283298 , n283299 , n283300 , n283301 , n283302 , n283303 , n283304 , n283305 , 
     n283306 , n283307 , n283308 , n283309 , n283310 , n283311 , n283312 , n283313 , n283314 , n283315 , 
     n283316 , n283317 , n283318 , n283319 , n283320 , n283321 , n283322 , n283323 , n283324 , n283325 , 
     n283326 , n283327 , n283328 , n283329 , n283330 , n283331 , n283332 , n283333 , n283334 , n283335 , 
     n283336 , n283337 , n283338 , n283339 , n283340 , n283341 , n283342 , n283343 , n283344 , n283345 , 
     n283346 , n283347 , n283348 , n283349 , n283350 , n283351 , n283352 , n283353 , n283354 , n283355 , 
     n283356 , n283357 , n283358 , n283359 , n283360 , n283361 , n283362 , n283363 , n283364 , n283365 , 
     n283366 , n283367 , n283368 , n283369 , n283370 , n283371 , n283372 , n283373 , n283374 , n283375 , 
     n283376 , n283377 , n283378 , n283379 , n283380 , n283381 , n283382 , n283383 , n283384 , n283385 , 
     n283386 , n283387 , n283388 , n283389 , n283390 , n283391 , n283392 , n283393 , n283394 , n283395 , 
     n283396 , n283397 , n283398 , n283399 , n283400 , n283401 , n283402 , n283403 , n283404 , n283405 , 
     n283406 , n283407 , n283408 , n283409 , n283410 , n283411 , n283412 , n283413 , n283414 , n283415 , 
     n283416 , n283417 , n283418 , n283419 , n283420 , n283421 , n283422 , n283423 , n283424 , n283425 , 
     n283426 , n283427 , n283428 , n283429 , n283430 , n283431 , n283432 , n283433 , n283434 , n283435 , 
     n283436 , n283437 , n283438 , n283439 , n283440 , n283441 , n283442 , n283443 , n283444 , n283445 , 
     n283446 , n283447 , n283448 , n283449 , n283450 , n283451 , n283452 , n283453 , n283454 , n283455 , 
     n283456 , n283457 , n283458 , n283459 , n283460 , n283461 , n283462 , n283463 , n283464 , n283465 , 
     n283466 , n283467 , n283468 , n283469 , n283470 , n283471 , n283472 , n283473 , n283474 , n283475 , 
     n283476 , n283477 , n283478 , n283479 , n283480 , n283481 , n283482 , n283483 , n283484 , n283485 , 
     n283486 , n283487 , n283488 , n283489 , n283490 , n283491 , n283492 , n283493 , n283494 , n283495 , 
     n283496 , n283497 , n283498 , n283499 , n283500 , n283501 , n283502 , n283503 , n283504 , n283505 , 
     n283506 , n283507 , n283508 , n283509 , n283510 , n283511 , n283512 , n283513 , n283514 , n283515 , 
     n283516 , n283517 , n283518 , n283519 , n283520 , n283521 , n283522 , n283523 , n283524 , n283525 , 
     n283526 , n283527 , n283528 , n283529 , n283530 , n283531 , n283532 , n283533 , n283534 , n283535 , 
     n283536 , n283537 , n283538 , n283539 , n283540 , n283541 , n283542 , n283543 , n283544 , n283545 , 
     n283546 , n283547 , n283548 , n283549 , n283550 , n283551 , n283552 , n283553 , n283554 , n283555 , 
     n283556 , n283557 , n283558 , n283559 , n283560 , n283561 , n283562 , n283563 , n283564 , n283565 , 
     n283566 , n283567 , n283568 , n283569 , n283570 , n283571 , n283572 , n283573 , n283574 , n283575 , 
     n283576 , n283577 , n283578 , n283579 , n283580 , n283581 , n283582 , n283583 , n283584 , n283585 , 
     n283586 , n283587 , n283588 , n283589 , n283590 , n283591 , n283592 , n283593 , n283594 , n283595 , 
     n283596 , n283597 , n283598 , n283599 , n283600 , n283601 , n283602 , n283603 , n283604 , n283605 , 
     n283606 , n283607 , n283608 , n283609 , n283610 , n283611 , n283612 , n283613 , n283614 , n283615 , 
     n283616 , n283617 , n283618 , n283619 , n283620 , n283621 , n283622 , n283623 , n283624 , n283625 , 
     n283626 , n283627 , n283628 , n283629 , n283630 , n283631 , n283632 , n283633 , n283634 , n283635 , 
     n283636 , n283637 , n283638 , n283639 , n283640 , n283641 , n283642 , n283643 , n283644 , n283645 , 
     n283646 , n283647 , n283648 , n283649 , n283650 , n283651 , n283652 , n283653 , n283654 , n283655 , 
     n283656 , n283657 , n283658 , n283659 , n283660 , n283661 , n283662 , n283663 , n283664 , n283665 , 
     n283666 , n283667 , n283668 , n283669 , n283670 , n283671 , n283672 , n283673 , n283674 , n283675 , 
     n283676 , n283677 , n283678 , n283679 , n283680 , n283681 , n283682 , n283683 , n283684 , n283685 , 
     n283686 , n283687 , n283688 , n283689 , n283690 , n283691 , n283692 , n283693 , n283694 , n283695 , 
     n283696 , n283697 , n283698 , n283699 , n283700 , n283701 , n283702 , n283703 , n283704 , n283705 , 
     n283706 , n283707 , n283708 , n283709 , n283710 , n283711 , n283712 , n283713 , n283714 , n283715 , 
     n283716 , n283717 , n283718 , n283719 , n283720 , n283721 , n283722 , n283723 , n283724 , n283725 , 
     n283726 , n283727 , n283728 , n283729 , n283730 , n283731 , n283732 , n283733 , n283734 , n283735 , 
     n283736 , n283737 , n283738 , n283739 , n283740 , n283741 , n283742 , n283743 , n283744 , n283745 , 
     n283746 , n283747 , n283748 , n283749 , n283750 , n283751 , n283752 , n283753 , n283754 , n283755 , 
     n283756 , n283757 , n283758 , n283759 , n283760 , n283761 , n283762 , n283763 , n283764 , n283765 , 
     n283766 , n283767 , n283768 , n283769 , n283770 , n283771 , n283772 , n283773 , n283774 , n283775 , 
     n283776 , n283777 , n283778 , n283779 , n283780 , n283781 , n283782 , n283783 , n283784 , n283785 , 
     n283786 , n283787 , n283788 , n283789 , n283790 , n283791 , n283792 , n283793 , n283794 , n283795 , 
     n283796 , n283797 , n283798 , n283799 , n283800 , n283801 , n283802 , n283803 , n283804 , n283805 , 
     n283806 , n283807 , n283808 , n283809 , n283810 , n283811 , n283812 , n283813 , n283814 , n283815 , 
     n283816 , n283817 , n283818 , n283819 , n283820 , n283821 , n283822 , n283823 , n283824 , n283825 , 
     n283826 , n283827 , n283828 , n283829 , n283830 , n283831 , n283832 , n283833 , n283834 , n283835 , 
     n283836 , n283837 , n283838 , n283839 , n283840 , n283841 , n283842 , n283843 , n283844 , n283845 , 
     n283846 , n283847 , n283848 , n283849 , n283850 , n283851 , n283852 , n283853 , n283854 , n283855 , 
     n283856 , n283857 , n283858 , n283859 , n283860 , n283861 , n283862 , n283863 , n283864 , n283865 , 
     n283866 , n283867 , n283868 , n283869 , n283870 , n283871 , n283872 , n283873 , n283874 , n283875 , 
     n283876 , n283877 , n283878 , n283879 , n283880 , n283881 , n283882 , n283883 , n283884 , n283885 , 
     n283886 , n283887 , n283888 , n283889 , n283890 , n283891 , n283892 , n283893 , n283894 , n283895 , 
     n283896 , n283897 , n283898 , n283899 , n283900 , n283901 , n283902 , n283903 , n283904 , n283905 , 
     n283906 , n283907 , n283908 , n283909 , n283910 , n283911 , n283912 , n283913 , n283914 , n283915 , 
     n283916 , n283917 , n283918 , n283919 , n283920 , n283921 , n283922 , n283923 , n283924 , n283925 , 
     n283926 , n283927 , n283928 , n283929 , n283930 , n283931 , n283932 , n283933 , n283934 , n283935 , 
     n283936 , n283937 , n283938 , n283939 , n283940 , n283941 , n283942 , n283943 , n283944 , n283945 , 
     n283946 , n283947 , n283948 , n283949 , n283950 , n283951 , n283952 , n283953 , n283954 , n283955 , 
     n283956 , n283957 , n283958 , n283959 , n283960 , n283961 , n283962 , n283963 , n283964 , n283965 , 
     n283966 , n283967 , n283968 , n283969 , n283970 , n283971 , n283972 , n283973 , n283974 , n283975 , 
     n283976 , n283977 , n283978 , n283979 , n283980 , n283981 , n283982 , n283983 , n283984 , n283985 , 
     n283986 , n283987 , n283988 , n283989 , n283990 , n283991 , n283992 , n283993 , n283994 , n283995 , 
     n283996 , n283997 , n283998 , n283999 , n284000 , n284001 , n284002 , n284003 , n284004 , n284005 , 
     n284006 , n284007 , n284008 , n284009 , n284010 , n284011 , n284012 , n284013 , n284014 , n284015 , 
     n284016 , n284017 , n284018 , n284019 , n284020 , n284021 , n284022 , n284023 , n284024 , n284025 , 
     n284026 , n284027 , n284028 , n284029 , n284030 , n284031 , n284032 , n284033 , n284034 , n284035 , 
     n284036 , n284037 , n284038 , n284039 , n284040 , n284041 , n284042 , n284043 , n284044 , n284045 , 
     n284046 , n284047 , n284048 , n284049 , n284050 , n284051 , n284052 , n284053 , n284054 , n284055 , 
     n284056 , n284057 , n284058 , n284059 , n284060 , n284061 , n284062 , n284063 , n284064 , n284065 , 
     n284066 , n284067 , n284068 , n284069 , n284070 , n284071 , n284072 , n284073 , n284074 , n284075 , 
     n284076 , n284077 , n284078 , n284079 , n284080 , n284081 , n284082 , n284083 , n284084 , n284085 , 
     n284086 , n284087 , n284088 , n284089 , n284090 , n284091 , n284092 , n284093 , n284094 , n284095 , 
     n284096 , n284097 , n284098 , n284099 , n284100 , n284101 , n284102 , n284103 , n284104 , n284105 , 
     n284106 , n284107 , n284108 , n284109 , n284110 , n284111 , n284112 , n284113 , n284114 , n284115 , 
     n284116 , n284117 , n284118 , n284119 , n284120 , n284121 , n284122 , n284123 , n284124 , n284125 , 
     n284126 , n284127 , n284128 , n284129 , n284130 , n284131 , n284132 , n284133 , n284134 , n284135 , 
     n284136 , n284137 , n284138 , n284139 , n284140 , n284141 , n284142 , n284143 , n284144 , n284145 , 
     n284146 , n284147 , n284148 , n284149 , n284150 , n284151 , n284152 , n284153 , n284154 , n284155 , 
     n284156 , n284157 , n284158 , n284159 , n284160 , n284161 , n284162 , n284163 , n284164 , n284165 , 
     n284166 , n284167 , n284168 , n284169 , n284170 , n284171 , n284172 , n284173 , n284174 , n284175 , 
     n284176 , n284177 , n284178 , n284179 , n284180 , n284181 , n284182 , n284183 , n284184 , n284185 , 
     n284186 , n284187 , n284188 , n284189 , n284190 , n284191 , n284192 , n284193 , n284194 , n284195 , 
     n284196 , n284197 , n284198 , n284199 , n284200 , n284201 , n284202 , n284203 , n284204 , n284205 , 
     n284206 , n284207 , n284208 , n284209 , n284210 , n284211 , n284212 , n284213 , n284214 , n284215 , 
     n284216 , n284217 , n284218 , n284219 , n284220 , n284221 , n284222 , n284223 , n284224 , n284225 , 
     n284226 , n284227 , n284228 , n284229 , n284230 , n284231 , n284232 , n284233 , n284234 , n284235 , 
     n284236 , n284237 , n284238 , n284239 , n284240 , n284241 , n284242 , n284243 , n284244 , n284245 , 
     n284246 , n284247 , n284248 , n284249 , n284250 , n284251 , n284252 , n284253 , n284254 , n284255 , 
     n284256 , n284257 , n284258 , n284259 , n284260 , n284261 , n284262 , n284263 , n284264 , n284265 , 
     n284266 , n284267 , n284268 , n284269 , n284270 , n284271 , n284272 , n284273 , n284274 , n284275 , 
     n284276 , n284277 , n284278 , n284279 , n284280 , n284281 , n284282 , n284283 , n284284 , n284285 , 
     n284286 , n284287 , n284288 , n284289 , n284290 , n284291 , n284292 , n284293 , n284294 , n284295 , 
     n284296 , n284297 , n284298 , n284299 , n284300 , n284301 , n284302 , n284303 , n284304 , n284305 , 
     n284306 , n284307 , n284308 , n284309 , n284310 , n284311 , n284312 , n284313 , n284314 , n284315 , 
     n284316 , n284317 , n284318 , n284319 , n284320 , n284321 , n284322 , n284323 , n284324 , n284325 , 
     n284326 , n284327 , n284328 , n284329 , n284330 , n284331 , n284332 , n284333 , n284334 , n284335 , 
     n284336 , n284337 , n284338 , n284339 , n284340 , n284341 , n284342 , n284343 , n284344 , n284345 , 
     n284346 , n284347 , n284348 , n284349 , n284350 , n284351 , n284352 , n284353 , n284354 , n284355 , 
     n284356 , n284357 , n284358 , n284359 , n284360 , n284361 , n284362 , n284363 , n284364 , n284365 , 
     n284366 , n284367 , n284368 , n284369 , n284370 , n284371 , n284372 , n284373 , n284374 , n284375 , 
     n284376 , n284377 , n284378 , n284379 , n284380 , n284381 , n284382 , n284383 , n284384 , n284385 , 
     n284386 , n284387 , n284388 , n284389 , n284390 , n284391 , n284392 , n284393 , n284394 , n284395 , 
     n284396 , n284397 , n284398 , n284399 , n284400 , n284401 , n284402 , n284403 , n284404 , n284405 , 
     n284406 , n284407 , n284408 , n284409 , n284410 , n284411 , n284412 , n284413 , n284414 , n284415 , 
     n284416 , n284417 , n284418 , n284419 , n284420 , n284421 , n284422 , n284423 , n284424 , n284425 , 
     n284426 , n284427 , n284428 , n284429 , n284430 , n284431 , n284432 , n284433 , n284434 , n284435 , 
     n284436 , n284437 , n284438 , n284439 , n284440 , n284441 , n284442 , n284443 , n284444 , n284445 , 
     n284446 , n284447 , n284448 , n284449 , n284450 , n284451 , n284452 , n284453 , n284454 , n284455 , 
     n284456 , n284457 , n284458 , n284459 , n284460 , n284461 , n284462 , n284463 , n284464 , n284465 , 
     n284466 , n284467 , n284468 , n284469 , n284470 , n284471 , n284472 , n284473 , n284474 , n284475 , 
     n284476 , n284477 , n284478 , n284479 , n284480 , n284481 , n284482 , n284483 , n284484 , n284485 , 
     n284486 , n284487 , n284488 , n284489 , n284490 , n284491 , n284492 , n284493 , n284494 , n284495 , 
     n284496 , n284497 , n284498 , n284499 , n284500 , n284501 , n284502 , n284503 , n284504 , n284505 , 
     n284506 , n284507 , n284508 , n284509 , n284510 , n284511 , n284512 , n284513 , n284514 , n284515 , 
     n284516 , n284517 , n284518 , n284519 , n284520 , n284521 , n284522 , n284523 , n284524 , n284525 , 
     n284526 , n284527 , n284528 , n284529 , n284530 , n284531 , n284532 , n284533 , n284534 , n284535 , 
     n284536 , n284537 , n284538 , n284539 , n284540 , n284541 , n284542 , n284543 , n284544 , n284545 , 
     n284546 , n284547 , n284548 , n284549 , n284550 , n284551 , n284552 , n284553 , n284554 , n284555 , 
     n284556 , n284557 , n284558 , n284559 , n284560 , n284561 , n284562 , n284563 , n284564 , n284565 , 
     n284566 , n284567 , n284568 , n284569 , n284570 , n284571 , n284572 , n284573 , n284574 , n284575 , 
     n284576 , n284577 , n284578 , n284579 , n284580 , n284581 , n284582 , n284583 , n284584 , n284585 , 
     n284586 , n284587 , n284588 , n284589 , n284590 , n284591 , n284592 , n284593 , n284594 , n284595 , 
     n284596 , n284597 , n284598 , n284599 , n284600 , n284601 , n284602 , n284603 , n284604 , n284605 , 
     n284606 , n284607 , n284608 , n284609 , n284610 , n284611 , n284612 , n284613 , n284614 , n284615 , 
     n284616 , n284617 , n284618 , n284619 , n284620 , n284621 , n284622 , n284623 , n284624 , n284625 , 
     n284626 , n284627 , n284628 , n284629 , n284630 , n284631 , n284632 , n284633 , n284634 , n284635 , 
     n284636 , n284637 , n284638 , n284639 , n284640 , n284641 , n284642 , n284643 , n284644 , n284645 , 
     n284646 , n284647 , n284648 , n284649 , n284650 , n284651 , n284652 , n284653 , n284654 , n284655 , 
     n284656 , n284657 , n284658 , n284659 , n284660 , n284661 , n284662 , n284663 , n284664 , n284665 , 
     n284666 , n284667 , n284668 , n284669 , n284670 , n284671 , n284672 , n284673 , n284674 , n284675 , 
     n284676 , n284677 , n284678 , n284679 , n284680 , n284681 , n284682 , n284683 , n284684 , n284685 , 
     n284686 , n284687 , n284688 , n284689 , n284690 , n284691 , n284692 , n284693 , n284694 , n284695 , 
     n284696 , n284697 , n284698 , n284699 , n284700 , n284701 , n284702 , n284703 , n284704 , n284705 , 
     n284706 , n284707 , n284708 , n284709 , n284710 , n284711 , n284712 , n284713 , n284714 , n284715 , 
     n284716 , n284717 , n284718 , n284719 , n284720 , n284721 , n284722 , n284723 , n284724 , n284725 , 
     n284726 , n284727 , n284728 , n284729 , n284730 , n284731 , n284732 , n284733 , n284734 , n284735 , 
     n284736 , n284737 , n284738 , n284739 , n284740 , n284741 , n284742 , n284743 , n284744 , n284745 , 
     n284746 , n284747 , n284748 , n284749 , n284750 , n284751 , n284752 , n284753 , n284754 , n284755 , 
     n284756 , n284757 , n284758 , n284759 , n284760 , n284761 , n284762 , n284763 , n284764 , n284765 , 
     n284766 , n284767 , n284768 , n284769 , n284770 , n284771 , n284772 , n284773 , n284774 , n284775 , 
     n284776 , n284777 , n284778 , n284779 , n284780 , n284781 , n284782 , n284783 , n284784 , n284785 , 
     n284786 , n284787 , n284788 , n284789 , n284790 , n284791 , n284792 , n284793 , n284794 , n284795 , 
     n284796 , n284797 , n284798 , n284799 , n284800 , n284801 , n284802 , n284803 , n284804 , n284805 , 
     n284806 , n284807 , n284808 , n284809 , n284810 , n284811 , n284812 , n284813 , n284814 , n284815 , 
     n284816 , n284817 , n284818 , n284819 , n284820 , n284821 , n284822 , n284823 , n284824 , n284825 , 
     n284826 , n284827 , n284828 , n284829 , n284830 , n284831 , n284832 , n284833 , n284834 , n284835 , 
     n284836 , n284837 , n284838 , n284839 , n284840 , n284841 , n284842 , n284843 , n284844 , n284845 , 
     n284846 , n284847 , n284848 , n284849 , n284850 , n284851 , n284852 , n284853 , n284854 , n284855 , 
     n284856 , n284857 , n284858 , n284859 , n284860 , n284861 , n284862 , n284863 , n284864 , n284865 , 
     n284866 , n284867 , n284868 , n284869 , n284870 , n284871 , n284872 , n284873 , n284874 , n284875 , 
     n284876 , n284877 , n284878 , n284879 , n284880 , n284881 , n284882 , n284883 , n284884 , n284885 , 
     n284886 , n284887 , n284888 , n284889 , n284890 , n284891 , n284892 , n284893 , n284894 , n284895 , 
     n284896 , n284897 , n284898 , n284899 , n284900 , n284901 , n284902 , n284903 , n284904 , n284905 , 
     n284906 , n284907 , n284908 , n284909 , n284910 , n284911 , n284912 , n284913 , n284914 , n284915 , 
     n284916 , n284917 , n284918 , n284919 , n284920 , n284921 , n284922 , n284923 , n284924 , n284925 , 
     n284926 , n284927 , n284928 , n284929 , n284930 , n284931 , n284932 , n284933 , n284934 , n284935 , 
     n284936 , n284937 , n284938 , n284939 , n284940 , n284941 , n284942 , n284943 , n284944 , n284945 , 
     n284946 , n284947 , n284948 , n284949 , n284950 , n284951 , n284952 , n284953 , n284954 , n284955 , 
     n284956 , n284957 , n284958 , n284959 , n284960 , n284961 , n284962 , n284963 , n284964 , n284965 , 
     n284966 , n284967 , n284968 , n284969 , n284970 , n284971 , n284972 , n284973 , n284974 , n284975 , 
     n284976 , n284977 , n284978 , n284979 , n284980 , n284981 , n284982 , n284983 , n284984 , n284985 , 
     n284986 , n284987 , n284988 , n284989 , n284990 , n284991 , n284992 , n284993 , n284994 , n284995 , 
     n284996 , n284997 , n284998 , n284999 , n285000 , n285001 , n285002 , n285003 , n285004 , n285005 , 
     n285006 , n285007 , n285008 , n285009 , n285010 , n285011 , n285012 , n285013 , n285014 , n285015 , 
     n285016 , n285017 , n285018 , n285019 , n285020 , n285021 , n285022 , n285023 , n285024 , n285025 , 
     n285026 , n285027 , n285028 , n285029 , n285030 , n285031 , n285032 , n285033 , n285034 , n285035 , 
     n285036 , n285037 , n285038 , n285039 , n285040 , n285041 , n285042 , n285043 , n285044 , n285045 , 
     n285046 , n285047 , n285048 , n285049 , n285050 , n285051 , n285052 , n285053 , n285054 , n285055 , 
     n285056 , n285057 , n285058 , n285059 , n285060 , n285061 , n285062 , n285063 , n285064 , n285065 , 
     n285066 , n285067 , n285068 , n285069 , n285070 , n285071 , n285072 , n285073 , n285074 , n285075 , 
     n285076 , n285077 , n285078 , n285079 , n285080 , n285081 , n285082 , n285083 , n285084 , n285085 , 
     n285086 , n285087 , n285088 , n285089 , n285090 , n285091 , n285092 , n285093 , n285094 , n285095 , 
     n285096 , n285097 , n285098 , n285099 , n285100 , n285101 , n285102 , n285103 , n285104 , n285105 , 
     n285106 , n285107 , n285108 , n285109 , n285110 , n285111 , n285112 , n285113 , n285114 , n285115 , 
     n285116 , n285117 , n285118 , n285119 , n285120 , n285121 , n285122 , n285123 , n285124 , n285125 , 
     n285126 , n285127 , n285128 , n285129 , n285130 , n285131 , n285132 , n285133 , n285134 , n285135 , 
     n285136 , n285137 , n285138 , n285139 , n285140 , n285141 , n285142 , n285143 , n285144 , n285145 , 
     n285146 , n285147 , n285148 , n285149 , n285150 , n285151 , n285152 , n285153 , n285154 , n285155 , 
     n285156 , n285157 , n285158 , n285159 , n285160 , n285161 , n285162 , n285163 , n285164 , n285165 , 
     n285166 , n285167 , n285168 , n285169 , n285170 , n285171 , n285172 , n285173 , n285174 , n285175 , 
     n285176 , n285177 , n285178 , n285179 , n285180 , n285181 , n285182 , n285183 , n285184 , n285185 , 
     n285186 , n285187 , n285188 , n285189 , n285190 , n285191 , n285192 , n285193 , n285194 , n285195 , 
     n285196 , n285197 , n285198 , n285199 , n285200 , n285201 , n285202 , n285203 , n285204 , n285205 , 
     n285206 , n285207 , n285208 , n285209 , n285210 , n285211 , n285212 , n285213 , n285214 , n285215 , 
     n285216 , n285217 , n285218 , n285219 , n285220 , n285221 , n285222 , n285223 , n285224 , n285225 , 
     n285226 , n285227 , n285228 , n285229 , n285230 , n285231 , n285232 , n285233 , n285234 , n285235 , 
     n285236 , n285237 , n285238 , n285239 , n285240 , n285241 , n285242 , n285243 , n285244 , n285245 , 
     n285246 , n285247 , n285248 , n285249 , n285250 , n285251 , n285252 , n285253 , n285254 , n285255 , 
     n285256 , n285257 , n285258 , n285259 , n285260 , n285261 , n285262 , n285263 , n285264 , n285265 , 
     n285266 , n285267 , n285268 , n285269 , n285270 , n285271 , n285272 , n285273 , n285274 , n285275 , 
     n285276 , n285277 , n285278 , n285279 , n285280 , n285281 , n285282 , n285283 , n285284 , n285285 , 
     n285286 , n285287 , n285288 , n285289 , n285290 , n285291 , n285292 , n285293 , n285294 , n285295 , 
     n285296 , n285297 , n285298 , n285299 , n285300 , n285301 , n285302 , n285303 , n285304 , n285305 , 
     n285306 , n285307 , n285308 , n285309 , n285310 , n285311 , n285312 , n285313 , n285314 , n285315 , 
     n285316 , n285317 , n285318 , n285319 , n285320 , n285321 , n285322 , n285323 , n285324 , n285325 , 
     n285326 , n285327 , n285328 , n285329 , n285330 , n285331 , n285332 , n285333 , n285334 , n285335 , 
     n285336 , n285337 , n285338 , n285339 , n285340 , n285341 , n285342 , n285343 , n285344 , n285345 , 
     n285346 , n285347 , n285348 , n285349 , n285350 , n285351 , n285352 , n285353 , n285354 , n285355 , 
     n285356 , n285357 , n285358 , n285359 , n285360 , n285361 , n285362 , n285363 , n285364 , n285365 , 
     n285366 , n285367 , n285368 , n285369 , n285370 , n285371 , n285372 , n285373 , n285374 , n285375 , 
     n285376 , n285377 , n285378 , n285379 , n285380 , n285381 , n285382 , n285383 , n285384 , n285385 , 
     n285386 , n285387 , n285388 , n285389 , n285390 , n285391 , n285392 , n285393 , n285394 , n285395 , 
     n285396 , n285397 , n285398 , n285399 , n285400 , n285401 , n285402 , n285403 , n285404 , n285405 , 
     n285406 , n285407 , n285408 , n285409 , n285410 , n285411 , n285412 , n285413 , n285414 , n285415 , 
     n285416 , n285417 , n285418 , n285419 , n285420 , n285421 , n285422 , n285423 , n285424 , n285425 , 
     n285426 , n285427 , n285428 , n285429 , n285430 , n285431 , n285432 , n285433 , n285434 , n285435 , 
     n285436 , n285437 , n285438 , n285439 , n285440 , n285441 , n285442 , n285443 , n285444 , n285445 , 
     n285446 , n285447 , n285448 , n285449 , n285450 , n285451 , n285452 , n285453 , n285454 , n285455 , 
     n285456 , n285457 , n285458 , n285459 , n285460 , n285461 , n285462 , n285463 , n285464 , n285465 , 
     n285466 , n285467 , n285468 , n285469 , n285470 , n285471 , n285472 , n285473 , n285474 , n285475 , 
     n285476 , n285477 , n285478 , n285479 , n285480 , n285481 , n285482 , n285483 , n285484 , n285485 , 
     n285486 , n285487 , n285488 , n285489 , n285490 , n285491 , n285492 , n285493 , n285494 , n285495 , 
     n285496 , n285497 , n285498 , n285499 , n285500 , n285501 , n285502 , n285503 , n285504 , n285505 , 
     n285506 , n285507 , n285508 , n285509 , n285510 , n285511 , n285512 , n285513 , n285514 , n285515 , 
     n285516 , n285517 , n285518 , n285519 , n285520 , n285521 , n285522 , n285523 , n285524 , n285525 , 
     n285526 , n285527 , n285528 , n285529 , n285530 , n285531 , n285532 , n285533 , n285534 , n285535 , 
     n285536 , n285537 , n285538 , n285539 , n285540 , n285541 , n285542 , n285543 , n285544 , n285545 , 
     n285546 , n285547 , n285548 , n285549 , n285550 , n285551 , n285552 , n285553 , n285554 , n285555 , 
     n285556 , n285557 , n285558 , n285559 , n285560 , n285561 , n285562 , n285563 , n285564 , n285565 , 
     n285566 , n285567 , n285568 , n285569 , n285570 , n285571 , n285572 , n285573 , n285574 , n285575 , 
     n285576 , n285577 , n285578 , n285579 , n285580 , n285581 , n285582 , n285583 , n285584 , n285585 , 
     n285586 , n285587 , n285588 , n285589 , n285590 , n285591 , n285592 , n285593 , n285594 , n285595 , 
     n285596 , n285597 , n285598 , n285599 , n285600 , n285601 , n285602 , n285603 , n285604 , n285605 , 
     n285606 , n285607 , n285608 , n285609 , n285610 , n285611 , n285612 , n285613 , n285614 , n285615 , 
     n285616 , n285617 , n285618 , n285619 , n285620 , n285621 , n285622 , n285623 , n285624 , n285625 , 
     n285626 , n285627 , n285628 , n285629 , n285630 , n285631 , n285632 , n285633 , n285634 , n285635 , 
     n285636 , n285637 , n285638 , n285639 , n285640 , n285641 , n285642 , n285643 , n285644 , n285645 , 
     n285646 , n285647 , n285648 , n285649 , n285650 , n285651 , n285652 , n285653 , n285654 , n285655 , 
     n285656 , n285657 , n285658 , n285659 , n285660 , n285661 , n285662 , n285663 , n285664 , n285665 , 
     n285666 , n285667 , n285668 , n285669 , n285670 , n285671 , n285672 , n285673 , n285674 , n285675 , 
     n285676 , n285677 , n285678 , n285679 , n285680 , n285681 , n285682 , n285683 , n285684 , n285685 , 
     n285686 , n285687 , n285688 , n285689 , n285690 , n285691 , n285692 , n285693 , n285694 , n285695 , 
     n285696 , n285697 , n285698 , n285699 , n285700 , n285701 , n285702 , n285703 , n285704 , n285705 , 
     n285706 , n285707 , n285708 , n285709 , n285710 , n285711 , n285712 , n285713 , n285714 , n285715 , 
     n285716 , n285717 , n285718 , n285719 , n285720 , n285721 , n285722 , n285723 , n285724 , n285725 , 
     n285726 , n285727 , n285728 , n285729 , n285730 , n285731 , n285732 , n285733 , n285734 , n285735 , 
     n285736 , n285737 , n285738 , n285739 , n285740 , n285741 , n285742 , n285743 , n285744 , n285745 , 
     n285746 , n285747 , n285748 , n285749 , n285750 , n285751 , n285752 , n285753 , n285754 , n285755 , 
     n285756 , n285757 , n285758 , n285759 , n285760 , n285761 , n285762 , n285763 , n285764 , n285765 , 
     n285766 , n285767 , n285768 , n285769 , n285770 , n285771 , n285772 , n285773 , n285774 , n285775 , 
     n285776 , n285777 , n285778 , n285779 , n285780 , n285781 , n285782 , n285783 , n285784 , n285785 , 
     n285786 , n285787 , n285788 , n285789 , n285790 , n285791 , n285792 , n285793 , n285794 , n285795 , 
     n285796 , n285797 , n285798 , n285799 , n285800 , n285801 , n285802 , n285803 , n285804 , n285805 , 
     n285806 , n285807 , n285808 , n285809 , n285810 , n285811 , n285812 , n285813 , n285814 , n285815 , 
     n285816 , n285817 , n285818 , n285819 , n285820 , n285821 , n285822 , n285823 , n285824 , n285825 , 
     n285826 , n285827 , n285828 , n285829 , n285830 , n285831 , n285832 , n285833 , n285834 , n285835 , 
     n285836 , n285837 , n285838 , n285839 , n285840 , n285841 , n285842 , n285843 , n285844 , n285845 , 
     n285846 , n285847 , n285848 , n285849 , n285850 , n285851 , n285852 , n285853 , n285854 , n285855 , 
     n285856 , n285857 , n285858 , n285859 , n285860 , n285861 , n285862 , n285863 , n285864 , n285865 , 
     n285866 , n285867 , n285868 , n285869 , n285870 , n285871 , n285872 , n285873 , n285874 , n285875 , 
     n285876 , n285877 , n285878 , n285879 , n285880 , n285881 , n285882 , n285883 , n285884 , n285885 , 
     n285886 , n285887 , n285888 , n285889 , n285890 , n285891 , n285892 , n285893 , n285894 , n285895 , 
     n285896 , n285897 , n285898 , n285899 , n285900 , n285901 , n285902 , n285903 , n285904 , n285905 , 
     n285906 , n285907 , n285908 , n285909 , n285910 , n285911 , n285912 , n285913 , n285914 , n285915 , 
     n285916 , n285917 , n285918 , n285919 , n285920 , n285921 , n285922 , n285923 , n285924 , n285925 , 
     n285926 , n285927 , n285928 , n285929 , n285930 , n285931 , n285932 , n285933 , n285934 , n285935 , 
     n285936 , n285937 , n285938 , n285939 , n285940 , n285941 , n285942 , n285943 , n285944 , n285945 , 
     n285946 , n285947 , n285948 , n285949 , n285950 , n285951 , n285952 , n285953 , n285954 , n285955 , 
     n285956 , n285957 , n285958 , n285959 , n285960 , n285961 , n285962 , n285963 , n285964 , n285965 , 
     n285966 , n285967 , n285968 , n285969 , n285970 , n285971 , n285972 , n285973 , n285974 , n285975 , 
     n285976 , n285977 , n285978 , n285979 , n285980 , n285981 , n285982 , n285983 , n285984 , n285985 , 
     n285986 , n285987 , n285988 , n285989 , n285990 , n285991 , n285992 , n285993 , n285994 , n285995 , 
     n285996 , n285997 , n285998 , n285999 , n286000 , n286001 , n286002 , n286003 , n286004 , n286005 , 
     n286006 , n286007 , n286008 , n286009 , n286010 , n286011 , n286012 , n286013 , n286014 , n286015 , 
     n286016 , n286017 , n286018 , n286019 , n286020 , n286021 , n286022 , n286023 , n286024 , n286025 , 
     n286026 , n286027 , n286028 , n286029 , n286030 , n286031 , n286032 , n286033 , n286034 , n286035 , 
     n286036 , n286037 , n286038 , n286039 , n286040 , n286041 , n286042 , n286043 , n286044 , n286045 , 
     n286046 , n286047 , n286048 , n286049 , n286050 , n286051 , n286052 , n286053 , n286054 , n286055 , 
     n286056 , n286057 , n286058 , n286059 , n286060 , n286061 , n286062 , n286063 , n286064 , n286065 , 
     n286066 , n286067 , n286068 , n286069 , n286070 , n286071 , n286072 , n286073 , n286074 , n286075 , 
     n286076 , n286077 , n286078 , n286079 , n286080 , n286081 , n286082 , n286083 , n286084 , n286085 , 
     n286086 , n286087 , n286088 , n286089 , n286090 , n286091 , n286092 , n286093 , n286094 , n286095 , 
     n286096 , n286097 , n286098 , n286099 , n286100 , n286101 , n286102 , n286103 , n286104 , n286105 , 
     n286106 , n286107 , n286108 , n286109 , n286110 , n286111 , n286112 , n286113 , n286114 , n286115 , 
     n286116 , n286117 , n286118 , n286119 , n286120 , n286121 , n286122 , n286123 , n286124 , n286125 , 
     n286126 , n286127 , n286128 , n286129 , n286130 , n286131 , n286132 , n286133 , n286134 , n286135 , 
     n286136 , n286137 , n286138 , n286139 , n286140 , n286141 , n286142 , n286143 , n286144 , n286145 , 
     n286146 , n286147 , n286148 , n286149 , n286150 , n286151 , n286152 , n286153 , n286154 , n286155 , 
     n286156 , n286157 , n286158 , n286159 , n286160 , n286161 , n286162 , n286163 , n286164 , n286165 , 
     n286166 , n286167 , n286168 , n286169 , n286170 , n286171 , n286172 , n286173 , n286174 , n286175 , 
     n286176 , n286177 , n286178 , n286179 , n286180 , n286181 , n286182 , n286183 , n286184 , n286185 , 
     n286186 , n286187 , n286188 , n286189 , n286190 , n286191 , n286192 , n286193 , n286194 , n286195 , 
     n286196 , n286197 , n286198 , n286199 , n286200 , n286201 , n286202 , n286203 , n286204 , n286205 , 
     n286206 , n286207 , n286208 , n286209 , n286210 , n286211 , n286212 , n286213 , n286214 , n286215 , 
     n286216 , n286217 , n286218 , n286219 , n286220 , n286221 , n286222 , n286223 , n286224 , n286225 , 
     n286226 , n286227 , n286228 , n286229 , n286230 , n286231 , n286232 , n286233 , n286234 , n286235 , 
     n286236 , n286237 , n286238 , n286239 , n286240 , n286241 , n286242 , n286243 , n286244 , n286245 , 
     n286246 , n286247 , n286248 , n286249 , n286250 , n286251 , n286252 , n286253 , n286254 , n286255 , 
     n286256 , n286257 , n286258 , n286259 , n286260 , n286261 , n286262 , n286263 , n286264 , n286265 , 
     n286266 , n286267 , n286268 , n286269 , n286270 , n286271 , n286272 , n286273 , n286274 , n286275 , 
     n286276 , n286277 , n286278 , n286279 , n286280 , n286281 , n286282 , n286283 , n286284 , n286285 , 
     n286286 , n286287 , n286288 , n286289 , n286290 , n286291 , n286292 , n286293 , n286294 , n286295 , 
     n286296 , n286297 , n286298 , n286299 , n286300 , n286301 , n286302 , n286303 , n286304 , n286305 , 
     n286306 , n286307 , n286308 , n286309 , n286310 , n286311 , n286312 , n286313 , n286314 , n286315 , 
     n286316 , n286317 , n286318 , n286319 , n286320 , n286321 , n286322 , n286323 , n286324 , n286325 , 
     n286326 , n286327 , n286328 , n286329 , n286330 , n286331 , n286332 , n286333 , n286334 , n286335 , 
     n286336 , n286337 , n286338 , n286339 , n286340 , n286341 , n286342 , n286343 , n286344 , n286345 , 
     n286346 , n286347 , n286348 , n286349 , n286350 , n286351 , n286352 , n286353 , n286354 , n286355 , 
     n286356 , n286357 , n286358 , n286359 , n286360 , n286361 , n286362 , n286363 , n286364 , n286365 , 
     n286366 , n286367 , n286368 , n286369 , n286370 , n286371 , n286372 , n286373 , n286374 , n286375 , 
     n286376 , n286377 , n286378 , n286379 , n286380 , n286381 , n286382 , n286383 , n286384 , n286385 , 
     n286386 , n286387 , n286388 , n286389 , n286390 , n286391 , n286392 , n286393 , n286394 , n286395 , 
     n286396 , n286397 , n286398 , n286399 , n286400 , n286401 , n286402 , n286403 , n286404 , n286405 , 
     n286406 , n286407 , n286408 , n286409 , n286410 , n286411 , n286412 , n286413 , n286414 , n286415 , 
     n286416 , n286417 , n286418 , n286419 , n286420 , n286421 , n286422 , n286423 , n286424 , n286425 , 
     n286426 , n286427 , n286428 , n286429 , n286430 , n286431 , n286432 , n286433 , n286434 , n286435 , 
     n286436 , n286437 , n286438 , n286439 , n286440 , n286441 , n286442 , n286443 , n286444 , n286445 , 
     n286446 , n286447 , n286448 , n286449 , n286450 , n286451 , n286452 , n286453 , n286454 , n286455 , 
     n286456 , n286457 , n286458 , n286459 , n286460 , n286461 , n286462 , n286463 , n286464 , n286465 , 
     n286466 , n286467 , n286468 , n286469 , n286470 , n286471 , n286472 , n286473 , n286474 , n286475 , 
     n286476 , n286477 , n286478 , n286479 , n286480 , n286481 , n286482 , n286483 , n286484 , n286485 , 
     n286486 , n286487 , n286488 , n286489 , n286490 , n286491 , n286492 , n286493 , n286494 , n286495 , 
     n286496 , n286497 , n286498 , n286499 , n286500 , n286501 , n286502 , n286503 , n286504 , n286505 , 
     n286506 , n286507 , n286508 , n286509 , n286510 , n286511 , n286512 , n286513 , n286514 , n286515 , 
     n286516 , n286517 , n286518 , n286519 , n286520 , n286521 , n286522 , n286523 , n286524 , n286525 , 
     n286526 , n286527 , n286528 , n286529 , n286530 , n286531 , n286532 , n286533 , n286534 , n286535 , 
     n286536 , n286537 , n286538 , n286539 , n286540 , n286541 , n286542 , n286543 , n286544 , n286545 , 
     n286546 , n286547 , n286548 , n286549 , n286550 , n286551 , n286552 , n286553 , n286554 , n286555 , 
     n286556 , n286557 , n286558 , n286559 , n286560 , n286561 , n286562 , n286563 , n286564 , n286565 , 
     n286566 , n286567 , n286568 , n286569 , n286570 , n286571 , n286572 , n286573 , n286574 , n286575 , 
     n286576 , n286577 , n286578 , n286579 , n286580 ;
buf ( RI19a22f70_2797 , n2 );
buf ( RI1754a798_67 , n3 );
buf ( RI19ad04a8_2209 , n5 );
buf ( RI19a23e70_2789 , n4 );
buf ( RI1754c610_2 , n6 );
buf ( RI19a23510_2794 , n1 );
buf ( RI19a859b8_2755 , n0 );
buf ( RI17534808_603 , n12 );
buf ( RI173f4d68_1562 , n453 );
buf ( RI173ac078_1917 , n452 );
buf ( RI17516358_697 , n454 );
buf ( RI1753aa78_586 , n9 );
buf ( RI19aad828_2471 , n449 );
buf ( RI17491398_1028 , n448 );
buf ( RI19ac0a40_2326 , n451 );
buf ( RI1751df18_673 , n450 );
buf ( RI173c95b0_1774 , n133 );
buf ( RI17340030_2129 , n132 );
buf ( RI174125e8_1418 , n134 );
buf ( RI19a8ffa8_2683 , n129 );
buf ( RI17465bf8_1240 , n128 );
buf ( RI19ac0680_2328 , n131 );
buf ( RI174ae8d0_885 , n130 );
buf ( RI1733be90_2149 , n455 );
buf ( RI173c9268_1775 , n461 );
buf ( RI173ff808_1510 , n460 );
buf ( RI173b67d0_1866 , n459 );
buf ( RI1752e610_622 , n458 );
buf ( RI1749baf0_977 , n456 );
buf ( RI19ab9a38_2383 , n457 );
buf ( RI173d4068_1722 , n467 );
buf ( RI1738b378_2077 , n466 );
buf ( RI1744bb40_1367 , n468 );
buf ( RI19a9c5f0_2595 , n463 );
buf ( RI17470350_1189 , n462 );
buf ( RI19acb828_2243 , n465 );
buf ( RI174b9460_834 , n464 );
buf ( RI173dd410_1677 , n469 );
buf ( RI173cee48_1747 , n475 );
buf ( RI17345580_2103 , n474 );
buf ( RI17446938_1392 , n476 );
buf ( RI19a8c498_2709 , n471 );
buf ( RI1746b148_1214 , n470 );
buf ( RI19abd890_2354 , n473 );
buf ( RI174b3e20_859 , n472 );
buf ( RI173ec398_1604 , n358 );
buf ( RI173a36a8_1959 , n357 );
buf ( RI1747e900_1119 , n359 );
buf ( RI19acf1d0_2217 , n356 );
buf ( RI17510160_716 , n355 );
buf ( RI19aa05b0_2566 , n354 );
buf ( RI17488680_1071 , n353 );
buf ( RI173895f0_2086 , n195 );
buf ( RI1740b9a0_1451 , n194 );
buf ( RI173c2cb0_1806 , n193 );
buf ( RI17339730_2161 , n192 );
buf ( RI174a7fd0_917 , n190 );
buf ( RI19ab3138_2431 , n191 );
buf ( RI19a95048_2647 , n617 );
buf ( RI1752a308_635 , n616 );
buf ( RI173ee468_1594 , n623 );
buf ( RI173a5778_1949 , n622 );
buf ( RI17493120_1019 , n624 );
buf ( RI19a9f548_2574 , n619 );
buf ( RI1748a750_1061 , n618 );
buf ( RI19ace168_2224 , n621 );
buf ( RI17513a18_705 , n620 );
buf ( RI173cd750_1754 , n638 );
buf ( RI173441d0_2109 , n637 );
buf ( RI17445588_1398 , n639 );
buf ( RI19a8dfc8_2697 , n634 );
buf ( RI17469d98_1220 , n633 );
buf ( RI19abeda8_2342 , n636 );
buf ( RI174b2a70_865 , n635 );
buf ( RI173bee58_1825 , n625 );
buf ( RI173f9250_1541 , n631 );
buf ( RI173b0560_1896 , n630 );
buf ( RI17389938_2085 , n632 );
buf ( RI19aadb70_2470 , n629 );
buf ( RI17524b60_652 , n628 );
buf ( RI19aab938_2485 , n627 );
buf ( RI17495880_1007 , n626 );
buf ( RI173e1268_1658 , n607 );
buf ( RI17398578_2013 , n606 );
buf ( RI17459088_1302 , n608 );
buf ( RI19a93d88_2655 , n603 );
buf ( RI1747d898_1124 , n602 );
buf ( RI19ac40a0_2299 , n605 );
buf ( RI174ce388_769 , n604 );
buf ( RI19a9e030_2584 , n601 );
buf ( RI1748be48_1054 , n600 );
buf ( RI173feae8_1514 , n614 );
buf ( RI173b5ab0_1870 , n613 );
buf ( RI173c0208_1819 , n615 );
buf ( RI19aa7c48_2511 , n610 );
buf ( RI1749add0_981 , n609 );
buf ( RI19a88e38_2732 , n612 );
buf ( RI1752d170_626 , n611 );
buf ( RI19a9bfd8_2598 , n484 );
buf ( RI1746f978_1192 , n483 );
buf ( RI1733b800_2151 , n255 );
buf ( RI173c4d80_1796 , n256 );
buf ( RI1740da70_1441 , n257 );
buf ( RI19ac21b0_2313 , n254 );
buf ( RI174aa0a0_907 , n253 );
buf ( RI19a91e98_2669 , n252 );
buf ( RI174613c8_1262 , n251 );
buf ( RI17399298_2009 , n262 );
buf ( RI173e1f88_1654 , n263 );
buf ( RI17459da8_1298 , n264 );
buf ( RI19a86c00_2747 , n261 );
buf ( RI174cf828_765 , n260 );
buf ( RI19aa5740_2526 , n259 );
buf ( RI1747e5b8_1120 , n258 );
buf ( RI173fda80_1519 , n567 );
buf ( RI173bc068_1839 , n565 );
buf ( RI17404d58_1484 , n566 );
buf ( RI17332ae8_2194 , n564 );
buf ( RI19ab5d48_2410 , n563 );
buf ( RI174a1040_951 , n562 );
buf ( RI173ad0e0_1912 , n554 );
buf ( RI173e7820_1627 , n560 );
buf ( RI1739e7e8_1983 , n559 );
buf ( RI1745f2f8_1272 , n561 );
buf ( RI19aa1d20_2554 , n556 );
buf ( RI17483b08_1094 , n555 );
buf ( RI19a82d30_2774 , n558 );
buf ( RI17508ac8_739 , n557 );
buf ( RI19a876c8_2742 , n539 );
buf ( RI174d1208_760 , n538 );
buf ( RI173d46f8_1720 , n545 );
buf ( RI1738ba08_2075 , n544 );
buf ( RI1744c1d0_1365 , n546 );
buf ( RI19a9ca28_2593 , n541 );
buf ( RI174709e0_1187 , n540 );
buf ( RI19acbc60_2241 , n543 );
buf ( RI174b9eb0_832 , n542 );
buf ( RI173a8f40_1932 , n551 );
buf ( RI173f1c30_1577 , n552 );
buf ( RI174b75e8_842 , n553 );
buf ( RI19ab0870_2450 , n548 );
buf ( RI1748df18_1044 , n547 );
buf ( RI19ac1d78_2315 , n550 );
buf ( RI175191c0_688 , n549 );
buf ( RI19abe6a0_2346 , n578 );
buf ( RI174b1d50_869 , n577 );
buf ( RI173db9d0_1685 , n590 );
buf ( RI17392ce0_2040 , n589 );
buf ( RI174534a8_1330 , n591 );
buf ( RI19ac7700_2274 , n588 );
buf ( RI174c5850_796 , n587 );
buf ( RI19a97820_2629 , n586 );
buf ( RI17478000_1151 , n585 );
buf ( RI174146b8_1408 , n584 );
buf ( RI17407170_1473 , n583 );
buf ( RI173be480_1828 , n582 );
buf ( RI17334f00_2183 , n581 );
buf ( RI174a3458_940 , n579 );
buf ( RI19ab4dd0_2417 , n580 );
buf ( RI1738ca70_2070 , n592 );
buf ( RI173c6b08_1787 , n598 );
buf ( RI1733d588_2142 , n597 );
buf ( RI1740f7f8_1432 , n599 );
buf ( RI19a90cc8_2677 , n594 );
buf ( RI17463150_1253 , n593 );
buf ( RI19ac1148_2322 , n596 );
buf ( RI174abe28_898 , n595 );
buf ( RI19aa48b8_2533 , n237 );
buf ( RI17480688_1110 , n236 );
buf ( RI19a85c10_2754 , n239 );
buf ( RI175019d0_755 , n238 );
buf ( RI173e4058_1644 , n241 );
buf ( RI1739b368_1999 , n240 );
buf ( RI1745be78_1288 , n242 );
buf ( RI19ab5f28_2409 , n569 );
buf ( RI174a1388_950 , n568 );
buf ( RI173f6460_1555 , n156 );
buf ( RI173ad770_1910 , n155 );
buf ( RI1752f060_620 , n157 );
buf ( RI19ab3c00_2425 , n154 );
buf ( RI17520330_666 , n153 );
buf ( RI19aac6d0_2480 , n152 );
buf ( RI17492a90_1021 , n151 );
buf ( RI173caca8_1767 , n575 );
buf ( RI17341728_2122 , n574 );
buf ( RI17413ce0_1411 , n576 );
buf ( RI19abf4b0_2338 , n573 );
buf ( RI174affc8_878 , n572 );
buf ( RI19a8e8b0_2693 , n571 );
buf ( RI174672f0_1233 , n570 );
buf ( RI19aac838_2479 , n346 );
buf ( RI17492dd8_1020 , n345 );
buf ( RI173e81f8_1624 , n531 );
buf ( RI1739f1c0_1980 , n530 );
buf ( RI1745fcd0_1269 , n532 );
buf ( RI19aa2248_2551 , n527 );
buf ( RI174844e0_1091 , n526 );
buf ( RI19a83438_2771 , n529 );
buf ( RI17509a40_736 , n528 );
buf ( RI174046c8_1486 , n537 );
buf ( RI17405730_1481 , n364 );
buf ( RI173bca40_1836 , n536 );
buf ( RI173334c0_2191 , n535 );
buf ( RI174a1a18_948 , n533 );
buf ( RI19ab63d8_2407 , n534 );
buf ( RI173a2cd0_1962 , n504 );
buf ( RI173dcd80_1679 , n510 );
buf ( RI17394090_2034 , n509 );
buf ( RI17454858_1324 , n511 );
buf ( RI19ac5e28_2285 , n508 );
buf ( RI174c7740_790 , n507 );
buf ( RI19a96038_2640 , n506 );
buf ( RI174793b0_1145 , n505 );
buf ( RI173fa2b8_1536 , n517 );
buf ( RI173b15c8_1891 , n516 );
buf ( RI17394db0_2030 , n518 );
buf ( RI19aa9d90_2497 , n513 );
buf ( RI174968e8_1002 , n512 );
buf ( RI19a9cc08_2592 , n515 );
buf ( RI17526528_647 , n514 );
buf ( RI19aa0358_2567 , n498 );
buf ( RI17488338_1072 , n497 );
buf ( RI19acef78_2218 , n500 );
buf ( RI1750fc38_717 , n499 );
buf ( RI173a3360_1960 , n501 );
buf ( RI173ec050_1605 , n502 );
buf ( RI1747c4e8_1130 , n503 );
buf ( RI19ac6080_2284 , n489 );
buf ( RI174c7c68_789 , n488 );
buf ( RI173ceb00_1748 , n495 );
buf ( RI17345238_2104 , n494 );
buf ( RI174465f0_1393 , n496 );
buf ( RI19abd6b0_2355 , n493 );
buf ( RI174b3ad8_860 , n492 );
buf ( RI19a8c240_2710 , n491 );
buf ( RI1746ae00_1215 , n490 );
buf ( RI19a8a2d8_2723 , n26 );
buf ( RI1746f630_1193 , n25 );
buf ( RI175361d0_598 , n482 );
buf ( RI1740d3e0_1443 , n481 );
buf ( RI173c46f0_1798 , n480 );
buf ( RI1733b170_2153 , n479 );
buf ( RI174a9a10_909 , n477 );
buf ( RI19ab1ef0_2440 , n478 );
buf ( RI173d3690_1725 , n486 );
buf ( RI1738a9a0_2080 , n485 );
buf ( RI1744b168_1370 , n487 );
buf ( RI19acb300_2246 , n250 );
buf ( RI174b8650_837 , n249 );
buf ( RI175385e8_592 , n521 );
buf ( RI17539218_590 , n520 );
buf ( RI17539e48_588 , n525 );
buf ( RI17537fd0_593 , n522 );
buf ( RI17536770_597 , n524 );
buf ( RI175379b8_594 , n523 );
buf ( RI17539830_589 , n519 );
buf ( RI174118c8_1422 , n723 );
buf ( RI173eda90_1597 , n729 );
buf ( RI17403318_1492 , n728 );
buf ( RI173ba628_1847 , n727 );
buf ( RI175342e0_604 , n726 );
buf ( RI19ab73c8_2400 , n725 );
buf ( RI1749f600_959 , n724 );
buf ( RI1744f650_1349 , n736 );
buf ( RI19a99f80_2612 , n731 );
buf ( RI17473e60_1171 , n730 );
buf ( RI19ac96e0_2259 , n733 );
buf ( RI174bf658_815 , n732 );
buf ( RI173d7b78_1704 , n735 );
buf ( RI1738ee88_2059 , n734 );
buf ( RI17400f00_1503 , n715 );
buf ( RI173f2608_1574 , n721 );
buf ( RI173a9918_1929 , n720 );
buf ( RI174be1b8_819 , n722 );
buf ( RI19aae7a0_2465 , n717 );
buf ( RI1748ec38_1040 , n716 );
buf ( RI19a23330_2795 , n719 );
buf ( RI1751a138_685 , n718 );
buf ( RI173ad428_1911 , n705 );
buf ( RI173e7b68_1626 , n709 );
buf ( RI1739eb30_1982 , n708 );
buf ( RI1745f640_1271 , n710 );
buf ( RI19a82f88_2773 , n143 );
buf ( RI17508ff0_738 , n142 );
buf ( RI19aa1f00_2553 , n707 );
buf ( RI17483e50_1093 , n706 );
buf ( RI173ffe98_1508 , n714 );
buf ( RI174050a0_1483 , n713 );
buf ( RI173bc3b0_1838 , n712 );
buf ( RI17332e30_2193 , n711 );
buf ( RI173e5750_1637 , n745 );
buf ( RI173f4048_1566 , n758 );
buf ( RI173ab358_1921 , n757 );
buf ( RI1750b408_731 , n759 );
buf ( RI19abcfa8_2359 , n756 );
buf ( RI1751ca78_677 , n755 );
buf ( RI19aad300_2474 , n754 );
buf ( RI17490678_1032 , n753 );
buf ( RI1744e5e8_1354 , n752 );
buf ( RI19acb120_2247 , n749 );
buf ( RI174bd768_821 , n748 );
buf ( RI19a9bd80_2599 , n747 );
buf ( RI17472df8_1176 , n746 );
buf ( RI173d6b10_1709 , n751 );
buf ( RI1738de20_2064 , n750 );
buf ( RI17497950_997 , n767 );
buf ( RI173eeaf8_1592 , n766 );
buf ( RI173a5e08_1947 , n765 );
buf ( RI19acc200_2238 , n764 );
buf ( RI17514468_703 , n763 );
buf ( RI19a9d400_2589 , n762 );
buf ( RI1748ade0_1059 , n761 );
buf ( RI173b2630_1886 , n760 );
buf ( RI173b6e60_1864 , n773 );
buf ( RI1740c030_1449 , n772 );
buf ( RI173c3340_1804 , n771 );
buf ( RI17339dc0_2159 , n770 );
buf ( RI19ab0ff0_2446 , n769 );
buf ( RI174a8660_915 , n768 );
buf ( RI1738cdb8_2069 , n737 );
buf ( RI173c7198_1785 , n743 );
buf ( RI1733dc18_2140 , n742 );
buf ( RI1740fe88_1430 , n744 );
buf ( RI19a90f20_2676 , n739 );
buf ( RI174637e0_1251 , n738 );
buf ( RI19ac12b0_2321 , n741 );
buf ( RI174ac4b8_896 , n740 );
buf ( RI173e43a0_1643 , n164 );
buf ( RI1739b6b0_1998 , n163 );
buf ( RI1745c1c0_1287 , n165 );
buf ( RI19a85e68_2753 , n162 );
buf ( RI17501ef8_754 , n161 );
buf ( RI19aa4a98_2532 , n160 );
buf ( RI174809d0_1109 , n159 );
buf ( RI173e4a30_1641 , n660 );
buf ( RI173f39b8_1568 , n666 );
buf ( RI173aacc8_1923 , n665 );
buf ( RI17502420_753 , n667 );
buf ( RI19a23150_2796 , n664 );
buf ( RI1751c028_679 , n663 );
buf ( RI19aaf628_2458 , n662 );
buf ( RI1748ffe8_1034 , n661 );
buf ( RI173c8200_1780 , n673 );
buf ( RI1733ec80_2135 , n672 );
buf ( RI17410ef0_1425 , n674 );
buf ( RI19ac1b98_2316 , n671 );
buf ( RI174ad520_891 , n670 );
buf ( RI19a919e8_2671 , n669 );
buf ( RI17464848_1246 , n668 );
buf ( RI173f6af0_1553 , n659 );
buf ( RI17404038_1488 , n658 );
buf ( RI173bb348_1843 , n657 );
buf ( RI17535780_600 , n656 );
buf ( RI174a0320_955 , n654 );
buf ( RI19ab7da0_2396 , n655 );
buf ( RI173f53f8_1560 , n653 );
buf ( RI173e6b00_1631 , n140 );
buf ( RI1739dac8_1987 , n139 );
buf ( RI1745e5d8_1276 , n141 );
buf ( RI19a84e00_2760 , n138 );
buf ( RI17507628_743 , n137 );
buf ( RI19aa3aa8_2540 , n136 );
buf ( RI17482de8_1098 , n135 );
buf ( RI173a3018_1961 , n640 );
buf ( RI173dd0c8_1678 , n644 );
buf ( RI173943d8_2033 , n643 );
buf ( RI17454ba0_1323 , n645 );
buf ( RI19a96290_2639 , n642 );
buf ( RI174796f8_1144 , n641 );
buf ( RI173b1910_1890 , n650 );
buf ( RI173fa600_1535 , n651 );
buf ( RI173971c8_2019 , n652 );
buf ( RI19a9e6c0_2581 , n649 );
buf ( RI17526a50_646 , n648 );
buf ( RI19aa9f70_2496 , n647 );
buf ( RI17496c30_1001 , n646 );
buf ( RI174a2dc8_942 , n704 );
buf ( RI173cf190_1746 , n695 );
buf ( RI173458c8_2102 , n694 );
buf ( RI17446c80_1391 , n696 );
buf ( RI19a8c6f0_2708 , n691 );
buf ( RI1746b490_1213 , n690 );
buf ( RI19abd9f8_2353 , n693 );
buf ( RI174b4168_858 , n692 );
buf ( RI173dd758_1676 , n689 );
buf ( RI173a39f0_1958 , n701 );
buf ( RI173ec6e0_1603 , n702 );
buf ( RI17480d18_1108 , n703 );
buf ( RI19acf428_2216 , n700 );
buf ( RI17510688_715 , n699 );
buf ( RI19aa0790_2565 , n698 );
buf ( RI174889c8_1070 , n697 );
buf ( RI1733c1d8_2148 , n675 );
buf ( RI173cb680_1764 , n681 );
buf ( RI173b6b18_1865 , n679 );
buf ( RI173ffb50_1509 , n680 );
buf ( RI1752eb38_621 , n678 );
buf ( RI1749be38_976 , n676 );
buf ( RI19ab9c18_2382 , n677 );
buf ( RI173d43b0_1721 , n687 );
buf ( RI1738b6c0_2076 , n686 );
buf ( RI1744be88_1366 , n688 );
buf ( RI19a9c848_2594 , n683 );
buf ( RI17470698_1188 , n682 );
buf ( RI19acba08_2242 , n685 );
buf ( RI174b9988_833 , n684 );
buf ( RI17450d48_1342 , n780 );
buf ( RI17408520_1467 , n779 );
buf ( RI173bf830_1822 , n778 );
buf ( RI173362b0_2177 , n777 );
buf ( RI174a4808_934 , n775 );
buf ( RI19ab34f8_2429 , n776 );
buf ( RI173ce470_1750 , n305 );
buf ( RI1744b7f8_1368 , n781 );
buf ( RI173c5410_1794 , n786 );
buf ( RI1740e100_1439 , n787 );
buf ( RI19a922d0_2667 , n783 );
buf ( RI17461a58_1260 , n782 );
buf ( RI19ac25e8_2311 , n785 );
buf ( RI174aa730_905 , n784 );
buf ( RI173e2960_1651 , n793 );
buf ( RI17399c70_2006 , n792 );
buf ( RI1745a780_1295 , n794 );
buf ( RI19a87218_2744 , n791 );
buf ( RI174d07a0_762 , n790 );
buf ( RI19aa5fb0_2523 , n789 );
buf ( RI1747ef90_1117 , n788 );
buf ( RI173ce128_1751 , n112 );
buf ( RI17344860_2107 , n111 );
buf ( RI17445c18_1396 , n113 );
buf ( RI19a8bbb0_2713 , n108 );
buf ( RI1746a428_1218 , n107 );
buf ( RI19abd188_2358 , n110 );
buf ( RI174b3100_863 , n109 );
buf ( RI173bf1a0_1824 , n774 );
buf ( RI19aabb90_2484 , n101 );
buf ( RI17495bc8_1006 , n100 );
buf ( RI19aaf448_2459 , n103 );
buf ( RI17525088_651 , n102 );
buf ( RI173f9598_1540 , n105 );
buf ( RI173b08a8_1895 , n104 );
buf ( RI1738bd50_2074 , n106 );
buf ( RI173fee30_1513 , n52 );
buf ( RI173b5df8_1869 , n51 );
buf ( RI173c2620_1808 , n53 );
buf ( RI1749b118_980 , n47 );
buf ( RI19aa7e28_2510 , n48 );
buf ( RI19a89e28_2725 , n50 );
buf ( RI1752d698_625 , n49 );
buf ( RI173a7500_1940 , n39 );
buf ( RI173988c0_2012 , n44 );
buf ( RI173e15b0_1657 , n45 );
buf ( RI174593d0_1301 , n46 );
buf ( RI19a93fe0_2654 , n41 );
buf ( RI1747dbe0_1123 , n40 );
buf ( RI19ac4280_2298 , n43 );
buf ( RI174ce8b0_768 , n42 );
buf ( RI17459a60_1299 , n38 );
buf ( RI17398f50_2010 , n36 );
buf ( RI173e1c40_1655 , n37 );
buf ( RI19a869a8_2748 , n35 );
buf ( RI174cf300_766 , n34 );
buf ( RI19aa5560_2527 , n33 );
buf ( RI1747e270_1121 , n32 );
buf ( RI173d3348_1726 , n30 );
buf ( RI1738a658_2081 , n29 );
buf ( RI1744ae20_1371 , n31 );
buf ( RI19abbe50_2368 , n28 );
buf ( RI174b8308_838 , n27 );
buf ( RI19ac4460_2297 , n24 );
buf ( RI174cedd8_767 , n23 );
buf ( RI173efea8_1586 , n15 );
buf ( RI17403660_1491 , n14 );
buf ( RI173ba970_1846 , n13 );
buf ( RI1749f948_958 , n10 );
buf ( RI19ab7530_2399 , n11 );
buf ( RI19a8fd50_2684 , n8 );
buf ( RI17465568_1242 , n7 );
buf ( RI1744f998_1348 , n22 );
buf ( RI19a9a160_2611 , n17 );
buf ( RI174741a8_1170 , n16 );
buf ( RI19ac9938_2258 , n19 );
buf ( RI174bfb80_814 , n18 );
buf ( RI173d7ec0_1703 , n21 );
buf ( RI1738f1d0_2058 , n20 );
buf ( RI17460d38_1264 , n98 );
buf ( RI17409f60_1459 , n97 );
buf ( RI173c1270_1814 , n96 );
buf ( RI17337cf0_2169 , n95 );
buf ( RI174a6590_925 , n93 );
buf ( RI19ab2148_2439 , n94 );
buf ( RI19aaa510_2493 , n85 );
buf ( RI17497608_998 , n84 );
buf ( RI173eca28_1602 , n91 );
buf ( RI173a3d38_1957 , n90 );
buf ( RI17483130_1097 , n92 );
buf ( RI19acf680_2215 , n89 );
buf ( RI17510bb0_714 , n88 );
buf ( RI19aa0970_2564 , n87 );
buf ( RI17488d10_1069 , n86 );
buf ( RI17335c20_2179 , n99 );
buf ( RI1745d570_1281 , n69 );
buf ( RI173d71a0_1707 , n75 );
buf ( RI1738e4b0_2062 , n74 );
buf ( RI1744ec78_1352 , n76 );
buf ( RI19a99698_2616 , n71 );
buf ( RI17473488_1174 , n70 );
buf ( RI19ac90c8_2262 , n73 );
buf ( RI174be6e0_818 , n72 );
buf ( RI173f4390_1565 , n82 );
buf ( RI173ab6a0_1920 , n81 );
buf ( RI1750ecc0_720 , n83 );
buf ( RI19abe2e0_2348 , n80 );
buf ( RI1751cfa0_676 , n79 );
buf ( RI19aad468_2473 , n78 );
buf ( RI174909c0_1031 , n77 );
buf ( RI19aa3238_2544 , n219 );
buf ( RI174820c8_1102 , n218 );
buf ( RI173d74e8_1706 , n225 );
buf ( RI1738e7f8_2061 , n224 );
buf ( RI1744efc0_1351 , n226 );
buf ( RI19ac92a8_2261 , n223 );
buf ( RI174bec08_817 , n222 );
buf ( RI19a998f0_2615 , n221 );
buf ( RI174737d0_1173 , n220 );
buf ( RI173f4a20_1563 , n232 );
buf ( RI173abd30_1918 , n231 );
buf ( RI17512aa0_708 , n233 );
buf ( RI19abf690_2337 , n230 );
buf ( RI1751d9f0_674 , n229 );
buf ( RI19aad648_2472 , n228 );
buf ( RI17491050_1029 , n227 );
buf ( RI173ddaa0_1675 , n248 );
buf ( RI174018d8_1500 , n247 );
buf ( RI173b8be8_1855 , n246 );
buf ( RI175319a0_612 , n245 );
buf ( RI1749dbc0_967 , n243 );
buf ( RI19ab8b38_2390 , n244 );
buf ( RI19a23678_2793 , n235 );
buf ( RI1751ab88_683 , n234 );
buf ( RI1744fce0_1347 , n203 );
buf ( RI173c98f8_1773 , n209 );
buf ( RI17340378_2128 , n208 );
buf ( RI17412930_1417 , n210 );
buf ( RI19a90188_2682 , n205 );
buf ( RI17465f40_1239 , n204 );
buf ( RI19ac0860_2327 , n207 );
buf ( RI174aec18_884 , n206 );
buf ( RI173e7190_1629 , n216 );
buf ( RI1739e158_1985 , n215 );
buf ( RI1745ec68_1274 , n217 );
buf ( RI19aa3c88_2539 , n212 );
buf ( RI17483478_1096 , n211 );
buf ( RI19a85058_2759 , n214 );
buf ( RI17508078_741 , n213 );
buf ( RI173cc6e8_1759 , n67 );
buf ( RI17343168_2114 , n66 );
buf ( RI17415720_1403 , n68 );
buf ( RI19a8d410_2702 , n63 );
buf ( RI17468d30_1225 , n62 );
buf ( RI19abe4c0_2347 , n65 );
buf ( RI174b1a08_870 , n64 );
buf ( RI1740fb40_1431 , n54 );
buf ( RI173f7ea0_1547 , n60 );
buf ( RI173af1b0_1902 , n59 );
buf ( RI1733d8d0_2141 , n61 );
buf ( RI19aa5a88_2525 , n58 );
buf ( RI17522c70_658 , n57 );
buf ( RI19aaac18_2490 , n56 );
buf ( RI174944d0_1013 , n55 );
buf ( RI17444ef8_1400 , n114 );
buf ( RI173dc060_1683 , n126 );
buf ( RI17393370_2038 , n125 );
buf ( RI17453b38_1328 , n127 );
buf ( RI19ac7b38_2272 , n124 );
buf ( RI174c62a0_794 , n123 );
buf ( RI19a97dc0_2627 , n122 );
buf ( RI17478690_1149 , n121 );
buf ( RI17447ce8_1386 , n120 );
buf ( RI17407800_1471 , n119 );
buf ( RI173beb10_1826 , n118 );
buf ( RI17335590_2181 , n117 );
buf ( RI174a3ae8_938 , n115 );
buf ( RI19ab52f8_2415 , n116 );
buf ( RI173d8f28_1698 , n149 );
buf ( RI17390238_2053 , n148 );
buf ( RI17450a00_1343 , n150 );
buf ( RI19a98630_2623 , n145 );
buf ( RI17475210_1165 , n144 );
buf ( RI19ac81c8_2269 , n147 );
buf ( RI174c1548_809 , n146 );
buf ( RI19ab4380_2422 , n173 );
buf ( RI174a5f00_927 , n172 );
buf ( RI173fac90_1533 , n179 );
buf ( RI173b1fa0_1888 , n178 );
buf ( RI1739b9f8_1997 , n180 );
buf ( RI19aa12d0_2559 , n177 );
buf ( RI175274a0_644 , n176 );
buf ( RI19aaa330_2494 , n175 );
buf ( RI174972c0_999 , n174 );
buf ( RI173cf820_1744 , n186 );
buf ( RI17345f58_2100 , n185 );
buf ( RI17447310_1389 , n187 );
buf ( RI19abddb8_2351 , n184 );
buf ( RI174b47f8_856 , n183 );
buf ( RI19a8cb28_2706 , n182 );
buf ( RI1746bb20_1211 , n181 );
buf ( RI19abcdc8_2360 , n189 );
buf ( RI174b6580_847 , n188 );
buf ( RI173e0200_1663 , n201 );
buf ( RI17397510_2018 , n200 );
buf ( RI17458020_1307 , n202 );
buf ( RI19ac3290_2305 , n199 );
buf ( RI174cc9c0_774 , n198 );
buf ( RI19a93068_2661 , n197 );
buf ( RI1747c830_1129 , n196 );
buf ( RI174c8be0_786 , n158 );
buf ( RI173dfeb8_1664 , n171 );
buf ( RI17401c20_1499 , n170 );
buf ( RI173b8f30_1854 , n169 );
buf ( RI17531ec8_611 , n168 );
buf ( RI1749df08_966 , n166 );
buf ( RI19ab8d90_2389 , n167 );
buf ( RI17453160_1331 , n291 );
buf ( RI17408868_1466 , n290 );
buf ( RI173bfb78_1821 , n289 );
buf ( RI173365f8_2176 , n288 );
buf ( RI174a4b50_933 , n286 );
buf ( RI19ab36d8_2428 , n287 );
buf ( RI173f9c28_1538 , n278 );
buf ( RI173eb330_1609 , n284 );
buf ( RI173a2640_1964 , n283 );
buf ( RI17475558_1164 , n285 );
buf ( RI19a9fae8_2571 , n280 );
buf ( RI17487618_1076 , n279 );
buf ( RI19ace870_2221 , n282 );
buf ( RI1750e798_721 , n281 );
buf ( RI173a7848_1939 , n265 );
buf ( RI17398c08_2011 , n268 );
buf ( RI173e18f8_1656 , n269 );
buf ( RI17459718_1300 , n270 );
buf ( RI19a94238_2653 , n267 );
buf ( RI1747df28_1122 , n266 );
buf ( RI174a9d58_908 , n277 );
buf ( RI173f0880_1583 , n276 );
buf ( RI173a7b90_1938 , n275 );
buf ( RI19aafad8_2456 , n272 );
buf ( RI1748cb68_1050 , n271 );
buf ( RI19a85508_2757 , n274 );
buf ( RI175172d0_694 , n273 );
buf ( RI17340a08_2126 , n307 );
buf ( RI173f8f08_1542 , n313 );
buf ( RI17404380_1487 , n312 );
buf ( RI173bb690_1842 , n311 );
buf ( RI17535ca8_599 , n310 );
buf ( RI174a0668_954 , n308 );
buf ( RI19ab7f80_2395 , n309 );
buf ( RI173d8be0_1699 , n319 );
buf ( RI1738fef0_2054 , n318 );
buf ( RI174506b8_1344 , n320 );
buf ( RI19a983d8_2624 , n315 );
buf ( RI17474ec8_1166 , n314 );
buf ( RI19ac7f70_2270 , n317 );
buf ( RI174c1020_810 , n316 );
buf ( RI173e2618_1652 , n334 );
buf ( RI17399928_2007 , n333 );
buf ( RI1745a438_1296 , n335 );
buf ( RI19a86fc0_2745 , n332 );
buf ( RI174d0278_763 , n331 );
buf ( RI19aa5dd0_2524 , n330 );
buf ( RI1747ec48_1118 , n329 );
buf ( RI173d39d8_1724 , n321 );
buf ( RI173c50c8_1795 , n327 );
buf ( RI1733bb48_2150 , n326 );
buf ( RI1740ddb8_1440 , n328 );
buf ( RI19ac2390_2312 , n325 );
buf ( RI174aa3e8_906 , n324 );
buf ( RI19a920f0_2668 , n323 );
buf ( RI17461710_1261 , n322 );
buf ( RI17335f68_2178 , n292 );
buf ( RI173b0bf0_1894 , n297 );
buf ( RI173f98e0_1539 , n298 );
buf ( RI1738e168_2063 , n299 );
buf ( RI19a981f8_2625 , n296 );
buf ( RI175255b0_650 , n295 );
buf ( RI19aa9688_2500 , n294 );
buf ( RI17495f10_1005 , n293 );
buf ( RI17344ba8_2106 , n304 );
buf ( RI17445f60_1395 , n306 );
buf ( RI19abd2f0_2357 , n303 );
buf ( RI174b3448_862 , n302 );
buf ( RI19a8be08_2712 , n301 );
buf ( RI1746a770_1217 , n300 );
buf ( RI173d2cb8_1728 , n441 );
buf ( RI17411f58_1420 , n447 );
buf ( RI173c4060_1800 , n445 );
buf ( RI1740cd50_1445 , n446 );
buf ( RI1733aae0_2155 , n444 );
buf ( RI174a9380_911 , n442 );
buf ( RI19ab1860_2442 , n443 );
buf ( RI173c39d0_1802 , n426 );
buf ( RI173fe110_1517 , n432 );
buf ( RI173b50d8_1873 , n431 );
buf ( RI173b95c0_1852 , n433 );
buf ( RI19a88460_2736 , n430 );
buf ( RI1752c1f8_629 , n429 );
buf ( RI19aa71f8_2515 , n428 );
buf ( RI1749a3f8_984 , n427 );
buf ( RI173d2970_1729 , n439 );
buf ( RI17389c80_2084 , n438 );
buf ( RI1744a448_1374 , n440 );
buf ( RI19a89888_2727 , n435 );
buf ( RI1746ec58_1196 , n434 );
buf ( RI19abb5e0_2372 , n437 );
buf ( RI174b7930_841 , n436 );
buf ( RI19a23858_2792 , n425 );
buf ( RI1751b0b0_682 , n424 );
buf ( RI173915e8_2047 , n394 );
buf ( RI173cb9c8_1763 , n400 );
buf ( RI17342448_2118 , n399 );
buf ( RI17414a00_1407 , n401 );
buf ( RI19a8f210_2689 , n396 );
buf ( RI17468010_1229 , n395 );
buf ( RI19abfc30_2334 , n398 );
buf ( RI174b0ce8_874 , n397 );
buf ( RI173e8f18_1620 , n407 );
buf ( RI1739fee0_1976 , n406 );
buf ( RI174609f0_1265 , n408 );
buf ( RI19aa2e78_2546 , n403 );
buf ( RI17485200_1087 , n402 );
buf ( RI19a83f78_2766 , n405 );
buf ( RI1750aee0_732 , n404 );
buf ( RI173e9f80_1615 , n409 );
buf ( RI173db340_1687 , n415 );
buf ( RI17392650_2042 , n414 );
buf ( RI17452e18_1332 , n416 );
buf ( RI19ac74a8_2275 , n413 );
buf ( RI174c4e00_798 , n412 );
buf ( RI19a976b8_2630 , n411 );
buf ( RI17477628_1154 , n410 );
buf ( RI173f8878_1544 , n422 );
buf ( RI173afb88_1899 , n421 );
buf ( RI17344518_2108 , n423 );
buf ( RI19aaa858_2492 , n420 );
buf ( RI17523be8_655 , n419 );
buf ( RI19aab410_2487 , n418 );
buf ( RI17494ea8_1010 , n417 );
buf ( RI19abaa28_2376 , n380 );
buf ( RI174b68c8_846 , n379 );
buf ( RI173a0228_1975 , n386 );
buf ( RI1740bce8_1450 , n385 );
buf ( RI173c2ff8_1805 , n384 );
buf ( RI17339a78_2160 , n383 );
buf ( RI19ab0e10_2447 , n382 );
buf ( RI174a8318_916 , n381 );
buf ( RI173e0548_1662 , n392 );
buf ( RI17397858_2017 , n391 );
buf ( RI17458368_1306 , n393 );
buf ( RI19ac34e8_2304 , n390 );
buf ( RI174ccee8_773 , n389 );
buf ( RI19a932c0_2660 , n388 );
buf ( RI1747cb78_1128 , n387 );
buf ( RI173b1c58_1889 , n352 );
buf ( RI174098d0_1461 , n362 );
buf ( RI173c0be0_1816 , n361 );
buf ( RI17337660_2171 , n360 );
buf ( RI1745c508_1286 , n363 );
buf ( RI173f6e38_1552 , n370 );
buf ( RI173ae148_1907 , n369 );
buf ( RI17332458_2196 , n371 );
buf ( RI19aaca18_2478 , n366 );
buf ( RI17493468_1018 , n365 );
buf ( RI19ab6cc0_2403 , n368 );
buf ( RI175212a8_663 , n367 );
buf ( RI173cb338_1765 , n377 );
buf ( RI17341db8_2120 , n376 );
buf ( RI17414370_1409 , n378 );
buf ( RI19a8efb8_2690 , n373 );
buf ( RI17467980_1231 , n372 );
buf ( RI19abfa50_2335 , n375 );
buf ( RI174b0658_876 , n374 );
buf ( RI19a831e0_2772 , n337 );
buf ( RI17509518_737 , n336 );
buf ( RI173d95b8_1696 , n343 );
buf ( RI173908c8_2051 , n342 );
buf ( RI17451090_1341 , n344 );
buf ( RI19ac8330_2268 , n341 );
buf ( RI174c1f98_807 , n340 );
buf ( RI19a98888_2622 , n339 );
buf ( RI174758a0_1163 , n338 );
buf ( RI19ab54d8_2414 , n348 );
buf ( RI17520858_665 , n347 );
buf ( RI173f67a8_1554 , n350 );
buf ( RI173adab8_1909 , n349 );
buf ( RI17532918_609 , n351 );
buf ( RI17411238_1424 , n817 );
buf ( RI173e9260_1619 , n823 );
buf ( RI17402c88_1494 , n822 );
buf ( RI173b9f98_1849 , n821 );
buf ( RI17533890_606 , n820 );
buf ( RI1749ef70_961 , n818 );
buf ( RI19ab7008_2402 , n819 );
buf ( RI17400870_1505 , n809 );
buf ( RI173c6478_1789 , n815 );
buf ( RI1733cef8_2144 , n814 );
buf ( RI1740f168_1434 , n816 );
buf ( RI19ac30b0_2306 , n813 );
buf ( RI174ab798_900 , n812 );
buf ( RI19a92e10_2662 , n811 );
buf ( RI17462ac0_1255 , n810 );
buf ( RI173acd98_1913 , n795 );
buf ( RI173e74d8_1628 , n801 );
buf ( RI1739e4a0_1984 , n800 );
buf ( RI1745efb0_1273 , n802 );
buf ( RI19aa3ee0_2538 , n797 );
buf ( RI174837c0_1095 , n796 );
buf ( RI19a852b0_2758 , n799 );
buf ( RI175085a0_740 , n798 );
buf ( RI173fb668_1530 , n808 );
buf ( RI17404a10_1485 , n807 );
buf ( RI173bbd20_1840 , n806 );
buf ( RI173327a0_2195 , n805 );
buf ( RI174a0cf8_952 , n803 );
buf ( RI19ab5a00_2411 , n804 );
buf ( RI1733f9a0_2131 , n866 );
buf ( RI173c8f20_1776 , n867 );
buf ( RI17411c10_1421 , n868 );
buf ( RI19ac04a0_2329 , n865 );
buf ( RI174ae240_887 , n864 );
buf ( RI173c6e50_1786 , n874 );
buf ( RI173b6488_1867 , n872 );
buf ( RI173ff4c0_1511 , n873 );
buf ( RI1752e0e8_623 , n871 );
buf ( RI1749b7a8_978 , n869 );
buf ( RI19ab98d0_2384 , n870 );
buf ( RI173d3d20_1723 , n880 );
buf ( RI1738b030_2078 , n879 );
buf ( RI19acb648_2244 , n878 );
buf ( RI174b8f38_835 , n877 );
buf ( RI19a9c398_2596 , n876 );
buf ( RI17470008_1190 , n875 );
buf ( RI173f22c0_1575 , n863 );
buf ( RI174039a8_1490 , n862 );
buf ( RI173bacb8_1845 , n861 );
buf ( RI17534d30_602 , n860 );
buf ( RI1749fc90_957 , n858 );
buf ( RI19ab7878_2398 , n859 );
buf ( RI173e6470_1633 , n856 );
buf ( RI1739d438_1989 , n855 );
buf ( RI1745df48_1278 , n857 );
buf ( RI19a84950_2762 , n854 );
buf ( RI17506bd8_745 , n853 );
buf ( RI19aa3580_2542 , n852 );
buf ( RI17482758_1100 , n851 );
buf ( RI173f9f70_1537 , n849 );
buf ( RI173b1280_1892 , n848 );
buf ( RI17392998_2041 , n850 );
buf ( RI19a9b420_2603 , n847 );
buf ( RI17526000_648 , n846 );
buf ( RI19aa9bb0_2498 , n845 );
buf ( RI174965a0_1003 , n844 );
buf ( RI173dca38_1680 , n842 );
buf ( RI17393d48_2035 , n841 );
buf ( RI17454510_1325 , n843 );
buf ( RI19a95de0_2641 , n838 );
buf ( RI17479068_1146 , n837 );
buf ( RI174c7218_791 , n839 );
buf ( RI19ac5bd0_2286 , n840 );
buf ( RI173ebd08_1606 , n835 );
buf ( RI1747a0d0_1141 , n836 );
buf ( RI19aa0100_2568 , n832 );
buf ( RI17487ff0_1073 , n831 );
buf ( RI19aced20_2219 , n834 );
buf ( RI1750f710_718 , n833 );
buf ( RI173ce7b8_1749 , n829 );
buf ( RI17344ef0_2105 , n828 );
buf ( RI174462a8_1394 , n830 );
buf ( RI19a8bfe8_2711 , n825 );
buf ( RI1746aab8_1216 , n824 );
buf ( RI19abd4d0_2356 , n827 );
buf ( RI174b3790_861 , n826 );
buf ( RI173cd408_1755 , n945 );
buf ( RI17343e88_2110 , n944 );
buf ( RI17445240_1399 , n946 );
buf ( RI19a8dd70_2698 , n941 );
buf ( RI17469a50_1221 , n940 );
buf ( RI19abebc8_2343 , n943 );
buf ( RI174b2728_866 , n942 );
buf ( RI173f8bc0_1543 , n938 );
buf ( RI173afed0_1898 , n937 );
buf ( RI17346930_2097 , n939 );
buf ( RI19aac388_2481 , n936 );
buf ( RI17524110_654 , n935 );
buf ( RI19aab5f0_2486 , n934 );
buf ( RI174951f0_1009 , n933 );
buf ( RI173dc6f0_1681 , n956 );
buf ( RI17393a00_2036 , n955 );
buf ( RI174541c8_1326 , n957 );
buf ( RI19a95b88_2642 , n952 );
buf ( RI17478d20_1147 , n951 );
buf ( RI19ac5978_2287 , n954 );
buf ( RI174c6cf0_792 , n953 );
buf ( RI17407e90_1469 , n949 );
buf ( RI1744c518_1364 , n950 );
buf ( RI19ab5820_2412 , n948 );
buf ( RI174a4178_936 , n947 );
buf ( RI17332110_2197 , n932 );
buf ( RI1740b658_1452 , n931 );
buf ( RI173c2968_1807 , n930 );
buf ( RI19ab2f58_2432 , n928 );
buf ( RI174a7c88_918 , n927 );
buf ( RI173393e8_2162 , n929 );
buf ( RI19a93518_2659 , n919 );
buf ( RI17529de0_636 , n918 );
buf ( RI173a5430_1950 , n924 );
buf ( RI173ee120_1595 , n925 );
buf ( RI17490d08_1030 , n926 );
buf ( RI19a9f368_2575 , n921 );
buf ( RI1748a408_1062 , n920 );
buf ( RI19acdf10_2225 , n923 );
buf ( RI175134f0_706 , n922 );
buf ( RI19a87470_2743 , n882 );
buf ( RI174d0cc8_761 , n881 );
buf ( RI173f18e8_1578 , n888 );
buf ( RI173a8bf8_1933 , n887 );
buf ( RI174b51d0_853 , n889 );
buf ( RI19ab0528_2451 , n884 );
buf ( RI1748dbd0_1045 , n883 );
buf ( RI19ab3a20_2426 , n886 );
buf ( RI17518c98_689 , n885 );
buf ( RI174122a0_1419 , n895 );
buf ( RI173be138_1829 , n893 );
buf ( RI17406e28_1474 , n894 );
buf ( RI17334bb8_2184 , n892 );
buf ( RI19ab4bf0_2418 , n891 );
buf ( RI174a3110_941 , n890 );
buf ( RI1738c728_2071 , n896 );
buf ( RI173c67c0_1788 , n902 );
buf ( RI1733d240_2143 , n901 );
buf ( RI1740f4b0_1433 , n903 );
buf ( RI19a90a70_2678 , n898 );
buf ( RI17462e08_1254 , n897 );
buf ( RI19ac0f68_2323 , n900 );
buf ( RI174abae0_899 , n899 );
buf ( RI173e3d10_1645 , n908 );
buf ( RI1739b020_2000 , n907 );
buf ( RI1745bb30_1289 , n909 );
buf ( RI175014a8_756 , n906 );
buf ( RI19aa46d8_2534 , n905 );
buf ( RI17480340_1111 , n904 );
buf ( RI173e50c0_1639 , n910 );
buf ( RI173d6480_1711 , n916 );
buf ( RI1738d790_2066 , n915 );
buf ( RI1744df58_1356 , n917 );
buf ( RI19acadd8_2249 , n914 );
buf ( RI174bcd18_823 , n913 );
buf ( RI19a9b8d0_2601 , n912 );
buf ( RI17472768_1178 , n911 );
buf ( RI17400bb8_1504 , n1002 );
buf ( RI173f1f78_1576 , n1008 );
buf ( RI173a9288_1931 , n1007 );
buf ( RI174ba3d8_831 , n1009 );
buf ( RI19ab0a50_2449 , n1004 );
buf ( RI1748e260_1043 , n1003 );
buf ( RI19ad0238_2210 , n1006 );
buf ( RI175196e8_687 , n1005 );
buf ( RI173eb678_1608 , n1016 );
buf ( RI173ba2e0_1848 , n1014 );
buf ( RI17402fd0_1493 , n1015 );
buf ( RI17533db8_605 , n1013 );
buf ( RI1749f2b8_960 , n1011 );
buf ( RI19ab71e8_2401 , n1012 );
buf ( RI17411580_1423 , n1010 );
buf ( RI173d7830_1705 , n1022 );
buf ( RI1738eb40_2060 , n1021 );
buf ( RI1744f308_1350 , n1023 );
buf ( RI19ac9500_2260 , n1020 );
buf ( RI174bf130_816 , n1019 );
buf ( RI19a99d28_2613 , n1018 );
buf ( RI17473b18_1172 , n1017 );
buf ( RI173b0218_1897 , n1039 );
buf ( RI173ee7b0_1593 , n1045 );
buf ( RI173a5ac0_1948 , n1044 );
buf ( RI17495538_1008 , n1046 );
buf ( RI19ace3c0_2223 , n1043 );
buf ( RI17513f40_704 , n1042 );
buf ( RI19a9f728_2573 , n1041 );
buf ( RI1748aa98_1060 , n1040 );
buf ( RI173e5408_1638 , n1024 );
buf ( RI173f3d00_1567 , n1037 );
buf ( RI173ab010_1922 , n1036 );
buf ( RI17507b50_742 , n1038 );
buf ( RI19aaf790_2457 , n1033 );
buf ( RI17490330_1033 , n1032 );
buf ( RI19a83b40_2768 , n1035 );
buf ( RI1751c550_678 , n1034 );
buf ( RI1744e2a0_1355 , n1031 );
buf ( RI173d67c8_1710 , n1030 );
buf ( RI1738dad8_2065 , n1029 );
buf ( RI19acaf40_2248 , n1028 );
buf ( RI174bd240_822 , n1027 );
buf ( RI19a9bb28_2600 , n1026 );
buf ( RI17472ab0_1177 , n1025 );
buf ( RI1744b4b0_1369 , n1052 );
buf ( RI1744e930_1353 , n1051 );
buf ( RI174081d8_1468 , n1050 );
buf ( RI173bf4e8_1823 , n1049 );
buf ( RI174a44c0_935 , n1047 );
buf ( RI19ab3318_2430 , n1048 );
buf ( RI173f50b0_1561 , n958 );
buf ( RI173e67b8_1632 , n964 );
buf ( RI1739d780_1988 , n963 );
buf ( RI1745e290_1277 , n965 );
buf ( RI19a84ba8_2761 , n962 );
buf ( RI17507100_744 , n961 );
buf ( RI19aa38c8_2541 , n960 );
buf ( RI17482aa0_1099 , n959 );
buf ( RI173f46d8_1564 , n971 );
buf ( RI17403cf0_1489 , n970 );
buf ( RI173bb000_1844 , n969 );
buf ( RI17535258_601 , n968 );
buf ( RI1749ffd8_956 , n966 );
buf ( RI19ab7a58_2397 , n967 );
buf ( RI173e22d0_1653 , n972 );
buf ( RI173f3670_1569 , n978 );
buf ( RI173aa980_1924 , n977 );
buf ( RI174cfd50_764 , n979 );
buf ( RI19a23c18_2790 , n976 );
buf ( RI1751bb00_680 , n975 );
buf ( RI19aaf268_2460 , n974 );
buf ( RI1748fca0_1035 , n973 );
buf ( RI173c7eb8_1781 , n985 );
buf ( RI1733e938_2136 , n984 );
buf ( RI17410ba8_1426 , n986 );
buf ( RI19a91808_2672 , n981 );
buf ( RI17464500_1247 , n980 );
buf ( RI19ac1a30_2317 , n983 );
buf ( RI174ad1d8_892 , n982 );
buf ( RI173e0f20_1659 , n993 );
buf ( RI17398230_2014 , n992 );
buf ( RI17458d40_1303 , n994 );
buf ( RI19ac3d58_2300 , n991 );
buf ( RI174cde60_770 , n990 );
buf ( RI19a93ba8_2656 , n989 );
buf ( RI1747d550_1125 , n988 );
buf ( RI174a09b0_953 , n987 );
buf ( RI173fe7a0_1515 , n1000 );
buf ( RI173b5768_1871 , n999 );
buf ( RI173bddf0_1830 , n1001 );
buf ( RI19a88be0_2733 , n998 );
buf ( RI1752cc48_627 , n997 );
buf ( RI19aa7a68_2512 , n996 );
buf ( RI1749aa88_982 , n995 );
buf ( RI173ac708_1915 , n1253 );
buf ( RI1751d4c8_675 , n1254 );
buf ( RI19ac36c8_2303 , n1252 );
buf ( RI1751e968_671 , n1251 );
buf ( RI19aadfa8_2468 , n1250 );
buf ( RI17491a28_1026 , n1249 );
buf ( RI173e2ff0_1649 , n1247 );
buf ( RI1739a300_2004 , n1246 );
buf ( RI1745ae10_1293 , n1248 );
buf ( RI19aa62f8_2521 , n1245 );
buf ( RI1747f620_1115 , n1244 );
buf ( RI173c5aa0_1792 , n1242 );
buf ( RI1733c520_2147 , n1241 );
buf ( RI1740e790_1437 , n1243 );
buf ( RI19a92708_2665 , n1238 );
buf ( RI174620e8_1258 , n1237 );
buf ( RI19ac2a98_2309 , n1240 );
buf ( RI174aadc0_903 , n1239 );
buf ( RI173d9900_1695 , n1235 );
buf ( RI17390c10_2050 , n1234 );
buf ( RI19ac8510_2267 , n1233 );
buf ( RI174c24c0_806 , n1232 );
buf ( RI19a98ae0_2621 , n1231 );
buf ( RI17475be8_1162 , n1230 );
buf ( RI174513d8_1340 , n1236 );
buf ( RI173413e0_2123 , n1229 );
buf ( RI17337318_2172 , n1180 );
buf ( RI1745a0f0_1297 , n1183 );
buf ( RI174a5bb8_928 , n1103 );
buf ( RI19ab4038_2423 , n1104 );
buf ( RI173c0898_1817 , n1181 );
buf ( RI17409588_1462 , n1182 );
buf ( RI173f1258_1580 , n1271 );
buf ( RI173a8568_1935 , n1270 );
buf ( RI174b09a0_875 , n1272 );
buf ( RI19a94df0_2648 , n1269 );
buf ( RI17518248_691 , n1268 );
buf ( RI19ab01e0_2453 , n1267 );
buf ( RI1748d540_1047 , n1266 );
buf ( RI173c5758_1793 , n1259 );
buf ( RI1740e448_1438 , n1260 );
buf ( RI19a92528_2666 , n1256 );
buf ( RI17461da0_1259 , n1255 );
buf ( RI19ac2840_2310 , n1258 );
buf ( RI174aaa78_904 , n1257 );
buf ( RI173e2ca8_1650 , n1264 );
buf ( RI17399fb8_2005 , n1263 );
buf ( RI1745aac8_1294 , n1265 );
buf ( RI19aa6190_2522 , n1262 );
buf ( RI1747f2d8_1116 , n1261 );
buf ( RI17336940_2175 , n1273 );
buf ( RI173c43a8_1799 , n1348 );
buf ( RI173c4a38_1797 , n1354 );
buf ( RI173ff178_1512 , n1353 );
buf ( RI173b6140_1868 , n1352 );
buf ( RI1752dbc0_624 , n1351 );
buf ( RI1749b460_979 , n1349 );
buf ( RI19ab96f0_2385 , n1350 );
buf ( RI1738ace8_2079 , n1359 );
buf ( RI19acb4e0_2245 , n1358 );
buf ( RI174b8a10_836 , n1357 );
buf ( RI19a9c1b8_2597 , n1356 );
buf ( RI1746fcc0_1191 , n1355 );
buf ( RI1739c3d0_1994 , n1340 );
buf ( RI1745cee0_1283 , n1341 );
buf ( RI19a864f8_2750 , n1339 );
buf ( RI17503398_750 , n1338 );
buf ( RI19aa5218_2529 , n1337 );
buf ( RI174816f0_1105 , n1336 );
buf ( RI17402940_1495 , n1346 );
buf ( RI173b9c50_1850 , n1345 );
buf ( RI17533368_607 , n1344 );
buf ( RI173e6e48_1630 , n1347 );
buf ( RI19ab9498_2386 , n1343 );
buf ( RI1749ec28_962 , n1342 );
buf ( RI19a838e8_2769 , n1138 );
buf ( RI1750a490_734 , n1137 );
buf ( RI173d9f90_1693 , n1278 );
buf ( RI173912a0_2048 , n1185 );
buf ( RI17451a68_1338 , n1279 );
buf ( RI19a98f90_2619 , n1275 );
buf ( RI17476278_1160 , n1274 );
buf ( RI19ac89c0_2265 , n1277 );
buf ( RI174c2f10_804 , n1276 );
buf ( RI173f74c8_1550 , n1285 );
buf ( RI173ae7d8_1905 , n1284 );
buf ( RI17336c88_2174 , n1286 );
buf ( RI19aacdd8_2476 , n1281 );
buf ( RI17493af8_1016 , n1280 );
buf ( RI19ab9df8_2381 , n1283 );
buf ( RI17521cf8_661 , n1282 );
buf ( RI173b2978_1885 , n1287 );
buf ( RI17485548_1086 , n1294 );
buf ( RI19a9e8a0_2580 , n1289 );
buf ( RI17489058_1068 , n1288 );
buf ( RI19acd358_2230 , n1291 );
buf ( RI175110d8_713 , n1290 );
buf ( RI173ecd70_1601 , n1293 );
buf ( RI173a4080_1956 , n1292 );
buf ( RI17477970_1153 , n1300 );
buf ( RI1740a2a8_1458 , n1299 );
buf ( RI173c15b8_1813 , n1298 );
buf ( RI17338038_2168 , n1297 );
buf ( RI174a68d8_924 , n1295 );
buf ( RI19ab2328_2438 , n1296 );
buf ( RI17406108_1478 , n1301 );
buf ( RI173aeb20_1904 , n1306 );
buf ( RI173f7810_1549 , n1307 );
buf ( RI173390a0_2163 , n1308 );
buf ( RI19aad120_2475 , n1303 );
buf ( RI17493e40_1015 , n1302 );
buf ( RI19abba90_2370 , n1305 );
buf ( RI17522220_660 , n1304 );
buf ( RI173cc058_1761 , n1314 );
buf ( RI17342ad8_2116 , n1313 );
buf ( RI17415090_1405 , n1315 );
buf ( RI19a8cd80_2705 , n1310 );
buf ( RI174686a0_1227 , n1309 );
buf ( RI19abdf98_2350 , n1312 );
buf ( RI174b1378_872 , n1311 );
buf ( RI19abb298_2373 , n1219 );
buf ( RI174b72a0_843 , n1218 );
buf ( RI173e46e8_1642 , n1320 );
buf ( RI1740c6c0_1447 , n1319 );
buf ( RI1733a450_2157 , n1318 );
buf ( RI174a8cf0_913 , n1316 );
buf ( RI19ab1518_2444 , n1317 );
buf ( RI17391fc0_2044 , n1321 );
buf ( RI173cc3a0_1760 , n1327 );
buf ( RI17342e20_2115 , n1326 );
buf ( RI174153d8_1404 , n1328 );
buf ( RI19a8cfd8_2704 , n1323 );
buf ( RI174689e8_1226 , n1322 );
buf ( RI19abe100_2349 , n1325 );
buf ( RI174b16c0_871 , n1324 );
buf ( RI173a0f48_1971 , n1333 );
buf ( RI173e9c38_1616 , n1193 );
buf ( RI174658b0_1241 , n1334 );
buf ( RI19acfd88_2212 , n1332 );
buf ( RI1750c380_728 , n1331 );
buf ( RI19aa0f10_2561 , n1330 );
buf ( RI17485f20_1083 , n1329 );
buf ( RI173ea958_1612 , n1335 );
buf ( RI173fa948_1534 , n1109 );
buf ( RI1744a100_1375 , n1360 );
buf ( RI19a8e220_2696 , n1362 );
buf ( RI17466918_1236 , n1361 );
buf ( RI173d8208_1702 , n1382 );
buf ( RI1738f518_2057 , n1381 );
buf ( RI19ac9b90_2257 , n1380 );
buf ( RI174c00a8_813 , n1379 );
buf ( RI19a9a3b8_2610 , n1378 );
buf ( RI174744f0_1169 , n1377 );
buf ( RI173f5740_1559 , n1388 );
buf ( RI173aca50_1914 , n1387 );
buf ( RI17520d80_664 , n1389 );
buf ( RI19aae110_2467 , n1384 );
buf ( RI17491d70_1025 , n1383 );
buf ( RI19ac4f28_2292 , n1386 );
buf ( RI1751ee90_670 , n1385 );
buf ( RI19aa8bc0_2505 , n1391 );
buf ( RI174989b8_992 , n1390 );
buf ( RI173a50e8_1951 , n1396 );
buf ( RI173eddd8_1596 , n1397 );
buf ( RI1748e8f0_1041 , n1398 );
buf ( RI19acdcb8_2226 , n1395 );
buf ( RI17512fc8_707 , n1394 );
buf ( RI19a9f188_2576 , n1393 );
buf ( RI1748a0c0_1063 , n1392 );
buf ( RI17512578_709 , n1404 );
buf ( RI1740afc8_1454 , n1403 );
buf ( RI173c22d8_1809 , n1402 );
buf ( RI17338d58_2164 , n1401 );
buf ( RI19ab2d78_2433 , n1400 );
buf ( RI174a75f8_920 , n1399 );
buf ( RI173c5de8_1791 , n1368 );
buf ( RI1733c868_2146 , n1367 );
buf ( RI1740ead8_1436 , n1369 );
buf ( RI19ac2cf0_2308 , n1366 );
buf ( RI174ab108_902 , n1365 );
buf ( RI19a92960_2664 , n1364 );
buf ( RI17462430_1257 , n1363 );
buf ( RI173e3338_1648 , n1375 );
buf ( RI1739a648_2003 , n1374 );
buf ( RI1745b158_1292 , n1376 );
buf ( RI19a87920_2741 , n1373 );
buf ( RI17500530_759 , n1372 );
buf ( RI19aa6640_2520 , n1371 );
buf ( RI1747f968_1114 , n1370 );
buf ( RI173f5a88_1558 , n1462 );
buf ( RI17524638_653 , n1463 );
buf ( RI19aae458_2466 , n1459 );
buf ( RI174920b8_1024 , n1458 );
buf ( RI19ac6878_2281 , n1461 );
buf ( RI1751f3b8_669 , n1460 );
buf ( RI17450028_1346 , n1090 );
buf ( RI19ac9de8_2256 , n1087 );
buf ( RI174c05d0_812 , n1086 );
buf ( RI19a9a610_2609 , n1085 );
buf ( RI17474838_1168 , n1084 );
buf ( RI173d8550_1701 , n1089 );
buf ( RI1738f860_2056 , n1088 );
buf ( RI173ca960_1768 , n1456 );
buf ( RI17413998_1412 , n1457 );
buf ( RI19abf2d0_2339 , n1455 );
buf ( RI174afc80_879 , n1454 );
buf ( RI19a8e6d0_2694 , n1453 );
buf ( RI17466fa8_1234 , n1452 );
buf ( RI173ca618_1769 , n1418 );
buf ( RI17341098_2124 , n1417 );
buf ( RI17413650_1413 , n1419 );
buf ( RI19abf0f0_2340 , n1416 );
buf ( RI174af938_880 , n1415 );
buf ( RI19a8e478_2695 , n1414 );
buf ( RI17466c60_1235 , n1413 );
buf ( RI173e7eb0_1625 , n1423 );
buf ( RI1739ee78_1981 , n1422 );
buf ( RI1745f988_1270 , n1424 );
buf ( RI19aa2068_2552 , n1421 );
buf ( RI17484198_1092 , n1420 );
buf ( RI17406450_1477 , n1405 );
buf ( RI173f7b58_1548 , n1411 );
buf ( RI173aee68_1903 , n1410 );
buf ( RI1733b4b8_2152 , n1412 );
buf ( RI19aaaa38_2491 , n1407 );
buf ( RI17494188_1014 , n1406 );
buf ( RI19aa4318_2536 , n1409 );
buf ( RI17522748_659 , n1408 );
buf ( RI19ab29b8_2435 , n1437 );
buf ( RI174a6f68_922 , n1436 );
buf ( RI173fc388_1526 , n1443 );
buf ( RI173b3350_1882 , n1442 );
buf ( RI173a71b8_1941 , n1444 );
buf ( RI19a90368_2681 , n1441 );
buf ( RI17529390_638 , n1440 );
buf ( RI19aa8878_2506 , n1439 );
buf ( RI17498670_993 , n1438 );
buf ( RI173d0bd0_1738 , n1450 );
buf ( RI17347308_2094 , n1449 );
buf ( RI174486c0_1383 , n1451 );
buf ( RI19a8af08_2718 , n1446 );
buf ( RI1746ced0_1205 , n1445 );
buf ( RI19abc8a0_2363 , n1448 );
buf ( RI174b5ba8_850 , n1447 );
buf ( RI1739ca60_1992 , n1434 );
buf ( RI173e5a98_1636 , n1435 );
buf ( RI19a841d0_2765 , n1433 );
buf ( RI17503de8_748 , n1432 );
buf ( RI19aa3058_2545 , n1143 );
buf ( RI17481d80_1103 , n1142 );
buf ( RI173eaca0_1611 , n1073 );
buf ( RI173dc3a8_1682 , n1430 );
buf ( RI173936b8_2037 , n1429 );
buf ( RI17453e80_1327 , n1431 );
buf ( RI19ac7d90_2271 , n1428 );
buf ( RI174c67c8_793 , n1427 );
buf ( RI19a98018_2626 , n1426 );
buf ( RI174789d8_1148 , n1425 );
buf ( RI173406c0_2127 , n1172 );
buf ( RI17450370_1345 , n1179 );
buf ( RI19aca040_2255 , n1176 );
buf ( RI174c0af8_811 , n1175 );
buf ( RI19a9a868_2608 , n1174 );
buf ( RI17474b80_1167 , n1173 );
buf ( RI173d8898_1700 , n1178 );
buf ( RI1738fba8_2055 , n1177 );
buf ( RI173a22f8_1965 , n1169 );
buf ( RI173eafe8_1610 , n1170 );
buf ( RI17473140_1175 , n1171 );
buf ( RI19a9f908_2572 , n1166 );
buf ( RI174872d0_1077 , n1165 );
buf ( RI19ace618_2222 , n1168 );
buf ( RI1750e270_722 , n1167 );
buf ( RI173fb320_1531 , n1228 );
buf ( RI1740ca08_1446 , n1227 );
buf ( RI173c3d18_1801 , n1226 );
buf ( RI1733a798_2156 , n1225 );
buf ( RI174a9038_912 , n1223 );
buf ( RI19ab16f8_2443 , n1224 );
buf ( RI173c3688_1803 , n1208 );
buf ( RI173fddc8_1518 , n1214 );
buf ( RI173b4d90_1874 , n1213 );
buf ( RI173b71a8_1863 , n1215 );
buf ( RI19a88208_2737 , n1212 );
buf ( RI1752bcd0_630 , n1211 );
buf ( RI19aa7090_2516 , n1210 );
buf ( RI1749a0b0_985 , n1209 );
buf ( RI173d22e0_1731 , n1221 );
buf ( RI173892a8_2087 , n1220 );
buf ( RI17449db8_1376 , n1222 );
buf ( RI19a89720_2728 , n1217 );
buf ( RI1746e5c8_1198 , n1216 );
buf ( RI173daff8_1688 , n1199 );
buf ( RI17392308_2043 , n1198 );
buf ( RI17452ad0_1333 , n1200 );
buf ( RI19ac7250_2276 , n1197 );
buf ( RI174c48d8_799 , n1196 );
buf ( RI19a97460_2631 , n1195 );
buf ( RI174772e0_1155 , n1194 );
buf ( RI173f8530_1545 , n1206 );
buf ( RI173af840_1900 , n1205 );
buf ( RI17342100_2119 , n1207 );
buf ( RI19aa8f80_2503 , n1204 );
buf ( RI175236c0_656 , n1203 );
buf ( RI19aab0c8_2488 , n1202 );
buf ( RI17494b60_1011 , n1201 );
buf ( RI173e8bd0_1621 , n1191 );
buf ( RI1739fb98_1977 , n1190 );
buf ( RI174606a8_1266 , n1192 );
buf ( RI19aa2c20_2547 , n1187 );
buf ( RI17484eb8_1088 , n1186 );
buf ( RI19a83d20_2767 , n1189 );
buf ( RI1750a9b8_733 , n1188 );
buf ( RI173caff0_1766 , n1133 );
buf ( RI17341a70_2121 , n1132 );
buf ( RI17414028_1410 , n1134 );
buf ( RI19a8ed60_2691 , n1129 );
buf ( RI17467638_1232 , n1128 );
buf ( RI19abf870_2336 , n1131 );
buf ( RI174b0310_877 , n1130 );
buf ( RI174053e8_1482 , n1184 );
buf ( RI173a6e70_1942 , n1067 );
buf ( RI173a1fb0_1966 , n1072 );
buf ( RI17470d28_1186 , n1074 );
buf ( RI19aa19d8_2555 , n1069 );
buf ( RI17486f88_1078 , n1068 );
buf ( RI19a82b50_2775 , n1071 );
buf ( RI1750dd48_723 , n1070 );
buf ( RI173f0538_1584 , n1065 );
buf ( RI19acd100_2231 , n1064 );
buf ( RI17516da8_695 , n1063 );
buf ( RI19a9e468_2582 , n1062 );
buf ( RI1748c820_1051 , n1061 );
buf ( RI174a7940_919 , n1066 );
buf ( RI173d3000_1727 , n1059 );
buf ( RI1738a310_2082 , n1058 );
buf ( RI1744aad8_1372 , n1060 );
buf ( RI19abbc70_2369 , n1057 );
buf ( RI174b7fc0_839 , n1056 );
buf ( RI19a8a080_2724 , n1055 );
buf ( RI1746f2e8_1194 , n1054 );
buf ( RI17457cd8_1308 , n1102 );
buf ( RI17409240_1463 , n1101 );
buf ( RI173c0550_1818 , n1100 );
buf ( RI17336fd0_2173 , n1099 );
buf ( RI174a5870_929 , n1097 );
buf ( RI19ab3de0_2424 , n1098 );
buf ( RI173f6118_1556 , n1095 );
buf ( RI1752b7a8_631 , n1096 );
buf ( RI19ab2508_2437 , n1094 );
buf ( RI1751fe08_667 , n1093 );
buf ( RI19aac040_2482 , n1092 );
buf ( RI17492748_1022 , n1091 );
buf ( RI173db688_1686 , n1150 );
buf ( RI173b88a0_1856 , n1148 );
buf ( RI17401590_1501 , n1149 );
buf ( RI17531478_613 , n1147 );
buf ( RI1749d878_968 , n1145 );
buf ( RI19ab8958_2391 , n1146 );
buf ( RI1751a660_684 , n1144 );
buf ( RI19a88028_2738 , n1154 );
buf ( RI1752b280_632 , n1153 );
buf ( RI19aa6d48_2517 , n1152 );
buf ( RI17499a20_987 , n1151 );
buf ( RI173fd738_1520 , n1156 );
buf ( RI173b4700_1876 , n1155 );
buf ( RI173b4a48_1875 , n1157 );
buf ( RI173d1f98_1732 , n1163 );
buf ( RI173599e0_2088 , n1162 );
buf ( RI17449a70_1377 , n1164 );
buf ( RI19a894c8_2729 , n1159 );
buf ( RI1746e280_1199 , n1158 );
buf ( RI19abaf50_2374 , n1161 );
buf ( RI174b6f58_844 , n1160 );
buf ( RI19abcbe8_2361 , n1119 );
buf ( RI174b6238_848 , n1118 );
buf ( RI173dfb70_1665 , n1125 );
buf ( RI17396e80_2020 , n1124 );
buf ( RI17457648_1310 , n1126 );
buf ( RI19a95930_2643 , n1121 );
buf ( RI1747c1a0_1131 , n1120 );
buf ( RI19ac5720_2288 , n1123 );
buf ( RI174cbf70_776 , n1122 );
buf ( RI17390f58_2049 , n1127 );
buf ( RI173e8888_1622 , n1140 );
buf ( RI1739f850_1978 , n1139 );
buf ( RI17460360_1267 , n1141 );
buf ( RI19aa27e8_2549 , n1136 );
buf ( RI17484b70_1089 , n1135 );
buf ( RI173cf4d8_1745 , n1116 );
buf ( RI17345c10_2101 , n1115 );
buf ( RI17446fc8_1390 , n1117 );
buf ( RI19a8c948_2707 , n1112 );
buf ( RI1746b7d8_1212 , n1111 );
buf ( RI19abdbd8_2352 , n1114 );
buf ( RI174b44b0_857 , n1113 );
buf ( RI173995e0_2008 , n1110 );
buf ( RI19a9fcc8_2570 , n1108 );
buf ( RI17526f78_645 , n1107 );
buf ( RI19aaa150_2495 , n1106 );
buf ( RI17496f78_1000 , n1105 );
buf ( RI173358d8_2180 , n1083 );
buf ( RI17409c18_1460 , n1081 );
buf ( RI173c0f28_1815 , n1080 );
buf ( RI173379a8_2170 , n1079 );
buf ( RI1745e920_1275 , n1082 );
buf ( RI174a6248_926 , n1077 );
buf ( RI19ab4560_2421 , n1078 );
buf ( RI19a8faf8_2685 , n1076 );
buf ( RI17465220_1243 , n1075 );
buf ( RI1740a5f0_1457 , n1464 );
buf ( RI173fc040_1527 , n1470 );
buf ( RI173b3008_1883 , n1469 );
buf ( RI173a4da0_1952 , n1471 );
buf ( RI19aa8530_2507 , n1466 );
buf ( RI17498328_994 , n1465 );
buf ( RI19a8eb08_2692 , n1468 );
buf ( RI17528e68_639 , n1467 );
buf ( RI173d0888_1739 , n1477 );
buf ( RI17346fc0_2095 , n1476 );
buf ( RI17448378_1384 , n1478 );
buf ( RI19a8acb0_2719 , n1473 );
buf ( RI1746cb88_1206 , n1472 );
buf ( RI19abc6c0_2364 , n1475 );
buf ( RI174b5860_851 , n1474 );
buf ( RI1733fce8_2130 , n1513 );
buf ( RI173eee40_1591 , n1512 );
buf ( RI173964a8_2023 , n1511 );
buf ( RI173cdde0_1752 , n1510 );
buf ( RI174001e0_1507 , n1509 );
buf ( RI173b74f0_1862 , n1508 );
buf ( RI1752f588_619 , n1507 );
buf ( RI1749c4c8_974 , n1505 );
buf ( RI19aba050_2380 , n1506 );
buf ( RI173d1c50_1733 , n1490 );
buf ( RI17359698_2089 , n1489 );
buf ( RI17449728_1378 , n1491 );
buf ( RI19a89270_2730 , n1486 );
buf ( RI1746df38_1200 , n1485 );
buf ( RI19abad70_2375 , n1488 );
buf ( RI174b6c10_845 , n1487 );
buf ( RI173fd3f0_1521 , n1484 );
buf ( RI173b43b8_1877 , n1483 );
buf ( RI19a87dd0_2739 , n1482 );
buf ( RI1752ad58_633 , n1481 );
buf ( RI19aa6b68_2518 , n1480 );
buf ( RI174996d8_988 , n1479 );
buf ( RI173c9f88_1771 , n1503 );
buf ( RI17412fc0_1415 , n1504 );
buf ( RI19ac0d88_2324 , n1502 );
buf ( RI174af2a8_882 , n1501 );
buf ( RI19a90818_2679 , n1500 );
buf ( RI174665d0_1237 , n1499 );
buf ( RI173ddde8_1674 , n1497 );
buf ( RI173950f8_2029 , n1496 );
buf ( RI174558c0_1319 , n1498 );
buf ( RI19a96bf0_2635 , n1493 );
buf ( RI1747a418_1140 , n1492 );
buf ( RI19ac69e0_2280 , n1495 );
buf ( RI174c9108_785 , n1494 );
buf ( RI173c8bd8_1777 , n1517 );
buf ( RI1733f658_2132 , n1516 );
buf ( RI19ac0338_2330 , n1515 );
buf ( RI174adef8_888 , n1514 );
buf ( RI17454ee8_1322 , n1518 );
buf ( RI17455578_1320 , n1523 );
buf ( RI17408bb0_1465 , n1522 );
buf ( RI173bfec0_1820 , n1521 );
buf ( RI174a4e98_932 , n1519 );
buf ( RI19ab3840_2427 , n1520 );
buf ( RI17394720_2032 , n1528 );
buf ( RI19a964e8_2638 , n1525 );
buf ( RI17479a40_1143 , n1524 );
buf ( RI19ac63c8_2283 , n1527 );
buf ( RI174c8190_788 , n1526 );
buf ( RI173d6e58_1708 , n1546 );
buf ( RI173b8210_1858 , n1545 );
buf ( RI17530a28_615 , n1544 );
buf ( RI1749d1e8_970 , n1542 );
buf ( RI19ab82c8_2394 , n1543 );
buf ( RI1739a990_2002 , n1539 );
buf ( RI173e3680_1647 , n1540 );
buf ( RI1745b4a0_1291 , n1541 );
buf ( RI19a87b78_2740 , n1538 );
buf ( RI17500a58_758 , n1537 );
buf ( RI19aa6988_2519 , n1536 );
buf ( RI1747fcb0_1113 , n1535 );
buf ( RI173b0f38_1893 , n1533 );
buf ( RI17390580_2052 , n1534 );
buf ( RI19a99ad0_2614 , n1532 );
buf ( RI17525ad8_649 , n1531 );
buf ( RI19aa9868_2499 , n1530 );
buf ( RI17496258_1004 , n1529 );
buf ( RI19aa7540_2514 , n1573 );
buf ( RI17523198_657 , n1572 );
buf ( RI17455230_1321 , n1571 );
buf ( RI19acd5b0_2229 , n1549 );
buf ( RI17511600_712 , n1548 );
buf ( RI17395ad0_2026 , n1554 );
buf ( RI173de7c0_1671 , n1555 );
buf ( RI17456298_1316 , n1556 );
buf ( RI19a946e8_2651 , n1551 );
buf ( RI1747adf0_1137 , n1550 );
buf ( RI19ac4910_2295 , n1553 );
buf ( RI174ca080_782 , n1552 );
buf ( RI1744a790_1373 , n1547 );
buf ( RI1749cb58_972 , n1569 );
buf ( RI19aba578_2378 , n1570 );
buf ( RI173a1290_1970 , n1561 );
buf ( RI17467cc8_1230 , n1562 );
buf ( RI19aa10f0_2560 , n1558 );
buf ( RI17486268_1082 , n1557 );
buf ( RI19acffe0_2211 , n1560 );
buf ( RI1750c8a8_727 , n1559 );
buf ( RI174458d0_1397 , n1568 );
buf ( RI174074b8_1472 , n1567 );
buf ( RI173be7c8_1827 , n1566 );
buf ( RI19ab5118_2416 , n1564 );
buf ( RI174a37a0_939 , n1563 );
buf ( RI17335248_2182 , n1565 );
buf ( RI1733f310_2133 , n1053 );
buf ( RI19a9e288_2583 , n1649 );
buf ( RI1748c4d8_1052 , n1648 );
buf ( RI19a96998_2636 , n1657 );
buf ( RI1752a830_634 , n1656 );
buf ( RI173ac3c0_1916 , n1585 );
buf ( RI17519c10_686 , n1586 );
buf ( RI19aadd50_2469 , n1582 );
buf ( RI174916e0_1027 , n1581 );
buf ( RI19ac1f58_2314 , n1584 );
buf ( RI1751e440_672 , n1583 );
buf ( RI17406ae0_1475 , n1708 );
buf ( RI17405a78_1480 , n1707 );
buf ( RI173bcd88_1835 , n1706 );
buf ( RI17333808_2190 , n1705 );
buf ( RI174a1d60_947 , n1703 );
buf ( RI19ab65b8_2406 , n1704 );
buf ( RI173e8540_1623 , n1701 );
buf ( RI1739f508_1979 , n1700 );
buf ( RI17460018_1268 , n1702 );
buf ( RI19aa24a0_2550 , n1697 );
buf ( RI17484828_1090 , n1696 );
buf ( RI19a83690_2770 , n1699 );
buf ( RI17509f68_735 , n1698 );
buf ( RI175373a0_595 , n1795 );
buf ( RI1753a460_587 , n1794 );
buf ( RI19abe808_2345 , n1777 );
buf ( RI174b2098_868 , n1776 );
buf ( RI173dbd18_1684 , n1803 );
buf ( RI17393028_2039 , n1802 );
buf ( RI174537f0_1329 , n1804 );
buf ( RI19a97b68_2628 , n1799 );
buf ( RI17478348_1150 , n1798 );
buf ( RI19ac7958_2273 , n1801 );
buf ( RI174c5d78_795 , n1800 );
buf ( RI19ab6090_2408 , n1797 );
buf ( RI174a16d0_949 , n1796 );
buf ( RI1744c860_1363 , n1793 );
buf ( RI19acbe40_2240 , n1790 );
buf ( RI174ba900_830 , n1789 );
buf ( RI19a9ce60_2591 , n1788 );
buf ( RI17471070_1185 , n1787 );
buf ( RI173d4d88_1718 , n1792 );
buf ( RI1738c098_2073 , n1791 );
buf ( RI173c9c40_1772 , n1669 );
buf ( RI17412c78_1416 , n1670 );
buf ( RI19ac0ba8_2325 , n1668 );
buf ( RI174aef60_883 , n1667 );
buf ( RI19a905c0_2680 , n1666 );
buf ( RI17466288_1238 , n1665 );
buf ( RI173d4a40_1719 , n1713 );
buf ( RI173b7ec8_1859 , n1712 );
buf ( RI17530500_616 , n1711 );
buf ( RI1749cea0_971 , n1709 );
buf ( RI19aba8c0_2377 , n1710 );
buf ( RI173d5418_1716 , n1718 );
buf ( RI1744cef0_1361 , n1719 );
buf ( RI19a9aac0_2607 , n1715 );
buf ( RI17471700_1183 , n1714 );
buf ( RI19aca298_2254 , n1717 );
buf ( RI174bb350_828 , n1716 );
buf ( RI173df198_1668 , n1734 );
buf ( RI19a9b1c8_2604 , n1728 );
buf ( RI174720d8_1180 , n1727 );
buf ( RI19aca9a0_2251 , n1730 );
buf ( RI174bc2c8_825 , n1729 );
buf ( RI173d5df0_1713 , n1732 );
buf ( RI1738d100_2068 , n1731 );
buf ( RI1744d8c8_1358 , n1733 );
buf ( RI173a4710_1954 , n1720 );
buf ( RI173deb08_1670 , n1725 );
buf ( RI17395e18_2025 , n1628 );
buf ( RI174565e0_1315 , n1726 );
buf ( RI19ac4b68_2294 , n1724 );
buf ( RI174ca5a8_781 , n1723 );
buf ( RI19a94940_2650 , n1722 );
buf ( RI1747b138_1136 , n1721 );
buf ( RI173cfb68_1743 , n1758 );
buf ( RI1744d238_1360 , n1759 );
buf ( RI17461080_1263 , n1741 );
buf ( RI173a08b8_1973 , n1739 );
buf ( RI173e95a8_1618 , n1740 );
buf ( RI19acf8d8_2214 , n1738 );
buf ( RI1750b930_730 , n1737 );
buf ( RI19aa0b50_2563 , n1736 );
buf ( RI17485890_1085 , n1735 );
buf ( RI173bdaa8_1831 , n1745 );
buf ( RI17406798_1476 , n1746 );
buf ( RI17334528_2186 , n1744 );
buf ( RI174a2a80_943 , n1742 );
buf ( RI19ab48a8_2419 , n1743 );
buf ( RI173c8548_1779 , n1579 );
buf ( RI1733efc8_2134 , n1578 );
buf ( RI19a8f648_2687 , n1575 );
buf ( RI17464b90_1245 , n1574 );
buf ( RI19abff78_2332 , n1577 );
buf ( RI174ad868_890 , n1576 );
buf ( RI19a8f8a0_2686 , n1748 );
buf ( RI17464ed8_1244 , n1747 );
buf ( RI19ac0158_2331 , n1750 );
buf ( RI174adbb0_889 , n1749 );
buf ( RI173c8890_1778 , n1580 );
buf ( RI173e6128_1634 , n1756 );
buf ( RI1739d0f0_1990 , n1755 );
buf ( RI1745dc00_1279 , n1757 );
buf ( RI19aa3418_2543 , n1752 );
buf ( RI17482410_1101 , n1751 );
buf ( RI19a846f8_2763 , n1754 );
buf ( RI175066b0_746 , n1753 );
buf ( RI1744d580_1359 , n1786 );
buf ( RI173d5760_1715 , n1764 );
buf ( RI19aca4f0_2253 , n1763 );
buf ( RI174bb878_827 , n1762 );
buf ( RI19a9ad18_2606 , n1761 );
buf ( RI17471a48_1182 , n1760 );
buf ( RI19ac5108_2291 , n1766 );
buf ( RI174caff8_779 , n1765 );
buf ( RI173ea2c8_1614 , n1772 );
buf ( RI173a15d8_1969 , n1771 );
buf ( RI1746a0e0_1219 , n1773 );
buf ( RI19aa1438_2558 , n1768 );
buf ( RI174865b0_1081 , n1767 );
buf ( RI19a82538_2778 , n1770 );
buf ( RI1750cdd0_726 , n1769 );
buf ( RI173ccd78_1757 , n1779 );
buf ( RI173437f8_2112 , n1778 );
buf ( RI17444bb0_1401 , n1780 );
buf ( RI19a8d8c0_2700 , n1775 );
buf ( RI174693c0_1223 , n1774 );
buf ( RI17394a68_2031 , n1785 );
buf ( RI19ac6620_2282 , n1784 );
buf ( RI174c86b8_787 , n1783 );
buf ( RI19a96740_2637 , n1782 );
buf ( RI17479d88_1142 , n1781 );
buf ( RI173a4a58_1953 , n1640 );
buf ( RI173ed748_1598 , n1641 );
buf ( RI1748c190_1053 , n1642 );
buf ( RI19a9efa8_2577 , n1637 );
buf ( RI17489a30_1065 , n1636 );
buf ( RI19acda60_2227 , n1639 );
buf ( RI17512050_710 , n1638 );
buf ( RI173d0540_1740 , n1634 );
buf ( RI17346c78_2096 , n1633 );
buf ( RI17448030_1385 , n1635 );
buf ( RI19a8aad0_2720 , n1630 );
buf ( RI1746c840_1207 , n1629 );
buf ( RI19abc4e0_2365 , n1632 );
buf ( RI174b5518_852 , n1631 );
buf ( RI19ac1670_2319 , n1627 );
buf ( RI174acb48_894 , n1626 );
buf ( RI173cfeb0_1742 , n1624 );
buf ( RI173465e8_2098 , n1623 );
buf ( RI174479a0_1387 , n1625 );
buf ( RI19a8a878_2721 , n1620 );
buf ( RI1746c1b0_1209 , n1619 );
buf ( RI19abc378_2366 , n1622 );
buf ( RI174b4e88_854 , n1621 );
buf ( RI173fb9b0_1529 , n1617 );
buf ( RI173a0570_1974 , n1618 );
buf ( RI19a8b958_2714 , n1616 );
buf ( RI17528418_641 , n1615 );
buf ( RI19aa8080_2509 , n1614 );
buf ( RI17497c98_996 , n1613 );
buf ( RI173a7ed8_1937 , n1612 );
buf ( RI173fafd8_1532 , n1610 );
buf ( RI173b22e8_1887 , n1609 );
buf ( RI1739de10_1986 , n1611 );
buf ( RI19aa29c8_2548 , n1608 );
buf ( RI175279c8_643 , n1607 );
buf ( RI173fe458_1516 , n1600 );
buf ( RI173b5420_1872 , n1599 );
buf ( RI173bb9d8_1841 , n1601 );
buf ( RI19a88a00_2734 , n1598 );
buf ( RI1752c720_628 , n1597 );
buf ( RI19aa7888_2513 , n1596 );
buf ( RI1749a740_983 , n1595 );
buf ( RI17389fc8_2083 , n1606 );
buf ( RI19abb748_2371 , n1605 );
buf ( RI174b7c78_840 , n1604 );
buf ( RI19a89bd0_2726 , n1603 );
buf ( RI1746efa0_1195 , n1602 );
buf ( RI173efb60_1587 , n1589 );
buf ( RI19accc50_2233 , n1588 );
buf ( RI17515e30_698 , n1587 );
buf ( RI17457990_1309 , n1594 );
buf ( RI1740d098_1444 , n1593 );
buf ( RI1733ae28_2154 , n1592 );
buf ( RI174a96c8_910 , n1590 );
buf ( RI19ab1ba8_2441 , n1591 );
buf ( RI1740d728_1442 , n1647 );
buf ( RI173bd760_1832 , n1646 );
buf ( RI173341e0_2187 , n1645 );
buf ( RI174a2738_944 , n1643 );
buf ( RI19ab4740_2420 , n1644 );
buf ( RI173fbcf8_1528 , n1680 );
buf ( RI173b2cc0_1884 , n1679 );
buf ( RI173a2988_1963 , n1681 );
buf ( RI19aa81e8_2508 , n1676 );
buf ( RI17497fe0_995 , n1675 );
buf ( RI19a8d230_2703 , n1678 );
buf ( RI17528940_640 , n1677 );
buf ( RI173e98f0_1617 , n1687 );
buf ( RI173a0c00_1972 , n1686 );
buf ( RI17463498_1252 , n1688 );
buf ( RI19acfb30_2213 , n1685 );
buf ( RI1750be58_729 , n1684 );
buf ( RI19aa0d30_2562 , n1683 );
buf ( RI17485bd8_1084 , n1682 );
buf ( RI173f15a0_1579 , n1694 );
buf ( RI173a88b0_1934 , n1693 );
buf ( RI174b2db8_864 , n1695 );
buf ( RI19aa40c0_2537 , n1692 );
buf ( RI17518770_690 , n1691 );
buf ( RI19ab03c0_2452 , n1690 );
buf ( RI1748d888_1046 , n1689 );
buf ( RI173d2628_1730 , n1674 );
buf ( RI173b7b80_1860 , n1673 );
buf ( RI1752ffd8_617 , n1672 );
buf ( RI1746e910_1197 , n1671 );
buf ( RI174a5528_930 , n1653 );
buf ( RI19accea8_2232 , n1651 );
buf ( RI17516880_696 , n1650 );
buf ( RI173f01f0_1585 , n1652 );
buf ( RI173fd0a8_1522 , n1659 );
buf ( RI173b4070_1878 , n1658 );
buf ( RI19aa9430_2501 , n1655 );
buf ( RI17499390_989 , n1654 );
buf ( RI173d1908_1734 , n1663 );
buf ( RI17359350_2090 , n1662 );
buf ( RI174493e0_1379 , n1664 );
buf ( RI19a89018_2731 , n1661 );
buf ( RI1746dbf0_1201 , n1660 );
buf ( RI17514990_702 , n1805 );
buf ( RI19a9ed50_2578 , n1913 );
buf ( RI174896e8_1066 , n1912 );
buf ( RI173bc6f8_1837 , n1914 );
buf ( RI17487960_1075 , n1930 );
buf ( RI173df4e0_1667 , n1926 );
buf ( RI173967f0_2022 , n1904 );
buf ( RI17456fb8_1312 , n1927 );
buf ( RI19a954f8_2645 , n1923 );
buf ( RI1747bb10_1133 , n1922 );
buf ( RI19ac52e8_2290 , n1925 );
buf ( RI174cb520_778 , n1924 );
buf ( RI174bdc90_820 , n1833 );
buf ( RI1740ac80_1455 , n1832 );
buf ( RI173c1f90_1810 , n1831 );
buf ( RI17338a10_2165 , n1830 );
buf ( RI174a72b0_921 , n1828 );
buf ( RI19ab2b98_2434 , n1829 );
buf ( RI19ac6e18_2278 , n1929 );
buf ( RI174c3e88_801 , n1928 );
buf ( RI173a8220_1936 , n1919 );
buf ( RI173f0f10_1581 , n1920 );
buf ( RI174ae588_886 , n1921 );
buf ( RI19a887a8_2735 , n1918 );
buf ( RI17517d20_692 , n1917 );
buf ( RI19ab0000_2454 , n1916 );
buf ( RI1748d1f8_1048 , n1915 );
buf ( RI17457300_1311 , n1940 );
buf ( RI19a8b4a8_2716 , n1942 );
buf ( RI1746d560_1203 , n1941 );
buf ( RI173d1278_1736 , n1944 );
buf ( RI17358cc0_2092 , n1943 );
buf ( RI17448d50_1381 , n1945 );
buf ( RI19abef88_2341 , n1865 );
buf ( RI174af5f0_881 , n1864 );
buf ( RI1740ee20_1435 , n1892 );
buf ( RI173d50d0_1717 , n1936 );
buf ( RI1738c3e0_2072 , n1935 );
buf ( RI1744cba8_1362 , n1937 );
buf ( RI19acc020_2239 , n1934 );
buf ( RI174bae28_829 , n1933 );
buf ( RI19a9d1a8_2590 , n1932 );
buf ( RI174713b8_1184 , n1931 );
buf ( RI173d0f18_1737 , n1910 );
buf ( RI17347650_2093 , n1909 );
buf ( RI17448a08_1382 , n1911 );
buf ( RI19abca80_2362 , n1908 );
buf ( RI174b5ef0_849 , n1907 );
buf ( RI19a8b250_2717 , n1906 );
buf ( RI1746d218_1204 , n1905 );
buf ( RI19acc5c0_2236 , n1939 );
buf ( RI17514eb8_701 , n1938 );
buf ( RI173e0890_1661 , n1882 );
buf ( RI17397ba0_2016 , n1881 );
buf ( RI174586b0_1305 , n1883 );
buf ( RI19ac3920_2302 , n1880 );
buf ( RI174cd410_772 , n1879 );
buf ( RI19a936f8_2658 , n1878 );
buf ( RI1747cec0_1127 , n1877 );
buf ( RI17530f50_614 , n1951 );
buf ( RI173f2950_1573 , n1817 );
buf ( RI173a9c60_1928 , n1816 );
buf ( RI174c1a70_808 , n1818 );
buf ( RI19aae980_2464 , n1815 );
buf ( RI1748ef80_1039 , n1814 );
buf ( RI173f2c98_1572 , n1846 );
buf ( RI19a97028_2633 , n1947 );
buf ( RI17476c50_1157 , n1946 );
buf ( RI173da968_1690 , n1949 );
buf ( RI17391c78_2045 , n1948 );
buf ( RI17452440_1335 , n1950 );
buf ( RI19ac6ff8_2277 , n1872 );
buf ( RI174c43b0_800 , n1871 );
buf ( RI173da620_1691 , n1972 );
buf ( RI17391930_2046 , n1971 );
buf ( RI174520f8_1336 , n1973 );
buf ( RI19ac8e70_2263 , n1970 );
buf ( RI174c3960_802 , n1969 );
buf ( RI19a99440_2617 , n1968 );
buf ( RI17476908_1158 , n1967 );
buf ( RI17405dc0_1479 , n1965 );
buf ( RI173bd0d0_1834 , n1964 );
buf ( RI17333b50_2189 , n1963 );
buf ( RI17408ef8_1464 , n1966 );
buf ( RI19ab6900_2405 , n1962 );
buf ( RI174a20a8_946 , n1961 );
buf ( RI19acc818_2235 , n1953 );
buf ( RI175153e0_700 , n1952 );
buf ( RI17397ee8_2015 , n1958 );
buf ( RI173e0bd8_1660 , n1959 );
buf ( RI174589f8_1304 , n1960 );
buf ( RI19ac3b00_2301 , n1957 );
buf ( RI174cd938_771 , n1956 );
buf ( RI19a93950_2657 , n1955 );
buf ( RI1747d208_1126 , n1954 );
buf ( RI17410860_1427 , n1806 );
buf ( RI17401f68_1498 , n1811 );
buf ( RI173b9278_1853 , n1810 );
buf ( RI175323f0_610 , n1809 );
buf ( RI1749e250_965 , n1807 );
buf ( RI19ab8f70_2388 , n1808 );
buf ( RI173d9270_1697 , n1813 );
buf ( RI173a1c68_1967 , n1812 );
buf ( RI173f81e8_1546 , n1837 );
buf ( RI173af4f8_1901 , n1836 );
buf ( RI19aaad80_2489 , n1835 );
buf ( RI17494818_1012 , n1834 );
buf ( RI173cca30_1758 , n1841 );
buf ( RI173434b0_2113 , n1840 );
buf ( RI17415a68_1402 , n1842 );
buf ( RI19a8d668_2701 , n1839 );
buf ( RI17469078_1224 , n1838 );
buf ( RI173d5aa8_1714 , n1823 );
buf ( RI19aca748_2252 , n1822 );
buf ( RI174bbda0_826 , n1821 );
buf ( RI19a9af70_2605 , n1820 );
buf ( RI17471d90_1181 , n1819 );
buf ( RI173f2fe0_1571 , n1827 );
buf ( RI173aa2f0_1926 , n1826 );
buf ( RI19aaeea8_2462 , n1825 );
buf ( RI1748f610_1037 , n1824 );
buf ( RI19a9d9a0_2587 , n1876 );
buf ( RI1748b470_1057 , n1875 );
buf ( RI17499d68_986 , n1855 );
buf ( RI19aabcf8_2483 , n1857 );
buf ( RI17492400_1023 , n1856 );
buf ( RI173a9fa8_1927 , n1845 );
buf ( RI174c5328_797 , n1847 );
buf ( RI19aaeb60_2463 , n1844 );
buf ( RI1748f2c8_1038 , n1843 );
buf ( RI173c74e0_1784 , n1853 );
buf ( RI1733df60_2139 , n1852 );
buf ( RI174101d0_1429 , n1854 );
buf ( RI19ac1490_2320 , n1851 );
buf ( RI174ac800_895 , n1850 );
buf ( RI19a91100_2675 , n1849 );
buf ( RI17463b28_1250 , n1848 );
buf ( RI174025f8_1496 , n1862 );
buf ( RI173b9908_1851 , n1861 );
buf ( RI17532e40_608 , n1860 );
buf ( RI19ab92b8_2387 , n1859 );
buf ( RI1749e8e0_963 , n1858 );
buf ( RI173dacb0_1689 , n1873 );
buf ( RI17452788_1334 , n1874 );
buf ( RI19a97208_2632 , n1870 );
buf ( RI17476f98_1156 , n1869 );
buf ( RI173ca2d0_1770 , n1867 );
buf ( RI17340d50_2125 , n1866 );
buf ( RI17413308_1414 , n1868 );
buf ( RI173a95d0_1930 , n1863 );
buf ( RI173c6130_1790 , n1891 );
buf ( RI1733cbb0_2145 , n1890 );
buf ( RI19a92bb8_2663 , n1887 );
buf ( RI17462778_1256 , n1886 );
buf ( RI19ac2f48_2307 , n1889 );
buf ( RI174ab450_901 , n1888 );
buf ( RI19aba398_2379 , n1885 );
buf ( RI1749c810_973 , n1884 );
buf ( RI173de130_1673 , n1898 );
buf ( RI17395440_2028 , n1897 );
buf ( RI17455c08_1318 , n1899 );
buf ( RI19ac6bc0_2279 , n1896 );
buf ( RI174c9630_784 , n1895 );
buf ( RI19a96e48_2634 , n1894 );
buf ( RI1747a760_1139 , n1893 );
buf ( RI173d01f8_1741 , n1903 );
buf ( RI17400528_1506 , n1902 );
buf ( RI173b7838_1861 , n1901 );
buf ( RI1752fab0_618 , n1900 );
buf ( RI173ef188_1590 , n1996 );
buf ( RI173a6498_1945 , n1995 );
buf ( RI1749c180_975 , n1997 );
buf ( RI173fcd60_1523 , n1993 );
buf ( RI173b3d28_1879 , n1992 );
buf ( RI173ade00_1908 , n1994 );
buf ( RI19aa90e8_2502 , n1991 );
buf ( RI17499048_990 , n1990 );
buf ( RI173cd0c0_1756 , n1985 );
buf ( RI17343b40_2111 , n1984 );
buf ( RI19a8db18_2699 , n1981 );
buf ( RI17469708_1222 , n1980 );
buf ( RI19abe9e8_2344 , n1983 );
buf ( RI174b23e0_867 , n1982 );
buf ( RI19a82970_2776 , n1989 );
buf ( RI1750d820_724 , n1988 );
buf ( RI19aa17f8_2556 , n1987 );
buf ( RI17486c40_1079 , n1986 );
buf ( RI1739c088_1995 , n1978 );
buf ( RI1745cb98_1284 , n1979 );
buf ( RI19a86318_2751 , n1977 );
buf ( RI17502e70_751 , n1976 );
buf ( RI19aa4ed0_2530 , n1975 );
buf ( RI174813a8_1106 , n1974 );
buf ( RI173df828_1666 , n2008 );
buf ( RI17396b38_2021 , n2007 );
buf ( RI19a95750_2644 , n2004 );
buf ( RI1747be58_1132 , n2003 );
buf ( RI19ac5540_2289 , n2006 );
buf ( RI174cba48_777 , n2005 );
buf ( RI173ef4d0_1589 , n2001 );
buf ( RI173a67e0_1944 , n2000 );
buf ( RI1749e598_964 , n2002 );
buf ( RI19a9dbf8_2586 , n1999 );
buf ( RI1748b7b8_1056 , n1998 );
buf ( RI173da2d8_1692 , n2013 );
buf ( RI17451db0_1337 , n2014 );
buf ( RI19ac8c18_2264 , n2012 );
buf ( RI174c3438_803 , n2011 );
buf ( RI19a991e8_2618 , n2010 );
buf ( RI174765c0_1159 , n2009 );
buf ( RI173d9c48_1694 , n2074 );
buf ( RI17451720_1339 , n2075 );
buf ( RI19ac8768_2266 , n2073 );
buf ( RI174c29e8_805 , n2072 );
buf ( RI19a98d38_2620 , n2071 );
buf ( RI17475f30_1161 , n2070 );
buf ( RI173f7180_1551 , n2042 );
buf ( RI173ae490_1906 , n2041 );
buf ( RI17334870_2185 , n2043 );
buf ( RI19aacbf8_2477 , n2038 );
buf ( RI174937b0_1017 , n2037 );
buf ( RI19ab8778_2392 , n2040 );
buf ( RI175217d0_662 , n2039 );
buf ( RI173f5dd0_1557 , n2047 );
buf ( RI17527ef0_642 , n2091 );
buf ( RI19ab0c30_2448 , n2090 );
buf ( RI1751f8e0_668 , n2089 );
buf ( RI173ef818_1588 , n2088 );
buf ( RI173a6b28_1943 , n2087 );
buf ( RI19acc9f8_2234 , n2086 );
buf ( RI17515908_699 , n2085 );
buf ( RI19a9de50_2585 , n2084 );
buf ( RI1748bb00_1055 , n2083 );
buf ( RI173f3328_1570 , n2081 );
buf ( RI173aa638_1925 , n2080 );
buf ( RI174cc498_775 , n2082 );
buf ( RI19aaf088_2461 , n2077 );
buf ( RI1748f958_1036 , n2076 );
buf ( RI19a23a38_2791 , n2079 );
buf ( RI1751b5d8_681 , n2078 );
buf ( RI173c7b70_1782 , n2069 );
buf ( RI1733e5f0_2137 , n2068 );
buf ( RI19ac1850_2318 , n2067 );
buf ( RI174ace90_893 , n2066 );
buf ( RI19a915b0_2673 , n2065 );
buf ( RI174641b8_1248 , n2064 );
buf ( RI173cbd10_1762 , n2097 );
buf ( RI17342790_2117 , n2096 );
buf ( RI17414d48_1406 , n2098 );
buf ( RI19a8f3f0_2688 , n2093 );
buf ( RI17468358_1228 , n2092 );
buf ( RI19abfd98_2333 , n2095 );
buf ( RI174b1030_873 , n2094 );
buf ( RI174022b0_1497 , n2106 );
buf ( RI17333178_2192 , n2105 );
buf ( RI17456c70_1313 , n2107 );
buf ( RI173eb9c0_1607 , n2103 );
buf ( RI17477cb8_1152 , n2104 );
buf ( RI19a9ff20_2569 , n2100 );
buf ( RI17487ca8_1074 , n2099 );
buf ( RI19aceac8_2220 , n2102 );
buf ( RI1750f1e8_719 , n2101 );
buf ( RI1740c378_1448 , n2028 );
buf ( RI173cda98_1753 , n2029 );
buf ( RI19ab11d0_2445 , n2026 );
buf ( RI174a89a8_914 , n2025 );
buf ( RI1733a108_2158 , n2027 );
buf ( RI173a6150_1946 , n2024 );
buf ( RI19acc3e0_2237 , n2023 );
buf ( RI19a9d658_2588 , n2022 );
buf ( RI1748b128_1058 , n2021 );
buf ( RI173f0bc8_1582 , n2019 );
buf ( RI174ac170_897 , n2020 );
buf ( RI19a86de0_2746 , n2018 );
buf ( RI175177f8_693 , n2017 );
buf ( RI19aafcb8_2455 , n2016 );
buf ( RI1748ceb0_1049 , n2015 );
buf ( RI19a85760_2756 , n2036 );
buf ( RI17500f80_757 , n2035 );
buf ( RI17407b48_1470 , n2046 );
buf ( RI19ab5640_2413 , n2045 );
buf ( RI174a3e30_937 , n2044 );
buf ( RI173bd418_1833 , n2033 );
buf ( RI17333e98_2188 , n2032 );
buf ( RI1740b310_1453 , n2034 );
buf ( RI174a23f0_945 , n2030 );
buf ( RI19ab6ae0_2404 , n2031 );
buf ( RI19a8a530_2722 , n2050 );
buf ( RI1746be68_1210 , n2049 );
buf ( RI19abc198_2367 , n2052 );
buf ( RI174b4b40_855 , n2051 );
buf ( RI173462a0_2099 , n2053 );
buf ( RI17447658_1388 , n2054 );
buf ( RI173de478_1672 , n2048 );
buf ( RI173ed0b8_1600 , n2058 );
buf ( RI173a43c8_1955 , n2057 );
buf ( RI19a9eaf8_2579 , n2056 );
buf ( RI174893a0_1067 , n2055 );
buf ( RI173c7828_1783 , n2062 );
buf ( RI1733e2a8_2138 , n2061 );
buf ( RI17410518_1428 , n2063 );
buf ( RI19a91358_2674 , n2060 );
buf ( RI17463e70_1249 , n2059 );
buf ( RI1739c718_1993 , n2121 );
buf ( RI1745d228_1282 , n2122 );
buf ( RI19aa53f8_2528 , n2118 );
buf ( RI17481a38_1104 , n2117 );
buf ( RI19a86750_2749 , n2120 );
buf ( RI175038c0_749 , n2119 );
buf ( RI19ac46b8_2296 , n2124 );
buf ( RI174c9b58_783 , n2123 );
buf ( RI19a94b98_2649 , n2126 );
buf ( RI1747b480_1135 , n2125 );
buf ( RI17395788_2027 , n2138 );
buf ( RI17455f50_1317 , n2139 );
buf ( RI19a94490_2652 , n2137 );
buf ( RI1747aaa8_1138 , n2136 );
buf ( RI1748e5a8_1042 , n2130 );
buf ( RI173c1900_1812 , n2116 );
buf ( RI17338380_2167 , n2129 );
buf ( RI174a6c20_923 , n2127 );
buf ( RI19ab2670_2436 , n2128 );
buf ( RI173dee50_1669 , n2134 );
buf ( RI17396160_2024 , n2133 );
buf ( RI17456928_1314 , n2135 );
buf ( RI19ac4dc0_2293 , n2132 );
buf ( RI174caad0_780 , n2131 );
buf ( RI1739acd8_2001 , n2142 );
buf ( RI173e39c8_1646 , n2143 );
buf ( RI1745b7e8_1290 , n2115 );
buf ( RI19aa44f8_2535 , n2141 );
buf ( RI1747fff8_1112 , n2140 );
buf ( RI173b8558_1857 , n2146 );
buf ( RI17401248_1502 , n2147 );
buf ( RI1749d530_969 , n2144 );
buf ( RI19ab8430_2393 , n2145 );
buf ( RI19a860c0_2752 , n2151 );
buf ( RI17502948_752 , n2150 );
buf ( RI19aa4cf0_2531 , n2149 );
buf ( RI17481060_1107 , n2148 );
buf ( RI173e4d78_1640 , n2153 );
buf ( RI1739bd40_1996 , n2152 );
buf ( RI1745c850_1285 , n2154 );
buf ( RI173d6138_1712 , n2113 );
buf ( RI1738d448_2067 , n2112 );
buf ( RI1744dc10_1357 , n2114 );
buf ( RI19a9b678_2602 , n2109 );
buf ( RI17472420_1179 , n2108 );
buf ( RI19acabf8_2250 , n2111 );
buf ( RI174bc7f0_824 , n2110 );
buf ( RI173ed400_1599 , n2157 );
buf ( RI17489d78_1064 , n2158 );
buf ( RI19acd808_2228 , n2156 );
buf ( RI17511b28_711 , n2155 );
buf ( RI19a952a0_2646 , n2160 );
buf ( RI1747b7c8_1134 , n2159 );
buf ( RI174a51e0_931 , n2164 );
buf ( RI1740a938_1456 , n2163 );
buf ( RI173c1c48_1811 , n2162 );
buf ( RI173386c8_2166 , n2161 );
buf ( RI17359008_2091 , n2165 );
buf ( RI173fc6d0_1525 , n2169 );
buf ( RI173b3698_1881 , n2168 );
buf ( RI19a91c40_2670 , n2167 );
buf ( RI175298b8_637 , n2166 );
buf ( RI173e5de0_1635 , n2179 );
buf ( RI1739cda8_1991 , n2178 );
buf ( RI1745d8b8_1280 , n2180 );
buf ( RI19a843b0_2764 , n2177 );
buf ( RI17506188_747 , n2176 );
buf ( RI173d15c0_1735 , n2175 );
buf ( RI173fca18_1524 , n2173 );
buf ( RI173b39e0_1880 , n2172 );
buf ( RI173ab9e8_1919 , n2174 );
buf ( RI19aa8da0_2504 , n2171 );
buf ( RI17498d00_991 , n2170 );
buf ( RI19a8b700_2715 , n2182 );
buf ( RI1746d8a8_1202 , n2181 );
buf ( RI173ea610_1613 , n2188 );
buf ( RI173a1920_1968 , n2187 );
buf ( RI1746c4f8_1208 , n2189 );
buf ( RI19a82790_2777 , n2184 );
buf ( RI1750d2f8_725 , n2183 );
buf ( RI19aa1618_2557 , n2186 );
buf ( RI174868f8_1080 , n2185 );
buf ( RI17449098_1380 , n2190 );
buf ( RI1754a6a8_69 , n2194 );
buf ( RI1754a720_68 , n2195 );
buf ( RI1754a630_70 , n2193 );
buf ( RI1754bad0_26 , n2191 );
buf ( RI1754a5b8_71 , n2192 );
buf ( RI17538c00_591 , n2196 );
buf ( RI19a25298_2780 , n2197 );
buf ( RI1754b788_33 , n2198 );
buf ( RI1754b878_31 , n2199 );
buf ( RI1754c430_6 , n2200 );
buf ( RI17536d88_596 , n2201 );
buf ( RI1754b800_32 , n2202 );
buf ( RI1754b530_38 , n2203 );
buf ( RI19a822e0_2779 , n2204 );
buf ( RI19ad0700_2208 , n2205 );
buf ( RI1754bcb0_22 , n2206 );
buf ( RI19a24ed8_2782 , n2207 );
buf ( RI19a250b8_2781 , n2208 );
buf ( RI1754be18_19 , n2209 );
buf ( RI1754b350_42 , n2210 );
buf ( RI1754c250_10 , n2211 );
buf ( RI1754b1e8_45 , n2212 );
buf ( RI19a24320_2787 , n2213 );
buf ( RI19a24578_2786 , n2214 );
buf ( RI1754b5a8_37 , n2215 );
buf ( RI19ad21b8_2198 , n2216 );
buf ( RI1754c160_12 , n2217 );
buf ( RI1754a900_64 , n2218 );
buf ( RI19a24c80_2783 , n2219 );
buf ( RI1754bf08_17 , n2220 );
buf ( RI1754ac48_57 , n2221 );
buf ( RI1754bf80_16 , n2222 );
buf ( RI1754bc38_23 , n2223 );
buf ( RI19a240c8_2788 , n2224 );
buf ( RI1754c070_14 , n2225 );
buf ( RI1754b3c8_41 , n2226 );
buf ( RI1754af18_51 , n2227 );
buf ( RI1754b080_48 , n2228 );
buf ( RI1754af90_50 , n2229 );
buf ( RI1754bda0_20 , n2230 );
buf ( RI1754aea0_52 , n2231 );
buf ( RI1754b260_44 , n2232 );
buf ( RI19ad0bb0_2206 , n2233 );
buf ( RI19a24a28_2784 , n2234 );
buf ( RI1754ae28_53 , n2235 );
buf ( RI1754a888_65 , n2236 );
buf ( RI1754bbc0_24 , n2237 );
buf ( RI19ad0e08_2205 , n2238 );
buf ( RI1754a810_66 , n2239 );
buf ( RI1754b440_40 , n2240 );
buf ( RI1754adb0_54 , n2241 );
buf ( RI1754c3b8_7 , n2242 );
buf ( RI19ad1060_2204 , n2243 );
buf ( RI1754ba58_27 , n2244 );
buf ( RI1754c340_8 , n2245 );
buf ( RI1754aa68_61 , n2246 );
buf ( RI1754ad38_55 , n2247 );
buf ( RI19ad12b8_2203 , n2248 );
buf ( RI1754be90_18 , n2249 );
buf ( RI1754c2c8_9 , n2250 );
buf ( RI1754c1d8_11 , n2251 );
buf ( RI19a247d0_2785 , n2252 );
buf ( RI1754b170_46 , n2253 );
buf ( RI1754aae0_60 , n2254 );
buf ( RI1754acc0_56 , n2255 );
buf ( RI1754a978_63 , n2256 );
buf ( RI19ad1588_2202 , n2257 );
buf ( RI1754b620_36 , n2258 );
buf ( RI1754bd28_21 , n2259 );
buf ( RI1754b9e0_28 , n2260 );
buf ( RI1754bb48_25 , n2261 );
buf ( RI1754ab58_59 , n2262 );
buf ( RI1754abd0_58 , n2263 );
buf ( RI1754b2d8_43 , n2264 );
buf ( RI1754c598_3 , n2265 );
buf ( RI19ad1858_2201 , n2266 );
buf ( RI1754b4b8_39 , n2267 );
buf ( RI1754b0f8_47 , n2268 );
buf ( RI1754c0e8_13 , n2269 );
buf ( RI1754bff8_15 , n2270 );
buf ( RI1754b698_35 , n2271 );
buf ( RI19ad1c18_2200 , n2272 );
buf ( RI1754c520_4 , n2273 );
buf ( RI1754b968_29 , n2274 );
buf ( RI19ad1ee8_2199 , n2275 );
buf ( RI1754b008_49 , n2276 );
buf ( RI1754c4a8_5 , n2277 );
buf ( RI1754b710_34 , n2278 );
buf ( RI1754a9f0_62 , n2279 );
buf ( RI1754b8f0_30 , n2280 );
buf ( RI19ad0958_2207 , n2281 );
buf ( n2282 , R_147ef_11ce6748 );
buf ( n2283 , R_5f38_10569f58 );
buf ( n2284 , R_13287_11ce6b08 );
buf ( n2285 , R_c94b_102f7608 );
buf ( n2286 , R_20a_1204ce78 );
buf ( n2287 , R_12f29_10571bb8 );
buf ( n2288 , R_13a43_13a1dec8 );
buf ( n2289 , R_1474d_1056fbd8 );
buf ( n2290 , R_14493_12657988 );
buf ( n2291 , R_11fd1_11ce17e8 );
buf ( n2292 , R_14705_1264d248 );
buf ( n2293 , R_105_f8cc2b8 );
buf ( n2294 , R_13cb9_11ce3c28 );
buf ( n2295 , R_138ee_13309fa8 );
buf ( n2296 , R_129dc_11543018 );
buf ( n2297 , R_10bcf_11ce1ba8 );
buf ( n2298 , R_13b6e_13a1e648 );
buf ( n2299 , R_14840_13a13ec8 );
buf ( n2300 , R_13482_10563838 );
buf ( n2301 , R_12d08_12650088 );
buf ( n2302 , R_10303_12b42dd8 );
buf ( n2303 , R_1437c_1056ac78 );
buf ( n2304 , R_87e9_1056cd98 );
buf ( n2305 , R_a30d_13320588 );
buf ( n2306 , R_144a2_133222e8 );
buf ( n2307 , R_1236b_13a1c8e8 );
buf ( n2308 , R_1396e_105627f8 );
buf ( n2309 , R_9ba7_10567258 );
buf ( n2310 , R_1f3_13797a68 );
buf ( n2311 , R_11c_13796528 );
buf ( n2312 , R_7a_1331e148 );
buf ( n2313 , R_117c9_1264ba88 );
buf ( n2314 , R_13b3f_1153ed38 );
buf ( n2315 , R_11abc_1264c2a8 );
buf ( n2316 , R_20d_137962a8 );
buf ( n2317 , R_207_1265a548 );
buf ( n2318 , R_14828_1207a118 );
buf ( n2319 , R_148eb_105aa7d8 );
buf ( n2320 , R_f3a4_10568bf8 );
buf ( n2321 , R_1b6_13799d68 );
buf ( n2322 , R_13429_1207f4d8 );
buf ( n2323 , R_14506_1056e878 );
buf ( n2324 , R_159_12b3d158 );
buf ( n2325 , R_108_105aaeb8 );
buf ( n2326 , R_102_13794cc8 );
buf ( n2327 , R_b1_12053638 );
buf ( n2328 , R_54_13309d28 );
buf ( n2329 , R_145d8_12b3ae58 );
buf ( n2330 , R_1278a_12083718 );
buf ( n2331 , R_13640_11cdeae8 );
buf ( n2332 , R_f706_11542578 );
buf ( n2333 , R_dc82_1153ebf8 );
buf ( n2334 , R_1491b_1265ef08 );
buf ( n2335 , R_14a05_10569738 );
buf ( n2336 , R_13fc5_102eac28 );
buf ( n2337 , R_1405a_115415d8 );
buf ( n2338 , R_136b3_126461c8 );
buf ( n2339 , R_1a0_132f9c88 );
buf ( n2340 , R_16f_1265bee8 );
buf ( n2341 , R_1480d_105a9dd8 );
buf ( n2342 , R_61_13304288 );
buf ( n2343 , R_e082_13798fa8 );
buf ( n2344 , R_10c7d_12082bd8 );
buf ( n2345 , R_14793_1379e188 );
buf ( n2346 , R_11ee1_102f4688 );
buf ( n2347 , R_128ba_12b27758 );
buf ( n2348 , R_70_120513d8 );
buf ( n2349 , R_129f0_12049bd8 );
buf ( n2350 , R_117e7_102f5588 );
buf ( n2351 , R_fee6_13309e68 );
buf ( n2352 , R_148f7_132f3ce8 );
buf ( n2353 , R_1362d_11ce39a8 );
buf ( n2354 , R_10693_126510c8 );
buf ( n2355 , R_11998_12656808 );
buf ( n2356 , R_143ec_11537df8 );
buf ( n2357 , R_138e8_1264afe8 );
buf ( n2358 , R_12650_12649b48 );
buf ( n2359 , R_137a1_105b63f8 );
buf ( n2360 , R_13afd_120772d8 );
buf ( n2361 , R_1490c_1264a7c8 );
buf ( n2362 , R_105e5_13306f88 );
buf ( n2363 , R_12e2b_132fa868 );
buf ( n2364 , R_144e7_12b38e78 );
buf ( n2365 , R_143e4_11cddf08 );
buf ( n2366 , R_1324a_1264c348 );
buf ( n2367 , R_1215a_11542ed8 );
buf ( n2368 , R_f685_11541678 );
buf ( n2369 , R_149ba_102ecb68 );
buf ( n2370 , R_135dc_12646088 );
buf ( n2371 , R_1476c_11cd7928 );
buf ( n2372 , R_146bd_11537998 );
buf ( n2373 , R_1df_12b39378 );
buf ( n2374 , R_13ee8_133069e8 );
buf ( n2375 , R_130_1265ac28 );
buf ( n2376 , R_65_12047c98 );
buf ( n2377 , R_13d75_1330d6a8 );
buf ( n2378 , R_13933_12081198 );
buf ( n2379 , R_133b5_12648388 );
buf ( n2380 , R_125a0_13311488 );
buf ( n2381 , R_8c_1379a808 );
buf ( n2382 , R_eadc_1207ead8 );
buf ( n2383 , R_134c7_126487e8 );
buf ( n2384 , R_11df5_1056e9b8 );
buf ( n2385 , R_144d5_102f8aa8 );
buf ( n2386 , R_12b2a_102eed28 );
buf ( n2387 , R_143d2_11538898 );
buf ( n2388 , R_1462c_102f8508 );
buf ( n2389 , R_13269_11543658 );
buf ( n2390 , R_f4_1331e0a8 );
buf ( n2391 , R_d7_132fde28 );
buf ( n2392 , R_238_1204ec78 );
buf ( n2393 , R_21b_1265e508 );
buf ( n2394 , R_12f3d_12b38b58 );
buf ( n2395 , R_112f1_1153c858 );
buf ( n2396 , R_f09_f8c93d8 );
buf ( n2397 , R_1487c_11cd99a8 );
buf ( n2398 , R_c08f_1207cb98 );
buf ( n2399 , R_923a_13a1ab88 );
buf ( n2400 , R_14042_102f2108 );
buf ( n2401 , R_143e8_102f3b48 );
buf ( n2402 , R_c2e7_13a19e68 );
buf ( n2403 , R_c175_12045118 );
buf ( n2404 , R_1450f_102f8b48 );
buf ( n2405 , R_12b14_12077238 );
buf ( n2406 , R_149e4_13a1c528 );
buf ( n2407 , R_12a04_11ce2968 );
buf ( n2408 , R_145ed_13a14e68 );
buf ( n2409 , R_13884_13796488 );
buf ( n2410 , R_13b0b_1330a688 );
buf ( n2411 , R_b5a4_102f4868 );
buf ( n2412 , R_14584_1056ec38 );
buf ( n2413 , R_13cee_12653148 );
buf ( n2414 , R_10bed_12080ab8 );
buf ( n2415 , R_117f0_102ef4a8 );
buf ( n2416 , R_10a2a_133048c8 );
buf ( n2417 , R_1be_137995e8 );
buf ( n2418 , R_151_12b448b8 );
buf ( n2419 , R_ef06_10563c98 );
buf ( n2420 , R_f9d4_1056b178 );
buf ( n2421 , R_e88a_13a13a68 );
buf ( n2422 , R_13c67_102f38c8 );
buf ( n2423 , R_128eb_10568dd8 );
buf ( n2424 , R_12eaf_f8c3118 );
buf ( n2425 , R_204_12039778 );
buf ( n2426 , R_14951_1265ebe8 );
buf ( n2427 , R_149c3_11ce5348 );
buf ( n2428 , R_1ad_12b28e78 );
buf ( n2429 , R_13f99_102f0da8 );
buf ( n2430 , R_162_12b25e58 );
buf ( n2431 , R_12003_11cdf628 );
buf ( n2432 , R_10b_11539478 );
buf ( n2433 , R_ff_1203c6f8 );
buf ( n2434 , R_1484f_1153ea18 );
buf ( n2435 , R_a8_12b425b8 );
buf ( n2436 , R_5d_13312068 );
buf ( n2437 , R_210_12043bd8 );
buf ( n2438 , R_13d84_102f4188 );
buf ( n2439 , R_142e1_10568658 );
buf ( n2440 , R_10f30_11cd9ae8 );
buf ( n2441 , R_1293d_12b43d78 );
buf ( n2442 , R_10b34_1056da18 );
buf ( n2443 , R_11a07_102eb4e8 );
buf ( n2444 , R_145b1_12082db8 );
buf ( n2445 , R_12c96_13a190a8 );
buf ( n2446 , R_d3b0_10565958 );
buf ( n2447 , R_13f2c_102f4b88 );
buf ( n2448 , R_fb8a_13a18608 );
buf ( n2449 , R_130d5_13319c88 );
buf ( n2450 , R_13f89_102f36e8 );
buf ( n2451 , R_146ff_13a1a4a8 );
buf ( n2452 , R_10ccb_1264f868 );
buf ( n2453 , R_124c3_1056f138 );
buf ( n2454 , R_10786_102f2568 );
buf ( n2455 , R_12a16_10568e78 );
buf ( n2456 , R_10726_102ef408 );
buf ( n2457 , R_137d3_12656da8 );
buf ( n2458 , R_13863_11cddb48 );
buf ( n2459 , R_14993_102f27e8 );
buf ( n2460 , R_bab1_1264a2c8 );
buf ( n2461 , R_1451e_10565818 );
buf ( n2462 , R_12a46_126515c8 );
buf ( n2463 , R_e7da_102f3508 );
buf ( n2464 , R_12756_13a1f0e8 );
buf ( n2465 , R_c4_13797ba8 );
buf ( n2466 , R_128da_1207ec18 );
buf ( n2467 , R_c282_12076838 );
buf ( n2468 , R_1272e_1056cbb8 );
buf ( n2469 , R_14a5f_120797b8 );
buf ( n2470 , R_14448_12663648 );
buf ( n2471 , R_c2_12048058 );
buf ( n2472 , R_1372d_11ce2aa8 );
buf ( n2473 , R_f878_1207c7d8 );
buf ( n2474 , R_13a76_13797888 );
buf ( n2475 , R_13a17_13796b68 );
buf ( n2476 , R_1cb_12044ad8 );
buf ( n2477 , R_14462_12b3f8b8 );
buf ( n2478 , R_6021_1379bd48 );
buf ( n2479 , R_144_13795128 );
buf ( n2480 , R_1383e_105671b8 );
buf ( n2481 , R_147ab_1056a6d8 );
buf ( n2482 , R_c6_1330e0a8 );
buf ( n2483 , R_249_12654368 );
buf ( n2484 , R_1305a_13796ca8 );
buf ( n2485 , R_12e4b_13307348 );
buf ( n2486 , R_14a38_137a1e28 );
buf ( n2487 , R_d1de_11cd9ea8 );
buf ( n2488 , R_138e2_11cd83c8 );
buf ( n2489 , R_13e62_1056dab8 );
buf ( n2490 , R_114a7_1331d748 );
buf ( n2491 , R_12f53_13319648 );
buf ( n2492 , R_f8a4_11543a18 );
buf ( n2493 , R_11ec3_13a157c8 );
buf ( n2494 , R_12c06_11cdac68 );
buf ( n2495 , R_12be8_12649788 );
buf ( n2496 , R_136c6_11cdc6a8 );
buf ( n2497 , R_1482e_13a1a228 );
buf ( n2498 , R_10ba7_115431f8 );
buf ( n2499 , R_89f2_11545098 );
buf ( n2500 , R_11953_1153c538 );
buf ( n2501 , R_9e64_11ce48a8 );
buf ( n2502 , R_e77d_11ce3ea8 );
buf ( n2503 , R_1091c_13a1a2c8 );
buf ( n2504 , R_114ec_12650628 );
buf ( n2505 , R_1286a_11cdcd88 );
buf ( n2506 , R_10d6d_1265db08 );
buf ( n2507 , R_1228f_1331f0e8 );
buf ( n2508 , R_1c5_126590a8 );
buf ( n2509 , R_14490_132f7d48 );
buf ( n2510 , R_1a1_1264a408 );
buf ( n2511 , R_976e_12056398 );
buf ( n2512 , R_6845_12648ec8 );
buf ( n2513 , R_16e_1379a3a8 );
buf ( n2514 , R_14a_12657528 );
buf ( n2515 , R_12718_10566fd8 );
buf ( n2516 , R_145c9_12075438 );
buf ( n2517 , R_c0_132fa5e8 );
buf ( n2518 , R_9c_12655f48 );
buf ( n2519 , R_d230_102edec8 );
buf ( n2520 , R_69_12658888 );
buf ( n2521 , R_13097_11ce5b68 );
buf ( n2522 , R_11051_1264a5e8 );
buf ( n2523 , R_145f0_11536818 );
buf ( n2524 , R_13ccd_132f9288 );
buf ( n2525 , R_e0_12661ac8 );
buf ( n2526 , R_22f_1331df68 );
buf ( n2527 , R_12a2a_11cd9f48 );
buf ( n2528 , R_10a54_11540458 );
buf ( n2529 , R_d027_13795628 );
buf ( n2530 , R_144d2_105677f8 );
buf ( n2531 , R_14638_11cd9228 );
buf ( n2532 , R_1454b_10568338 );
buf ( n2533 , R_147fe_1265bb28 );
buf ( n2534 , R_e861_12650448 );
buf ( n2535 , R_c03c_137931e8 );
buf ( n2536 , R_13574_102f97c8 );
buf ( n2537 , R_10e6d_102ec0c8 );
buf ( n2538 , R_c8_1331c348 );
buf ( n2539 , R_247_12b3bad8 );
buf ( n2540 , R_77_126636e8 );
buf ( n2541 , R_13a50_1056bb78 );
buf ( n2542 , R_129a5_11543798 );
buf ( n2543 , R_ef35_102f6d48 );
buf ( n2544 , R_1028c_137951c8 );
buf ( n2545 , R_1348b_12051838 );
buf ( n2546 , R_11f8b_11cdc428 );
buf ( n2547 , R_1452d_f8c5878 );
buf ( n2548 , R_12a3b_12650308 );
buf ( n2549 , R_13fd5_12079d58 );
buf ( n2550 , R_dd89_13302de8 );
buf ( n2551 , R_13dcc_102f7ec8 );
buf ( n2552 , R_14822_102f5768 );
buf ( n2553 , R_baf1_12084e38 );
buf ( n2554 , R_1315c_11ce75a8 );
buf ( n2555 , R_df0e_12654d68 );
buf ( n2556 , R_efea_11cdc248 );
buf ( n2557 , R_fe90_13a14a08 );
buf ( n2558 , R_1453c_102ec208 );
buf ( n2559 , R_aaa7_102edba8 );
buf ( n2560 , R_13c4e_13a1c988 );
buf ( n2561 , R_f758_13a13d88 );
buf ( n2562 , R_1485e_12b38f18 );
buf ( n2563 , R_ece9_1264c488 );
buf ( n2564 , R_14a35_12037f18 );
buf ( n2565 , R_1190c_102ecfc8 );
buf ( n2566 , R_12810_12650d08 );
buf ( n2567 , R_f016_12044df8 );
buf ( n2568 , R_1494e_13a14f08 );
buf ( n2569 , R_14344_1264eaa8 );
buf ( n2570 , R_10e_1265af48 );
buf ( n2571 , R_13f62_12075758 );
buf ( n2572 , R_fc_133201c8 );
buf ( n2573 , R_1378e_11cdd8c8 );
buf ( n2574 , R_147eb_120847f8 );
buf ( n2575 , R_13331_13308ec8 );
buf ( n2576 , R_213_12654f48 );
buf ( n2577 , R_146ae_1265dc48 );
buf ( n2578 , R_201_1153b138 );
buf ( n2579 , R_11d47_f8cc0d8 );
buf ( n2580 , R_c820_13a19328 );
buf ( n2581 , R_edbe_132fbd08 );
buf ( n2582 , R_be_132f4148 );
buf ( n2583 , R_a1_12043c78 );
buf ( n2584 , R_131b9_102f29c8 );
buf ( n2585 , R_12eb9_1153f738 );
buf ( n2586 , R_146e1_1153fb98 );
buf ( n2587 , R_1487f_13a173e8 );
buf ( n2588 , R_13fb4_11544af8 );
buf ( n2589 , R_1446b_10568798 );
buf ( n2590 , R_ef60_1264cf28 );
buf ( n2591 , R_1463b_1207bd38 );
buf ( n2592 , R_13166_1153aff8 );
buf ( n2593 , R_10a4b_10565bd8 );
buf ( n2594 , R_14599_12080c98 );
buf ( n2595 , R_10b18_12080018 );
buf ( n2596 , R_7254_12055078 );
buf ( n2597 , R_db04_1207b3d8 );
buf ( n2598 , R_149f9_10570cb8 );
buf ( n2599 , R_14a4a_1265d608 );
buf ( n2600 , R_14796_1264b808 );
buf ( n2601 , R_120d3_1379f3a8 );
buf ( n2602 , R_119cb_102f2068 );
buf ( n2603 , R_12acb_10565458 );
buf ( n2604 , R_145b4_12083358 );
buf ( n2605 , R_11ae9_12651528 );
buf ( n2606 , R_13af6_f8ce6f8 );
buf ( n2607 , R_13451_102f0128 );
buf ( n2608 , R_ef8c_1204e098 );
buf ( n2609 , R_ca_12b3e058 );
buf ( n2610 , R_245_f8c5ff8 );
buf ( n2611 , R_af_12b2a8b8 );
buf ( n2612 , R_10e57_11544eb8 );
buf ( n2613 , R_b243_f8c5698 );
buf ( n2614 , R_13633_13a13248 );
buf ( n2615 , R_11c97_10562078 );
buf ( n2616 , R_13838_102f5e48 );
buf ( n2617 , R_efb7_13a1bc68 );
buf ( n2618 , R_d4db_10566038 );
buf ( n2619 , R_10bc8_11ce66a8 );
buf ( n2620 , R_c9c0_102eee68 );
buf ( n2621 , R_13608_10563798 );
buf ( n2622 , R_8f_12b299b8 );
buf ( n2623 , R_59_133089c8 );
buf ( n2624 , R_134f1_102ebf88 );
buf ( n2625 , R_10499_1331e828 );
buf ( n2626 , R_14424_102f8f08 );
buf ( n2627 , R_1d6_133209e8 );
buf ( n2628 , R_ebe2_13a18568 );
buf ( n2629 , R_139_12b44ef8 );
buf ( n2630 , R_97_13792c48 );
buf ( n2631 , R_144ed_105660d8 );
buf ( n2632 , R_120c8_11541d58 );
buf ( n2633 , R_11736_11cde408 );
buf ( n2634 , R_149a8_13317528 );
buf ( n2635 , R_1450c_1056eff8 );
buf ( n2636 , R_147d9_120828b8 );
buf ( n2637 , R_11ea5_1264a9a8 );
buf ( n2638 , R_11425_1207c918 );
buf ( n2639 , R_d53e_1207c2d8 );
buf ( n2640 , R_14787_12b352b8 );
buf ( n2641 , R_13cf3_10571078 );
buf ( n2642 , R_13f36_1330ebe8 );
buf ( n2643 , R_d00d_102ee968 );
buf ( n2644 , R_a1e6_11cde368 );
buf ( n2645 , R_13f77_13a19648 );
buf ( n2646 , R_118_132f5f48 );
buf ( n2647 , R_13688_120832b8 );
buf ( n2648 , R_1f7_105a9978 );
buf ( n2649 , R_f630_1056b858 );
buf ( n2650 , R_136a1_1153fa58 );
buf ( n2651 , R_1b7_126577a8 );
buf ( n2652 , R_158_12b27938 );
buf ( n2653 , R_ec_1330a868 );
buf ( n2654 , R_223_f8c32f8 );
buf ( n2655 , R_133bf_11543338 );
buf ( n2656 , R_f2a8_102f47c8 );
buf ( n2657 , R_e112_12076e78 );
buf ( n2658 , R_12b72_1056c6b8 );
buf ( n2659 , R_2f00_102f3d28 );
buf ( n2660 , R_14819_1331de28 );
buf ( n2661 , R_e809_13313c48 );
buf ( n2662 , R_14358_11cd8788 );
buf ( n2663 , R_1473e_11543b58 );
buf ( n2664 , R_139c7_102ed1a8 );
buf ( n2665 , R_13d65_12036a78 );
buf ( n2666 , R_12c10_102ea548 );
buf ( n2667 , R_13870_11ce5e88 );
buf ( n2668 , R_dede_13a16448 );
buf ( n2669 , R_12c49_12b27438 );
buf ( n2670 , R_1192b_12645e08 );
buf ( n2671 , R_bd66_126533c8 );
buf ( n2672 , R_13fa2_1379f6c8 );
buf ( n2673 , R_13407_1056df18 );
buf ( n2674 , R_118b0_1204acb8 );
buf ( n2675 , R_13c3e_126496e8 );
buf ( n2676 , R_1438a_11cda268 );
buf ( n2677 , R_11e51_102fa268 );
buf ( n2678 , R_102b9_132f6588 );
buf ( n2679 , R_d9_1330dec8 );
buf ( n2680 , R_bc_13799c28 );
buf ( n2681 , R_236_13795f88 );
buf ( n2682 , R_ffee_1264d568 );
buf ( n2683 , R_10ea9_102f8788 );
buf ( n2684 , R_14852_13a154a8 );
buf ( n2685 , R_e696_11cdce28 );
buf ( n2686 , R_1ae_1203c3d8 );
buf ( n2687 , R_1457e_133027e8 );
buf ( n2688 , R_161_12656c68 );
buf ( n2689 , R_127_12b3cc58 );
buf ( n2690 , R_ea26_1265a4a8 );
buf ( n2691 , R_1e8_11539298 );
buf ( n2692 , R_139e4_102f59e8 );
buf ( n2693 , R_1477b_1204f218 );
buf ( n2694 , R_1459c_12056a78 );
buf ( n2695 , R_1336e_11545138 );
buf ( n2696 , R_108cd_102f7ce8 );
buf ( n2697 , R_13b4f_13305c28 );
buf ( n2698 , R_1a2_12b423d8 );
buf ( n2699 , R_16d_12664c28 );
buf ( n2700 , R_14656_11ce6ce8 );
buf ( n2701 , R_827e_1207e998 );
buf ( n2702 , R_11ab0_1204a358 );
buf ( n2703 , R_144ab_12b39af8 );
buf ( n2704 , R_144c3_12080338 );
buf ( n2705 , R_12794_102f5b28 );
buf ( n2706 , R_13149_102f7888 );
buf ( n2707 , R_144e4_12b28838 );
buf ( n2708 , R_13e_12660da8 );
buf ( n2709 , R_123_1330d888 );
buf ( n2710 , R_e7_137956c8 );
buf ( n2711 , R_cc_12038918 );
buf ( n2712 , R_137c7_102f79c8 );
buf ( n2713 , R_243_13796d48 );
buf ( n2714 , R_13795_13795588 );
buf ( n2715 , R_228_10570c18 );
buf ( n2716 , R_13f01_1056e2d8 );
buf ( n2717 , R_13d8e_11cd77e8 );
buf ( n2718 , R_1ec_12039ef8 );
buf ( n2719 , R_f175_13a17ca8 );
buf ( n2720 , R_1d1_126540e8 );
buf ( n2721 , R_14409_12b434b8 );
buf ( n2722 , R_138b2_102f06c8 );
buf ( n2723 , R_14653_1207e0d8 );
buf ( n2724 , R_13044_102f7a68 );
buf ( n2725 , R_13133_13a1ae08 );
buf ( n2726 , R_10b8f_1265ad68 );
buf ( n2727 , R_12e35_12b3b858 );
buf ( n2728 , R_12df0_12050bb8 );
buf ( n2729 , R_fc88_1207be78 );
buf ( n2730 , R_13804_102ef548 );
buf ( n2731 , R_13b68_137a1ba8 );
buf ( n2732 , R_134_13312b68 );
buf ( n2733 , R_14990_1331ae08 );
buf ( n2734 , R_1db_12043db8 );
buf ( n2735 , R_ccdc_102f6488 );
buf ( n2736 , R_1494b_11ce61a8 );
buf ( n2737 , R_12c39_10562ed8 );
buf ( n2738 , R_131c2_11ce4b28 );
buf ( n2739 , R_12d97_126626a8 );
buf ( n2740 , R_12d59_12b26b78 );
buf ( n2741 , R_1352d_13315188 );
buf ( n2742 , R_12c4f_13321d48 );
buf ( n2743 , R_1343e_10562d98 );
buf ( n2744 , R_1345b_102fa088 );
buf ( n2745 , R_1167d_115410d8 );
buf ( n2746 , R_14008_1264dec8 );
buf ( n2747 , R_11bc8_11544e18 );
buf ( n2748 , R_13c9a_1207e178 );
buf ( n2749 , R_148be_12b27f78 );
buf ( n2750 , R_14360_105ad078 );
buf ( n2751 , R_13aa3_12078138 );
buf ( n2752 , R_116da_13a1a7c8 );
buf ( n2753 , R_14732_102f5448 );
buf ( n2754 , R_cec6_132f3608 );
buf ( n2755 , R_133dc_13a1ea08 );
buf ( n2756 , R_14942_f8c5058 );
buf ( n2757 , R_13a0f_10563018 );
buf ( n2758 , R_bd10_f8ce978 );
buf ( n2759 , R_12da1_12647528 );
buf ( n2760 , R_12af5_12052418 );
buf ( n2761 , R_13cf9_13a1c0c8 );
buf ( n2762 , R_13658_12646628 );
buf ( n2763 , R_149bd_1204adf8 );
buf ( n2764 , R_13233_11cde908 );
buf ( n2765 , R_12585_1207a898 );
buf ( n2766 , R_118e9_10564a58 );
buf ( n2767 , R_1359a_13a18928 );
buf ( n2768 , R_12451_13a1d568 );
buf ( n2769 , R_dcbb_1265bf88 );
buf ( n2770 , R_f424_13a1b948 );
buf ( n2771 , R_1226a_11cdef48 );
buf ( n2772 , R_14641_13a12d48 );
buf ( n2773 , R_1257c_11ce4448 );
buf ( n2774 , R_e309_120806f8 );
buf ( n2775 , R_11ccc_13314be8 );
buf ( n2776 , R_146c0_13a15908 );
buf ( n2777 , R_14843_13a196e8 );
buf ( n2778 , R_11d00_1207f9d8 );
buf ( n2779 , R_14a1d_13a14c88 );
buf ( n2780 , R_13d54_11ce00c8 );
buf ( n2781 , R_135b5_132fdd88 );
buf ( n2782 , R_d40b_10569058 );
buf ( n2783 , R_145f9_102ee148 );
buf ( n2784 , R_14882_1056d838 );
buf ( n2785 , R_101a4_f8c2ad8 );
buf ( n2786 , R_13abf_13a15188 );
buf ( n2787 , R_eab3_126509e8 );
buf ( n2788 , R_8296_13322608 );
buf ( n2789 , R_6d_12036618 );
buf ( n2790 , R_50_12b3c118 );
buf ( n2791 , R_11b19_102ee508 );
buf ( n2792 , R_de1d_13a193c8 );
buf ( n2793 , R_14477_11cdcc48 );
buf ( n2794 , R_1195d_12038198 );
buf ( n2795 , R_14527_102eb6c8 );
buf ( n2796 , R_be8c_126504e8 );
buf ( n2797 , R_11e87_12b3c398 );
buf ( n2798 , R_14a02_13309aa8 );
buf ( n2799 , R_12b_1203e6d8 );
buf ( n2800 , R_f1_13799ea8 );
buf ( n2801 , R_21e_126608a8 );
buf ( n2802 , R_1e4_12b28338 );
buf ( n2803 , R_115ff_13304148 );
buf ( n2804 , R_10d8e_1264cfc8 );
buf ( n2805 , R_11500_12083c18 );
buf ( n2806 , R_c4bc_137945e8 );
buf ( n2807 , R_1465c_10568f18 );
buf ( n2808 , R_133e6_11cd9048 );
buf ( n2809 , R_7c4f_11ce4a88 );
buf ( n2810 , R_11f78_12b2c118 );
buf ( n2811 , R_1013a_132f59a8 );
buf ( n2812 , R_149e1_105b62b8 );
buf ( n2813 , R_150_1330cac8 );
buf ( n2814 , R_111_12b3e238 );
buf ( n2815 , R_f9_1204ba78 );
buf ( n2816 , R_ba_1331bc68 );
buf ( n2817 , R_4b_1264c028 );
buf ( n2818 , R_216_1204a038 );
buf ( n2819 , R_13733_f8d0098 );
buf ( n2820 , R_1fe_120539f8 );
buf ( n2821 , R_146de_12648748 );
buf ( n2822 , R_1bf_1265cd48 );
buf ( n2823 , R_74_1331da68 );
buf ( n2824 , R_f5c3_1264d108 );
buf ( n2825 , R_f1f7_120367f8 );
buf ( n2826 , R_e338_13301ac8 );
buf ( n2827 , R_1486d_1056e558 );
buf ( n2828 , R_13e2d_12047fb8 );
buf ( n2829 , R_12344_137a0de8 );
buf ( n2830 , R_14729_10570178 );
buf ( n2831 , R_13364_105717f8 );
buf ( n2832 , R_11160_1153e298 );
buf ( n2833 , R_10a01_11cde228 );
buf ( n2834 , R_13c6f_12041658 );
buf ( n2835 , R_148c4_10568978 );
buf ( n2836 , R_11c81_132f7348 );
buf ( n2837 , R_10ec5_11cdb028 );
buf ( n2838 , R_14441_12659008 );
buf ( n2839 , R_cbab_105a9a18 );
buf ( n2840 , R_1238a_126482e8 );
buf ( n2841 , R_a6_12660448 );
buf ( n2842 , R_12b36_11ce6428 );
buf ( n2843 , R_dc46_10566498 );
buf ( n2844 , R_11f_137936e8 );
buf ( n2845 , R_ce_12055fd8 );
buf ( n2846 , R_241_132fd748 );
buf ( n2847 , R_147f8_1207ccd8 );
buf ( n2848 , R_1f0_13798a08 );
buf ( n2849 , R_1467d_1056bcb8 );
buf ( n2850 , R_14668_11546178 );
buf ( n2851 , R_132cc_1153edd8 );
buf ( n2852 , R_136ba_11ce37c8 );
buf ( n2853 , R_12c23_102f1d48 );
buf ( n2854 , R_106be_1264edc8 );
buf ( n2855 , R_11bde_10564878 );
buf ( n2856 , R_11a1a_11cd9a48 );
buf ( n2857 , R_9548_11ce6ba8 );
buf ( n2858 , R_f451_11542438 );
buf ( n2859 , R_119b7_105663f8 );
buf ( n2860 , R_142e5_102f2388 );
buf ( n2861 , R_147e4_13a19dc8 );
buf ( n2862 , R_d862_12661348 );
buf ( n2863 , R_d940_13a19d28 );
buf ( n2864 , R_eb8c_13a19288 );
buf ( n2865 , R_1175e_11cda088 );
buf ( n2866 , R_146f9_11ce4768 );
buf ( n2867 , R_14551_102eae08 );
buf ( n2868 , R_14578_12b3a6d8 );
buf ( n2869 , R_1467a_13a13568 );
buf ( n2870 , R_1130e_1056bfd8 );
buf ( n2871 , R_1493f_1056d3d8 );
buf ( n2872 , R_14948_102f76a8 );
buf ( n2873 , R_10230_1153d1b8 );
buf ( n2874 , R_f4d1_13a17848 );
buf ( n2875 , R_14772_11cda8a8 );
buf ( n2876 , R_1466e_1203e138 );
buf ( n2877 , R_14999_120382d8 );
buf ( n2878 , R_9d72_102f18e8 );
buf ( n2879 , R_eeaf_10566f38 );
buf ( n2880 , R_13083_12b3ff98 );
buf ( n2881 , R_e288_11541fd8 );
buf ( n2882 , R_13969_102ea408 );
buf ( n2883 , R_13825_1264d928 );
buf ( n2884 , R_134a8_13a13c48 );
buf ( n2885 , R_fcde_115390b8 );
buf ( n2886 , R_14566_102f6988 );
buf ( n2887 , R_f5eb_11544558 );
buf ( n2888 , R_12318_102ec348 );
buf ( n2889 , R_d2c9_11cd9408 );
buf ( n2890 , R_16c_132f7ca8 );
buf ( n2891 , R_d894_1056f778 );
buf ( n2892 , R_12323_102ec8e8 );
buf ( n2893 , R_1a3_13303108 );
buf ( n2894 , R_118ba_13307ac8 );
buf ( n2895 , R_12704_10562938 );
buf ( n2896 , R_148c7_1264d888 );
buf ( n2897 , R_148bb_12661d48 );
buf ( n2898 , R_1221a_13a1d248 );
buf ( n2899 , R_135b0_12651348 );
buf ( n2900 , R_1470e_10562898 );
buf ( n2901 , R_efa_1207d1d8 );
buf ( n2902 , R_ce1e_102f95e8 );
buf ( n2903 , R_126e3_105b5c78 );
buf ( n2904 , R_14026_102ecd48 );
buf ( n2905 , R_11e36_102ed608 );
buf ( n2906 , R_11515_12039318 );
buf ( n2907 , R_108e3_1056dd38 );
buf ( n2908 , R_128f4_1207aa78 );
buf ( n2909 , R_147ae_1207ce18 );
buf ( n2910 , R_12235_12650e48 );
buf ( n2911 , R_12183_12052eb8 );
buf ( n2912 , R_14647_102f04e8 );
buf ( n2913 , R_13aef_11cdd968 );
buf ( n2914 , R_1249f_102f9368 );
buf ( n2915 , R_f34d_13a18ec8 );
buf ( n2916 , R_12c3f_f8cfd78 );
buf ( n2917 , R_13d5d_1153d4d8 );
buf ( n2918 , R_12126_102ef228 );
buf ( n2919 , R_ad_12b3b358 );
buf ( n2920 , R_92_13312d48 );
buf ( n2921 , R_113db_f8cb4f8 );
buf ( n2922 , R_10d98_f8c6318 );
buf ( n2923 , R_1481f_1264dce8 );
buf ( n2924 , R_ad98_102f3aa8 );
buf ( n2925 , R_55_132f50e8 );
buf ( n2926 , R_102d5_f8ced38 );
buf ( n2927 , R_144ae_11545ef8 );
buf ( n2928 , R_a3e0_12655308 );
buf ( n2929 , R_5dbf_13a15f48 );
buf ( n2930 , R_e2_1203f858 );
buf ( n2931 , R_22d_1379de68 );
buf ( n2932 , R_135c4_105b5bd8 );
buf ( n2933 , R_13cff_13a16308 );
buf ( n2934 , R_12692_102eb8a8 );
buf ( n2935 , R_13375_13794a48 );
buf ( n2936 , R_12f6a_10562438 );
buf ( n2937 , R_128c4_102ea5e8 );
buf ( n2938 , R_122f0_12650f88 );
buf ( n2939 , R_14855_12056f78 );
buf ( n2940 , R_14885_13795a88 );
buf ( n2941 , R_bb92_11ce0ca8 );
buf ( n2942 , R_8b04_1265cf28 );
buf ( n2943 , R_e71c_115426b8 );
buf ( n2944 , R_14a23_120545d8 );
buf ( n2945 , R_149_1330f408 );
buf ( n2946 , R_b8_13305048 );
buf ( n2947 , R_1c6_1379cce8 );
buf ( n2948 , R_e13d_102eb448 );
buf ( n2949 , R_14617_11ce2f08 );
buf ( n2950 , R_13557_11545778 );
buf ( n2951 , R_148cd_12082c78 );
buf ( n2952 , R_11768_1264ffe8 );
buf ( n2953 , R_12503_11cdd008 );
buf ( n2954 , R_1239d_1330d1a8 );
buf ( n2955 , R_1448c_105662b8 );
buf ( n2956 , R_160_f8c0d78 );
buf ( n2957 , R_143_13795e48 );
buf ( n2958 , R_1252c_102f1208 );
buf ( n2959 , R_1cc_f8cc858 );
buf ( n2960 , R_149de_11cde7c8 );
buf ( n2961 , R_1af_12b40678 );
buf ( n2962 , R_a28f_11ce5708 );
buf ( n2963 , R_f7ae_11ce57a8 );
buf ( n2964 , R_1243d_10571118 );
buf ( n2965 , R_d0df_126478e8 );
buf ( n2966 , R_1498d_1153fe18 );
buf ( n2967 , R_10350_11cda6c8 );
buf ( n2968 , R_103a6_10569878 );
buf ( n2969 , R_128b0_1056c118 );
buf ( n2970 , R_14936_10561e98 );
buf ( n2971 , R_10d1b_11cd7748 );
buf ( n2972 , R_ed92_102eea08 );
buf ( n2973 , R_145d2_11cdb208 );
buf ( n2974 , R_109f6_1153ca38 );
buf ( n2975 , R_cc46_1207b298 );
buf ( n2976 , R_11006_126501c8 );
buf ( n2977 , R_188_1265c348 );
buf ( n2978 , R_187_12b25d18 );
buf ( n2979 , R_12f_1379dbe8 );
buf ( n2980 , R_db_12663f08 );
buf ( n2981 , R_84_12652ce8 );
buf ( n2982 , R_81_12042a58 );
buf ( n2983 , R_234_12b43af8 );
buf ( n2984 , R_1e0_133037e8 );
buf ( n2985 , R_13ed7_1207ad98 );
buf ( n2986 , R_189_f8c6458 );
buf ( n2987 , R_186_126553a8 );
buf ( n2988 , R_157_132f7a28 );
buf ( n2989 , R_d0_105aa238 );
buf ( n2990 , R_23f_13307848 );
buf ( n2991 , R_11399_12b3c1b8 );
buf ( n2992 , R_1b8_11537358 );
buf ( n2993 , R_f82c_f8cdc58 );
buf ( n2994 , R_d9ca_10562bb8 );
buf ( n2995 , R_145f6_f8c3398 );
buf ( n2996 , R_1449c_11ce71e8 );
buf ( n2997 , R_13850_13a1fe08 );
buf ( n2998 , R_135e3_13306da8 );
buf ( n2999 , R_ec0b_132fa368 );
buf ( n3000 , R_147e0_13a12fc8 );
buf ( n3001 , R_13add_132ff728 );
buf ( n3002 , R_f65b_12084578 );
buf ( n3003 , R_10cb4_11cdf9e8 );
buf ( n3004 , R_18a_133173e8 );
buf ( n3005 , R_185_12042cd8 );
buf ( n3006 , R_134d0_12651028 );
buf ( n3007 , R_144f3_102f3fa8 );
buf ( n3008 , R_12dd1_f8c52d8 );
buf ( n3009 , R_135a9_10567938 );
buf ( n3010 , R_11b39_102ec988 );
buf ( n3011 , R_1386a_102ebda8 );
buf ( n3012 , R_14747_12042b98 );
buf ( n3013 , R_148d0_137a0a28 );
buf ( n3014 , R_11f4d_137986e8 );
buf ( n3015 , R_13d05_12081378 );
buf ( n3016 , R_f56e_102f2608 );
buf ( n3017 , R_62_12b26498 );
buf ( n3018 , R_10e0b_1056abd8 );
buf ( n3019 , R_ba73_1264c8e8 );
buf ( n3020 , R_14888_12653288 );
buf ( n3021 , R_fc34_1379c428 );
buf ( n3022 , R_18b_12663fa8 );
buf ( n3023 , R_184_1153acd8 );
buf ( n3024 , R_119d5_1331dc48 );
buf ( n3025 , R_122b5_13305688 );
buf ( n3026 , R_e051_12649f08 );
buf ( n3027 , R_ca0a_10567438 );
buf ( n3028 , R_10a84_115427f8 );
buf ( n3029 , R_668e_10563f18 );
buf ( n3030 , R_14539_102f7108 );
buf ( n3031 , R_c3d6_11cdb7a8 );
buf ( n3032 , R_11703_132fa728 );
buf ( n3033 , R_1472f_105708f8 );
buf ( n3034 , R_1307a_11cdc1a8 );
buf ( n3035 , R_fdae_1153d258 );
buf ( n3036 , R_13ac5_102ee3c8 );
buf ( n3037 , R_120bd_1153ff58 );
buf ( n3038 , R_13f6e_12649dc8 );
buf ( n3039 , R_1177b_1207fbb8 );
buf ( n3040 , R_f804_1379efe8 );
buf ( n3041 , R_111d5_13a17c08 );
buf ( n3042 , R_14750_13304008 );
buf ( n3043 , R_137d9_12055e98 );
buf ( n3044 , R_87_132ffa48 );
buf ( n3045 , R_7e_137949a8 );
buf ( n3046 , R_f140_1056f598 );
buf ( n3047 , R_d43f_12079678 );
buf ( n3048 , R_11900_1056f6d8 );
buf ( n3049 , R_18c_12660e48 );
buf ( n3050 , R_c969_1330f9a8 );
buf ( n3051 , R_183_126587e8 );
buf ( n3052 , R_11093_102f60c8 );
buf ( n3053 , R_f31e_120770f8 );
buf ( n3054 , R_f06_1265f728 );
buf ( n3055 , R_d5cf_102f5128 );
buf ( n3056 , R_10874_12037838 );
buf ( n3057 , R_11324_13a1f228 );
buf ( n3058 , R_13621_120823b8 );
buf ( n3059 , R_120dd_f8cdcf8 );
buf ( n3060 , R_148d3_12049a98 );
buf ( n3061 , R_13e42_12648888 );
buf ( n3062 , R_144c0_12078db8 );
buf ( n3063 , R_12978_13316d08 );
buf ( n3064 , R_11b5e_13a1b088 );
buf ( n3065 , R_13025_13a1ef08 );
buf ( n3066 , R_e615_12084bb8 );
buf ( n3067 , R_149b7_102ea4a8 );
buf ( n3068 , R_1497e_1207ef38 );
buf ( n3069 , R_11fee_12b2a3b8 );
buf ( n3070 , R_11b_12b43198 );
buf ( n3071 , R_5e_126647c8 );
buf ( n3072 , R_1f4_1265d108 );
buf ( n3073 , R_1445f_13792888 );
buf ( n3074 , R_13981_13798aa8 );
buf ( n3075 , R_14569_11cdbfc8 );
buf ( n3076 , R_114_12b3e4b8 );
buf ( n3077 , R_f6_12664188 );
buf ( n3078 , R_9f_12054d58 );
buf ( n3079 , R_66_13308068 );
buf ( n3080 , R_219_1203c338 );
buf ( n3081 , R_132a5_12654868 );
buf ( n3082 , R_f9aa_11cdd5a8 );
buf ( n3083 , R_1fb_126610c8 );
buf ( n3084 , R_1a4_13798648 );
buf ( n3085 , R_16b_1331a2c8 );
buf ( n3086 , R_9a_12658568 );
buf ( n3087 , R_13c54_102f6e88 );
buf ( n3088 , R_14933_1207e5d8 );
buf ( n3089 , R_a6b7_1264b588 );
buf ( n3090 , R_10fad_13a15548 );
buf ( n3091 , R_18d_13321a28 );
buf ( n3092 , R_182_13315cc8 );
buf ( n3093 , R_14a58_102f65c8 );
buf ( n3094 , R_c8f6_132f4a08 );
buf ( n3095 , R_1458d_13a17ac8 );
buf ( n3096 , R_126d9_11545598 );
buf ( n3097 , R_10942_102f85a8 );
buf ( n3098 , R_14a32_12654ea8 );
buf ( n3099 , R_b7bc_12b28798 );
buf ( n3100 , R_1389f_11cda3a8 );
buf ( n3101 , R_14602_102ed7e8 );
buf ( n3102 , R_100bf_1330b9e8 );
buf ( n3103 , R_112eb_115386b8 );
buf ( n3104 , R_146d5_105b59f8 );
buf ( n3105 , R_1206a_1207c878 );
buf ( n3106 , R_e2de_1264ce88 );
buf ( n3107 , R_13b3a_11cddaa8 );
buf ( n3108 , R_13739_10563bf8 );
buf ( n3109 , R_148d6_11cd86e8 );
buf ( n3110 , R_1319d_11544918 );
buf ( n3111 , R_12f7f_12077eb8 );
buf ( n3112 , R_1242c_f8cda78 );
buf ( n3113 , R_14483_12054fd8 );
buf ( n3114 , R_14456_102ea728 );
buf ( n3115 , R_6b42_120790d8 );
buf ( n3116 , R_1186d_f8cbb38 );
buf ( n3117 , R_147d3_12648e28 );
buf ( n3118 , R_11add_1056c4d8 );
buf ( n3119 , R_13c18_1264df68 );
buf ( n3120 , R_13e19_132f7c08 );
buf ( n3121 , R_b6_1265e148 );
buf ( n3122 , R_13bb8_1265edc8 );
buf ( n3123 , R_146a8_12050118 );
buf ( n3124 , R_18e_12043ef8 );
buf ( n3125 , R_181_12647a28 );
buf ( n3126 , R_b677_12083178 );
buf ( n3127 , R_1176f_1379f8a8 );
buf ( n3128 , R_11d7b_102f2d88 );
buf ( n3129 , R_145bd_1207cff8 );
buf ( n3130 , R_13bae_105700d8 );
buf ( n3131 , R_10fed_1330ad68 );
buf ( n3132 , R_1479f_11cde4a8 );
buf ( n3133 , R_71_1265e8c8 );
buf ( n3134 , R_3ca5_102eebe8 );
buf ( n3135 , R_14769_1056b718 );
buf ( n3136 , R_139ba_11ce35e8 );
buf ( n3137 , R_ccf5_13a128e8 );
buf ( n3138 , R_13964_1207def8 );
buf ( n3139 , R_13920_133128e8 );
buf ( n3140 , R_13b74_11cd8dc8 );
buf ( n3141 , R_13e6d_11cd90e8 );
buf ( n3142 , R_13ae8_11545db8 );
buf ( n3143 , R_e946_13796668 );
buf ( n3144 , R_12db3_10562b18 );
buf ( n3145 , R_7b5f_1264bc68 );
buf ( n3146 , R_139f5_132fc348 );
buf ( n3147 , R_cd6e_10562a78 );
buf ( n3148 , R_13626_12077cd8 );
buf ( n3149 , R_148dc_102f3c88 );
buf ( n3150 , R_11db0_13302748 );
buf ( n3151 , R_1470b_115413f8 );
buf ( n3152 , R_fd8e_120835d8 );
buf ( n3153 , R_142aa_102f2a68 );
buf ( n3154 , R_1267b_1056b538 );
buf ( n3155 , R_10df7_1264ae08 );
buf ( n3156 , R_b753_102ebe48 );
buf ( n3157 , R_14a47_102eeb48 );
buf ( n3158 , R_12f94_1379c068 );
buf ( n3159 , R_f3d0_1264e3c8 );
buf ( n3160 , R_13cd6_10565638 );
buf ( n3161 , R_123b1_12b3e378 );
buf ( n3162 , R_144cf_f8c96f8 );
buf ( n3163 , R_13d0c_102f6168 );
buf ( n3164 , R_13c61_12081d78 );
buf ( n3165 , R_134f6_11ce6608 );
buf ( n3166 , R_112c2_12b294b8 );
buf ( n3167 , R_11922_1056c898 );
buf ( n3168 , R_11971_1207dbd8 );
buf ( n3169 , R_138_1265b308 );
buf ( n3170 , R_d2_12654c28 );
buf ( n3171 , R_23d_12656088 );
buf ( n3172 , R_8a_1379cba8 );
buf ( n3173 , R_38ad_12048418 );
buf ( n3174 , R_7b_12651de8 );
buf ( n3175 , R_13889_10564918 );
buf ( n3176 , R_13188_12079c18 );
buf ( n3177 , R_13b8c_13a15728 );
buf ( n3178 , R_947f_1056eaf8 );
buf ( n3179 , R_1d7_12649648 );
buf ( n3180 , R_149db_102f1668 );
buf ( n3181 , R_ac1d_120826d8 );
buf ( n3182 , R_13a06_105668f8 );
buf ( n3183 , R_18f_132fc988 );
buf ( n3184 , R_180_1265fea8 );
buf ( n3185 , R_10e36_11ce6d88 );
buf ( n3186 , R_136a7_12035cb8 );
buf ( n3187 , R_148df_13a1d608 );
buf ( n3188 , R_1380f_12080838 );
buf ( n3189 , R_1485b_1265a688 );
buf ( n3190 , R_14930_102f1a28 );
buf ( n3191 , R_10044_102f1c08 );
buf ( n3192 , R_d2a3_1207bbf8 );
buf ( n3193 , R_1c0_1203c0b8 );
buf ( n3194 , R_14f_12b25778 );
buf ( n3195 , R_8472_126654e8 );
buf ( n3196 , R_1483d_11ce0d48 );
buf ( n3197 , R_12b67_11cdf3a8 );
buf ( n3198 , R_11346_12655448 );
buf ( n3199 , R_13893_12084d98 );
buf ( n3200 , R_103f0_1207ecb8 );
buf ( n3201 , R_1308d_1379eea8 );
buf ( n3202 , R_f8ce_102f10c8 );
buf ( n3203 , R_13f82_11543978 );
buf ( n3204 , R_12359_133022e8 );
buf ( n3205 , R_12cd3_13a1f728 );
buf ( n3206 , R_13546_1153efb8 );
buf ( n3207 , R_143b6_115408b8 );
buf ( n3208 , R_148e5_10568518 );
buf ( n3209 , R_10a79_11545278 );
buf ( n3210 , R_1368d_102f3be8 );
buf ( n3211 , R_14002_12047518 );
buf ( n3212 , R_febc_1207caf8 );
buf ( n3213 , R_14987_10571d98 );
buf ( n3214 , R_14894_126569e8 );
buf ( n3215 , R_13e23_102f1708 );
buf ( n3216 , R_12304_10569e18 );
buf ( n3217 , R_12daa_f8cc218 );
buf ( n3218 , R_1289e_13316128 );
buf ( n3219 , R_146ea_132fd6a8 );
buf ( n3220 , R_104_12b414d8 );
buf ( n3221 , R_e9_12055a78 );
buf ( n3222 , R_226_12652568 );
buf ( n3223 , R_20b_12656bc8 );
buf ( n3224 , R_1484c_1056c078 );
buf ( n3225 , R_149fc_12077a58 );
buf ( n3226 , R_143f0_120442b8 );
buf ( n3227 , R_107_1203f538 );
buf ( n3228 , R_208_12b260d8 );
buf ( n3229 , R_1d2_1203ce78 );
buf ( n3230 , R_1442a_102f6668 );
buf ( n3231 , R_13d_1379c568 );
buf ( n3232 , R_134be_13a19148 );
buf ( n3233 , R_145cf_13304328 );
buf ( n3234 , R_12fa4_1153e0b8 );
buf ( n3235 , R_1053d_12079858 );
buf ( n3236 , R_ee_f8c86b8 );
buf ( n3237 , R_221_12652888 );
buf ( n3238 , R_13eb5_132f7ac8 );
buf ( n3239 , R_190_133178e8 );
buf ( n3240 , R_17f_115396f8 );
buf ( n3241 , R_137af_11ce6e28 );
buf ( n3242 , R_1455a_102ed748 );
buf ( n3243 , R_10db8_102f74c8 );
buf ( n3244 , R_ab_1264cde8 );
buf ( n3245 , R_1187e_12077698 );
buf ( n3246 , R_5a_126653a8 );
buf ( n3247 , R_7e57_13a1a188 );
buf ( n3248 , R_146ed_1153a238 );
buf ( n3249 , R_1b0_12b29918 );
buf ( n3250 , R_15f_1265f188 );
buf ( n3251 , R_138b8_1264a368 );
buf ( n3252 , R_13bd6_102f9188 );
buf ( n3253 , R_14a17_102f0ee8 );
buf ( n3254 , R_143a6_133121a8 );
buf ( n3255 , R_11f57_12649328 );
buf ( n3256 , R_14972_13302608 );
buf ( n3257 , R_10701_1207f1b8 );
buf ( n3258 , R_14503_1203e3b8 );
buf ( n3259 , R_a4_12b36e98 );
buf ( n3260 , R_6a_12b40178 );
buf ( n3261 , R_aeba_105624d8 );
buf ( n3262 , R_1379b_11ce6ec8 );
buf ( n3263 , R_134e2_13a1e3c8 );
buf ( n3264 , R_10973_12663008 );
buf ( n3265 , R_11c66_102f7ba8 );
buf ( n3266 , R_1325f_126468a8 );
buf ( n3267 , R_1327d_10570d58 );
buf ( n3268 , R_13417_102f3968 );
buf ( n3269 , R_101_1264f048 );
buf ( n3270 , R_95_133017a8 );
buf ( n3271 , R_20e_1265e788 );
buf ( n3272 , R_13c59_105b5638 );
buf ( n3273 , R_13ca1_12652f68 );
buf ( n3274 , R_1481c_11cdb988 );
buf ( n3275 , R_14611_11545458 );
buf ( n3276 , R_12fae_102f7388 );
buf ( n3277 , R_1469f_1207d138 );
buf ( n3278 , R_142dd_13314828 );
buf ( n3279 , R_1279d_12079fd8 );
buf ( n3280 , R_12646_1056b2b8 );
buf ( n3281 , R_11486_102ee788 );
buf ( n3282 , R_13389_1207fb18 );
buf ( n3283 , R_1492d_11ce64c8 );
buf ( n3284 , R_12d46_12648928 );
buf ( n3285 , R_145b7_12b3d5b8 );
buf ( n3286 , R_b211_12048c38 );
buf ( n3287 , R_143aa_13795c68 );
buf ( n3288 , R_1110c_11cdc928 );
buf ( n3289 , R_1a5_12b3c618 );
buf ( n3290 , R_16a_137a1248 );
buf ( n3291 , R_df67_1207b8d8 );
buf ( n3292 , R_124f6_1264f2c8 );
buf ( n3293 , R_12b54_102f2248 );
buf ( n3294 , R_d7dc_13a17de8 );
buf ( n3295 , R_1247b_11ce4808 );
buf ( n3296 , R_149ea_11540598 );
buf ( n3297 , R_10a_12b30678 );
buf ( n3298 , R_13c77_13a1cc08 );
buf ( n3299 , R_205_12653dc8 );
buf ( n3300 , R_14753_1264efa8 );
buf ( n3301 , R_191_12043d18 );
buf ( n3302 , R_17e_132f8568 );
buf ( n3303 , R_11c4b_13a15c28 );
buf ( n3304 , R_13208_11542758 );
buf ( n3305 , R_e0ad_133021a8 );
buf ( n3306 , R_11a3f_12b3e9b8 );
buf ( n3307 , R_1230e_f8cb598 );
buf ( n3308 , R_eee_1056adb8 );
buf ( n3309 , R_14444_12648108 );
buf ( n3310 , R_1dc_11538d98 );
buf ( n3311 , R_12b7a_1264f188 );
buf ( n3312 , R_133_13313888 );
buf ( n3313 , R_147b1_105b5a98 );
buf ( n3314 , R_f116_11ce1068 );
buf ( n3315 , R_13a5c_1379a268 );
buf ( n3316 , R_14340_12078458 );
buf ( n3317 , R_e522_1330ed28 );
buf ( n3318 , R_146f0_1153da78 );
buf ( n3319 , R_136f4_12649148 );
buf ( n3320 , R_119e8_1153e798 );
buf ( n3321 , R_1391b_12b277f8 );
buf ( n3322 , R_fd37_120394f8 );
buf ( n3323 , R_1461d_11539dd8 );
buf ( n3324 , R_ee50_102eb9e8 );
buf ( n3325 , R_dd_132f61c8 );
buf ( n3326 , R_232_105afa58 );
buf ( n3327 , R_4c_12652b08 );
buf ( n3328 , R_135a0_1153f0f8 );
buf ( n3329 , R_125d0_12b3f6d8 );
buf ( n3330 , R_b4_13302988 );
buf ( n3331 , R_51_13309648 );
buf ( n3332 , R_f925_12048b98 );
buf ( n3333 , R_14034_f8cf198 );
buf ( n3334 , R_123e9_f8c0eb8 );
buf ( n3335 , R_14726_1203bc58 );
buf ( n3336 , R_10894_1153ad78 );
buf ( n3337 , R_1b9_1379b7a8 );
buf ( n3338 , R_156_137927e8 );
buf ( n3339 , R_1471a_1379da08 );
buf ( n3340 , R_13d4e_11544f58 );
buf ( n3341 , R_112ae_115429d8 );
buf ( n3342 , R_dcb0_10564e18 );
buf ( n3343 , R_13ae3_12083498 );
buf ( n3344 , R_11a90_13a1ba88 );
buf ( n3345 , R_13f1a_10566998 );
buf ( n3346 , R_fdd5_1264d068 );
buf ( n3347 , R_13acb_13a17988 );
buf ( n3348 , R_ef1_13a16ee8 );
buf ( n3349 , R_145e1_12b40d58 );
buf ( n3350 , R_14915_102f7748 );
buf ( n3351 , R_ed3c_120760b8 );
buf ( n3352 , R_13cdc_11542398 );
buf ( n3353 , R_f544_102f5d08 );
buf ( n3354 , R_147e7_13793fa8 );
buf ( n3355 , R_e4_133095a8 );
buf ( n3356 , R_8d_1153d078 );
buf ( n3357 , R_78_12044178 );
buf ( n3358 , R_22b_12b3b538 );
buf ( n3359 , R_128ff_105b6178 );
buf ( n3360 , R_148ac_102f0f88 );
buf ( n3361 , R_1e9_133208a8 );
buf ( n3362 , R_192_12b44a98 );
buf ( n3363 , R_17d_12661f28 );
buf ( n3364 , R_12b83_13305e08 );
buf ( n3365 , R_fbb3_10567078 );
buf ( n3366 , R_126_12660588 );
buf ( n3367 , R_cfc6_1264a868 );
buf ( n3368 , R_1492a_13a1e1e8 );
buf ( n3369 , R_116bb_1207d6d8 );
buf ( n3370 , R_144d8_1330d9c8 );
buf ( n3371 , R_e6f2_102ecc08 );
buf ( n3372 , R_14a14_1207bdd8 );
buf ( n3373 , R_10f70_11544a58 );
buf ( n3374 , R_119fa_1207f2f8 );
buf ( n3375 , R_cef5_1265b6c8 );
buf ( n3376 , R_115b3_12082458 );
buf ( n3377 , R_211_1265c028 );
buf ( n3378 , R_146cc_11542618 );
buf ( n3379 , R_fe_120448f8 );
buf ( n3380 , R_119df_1056bad8 );
buf ( n3381 , R_13787_11ce21e8 );
buf ( n3382 , R_147dd_11ce6068 );
buf ( n3383 , R_14695_11cdf8a8 );
buf ( n3384 , R_149b1_102fa128 );
buf ( n3385 , R_110af_1379aee8 );
buf ( n3386 , R_14560_1330b3a8 );
buf ( n3387 , R_143ff_11cdca68 );
buf ( n3388 , R_d4_12654a48 );
buf ( n3389 , R_23b_13799408 );
buf ( n3390 , R_1c7_132fc0c8 );
buf ( n3391 , R_148_105aacd8 );
buf ( n3392 , R_13d6d_13a17668 );
buf ( n3393 , R_ce64_1056f9f8 );
buf ( n3394 , R_14474_13307a28 );
buf ( n3395 , R_12bde_102f62a8 );
buf ( n3396 , R_1436a_102eefa8 );
buf ( n3397 , R_14957_11540db8 );
buf ( n3398 , R_b634_11cdc068 );
buf ( n3399 , R_1460e_11ce2dc8 );
buf ( n3400 , R_f24f_11ce2fa8 );
buf ( n3401 , R_13763_105679d8 );
buf ( n3402 , R_f0b2_102f7f68 );
buf ( n3403 , R_14620_11ce6108 );
buf ( n3404 , R_131f5_12084618 );
buf ( n3405 , R_1490f_12651e88 );
buf ( n3406 , R_136cc_1264fcc8 );
buf ( n3407 , R_f227_1207a398 );
buf ( n3408 , R_13959_1153f918 );
buf ( n3409 , R_142cf_12659aa8 );
buf ( n3410 , R_f6b2_11cdfb28 );
buf ( n3411 , R_1ed_1203f5d8 );
buf ( n3412 , R_a2f6_11cdb3e8 );
buf ( n3413 , R_fc5e_13a18888 );
buf ( n3414 , R_122_12663d28 );
buf ( n3415 , R_13f67_12083b78 );
buf ( n3416 , R_13740_11cdb348 );
buf ( n3417 , R_146c9_1153fd78 );
buf ( n3418 , R_145db_13a12b68 );
buf ( n3419 , R_101ae_13a1fae8 );
buf ( n3420 , R_bb03_12b29ff8 );
buf ( n3421 , R_1101b_12045f38 );
buf ( n3422 , R_12bfd_10564b98 );
buf ( n3423 , R_121a5_1056a138 );
buf ( n3424 , R_127df_1330a728 );
buf ( n3425 , R_11617_105656d8 );
buf ( n3426 , R_13f90_12080518 );
buf ( n3427 , R_13be9_12662388 );
buf ( n3428 , R_12760_1331ab88 );
buf ( n3429 , R_126bb_10563b58 );
buf ( n3430 , R_147c6_12081cd8 );
buf ( n3431 , R_21c_12b41398 );
buf ( n3432 , R_13b33_102f0588 );
buf ( n3433 , R_1f8_132f5fe8 );
buf ( n3434 , R_11d2f_105665d8 );
buf ( n3435 , R_1227d_1265f2c8 );
buf ( n3436 , R_11a35_102f44a8 );
buf ( n3437 , R_1479c_1056c758 );
buf ( n3438 , R_116e4_12659828 );
buf ( n3439 , R_14662_1207ceb8 );
buf ( n3440 , R_14515_12079ad8 );
buf ( n3441 , R_117_12650c68 );
buf ( n3442 , R_115ca_11ce5fc8 );
buf ( n3443 , R_f3_1379bde8 );
buf ( n3444 , R_e229_102ecca8 );
buf ( n3445 , R_202_12b3f098 );
buf ( n3446 , R_1e5_1203a218 );
buf ( n3447 , R_12a_1331fea8 );
buf ( n3448 , R_10d_1330bda8 );
buf ( n3449 , R_135d6_1056fef8 );
buf ( n3450 , R_14918_13a1d888 );
buf ( n3451 , R_1452a_10564378 );
buf ( n3452 , R_14984_1056bc18 );
buf ( n3453 , R_1cd_1265c8e8 );
buf ( n3454 , R_eb34_11cda628 );
buf ( n3455 , R_125ac_11ce4308 );
buf ( n3456 , R_193_f8c7cb8 );
buf ( n3457 , R_1216d_1264d7e8 );
buf ( n3458 , R_17c_132fe648 );
buf ( n3459 , R_142_13792ce8 );
buf ( n3460 , R_cdb8_102f4f48 );
buf ( n3461 , R_144bd_11cdeb88 );
buf ( n3462 , R_131ae_1056bd58 );
buf ( n3463 , R_14909_1379f768 );
buf ( n3464 , R_14924_12b3adb8 );
buf ( n3465 , R_102a2_12b41e38 );
buf ( n3466 , R_13aa8_120525f8 );
buf ( n3467 , R_d3ca_102ef7c8 );
buf ( n3468 , R_1459f_120792b8 );
buf ( n3469 , R_120b3_12b407b8 );
buf ( n3470 , R_127a7_105683d8 );
buf ( n3471 , R_14545_1056b218 );
buf ( n3472 , R_12056_1204f178 );
buf ( n3473 , R_11f2a_10563ab8 );
buf ( n3474 , R_e021_12b26718 );
buf ( n3475 , R_f377_1056d1f8 );
buf ( n3476 , R_127ca_13a16da8 );
buf ( n3477 , R_14689_120838f8 );
buf ( n3478 , R_11be7_1207a6b8 );
buf ( n3479 , R_139a1_1264c668 );
buf ( n3480 , R_14536_12b42978 );
buf ( n3481 , R_13c2d_11cdd828 );
buf ( n3482 , R_14906_11544ff8 );
buf ( n3483 , R_11a5d_132f52c8 );
buf ( n3484 , R_ca63_1331c8e8 );
buf ( n3485 , R_14714_102f77e8 );
buf ( n3486 , R_14799_137933c8 );
buf ( n3487 , R_1390f_13a14828 );
buf ( n3488 , R_1234f_12083858 );
buf ( n3489 , R_142c6_12081738 );
buf ( n3490 , R_127ae_12b3ccf8 );
buf ( n3491 , R_13590_12079a38 );
buf ( n3492 , R_148b8_102eaa48 );
buf ( n3493 , R_5735_137a0988 );
buf ( n3494 , R_1a6_12038698 );
buf ( n3495 , R_169_1203e458 );
buf ( n3496 , R_127c1_12082638 );
buf ( n3497 , R_1288a_137a1ec8 );
buf ( n3498 , R_1488e_102f6708 );
buf ( n3499 , R_113b9_1264ea08 );
buf ( n3500 , R_1430f_11cd8fa8 );
buf ( n3501 , R_f97f_13304dc8 );
buf ( n3502 , R_104fa_120761f8 );
buf ( n3503 , R_119ae_11cdfa88 );
buf ( n3504 , R_12c78_1207ca58 );
buf ( n3505 , R_d606_11ce46c8 );
buf ( n3506 , R_146a5_102f90e8 );
buf ( n3507 , R_14900_120781d8 );
buf ( n3508 , R_1374f_13a16808 );
buf ( n3509 , R_ff3c_11ce1f68 );
buf ( n3510 , R_e834_10564238 );
buf ( n3511 , R_14a5e_105aa4b8 );
buf ( n3512 , R_13465_13316bc8 );
buf ( n3513 , R_13d25_11540b38 );
buf ( n3514 , R_56_13308248 );
buf ( n3515 , R_ef7_1153e838 );
buf ( n3516 , R_13193_102ec7a8 );
buf ( n3517 , R_132f1_13a145a8 );
buf ( n3518 , R_1291e_1056ee18 );
buf ( n3519 , R_14921_105640f8 );
buf ( n3520 , R_1371a_12083fd8 );
buf ( n3521 , R_14837_132f32e8 );
buf ( n3522 , R_13a37_12b3d338 );
buf ( n3523 , R_dad2_1379c6a8 );
buf ( n3524 , R_1495d_12b43878 );
buf ( n3525 , R_149f3_12b27c58 );
buf ( n3526 , R_107c6_1203f998 );
buf ( n3527 , R_1456c_12b437d8 );
buf ( n3528 , R_11888_13794868 );
buf ( n3529 , R_13b62_13a13428 );
buf ( n3530 , R_1360f_10563158 );
buf ( n3531 , R_1b1_12657ac8 );
buf ( n3532 , R_10844_1153e1f8 );
buf ( n3533 , R_194_1331d4c8 );
buf ( n3534 , R_17b_1265ea08 );
buf ( n3535 , R_15e_126544a8 );
buf ( n3536 , R_be25_102ec028 );
buf ( n3537 , R_148fd_102eb768 );
buf ( n3538 , R_14683_13a1d9c8 );
buf ( n3539 , R_a069_12080298 );
buf ( n3540 , R_1233a_13a143c8 );
buf ( n3541 , R_6e_13304b48 );
buf ( n3542 , R_1334f_1204e598 );
buf ( n3543 , R_121e7_1207ff78 );
buf ( n3544 , R_12bb7_102f3e68 );
buf ( n3545 , R_12bcc_12652608 );
buf ( n3546 , R_f783_13797b08 );
buf ( n3547 , R_14680_12076fb8 );
buf ( n3548 , R_13d2b_12085338 );
buf ( n3549 , R_11bbe_1153de38 );
buf ( n3550 , R_148e8_1264bda8 );
buf ( n3551 , R_148fa_102f5948 );
buf ( n3552 , R_149d8_132fc168 );
buf ( n3553 , R_148ee_120808d8 );
buf ( n3554 , R_148f4_11cd8468 );
buf ( n3555 , R_ff98_12b41618 );
buf ( n3556 , R_13bc3_102f8d28 );
buf ( n3557 , R_12b1f_120564d8 );
buf ( n3558 , R_c961_12080f18 );
buf ( n3559 , R_214_12655588 );
buf ( n3560 , R_dff5_102ed9c8 );
buf ( n3561 , R_13d49_13a16bc8 );
buf ( n3562 , R_fb_1379f808 );
buf ( n3563 , R_12958_102f1848 );
buf ( n3564 , R_12220_1379e908 );
buf ( n3565 , R_144de_12076798 );
buf ( n3566 , R_c6d1_10566178 );
buf ( n3567 , R_11547_1264cc08 );
buf ( n3568 , R_138ac_102eb128 );
buf ( n3569 , R_12853_105b58b8 );
buf ( n3570 , R_1f1_12655268 );
buf ( n3571 , R_11e_12b29b98 );
buf ( n3572 , R_13d30_1207b658 );
buf ( n3573 , R_b2_105aa0f8 );
buf ( n3574 , R_d5a1_105690f8 );
buf ( n3575 , R_c700_13304788 );
buf ( n3576 , R_a359_12662888 );
buf ( n3577 , R_1449f_12055898 );
buf ( n3578 , R_14587_10565ef8 );
buf ( n3579 , R_14759_1056e378 );
buf ( n3580 , R_1385d_1056ab38 );
buf ( n3581 , R_1401f_132fb588 );
buf ( n3582 , R_1245b_12658f68 );
buf ( n3583 , R_fe3a_11cdb168 );
buf ( n3584 , R_a47d_13a18f68 );
buf ( n3585 , R_145ea_1056c438 );
buf ( n3586 , R_99a4_102f5bc8 );
buf ( n3587 , R_1491e_12661528 );
buf ( n3588 , R_1c1_126618e8 );
buf ( n3589 , R_b180_12039a98 );
buf ( n3590 , R_14e_12b29e18 );
buf ( n3591 , R_13b1f_12052c38 );
buf ( n3592 , R_146e4_f8cb638 );
buf ( n3593 , R_14581_10571b18 );
buf ( n3594 , R_1354d_12040078 );
buf ( n3595 , R_13508_120842f8 );
buf ( n3596 , R_148d9_13a14d28 );
buf ( n3597 , R_149c0_102ed068 );
buf ( n3598 , R_1477e_10568fb8 );
buf ( n3599 , R_14735_105680b8 );
buf ( n3600 , R_13d35_11ce1108 );
buf ( n3601 , R_4d49_102f8dc8 );
buf ( n3602 , R_133aa_11545b38 );
buf ( n3603 , R_14518_102f67a8 );
buf ( n3604 , R_bf1d_1153d618 );
buf ( n3605 , R_a9_1204d4b8 );
buf ( n3606 , R_14702_12b3d0b8 );
buf ( n3607 , R_1431c_11cde188 );
buf ( n3608 , R_9323_1331d068 );
buf ( n3609 , R_14a2f_12075ed8 );
buf ( n3610 , R_1e1_13321ca8 );
buf ( n3611 , R_12e_105af9b8 );
buf ( n3612 , R_9d_1379c9c8 );
buf ( n3613 , R_12caa_126508a8 );
buf ( n3614 , R_115df_10566c18 );
buf ( n3615 , R_144fd_102f1b68 );
buf ( n3616 , R_127f1_12b2a098 );
buf ( n3617 , R_137eb_12082138 );
buf ( n3618 , R_11b9a_12b3f278 );
buf ( n3619 , R_1483a_12081f58 );
buf ( n3620 , R_7d2b_11ce4948 );
buf ( n3621 , R_13a49_102f8e68 );
buf ( n3622 , R_1493c_11cdc568 );
buf ( n3623 , R_14a3e_102ed428 );
buf ( n3624 , R_195_12045cb8 );
buf ( n3625 , R_14489_12b3fe58 );
buf ( n3626 , R_17a_1330dc48 );
buf ( n3627 , R_1066b_1264a228 );
buf ( n3628 , R_139b5_11536318 );
buf ( n3629 , R_12775_126513e8 );
buf ( n3630 , R_13d43_13a1c168 );
buf ( n3631 , R_13e78_1056a598 );
buf ( n3632 , R_90_f8cccb8 );
buf ( n3633 , R_75_12b443b8 );
buf ( n3634 , R_14816_10565db8 );
buf ( n3635 , R_e4c7_10571398 );
buf ( n3636 , R_14354_13317348 );
buf ( n3637 , R_146c3_12b3bfd8 );
buf ( n3638 , R_db95_12b2ff98 );
buf ( n3639 , R_b45b_11ce7508 );
buf ( n3640 , R_145de_1056b5d8 );
buf ( n3641 , R_13c7d_1056d798 );
buf ( n3642 , R_c7c0_102ed4c8 );
buf ( n3643 , R_1ff_13315c28 );
buf ( n3644 , R_1361a_102f01c8 );
buf ( n3645 , R_110_1204b938 );
buf ( n3646 , R_10c17_13a13888 );
buf ( n3647 , R_d6_1264b1c8 );
buf ( n3648 , R_239_12b2a958 );
buf ( n3649 , R_144a8_115369f8 );
buf ( n3650 , R_12516_13305188 );
buf ( n3651 , R_14699_10567e38 );
buf ( n3652 , R_12de4_12045b18 );
buf ( n3653 , R_10fd9_11ce1928 );
buf ( n3654 , R_145c6_13a1cb68 );
buf ( n3655 , R_147c3_13a177a8 );
buf ( n3656 , R_1313e_1207a1b8 );
buf ( n3657 , R_e9a6_1153dcf8 );
buf ( n3658 , R_123a6_12077418 );
buf ( n3659 , R_e669_1056eb98 );
buf ( n3660 , R_eea5_13793c88 );
buf ( n3661 , R_8e12_f8c7538 );
buf ( n3662 , R_11a2c_12b3f1d8 );
buf ( n3663 , R_bc89_12664548 );
buf ( n3664 , R_b132_13300a88 );
buf ( n3665 , R_14626_102f4ae8 );
buf ( n3666 , R_125c9_11ce5c08 );
buf ( n3667 , R_14891_1265e0a8 );
buf ( n3668 , R_13ba9_1056f4f8 );
buf ( n3669 , R_11299_1056a4f8 );
buf ( n3670 , R_1395f_1207ba18 );
buf ( n3671 , R_1085f_13312a28 );
buf ( n3672 , R_c642_12b41b18 );
buf ( n3673 , R_1445c_f8ce478 );
buf ( n3674 , R_14981_12b3f598 );
buf ( n3675 , R_148e2_12650b28 );
buf ( n3676 , R_988f_13a1e968 );
buf ( n3677 , R_962b_105647d8 );
buf ( n3678 , R_124a7_12079498 );
buf ( n3679 , R_fe64_1153f378 );
buf ( n3680 , R_11f16_102eb088 );
buf ( n3681 , R_13e03_1379bf28 );
buf ( n3682 , R_14927_11cdf808 );
buf ( n3683 , R_1ba_1330eb48 );
buf ( n3684 , R_14471_13793be8 );
buf ( n3685 , R_121fd_11ce3048 );
buf ( n3686 , R_14499_1207a9d8 );
buf ( n3687 , R_155_12b43f58 );
buf ( n3688 , R_98_12048af8 );
buf ( n3689 , R_e916_105699b8 );
buf ( n3690 , R_e1ea_1056b998 );
buf ( n3691 , R_11af3_13793788 );
buf ( n3692 , R_13bcf_12650948 );
buf ( n3693 , R_10070_12077e18 );
buf ( n3694 , R_f2f6_126613e8 );
buf ( n3695 , R_104a3_11542d98 );
buf ( n3696 , R_149ae_10565138 );
buf ( n3697 , R_1430b_1204c8d8 );
buf ( n3698 , R_ede8_1056dfb8 );
buf ( n3699 , R_13495_13a1e008 );
buf ( n3700 , R_df_132f6808 );
buf ( n3701 , R_230_12664a48 );
buf ( n3702 , R_136ac_102eacc8 );
buf ( n3703 , R_dd20_137974c8 );
buf ( n3704 , R_14741_132f2c08 );
buf ( n3705 , R_137c1_11543dd8 );
buf ( n3706 , R_14364_11ce6568 );
buf ( n3707 , R_11d60_132fc8e8 );
buf ( n3708 , R_14a44_105b60d8 );
buf ( n3709 , R_13749_11543518 );
buf ( n3710 , R_854a_1207fed8 );
buf ( n3711 , R_14a11_12045a78 );
buf ( n3712 , R_1a7_12659b48 );
buf ( n3713 , R_168_105b3158 );
buf ( n3714 , R_f03_13a17208 );
buf ( n3715 , R_1274c_12653fa8 );
buf ( n3716 , R_147b7_12079df8 );
buf ( n3717 , R_a2_1379e228 );
buf ( n3718 , R_63_f8c7b78 );
buf ( n3719 , R_13c49_102ecac8 );
buf ( n3720 , R_d68f_12078a98 );
buf ( n3721 , R_148f1_11cde688 );
buf ( n3722 , R_196_11536778 );
buf ( n3723 , R_179_13301c08 );
buf ( n3724 , R_11c1b_120757f8 );
buf ( n3725 , R_1181a_10565098 );
buf ( n3726 , R_14912_13300628 );
buf ( n3727 , R_10c93_13310768 );
buf ( n3728 , R_147f2_10571618 );
buf ( n3729 , R_c832_12075f78 );
buf ( n3730 , R_14530_11540778 );
buf ( n3731 , R_e8ba_11ce3b88 );
buf ( n3732 , R_14903_11ce50c8 );
buf ( n3733 , R_14629_115412b8 );
buf ( n3734 , R_11966_10562118 );
buf ( n3735 , R_f8fa_105b4d78 );
buf ( n3736 , R_1d8_1331f5e8 );
buf ( n3737 , R_1281b_1207f6b8 );
buf ( n3738 , R_137_1331a7c8 );
buf ( n3739 , R_5f_12b428d8 );
buf ( n3740 , R_12288_126495a8 );
buf ( n3741 , R_a469_13a14648 );
buf ( n3742 , R_130cc_13a17348 );
buf ( n3743 , R_136e6_11cdcb08 );
buf ( n3744 , R_d806_102f5a88 );
buf ( n3745 , R_fd98_12052d78 );
buf ( n3746 , R_144b4_1153eab8 );
buf ( n3747 , R_1482b_12b3b3f8 );
buf ( n3748 , R_13858_12081e18 );
buf ( n3749 , R_1d3_1265ae08 );
buf ( n3750 , R_13c_1265b1c8 );
buf ( n3751 , R_14596_12048558 );
buf ( n3752 , R_eb_1153bf98 );
buf ( n3753 , R_224_12b29698 );
buf ( n3754 , R_13d3c_132f70c8 );
buf ( n3755 , R_c353_102f31e8 );
buf ( n3756 , R_1092e_13a140a8 );
buf ( n3757 , R_1018e_10563478 );
buf ( n3758 , R_12875_1153eb58 );
buf ( n3759 , R_13693_13795448 );
buf ( n3760 , R_123bb_11ce7008 );
buf ( n3761 , R_dfc9_12647208 );
buf ( n3762 , R_da6d_12082098 );
buf ( n3763 , R_1198e_1153d758 );
buf ( n3764 , R_149ff_1264c848 );
buf ( n3765 , R_1180e_12648248 );
buf ( n3766 , R_12535_126604e8 );
buf ( n3767 , R_12780_10568b58 );
buf ( n3768 , R_9dc0_102f6f28 );
buf ( n3769 , R_c4a7_1330a908 );
buf ( n3770 , R_11bfb_12649968 );
buf ( n3771 , R_13fe4_105622f8 );
buf ( n3772 , R_12e0c_13797388 );
buf ( n3773 , R_1454e_11ce1c48 );
buf ( n3774 , R_14069_1153db18 );
buf ( n3775 , R_10c0e_120464d8 );
buf ( n3776 , R_13c1f_f8c8938 );
buf ( n3777 , R_d910_1056e418 );
buf ( n3778 , R_cfae_13a15368 );
buf ( n3779 , R_10806_1264d608 );
buf ( n3780 , R_13706_13319b48 );
buf ( n3781 , R_12e21_1330cb68 );
buf ( n3782 , R_f8_12665808 );
buf ( n3783 , R_67_105aac38 );
buf ( n3784 , R_217_105b3fb8 );
buf ( n3785 , R_12a8e_1264ef08 );
buf ( n3786 , R_e5ea_115436f8 );
buf ( n3787 , R_14858_10571c58 );
buf ( n3788 , R_111b8_102ebbc8 );
buf ( n3789 , R_12ba4_12b28ab8 );
buf ( n3790 , R_108f1_102f35a8 );
buf ( n3791 , R_138a5_1264e468 );
buf ( n3792 , R_131ff_13a1eaa8 );
buf ( n3793 , R_11448_11ce41c8 );
buf ( n3794 , R_11534_13a13ce8 );
buf ( n3795 , R_12d1d_1207c238 );
buf ( n3796 , R_134e8_13a1e8c8 );
buf ( n3797 , R_b82e_1153c2b8 );
buf ( n3798 , R_11572_11ce43a8 );
buf ( n3799 , R_14897_1265c988 );
buf ( n3800 , R_125fa_1265b128 );
buf ( n3801 , R_b95d_102f8008 );
buf ( n3802 , R_14436_10570718 );
buf ( n3803 , R_f951_132fcde8 );
buf ( n3804 , R_10246_1056ae58 );
buf ( n3805 , R_12041_11ce0ac8 );
buf ( n3806 , R_138cd_1153e018 );
buf ( n3807 , R_1b2_12660f88 );
buf ( n3808 , R_197_1379a768 );
buf ( n3809 , R_121dd_12659328 );
buf ( n3810 , R_178_12658d88 );
buf ( n3811 , R_15d_133195a8 );
buf ( n3812 , R_13f24_13318428 );
buf ( n3813 , R_146f6_132fbc68 );
buf ( n3814 , R_b880_12083d58 );
buf ( n3815 , R_12ab4_132f57c8 );
buf ( n3816 , R_ed14_133110c8 );
buf ( n3817 , R_144f0_132ff0e8 );
buf ( n3818 , R_10aa5_12053f98 );
buf ( n3819 , R_1290a_11ce1388 );
buf ( n3820 , R_9d4e_11cddbe8 );
buf ( n3821 , R_e6_12b344f8 );
buf ( n3822 , R_b0_12b3f458 );
buf ( n3823 , R_229_126659e8 );
buf ( n3824 , R_12b3f_105b6538 );
buf ( n3825 , R_1f5_1203e958 );
buf ( n3826 , R_f624_1265b808 );
buf ( n3827 , R_14711_11ce2828 );
buf ( n3828 , R_fe05_102f9548 );
buf ( n3829 , R_1118b_11cdb8e8 );
buf ( n3830 , R_1c8_f8c6b38 );
buf ( n3831 , R_147_12b38c98 );
buf ( n3832 , R_11a_1204b438 );
buf ( n3833 , R_14778_13a1f688 );
buf ( n3834 , R_137fd_11544418 );
buf ( n3835 , R_f0_13795d08 );
buf ( n3836 , R_c3_132ff188 );
buf ( n3837 , R_21f_1265a2c8 );
buf ( n3838 , R_12e60_132f3a68 );
buf ( n3839 , R_4a02_12646e48 );
buf ( n3840 , R_c5_12657e88 );
buf ( n3841 , R_132ae_1056ef58 );
buf ( n3842 , R_d400_133126a8 );
buf ( n3843 , R_128a8_f8c9978 );
buf ( n3844 , R_ecbd_12040a78 );
buf ( n3845 , R_146ba_11cd8c88 );
buf ( n3846 , R_ea59_102f5088 );
buf ( n3847 , R_1183a_1204a498 );
buf ( n3848 , R_13d1f_1207ddb8 );
buf ( n3849 , R_136e0_11ce7148 );
buf ( n3850 , R_ddb7_12078b38 );
buf ( n3851 , R_14575_13307c08 );
buf ( n3852 , R_14864_13a1b768 );
buf ( n3853 , R_1471d_12040bb8 );
buf ( n3854 , R_11237_1056f958 );
buf ( n3855 , R_13fee_12663288 );
buf ( n3856 , R_c1_1204fd58 );
buf ( n3857 , R_14632_11cd85a8 );
buf ( n3858 , R_4d_12662d88 );
buf ( n3859 , R_b895_1264a4a8 );
buf ( n3860 , R_11b87_12648b08 );
buf ( n3861 , R_111c4_12076658 );
buf ( n3862 , R_a534_12b3d018 );
buf ( n3863 , R_11805_12b41578 );
buf ( n3864 , R_c901_126603a8 );
buf ( n3865 , R_13bde_13a1bbc8 );
buf ( n3866 , R_149b4_10564d78 );
buf ( n3867 , R_c7_126589c8 );
buf ( n3868 , R_248_1331ef08 );
buf ( n3869 , R_5b_12655088 );
buf ( n3870 , R_13720_102f3f08 );
buf ( n3871 , R_b9b1_1056c9d8 );
buf ( n3872 , R_f1cc_10567ed8 );
buf ( n3873 , R_cd0b_11542f78 );
buf ( n3874 , R_1497b_11cdfda8 );
buf ( n3875 , R_12d6f_13799b88 );
buf ( n3876 , R_14305_120844d8 );
buf ( n3877 , R_145ae_102efe08 );
buf ( n3878 , R_147d6_12b27b18 );
buf ( n3879 , R_13dc3_11cdbf28 );
buf ( n3880 , R_dc22_1153d438 );
buf ( n3881 , R_5970_11cdbe88 );
buf ( n3882 , R_113_1265c528 );
buf ( n3883 , R_82_f8cbc78 );
buf ( n3884 , R_1fc_12050078 );
buf ( n3885 , R_b00a_1153e658 );
buf ( n3886 , R_1346e_10567bb8 );
buf ( n3887 , R_1dd_12b395f8 );
buf ( n3888 , R_10390_1207ed58 );
buf ( n3889 , R_12cf4_13310ee8 );
buf ( n3890 , R_10675_1203cab8 );
buf ( n3891 , R_1399b_1264c3e8 );
buf ( n3892 , R_132_120518d8 );
buf ( n3893 , R_d8_12b3c938 );
buf ( n3894 , R_237_105a9fb8 );
buf ( n3895 , R_d4b2_1265bda8 );
buf ( n3896 , R_14453_12649d28 );
buf ( n3897 , R_10e2c_102ecde8 );
buf ( n3898 , R_52_13799868 );
buf ( n3899 , R_143dc_120824f8 );
buf ( n3900 , R_13ebe_11ce4128 );
buf ( n3901 , R_14053_102f21a8 );
buf ( n3902 , R_10960_133050e8 );
buf ( n3903 , R_1037b_1264a048 );
buf ( n3904 , R_7fe6_12b3f638 );
buf ( n3905 , R_12685_11cdf088 );
buf ( n3906 , R_135e9_11ce0de8 );
buf ( n3907 , R_bf_1379fa88 );
buf ( n3908 , R_85_12b41898 );
buf ( n3909 , R_149d5_11541358 );
buf ( n3910 , R_13f4d_10561fd8 );
buf ( n3911 , R_d0f1_1056a1d8 );
buf ( n3912 , R_a3f3_12646da8 );
buf ( n3913 , R_1311d_13a131a8 );
buf ( n3914 , R_1026e_11541ad8 );
buf ( n3915 , R_139de_13310588 );
buf ( n3916 , R_144cc_11ce23c8 );
buf ( n3917 , R_1403a_1331cc08 );
buf ( n3918 , R_1ce_12656628 );
buf ( n3919 , R_198_12b3fdb8 );
buf ( n3920 , R_d37f_1379a1c8 );
buf ( n3921 , R_177_1330de28 );
buf ( n3922 , R_141_12b3cf78 );
buf ( n3923 , R_14500_102f92c8 );
buf ( n3924 , R_c9_12b28fb8 );
buf ( n3925 , R_246_1203df58 );
buf ( n3926 , R_93_12659be8 );
buf ( n3927 , R_72_132fe788 );
buf ( n3928 , R_125bf_105685b8 );
buf ( n3929 , R_1a8_137a0d48 );
buf ( n3930 , R_147a5_1264a728 );
buf ( n3931 , R_167_1204f678 );
buf ( n3932 , R_7f_105ac998 );
buf ( n3933 , R_149f0_13a1fea8 );
buf ( n3934 , R_12210_13793aa8 );
buf ( n3935 , R_13db7_11ce11a8 );
buf ( n3936 , R_100e9_132f3ec8 );
buf ( n3937 , R_5362_13a18108 );
buf ( n3938 , R_124d7_13a18e28 );
buf ( n3939 , R_14a55_133001c8 );
buf ( n3940 , R_12419_1153d398 );
buf ( n3941 , R_108b6_1264e0a8 );
buf ( n3942 , R_10d4d_11cded68 );
buf ( n3943 , R_1464a_13a15b88 );
buf ( n3944 , R_c7f2_11cdc748 );
buf ( n3945 , R_13c83_11544698 );
buf ( n3946 , R_1489a_f8c6c78 );
buf ( n3947 , R_125b6_12040b18 );
buf ( n3948 , R_c00b_12079718 );
buf ( n3949 , R_eeb_13a13608 );
buf ( n3950 , R_f088_1330ba88 );
buf ( n3951 , R_1365e_1207b838 );
buf ( n3952 , R_fa81_12052198 );
buf ( n3953 , R_145f3_13a14788 );
buf ( n3954 , R_10995_102f3148 );
buf ( n3955 , R_123f8_13a13388 );
buf ( n3956 , R_6358_1204fe98 );
buf ( n3957 , R_14763_11ce4c68 );
buf ( n3958 , R_1433c_12077c38 );
buf ( n3959 , R_dde7_13a141e8 );
buf ( n3960 , R_13ef9_1204a858 );
buf ( n3961 , R_14810_1056db58 );
buf ( n3962 , R_13fdc_102f15c8 );
buf ( n3963 , R_d995_11ce0fc8 );
buf ( n3964 , R_117fc_12056078 );
buf ( n3965 , R_8d57_11ce53e8 );
buf ( n3966 , R_11bb4_12b39cd8 );
buf ( n3967 , R_13b97_1207a438 );
buf ( n3968 , R_14068_11cdc108 );
buf ( n3969 , R_1335a_105b5ef8 );
buf ( n3970 , R_1043d_13a1c5c8 );
buf ( n3971 , R_128cf_11cdabc8 );
buf ( n3972 , R_1219b_1207a938 );
buf ( n3973 , R_10dce_105631f8 );
buf ( n3974 , R_bbfa_10564418 );
buf ( n3975 , R_11864_12b44318 );
buf ( n3976 , R_12435_11ce4088 );
buf ( n3977 , R_a7_1265a5e8 );
buf ( n3978 , R_111f4_11cdf6c8 );
buf ( n3979 , R_135cf_1207eb78 );
buf ( n3980 , R_102ef_1153c218 );
buf ( n3981 , R_12ca0_11ce0668 );
buf ( n3982 , R_1c2_1330f228 );
buf ( n3983 , R_c6f4_12056438 );
buf ( n3984 , R_1404f_12b3e738 );
buf ( n3985 , R_ee7b_1379a628 );
buf ( n3986 , R_127e9_f8c8078 );
buf ( n3987 , R_14d_1203cbf8 );
buf ( n3988 , R_bd_1203f3f8 );
buf ( n3989 , R_48_13301848 );
buf ( n3990 , R_10afa_13a15d68 );
buf ( n3991 , R_ed66_11ce3368 );
buf ( n3992 , R_13a92_102f0bc8 );
buf ( n3993 , R_e9fb_12646268 );
buf ( n3994 , R_10d30_12084078 );
buf ( n3995 , R_149ab_1153d7f8 );
buf ( n3996 , R_88_13300d08 );
buf ( n3997 , R_6b_105aaff8 );
buf ( n3998 , R_11c31_115418f8 );
buf ( n3999 , R_13677_102f9868 );
buf ( n4000 , R_133f2_1379f088 );
buf ( n4001 , R_13edf_120837b8 );
buf ( n4002 , R_d399_137980a8 );
buf ( n4003 , R_1446e_1207d958 );
buf ( n4004 , R_1382d_1207d9f8 );
buf ( n4005 , R_cb_1331fa48 );
buf ( n4006 , R_244_1264c708 );
buf ( n4007 , R_12dc8_13a1f548 );
buf ( n4008 , R_12299_1265d1a8 );
buf ( n4009 , R_1474a_12076dd8 );
buf ( n4010 , R_13844_12663aa8 );
buf ( n4011 , R_13c11_1153d578 );
buf ( n4012 , R_14650_1056f278 );
buf ( n4013 , R_146fc_12647848 );
buf ( n4014 , R_10f84_1207bab8 );
buf ( n4015 , R_131cc_12b272f8 );
buf ( n4016 , R_1451b_10567cf8 );
buf ( n4017 , R_14390_10567c58 );
buf ( n4018 , R_13754_12082318 );
buf ( n4019 , R_1bb_12664868 );
buf ( n4020 , R_154_1204e1d8 );
buf ( n4021 , R_14831_1264f408 );
buf ( n4022 , R_7c_105b1cb8 );
buf ( n4023 , R_f1a0_12075938 );
buf ( n4024 , R_e9d0_1153f558 );
buf ( n4025 , R_f0eb_102f7568 );
buf ( n4026 , R_fb0c_1331a368 );
buf ( n4027 , R_1397b_1331b268 );
buf ( n4028 , R_e589_1379bb68 );
buf ( n4029 , R_1381a_120547b8 );
buf ( n4030 , R_1463e_105703f8 );
buf ( n4031 , R_12e76_11cd9908 );
buf ( n4032 , R_199_132fb3a8 );
buf ( n4033 , R_176_12b265d8 );
buf ( n4034 , R_125_13798008 );
buf ( n4035 , R_11ad2_102ed108 );
buf ( n4036 , R_1ea_1265a868 );
buf ( n4037 , R_10764_11cd9548 );
buf ( n4038 , R_14563_1264d6a8 );
buf ( n4039 , R_12c1a_102f0268 );
buf ( n4040 , R_146d2_1203a998 );
buf ( n4041 , R_147bd_102f9048 );
buf ( n4042 , R_fa57_1207f398 );
buf ( n4043 , R_c5a3_120849d8 );
buf ( n4044 , R_11dc9_f8c9b58 );
buf ( n4045 , R_11d95_1153f198 );
buf ( n4046 , R_1329b_11cd95e8 );
buf ( n4047 , R_14861_f8c41f8 );
buf ( n4048 , R_1064a_10561f38 );
buf ( n4049 , R_ce07_f8c8f78 );
buf ( n4050 , R_14720_11ce07a8 );
buf ( n4051 , R_13ca7_12078098 );
buf ( n4052 , R_147f5_1207a078 );
buf ( n4053 , R_142d3_12036758 );
buf ( n4054 , R_13dee_12083a38 );
buf ( n4055 , R_ec91_126490a8 );
buf ( n4056 , R_13421_11544c38 );
buf ( n4057 , R_cf92_11cdfee8 );
buf ( n4058 , R_4c49_13a1d748 );
buf ( n4059 , R_114d1_13307de8 );
buf ( n4060 , R_cff7_12076bf8 );
buf ( n4061 , R_142ff_11ce1b08 );
buf ( n4062 , R_139c0_13a1e5a8 );
buf ( n4063 , R_143cc_1056e738 );
buf ( n4064 , R_ba4e_13a1d388 );
buf ( n4065 , R_12485_105b6358 );
buf ( n4066 , R_11f0c_13a1aea8 );
buf ( n4067 , R_14867_12054b78 );
buf ( n4068 , R_137b5_10569cd8 );
buf ( n4069 , R_11d1b_12649288 );
buf ( n4070 , R_13d7b_102f56c8 );
buf ( n4071 , R_14a2c_102f12a8 );
buf ( n4072 , R_14608_13a155e8 );
buf ( n4073 , R_144c9_10571578 );
buf ( n4074 , R_fc0a_11541858 );
buf ( n4075 , R_144fa_120775f8 );
buf ( n4076 , R_129_1331c988 );
buf ( n4077 , R_13561_1330d068 );
buf ( n4078 , R_e1_12661708 );
buf ( n4079 , R_1299a_1207b158 );
buf ( n4080 , R_1489d_105686f8 );
buf ( n4081 , R_22e_132f2ac8 );
buf ( n4082 , R_6d01_102f72e8 );
buf ( n4083 , R_ffc3_12656e48 );
buf ( n4084 , R_1496f_102f9908 );
buf ( n4085 , R_1e6_13792a68 );
buf ( n4086 , R_14760_11ce3868 );
buf ( n4087 , R_d2d1_13793468 );
buf ( n4088 , R_12145_1207b978 );
buf ( n4089 , R_f5_11537038 );
buf ( n4090 , R_bb_13799cc8 );
buf ( n4091 , R_21a_1265b088 );
buf ( n4092 , R_14975_11541998 );
buf ( n4093 , R_147c0_11ce20a8 );
buf ( n4094 , R_13b7f_1153a198 );
buf ( n4095 , R_13615_12084c58 );
buf ( n4096 , R_14a29_10571438 );
buf ( n4097 , R_13526_102f49a8 );
buf ( n4098 , R_11215_12075b18 );
buf ( n4099 , R_10e4c_13a169e8 );
buf ( n4100 , R_13d97_105651d8 );
buf ( n4101 , R_1b3_1379b348 );
buf ( n4102 , R_13fab_11538758 );
buf ( n4103 , R_10ff9_105aad78 );
buf ( n4104 , R_145c0_11cd7f68 );
buf ( n4105 , R_145fc_120476f8 );
buf ( n4106 , R_15c_137992c8 );
buf ( n4107 , R_67bc_13311028 );
buf ( n4108 , R_efc2_11cdefe8 );
buf ( n4109 , R_145cc_132f8388 );
buf ( n4110 , R_ae_1379c1a8 );
buf ( n4111 , R_1263c_11cdf768 );
buf ( n4112 , R_57_126522e8 );
buf ( n4113 , R_14659_1264e1e8 );
buf ( n4114 , R_13899_133075c8 );
buf ( n4115 , R_125e5_13311348 );
buf ( n4116 , R_113fb_11ce7288 );
buf ( n4117 , R_11e0e_102f4908 );
buf ( n4118 , R_11270_12b29a58 );
buf ( n4119 , R_f61a_13305cc8 );
buf ( n4120 , R_1499f_133198c8 );
buf ( n4121 , R_121_13795808 );
buf ( n4122 , R_106_12b25a98 );
buf ( n4123 , R_1458a_102eb268 );
buf ( n4124 , R_126cf_13a19788 );
buf ( n4125 , R_209_1379cb08 );
buf ( n4126 , R_1ee_12656268 );
buf ( n4127 , R_12c5a_102ef688 );
buf ( n4128 , R_1270e_11cdb708 );
buf ( n4129 , R_e437_102f2c48 );
buf ( n4130 , R_147cf_11ce5168 );
buf ( n4131 , R_e233_1056d338 );
buf ( n4132 , R_13bbe_11ce55c8 );
buf ( n4133 , R_11e6b_1207d458 );
buf ( n4134 , R_13f0b_12b42f18 );
buf ( n4135 , R_103_12b41c58 );
buf ( n4136 , R_cd_12b39a58 );
buf ( n4137 , R_242_12654688 );
buf ( n4138 , R_20c_12b43c38 );
buf ( n4139 , R_11ce5_1379e048 );
buf ( n4140 , R_ef4_1056dc98 );
buf ( n4141 , R_11823_13a15fe8 );
buf ( n4142 , R_130b8_13a12988 );
buf ( n4143 , R_12baf_12648ba8 );
buf ( n4144 , R_119a4_102f3288 );
buf ( n4145 , R_f4e5_1264b308 );
buf ( n4146 , R_12c6f_11cdea48 );
buf ( n4147 , R_1473b_102fa308 );
buf ( n4148 , R_8b_132f8608 );
buf ( n4149 , R_11467_105659f8 );
buf ( n4150 , R_11b4a_11ce1568 );
buf ( n4151 , R_137f7_12077878 );
buf ( n4152 , R_e5b5_1153d938 );
buf ( n4153 , R_14775_13a1bda8 );
buf ( n4154 , R_14671_1264ab88 );
buf ( n4155 , R_14066_12084258 );
buf ( n4156 , R_13954_12076518 );
buf ( n4157 , R_de4d_12b26538 );
buf ( n4158 , R_149f6_11cda308 );
buf ( n4159 , R_aff6_102f4a48 );
buf ( n4160 , R_d75d_1207c0f8 );
buf ( n4161 , R_10f46_12081ff8 );
buf ( n4162 , R_c50b_11cdd3c8 );
buf ( n4163 , R_136ed_12082ef8 );
buf ( n4164 , R_101d1_1056e198 );
buf ( n4165 , R_1a9_12037658 );
buf ( n4166 , R_166_120507f8 );
buf ( n4167 , R_9b_12b3b178 );
buf ( n4168 , R_bb16_12650268 );
buf ( n4169 , R_1265a_105635b8 );
buf ( n4170 , R_b802_1265dba8 );
buf ( n4171 , R_131ea_102f4cc8 );
buf ( n4172 , R_14a0e_10570e98 );
buf ( n4173 , R_19a_12662068 );
buf ( n4174 , R_175_12b3fc78 );
buf ( n4175 , R_109_12b2c7f8 );
buf ( n4176 , R_206_105b5b38 );
buf ( n4177 , R_146b4_1153fcd8 );
buf ( n4178 , R_11e21_11cd9e08 );
buf ( n4179 , R_104ba_f8c7218 );
buf ( n4180 , R_13fbc_11541218 );
buf ( n4181 , R_144ba_102f8c88 );
buf ( n4182 , R_11622_102ed388 );
buf ( n4183 , R_13c02_12b29198 );
buf ( n4184 , R_13ba3_105626b8 );
buf ( n4185 , R_ff0f_12081918 );
buf ( n4186 , R_123d6_11541e98 );
buf ( n4187 , R_fd64_102f3328 );
buf ( n4188 , R_14486_102ef728 );
buf ( n4189 , R_13776_1379fd08 );
buf ( n4190 , R_14665_132f5ae8 );
buf ( n4191 , R_10098_13793968 );
buf ( n4192 , R_11072_13a1ed28 );
buf ( n4193 , R_14554_10565778 );
buf ( n4194 , R_137a8_1056b678 );
buf ( n4195 , R_11b55_12649a08 );
buf ( n4196 , R_14411_12663508 );
buf ( n4197 , R_84a7_12b40fd8 );
buf ( n4198 , R_133fc_1153ee78 );
buf ( n4199 , R_da_1331b088 );
buf ( n4200 , R_a0_1379b2a8 );
buf ( n4201 , R_235_1264d4c8 );
buf ( n4202 , R_1333b_11542c58 );
buf ( n4203 , R_132e7_11ce28c8 );
buf ( n4204 , R_1357d_1153feb8 );
buf ( n4205 , R_14644_1056d978 );
buf ( n4206 , R_100_1265f0e8 );
buf ( n4207 , R_79_137a1388 );
buf ( n4208 , R_e0d7_126556c8 );
buf ( n4209 , R_11b42_1264b6c8 );
buf ( n4210 , R_20f_12b28018 );
buf ( n4211 , R_f4db_1207bfb8 );
buf ( n4212 , R_1193e_13a19968 );
buf ( n4213 , R_138d5_1379b848 );
buf ( n4214 , R_13e4c_1207f118 );
buf ( n4215 , R_13a7e_102f6ac8 );
buf ( n4216 , R_12d79_102ee468 );
buf ( n4217 , R_116a8_12084398 );
buf ( n4218 , R_116_1265f868 );
buf ( n4219 , R_148a3_11cdecc8 );
buf ( n4220 , R_13273_13a1a688 );
buf ( n4221 , R_1f9_1379ddc8 );
buf ( n4222 , R_1025b_1330bee8 );
buf ( n4223 , R_122e8_12b39878 );
buf ( n4224 , R_11ba2_11544738 );
buf ( n4225 , R_12521_1056c258 );
buf ( n4226 , R_e8e6_f8cf4b8 );
buf ( n4227 , R_8cd2_1264ac28 );
buf ( n4228 , R_11a11_126477a8 );
buf ( n4229 , R_143c6_120850b8 );
buf ( n4230 , R_13e99_12039e58 );
buf ( n4231 , R_1466b_13306808 );
buf ( n4232 , R_14465_1207a758 );
buf ( n4233 , R_134b3_102f3468 );
buf ( n4234 , R_11fe7_1330c3e8 );
buf ( n4235 , R_1258d_13a14dc8 );
buf ( n4236 , R_14677_105712f8 );
buf ( n4237 , R_1367d_102eb628 );
buf ( n4238 , R_1e2_12663c88 );
buf ( n4239 , R_b9_12661848 );
buf ( n4240 , R_12d_12660268 );
buf ( n4241 , R_f47c_1153ded8 );
buf ( n4242 , R_1468c_13a1aae8 );
buf ( n4243 , R_145ba_120815f8 );
buf ( n4244 , R_14790_11cd9cc8 );
buf ( n4245 , R_14419_12048f58 );
buf ( n4246 , R_13bb3_1207b6f8 );
buf ( n4247 , R_1046b_105688d8 );
buf ( n4248 , R_1232e_13314008 );
buf ( n4249 , R_1170d_1264c528 );
buf ( n4250 , R_14a41_1056fa98 );
buf ( n4251 , R_14459_11cd92c8 );
buf ( n4252 , R_14480_11cdcf68 );
buf ( n4253 , R_13a88_11ce3f48 );
buf ( n4254 , R_c8f0_102f0d08 );
buf ( n4255 , R_134ff_1056bf38 );
buf ( n4256 , R_aac5_13a18748 );
buf ( n4257 , R_14509_13a1e148 );
buf ( n4258 , R_cebc_12039d18 );
buf ( n4259 , R_135bd_12081058 );
buf ( n4260 , R_147ba_12078ef8 );
buf ( n4261 , R_f4a6_105654f8 );
buf ( n4262 , R_1182e_13a19aa8 );
buf ( n4263 , R_142eb_11cdec28 );
buf ( n4264 , R_13bf5_10568ab8 );
buf ( n4265 , R_12093_12077058 );
buf ( n4266 , R_13dac_13a15688 );
buf ( n4267 , R_dc51_13304f08 );
buf ( n4268 , R_13e8f_1264a0e8 );
buf ( n4269 , R_13c89_12b39f58 );
buf ( n4270 , R_f0be_102f1de8 );
buf ( n4271 , R_9373_10563e78 );
buf ( n4272 , R_11a48_13a195a8 );
buf ( n4273 , R_f3f9_1153f9b8 );
buf ( n4274 , R_1d4_12b42fb8 );
buf ( n4275 , R_e3f1_12b25bd8 );
buf ( n4276 , R_13c27_13309b48 );
buf ( n4277 , R_240_105ab4f8 );
buf ( n4278 , R_cf_13311a28 );
buf ( n4279 , R_13c38_1204a3f8 );
buf ( n4280 , R_13b_13300f88 );
buf ( n4281 , R_11ef6_11cd7888 );
buf ( n4282 , R_135c9_11ce6888 );
buf ( n4283 , R_116d1_1153d898 );
buf ( n4284 , R_149d2_12080158 );
buf ( n4285 , R_ba5b_12b403f8 );
buf ( n4286 , R_ea84_1330ca28 );
buf ( n4287 , R_f59a_11ce3908 );
buf ( n4288 , R_1496c_1331e968 );
buf ( n4289 , R_12bd5_11ce3fe8 );
buf ( n4290 , R_1253e_105b6678 );
buf ( n4291 , R_14873_11cd79c8 );
buf ( n4292 , R_149a5_132ff868 );
buf ( n4293 , R_14512_11540bd8 );
buf ( n4294 , R_14756_10565318 );
buf ( n4295 , R_1c9_13313a68 );
buf ( n4296 , R_d09b_12660948 );
buf ( n4297 , R_203_12050cf8 );
buf ( n4298 , R_10c_12038058 );
buf ( n4299 , R_146_12b42298 );
buf ( n4300 , R_136c1_12b276b8 );
buf ( n4301 , R_1480a_12649e68 );
buf ( n4302 , R_1d9_1379e7c8 );
buf ( n4303 , R_13e84_1056ad18 );
buf ( n4304 , R_1021c_1056fc78 );
buf ( n4305 , R_136_132fe6e8 );
buf ( n4306 , R_145ff_102ef2c8 );
buf ( n4307 , R_19b_12b28dd8 );
buf ( n4308 , R_1031a_11540e58 );
buf ( n4309 , R_1f2_11538438 );
buf ( n4310 , R_13114_102f3648 );
buf ( n4311 , R_ec36_12042af8 );
buf ( n4312 , R_222_133189c8 );
buf ( n4313 , R_6f_12b3a458 );
buf ( n4314 , R_96_1203c838 );
buf ( n4315 , R_ed_1203deb8 );
buf ( n4316 , R_11d_1204c838 );
buf ( n4317 , R_174_13318928 );
buf ( n4318 , R_119f1_13316588 );
buf ( n4319 , R_1486a_13a1d428 );
buf ( n4320 , R_11717_1207d778 );
buf ( n4321 , R_14781_115447d8 );
buf ( n4322 , R_13995_12038738 );
buf ( n4323 , R_e4f5_12049598 );
buf ( n4324 , R_74a9_12645d68 );
buf ( n4325 , R_10208_12038558 );
buf ( n4326 , R_145ab_12b3f9f8 );
buf ( n4327 , R_227_1331e508 );
buf ( n4328 , R_e8_133028e8 );
buf ( n4329 , R_13809_1153faf8 );
buf ( n4330 , R_f732_12649008 );
buf ( n4331 , R_14524_137968e8 );
buf ( n4332 , R_146d8_11cd94a8 );
buf ( n4333 , R_14064_1264d2e8 );
buf ( n4334 , R_12dfa_11cd88c8 );
buf ( n4335 , R_135ef_102f0a88 );
buf ( n4336 , R_10ee5_12047798 );
buf ( n4337 , R_14548_120493b8 );
buf ( n4338 , R_11030_11cdbca8 );
buf ( n4339 , R_1400f_13a1a368 );
buf ( n4340 , R_f051_1264e6e8 );
buf ( n4341 , R_de7c_102eafe8 );
buf ( n4342 , R_13538_120754d8 );
buf ( n4343 , R_13e56_12b297d8 );
buf ( n4344 , R_84eb_1331c2a8 );
buf ( n4345 , R_1498a_1207e3f8 );
buf ( n4346 , R_148a6_115459f8 );
buf ( n4347 , R_212_1330bd08 );
buf ( n4348 , R_fd_13307d48 );
buf ( n4349 , R_144a5_13a1c028 );
buf ( n4350 , R_10110_120369d8 );
buf ( n4351 , R_12b5e_12651208 );
buf ( n4352 , R_149ed_13303428 );
buf ( n4353 , R_144db_12078598 );
buf ( n4354 , R_bf9f_11cd9b88 );
buf ( n4355 , R_14017_f8c20d8 );
buf ( n4356 , R_13a3d_f8ca918 );
buf ( n4357 , R_13b2d_120830d8 );
buf ( n4358 , R_8e_132f37e8 );
buf ( n4359 , R_12aeb_120810f8 );
buf ( n4360 , R_a23e_11ce5ca8 );
buf ( n4361 , R_12ce9_12081c38 );
buf ( n4362 , R_f00_1207c058 );
buf ( n4363 , R_c1fe_1264be48 );
buf ( n4364 , R_f2d2_11cdf948 );
buf ( n4365 , R_14385_12044c18 );
buf ( n4366 , R_143c0_1265fb88 );
buf ( n4367 , R_14496_13a1c668 );
buf ( n4368 , R_14738_12b28bf8 );
buf ( n4369 , R_cab9_102f99a8 );
buf ( n4370 , R_1255c_f8c61d8 );
buf ( n4371 , R_143ba_11cde868 );
buf ( n4372 , R_147c9_13a18ce8 );
buf ( n4373 , R_13311_13a198c8 );
buf ( n4374 , R_147a2_102f2ce8 );
buf ( n4375 , R_fbe0_13a1b628 );
buf ( n4376 , R_dcc6_12664ae8 );
buf ( n4377 , R_103cf_12085158 );
buf ( n4378 , R_13909_1204f5d8 );
buf ( n4379 , R_1197b_115433d8 );
buf ( n4380 , R_144e1_13a1f4a8 );
buf ( n4381 , R_145a2_11cd7ce8 );
buf ( n4382 , R_12d50_120851f8 );
buf ( n4383 , R_12380_10563338 );
buf ( n4384 , R_107a7_1379f9e8 );
buf ( n4385 , R_10e8a_102ea688 );
buf ( n4386 , R_122fb_13a17708 );
buf ( n4387 , R_12aa7_12037798 );
buf ( n4388 , R_12107_1264d428 );
buf ( n4389 , R_14533_1330c8e8 );
buf ( n4390 , R_14542_120759d8 );
buf ( n4391 , R_4276_102effe8 );
buf ( n4392 , R_1478d_115453b8 );
buf ( n4393 , R_130c1_11542258 );
buf ( n4394 , R_13ff8_102f9fe8 );
buf ( n4395 , R_1aa_13795268 );
buf ( n4396 , R_116b1_13a159a8 );
buf ( n4397 , R_1bc_126536e8 );
buf ( n4398 , R_b76e_1153c8f8 );
buf ( n4399 , R_4e_13792e28 );
buf ( n4400 , R_60_12b44bd8 );
buf ( n4401 , R_a5_13311668 );
buf ( n4402 , R_b7_1379f948 );
buf ( n4403 , R_153_13793288 );
buf ( n4404 , R_165_13306948 );
buf ( n4405 , R_f9fe_102f9408 );
buf ( n4406 , R_14431_12080478 );
buf ( n4407 , R_1c3_12047158 );
buf ( n4408 , R_64_f8c1bd8 );
buf ( n4409 , R_14c_120387d8 );
buf ( n4410 , R_12471_102f7068 );
buf ( n4411 , R_148c1_13316f88 );
buf ( n4412 , R_11433_1265f048 );
buf ( n4413 , R_13ce2_1264aa48 );
buf ( n4414 , R_121bd_115449b8 );
buf ( n4415 , R_14813_10566d58 );
buf ( n4416 , R_147fb_102f83c8 );
buf ( n4417 , R_146ab_12051658 );
buf ( n4418 , R_12c65_1264cb68 );
buf ( n4419 , R_e2b4_f8c0f58 );
buf ( n4420 , R_10c61_120805b8 );
buf ( n4421 , R_10f1d_10566df8 );
buf ( n4422 , R_10de4_1379b5c8 );
buf ( n4423 , R_ae51_105ab098 );
buf ( n4424 , R_146f3_12659d28 );
buf ( n4425 , R_d03f_126484c8 );
buf ( n4426 , R_9fe2_11543fb8 );
buf ( n4427 , R_10b79_12657028 );
buf ( n4428 , R_64c2_12662748 );
buf ( n4429 , R_139d0_102f1fc8 );
buf ( n4430 , R_13639_1207f578 );
buf ( n4431 , R_1b4_12654728 );
buf ( n4432 , R_1cf_133184c8 );
buf ( n4433 , R_e214_1207ae38 );
buf ( n4434 , R_140_12665448 );
buf ( n4435 , R_15b_f8c0378 );
buf ( n4436 , R_1435c_13304d28 );
buf ( n4437 , R_10745_12056898 );
buf ( n4438 , R_1044f_120557f8 );
buf ( n4439 , R_10824_11ce3188 );
buf ( n4440 , R_13820_12b41438 );
buf ( n4441 , R_69b8_11cdc888 );
buf ( n4442 , R_124b9_1056d658 );
buf ( n4443 , R_143f4_102edd88 );
buf ( n4444 , R_142f5_1264a908 );
buf ( n4445 , R_76_f8ca198 );
buf ( n4446 , R_ac_12660a88 );
buf ( n4447 , R_1269b_11cd9368 );
buf ( n4448 , R_147b4_120766f8 );
buf ( n4449 , R_14834_13a16a88 );
buf ( n4450 , R_12e88_102f8a08 );
buf ( n4451 , R_f021_102ec168 );
buf ( n4452 , R_f6dd_13a163a8 );
buf ( n4453 , R_145e4_126463a8 );
buf ( n4454 , R_14723_1264db08 );
buf ( n4455 , R_173_f8c3438 );
buf ( n4456 , R_19c_12b40218 );
buf ( n4457 , R_11142_10562f78 );
buf ( n4458 , R_23e_1265bc68 );
buf ( n4459 , R_d1_13311f28 );
buf ( n4460 , R_13512_12080dd8 );
buf ( n4461 , R_7859_11cdaee8 );
buf ( n4462 , R_14593_115458b8 );
buf ( n4463 , R_148a9_12647ac8 );
buf ( n4464 , R_10577_11545318 );
buf ( n4465 , R_133ca_1203e098 );
buf ( n4466 , R_13b92_13a14be8 );
buf ( n4467 , R_10efd_102ec3e8 );
buf ( n4468 , R_f0b_1153f4b8 );
buf ( n4469 , R_12e15_10568018 );
buf ( n4470 , R_200_12b29eb8 );
buf ( n4471 , R_21d_137a03e8 );
buf ( n4472 , R_f2_12652ec8 );
buf ( n4473 , R_10f_12b3e5f8 );
buf ( n4474 , R_ca13_11ce4628 );
buf ( n4475 , R_14966_11546218 );
buf ( n4476 , R_13ad8_1203a358 );
buf ( n4477 , R_12d8d_105b5db8 );
buf ( n4478 , R_10165_1264cac8 );
buf ( n4479 , R_1337f_13a12c08 );
buf ( n4480 , R_53_f8c2a38 );
buf ( n4481 , R_149c9_132f4fa8 );
buf ( n4482 , R_10aae_1207c558 );
buf ( n4483 , R_13aad_11541a38 );
buf ( n4484 , R_12362_10563dd8 );
buf ( n4485 , R_5c4e_1056ced8 );
buf ( n4486 , R_130f5_1056a098 );
buf ( n4487 , R_12a7c_11cdde68 );
buf ( n4488 , R_14415_12b2a318 );
buf ( n4489 , R_1488b_13a189c8 );
buf ( n4490 , R_14062_1204cf18 );
buf ( n4491 , R_14784_11cd8508 );
buf ( n4492 , R_1032f_10570f38 );
buf ( n4493 , R_9bdf_102ee5a8 );
buf ( n4494 , R_13bf0_1331c528 );
buf ( n4495 , R_11b90_11ce0208 );
buf ( n4496 , R_149cf_13a17b68 );
buf ( n4497 , R_12021_11ce25a8 );
buf ( n4498 , R_1de_12056d98 );
buf ( n4499 , R_49_1331f4a8 );
buf ( n4500 , R_131_105ab3b8 );
buf ( n4501 , R_1462f_13794688 );
buf ( n4502 , R_10628_1203d2d8 );
buf ( n4503 , R_122bf_10570038 );
buf ( n4504 , R_11387_11540d18 );
buf ( n4505 , R_11fa6_13306308 );
buf ( n4506 , R_85b5_120819b8 );
buf ( n4507 , R_142ef_102eec88 );
buf ( n4508 , R_1434c_102f13e8 );
buf ( n4509 , R_22c_1379b708 );
buf ( n4510 , R_5c_137944a8 );
buf ( n4511 , R_e3_1203e778 );
buf ( n4512 , R_b948_1153a5f8 );
buf ( n4513 , R_e169_11cd7a68 );
buf ( n4514 , R_d051_11536ef8 );
buf ( n4515 , R_10e01_120551b8 );
buf ( n4516 , R_233_12b392d8 );
buf ( n4517 , R_68_12b283d8 );
buf ( n4518 , R_dc_13300768 );
buf ( n4519 , R_13bfb_13316a88 );
buf ( n4520 , R_10ad6_10565598 );
buf ( n4521 , R_14870_10570538 );
buf ( n4522 , R_12260_13a1b268 );
buf ( n4523 , R_d661_1265cfc8 );
buf ( n4524 , R_14572_11cd9d68 );
buf ( n4525 , R_130ff_12078318 );
buf ( n4526 , R_a98a_11cdaf88 );
buf ( n4527 , R_14978_12b321f8 );
buf ( n4528 , R_14a1a_115445f8 );
buf ( n4529 , R_14a26_13792568 );
buf ( n4530 , R_b327_12648568 );
buf ( n4531 , R_108fb_105b5e58 );
buf ( n4532 , R_1440d_11544238 );
buf ( n4533 , R_10cff_13a1dc48 );
buf ( n4534 , R_139ae_11cd8b48 );
buf ( n4535 , R_14338_11cda808 );
buf ( n4536 , R_106b3_13a16088 );
buf ( n4537 , R_c4f8_11ce12e8 );
buf ( n4538 , R_215_1265b948 );
buf ( n4539 , R_fa_133070c8 );
buf ( n4540 , R_11b68_1264ec88 );
buf ( n4541 , R_129b1_1056f098 );
buf ( n4542 , R_13670_10564558 );
buf ( n4543 , R_1439c_11cdd148 );
buf ( n4544 , R_107e6_11cdbc08 );
buf ( n4545 , R_f279_13a1acc8 );
buf ( n4546 , R_12ed9_102edf68 );
buf ( n4547 , R_12bc1_13a1f048 );
buf ( n4548 , R_13b19_12b2ba38 );
buf ( n4549 , R_e361_120812d8 );
buf ( n4550 , R_bef9_11ce0528 );
buf ( n4551 , R_13ce8_120793f8 );
buf ( n4552 , R_a235_12084a78 );
buf ( n4553 , R_14521_1264f228 );
buf ( n4554 , R_13cad_13a1edc8 );
buf ( n4555 , R_148af_11540098 );
buf ( n4556 , R_10968_13304968 );
buf ( n4557 , R_13fcb_102f0c68 );
buf ( n4558 , R_11645_13304e68 );
buf ( n4559 , R_bf09_1056b498 );
buf ( n4560 , R_12553_13310308 );
buf ( n4561 , R_145d5_132fa228 );
buf ( n4562 , R_146a2_1207bf18 );
buf ( n4563 , R_136fc_12076018 );
buf ( n4564 , R_149a2_1264d1a8 );
buf ( n4565 , R_12b9a_13a14968 );
buf ( n4566 , R_137cc_10569af8 );
buf ( n4567 , R_c5ef_12081238 );
buf ( n4568 , R_1184d_11cd9188 );
buf ( n4569 , R_13c8f_102ed568 );
buf ( n4570 , R_109bf_1379c248 );
buf ( n4571 , R_14326_13301528 );
buf ( n4572 , R_11123_12045258 );
buf ( n4573 , R_e197_11ce3228 );
buf ( n4574 , R_172_126656c8 );
buf ( n4575 , R_19d_132ffb88 );
buf ( n4576 , R_c306_f8c5418 );
buf ( n4577 , R_b5_133157c8 );
buf ( n4578 , R_13902_13799ae8 );
buf ( n4579 , R_14348_1056c398 );
buf ( n4580 , R_1457b_102f5628 );
buf ( n4581 , R_14766_105674d8 );
buf ( n4582 , R_d2c1_12036e38 );
buf ( n4583 , R_1f6_1330dce8 );
buf ( n4584 , R_10c28_12080e78 );
buf ( n4585 , R_119_133166c8 );
buf ( n4586 , R_1300e_12646bc8 );
buf ( n4587 , R_13129_10567b18 );
buf ( n4588 , R_1394d_1056f318 );
buf ( n4589 , R_14846_13798b48 );
buf ( n4590 , R_146cf_1379e868 );
buf ( n4591 , R_10019_11542118 );
buf ( n4592 , R_fb35_132fb4e8 );
buf ( n4593 , R_11a23_126506c8 );
buf ( n4594 , R_9aae_1056dbf8 );
buf ( n4595 , R_14468_1264aea8 );
buf ( n4596 , R_7aaf_f8c22b8 );
buf ( n4597 , R_b5af_1264e508 );
buf ( n4598 , R_13f11_11cd7b08 );
buf ( n4599 , R_e6c6_12075cf8 );
buf ( n4600 , R_14374_102f0768 );
buf ( n4601 , R_14605_13a182e8 );
buf ( n4602 , R_13de4_102f94a8 );
buf ( n4603 , R_102c2_1264ed28 );
buf ( n4604 , R_91_13799548 );
buf ( n4605 , R_135f5_11cda4e8 );
buf ( n4606 , R_14807_1331e288 );
buf ( n4607 , R_14a08_11cdc388 );
buf ( n4608 , R_cb44_12b3ee18 );
buf ( n4609 , R_13a63_11544198 );
buf ( n4610 , R_109ca_1264cd48 );
buf ( n4611 , R_12e41_10569198 );
buf ( n4612 , R_e46a_13a181a8 );
buf ( n4613 , R_12963_13a1afe8 );
buf ( n4614 , R_14a5a_12b42158 );
buf ( n4615 , R_13e38_1207efd8 );
buf ( n4616 , R_144ea_1264f5e8 );
buf ( n4617 , R_11668_137a1d88 );
buf ( n4618 , R_13ec7_11540318 );
buf ( n4619 , R_ff67_13799688 );
buf ( n4620 , R_13b27_102eb588 );
buf ( n4621 , R_fa2a_1056e0f8 );
buf ( n4622 , R_145a5_132f4dc8 );
buf ( n4623 , R_14060_13a15ae8 );
buf ( n4624 , R_164_12b27118 );
buf ( n4625 , R_104d9_120779b8 );
buf ( n4626 , R_1ab_f8c2998 );
buf ( n4627 , R_23c_13319328 );
buf ( n4628 , R_bbdf_133063a8 );
buf ( n4629 , R_d3_12659968 );
buf ( n4630 , R_cc7b_13a1b128 );
buf ( n4631 , R_12ffe_1331cd48 );
buf ( n4632 , R_1323e_126561c8 );
buf ( n4633 , R_1207f_133190a8 );
buf ( n4634 , R_10f99_126549a8 );
buf ( n4635 , R_913d_12646b28 );
buf ( n4636 , R_c3ee_102f6848 );
buf ( n4637 , R_13b12_13a1a728 );
buf ( n4638 , R_10a0c_11cdf1c8 );
buf ( n4639 , R_13974_13a19008 );
buf ( n4640 , R_13602_126635a8 );
buf ( n4641 , R_124e1_11cdb668 );
buf ( n4642 , R_142d7_12b30d58 );
buf ( n4643 , R_14960_105b5598 );
buf ( n4644 , R_f86d_120385f8 );
buf ( n4645 , R_148a0_12b38ab8 );
buf ( n4646 , R_e63f_f8cb9f8 );
buf ( n4647 , R_12741_105642d8 );
buf ( n4648 , R_684e_1056aa98 );
buf ( n4649 , R_13b04_12081558 );
buf ( n4650 , R_1453f_11ce2328 );
buf ( n4651 , R_148b5_1207f898 );
buf ( n4652 , R_1499c_12080658 );
buf ( n4653 , R_128e2_12647668 );
buf ( n4654 , R_13345_11ce0988 );
buf ( n4655 , R_cd4f_102f2f68 );
buf ( n4656 , R_13dd3_1204cd38 );
buf ( n4657 , R_13ea4_11ce0708 );
buf ( n4658 , R_f16b_11cda448 );
buf ( n4659 , R_139fe_1153e5b8 );
buf ( n4660 , R_12eed_102ee1e8 );
buf ( n4661 , R_13479_13306b28 );
buf ( n4662 , R_1135b_1056d158 );
buf ( n4663 , R_131a5_1153dc58 );
buf ( n4664 , R_14744_1264b3a8 );
buf ( n4665 , R_144c6_1056d5b8 );
buf ( n4666 , R_13109_f8c4798 );
buf ( n4667 , R_137bb_10564058 );
buf ( n4668 , R_146db_1056a818 );
buf ( n4669 , R_119c2_13a1a548 );
buf ( n4670 , R_eb5e_1056d018 );
buf ( n4671 , R_b0d7_1153e3d8 );
buf ( n4672 , R_13b9e_12083038 );
buf ( n4673 , R_1116a_13a15868 );
buf ( n4674 , R_12a65_10564c38 );
buf ( n4675 , R_14969_11cdb2a8 );
buf ( n4676 , R_1464d_12075618 );
buf ( n4677 , R_e3c5_12080a18 );
buf ( n4678 , R_1469c_120511f8 );
buf ( n4679 , R_d50f_12663828 );
buf ( n4680 , R_137f0_12079358 );
buf ( n4681 , R_11593_1207a258 );
buf ( n4682 , R_14350_1207d8b8 );
buf ( n4683 , R_cbe2_11536a98 );
buf ( n4684 , R_110ed_10563d38 );
buf ( n4685 , R_1125d_102f86e8 );
buf ( n4686 , R_13c09_11ce4268 );
buf ( n4687 , R_135fc_13795948 );
buf ( n4688 , R_14557_11cdcec8 );
buf ( n4689 , R_112_13312248 );
buf ( n4690 , R_1fd_133221a8 );
buf ( n4691 , R_9e_11539838 );
buf ( n4692 , R_143b2_11cddd28 );
buf ( n4693 , R_12fec_102efea8 );
buf ( n4694 , R_c4d7_13a1f408 );
buf ( n4695 , R_1398e_13320bc8 );
buf ( n4696 , R_12894_11ce1428 );
buf ( n4697 , R_b6f4_102f9ea8 );
buf ( n4698 , R_fcb3_12649be8 );
buf ( n4699 , R_12375_1207edf8 );
buf ( n4700 , R_146b1_102ed248 );
buf ( n4701 , R_11b11_11545818 );
buf ( n4702 , R_58_13317a28 );
buf ( n4703 , R_73_12b3e0f8 );
buf ( n4704 , R_bd7c_11ce2be8 );
buf ( n4705 , R_12fd8_10565278 );
buf ( n4706 , R_14876_12054678 );
buf ( n4707 , R_138da_1153dbb8 );
buf ( n4708 , R_14825_12647168 );
buf ( n4709 , R_14a4d_12646ee8 );
buf ( n4710 , R_124_1203edb8 );
buf ( n4711 , R_15a_f8c6958 );
buf ( n4712 , R_1b5_1331afe8 );
buf ( n4713 , R_1eb_12038d78 );
buf ( n4714 , R_1475d_11546038 );
buf ( n4715 , R_171_105aa5f8 );
buf ( n4716 , R_106ea_102f6528 );
buf ( n4717 , R_19e_1331e788 );
buf ( n4718 , R_11a86_1204ffd8 );
buf ( n4719 , R_fad7_102f5ee8 );
buf ( n4720 , R_e21e_1056b7b8 );
buf ( n4721 , R_12933_11cd7c48 );
buf ( n4722 , R_6c_12040938 );
buf ( n4723 , R_99_12b27618 );
buf ( n4724 , R_1353d_1153d9d8 );
buf ( n4725 , R_b283_1330acc8 );
buf ( n4726 , R_143ae_13a1cca8 );
buf ( n4727 , R_14801_11540c78 );
buf ( n4728 , R_149e7_10568298 );
buf ( n4729 , R_14708_1203c018 );
buf ( n4730 , R_14450_13a17028 );
buf ( n4731 , R_128_12b43b98 );
buf ( n4732 , R_145_1265aa48 );
buf ( n4733 , R_1ca_1265ff48 );
buf ( n4734 , R_1e7_12b3d798 );
buf ( n4735 , R_7741_13a16128 );
buf ( n4736 , R_da39_12b40718 );
buf ( n4737 , R_e38d_12651168 );
buf ( n4738 , R_12fc4_11544878 );
buf ( n4739 , R_145e7_11544058 );
buf ( n4740 , R_1465f_105676b8 );
buf ( n4741 , R_10fc1_12078638 );
buf ( n4742 , R_704f_11ce4da8 );
buf ( n4743 , R_13a8d_13318108 );
buf ( n4744 , R_145c3_1264da68 );
buf ( n4745 , R_faad_13a1fd68 );
buf ( n4746 , R_12738_10570678 );
buf ( n4747 , R_11935_13a1ff48 );
buf ( n4748 , R_11720_1330eaa8 );
buf ( n4749 , R_d16a_11ce5de8 );
buf ( n4750 , R_13e0d_13a1b4e8 );
buf ( n4751 , R_1447d_11ce3a48 );
buf ( n4752 , R_152_12b3c4d8 );
buf ( n4753 , R_105ba_13306bc8 );
buf ( n4754 , R_b1aa_12649468 );
buf ( n4755 , R_1bd_12653be8 );
buf ( n4756 , R_14a50_13a161c8 );
buf ( n4757 , R_13a83_10567a78 );
buf ( n4758 , R_123c2_13797108 );
buf ( n4759 , R_144b7_13305d68 );
buf ( n4760 , R_13814_137926a8 );
buf ( n4761 , R_12cbd_13a14328 );
buf ( n4762 , R_11bab_120768d8 );
buf ( n4763 , R_c07e_13a18b08 );
buf ( n4764 , R_142f9_11545e58 );
buf ( n4765 , R_1478a_12652928 );
buf ( n4766 , R_14a3b_11ce2d28 );
buf ( n4767 , R_c3a2_13a19508 );
buf ( n4768 , R_aa_126535a8 );
buf ( n4769 , R_146e7_10566538 );
buf ( n4770 , R_138fb_12082778 );
buf ( n4771 , R_13988_133186a8 );
buf ( n4772 , R_13c43_1264cca8 );
buf ( n4773 , R_14590_132f3b08 );
buf ( n4774 , R_110cf_137940e8 );
buf ( n4775 , R_13326_12648d88 );
buf ( n4776 , R_13153_10567118 );
buf ( n4777 , R_1405e_f8c95b8 );
buf ( n4778 , R_1051f_13793b48 );
buf ( n4779 , R_f518_12075bb8 );
buf ( n4780 , R_143a2_12079038 );
buf ( n4781 , R_147a8_12657de8 );
buf ( n4782 , R_13cb3_102f6fc8 );
buf ( n4783 , R_10c3d_f8c5b98 );
buf ( n4784 , R_e7ab_1264f7c8 );
buf ( n4785 , R_13449_12077378 );
buf ( n4786 , R_14403_12b29418 );
buf ( n4787 , R_148b2_132fc708 );
buf ( n4788 , R_1468f_10562cf8 );
buf ( n4789 , R_f7_13309828 );
buf ( n4790 , R_13f54_102f4e08 );
buf ( n4791 , R_218_12050258 );
buf ( n4792 , R_83_1379cd88 );
buf ( n4793 , R_12f16_137a0b68 );
buf ( n4794 , R_10598_102ead68 );
buf ( n4795 , R_10365_12051478 );
buf ( n4796 , R_13ab4_13a12ca8 );
buf ( n4797 , R_13393_10568a18 );
buf ( n4798 , R_13683_1207cf58 );
buf ( n4799 , R_13a_105ac2b8 );
buf ( n4800 , R_127d5_11cdf268 );
buf ( n4801 , R_11917_11ce1248 );
buf ( n4802 , R_1d5_1265e468 );
buf ( n4803 , R_12e98_1204e778 );
buf ( n4804 , R_b3_12655ea8 );
buf ( n4805 , R_149cc_10564cd8 );
buf ( n4806 , R_134d9_10565f98 );
buf ( n4807 , R_fd0b_102ec488 );
buf ( n4808 , R_af25_133136a8 );
buf ( n4809 , R_11948_12b288d8 );
buf ( n4810 , R_149c6_1207b018 );
buf ( n4811 , R_14b_12b28a18 );
buf ( n4812 , R_1c4_12652e28 );
buf ( n4813 , R_10199_13a1f368 );
buf ( n4814 , R_80_12055438 );
buf ( n4815 , R_10b70_f8cd438 );
buf ( n4816 , R_10cdf_115401d8 );
buf ( n4817 , R_11a66_1207dc78 );
buf ( n4818 , R_132fc_13307708 );
buf ( n4819 , R_8c7b_12076b58 );
buf ( n4820 , R_1495a_1207a2f8 );
buf ( n4821 , R_1201a_10570218 );
buf ( n4822 , R_132d6_11ce0348 );
buf ( n4823 , R_14963_13304be8 );
buf ( n4824 , R_1285e_11545c78 );
buf ( n4825 , R_130de_102f58a8 );
buf ( n4826 , R_fb5f_13a1e288 );
buf ( n4827 , R_13ecf_1207c5f8 );
buf ( n4828 , R_1456f_13a1f5e8 );
buf ( n4829 , R_ea_1331a9a8 );
buf ( n4830 , R_120_12b400d8 );
buf ( n4831 , R_13eac_11ce2a08 );
buf ( n4832 , R_12568_1056b0d8 );
buf ( n4833 , R_e3ba_1207df98 );
buf ( n4834 , R_dcf2_12085298 );
buf ( n4835 , R_1ef_f8c2cb8 );
buf ( n4836 , R_225_12b3a318 );
buf ( n4837 , R_f7da_1204e9f8 );
buf ( n4838 , R_f857_13a13748 );
buf ( n4839 , R_1461a_13301988 );
buf ( n4840 , R_146b7_13a15228 );
buf ( n4841 , R_1384a_126503a8 );
buf ( n4842 , R_c8e7_105b6498 );
buf ( n4843 , R_86_137a1a68 );
buf ( n4844 , R_a3_126621a8 );
buf ( n4845 , R_f862_13a1a908 );
buf ( n4846 , R_10ab7_102f7b08 );
buf ( n4847 , R_11890_102eb308 );
buf ( n4848 , R_df3c_120774b8 );
buf ( n4849 , R_1369b_1330c2a8 );
buf ( n4850 , R_12e03_132ff368 );
buf ( n4851 , R_1356b_102f5da8 );
buf ( n4852 , R_10e42_1207e718 );
buf ( n4853 , R_10f59_f8c2c18 );
buf ( n4854 , R_127b6_12b412f8 );
buf ( n4855 , R_120e7_12b44818 );
buf ( n4856 , R_12492_1265b9e8 );
buf ( n4857 , R_10d12_13792b08 );
buf ( n4858 , R_130ae_12044b78 );
buf ( n4859 , R_13652_11ce1ce8 );
buf ( n4860 , R_117a7_12080fb8 );
buf ( n4861 , R_14674_13a13ba8 );
buf ( n4862 , R_11306_11540638 );
buf ( n4863 , R_d5_126617a8 );
buf ( n4864 , R_de_1265ce88 );
buf ( n4865 , R_12c_1379b488 );
buf ( n4866 , R_135_f8c6f98 );
buf ( n4867 , R_1da_12664b88 );
buf ( n4868 , R_1e3_1153c498 );
buf ( n4869 , R_122dd_13a1b6c8 );
buf ( n4870 , R_231_1379a6c8 );
buf ( n4871 , R_23a_12660b28 );
buf ( n4872 , R_1240e_13a150e8 );
buf ( n4873 , R_14686_13a137e8 );
buf ( n4874 , R_146c6_f8cf918 );
buf ( n4875 , R_13f5b_1207c738 );
buf ( n4876 , R_ebb7_102efd68 );
buf ( n4877 , R_1447a_105697d8 );
buf ( n4878 , R_13c95_12650ee8 );
buf ( n4879 , R_11de0_12083cb8 );
buf ( n4880 , R_11552_12648c48 );
buf ( n4881 , R_11cb2_1207ab18 );
buf ( n4882 , R_14849_11ce0028 );
buf ( n4883 , R_13f45_13a134c8 );
buf ( n4884 , R_13726_12084f78 );
buf ( n4885 , R_121f2_102f30a8 );
buf ( n4886 , R_ef_1379b0c8 );
buf ( n4887 , R_163_12b38a18 );
buf ( n4888 , R_1ac_12b29558 );
buf ( n4889 , R_220_12b25638 );
buf ( n4890 , R_14623_13a12a28 );
buf ( n4891 , R_1393a_11ce3408 );
buf ( n4892 , R_139ea_11cd8828 );
buf ( n4893 , R_cf49_11541718 );
buf ( n4894 , R_b889_1056a458 );
buf ( n4895 , R_1349f_1204fdf8 );
buf ( n4896 , R_170_120440d8 );
buf ( n4897 , R_19f_133087e8 );
buf ( n4898 , R_a9d8_102f22e8 );
buf ( n4899 , R_7d_12660308 );
buf ( n4900 , R_1460b_10569a58 );
buf ( n4901 , R_11983_13318568 );
buf ( n4902 , R_a6e4_13314648 );
buf ( n4903 , R_144b1_1207b478 );
buf ( n4904 , R_14614_12664f48 );
buf ( n4905 , R_139d7_132fda68 );
buf ( n4906 , R_ec64_11ce6248 );
buf ( n4907 , R_12d32_115454f8 );
buf ( n4908 , R_82bb_1204a678 );
buf ( n4909 , R_1472c_13a139c8 );
buf ( n4910 , R_144f7_10565e58 );
buf ( n4911 , R_10dad_12082f98 );
buf ( n4912 , R_b05c_1330b4e8 );
buf ( n4913 , R_13ef1_105714d8 );
buf ( n4914 , R_14635_12b3b038 );
buf ( n4915 , R_117b5_1056fdb8 );
buf ( n4916 , R_14692_11cdf128 );
buf ( n4917 , R_13f_1203dd78 );
buf ( n4918 , R_1055c_105672f8 );
buf ( n4919 , R_1d0_12040258 );
buf ( n4920 , R_13aba_1265cde8 );
buf ( n4921 , R_131e1_102f2ec8 );
buf ( n4922 , R_eb07_1153ef18 );
buf ( n4923 , R_9c9a_1056c578 );
buf ( n4924 , R_10605_11545d18 );
buf ( n4925 , R_13a97_12079218 );
buf ( n4926 , R_1331b_102efc28 );
buf ( n4927 , R_14879_11ce58e8 );
buf ( n4928 , R_14996_102eb3a8 );
buf ( n4929 , R_1405c_11ce34a8 );
buf ( n4930 , R_14945_1056e238 );
buf ( n4931 , R_b65f_11cdba28 );
buf ( n4932 , R_13f3e_13a1e508 );
buf ( n4933 , R_dbc0_132fb9e8 );
buf ( n4934 , R_1351c_13797068 );
buf ( n4935 , R_14804_120788b8 );
buf ( n4936 , R_14a0b_133206c8 );
buf ( n4937 , R_89_126595a8 );
buf ( n4938 , R_13c33_11ce3688 );
buf ( n4939 , R_4f_12b44d18 );
buf ( n4940 , R_cb5a_12b256d8 );
buf ( n4941 , R_13b85_10571258 );
buf ( n4942 , R_138f4_1330a9a8 );
buf ( n4943 , R_ee1a_1264fae8 );
buf ( n4944 , R_10411_102f8828 );
buf ( n4945 , R_14331_1056be98 );
buf ( n4946 , R_14717_1153a378 );
buf ( n4947 , R_94_1330ee68 );
buf ( n4948 , R_e5_1153cfd8 );
buf ( n4949 , R_22a_12b43698 );
buf ( n4950 , R_cba1_13a16e48 );
buf ( n4951 , R_129d1_12047978 );
buf ( n4952 , R_143d8_11cdc2e8 );
buf ( n4953 , R_13070_1264b268 );
buf ( n4954 , R_12915_1056d518 );
buf ( n4955 , R_12942_11cdd0a8 );
buf ( n4956 , R_145a8_12662608 );
buf ( n4957 , R_fda2_1264e328 );
buf ( n4958 , R_ee25_13a16588 );
buf ( n4959 , R_13a1f_11cde2c8 );
buf ( n4960 , R_1432d_11cdddc8 );
buf ( n4961 , R_13be3_12036bb8 );
buf ( n4962 , R_fe10_13a14468 );
buf ( n4963 , R_12610_1204bcf8 );
buf ( n4964 , R_13701_11cdc608 );
buf ( n4965 , R_12597_105711b8 );
buf ( n4966 , R_1441d_12035d58 );
buf ( n4967 , R_1443c_137979c8 );
buf ( n4968 , R_139a7_11ce70a8 );
buf ( n4969 , R_13ad3_1056bdf8 );
buf ( n4970 , R_143e0_102efcc8 );
buf ( n4971 , R_147cc_13315ae8 );
buf ( n4972 , R_1444b_11cdad08 );
buf ( n4973 , R_12631_12036c58 );
buf ( n4974 , R_13dda_102f4fe8 );
buf ( n4975 , R_efd_13a14fa8 );
buf ( n4976 , R_14954_12054358 );
buf ( n4977 , R_1287f_115422f8 );
buf ( n4978 , R_1169f_102f8968 );
buf ( n4979 , R_13a2b_1264b628 );
buf ( n4980 , R_11285_102f9e08 );
buf ( n4981 , R_12548_1056ce38 );
buf ( n4982 , R_1173e_12649fa8 );
buf ( n4983 , R_10b51_13a18a68 );
buf ( n4984 , R_148ca_13a18c48 );
buf ( n4985 , R_12c82_102f0448 );
buf ( n4986 , R_13b79_11543d38 );
buf ( n4987 , R_14057_f8cd618 );
buf ( n4988 , R_a2e4_1056c618 );
buf ( n4989 , R_101e6_1330c7a8 );
buf ( n4990 , R_13a56_f8c0a58 );
buf ( n4991 , R_d6bc_13a1ca28 );
buf ( n4992 , R_4a_1265e648 );
buf ( n4993 , R_115_13316c68 );
buf ( n4994 , R_1224c_12b3d478 );
buf ( n4995 , R_1fa_1265d388 );
buf ( n4996 , R_eeda_11cd81e8 );
buf ( n4997 , R_1455d_11cd9fe8 );
buf ( n4998 , R_1402e_1264dc48 );
buf ( n4999 , R_c753_12039098 );
buf ( n5000 , R_1283c_13a1da68 );
buf ( n5001 , R_aeda_13a1d6a8 );
buf ( n5002 , R_14939_1379f448 );
buf ( n5003 , R_14a20_13a13e28 );
buf ( n5004 , R_13a9d_12081698 );
buf ( n5005 , R_117c0_11ce3e08 );
buf ( n5006 , R_114e1_132f28e8 );
buf ( n5007 , R_1476f_132fb768 );
buf ( R_147ef_11ce6748 , n25340 );
buf ( R_5f38_10569f58 , n31580 );
buf ( R_13287_11ce6b08 , n35435 );
buf ( R_c94b_102f7608 , n37731 );
buf ( R_20a_1204ce78 , n37733 );
buf ( R_12f29_10571bb8 , n39770 );
buf ( R_13a43_13a1dec8 , n41948 );
buf ( R_1474d_1056fbd8 , n41954 );
buf ( R_14493_12657988 , n41960 );
buf ( R_11fd1_11ce17e8 , n43523 );
buf ( R_14705_1264d248 , n43529 );
buf ( R_105_f8cc2b8 , n221291 );
buf ( R_13cb9_11ce3c28 , n44777 );
buf ( R_138ee_13309fa8 , n223848 );
buf ( R_129dc_11543018 , n47179 );
buf ( R_10bcf_11ce1ba8 , n48254 );
buf ( R_13b6e_13a1e648 , n226818 );
buf ( R_14840_13a13ec8 , n49065 );
buf ( R_13482_10563838 , n49964 );
buf ( R_12d08_12650088 , n228379 );
buf ( R_10303_12b42dd8 , n229122 );
buf ( R_1437c_1056ac78 , n229140 );
buf ( R_87e9_1056cd98 , n52240 );
buf ( R_a30d_13320588 , n53008 );
buf ( R_144a2_133222e8 , n53014 );
buf ( R_1236b_13a1c8e8 , n53686 );
buf ( R_1396e_105627f8 , n54207 );
buf ( R_9ba7_10567258 , n54337 );
buf ( R_1f3_13797a68 , n54338 );
buf ( R_11c_13796528 , n54339 );
buf ( R_7a_1331e148 , n232101 );
buf ( R_117c9_1264ba88 , n55113 );
buf ( R_13b3f_1153ed38 , n55157 );
buf ( R_11abc_1264c2a8 , n55743 );
buf ( R_20d_137962a8 , n55744 );
buf ( R_207_1265a548 , n55745 );
buf ( R_14828_1207a118 , n233513 );
buf ( R_148eb_105aa7d8 , n233519 );
buf ( R_f3a4_10568bf8 , n233844 );
buf ( R_1b6_13799d68 , n233845 );
buf ( R_13429_1207f4d8 , n234027 );
buf ( R_14506_1056e878 , n234033 );
buf ( R_159_12b3d158 , n234034 );
buf ( R_108_105aaeb8 , n234035 );
buf ( R_102_13794cc8 , n234037 );
buf ( R_b1_12053638 , n234038 );
buf ( R_54_13309d28 , n234039 );
buf ( R_145d8_12b3ae58 , n234045 );
buf ( R_1278a_12083718 , n234319 );
buf ( R_13640_11cdeae8 , n234451 );
buf ( R_f706_11542578 , n234821 );
buf ( R_dc82_1153ebf8 , n235055 );
buf ( R_1491b_1265ef08 , n235061 );
buf ( R_14a05_10569738 , n235067 );
buf ( R_13fc5_102eac28 , n235737 );
buf ( R_1405a_115415d8 , n235740 );
buf ( R_136b3_126461c8 , n235900 );
buf ( R_1a0_132f9c88 , n235901 );
buf ( R_16f_1265bee8 , n235902 );
buf ( R_1480d_105a9dd8 , n235908 );
buf ( R_61_13304288 , n235909 );
buf ( R_e082_13798fa8 , n236516 );
buf ( R_10c7d_12082bd8 , n236801 );
buf ( R_14793_1379e188 , n236807 );
buf ( R_11ee1_102f4688 , n237364 );
buf ( R_128ba_12b27758 , n237717 );
buf ( R_70_120513d8 , n237718 );
buf ( R_129f0_12049bd8 , n237884 );
buf ( R_117e7_102f5588 , n238117 );
buf ( R_fee6_13309e68 , n238226 );
buf ( R_148f7_132f3ce8 , n238232 );
buf ( R_1362d_11ce39a8 , n238641 );
buf ( R_10693_126510c8 , n239243 );
buf ( R_11998_12656808 , n239792 );
buf ( R_143ec_11537df8 , n239798 );
buf ( R_138e8_1264afe8 , n240085 );
buf ( R_12650_12649b48 , n240532 );
buf ( R_137a1_105b63f8 , n241071 );
buf ( R_13afd_120772d8 , n241381 );
buf ( R_1490c_1264a7c8 , n241387 );
buf ( R_105e5_13306f88 , n241690 );
buf ( R_12e2b_132fa868 , n241979 );
buf ( R_144e7_12b38e78 , n241985 );
buf ( R_143e4_11cddf08 , n241990 );
buf ( R_1324a_1264c348 , n242093 );
buf ( R_1215a_11542ed8 , n242396 );
buf ( R_f685_11541678 , n242602 );
buf ( R_149ba_102ecb68 , n242608 );
buf ( R_135dc_12646088 , n242876 );
buf ( R_1476c_11cd7928 , n242882 );
buf ( R_146bd_11537998 , n242888 );
buf ( R_1df_12b39378 , n242889 );
buf ( R_13ee8_133069e8 , n243211 );
buf ( R_130_1265ac28 , n243212 );
buf ( R_65_12047c98 , n243213 );
buf ( R_13d75_1330d6a8 , n243273 );
buf ( R_13933_12081198 , n243443 );
buf ( R_133b5_12648388 , n243675 );
buf ( R_125a0_13311488 , n244070 );
buf ( R_8c_1379a808 , n244071 );
buf ( R_eadc_1207ead8 , n244220 );
buf ( R_134c7_126487e8 , n244404 );
buf ( R_11df5_1056e9b8 , n244487 );
buf ( R_144d5_102f8aa8 , n244493 );
buf ( R_12b2a_102eed28 , n244604 );
buf ( R_143d2_11538898 , n244615 );
buf ( R_1462c_102f8508 , n244620 );
buf ( R_13269_11543658 , n244792 );
buf ( R_f4_1331e0a8 , n244793 );
buf ( R_d7_132fde28 , n244794 );
buf ( R_238_1204ec78 , n244795 );
buf ( R_21b_1265e508 , n244796 );
buf ( R_12f3d_12b38b58 , n244843 );
buf ( R_112f1_1153c858 , n244990 );
buf ( R_f09_f8c93d8 , n244993 );
buf ( R_1487c_11cd99a8 , n244999 );
buf ( R_c08f_1207cb98 , n245224 );
buf ( R_923a_13a1ab88 , n245417 );
buf ( R_14042_102f2108 , n245693 );
buf ( R_143e8_102f3b48 , n245699 );
buf ( R_c2e7_13a19e68 , n245941 );
buf ( R_c175_12045118 , n246094 );
buf ( R_1450f_102f8b48 , n246100 );
buf ( R_12b14_12077238 , n246220 );
buf ( R_149e4_13a1c528 , n246226 );
buf ( R_12a04_11ce2968 , n246463 );
buf ( R_145ed_13a14e68 , n246469 );
buf ( R_13884_13796488 , n246685 );
buf ( R_13b0b_1330a688 , n246902 );
buf ( R_b5a4_102f4868 , n247222 );
buf ( R_14584_1056ec38 , n247228 );
buf ( R_13cee_12653148 , n247281 );
buf ( R_10bed_12080ab8 , n247426 );
buf ( R_117f0_102ef4a8 , n247588 );
buf ( R_10a2a_133048c8 , n247747 );
buf ( R_1be_137995e8 , n247748 );
buf ( R_151_12b448b8 , n247749 );
buf ( R_ef06_10563c98 , n247885 );
buf ( R_f9d4_1056b178 , n248088 );
buf ( R_e88a_13a13a68 , n248294 );
buf ( R_13c67_102f38c8 , n248492 );
buf ( R_128eb_10568dd8 , n248775 );
buf ( R_12eaf_f8c3118 , n248821 );
buf ( R_204_12039778 , n248822 );
buf ( R_14951_1265ebe8 , n248828 );
buf ( R_149c3_11ce5348 , n248834 );
buf ( R_1ad_12b28e78 , n248835 );
buf ( R_13f99_102f0da8 , n248998 );
buf ( R_162_12b25e58 , n248999 );
buf ( R_12003_11cdf628 , n249035 );
buf ( R_10b_11539478 , n249036 );
buf ( R_ff_1203c6f8 , n249037 );
buf ( R_1484f_1153ea18 , n249043 );
buf ( R_a8_12b425b8 , n249044 );
buf ( R_5d_13312068 , n249045 );
buf ( R_210_12043bd8 , n249046 );
buf ( R_13d84_102f4188 , n249122 );
buf ( R_142e1_10568658 , n249134 );
buf ( R_10f30_11cd9ae8 , n249223 );
buf ( R_1293d_12b43d78 , n249410 );
buf ( R_10b34_1056da18 , n249514 );
buf ( R_11a07_102eb4e8 , n249625 );
buf ( R_145b1_12082db8 , n249631 );
buf ( R_12c96_13a190a8 , n249782 );
buf ( R_d3b0_10565958 , n249875 );
buf ( R_13f2c_102f4b88 , n249979 );
buf ( R_fb8a_13a18608 , n250071 );
buf ( R_130d5_13319c88 , n250246 );
buf ( R_13f89_102f36e8 , n250286 );
buf ( R_146ff_13a1a4a8 , n250292 );
buf ( R_10ccb_1264f868 , n250388 );
buf ( R_124c3_1056f138 , n250436 );
buf ( R_10786_102f2568 , n250604 );
buf ( R_12a16_10568e78 , n250735 );
buf ( R_10726_102ef408 , n250837 );
buf ( R_137d3_12656da8 , n250919 );
buf ( R_13863_11cddb48 , n250974 );
buf ( R_14993_102f27e8 , n250980 );
buf ( R_bab1_1264a2c8 , n251101 );
buf ( R_1451e_10565818 , n251107 );
buf ( R_12a46_126515c8 , n251195 );
buf ( R_e7da_102f3508 , n251246 );
buf ( R_12756_13a1f0e8 , n251366 );
buf ( R_c4_13797ba8 , n251367 );
buf ( R_128da_1207ec18 , n251468 );
buf ( R_c282_12076838 , n251501 );
buf ( R_1272e_1056cbb8 , n251560 );
buf ( R_14a5f_120797b8 , n251564 );
buf ( R_14448_12663648 , n251570 );
buf ( R_c2_12048058 , n251571 );
buf ( R_1372d_11ce2aa8 , n251715 );
buf ( R_f878_1207c7d8 , n251761 );
buf ( R_13a76_13797888 , n251867 );
buf ( R_13a17_13796b68 , n251914 );
buf ( R_1cb_12044ad8 , n251915 );
buf ( R_14462_12b3f8b8 , n251921 );
buf ( R_6021_1379bd48 , n252075 );
buf ( R_144_13795128 , n252076 );
buf ( R_1383e_105671b8 , n252205 );
buf ( R_147ab_1056a6d8 , n252211 );
buf ( R_c6_1330e0a8 , n252212 );
buf ( R_249_12654368 , n252214 );
buf ( R_1305a_13796ca8 , n252269 );
buf ( R_12e4b_13307348 , n252363 );
buf ( R_14a38_137a1e28 , n252369 );
buf ( R_d1de_11cd9ea8 , n252474 );
buf ( R_138e2_11cd83c8 , n252585 );
buf ( R_13e62_1056dab8 , n252668 );
buf ( R_114a7_1331d748 , n252714 );
buf ( R_12f53_13319648 , n252759 );
buf ( R_f8a4_11543a18 , n252862 );
buf ( R_11ec3_13a157c8 , n252949 );
buf ( R_12c06_11cdac68 , n253092 );
buf ( R_12be8_12649788 , n253128 );
buf ( R_136c6_11cdc6a8 , n253218 );
buf ( R_1482e_13a1a228 , n253224 );
buf ( R_10ba7_115431f8 , n253316 );
buf ( R_89f2_11545098 , n253361 );
buf ( R_11953_1153c538 , n253405 );
buf ( R_9e64_11ce48a8 , n253489 );
buf ( R_e77d_11ce3ea8 , n253547 );
buf ( R_1091c_13a1a2c8 , n253601 );
buf ( R_114ec_12650628 , n253703 );
buf ( R_1286a_11cdcd88 , n253760 );
buf ( R_10d6d_1265db08 , n253888 );
buf ( R_1228f_1331f0e8 , n253909 );
buf ( R_1c5_126590a8 , n253910 );
buf ( R_14490_132f7d48 , n253915 );
buf ( R_1a1_1264a408 , n253916 );
buf ( R_976e_12056398 , n253965 );
buf ( R_6845_12648ec8 , n253998 );
buf ( R_16e_1379a3a8 , n253999 );
buf ( R_14a_12657528 , n254000 );
buf ( R_12718_10566fd8 , n254045 );
buf ( R_145c9_12075438 , n254051 );
buf ( R_c0_132fa5e8 , n254052 );
buf ( R_9c_12655f48 , n254053 );
buf ( R_d230_102edec8 , n254108 );
buf ( R_69_12658888 , n254109 );
buf ( R_13097_11ce5b68 , n254139 );
buf ( R_11051_1264a5e8 , n254184 );
buf ( R_145f0_11536818 , n254190 );
buf ( R_13ccd_132f9288 , n254211 );
buf ( R_e0_12661ac8 , n254212 );
buf ( R_22f_1331df68 , n254213 );
buf ( R_12a2a_11cd9f48 , n254260 );
buf ( R_10a54_11540458 , n254366 );
buf ( R_d027_13795628 , n254415 );
buf ( R_144d2_105677f8 , n254421 );
buf ( R_14638_11cd9228 , n254427 );
buf ( R_1454b_10568338 , n254433 );
buf ( R_147fe_1265bb28 , n254439 );
buf ( R_e861_12650448 , n254473 );
buf ( R_c03c_137931e8 , n254518 );
buf ( R_13574_102f97c8 , n254623 );
buf ( R_10e6d_102ec0c8 , n254671 );
buf ( R_c8_1331c348 , n254672 );
buf ( R_247_12b3bad8 , n254673 );
buf ( R_77_126636e8 , n254674 );
buf ( R_13a50_1056bb78 , n254745 );
buf ( R_129a5_11543798 , n254801 );
buf ( R_ef35_102f6d48 , n254885 );
buf ( R_1028c_137951c8 , n254932 );
buf ( R_1348b_12051838 , n254998 );
buf ( R_11f8b_11cdc428 , n255019 );
buf ( R_1452d_f8c5878 , n255025 );
buf ( R_12a3b_12650308 , n255056 );
buf ( R_13fd5_12079d58 , n255114 );
buf ( R_dd89_13302de8 , n255138 );
buf ( R_13dcc_102f7ec8 , n255188 );
buf ( R_14822_102f5768 , n255194 );
buf ( R_baf1_12084e38 , n255239 );
buf ( R_1315c_11ce75a8 , n255283 );
buf ( R_df0e_12654d68 , n255334 );
buf ( R_efea_11cdc248 , n255377 );
buf ( R_fe90_13a14a08 , n255475 );
buf ( R_1453c_102ec208 , n255480 );
buf ( R_aaa7_102edba8 , n255536 );
buf ( R_13c4e_13a1c988 , n255634 );
buf ( R_f758_13a13d88 , n255656 );
buf ( R_1485e_12b38f18 , n255662 );
buf ( R_ece9_1264c488 , n255710 );
buf ( R_14a35_12037f18 , n255716 );
buf ( R_1190c_102ecfc8 , n255901 );
buf ( R_12810_12650d08 , n255945 );
buf ( R_f016_12044df8 , n255970 );
buf ( R_1494e_13a14f08 , n255975 );
buf ( R_14344_1264eaa8 , n255982 );
buf ( R_10e_1265af48 , n255983 );
buf ( R_13f62_12075758 , n256034 );
buf ( R_fc_133201c8 , n256035 );
buf ( R_1378e_11cdd8c8 , n256054 );
buf ( R_147eb_120847f8 , n256060 );
buf ( R_13331_13308ec8 , n256083 );
buf ( R_213_12654f48 , n256084 );
buf ( R_146ae_1265dc48 , n256090 );
buf ( R_201_1153b138 , n256091 );
buf ( R_11d47_f8cc0d8 , n256115 );
buf ( R_c820_13a19328 , n256167 );
buf ( R_edbe_132fbd08 , n256217 );
buf ( R_be_132f4148 , n256218 );
buf ( R_a1_12043c78 , n256219 );
buf ( R_131b9_102f29c8 , n256262 );
buf ( R_12eb9_1153f738 , n256295 );
buf ( R_146e1_1153fb98 , n256301 );
buf ( R_1487f_13a173e8 , n256307 );
buf ( R_13fb4_11544af8 , n256328 );
buf ( R_1446b_10568798 , n256332 );
buf ( R_ef60_1264cf28 , n256379 );
buf ( R_1463b_1207bd38 , n256385 );
buf ( R_13166_1153aff8 , n256407 );
buf ( R_10a4b_10565bd8 , n256418 );
buf ( R_14599_12080c98 , n256424 );
buf ( R_10b18_12080018 , n256469 );
buf ( R_7254_12055078 , n256516 );
buf ( R_db04_1207b3d8 , n256561 );
buf ( R_149f9_10570cb8 , n256567 );
buf ( R_14a4a_1265d608 , n256573 );
buf ( R_14796_1264b808 , n256579 );
buf ( R_120d3_1379f3a8 , n256595 );
buf ( R_119cb_102f2068 , n256639 );
buf ( R_12acb_10565458 , n256676 );
buf ( R_145b4_12083358 , n256682 );
buf ( R_11ae9_12651528 , n256732 );
buf ( R_13af6_f8ce6f8 , n256788 );
buf ( R_13451_102f0128 , n256818 );
buf ( R_ef8c_1204e098 , n256918 );
buf ( R_ca_12b3e058 , n256919 );
buf ( R_245_f8c5ff8 , n256920 );
buf ( R_af_12b2a8b8 , n256921 );
buf ( R_10e57_11544eb8 , n256945 );
buf ( R_b243_f8c5698 , n256990 );
buf ( R_13633_13a13248 , n257031 );
buf ( R_11c97_10562078 , n257076 );
buf ( R_13838_102f5e48 , n257103 );
buf ( R_efb7_13a1bc68 , n257139 );
buf ( R_d4db_10566038 , n257177 );
buf ( R_10bc8_11ce66a8 , n257225 );
buf ( R_c9c0_102eee68 , n257252 );
buf ( R_13608_10563798 , n257294 );
buf ( R_8f_12b299b8 , n257295 );
buf ( R_59_133089c8 , n257296 );
buf ( R_134f1_102ebf88 , n257321 );
buf ( R_10499_1331e828 , n257344 );
buf ( R_14424_102f8f08 , n257355 );
buf ( R_1d6_133209e8 , n257356 );
buf ( R_ebe2_13a18568 , n257403 );
buf ( R_139_12b44ef8 , n257404 );
buf ( R_97_13792c48 , n257405 );
buf ( R_144ed_105660d8 , n257411 );
buf ( R_120c8_11541d58 , n257443 );
buf ( R_11736_11cde408 , n257467 );
buf ( R_149a8_13317528 , n257472 );
buf ( R_1450c_1056eff8 , n257477 );
buf ( R_147d9_120828b8 , n257482 );
buf ( R_11ea5_1264a9a8 , n257515 );
buf ( R_11425_1207c918 , n257560 );
buf ( R_d53e_1207c2d8 , n257604 );
buf ( R_14787_12b352b8 , n257610 );
buf ( R_13cf3_10571078 , n257650 );
buf ( R_13f36_1330ebe8 , n257674 );
buf ( R_d00d_102ee968 , n257719 );
buf ( R_a1e6_11cde368 , n257767 );
buf ( R_13f77_13a19648 , n257790 );
buf ( R_118_132f5f48 , n257791 );
buf ( R_13688_120832b8 , n257808 );
buf ( R_1f7_105a9978 , n257809 );
buf ( R_f630_1056b858 , n257854 );
buf ( R_136a1_1153fa58 , n257874 );
buf ( R_1b7_126577a8 , n257875 );
buf ( R_158_12b27938 , n257876 );
buf ( R_ec_1330a868 , n257877 );
buf ( R_223_f8c32f8 , n257878 );
buf ( R_133bf_11543338 , n257978 );
buf ( R_f2a8_102f47c8 , n258025 );
buf ( R_e112_12076e78 , n258051 );
buf ( R_12b72_1056c6b8 , n258098 );
buf ( R_2f00_102f3d28 , n258132 );
buf ( R_14819_1331de28 , n258137 );
buf ( R_e809_13313c48 , n258182 );
buf ( R_14358_11cd8788 , n258188 );
buf ( R_1473e_11543b58 , n258194 );
buf ( R_139c7_102ed1a8 , n258216 );
buf ( R_13d65_12036a78 , n258247 );
buf ( R_12c10_102ea548 , n258276 );
buf ( R_13870_11ce5e88 , n258285 );
buf ( R_dede_13a16448 , n258331 );
buf ( R_12c49_12b27438 , n258374 );
buf ( R_1192b_12645e08 , n258417 );
buf ( R_bd66_126533c8 , n258425 );
buf ( R_13fa2_1379f6c8 , n258445 );
buf ( R_13407_1056df18 , n258537 );
buf ( R_118b0_1204acb8 , n258636 );
buf ( R_13c3e_126496e8 , n258652 );
buf ( R_1438a_11cda268 , n258662 );
buf ( R_11e51_102fa268 , n258699 );
buf ( R_102b9_132f6588 , n258746 );
buf ( R_d9_1330dec8 , n258747 );
buf ( R_bc_13799c28 , n258748 );
buf ( R_236_13795f88 , n258749 );
buf ( R_ffee_1264d568 , n258762 );
buf ( R_10ea9_102f8788 , n258784 );
buf ( R_14852_13a154a8 , n258790 );
buf ( R_e696_11cdce28 , n258833 );
buf ( R_1ae_1203c3d8 , n258834 );
buf ( R_1457e_133027e8 , n258838 );
buf ( R_161_12656c68 , n258839 );
buf ( R_127_12b3cc58 , n258840 );
buf ( R_ea26_1265a4a8 , n258883 );
buf ( R_1e8_11539298 , n258884 );
buf ( R_139e4_102f59e8 , n258905 );
buf ( R_1477b_1204f218 , n258911 );
buf ( R_1459c_12056a78 , n258917 );
buf ( R_1336e_11545138 , n258952 );
buf ( R_108cd_102f7ce8 , n258998 );
buf ( R_13b4f_13305c28 , n259038 );
buf ( R_1a2_12b423d8 , n259039 );
buf ( R_16d_12664c28 , n259040 );
buf ( R_14656_11ce6ce8 , n259045 );
buf ( R_827e_1207e998 , n259090 );
buf ( R_11ab0_1204a358 , n259134 );
buf ( R_144ab_12b39af8 , n259139 );
buf ( R_144c3_12080338 , n259145 );
buf ( R_12794_102f5b28 , n259184 );
buf ( R_13149_102f7888 , n259240 );
buf ( R_144e4_12b28838 , n259246 );
buf ( R_13e_12660da8 , n259247 );
buf ( R_123_1330d888 , n259248 );
buf ( R_e7_137956c8 , n259249 );
buf ( R_cc_12038918 , n259250 );
buf ( R_137c7_102f79c8 , n259288 );
buf ( R_243_13796d48 , n259289 );
buf ( R_13795_13795588 , n259329 );
buf ( R_228_10570c18 , n259330 );
buf ( R_13f01_1056e2d8 , n259365 );
buf ( R_13d8e_11cd77e8 , n259415 );
buf ( R_1ec_12039ef8 , n259416 );
buf ( R_f175_13a17ca8 , n259428 );
buf ( R_1d1_126540e8 , n259429 );
buf ( R_14409_12b434b8 , n259438 );
buf ( R_138b2_102f06c8 , n259446 );
buf ( R_14653_1207e0d8 , n259451 );
buf ( R_13044_102f7a68 , n259476 );
buf ( R_13133_13a1ae08 , n259520 );
buf ( R_10b8f_1265ad68 , n259568 );
buf ( R_12e35_12b3b858 , n259618 );
buf ( R_12df0_12050bb8 , n259631 );
buf ( R_fc88_1207be78 , n259654 );
buf ( R_13804_102ef548 , n259682 );
buf ( R_13b68_137a1ba8 , n259712 );
buf ( R_134_13312b68 , n259713 );
buf ( R_14990_1331ae08 , n259719 );
buf ( R_1db_12043db8 , n259720 );
buf ( R_ccdc_102f6488 , n259765 );
buf ( R_1494b_11ce61a8 , n259771 );
buf ( R_12c39_10562ed8 , n259795 );
buf ( R_131c2_11ce4b28 , n259806 );
buf ( R_12d97_126626a8 , n259836 );
buf ( R_12d59_12b26b78 , n259881 );
buf ( R_1352d_13315188 , n259921 );
buf ( R_12c4f_13321d48 , n259948 );
buf ( R_1343e_10562d98 , n259991 );
buf ( R_1345b_102fa088 , n260034 );
buf ( R_1167d_115410d8 , n260075 );
buf ( R_14008_1264dec8 , n260147 );
buf ( R_11bc8_11544e18 , n260169 );
buf ( R_13c9a_1207e178 , n260177 );
buf ( R_148be_12b27f78 , n260183 );
buf ( R_14360_105ad078 , n260188 );
buf ( R_13aa3_12078138 , n260207 );
buf ( R_116da_13a1a7c8 , n260240 );
buf ( R_14732_102f5448 , n260246 );
buf ( R_cec6_132f3608 , n260268 );
buf ( R_133dc_13a1ea08 , n260288 );
buf ( R_14942_f8c5058 , n260293 );
buf ( R_13a0f_10563018 , n260325 );
buf ( R_bd10_f8ce978 , n260332 );
buf ( R_12da1_12647528 , n260362 );
buf ( R_12af5_12052418 , n260415 );
buf ( R_13cf9_13a1c0c8 , n260433 );
buf ( R_13658_12646628 , n260455 );
buf ( R_149bd_1204adf8 , n260460 );
buf ( R_13233_11cde908 , n260484 );
buf ( R_12585_1207a898 , n260572 );
buf ( R_118e9_10564a58 , n260619 );
buf ( R_1359a_13a18928 , n260668 );
buf ( R_12451_13a1d568 , n260700 );
buf ( R_dcbb_1265bf88 , n260724 );
buf ( R_f424_13a1b948 , n260763 );
buf ( R_1226a_11cdef48 , n260786 );
buf ( R_14641_13a12d48 , n260792 );
buf ( R_1257c_11ce4448 , n260839 );
buf ( R_e309_120806f8 , n260864 );
buf ( R_11ccc_13314be8 , n260900 );
buf ( R_146c0_13a15908 , n260905 );
buf ( R_14843_13a196e8 , n260910 );
buf ( R_11d00_1207f9d8 , n260923 );
buf ( R_14a1d_13a14c88 , n260929 );
buf ( R_13d54_11ce00c8 , n260938 );
buf ( R_135b5_132fdd88 , n260979 );
buf ( R_d40b_10569058 , n261012 );
buf ( R_145f9_102ee148 , n261018 );
buf ( R_14882_1056d838 , n261024 );
buf ( R_101a4_f8c2ad8 , n261070 );
buf ( R_13abf_13a15188 , n261088 );
buf ( R_eab3_126509e8 , n261121 );
buf ( R_8296_13322608 , n261167 );
buf ( R_6d_12036618 , n261168 );
buf ( R_50_12b3c118 , n261169 );
buf ( R_11b19_102ee508 , n261211 );
buf ( R_de1d_13a193c8 , n261222 );
buf ( R_14477_11cdcc48 , n261227 );
buf ( R_1195d_12038198 , n261250 );
buf ( R_14527_102eb6c8 , n261256 );
buf ( R_be8c_126504e8 , n261285 );
buf ( R_11e87_12b3c398 , n261333 );
buf ( R_14a02_13309aa8 , n261339 );
buf ( R_12b_1203e6d8 , n261340 );
buf ( R_f1_13799ea8 , n261341 );
buf ( R_21e_126608a8 , n261342 );
buf ( R_1e4_12b28338 , n261343 );
buf ( R_115ff_13304148 , n261376 );
buf ( R_10d8e_1264cfc8 , n261398 );
buf ( R_11500_12083c18 , n261409 );
buf ( R_c4bc_137945e8 , n261447 );
buf ( R_1465c_10568f18 , n261453 );
buf ( R_133e6_11cd9048 , n261497 );
buf ( R_7c4f_11ce4a88 , n261537 );
buf ( R_11f78_12b2c118 , n261588 );
buf ( R_1013a_132f59a8 , n261611 );
buf ( R_149e1_105b62b8 , n261616 );
buf ( R_150_1330cac8 , n261617 );
buf ( R_111_12b3e238 , n261618 );
buf ( R_f9_1204ba78 , n261619 );
buf ( R_ba_1331bc68 , n261620 );
buf ( R_4b_1264c028 , n261621 );
buf ( R_216_1204a038 , n261622 );
buf ( R_13733_f8d0098 , n261641 );
buf ( R_1fe_120539f8 , n261642 );
buf ( R_146de_12648748 , n261647 );
buf ( R_1bf_1265cd48 , n261648 );
buf ( R_74_1331da68 , n261649 );
buf ( R_f5c3_1264d108 , n261681 );
buf ( R_f1f7_120367f8 , n261725 );
buf ( R_e338_13301ac8 , n261747 );
buf ( R_1486d_1056e558 , n261753 );
buf ( R_13e2d_12047fb8 , n261786 );
buf ( R_12344_137a0de8 , n261818 );
buf ( R_14729_10570178 , n261824 );
buf ( R_13364_105717f8 , n261876 );
buf ( R_11160_1153e298 , n261907 );
buf ( R_10a01_11cde228 , n261928 );
buf ( R_13c6f_12041658 , n261956 );
buf ( R_148c4_10568978 , n261961 );
buf ( R_11c81_132f7348 , n262010 );
buf ( R_10ec5_11cdb028 , n262038 );
buf ( R_14441_12659008 , n262046 );
buf ( R_cbab_105a9a18 , n262057 );
buf ( R_1238a_126482e8 , n262090 );
buf ( R_a6_12660448 , n262091 );
buf ( R_12b36_11ce6428 , n262103 );
buf ( R_dc46_10566498 , n262127 );
buf ( R_11f_137936e8 , n262128 );
buf ( R_ce_12055fd8 , n262129 );
buf ( R_241_132fd748 , n262130 );
buf ( R_147f8_1207ccd8 , n262135 );
buf ( R_1f0_13798a08 , n262136 );
buf ( R_1467d_1056bcb8 , n262142 );
buf ( R_14668_11546178 , n262147 );
buf ( R_132cc_1153edd8 , n262190 );
buf ( R_136ba_11ce37c8 , n262210 );
buf ( R_12c23_102f1d48 , n262234 );
buf ( R_106be_1264edc8 , n262257 );
buf ( R_11bde_10564878 , n262279 );
buf ( R_11a1a_11cd9a48 , n262302 );
buf ( R_9548_11ce6ba8 , n262324 );
buf ( R_f451_11542438 , n262347 );
buf ( R_119b7_105663f8 , n262392 );
buf ( R_142e5_102f2388 , n262397 );
buf ( R_147e4_13a19dc8 , n262403 );
buf ( R_d862_12661348 , n262446 );
buf ( R_d940_13a19d28 , n262468 );
buf ( R_eb8c_13a19288 , n262505 );
buf ( R_1175e_11cda088 , n262539 );
buf ( R_146f9_11ce4768 , n262544 );
buf ( R_14551_102eae08 , n262550 );
buf ( R_14578_12b3a6d8 , n262555 );
buf ( R_1467a_13a13568 , n262560 );
buf ( R_1130e_1056bfd8 , n262580 );
buf ( R_1493f_1056d3d8 , n262586 );
buf ( R_14948_102f76a8 , n262592 );
buf ( R_10230_1153d1b8 , n262644 );
buf ( R_f4d1_13a17848 , n262666 );
buf ( R_14772_11cda8a8 , n262672 );
buf ( R_1466e_1203e138 , n262677 );
buf ( R_14999_120382d8 , n262682 );
buf ( R_9d72_102f18e8 , n262724 );
buf ( R_eeaf_10566f38 , n262765 );
buf ( R_13083_12b3ff98 , n262810 );
buf ( R_e288_11541fd8 , n262852 );
buf ( R_13969_102ea408 , n262870 );
buf ( R_13825_1264d928 , n262907 );
buf ( R_134a8_13a13c48 , n262941 );
buf ( R_fcde_115390b8 , n262965 );
buf ( R_14566_102f6988 , n262970 );
buf ( R_f5eb_11544558 , n262991 );
buf ( R_12318_102ec348 , n263031 );
buf ( R_d2c9_11cd9408 , n263074 );
buf ( R_16c_132f7ca8 , n263075 );
buf ( R_d894_1056f778 , n263098 );
buf ( R_12323_102ec8e8 , n263142 );
buf ( R_1a3_13303108 , n263143 );
buf ( R_118ba_13307ac8 , n263165 );
buf ( R_12704_10562938 , n263187 );
buf ( R_148c7_1264d888 , n263193 );
buf ( R_148bb_12661d48 , n263199 );
buf ( R_1221a_13a1d248 , n263248 );
buf ( R_135b0_12651348 , n263257 );
buf ( R_1470e_10562898 , n263263 );
buf ( R_efa_1207d1d8 , n263266 );
buf ( R_ce1e_102f95e8 , n263289 );
buf ( R_126e3_105b5c78 , n263333 );
buf ( R_14026_102ecd48 , n263375 );
buf ( R_11e36_102ed608 , n263398 );
buf ( R_11515_12039318 , n263409 );
buf ( R_108e3_1056dd38 , n263452 );
buf ( R_128f4_1207aa78 , n263462 );
buf ( R_147ae_1207ce18 , n263468 );
buf ( R_12235_12650e48 , n263510 );
buf ( R_12183_12052eb8 , n263543 );
buf ( R_14647_102f04e8 , n263549 );
buf ( R_13aef_11cdd968 , n263578 );
buf ( R_1249f_102f9368 , n263601 );
buf ( R_f34d_13a18ec8 , n263633 );
buf ( R_12c3f_f8cfd78 , n263661 );
buf ( R_13d5d_1153d4d8 , n263705 );
buf ( R_12126_102ef228 , n263727 );
buf ( R_ad_12b3b358 , n263728 );
buf ( R_92_13312d48 , n263729 );
buf ( R_113db_f8cb4f8 , n263764 );
buf ( R_10d98_f8c6318 , n263812 );
buf ( R_1481f_1264dce8 , n263817 );
buf ( R_ad98_102f3aa8 , n263840 );
buf ( R_55_132f50e8 , n263841 );
buf ( R_102d5_f8ced38 , n263871 );
buf ( R_144ae_11545ef8 , n263877 );
buf ( R_a3e0_12655308 , n263892 );
buf ( R_5dbf_13a15f48 , n263914 );
buf ( R_e2_1203f858 , n263915 );
buf ( R_22d_1379de68 , n263916 );
buf ( R_135c4_105b5bd8 , n263955 );
buf ( R_13cff_13a16308 , n263976 );
buf ( R_12692_102eb8a8 , n264001 );
buf ( R_13375_13794a48 , n264043 );
buf ( R_12f6a_10562438 , n264090 );
buf ( R_128c4_102ea5e8 , n264123 );
buf ( R_122f0_12650f88 , n264132 );
buf ( R_14855_12056f78 , n264138 );
buf ( R_14885_13795a88 , n264144 );
buf ( R_bb92_11ce0ca8 , n264152 );
buf ( R_8b04_1265cf28 , n264174 );
buf ( R_e71c_115426b8 , n264218 );
buf ( R_14a23_120545d8 , n264223 );
buf ( R_149_1330f408 , n264224 );
buf ( R_b8_13305048 , n264225 );
buf ( R_1c6_1379cce8 , n264226 );
buf ( R_e13d_102eb448 , n264260 );
buf ( R_14617_11ce2f08 , n264265 );
buf ( R_13557_11545778 , n264286 );
buf ( R_148cd_12082c78 , n264292 );
buf ( R_11768_1264ffe8 , n264302 );
buf ( R_12503_11cdd008 , n264347 );
buf ( R_1239d_1330d1a8 , n264358 );
buf ( R_1448c_105662b8 , n264363 );
buf ( R_160_f8c0d78 , n264364 );
buf ( R_143_13795e48 , n264365 );
buf ( R_1252c_102f1208 , n264398 );
buf ( R_1cc_f8cc858 , n264399 );
buf ( R_149de_11cde7c8 , n264405 );
buf ( R_1af_12b40678 , n264406 );
buf ( R_a28f_11ce5708 , n264437 );
buf ( R_f7ae_11ce57a8 , n264472 );
buf ( R_1243d_10571118 , n264502 );
buf ( R_d0df_126478e8 , n264541 );
buf ( R_1498d_1153fe18 , n264546 );
buf ( R_10350_11cda6c8 , n264579 );
buf ( R_103a6_10569878 , n264591 );
buf ( R_128b0_1056c118 , n264636 );
buf ( R_14936_10561e98 , n264642 );
buf ( R_10d1b_11cd7748 , n264687 );
buf ( R_ed92_102eea08 , n264733 );
buf ( R_145d2_11cdb208 , n264739 );
buf ( R_109f6_1153ca38 , n264762 );
buf ( R_cc46_1207b298 , n264784 );
buf ( R_11006_126501c8 , n264808 );
buf ( R_188_1265c348 , n264809 );
buf ( R_187_12b25d18 , n264810 );
buf ( R_12f_1379dbe8 , n264811 );
buf ( R_db_12663f08 , n264812 );
buf ( R_84_12652ce8 , n264813 );
buf ( R_81_12042a58 , n264814 );
buf ( R_234_12b43af8 , n264815 );
buf ( R_1e0_133037e8 , n264816 );
buf ( R_13ed7_1207ad98 , n264844 );
buf ( R_189_f8c6458 , n264845 );
buf ( R_186_126553a8 , n264846 );
buf ( R_157_132f7a28 , n264847 );
buf ( R_d0_105aa238 , n264848 );
buf ( R_23f_13307848 , n264849 );
buf ( R_11399_12b3c1b8 , n264868 );
buf ( R_1b8_11537358 , n264869 );
buf ( R_f82c_f8cdc58 , n264912 );
buf ( R_d9ca_10562bb8 , n264955 );
buf ( R_145f6_f8c3398 , n264960 );
buf ( R_1449c_11ce71e8 , n264966 );
buf ( R_13850_13a1fe08 , n264987 );
buf ( R_135e3_13306da8 , n265005 );
buf ( R_ec0b_132fa368 , n265017 );
buf ( R_147e0_13a12fc8 , n265023 );
buf ( R_13add_132ff728 , n265061 );
buf ( R_f65b_12084578 , n265084 );
buf ( R_10cb4_11cdf9e8 , n265117 );
buf ( R_18a_133173e8 , n265118 );
buf ( R_185_12042cd8 , n265119 );
buf ( R_134d0_12651028 , n265140 );
buf ( R_144f3_102f3fa8 , n265145 );
buf ( R_12dd1_f8c52d8 , n265156 );
buf ( R_135a9_10567938 , n265199 );
buf ( R_11b39_102ec988 , n265242 );
buf ( R_1386a_102ebda8 , n265251 );
buf ( R_14747_12042b98 , n265257 );
buf ( R_148d0_137a0a28 , n265263 );
buf ( R_11f4d_137986e8 , n265298 );
buf ( R_13d05_12081378 , n265326 );
buf ( R_f56e_102f2608 , n265338 );
buf ( R_62_12b26498 , n265339 );
buf ( R_10e0b_1056abd8 , n265371 );
buf ( R_ba73_1264c8e8 , n265414 );
buf ( R_14888_12653288 , n265420 );
buf ( R_fc34_1379c428 , n265464 );
buf ( R_18b_12663fa8 , n265465 );
buf ( R_184_1153acd8 , n265466 );
buf ( R_119d5_1331dc48 , n265489 );
buf ( R_122b5_13305688 , n265529 );
buf ( R_e051_12649f08 , n265553 );
buf ( R_ca0a_10567438 , n265583 );
buf ( R_10a84_115427f8 , n265604 );
buf ( R_668e_10563f18 , n265611 );
buf ( R_14539_102f7108 , n265616 );
buf ( R_c3d6_11cdb7a8 , n265659 );
buf ( R_11703_132fa728 , n265677 );
buf ( R_1472f_105708f8 , n265682 );
buf ( R_1307a_11cdc1a8 , n265705 );
buf ( R_fdae_1153d258 , n265730 );
buf ( R_13ac5_102ee3c8 , n265759 );
buf ( R_120bd_1153ff58 , n265804 );
buf ( R_13f6e_12649dc8 , n265825 );
buf ( R_1177b_1207fbb8 , n265870 );
buf ( R_f804_1379efe8 , n265893 );
buf ( R_111d5_13a17c08 , n265911 );
buf ( R_14750_13304008 , n265916 );
buf ( R_137d9_12055e98 , n265922 );
buf ( R_87_132ffa48 , n265923 );
buf ( R_7e_137949a8 , n265924 );
buf ( R_f140_1056f598 , n265946 );
buf ( R_d43f_12079678 , n265959 );
buf ( R_11900_1056f6d8 , n266004 );
buf ( R_18c_12660e48 , n266005 );
buf ( R_c969_1330f9a8 , n266036 );
buf ( R_183_126587e8 , n266037 );
buf ( R_11093_102f60c8 , n266060 );
buf ( R_f31e_120770f8 , n266071 );
buf ( R_f06_1265f728 , n266074 );
buf ( R_d5cf_102f5128 , n266120 );
buf ( R_10874_12037838 , n266132 );
buf ( R_11324_13a1f228 , n266144 );
buf ( R_13621_120823b8 , n266179 );
buf ( R_120dd_f8cdcf8 , n266211 );
buf ( R_148d3_12049a98 , n266217 );
buf ( R_13e42_12648888 , n266239 );
buf ( R_144c0_12078db8 , n266245 );
buf ( R_12978_13316d08 , n266267 );
buf ( R_11b5e_13a1b088 , n266300 );
buf ( R_13025_13a1ef08 , n266344 );
buf ( R_e615_12084bb8 , n266357 );
buf ( R_149b7_102ea4a8 , n266363 );
buf ( R_1497e_1207ef38 , n266368 );
buf ( R_11fee_12b2a3b8 , n266408 );
buf ( R_11b_12b43198 , n266409 );
buf ( R_5e_126647c8 , n266410 );
buf ( R_1f4_1265d108 , n266411 );
buf ( R_1445f_13792888 , n266416 );
buf ( R_13981_13798aa8 , n266445 );
buf ( R_14569_11cdbfc8 , n266451 );
buf ( R_114_12b3e4b8 , n266452 );
buf ( R_f6_12664188 , n266453 );
buf ( R_9f_12054d58 , n266454 );
buf ( R_66_13308068 , n266455 );
buf ( R_219_1203c338 , n266456 );
buf ( R_132a5_12654868 , n266490 );
buf ( R_f9aa_11cdd5a8 , n266534 );
buf ( R_1fb_126610c8 , n266535 );
buf ( R_1a4_13798648 , n266536 );
buf ( R_16b_1331a2c8 , n266537 );
buf ( R_9a_12658568 , n266538 );
buf ( R_13c54_102f6e88 , n266580 );
buf ( R_14933_1207e5d8 , n266585 );
buf ( R_a6b7_1264b588 , n266607 );
buf ( R_10fad_13a15548 , n266628 );
buf ( R_18d_13321a28 , n266629 );
buf ( R_182_13315cc8 , n266630 );
buf ( R_14a58_102f65c8 , n266638 );
buf ( R_c8f6_132f4a08 , n266656 );
buf ( R_1458d_13a17ac8 , n266661 );
buf ( R_126d9_11545598 , n266682 );
buf ( R_10942_102f85a8 , n266715 );
buf ( R_14a32_12654ea8 , n266721 );
buf ( R_b7bc_12b28798 , n266752 );
buf ( R_1389f_11cda3a8 , n266768 );
buf ( R_14602_102ed7e8 , n266774 );
buf ( R_100bf_1330b9e8 , n266795 );
buf ( R_112eb_115386b8 , n266806 );
buf ( R_146d5_105b59f8 , n266812 );
buf ( R_1206a_1207c878 , n266823 );
buf ( R_e2de_1264ce88 , n266848 );
buf ( R_13b3a_11cddaa8 , n266867 );
buf ( R_13739_10563bf8 , n266875 );
buf ( R_148d6_11cd86e8 , n266881 );
buf ( R_1319d_11544918 , n266893 );
buf ( R_12f7f_12077eb8 , n266916 );
buf ( R_1242c_f8cda78 , n266936 );
buf ( R_14483_12054fd8 , n266941 );
buf ( R_14456_102ea728 , n266947 );
buf ( R_6b42_120790d8 , n266965 );
buf ( R_1186d_f8cbb38 , n266985 );
buf ( R_147d3_12648e28 , n266991 );
buf ( R_11add_1056c4d8 , n267016 );
buf ( R_13c18_1264df68 , n267053 );
buf ( R_13e19_132f7c08 , n267084 );
buf ( R_b6_1265e148 , n267085 );
buf ( R_13bb8_1265edc8 , n267104 );
buf ( R_146a8_12050118 , n267109 );
buf ( R_18e_12043ef8 , n267110 );
buf ( R_181_12647a28 , n267111 );
buf ( R_b677_12083178 , n267155 );
buf ( R_1176f_1379f8a8 , n267186 );
buf ( R_11d7b_102f2d88 , n267214 );
buf ( R_145bd_1207cff8 , n267219 );
buf ( R_13bae_105700d8 , n267237 );
buf ( R_10fed_1330ad68 , n267260 );
buf ( R_1479f_11cde4a8 , n267265 );
buf ( R_71_1265e8c8 , n267266 );
buf ( R_3ca5_102eebe8 , n267288 );
buf ( R_14769_1056b718 , n267294 );
buf ( R_139ba_11ce35e8 , n267301 );
buf ( R_ccf5_13a128e8 , n267332 );
buf ( R_13964_1207def8 , n267351 );
buf ( R_13920_133128e8 , n267369 );
buf ( R_13b74_11cd8dc8 , n267406 );
buf ( R_13e6d_11cd90e8 , n267418 );
buf ( R_13ae8_11545db8 , n267435 );
buf ( R_e946_13796668 , n267457 );
buf ( R_12db3_10562b18 , n267479 );
buf ( R_7b5f_1264bc68 , n267500 );
buf ( R_139f5_132fc348 , n267546 );
buf ( R_cd6e_10562a78 , n267572 );
buf ( R_13626_12077cd8 , n267599 );
buf ( R_148dc_102f3c88 , n267604 );
buf ( R_11db0_13302748 , n267619 );
buf ( R_1470b_115413f8 , n267624 );
buf ( R_fd8e_120835d8 , n267647 );
buf ( R_142aa_102f2a68 , n267652 );
buf ( R_1267b_1056b538 , n267698 );
buf ( R_10df7_1264ae08 , n267711 );
buf ( R_b753_102ebe48 , n267742 );
buf ( R_14a47_102eeb48 , n267748 );
buf ( R_12f94_1379c068 , n267790 );
buf ( R_f3d0_1264e3c8 , n267812 );
buf ( R_13cd6_10565638 , n267832 );
buf ( R_123b1_12b3e378 , n267842 );
buf ( R_144cf_f8c96f8 , n267848 );
buf ( R_13d0c_102f6168 , n267878 );
buf ( R_13c61_12081d78 , n267903 );
buf ( R_134f6_11ce6608 , n267910 );
buf ( R_112c2_12b294b8 , n267949 );
buf ( R_11922_1056c898 , n267992 );
buf ( R_11971_1207dbd8 , n268017 );
buf ( R_138_1265b308 , n268018 );
buf ( R_d2_12654c28 , n268019 );
buf ( R_23d_12656088 , n268020 );
buf ( R_8a_1379cba8 , n268021 );
buf ( R_38ad_12048418 , n268033 );
buf ( R_7b_12651de8 , n268034 );
buf ( R_13889_10564918 , n268052 );
buf ( R_13188_12079c18 , n268064 );
buf ( R_13b8c_13a15728 , n268107 );
buf ( R_947f_1056eaf8 , n268130 );
buf ( R_1d7_12649648 , n268131 );
buf ( R_149db_102f1668 , n268136 );
buf ( R_ac1d_120826d8 , n268171 );
buf ( R_13a06_105668f8 , n268215 );
buf ( R_18f_132fc988 , n268216 );
buf ( R_180_1265fea8 , n268217 );
buf ( R_10e36_11ce6d88 , n268261 );
buf ( R_136a7_12035cb8 , n268292 );
buf ( R_148df_13a1d608 , n268296 );
buf ( R_1380f_12080838 , n268336 );
buf ( R_1485b_1265a688 , n268342 );
buf ( R_14930_102f1a28 , n268347 );
buf ( R_10044_102f1c08 , n268370 );
buf ( R_d2a3_1207bbf8 , n268388 );
buf ( R_1c0_1203c0b8 , n268389 );
buf ( R_14f_12b25778 , n268390 );
buf ( R_8472_126654e8 , n268423 );
buf ( R_1483d_11ce0d48 , n268427 );
buf ( R_12b67_11cdf3a8 , n268449 );
buf ( R_11346_12655448 , n268463 );
buf ( R_13893_12084d98 , n268508 );
buf ( R_103f0_1207ecb8 , n268520 );
buf ( R_1308d_1379eea8 , n268542 );
buf ( R_f8ce_102f10c8 , n268564 );
buf ( R_13f82_11543978 , n268588 );
buf ( R_12359_133022e8 , n268610 );
buf ( R_12cd3_13a1f728 , n268658 );
buf ( R_13546_1153efb8 , n268703 );
buf ( R_143b6_115408b8 , n268708 );
buf ( R_148e5_10568518 , n268713 );
buf ( R_10a79_11545278 , n268726 );
buf ( R_1368d_102f3be8 , n268744 );
buf ( R_14002_12047518 , n268785 );
buf ( R_febc_1207caf8 , n268829 );
buf ( R_14987_10571d98 , n268835 );
buf ( R_14894_126569e8 , n268841 );
buf ( R_13e23_102f1708 , n268863 );
buf ( R_12304_10569e18 , n268873 );
buf ( R_12daa_f8cc218 , n268916 );
buf ( R_1289e_13316128 , n268937 );
buf ( R_146ea_132fd6a8 , n268943 );
buf ( R_104_12b414d8 , n268944 );
buf ( R_e9_12055a78 , n268945 );
buf ( R_226_12652568 , n268946 );
buf ( R_20b_12656bc8 , n268947 );
buf ( R_1484c_1056c078 , n268953 );
buf ( R_149fc_12077a58 , n268958 );
buf ( R_143f0_120442b8 , n268964 );
buf ( R_107_1203f538 , n268965 );
buf ( R_208_12b260d8 , n268966 );
buf ( R_1d2_1203ce78 , n268967 );
buf ( R_1442a_102f6668 , n268974 );
buf ( R_13d_1379c568 , n268975 );
buf ( R_134be_13a19148 , n268997 );
buf ( R_145cf_13304328 , n269002 );
buf ( R_12fa4_1153e0b8 , n269011 );
buf ( R_1053d_12079858 , n269041 );
buf ( R_ee_f8c86b8 , n269042 );
buf ( R_221_12652888 , n269043 );
buf ( R_13eb5_132f7ac8 , n269063 );
buf ( R_190_133178e8 , n269064 );
buf ( R_17f_115396f8 , n269065 );
buf ( R_137af_11ce6e28 , n269073 );
buf ( R_1455a_102ed748 , n269078 );
buf ( R_10db8_102f74c8 , n269111 );
buf ( R_ab_1264cde8 , n269112 );
buf ( R_1187e_12077698 , n269152 );
buf ( R_5a_126653a8 , n269153 );
buf ( R_7e57_13a1a188 , n269172 );
buf ( R_146ed_1153a238 , n269178 );
buf ( R_1b0_12b29918 , n269179 );
buf ( R_15f_1265f188 , n269180 );
buf ( R_138b8_1264a368 , n269199 );
buf ( R_13bd6_102f9188 , n269221 );
buf ( R_14a17_102f0ee8 , n269227 );
buf ( R_143a6_133121a8 , n269232 );
buf ( R_11f57_12649328 , n269254 );
buf ( R_14972_13302608 , n269260 );
buf ( R_10701_1207f1b8 , n269273 );
buf ( R_14503_1203e3b8 , n269279 );
buf ( R_a4_12b36e98 , n269280 );
buf ( R_6a_12b40178 , n269281 );
buf ( R_aeba_105624d8 , n269303 );
buf ( R_1379b_11ce6ec8 , n269322 );
buf ( R_134e2_13a1e3c8 , n269332 );
buf ( R_10973_12663008 , n269343 );
buf ( R_11c66_102f7ba8 , n269358 );
buf ( R_1325f_126468a8 , n269370 );
buf ( R_1327d_10570d58 , n269392 );
buf ( R_13417_102f3968 , n269413 );
buf ( R_101_1264f048 , n269414 );
buf ( R_95_133017a8 , n269415 );
buf ( R_20e_1265e788 , n269416 );
buf ( R_13c59_105b5638 , n269458 );
buf ( R_13ca1_12652f68 , n269480 );
buf ( R_1481c_11cdb988 , n269485 );
buf ( R_14611_11545458 , n269491 );
buf ( R_12fae_102f7388 , n269533 );
buf ( R_1469f_1207d138 , n269538 );
buf ( R_142dd_13314828 , n269548 );
buf ( R_1279d_12079fd8 , n269570 );
buf ( R_12646_1056b2b8 , n269592 );
buf ( R_11486_102ee788 , n269624 );
buf ( R_13389_1207fb18 , n269634 );
buf ( R_1492d_11ce64c8 , n269639 );
buf ( R_12d46_12648928 , n269660 );
buf ( R_145b7_12b3d5b8 , n269665 );
buf ( R_b211_12048c38 , n269687 );
buf ( R_143aa_13795c68 , n269692 );
buf ( R_1110c_11cdc928 , n269713 );
buf ( R_1a5_12b3c618 , n269714 );
buf ( R_16a_137a1248 , n269715 );
buf ( R_df67_1207b8d8 , n269758 );
buf ( R_124f6_1264f2c8 , n269790 );
buf ( R_12b54_102f2248 , n269812 );
buf ( R_d7dc_13a17de8 , n269825 );
buf ( R_1247b_11ce4808 , n269836 );
buf ( R_149ea_11540598 , n269842 );
buf ( R_10a_12b30678 , n269843 );
buf ( R_13c77_13a1cc08 , n269853 );
buf ( R_205_12653dc8 , n269854 );
buf ( R_14753_1264efa8 , n269860 );
buf ( R_191_12043d18 , n269861 );
buf ( R_17e_132f8568 , n269862 );
buf ( R_11c4b_13a15c28 , n269874 );
buf ( R_13208_11542758 , n269885 );
buf ( R_e0ad_133021a8 , n269897 );
buf ( R_11a3f_12b3e9b8 , n269908 );
buf ( R_1230e_f8cb598 , n269944 );
buf ( R_eee_1056adb8 , n269946 );
buf ( R_14444_12648108 , n269951 );
buf ( R_1dc_11538d98 , n269952 );
buf ( R_12b7a_1264f188 , n269995 );
buf ( R_133_13313888 , n269996 );
buf ( R_147b1_105b5a98 , n270002 );
buf ( R_f116_11ce1068 , n270025 );
buf ( R_13a5c_1379a268 , n270054 );
buf ( R_14340_12078458 , n270059 );
buf ( R_e522_1330ed28 , n270093 );
buf ( R_146f0_1153da78 , n270098 );
buf ( R_136f4_12649148 , n270119 );
buf ( R_119e8_1153e798 , n270141 );
buf ( R_1391b_12b277f8 , n270188 );
buf ( R_fd37_120394f8 , n270210 );
buf ( R_1461d_11539dd8 , n270216 );
buf ( R_ee50_102eb9e8 , n270229 );
buf ( R_dd_132f61c8 , n270230 );
buf ( R_232_105afa58 , n270231 );
buf ( R_4c_12652b08 , n270232 );
buf ( R_135a0_1153f0f8 , n270263 );
buf ( R_125d0_12b3f6d8 , n270291 );
buf ( R_b4_13302988 , n270292 );
buf ( R_51_13309648 , n270293 );
buf ( R_f925_12048b98 , n270315 );
buf ( R_14034_f8cf198 , n270322 );
buf ( R_123e9_f8c0eb8 , n270331 );
buf ( R_14726_1203bc58 , n270337 );
buf ( R_10894_1153ad78 , n270359 );
buf ( R_1b9_1379b7a8 , n270360 );
buf ( R_156_137927e8 , n270361 );
buf ( R_1471a_1379da08 , n270367 );
buf ( R_13d4e_11544f58 , n270384 );
buf ( R_112ae_115429d8 , n270406 );
buf ( R_dcb0_10564e18 , n270419 );
buf ( R_13ae3_12083498 , n270437 );
buf ( R_11a90_13a1ba88 , n270448 );
buf ( R_13f1a_10566998 , n270470 );
buf ( R_fdd5_1264d068 , n270483 );
buf ( R_13acb_13a17988 , n270503 );
buf ( R_ef1_13a16ee8 , n270505 );
buf ( R_145e1_12b40d58 , n270511 );
buf ( R_14915_102f7748 , n270515 );
buf ( R_ed3c_120760b8 , n270537 );
buf ( R_13cdc_11542398 , n270565 );
buf ( R_f544_102f5d08 , n270610 );
buf ( R_147e7_13793fa8 , n270615 );
buf ( R_e4_133095a8 , n270616 );
buf ( R_8d_1153d078 , n270617 );
buf ( R_78_12044178 , n270618 );
buf ( R_22b_12b3b538 , n270619 );
buf ( R_128ff_105b6178 , n270632 );
buf ( R_148ac_102f0f88 , n270637 );
buf ( R_1e9_133208a8 , n270638 );
buf ( R_192_12b44a98 , n270639 );
buf ( R_17d_12661f28 , n270640 );
buf ( R_12b83_13305e08 , n270650 );
buf ( R_fbb3_10567078 , n270672 );
buf ( R_126_12660588 , n270673 );
buf ( R_cfc6_1264a868 , n270715 );
buf ( R_1492a_13a1e1e8 , n270720 );
buf ( R_116bb_1207d6d8 , n270743 );
buf ( R_144d8_1330d9c8 , n270747 );
buf ( R_e6f2_102ecc08 , n270790 );
buf ( R_14a14_1207bdd8 , n270795 );
buf ( R_10f70_11544a58 , n270819 );
buf ( R_119fa_1207f2f8 , n270839 );
buf ( R_cef5_1265b6c8 , n270850 );
buf ( R_115b3_12082458 , n270872 );
buf ( R_211_1265c028 , n270873 );
buf ( R_146cc_11542618 , n270879 );
buf ( R_fe_120448f8 , n270880 );
buf ( R_119df_1056bad8 , n270890 );
buf ( R_13787_11ce21e8 , n270921 );
buf ( R_147dd_11ce6068 , n270926 );
buf ( R_14695_11cdf8a8 , n270932 );
buf ( R_149b1_102fa128 , n270938 );
buf ( R_110af_1379aee8 , n270945 );
buf ( R_14560_1330b3a8 , n270951 );
buf ( R_143ff_11cdca68 , n270958 );
buf ( R_d4_12654a48 , n270959 );
buf ( R_23b_13799408 , n270960 );
buf ( R_1c7_132fc0c8 , n270961 );
buf ( R_148_105aacd8 , n270962 );
buf ( R_13d6d_13a17668 , n270973 );
buf ( R_ce64_1056f9f8 , n270996 );
buf ( R_14474_13307a28 , n271000 );
buf ( R_12bde_102f62a8 , n271033 );
buf ( R_1436a_102eefa8 , n271038 );
buf ( R_14957_11540db8 , n271043 );
buf ( R_b634_11cdc068 , n271086 );
buf ( R_1460e_11ce2dc8 , n271091 );
buf ( R_f24f_11ce2fa8 , n271104 );
buf ( R_13763_105679d8 , n271120 );
buf ( R_f0b2_102f7f68 , n271142 );
buf ( R_14620_11ce6108 , n271147 );
buf ( R_131f5_12084618 , n271188 );
buf ( R_1490f_12651e88 , n271193 );
buf ( R_136cc_1264fcc8 , n271210 );
buf ( R_f227_1207a398 , n271233 );
buf ( R_13959_1153f918 , n271250 );
buf ( R_142cf_12659aa8 , n271255 );
buf ( R_f6b2_11cdfb28 , n271267 );
buf ( R_1ed_1203f5d8 , n271268 );
buf ( R_a2f6_11cdb3e8 , n271275 );
buf ( R_fc5e_13a18888 , n271286 );
buf ( R_122_12663d28 , n271287 );
buf ( R_13f67_12083b78 , n271305 );
buf ( R_13740_11cdb348 , n271312 );
buf ( R_146c9_1153fd78 , n271317 );
buf ( R_145db_13a12b68 , n271322 );
buf ( R_101ae_13a1fae8 , n271360 );
buf ( R_bb03_12b29ff8 , n271368 );
buf ( R_1101b_12045f38 , n271390 );
buf ( R_12bfd_10564b98 , n271404 );
buf ( R_121a5_1056a138 , n271415 );
buf ( R_127df_1330a728 , n271427 );
buf ( R_11617_105656d8 , n271437 );
buf ( R_13f90_12080518 , n271447 );
buf ( R_13be9_12662388 , n271487 );
buf ( R_12760_1331ab88 , n271522 );
buf ( R_126bb_10563b58 , n271534 );
buf ( R_147c6_12081cd8 , n271540 );
buf ( R_21c_12b41398 , n271541 );
buf ( R_13b33_102f0588 , n271559 );
buf ( R_1f8_132f5fe8 , n271560 );
buf ( R_11d2f_105665d8 , n271582 );
buf ( R_1227d_1265f2c8 , n271593 );
buf ( R_11a35_102f44a8 , n271603 );
buf ( R_1479c_1056c758 , n271609 );
buf ( R_116e4_12659828 , n271630 );
buf ( R_14662_1207ceb8 , n271634 );
buf ( R_14515_12079ad8 , n271638 );
buf ( R_117_12650c68 , n271639 );
buf ( R_115ca_11ce5fc8 , n271650 );
buf ( R_f3_1379bde8 , n271651 );
buf ( R_e229_102ecca8 , n271674 );
buf ( R_202_12b3f098 , n271675 );
buf ( R_1e5_1203a218 , n271676 );
buf ( R_12a_1331fea8 , n271677 );
buf ( R_10d_1330bda8 , n271678 );
buf ( R_135d6_1056fef8 , n271699 );
buf ( R_14918_13a1d888 , n271704 );
buf ( R_1452a_10564378 , n271710 );
buf ( R_14984_1056bc18 , n271715 );
buf ( R_1cd_1265c8e8 , n271716 );
buf ( R_eb34_11cda628 , n271762 );
buf ( R_125ac_11ce4308 , n271784 );
buf ( R_193_f8c7cb8 , n271785 );
buf ( R_1216d_1264d7e8 , n271829 );
buf ( R_17c_132fe648 , n271830 );
buf ( R_142_13792ce8 , n271831 );
buf ( R_cdb8_102f4f48 , n271851 );
buf ( R_144bd_11cdeb88 , n271856 );
buf ( R_131ae_1056bd58 , n271867 );
buf ( R_14909_1379f768 , n271873 );
buf ( R_14924_12b3adb8 , n271879 );
buf ( R_102a2_12b41e38 , n271912 );
buf ( R_13aa8_120525f8 , n271929 );
buf ( R_d3ca_102ef7c8 , n271940 );
buf ( R_1459f_120792b8 , n271946 );
buf ( R_120b3_12b407b8 , n271957 );
buf ( R_127a7_105683d8 , n272002 );
buf ( R_14545_1056b218 , n272008 );
buf ( R_12056_1204f178 , n272032 );
buf ( R_11f2a_10563ab8 , n272054 );
buf ( R_e021_12b26718 , n272065 );
buf ( R_f377_1056d1f8 , n272086 );
buf ( R_127ca_13a16da8 , n272096 );
buf ( R_14689_120838f8 , n272100 );
buf ( R_11be7_1207a6b8 , n272120 );
buf ( R_139a1_1264c668 , n272127 );
buf ( R_14536_12b42978 , n272131 );
buf ( R_13c2d_11cdd828 , n272171 );
buf ( R_14906_11544ff8 , n272177 );
buf ( R_11a5d_132f52c8 , n272187 );
buf ( R_ca63_1331c8e8 , n272211 );
buf ( R_14714_102f77e8 , n272216 );
buf ( R_14799_137933c8 , n272222 );
buf ( R_1390f_13a14828 , n272242 );
buf ( R_1234f_12083858 , n272265 );
buf ( R_142c6_12081738 , n272272 );
buf ( R_127ae_12b3ccf8 , n272291 );
buf ( R_13590_12079a38 , n272301 );
buf ( R_148b8_102eaa48 , n272306 );
buf ( R_5735_137a0988 , n272316 );
buf ( R_1a6_12038698 , n272317 );
buf ( R_169_1203e458 , n272318 );
buf ( R_127c1_12082638 , n272329 );
buf ( R_1288a_137a1ec8 , n272351 );
buf ( R_1488e_102f6708 , n272356 );
buf ( R_113b9_1264ea08 , n272388 );
buf ( R_1430f_11cd8fa8 , n272393 );
buf ( R_f97f_13304dc8 , n272406 );
buf ( R_104fa_120761f8 , n272419 );
buf ( R_119ae_11cdfa88 , n272429 );
buf ( R_12c78_1207ca58 , n272459 );
buf ( R_d606_11ce46c8 , n272482 );
buf ( R_146a5_102f90e8 , n272487 );
buf ( R_14900_120781d8 , n272492 );
buf ( R_1374f_13a16808 , n272500 );
buf ( R_ff3c_11ce1f68 , n272523 );
buf ( R_e834_10564238 , n272536 );
buf ( R_14a5e_105aa4b8 , n272541 );
buf ( R_13465_13316bc8 , n272571 );
buf ( R_13d25_11540b38 , n272601 );
buf ( R_56_13308248 , n272602 );
buf ( R_ef7_1153e838 , n272605 );
buf ( R_13193_102ec7a8 , n272617 );
buf ( R_132f1_13a145a8 , n272639 );
buf ( R_1291e_1056ee18 , n272649 );
buf ( R_14921_105640f8 , n272654 );
buf ( R_1371a_12083fd8 , n272662 );
buf ( R_14837_132f32e8 , n272668 );
buf ( R_13a37_12b3d338 , n272717 );
buf ( R_dad2_1379c6a8 , n272730 );
buf ( R_1495d_12b43878 , n272736 );
buf ( R_149f3_12b27c58 , n272740 );
buf ( R_107c6_1203f998 , n272750 );
buf ( R_1456c_12b437d8 , n272756 );
buf ( R_11888_13794868 , n272779 );
buf ( R_13b62_13a13428 , n272787 );
buf ( R_1360f_10563158 , n272828 );
buf ( R_1b1_12657ac8 , n272829 );
buf ( R_10844_1153e1f8 , n272862 );
buf ( R_194_1331d4c8 , n272863 );
buf ( R_17b_1265ea08 , n272864 );
buf ( R_15e_126544a8 , n272865 );
buf ( R_be25_102ec028 , n272872 );
buf ( R_148fd_102eb768 , n272877 );
buf ( R_14683_13a1d9c8 , n272881 );
buf ( R_a069_12080298 , n272898 );
buf ( R_1233a_13a143c8 , n272921 );
buf ( R_6e_13304b48 , n272922 );
buf ( R_1334f_1204e598 , n272932 );
buf ( R_121e7_1207ff78 , n272943 );
buf ( R_12bb7_102f3e68 , n272988 );
buf ( R_12bcc_12652608 , n273000 );
buf ( R_f783_13797b08 , n273022 );
buf ( R_14680_12076fb8 , n273028 );
buf ( R_13d2b_12085338 , n273059 );
buf ( R_11bbe_1153de38 , n273078 );
buf ( R_148e8_1264bda8 , n273083 );
buf ( R_148fa_102f5948 , n273088 );
buf ( R_149d8_132fc168 , n273093 );
buf ( R_148ee_120808d8 , n273099 );
buf ( R_148f4_11cd8468 , n273104 );
buf ( R_ff98_12b41618 , n273117 );
buf ( R_13bc3_102f8d28 , n273133 );
buf ( R_12b1f_120564d8 , n273155 );
buf ( R_c961_12080f18 , n273175 );
buf ( R_214_12655588 , n273176 );
buf ( R_dff5_102ed9c8 , n273206 );
buf ( R_13d49_13a16bc8 , n273226 );
buf ( R_fb_1379f808 , n273227 );
buf ( R_12958_102f1848 , n273272 );
buf ( R_12220_1379e908 , n273278 );
buf ( R_144de_12076798 , n273282 );
buf ( R_c6d1_10566178 , n273326 );
buf ( R_11547_1264cc08 , n273336 );
buf ( R_138ac_102eb128 , n273379 );
buf ( R_12853_105b58b8 , n273412 );
buf ( R_1f1_12655268 , n273413 );
buf ( R_11e_12b29b98 , n273414 );
buf ( R_13d30_1207b658 , n273442 );
buf ( R_b2_105aa0f8 , n273443 );
buf ( R_d5a1_105690f8 , n273466 );
buf ( R_c700_13304788 , n273478 );
buf ( R_a359_12662888 , n273487 );
buf ( R_1449f_12055898 , n273493 );
buf ( R_14587_10565ef8 , n273498 );
buf ( R_14759_1056e378 , n273503 );
buf ( R_1385d_1056ab38 , n273510 );
buf ( R_1401f_132fb588 , n273532 );
buf ( R_1245b_12658f68 , n273553 );
buf ( R_fe3a_11cdb168 , n273574 );
buf ( R_a47d_13a18f68 , n273582 );
buf ( R_145ea_1056c438 , n273588 );
buf ( R_99a4_102f5bc8 , n273606 );
buf ( R_1491e_12661528 , n273611 );
buf ( R_1c1_126618e8 , n273612 );
buf ( R_b180_12039a98 , n273655 );
buf ( R_14e_12b29e18 , n273656 );
buf ( R_13b1f_12052c38 , n273685 );
buf ( R_146e4_f8cb638 , n273691 );
buf ( R_14581_10571b18 , n273697 );
buf ( R_1354d_12040078 , n273716 );
buf ( R_13508_120842f8 , n273726 );
buf ( R_148d9_13a14d28 , n273732 );
buf ( R_149c0_102ed068 , n273736 );
buf ( R_1477e_10568fb8 , n273741 );
buf ( R_14735_105680b8 , n273745 );
buf ( R_13d35_11ce1108 , n273762 );
buf ( R_4d49_102f8dc8 , n273769 );
buf ( R_133aa_11545b38 , n273793 );
buf ( R_14518_102f67a8 , n273798 );
buf ( R_bf1d_1153d618 , n273839 );
buf ( R_a9_1204d4b8 , n273840 );
buf ( R_14702_12b3d0b8 , n273846 );
buf ( R_1431c_11cde188 , n273857 );
buf ( R_9323_1331d068 , n273869 );
buf ( R_14a2f_12075ed8 , n273874 );
buf ( R_1e1_13321ca8 , n273875 );
buf ( R_12e_105af9b8 , n273876 );
buf ( R_9d_1379c9c8 , n273877 );
buf ( R_12caa_126508a8 , n273898 );
buf ( R_115df_10566c18 , n273920 );
buf ( R_144fd_102f1b68 , n273926 );
buf ( R_127f1_12b2a098 , n273945 );
buf ( R_137eb_12082138 , n273964 );
buf ( R_11b9a_12b3f278 , n273986 );
buf ( R_1483a_12081f58 , n273992 );
buf ( R_7d2b_11ce4948 , n274000 );
buf ( R_13a49_102f8e68 , n274028 );
buf ( R_1493c_11cdc568 , n274033 );
buf ( R_14a3e_102ed428 , n274038 );
buf ( R_195_12045cb8 , n274039 );
buf ( R_14489_12b3fe58 , n274045 );
buf ( R_17a_1330dc48 , n274046 );
buf ( R_1066b_1264a228 , n274057 );
buf ( R_139b5_11536318 , n274065 );
buf ( R_12775_126513e8 , n274077 );
buf ( R_13d43_13a1c168 , n274095 );
buf ( R_13e78_1056a598 , n274107 );
buf ( R_90_f8cccb8 , n274108 );
buf ( R_75_12b443b8 , n274109 );
buf ( R_14816_10565db8 , n274115 );
buf ( R_e4c7_10571398 , n274159 );
buf ( R_14354_13317348 , n274164 );
buf ( R_146c3_12b3bfd8 , n274169 );
buf ( R_db95_12b2ff98 , n274180 );
buf ( R_b45b_11ce7508 , n274191 );
buf ( R_145de_1056b5d8 , n274196 );
buf ( R_13c7d_1056d798 , n274206 );
buf ( R_c7c0_102ed4c8 , n274234 );
buf ( R_1ff_13315c28 , n274235 );
buf ( R_1361a_102f01c8 , n274242 );
buf ( R_110_1204b938 , n274243 );
buf ( R_10c17_13a13888 , n274275 );
buf ( R_d6_1264b1c8 , n274276 );
buf ( R_239_12b2a958 , n274277 );
buf ( R_144a8_115369f8 , n274281 );
buf ( R_12516_13305188 , n274301 );
buf ( R_14699_10567e38 , n274307 );
buf ( R_12de4_12045b18 , n274315 );
buf ( R_10fd9_11ce1928 , n274338 );
buf ( R_145c6_13a1cb68 , n274343 );
buf ( R_147c3_13a177a8 , n274348 );
buf ( R_1313e_1207a1b8 , n274371 );
buf ( R_e9a6_1153dcf8 , n274383 );
buf ( R_123a6_12077418 , n274426 );
buf ( R_e669_1056eb98 , n274437 );
buf ( R_eea5_13793c88 , n274449 );
buf ( R_8e12_f8c7538 , n274466 );
buf ( R_11a2c_12b3f1d8 , n274498 );
buf ( R_bc89_12664548 , n274519 );
buf ( R_b132_13300a88 , n274541 );
buf ( R_14626_102f4ae8 , n274547 );
buf ( R_125c9_11ce5c08 , n274558 );
buf ( R_14891_1265e0a8 , n274562 );
buf ( R_13ba9_1056f4f8 , n274599 );
buf ( R_11299_1056a4f8 , n274620 );
buf ( R_1395f_1207ba18 , n274659 );
buf ( R_1085f_13312a28 , n274687 );
buf ( R_c642_12b41b18 , n274699 );
buf ( R_1445c_f8ce478 , n274703 );
buf ( R_14981_12b3f598 , n274707 );
buf ( R_148e2_12650b28 , n274712 );
buf ( R_988f_13a1e968 , n274755 );
buf ( R_962b_105647d8 , n274800 );
buf ( R_124a7_12079498 , n274840 );
buf ( R_fe64_1153f378 , n274872 );
buf ( R_11f16_102eb088 , n274894 );
buf ( R_13e03_1379bf28 , n274916 );
buf ( R_14927_11cdf808 , n274921 );
buf ( R_1ba_1330eb48 , n274922 );
buf ( R_14471_13793be8 , n274927 );
buf ( R_121fd_11ce3048 , n274939 );
buf ( R_14499_1207a9d8 , n274945 );
buf ( R_155_12b43f58 , n274946 );
buf ( R_98_12048af8 , n274947 );
buf ( R_e916_105699b8 , n274968 );
buf ( R_e1ea_1056b998 , n275001 );
buf ( R_11af3_13793788 , n275010 );
buf ( R_13bcf_12650948 , n275021 );
buf ( R_10070_12077e18 , n275034 );
buf ( R_f2f6_126613e8 , n275054 );
buf ( R_104a3_11542d98 , n275065 );
buf ( R_149ae_10565138 , n275069 );
buf ( R_1430b_1204c8d8 , n275076 );
buf ( R_ede8_1056dfb8 , n275088 );
buf ( R_13495_13a1e008 , n275109 );
buf ( R_df_132f6808 , n275110 );
buf ( R_230_12664a48 , n275111 );
buf ( R_136ac_102eacc8 , n275142 );
buf ( R_dd20_137974c8 , n275164 );
buf ( R_14741_132f2c08 , n275170 );
buf ( R_137c1_11543dd8 , n275178 );
buf ( R_14364_11ce6568 , n275183 );
buf ( R_11d60_132fc8e8 , n275196 );
buf ( R_14a44_105b60d8 , n275200 );
buf ( R_13749_11543518 , n275223 );
buf ( R_854a_1207fed8 , n275235 );
buf ( R_14a11_12045a78 , n275239 );
buf ( R_1a7_12659b48 , n275240 );
buf ( R_168_105b3158 , n275241 );
buf ( R_f03_13a17208 , n275243 );
buf ( R_1274c_12653fa8 , n275274 );
buf ( R_147b7_12079df8 , n275278 );
buf ( R_a2_1379e228 , n275279 );
buf ( R_63_f8c7b78 , n275280 );
buf ( R_13c49_102ecac8 , n275288 );
buf ( R_d68f_12078a98 , n275310 );
buf ( R_148f1_11cde688 , n275315 );
buf ( R_196_11536778 , n275316 );
buf ( R_179_13301c08 , n275317 );
buf ( R_11c1b_120757f8 , n275327 );
buf ( R_1181a_10565098 , n275340 );
buf ( R_14912_13300628 , n275346 );
buf ( R_10c93_13310768 , n275379 );
buf ( R_147f2_10571618 , n275383 );
buf ( R_c832_12075f78 , n275395 );
buf ( R_14530_11540778 , n275400 );
buf ( R_e8ba_11ce3b88 , n275411 );
buf ( R_14903_11ce50c8 , n275417 );
buf ( R_14629_115412b8 , n275423 );
buf ( R_11966_10562118 , n275445 );
buf ( R_f8fa_105b4d78 , n275457 );
buf ( R_1d8_1331f5e8 , n275458 );
buf ( R_1281b_1207f6b8 , n275470 );
buf ( R_137_1331a7c8 , n275471 );
buf ( R_5f_12b428d8 , n275472 );
buf ( R_12288_126495a8 , n275484 );
buf ( R_a469_13a14648 , n275505 );
buf ( R_130cc_13a17348 , n275526 );
buf ( R_136e6_11cdcb08 , n275554 );
buf ( R_d806_102f5a88 , n275575 );
buf ( R_fd98_12052d78 , n275598 );
buf ( R_144b4_1153eab8 , n275603 );
buf ( R_1482b_12b3b3f8 , n275608 );
buf ( R_13858_12081e18 , n275616 );
buf ( R_1d3_1265ae08 , n275617 );
buf ( R_13c_1265b1c8 , n275618 );
buf ( R_14596_12048558 , n275624 );
buf ( R_eb_1153bf98 , n275625 );
buf ( R_224_12b29698 , n275626 );
buf ( R_13d3c_132f70c8 , n275634 );
buf ( R_c353_102f31e8 , n275646 );
buf ( R_1092e_13a140a8 , n275652 );
buf ( R_1018e_10563478 , n275694 );
buf ( R_12875_1153eb58 , n275716 );
buf ( R_13693_13795448 , n275723 );
buf ( R_123bb_11ce7008 , n275734 );
buf ( R_dfc9_12647208 , n275745 );
buf ( R_da6d_12082098 , n275756 );
buf ( R_1198e_1153d758 , n275792 );
buf ( R_149ff_1264c848 , n275796 );
buf ( R_1180e_12648248 , n275828 );
buf ( R_12535_126604e8 , n275862 );
buf ( R_12780_10568b58 , n275873 );
buf ( R_9dc0_102f6f28 , n275894 );
buf ( R_c4a7_1330a908 , n275937 );
buf ( R_11bfb_12649968 , n275957 );
buf ( R_13fe4_105622f8 , n275979 );
buf ( R_12e0c_13797388 , n276001 );
buf ( R_1454e_11ce1c48 , n276005 );
buf ( R_14069_1153db18 , n276008 );
buf ( R_10c0e_120464d8 , n276019 );
buf ( R_13c1f_f8c8938 , n276027 );
buf ( R_d910_1056e418 , n276039 );
buf ( R_cfae_13a15368 , n276050 );
buf ( R_10806_1264d608 , n276062 );
buf ( R_13706_13319b48 , n276103 );
buf ( R_12e21_1330cb68 , n276139 );
buf ( R_f8_12665808 , n276140 );
buf ( R_67_105aac38 , n276141 );
buf ( R_217_105b3fb8 , n276142 );
buf ( R_12a8e_1264ef08 , n276152 );
buf ( R_e5ea_115436f8 , n276164 );
buf ( R_14858_10571c58 , n276169 );
buf ( R_111b8_102ebbc8 , n276190 );
buf ( R_12ba4_12b28ab8 , n276212 );
buf ( R_108f1_102f35a8 , n276231 );
buf ( R_138a5_1264e468 , n276260 );
buf ( R_131ff_13a1eaa8 , n276270 );
buf ( R_11448_11ce41c8 , n276282 );
buf ( R_11534_13a13ce8 , n276294 );
buf ( R_12d1d_1207c238 , n276316 );
buf ( R_134e8_13a1e8c8 , n276323 );
buf ( R_b82e_1153c2b8 , n276356 );
buf ( R_11572_11ce43a8 , n276379 );
buf ( R_14897_1265c988 , n276383 );
buf ( R_125fa_1265b128 , n276404 );
buf ( R_b95d_102f8008 , n276425 );
buf ( R_14436_10570718 , n276432 );
buf ( R_f951_132fcde8 , n276443 );
buf ( R_10246_1056ae58 , n276464 );
buf ( R_12041_11ce0ac8 , n276475 );
buf ( R_138cd_1153e018 , n276485 );
buf ( R_1b2_12660f88 , n276486 );
buf ( R_197_1379a768 , n276487 );
buf ( R_121dd_12659328 , n276499 );
buf ( R_178_12658d88 , n276500 );
buf ( R_15d_133195a8 , n276501 );
buf ( R_13f24_13318428 , n276514 );
buf ( R_146f6_132fbc68 , n276520 );
buf ( R_b880_12083d58 , n276531 );
buf ( R_12ab4_132f57c8 , n276544 );
buf ( R_ed14_133110c8 , n276556 );
buf ( R_144f0_132ff0e8 , n276562 );
buf ( R_10aa5_12053f98 , n276573 );
buf ( R_1290a_11ce1388 , n276586 );
buf ( R_9d4e_11cddbe8 , n276597 );
buf ( R_e6_12b344f8 , n276598 );
buf ( R_b0_12b3f458 , n276599 );
buf ( R_229_126659e8 , n276600 );
buf ( R_12b3f_105b6538 , n276609 );
buf ( R_1f5_1203e958 , n276610 );
buf ( R_f624_1265b808 , n276633 );
buf ( R_14711_11ce2828 , n276639 );
buf ( R_fe05_102f9548 , n276651 );
buf ( R_1118b_11cdb8e8 , n276665 );
buf ( R_1c8_f8c6b38 , n276666 );
buf ( R_147_12b38c98 , n276667 );
buf ( R_11a_1204b438 , n276668 );
buf ( R_14778_13a1f688 , n276672 );
buf ( R_137fd_11544418 , n276678 );
buf ( R_f0_13795d08 , n276679 );
buf ( R_c3_132ff188 , n276680 );
buf ( R_21f_1265a2c8 , n276681 );
buf ( R_12e60_132f3a68 , n276713 );
buf ( R_4a02_12646e48 , n276725 );
buf ( R_c5_12657e88 , n276726 );
buf ( R_132ae_1056ef58 , n276736 );
buf ( R_d400_133126a8 , n276781 );
buf ( R_128a8_f8c9978 , n276792 );
buf ( R_ecbd_12040a78 , n276815 );
buf ( R_146ba_11cd8c88 , n276820 );
buf ( R_ea59_102f5088 , n276856 );
buf ( R_1183a_1204a498 , n276891 );
buf ( R_13d1f_1207ddb8 , n276899 );
buf ( R_136e0_11ce7148 , n276941 );
buf ( R_ddb7_12078b38 , n276953 );
buf ( R_14575_13307c08 , n276957 );
buf ( R_14864_13a1b768 , n276961 );
buf ( R_1471d_12040bb8 , n276967 );
buf ( R_11237_1056f958 , n276978 );
buf ( R_13fee_12663288 , n276989 );
buf ( R_c1_1204fd58 , n276990 );
buf ( R_14632_11cd85a8 , n276994 );
buf ( R_4d_12662d88 , n276995 );
buf ( R_b895_1264a4a8 , n277004 );
buf ( R_11b87_12648b08 , n277034 );
buf ( R_111c4_12076658 , n277058 );
buf ( R_a534_12b3d018 , n277070 );
buf ( R_11805_12b41578 , n277079 );
buf ( R_c901_126603a8 , n277103 );
buf ( R_13bde_13a1bbc8 , n277113 );
buf ( R_149b4_10564d78 , n277118 );
buf ( R_c7_126589c8 , n277119 );
buf ( R_248_1331ef08 , n277120 );
buf ( R_5b_12655088 , n277121 );
buf ( R_13720_102f3f08 , n277141 );
buf ( R_b9b1_1056c9d8 , n277152 );
buf ( R_f1cc_10567ed8 , n277165 );
buf ( R_cd0b_11542f78 , n277176 );
buf ( R_1497b_11cdfda8 , n277180 );
buf ( R_12d6f_13799b88 , n277192 );
buf ( R_14305_120844d8 , n277199 );
buf ( R_145ae_102efe08 , n277205 );
buf ( R_147d6_12b27b18 , n277210 );
buf ( R_13dc3_11cdbf28 , n277222 );
buf ( R_dc22_1153d438 , n277233 );
buf ( R_5970_11cdbe88 , n277245 );
buf ( R_113_1265c528 , n277246 );
buf ( R_82_f8cbc78 , n277247 );
buf ( R_1fc_12050078 , n277248 );
buf ( R_b00a_1153e658 , n277259 );
buf ( R_1346e_10567bb8 , n277279 );
buf ( R_1dd_12b395f8 , n277280 );
buf ( R_10390_1207ed58 , n277292 );
buf ( R_12cf4_13310ee8 , n277304 );
buf ( R_10675_1203cab8 , n277316 );
buf ( R_1399b_1264c3e8 , n277326 );
buf ( R_132_120518d8 , n277327 );
buf ( R_d8_12b3c938 , n277328 );
buf ( R_237_105a9fb8 , n277329 );
buf ( R_d4b2_1265bda8 , n277352 );
buf ( R_14453_12649d28 , n277357 );
buf ( R_10e2c_102ecde8 , n277369 );
buf ( R_52_13799868 , n277370 );
buf ( R_143dc_120824f8 , n277376 );
buf ( R_13ebe_11ce4128 , n277398 );
buf ( R_14053_102f21a8 , n277412 );
buf ( R_10960_133050e8 , n277434 );
buf ( R_1037b_1264a048 , n277444 );
buf ( R_7fe6_12b3f638 , n277465 );
buf ( R_12685_11cdf088 , n277476 );
buf ( R_135e9_11ce0de8 , n277494 );
buf ( R_bf_1379fa88 , n277495 );
buf ( R_85_12b41898 , n277496 );
buf ( R_149d5_11541358 , n277502 );
buf ( R_13f4d_10561fd8 , n277510 );
buf ( R_d0f1_1056a1d8 , n277518 );
buf ( R_a3f3_12646da8 , n277536 );
buf ( R_1311d_13a131a8 , n277557 );
buf ( R_1026e_11541ad8 , n277567 );
buf ( R_139de_13310588 , n277576 );
buf ( R_144cc_11ce23c8 , n277582 );
buf ( R_1403a_1331cc08 , n277601 );
buf ( R_1ce_12656628 , n277602 );
buf ( R_198_12b3fdb8 , n277603 );
buf ( R_d37f_1379a1c8 , n277620 );
buf ( R_177_1330de28 , n277621 );
buf ( R_141_12b3cf78 , n277622 );
buf ( R_14500_102f92c8 , n277627 );
buf ( R_c9_12b28fb8 , n277628 );
buf ( R_246_1203df58 , n277629 );
buf ( R_93_12659be8 , n277630 );
buf ( R_72_132fe788 , n277631 );
buf ( R_125bf_105685b8 , n277641 );
buf ( R_1a8_137a0d48 , n277642 );
buf ( R_147a5_1264a728 , n277647 );
buf ( R_167_1204f678 , n277648 );
buf ( R_7f_105ac998 , n277649 );
buf ( R_149f0_13a1fea8 , n277653 );
buf ( R_12210_13793aa8 , n277673 );
buf ( R_13db7_11ce11a8 , n277686 );
buf ( R_100e9_132f3ec8 , n277698 );
buf ( R_5362_13a18108 , n277707 );
buf ( R_124d7_13a18e28 , n277717 );
buf ( R_14a55_133001c8 , n277723 );
buf ( R_12419_1153d398 , n277735 );
buf ( R_108b6_1264e0a8 , n277747 );
buf ( R_10d4d_11cded68 , n277758 );
buf ( R_1464a_13a15b88 , n277764 );
buf ( R_c7f2_11cdc748 , n277774 );
buf ( R_13c83_11544698 , n277782 );
buf ( R_1489a_f8c6c78 , n277786 );
buf ( R_125b6_12040b18 , n277797 );
buf ( R_c00b_12079718 , n277809 );
buf ( R_eeb_13a13608 , n277815 );
buf ( R_f088_1330ba88 , n277828 );
buf ( R_1365e_1207b838 , n277847 );
buf ( R_fa81_12052198 , n277859 );
buf ( R_145f3_13a14788 , n277863 );
buf ( R_10995_102f3148 , n277884 );
buf ( R_123f8_13a13388 , n277890 );
buf ( R_6358_1204fe98 , n277914 );
buf ( R_14763_11ce4c68 , n277920 );
buf ( R_1433c_12077c38 , n277925 );
buf ( R_dde7_13a141e8 , n277937 );
buf ( R_13ef9_1204a858 , n277946 );
buf ( R_14810_1056db58 , n277951 );
buf ( R_13fdc_102f15c8 , n277971 );
buf ( R_d995_11ce0fc8 , n277982 );
buf ( R_117fc_12056078 , n277994 );
buf ( R_8d57_11ce53e8 , n278006 );
buf ( R_11bb4_12b39cd8 , n278015 );
buf ( R_13b97_1207a438 , n278043 );
buf ( R_14068_11cdc108 , n278046 );
buf ( R_1335a_105b5ef8 , n278067 );
buf ( R_1043d_13a1c5c8 , n278078 );
buf ( R_128cf_11cdabc8 , n278111 );
buf ( R_1219b_1207a938 , n278134 );
buf ( R_10dce_105631f8 , n278146 );
buf ( R_bbfa_10564418 , n278154 );
buf ( R_11864_12b44318 , n278165 );
buf ( R_12435_11ce4088 , n278186 );
buf ( R_a7_1265a5e8 , n278187 );
buf ( R_111f4_11cdf6c8 , n278216 );
buf ( R_135cf_1207eb78 , n278223 );
buf ( R_102ef_1153c218 , n278236 );
buf ( R_12ca0_11ce0668 , n278259 );
buf ( R_1c2_1330f228 , n278260 );
buf ( R_c6f4_12056438 , n278282 );
buf ( R_1404f_12b3e738 , n278289 );
buf ( R_ee7b_1379a628 , n278301 );
buf ( R_127e9_f8c8078 , n278312 );
buf ( R_14d_1203cbf8 , n278313 );
buf ( R_bd_1203f3f8 , n278314 );
buf ( R_48_13301848 , n278315 );
buf ( R_10afa_13a15d68 , n278327 );
buf ( R_ed66_11ce3368 , n278339 );
buf ( R_13a92_102f0bc8 , n278346 );
buf ( R_e9fb_12646268 , n278367 );
buf ( R_10d30_12084078 , n278378 );
buf ( R_149ab_1153d7f8 , n278382 );
buf ( R_88_13300d08 , n278383 );
buf ( R_6b_105aaff8 , n278384 );
buf ( R_11c31_115418f8 , n278396 );
buf ( R_13677_102f9868 , n278405 );
buf ( R_133f2_1379f088 , n278431 );
buf ( R_13edf_120837b8 , n278453 );
buf ( R_d399_137980a8 , n278476 );
buf ( R_1446e_1207d958 , n278480 );
buf ( R_1382d_1207d9f8 , n278488 );
buf ( R_cb_1331fa48 , n278489 );
buf ( R_244_1264c708 , n278490 );
buf ( R_12dc8_13a1f548 , n278501 );
buf ( R_12299_1265d1a8 , n278523 );
buf ( R_1474a_12076dd8 , n278528 );
buf ( R_13844_12663aa8 , n278549 );
buf ( R_13c11_1153d578 , n278568 );
buf ( R_14650_1056f278 , n278572 );
buf ( R_146fc_12647848 , n278578 );
buf ( R_10f84_1207bab8 , n278588 );
buf ( R_131cc_12b272f8 , n278608 );
buf ( R_1451b_10567cf8 , n278613 );
buf ( R_14390_10567c58 , n278621 );
buf ( R_13754_12082318 , n278627 );
buf ( R_1bb_12664868 , n278628 );
buf ( R_154_1204e1d8 , n278629 );
buf ( R_14831_1264f408 , n278635 );
buf ( R_7c_105b1cb8 , n278636 );
buf ( R_f1a0_12075938 , n278648 );
buf ( R_e9d0_1153f558 , n278660 );
buf ( R_f0eb_102f7568 , n278692 );
buf ( R_fb0c_1331a368 , n278704 );
buf ( R_1397b_1331b268 , n278712 );
buf ( R_e589_1379bb68 , n278724 );
buf ( R_1381a_120547b8 , n278731 );
buf ( R_1463e_105703f8 , n278736 );
buf ( R_12e76_11cd9908 , n278746 );
buf ( R_199_132fb3a8 , n278747 );
buf ( R_176_12b265d8 , n278748 );
buf ( R_125_13798008 , n278749 );
buf ( R_11ad2_102ed108 , n278772 );
buf ( R_1ea_1265a868 , n278773 );
buf ( R_10764_11cd9548 , n278794 );
buf ( R_14563_1264d6a8 , n278800 );
buf ( R_12c1a_102f0268 , n278831 );
buf ( R_146d2_1203a998 , n278835 );
buf ( R_147bd_102f9048 , n278839 );
buf ( R_fa57_1207f398 , n278851 );
buf ( R_c5a3_120849d8 , n278883 );
buf ( R_11dc9_f8c9b58 , n278908 );
buf ( R_11d95_1153f198 , n278935 );
buf ( R_1329b_11cd95e8 , n278946 );
buf ( R_14861_f8c41f8 , n278951 );
buf ( R_1064a_10561f38 , n278962 );
buf ( R_ce07_f8c8f78 , n278973 );
buf ( R_14720_11ce07a8 , n278978 );
buf ( R_13ca7_12078098 , n278987 );
buf ( R_147f5_1207a078 , n278992 );
buf ( R_142d3_12036758 , n278997 );
buf ( R_13dee_12083a38 , n279019 );
buf ( R_ec91_126490a8 , n279031 );
buf ( R_13421_11544c38 , n279042 );
buf ( R_cf92_11cdfee8 , n279051 );
buf ( R_4c49_13a1d748 , n279063 );
buf ( R_114d1_13307de8 , n279075 );
buf ( R_cff7_12076bf8 , n279086 );
buf ( R_142ff_11ce1b08 , n279093 );
buf ( R_139c0_13a1e5a8 , n279115 );
buf ( R_143cc_1056e738 , n279122 );
buf ( R_ba4e_13a1d388 , n279143 );
buf ( R_12485_105b6358 , n279165 );
buf ( R_11f0c_13a1aea8 , n279176 );
buf ( R_14867_12054b78 , n279180 );
buf ( R_137b5_10569cd8 , n279186 );
buf ( R_11d1b_12649288 , n279199 );
buf ( R_13d7b_102f56c8 , n279218 );
buf ( R_14a2c_102f12a8 , n279224 );
buf ( R_14608_13a155e8 , n279229 );
buf ( R_144c9_10571578 , n279234 );
buf ( R_fc0a_11541858 , n279256 );
buf ( R_144fa_120775f8 , n279260 );
buf ( R_129_1331c988 , n279261 );
buf ( R_13561_1330d068 , n279272 );
buf ( R_e1_12661708 , n279273 );
buf ( R_1299a_1207b158 , n279285 );
buf ( R_1489d_105686f8 , n279290 );
buf ( R_22e_132f2ac8 , n279291 );
buf ( R_6d01_102f72e8 , n279302 );
buf ( R_ffc3_12656e48 , n279314 );
buf ( R_1496f_102f9908 , n279320 );
buf ( R_1e6_13792a68 , n279321 );
buf ( R_14760_11ce3868 , n279325 );
buf ( R_d2d1_13793468 , n279354 );
buf ( R_12145_1207b978 , n279365 );
buf ( R_f5_11537038 , n279366 );
buf ( R_bb_13799cc8 , n279367 );
buf ( R_21a_1265b088 , n279368 );
buf ( R_14975_11541998 , n279372 );
buf ( R_147c0_11ce20a8 , n279376 );
buf ( R_13b7f_1153a198 , n279384 );
buf ( R_13615_12084c58 , n279393 );
buf ( R_14a29_10571438 , n279397 );
buf ( R_13526_102f49a8 , n279408 );
buf ( R_11215_12075b18 , n279420 );
buf ( R_10e4c_13a169e8 , n279430 );
buf ( R_13d97_105651d8 , n279441 );
buf ( R_1b3_1379b348 , n279442 );
buf ( R_13fab_11538758 , n279452 );
buf ( R_10ff9_105aad78 , n279462 );
buf ( R_145c0_11cd7f68 , n279467 );
buf ( R_145fc_120476f8 , n279471 );
buf ( R_15c_137992c8 , n279472 );
buf ( R_67bc_13311028 , n279479 );
buf ( R_efc2_11cdefe8 , n279491 );
buf ( R_145cc_132f8388 , n279495 );
buf ( R_ae_1379c1a8 , n279496 );
buf ( R_1263c_11cdf768 , n279508 );
buf ( R_57_126522e8 , n279509 );
buf ( R_14659_1264e1e8 , n279515 );
buf ( R_13899_133075c8 , n279533 );
buf ( R_125e5_13311348 , n279566 );
buf ( R_113fb_11ce7288 , n279587 );
buf ( R_11e0e_102f4908 , n279599 );
buf ( R_11270_12b29a58 , n279607 );
buf ( R_f61a_13305cc8 , n279618 );
buf ( R_1499f_133198c8 , n279623 );
buf ( R_121_13795808 , n279624 );
buf ( R_106_12b25a98 , n279625 );
buf ( R_1458a_102eb268 , n279629 );
buf ( R_126cf_13a19788 , n279640 );
buf ( R_209_1379cb08 , n279641 );
buf ( R_1ee_12656268 , n279642 );
buf ( R_12c5a_102ef688 , n279654 );
buf ( R_1270e_11cdb708 , n279666 );
buf ( R_e437_102f2c48 , n279679 );
buf ( R_147cf_11ce5168 , n279685 );
buf ( R_e233_1056d338 , n279696 );
buf ( R_13bbe_11ce55c8 , n279726 );
buf ( R_11e6b_1207d458 , n279740 );
buf ( R_13f0b_12b42f18 , n279751 );
buf ( R_103_12b41c58 , n279752 );
buf ( R_cd_12b39a58 , n279753 );
buf ( R_242_12654688 , n279754 );
buf ( R_20c_12b43c38 , n279755 );
buf ( R_11ce5_1379e048 , n279765 );
buf ( R_ef4_1056dc98 , n279768 );
buf ( R_11823_13a15fe8 , n279778 );
buf ( R_130b8_13a12988 , n279790 );
buf ( R_12baf_12648ba8 , n279812 );
buf ( R_119a4_102f3288 , n279823 );
buf ( R_f4e5_1264b308 , n279834 );
buf ( R_12c6f_11cdea48 , n279845 );
buf ( R_1473b_102fa308 , n279849 );
buf ( R_8b_132f8608 , n279850 );
buf ( R_11467_105659f8 , n279861 );
buf ( R_11b4a_11ce1568 , n279870 );
buf ( R_137f7_12077878 , n279889 );
buf ( R_e5b5_1153d938 , n279900 );
buf ( R_14775_13a1bda8 , n279906 );
buf ( R_14671_1264ab88 , n279911 );
buf ( R_14066_12084258 , n279914 );
buf ( R_13954_12076518 , n279923 );
buf ( R_de4d_12b26538 , n279947 );
buf ( R_149f6_11cda308 , n279951 );
buf ( R_aff6_102f4a48 , n279963 );
buf ( R_d75d_1207c0f8 , n279974 );
buf ( R_10f46_12081ff8 , n279986 );
buf ( R_c50b_11cdd3c8 , n280006 );
buf ( R_136ed_12082ef8 , n280015 );
buf ( R_101d1_1056e198 , n280037 );
buf ( R_1a9_12037658 , n280038 );
buf ( R_166_120507f8 , n280039 );
buf ( R_9b_12b3b178 , n280040 );
buf ( R_bb16_12650268 , n280058 );
buf ( R_1265a_105635b8 , n280068 );
buf ( R_b802_1265dba8 , n280078 );
buf ( R_131ea_102f4cc8 , n280098 );
buf ( R_14a0e_10570e98 , n280102 );
buf ( R_19a_12662068 , n280103 );
buf ( R_175_12b3fc78 , n280104 );
buf ( R_109_12b2c7f8 , n280105 );
buf ( R_206_105b5b38 , n280106 );
buf ( R_146b4_1153fcd8 , n280111 );
buf ( R_11e21_11cd9e08 , n280126 );
buf ( R_104ba_f8c7218 , n280150 );
buf ( R_13fbc_11541218 , n280159 );
buf ( R_144ba_102f8c88 , n280164 );
buf ( R_11622_102ed388 , n280184 );
buf ( R_13c02_12b29198 , n280192 );
buf ( R_13ba3_105626b8 , n280209 );
buf ( R_ff0f_12081918 , n280231 );
buf ( R_123d6_11541e98 , n280242 );
buf ( R_fd64_102f3328 , n280255 );
buf ( R_14486_102ef728 , n280259 );
buf ( R_13776_1379fd08 , n280267 );
buf ( R_14665_132f5ae8 , n280271 );
buf ( R_10098_13793968 , n280283 );
buf ( R_11072_13a1ed28 , n280294 );
buf ( R_14554_10565778 , n280298 );
buf ( R_137a8_1056b678 , n280340 );
buf ( R_11b55_12649a08 , n280351 );
buf ( R_14411_12663508 , n280356 );
buf ( R_84a7_12b40fd8 , n280376 );
buf ( R_133fc_1153ee78 , n280387 );
buf ( R_da_1331b088 , n280388 );
buf ( R_a0_1379b2a8 , n280389 );
buf ( R_235_1264d4c8 , n280390 );
buf ( R_1333b_11542c58 , n280409 );
buf ( R_132e7_11ce28c8 , n280419 );
buf ( R_1357d_1153feb8 , n280428 );
buf ( R_14644_1056d978 , n280433 );
buf ( R_100_1265f0e8 , n280434 );
buf ( R_79_137a1388 , n280435 );
buf ( R_e0d7_126556c8 , n280468 );
buf ( R_11b42_1264b6c8 , n280479 );
buf ( R_20f_12b28018 , n280480 );
buf ( R_f4db_1207bfb8 , n280492 );
buf ( R_1193e_13a19968 , n280502 );
buf ( R_138d5_1379b848 , n280511 );
buf ( R_13e4c_1207f118 , n280534 );
buf ( R_13a7e_102f6ac8 , n280543 );
buf ( R_12d79_102ee468 , n280554 );
buf ( R_116a8_12084398 , n280563 );
buf ( R_116_1265f868 , n280564 );
buf ( R_148a3_11cdecc8 , n280569 );
buf ( R_13273_13a1a688 , n280590 );
buf ( R_1f9_1379ddc8 , n280591 );
buf ( R_1025b_1330bee8 , n280600 );
buf ( R_122e8_12b39878 , n280612 );
buf ( R_11ba2_11544738 , n280633 );
buf ( R_12521_1056c258 , n280668 );
buf ( R_e8e6_f8cf4b8 , n280680 );
buf ( R_8cd2_1264ac28 , n280693 );
buf ( R_11a11_126477a8 , n280702 );
buf ( R_143c6_120850b8 , n280709 );
buf ( R_13e99_12039e58 , n280720 );
buf ( R_1466b_13306808 , n280724 );
buf ( R_14465_1207a758 , n280729 );
buf ( R_134b3_102f3468 , n280739 );
buf ( R_11fe7_1330c3e8 , n280751 );
buf ( R_1258d_13a14dc8 , n280771 );
buf ( R_14677_105712f8 , n280777 );
buf ( R_1367d_102eb628 , n280785 );
buf ( R_1e2_12663c88 , n280786 );
buf ( R_b9_12661848 , n280787 );
buf ( R_12d_12660268 , n280788 );
buf ( R_f47c_1153ded8 , n280810 );
buf ( R_1468c_13a1aae8 , n280815 );
buf ( R_145ba_120815f8 , n280819 );
buf ( R_14790_11cd9cc8 , n280824 );
buf ( R_14419_12048f58 , n280829 );
buf ( R_13bb3_1207b6f8 , n280836 );
buf ( R_1046b_105688d8 , n280843 );
buf ( R_1232e_13314008 , n280855 );
buf ( R_1170d_1264c528 , n280866 );
buf ( R_14a41_1056fa98 , n280870 );
buf ( R_14459_11cd92c8 , n280874 );
buf ( R_14480_11cdcf68 , n280880 );
buf ( R_13a88_11ce3f48 , n280887 );
buf ( R_c8f0_102f0d08 , n280896 );
buf ( R_134ff_1056bf38 , n280906 );
buf ( R_aac5_13a18748 , n280928 );
buf ( R_14509_13a1e148 , n280933 );
buf ( R_cebc_12039d18 , n280954 );
buf ( R_135bd_12081058 , n280963 );
buf ( R_147ba_12078ef8 , n280968 );
buf ( R_f4a6_105654f8 , n280979 );
buf ( R_1182e_13a19aa8 , n280988 );
buf ( R_142eb_11cdec28 , n280995 );
buf ( R_13bf5_10568ab8 , n281001 );
buf ( R_12093_12077058 , n281011 );
buf ( R_13dac_13a15688 , n281022 );
buf ( R_dc51_13304f08 , n281044 );
buf ( R_13e8f_1264a0e8 , n281056 );
buf ( R_13c89_12b39f58 , n281073 );
buf ( R_f0be_102f1de8 , n281086 );
buf ( R_9373_10563e78 , n281111 );
buf ( R_11a48_13a195a8 , n281120 );
buf ( R_f3f9_1153f9b8 , n281132 );
buf ( R_1d4_12b42fb8 , n281133 );
buf ( R_e3f1_12b25bd8 , n281145 );
buf ( R_13c27_13309b48 , n281154 );
buf ( R_240_105ab4f8 , n281155 );
buf ( R_cf_13311a28 , n281156 );
buf ( R_13c38_1204a3f8 , n281162 );
buf ( R_13b_13300f88 , n281163 );
buf ( R_11ef6_11cd7888 , n281174 );
buf ( R_135c9_11ce6888 , n281182 );
buf ( R_116d1_1153d898 , n281192 );
buf ( R_149d2_12080158 , n281198 );
buf ( R_ba5b_12b403f8 , n281211 );
buf ( R_ea84_1330ca28 , n281222 );
buf ( R_f59a_11ce3908 , n281234 );
buf ( R_1496c_1331e968 , n281239 );
buf ( R_12bd5_11ce3fe8 , n281249 );
buf ( R_1253e_105b6678 , n281259 );
buf ( R_14873_11cd79c8 , n281264 );
buf ( R_149a5_132ff868 , n281268 );
buf ( R_14512_11540bd8 , n281272 );
buf ( R_14756_10565318 , n281277 );
buf ( R_1c9_13313a68 , n281278 );
buf ( R_d09b_12660948 , n281284 );
buf ( R_203_12050cf8 , n281285 );
buf ( R_10c_12038058 , n281286 );
buf ( R_146_12b42298 , n281287 );
buf ( R_136c1_12b276b8 , n281295 );
buf ( R_1480a_12649e68 , n281301 );
buf ( R_1d9_1379e7c8 , n281302 );
buf ( R_13e84_1056ad18 , n281315 );
buf ( R_1021c_1056fc78 , n281326 );
buf ( R_136_132fe6e8 , n281327 );
buf ( R_145ff_102ef2c8 , n281331 );
buf ( R_19b_12b28dd8 , n281332 );
buf ( R_1031a_11540e58 , n281345 );
buf ( R_1f2_11538438 , n281346 );
buf ( R_13114_102f3648 , n281358 );
buf ( R_ec36_12042af8 , n281381 );
buf ( R_222_133189c8 , n281382 );
buf ( R_6f_12b3a458 , n281383 );
buf ( R_96_1203c838 , n281384 );
buf ( R_ed_1203deb8 , n281385 );
buf ( R_11d_1204c838 , n281386 );
buf ( R_174_13318928 , n281387 );
buf ( R_119f1_13316588 , n281406 );
buf ( R_1486a_13a1d428 , n281410 );
buf ( R_11717_1207d778 , n281420 );
buf ( R_14781_115447d8 , n281424 );
buf ( R_13995_12038738 , n281432 );
buf ( R_e4f5_12049598 , n281443 );
buf ( R_74a9_12645d68 , n281452 );
buf ( R_10208_12038558 , n281474 );
buf ( R_145ab_12b3f9f8 , n281479 );
buf ( R_227_1331e508 , n281480 );
buf ( R_e8_133028e8 , n281481 );
buf ( R_13809_1153faf8 , n281488 );
buf ( R_f732_12649008 , n281499 );
buf ( R_14524_137968e8 , n281504 );
buf ( R_146d8_11cd94a8 , n281509 );
buf ( R_14064_1264d2e8 , n281512 );
buf ( R_12dfa_11cd88c8 , n281523 );
buf ( R_135ef_102f0a88 , n281530 );
buf ( R_10ee5_12047798 , n281539 );
buf ( R_14548_120493b8 , n281544 );
buf ( R_11030_11cdbca8 , n281554 );
buf ( R_1400f_13a1a368 , n281563 );
buf ( R_f051_1264e6e8 , n281576 );
buf ( R_de7c_102eafe8 , n281599 );
buf ( R_13538_120754d8 , n281611 );
buf ( R_13e56_12b297d8 , n281633 );
buf ( R_84eb_1331c2a8 , n281640 );
buf ( R_1498a_1207e3f8 , n281644 );
buf ( R_148a6_115459f8 , n281648 );
buf ( R_212_1330bd08 , n281649 );
buf ( R_fd_13307d48 , n281650 );
buf ( R_144a5_13a1c028 , n281654 );
buf ( R_10110_120369d8 , n281665 );
buf ( R_12b5e_12651208 , n281675 );
buf ( R_149ed_13303428 , n281679 );
buf ( R_144db_12078598 , n281683 );
buf ( R_bf9f_11cd9b88 , n281703 );
buf ( R_14017_f8c20d8 , n281712 );
buf ( R_13a3d_f8ca918 , n281720 );
buf ( R_13b2d_120830d8 , n281727 );
buf ( R_8e_132f37e8 , n281728 );
buf ( R_12aeb_120810f8 , n281737 );
buf ( R_a23e_11ce5ca8 , n281744 );
buf ( R_12ce9_12081c38 , n281755 );
buf ( R_f00_1207c058 , n281758 );
buf ( R_c1fe_1264be48 , n281770 );
buf ( R_f2d2_11cdf948 , n281793 );
buf ( R_14385_12044c18 , n281803 );
buf ( R_143c0_1265fb88 , n281810 );
buf ( R_14496_13a1c668 , n281814 );
buf ( R_14738_12b28bf8 , n281820 );
buf ( R_cab9_102f99a8 , n281832 );
buf ( R_1255c_f8c61d8 , n281842 );
buf ( R_143ba_11cde868 , n281847 );
buf ( R_147c9_13a18ce8 , n281852 );
buf ( R_13311_13a198c8 , n281863 );
buf ( R_147a2_102f2ce8 , n281867 );
buf ( R_fbe0_13a1b628 , n281880 );
buf ( R_dcc6_12664ae8 , n281892 );
buf ( R_103cf_12085158 , n281902 );
buf ( R_13909_1204f5d8 , n281910 );
buf ( R_1197b_115433d8 , n281921 );
buf ( R_144e1_13a1f4a8 , n281926 );
buf ( R_145a2_11cd7ce8 , n281930 );
buf ( R_12d50_120851f8 , n281939 );
buf ( R_12380_10563338 , n281951 );
buf ( R_107a7_1379f9e8 , n281960 );
buf ( R_10e8a_102ea688 , n281967 );
buf ( R_122fb_13a17708 , n281979 );
buf ( R_12aa7_12037798 , n281990 );
buf ( R_12107_1264d428 , n282001 );
buf ( R_14533_1330c8e8 , n282005 );
buf ( R_14542_120759d8 , n282011 );
buf ( R_4276_102effe8 , n282022 );
buf ( R_1478d_115453b8 , n282028 );
buf ( R_130c1_11542258 , n282037 );
buf ( R_13ff8_102f9fe8 , n282048 );
buf ( R_1aa_13795268 , n282049 );
buf ( R_116b1_13a159a8 , n282058 );
buf ( R_1bc_126536e8 , n282059 );
buf ( R_b76e_1153c8f8 , n282069 );
buf ( R_4e_13792e28 , n282070 );
buf ( R_60_12b44bd8 , n282071 );
buf ( R_a5_13311668 , n282072 );
buf ( R_b7_1379f948 , n282073 );
buf ( R_153_13793288 , n282074 );
buf ( R_165_13306948 , n282075 );
buf ( R_f9fe_102f9408 , n282087 );
buf ( R_14431_12080478 , n282094 );
buf ( R_1c3_12047158 , n282095 );
buf ( R_64_f8c1bd8 , n282096 );
buf ( R_14c_120387d8 , n282097 );
buf ( R_12471_102f7068 , n282108 );
buf ( R_148c1_13316f88 , n282113 );
buf ( R_11433_1265f048 , n282149 );
buf ( R_13ce2_1264aa48 , n282156 );
buf ( R_121bd_115449b8 , n282166 );
buf ( R_14813_10566d58 , n282171 );
buf ( R_147fb_102f83c8 , n282175 );
buf ( R_146ab_12051658 , n282180 );
buf ( R_12c65_1264cb68 , n282191 );
buf ( R_e2b4_f8c0f58 , n282202 );
buf ( R_10c61_120805b8 , n282213 );
buf ( R_10f1d_10566df8 , n282223 );
buf ( R_10de4_1379b5c8 , n282235 );
buf ( R_ae51_105ab098 , n282248 );
buf ( R_146f3_12659d28 , n282253 );
buf ( R_d03f_126484c8 , n282264 );
buf ( R_9fe2_11543fb8 , n282274 );
buf ( R_10b79_12657028 , n282295 );
buf ( R_64c2_12662748 , n282302 );
buf ( R_139d0_102f1fc8 , n282314 );
buf ( R_13639_1207f578 , n282321 );
buf ( R_1b4_12654728 , n282322 );
buf ( R_1cf_133184c8 , n282323 );
buf ( R_e214_1207ae38 , n282334 );
buf ( R_140_12665448 , n282335 );
buf ( R_15b_f8c0378 , n282336 );
buf ( R_1435c_13304d28 , n282341 );
buf ( R_10745_12056898 , n282351 );
buf ( R_1044f_120557f8 , n282360 );
buf ( R_10824_11ce3188 , n282369 );
buf ( R_13820_12b41438 , n282376 );
buf ( R_69b8_11cdc888 , n282386 );
buf ( R_124b9_1056d658 , n282393 );
buf ( R_143f4_102edd88 , n282398 );
buf ( R_142f5_1264a908 , n282405 );
buf ( R_76_f8ca198 , n282406 );
buf ( R_ac_12660a88 , n282407 );
buf ( R_1269b_11cd9368 , n282416 );
buf ( R_147b4_120766f8 , n282420 );
buf ( R_14834_13a16a88 , n282425 );
buf ( R_12e88_102f8a08 , n282431 );
buf ( R_f021_102ec168 , n282443 );
buf ( R_f6dd_13a163a8 , n282454 );
buf ( R_145e4_126463a8 , n282459 );
buf ( R_14723_1264db08 , n282464 );
buf ( R_173_f8c3438 , n282465 );
buf ( R_19c_12b40218 , n282466 );
buf ( R_11142_10562f78 , n282475 );
buf ( R_23e_1265bc68 , n282476 );
buf ( R_d1_13311f28 , n282477 );
buf ( R_13512_12080dd8 , n282488 );
buf ( R_7859_11cdaee8 , n282499 );
buf ( R_14593_115458b8 , n282504 );
buf ( R_148a9_12647ac8 , n282508 );
buf ( R_10577_11545318 , n282514 );
buf ( R_133ca_1203e098 , n282526 );
buf ( R_13b92_13a14be8 , n282544 );
buf ( R_10efd_102ec3e8 , n282554 );
buf ( R_f0b_1153f4b8 , n282557 );
buf ( R_12e15_10568018 , n282567 );
buf ( R_200_12b29eb8 , n282568 );
buf ( R_21d_137a03e8 , n282569 );
buf ( R_f2_12652ec8 , n282570 );
buf ( R_10f_12b3e5f8 , n282571 );
buf ( R_ca13_11ce4628 , n282579 );
buf ( R_14966_11546218 , n282583 );
buf ( R_13ad8_1203a358 , n282589 );
buf ( R_12d8d_105b5db8 , n282600 );
buf ( R_10165_1264cac8 , n282612 );
buf ( R_1337f_13a12c08 , n282623 );
buf ( R_53_f8c2a38 , n282624 );
buf ( R_149c9_132f4fa8 , n282628 );
buf ( R_10aae_1207c558 , n282635 );
buf ( R_13aad_11541a38 , n282641 );
buf ( R_12362_10563dd8 , n282651 );
buf ( R_5c4e_1056ced8 , n282660 );
buf ( R_130f5_1056a098 , n282672 );
buf ( R_12a7c_11cdde68 , n282684 );
buf ( R_14415_12b2a318 , n282689 );
buf ( R_1488b_13a189c8 , n282694 );
buf ( R_14062_1204cf18 , n282697 );
buf ( R_14784_11cd8508 , n282702 );
buf ( R_1032f_10570f38 , n282711 );
buf ( R_9bdf_102ee5a8 , n282722 );
buf ( R_13bf0_1331c528 , n282731 );
buf ( R_11b90_11ce0208 , n282741 );
buf ( R_149cf_13a17b68 , n282745 );
buf ( R_12021_11ce25a8 , n282754 );
buf ( R_1de_12056d98 , n282755 );
buf ( R_49_1331f4a8 , n282756 );
buf ( R_131_105ab3b8 , n282757 );
buf ( R_1462f_13794688 , n282761 );
buf ( R_10628_1203d2d8 , n282773 );
buf ( R_122bf_10570038 , n282784 );
buf ( R_11387_11540d18 , n282795 );
buf ( R_11fa6_13306308 , n282804 );
buf ( R_85b5_120819b8 , n282816 );
buf ( R_142ef_102eec88 , n282821 );
buf ( R_1434c_102f13e8 , n282826 );
buf ( R_22c_1379b708 , n282827 );
buf ( R_5c_137944a8 , n282828 );
buf ( R_e3_1203e778 , n282829 );
buf ( R_b948_1153a5f8 , n282838 );
buf ( R_e169_11cd7a68 , n282849 );
buf ( R_d051_11536ef8 , n282855 );
buf ( R_10e01_120551b8 , n282866 );
buf ( R_233_12b392d8 , n282867 );
buf ( R_68_12b283d8 , n282868 );
buf ( R_dc_13300768 , n282869 );
buf ( R_13bfb_13316a88 , n282877 );
buf ( R_10ad6_10565598 , n282887 );
buf ( R_14870_10570538 , n282892 );
buf ( R_12260_13a1b268 , n282903 );
buf ( R_d661_1265cfc8 , n282914 );
buf ( R_14572_11cd9d68 , n282919 );
buf ( R_130ff_12078318 , n282930 );
buf ( R_a98a_11cdaf88 , n282938 );
buf ( R_14978_12b321f8 , n282942 );
buf ( R_14a1a_115445f8 , n282947 );
buf ( R_14a26_13792568 , n282951 );
buf ( R_b327_12648568 , n282963 );
buf ( R_108fb_105b5e58 , n282973 );
buf ( R_1440d_11544238 , n282979 );
buf ( R_10cff_13a1dc48 , n282990 );
buf ( R_139ae_11cd8b48 , n282998 );
buf ( R_14338_11cda808 , n283003 );
buf ( R_106b3_13a16088 , n283013 );
buf ( R_c4f8_11ce12e8 , n283023 );
buf ( R_215_1265b948 , n283024 );
buf ( R_fa_133070c8 , n283025 );
buf ( R_11b68_1264ec88 , n283036 );
buf ( R_129b1_1056f098 , n283048 );
buf ( R_13670_10564558 , n283054 );
buf ( R_1439c_11cdd148 , n283064 );
buf ( R_107e6_11cdbc08 , n283074 );
buf ( R_f279_13a1acc8 , n283086 );
buf ( R_12ed9_102edf68 , n283099 );
buf ( R_12bc1_13a1f048 , n283110 );
buf ( R_13b19_12b2ba38 , n283118 );
buf ( R_e361_120812d8 , n283129 );
buf ( R_bef9_11ce0528 , n283137 );
buf ( R_13ce8_120793f8 , n283145 );
buf ( R_a235_12084a78 , n283154 );
buf ( R_14521_1264f228 , n283158 );
buf ( R_13cad_13a1edc8 , n283165 );
buf ( R_148af_11540098 , n283170 );
buf ( R_10968_13304968 , n283179 );
buf ( R_13fcb_102f0c68 , n283186 );
buf ( R_11645_13304e68 , n283198 );
buf ( R_bf09_1056b498 , n283204 );
buf ( R_12553_13310308 , n283214 );
buf ( R_145d5_132fa228 , n283218 );
buf ( R_146a2_1207bf18 , n283222 );
buf ( R_136fc_12076018 , n283231 );
buf ( R_149a2_1264d1a8 , n283236 );
buf ( R_12b9a_13a14968 , n283249 );
buf ( R_137cc_10569af8 , n283256 );
buf ( R_c5ef_12081238 , n283279 );
buf ( R_1184d_11cd9188 , n283288 );
buf ( R_13c8f_102ed568 , n283297 );
buf ( R_109bf_1379c248 , n283306 );
buf ( R_14326_13301528 , n283317 );
buf ( R_11123_12045258 , n283327 );
buf ( R_e197_11ce3228 , n283339 );
buf ( R_172_126656c8 , n283340 );
buf ( R_19d_132ffb88 , n283341 );
buf ( R_c306_f8c5418 , n283354 );
buf ( R_b5_133157c8 , n283355 );
buf ( R_13902_13799ae8 , n283363 );
buf ( R_14348_1056c398 , n283368 );
buf ( R_1457b_102f5628 , n283373 );
buf ( R_14766_105674d8 , n283377 );
buf ( R_d2c1_12036e38 , n283388 );
buf ( R_1f6_1330dce8 , n283389 );
buf ( R_10c28_12080e78 , n283398 );
buf ( R_119_133166c8 , n283399 );
buf ( R_1300e_12646bc8 , n283405 );
buf ( R_13129_10567b18 , n283417 );
buf ( R_1394d_1056f318 , n283425 );
buf ( R_14846_13798b48 , n283429 );
buf ( R_146cf_1379e868 , n283434 );
buf ( R_10019_11542118 , n283445 );
buf ( R_fb35_132fb4e8 , n283457 );
buf ( R_11a23_126506c8 , n283465 );
buf ( R_9aae_1056dbf8 , n283476 );
buf ( R_14468_1264aea8 , n283481 );
buf ( R_7aaf_f8c22b8 , n283490 );
buf ( R_b5af_1264e508 , n283511 );
buf ( R_13f11_11cd7b08 , n283518 );
buf ( R_e6c6_12075cf8 , n283530 );
buf ( R_14374_102f0768 , n283537 );
buf ( R_14605_13a182e8 , n283541 );
buf ( R_13de4_102f94a8 , n283552 );
buf ( R_102c2_1264ed28 , n283574 );
buf ( R_91_13799548 , n283575 );
buf ( R_135f5_11cda4e8 , n283583 );
buf ( R_14807_1331e288 , n283588 );
buf ( R_14a08_11cdc388 , n283592 );
buf ( R_cb44_12b3ee18 , n283604 );
buf ( R_13a63_11544198 , n283636 );
buf ( R_109ca_1264cd48 , n283647 );
buf ( R_12e41_10569198 , n283659 );
buf ( R_e46a_13a181a8 , n283671 );
buf ( R_12963_13a1afe8 , n283683 );
buf ( R_14a5a_12b42158 , n283687 );
buf ( R_13e38_1207efd8 , n283699 );
buf ( R_144ea_1264f5e8 , n283703 );
buf ( R_11668_137a1d88 , n283726 );
buf ( R_13ec7_11540318 , n283736 );
buf ( R_ff67_13799688 , n283747 );
buf ( R_13b27_102eb588 , n283756 );
buf ( R_fa2a_1056e0f8 , n283767 );
buf ( R_145a5_132f4dc8 , n283771 );
buf ( R_14060_13a15ae8 , n283774 );
buf ( R_164_12b27118 , n283775 );
buf ( R_104d9_120779b8 , n283786 );
buf ( R_1ab_f8c2998 , n283787 );
buf ( R_23c_13319328 , n283788 );
buf ( R_bbdf_133063a8 , n283795 );
buf ( R_d3_12659968 , n283796 );
buf ( R_cc7b_13a1b128 , n283807 );
buf ( R_12ffe_1331cd48 , n283816 );
buf ( R_1323e_126561c8 , n283828 );
buf ( R_1207f_133190a8 , n283839 );
buf ( R_10f99_126549a8 , n283850 );
buf ( R_913d_12646b28 , n283861 );
buf ( R_c3ee_102f6848 , n283873 );
buf ( R_13b12_13a1a728 , n283882 );
buf ( R_10a0c_11cdf1c8 , n283893 );
buf ( R_13974_13a19008 , n283900 );
buf ( R_13602_126635a8 , n283907 );
buf ( R_124e1_11cdb668 , n283918 );
buf ( R_142d7_12b30d58 , n283923 );
buf ( R_14960_105b5598 , n283927 );
buf ( R_f86d_120385f8 , n283940 );
buf ( R_148a0_12b38ab8 , n283945 );
buf ( R_e63f_f8cb9f8 , n283957 );
buf ( R_12741_105642d8 , n283968 );
buf ( R_684e_1056aa98 , n283974 );
buf ( R_13b04_12081558 , n283982 );
buf ( R_1453f_11ce2328 , n283987 );
buf ( R_148b5_1207f898 , n283991 );
buf ( R_1499c_12080658 , n283996 );
buf ( R_128e2_12647668 , n284005 );
buf ( R_13345_11ce0988 , n284016 );
buf ( R_cd4f_102f2f68 , n284026 );
buf ( R_13dd3_1204cd38 , n284034 );
buf ( R_13ea4_11ce0708 , n284046 );
buf ( R_f16b_11cda448 , n284058 );
buf ( R_139fe_1153e5b8 , n284068 );
buf ( R_12eed_102ee1e8 , n284078 );
buf ( R_13479_13306b28 , n284090 );
buf ( R_1135b_1056d158 , n284101 );
buf ( R_131a5_1153dc58 , n284109 );
buf ( R_14744_1264b3a8 , n284113 );
buf ( R_144c6_1056d5b8 , n284117 );
buf ( R_13109_f8c4798 , n284128 );
buf ( R_137bb_10564058 , n284137 );
buf ( R_146db_1056a818 , n284141 );
buf ( R_119c2_13a1a548 , n284153 );
buf ( R_eb5e_1056d018 , n284164 );
buf ( R_b0d7_1153e3d8 , n284176 );
buf ( R_13b9e_12083038 , n284184 );
buf ( R_1116a_13a15868 , n284195 );
buf ( R_12a65_10564c38 , n284206 );
buf ( R_14969_11cdb2a8 , n284210 );
buf ( R_1464d_12075618 , n284215 );
buf ( R_e3c5_12080a18 , n284227 );
buf ( R_1469c_120511f8 , n284231 );
buf ( R_d50f_12663828 , n284243 );
buf ( R_137f0_12079358 , n284249 );
buf ( R_11593_1207a258 , n284259 );
buf ( R_14350_1207d8b8 , n284264 );
buf ( R_cbe2_11536a98 , n284275 );
buf ( R_110ed_10563d38 , n284285 );
buf ( R_1125d_102f86e8 , n284293 );
buf ( R_13c09_11ce4268 , n284301 );
buf ( R_135fc_13795948 , n284309 );
buf ( R_14557_11cdcec8 , n284313 );
buf ( R_112_13312248 , n284314 );
buf ( R_1fd_133221a8 , n284315 );
buf ( R_9e_11539838 , n284316 );
buf ( R_143b2_11cddd28 , n284321 );
buf ( R_12fec_102efea8 , n284331 );
buf ( R_c4d7_13a1f408 , n284342 );
buf ( R_1398e_13320bc8 , n284348 );
buf ( R_12894_11ce1428 , n284359 );
buf ( R_b6f4_102f9ea8 , n284369 );
buf ( R_fcb3_12649be8 , n284380 );
buf ( R_12375_1207edf8 , n284391 );
buf ( R_146b1_102ed248 , n284396 );
buf ( R_11b11_11545818 , n284406 );
buf ( R_58_13317a28 , n284407 );
buf ( R_73_12b3e0f8 , n284408 );
buf ( R_bd7c_11ce2be8 , n284415 );
buf ( R_12fd8_10565278 , n284425 );
buf ( R_14876_12054678 , n284430 );
buf ( R_138da_1153dbb8 , n284436 );
buf ( R_14825_12647168 , n284440 );
buf ( R_14a4d_12646ee8 , n284444 );
buf ( R_124_1203edb8 , n284445 );
buf ( R_15a_f8c6958 , n284446 );
buf ( R_1b5_1331afe8 , n284447 );
buf ( R_1eb_12038d78 , n284448 );
buf ( R_1475d_11546038 , n284453 );
buf ( R_171_105aa5f8 , n284454 );
buf ( R_106ea_102f6528 , n284466 );
buf ( R_19e_1331e788 , n284467 );
buf ( R_11a86_1204ffd8 , n284487 );
buf ( R_fad7_102f5ee8 , n284500 );
buf ( R_e21e_1056b7b8 , n284512 );
buf ( R_12933_11cd7c48 , n284523 );
buf ( R_6c_12040938 , n284524 );
buf ( R_99_12b27618 , n284525 );
buf ( R_1353d_1153d9d8 , n284533 );
buf ( R_b283_1330acc8 , n284542 );
buf ( R_143ae_13a1cca8 , n284547 );
buf ( R_14801_11540c78 , n284551 );
buf ( R_149e7_10568298 , n284555 );
buf ( R_14708_1203c018 , n284560 );
buf ( R_14450_13a17028 , n284565 );
buf ( R_128_12b43b98 , n284566 );
buf ( R_145_1265aa48 , n284567 );
buf ( R_1ca_1265ff48 , n284568 );
buf ( R_1e7_12b3d798 , n284569 );
buf ( R_7741_13a16128 , n284579 );
buf ( R_da39_12b40718 , n284591 );
buf ( R_e38d_12651168 , n284603 );
buf ( R_12fc4_11544878 , n284614 );
buf ( R_145e7_11544058 , n284618 );
buf ( R_1465f_105676b8 , n284623 );
buf ( R_10fc1_12078638 , n284632 );
buf ( R_704f_11ce4da8 , n284640 );
buf ( R_13a8d_13318108 , n284646 );
buf ( R_145c3_1264da68 , n284650 );
buf ( R_faad_13a1fd68 , n284661 );
buf ( R_12738_10570678 , n284670 );
buf ( R_11935_13a1ff48 , n284680 );
buf ( R_11720_1330eaa8 , n284688 );
buf ( R_d16a_11ce5de8 , n284706 );
buf ( R_13e0d_13a1b4e8 , n284717 );
buf ( R_1447d_11ce3a48 , n284721 );
buf ( R_152_12b3c4d8 , n284722 );
buf ( R_105ba_13306bc8 , n284734 );
buf ( R_b1aa_12649468 , n284740 );
buf ( R_1bd_12653be8 , n284741 );
buf ( R_14a50_13a161c8 , n284746 );
buf ( R_13a83_10567a78 , n284752 );
buf ( R_123c2_13797108 , n284758 );
buf ( R_144b7_13305d68 , n284762 );
buf ( R_13814_137926a8 , n284768 );
buf ( R_12cbd_13a14328 , n284778 );
buf ( R_11bab_120768d8 , n284786 );
buf ( R_c07e_13a18b08 , n284797 );
buf ( R_142f9_11545e58 , n284802 );
buf ( R_1478a_12652928 , n284806 );
buf ( R_14a3b_11ce2d28 , n284810 );
buf ( R_c3a2_13a19508 , n284821 );
buf ( R_aa_126535a8 , n284822 );
buf ( R_146e7_10566538 , n284827 );
buf ( R_138fb_12082778 , n284836 );
buf ( R_13988_133186a8 , n284844 );
buf ( R_13c43_1264cca8 , n284850 );
buf ( R_14590_132f3b08 , n284854 );
buf ( R_110cf_137940e8 , n284863 );
buf ( R_13326_12648d88 , n284874 );
buf ( R_13153_10567118 , n284885 );
buf ( R_1405e_f8c95b8 , n284888 );
buf ( R_1051f_13793b48 , n284913 );
buf ( R_f518_12075bb8 , n284925 );
buf ( R_143a2_12079038 , n284932 );
buf ( R_147a8_12657de8 , n284936 );
buf ( R_13cb3_102f6fc8 , n284943 );
buf ( R_10c3d_f8c5b98 , n284952 );
buf ( R_e7ab_1264f7c8 , n284963 );
buf ( R_13449_12077378 , n284976 );
buf ( R_14403_12b29418 , n284981 );
buf ( R_148b2_132fc708 , n284986 );
buf ( R_1468f_10562cf8 , n284990 );
buf ( R_f7_13309828 , n284991 );
buf ( R_13f54_102f4e08 , n284999 );
buf ( R_218_12050258 , n285000 );
buf ( R_83_1379cd88 , n285001 );
buf ( R_12f16_137a0b68 , n285010 );
buf ( R_10598_102ead68 , n285018 );
buf ( R_10365_12051478 , n285028 );
buf ( R_13ab4_13a12ca8 , n285036 );
buf ( R_13393_10568a18 , n285048 );
buf ( R_13683_1207cf58 , n285055 );
buf ( R_13a_105ac2b8 , n285056 );
buf ( R_127d5_11cdf268 , n285068 );
buf ( R_11917_11ce1248 , n285079 );
buf ( R_1d5_1265e468 , n285080 );
buf ( R_12e98_1204e778 , n285087 );
buf ( R_b3_12655ea8 , n285088 );
buf ( R_149cc_10564cd8 , n285093 );
buf ( R_134d9_10565f98 , n285103 );
buf ( R_fd0b_102ec488 , n285115 );
buf ( R_af25_133136a8 , n285127 );
buf ( R_11948_12b288d8 , n285138 );
buf ( R_149c6_1207b018 , n285142 );
buf ( R_14b_12b28a18 , n285143 );
buf ( R_1c4_12652e28 , n285144 );
buf ( R_10199_13a1f368 , n285155 );
buf ( R_80_12055438 , n285156 );
buf ( R_10b70_f8cd438 , n285165 );
buf ( R_10cdf_115401d8 , n285175 );
buf ( R_11a66_1207dc78 , n285183 );
buf ( R_132fc_13307708 , n285195 );
buf ( R_8c7b_12076b58 , n285206 );
buf ( R_1495a_1207a2f8 , n285210 );
buf ( R_1201a_10570218 , n285222 );
buf ( R_132d6_11ce0348 , n285233 );
buf ( R_14963_13304be8 , n285237 );
buf ( R_1285e_11545c78 , n285247 );
buf ( R_130de_102f58a8 , n285256 );
buf ( R_fb5f_13a1e288 , n285269 );
buf ( R_13ecf_1207c5f8 , n285278 );
buf ( R_1456f_13a1f5e8 , n285282 );
buf ( R_ea_1331a9a8 , n285283 );
buf ( R_120_12b400d8 , n285284 );
buf ( R_13eac_11ce2a08 , n285307 );
buf ( R_12568_1056b0d8 , n285318 );
buf ( R_e3ba_1207df98 , n285330 );
buf ( R_dcf2_12085298 , n285342 );
buf ( R_1ef_f8c2cb8 , n285343 );
buf ( R_225_12b3a318 , n285344 );
buf ( R_f7da_1204e9f8 , n285355 );
buf ( R_f857_13a13748 , n285366 );
buf ( R_1461a_13301988 , n285371 );
buf ( R_146b7_13a15228 , n285375 );
buf ( R_1384a_126503a8 , n285382 );
buf ( R_c8e7_105b6498 , n285391 );
buf ( R_86_137a1a68 , n285392 );
buf ( R_a3_126621a8 , n285393 );
buf ( R_f862_13a1a908 , n285405 );
buf ( R_10ab7_102f7b08 , n285415 );
buf ( R_11890_102eb308 , n285423 );
buf ( R_df3c_120774b8 , n285436 );
buf ( R_1369b_1330c2a8 , n285445 );
buf ( R_12e03_132ff368 , n285455 );
buf ( R_1356b_102f5da8 , n285466 );
buf ( R_10e42_1207e718 , n285478 );
buf ( R_10f59_f8c2c18 , n285486 );
buf ( R_127b6_12b412f8 , n285493 );
buf ( R_120e7_12b44818 , n285503 );
buf ( R_12492_1265b9e8 , n285515 );
buf ( R_10d12_13792b08 , n285523 );
buf ( R_130ae_12044b78 , n285536 );
buf ( R_13652_11ce1ce8 , n285542 );
buf ( R_117a7_12080fb8 , n285551 );
buf ( R_14674_13a13ba8 , n285555 );
buf ( R_11306_11540638 , n285566 );
buf ( R_d5_126617a8 , n285567 );
buf ( R_de_1265ce88 , n285568 );
buf ( R_12c_1379b488 , n285569 );
buf ( R_135_f8c6f98 , n285570 );
buf ( R_1da_12664b88 , n285571 );
buf ( R_1e3_1153c498 , n285572 );
buf ( R_122dd_13a1b6c8 , n285582 );
buf ( R_231_1379a6c8 , n285583 );
buf ( R_23a_12660b28 , n285584 );
buf ( R_1240e_13a150e8 , n285594 );
buf ( R_14686_13a137e8 , n285598 );
buf ( R_146c6_f8cf918 , n285603 );
buf ( R_13f5b_1207c738 , n285611 );
buf ( R_ebb7_102efd68 , n285622 );
buf ( R_1447a_105697d8 , n285627 );
buf ( R_13c95_12650ee8 , n285634 );
buf ( R_11de0_12083cb8 , n285646 );
buf ( R_11552_12648c48 , n285658 );
buf ( R_11cb2_1207ab18 , n285669 );
buf ( R_14849_11ce0028 , n285673 );
buf ( R_13f45_13a134c8 , n285681 );
buf ( R_13726_12084f78 , n285688 );
buf ( R_121f2_102f30a8 , n285699 );
buf ( R_ef_1379b0c8 , n285700 );
buf ( R_163_12b38a18 , n285701 );
buf ( R_1ac_12b29558 , n285702 );
buf ( R_220_12b25638 , n285703 );
buf ( R_14623_13a12a28 , n285707 );
buf ( R_1393a_11ce3408 , n285715 );
buf ( R_139ea_11cd8828 , n285722 );
buf ( R_cf49_11541718 , n285733 );
buf ( R_b889_1056a458 , n285743 );
buf ( R_1349f_1204fdf8 , n285754 );
buf ( R_170_120440d8 , n285755 );
buf ( R_19f_133087e8 , n285756 );
buf ( R_a9d8_102f22e8 , n285769 );
buf ( R_7d_12660308 , n285770 );
buf ( R_1460b_10569a58 , n285774 );
buf ( R_11983_13318568 , n285782 );
buf ( R_a6e4_13314648 , n285794 );
buf ( R_144b1_1207b478 , n285798 );
buf ( R_14614_12664f48 , n285802 );
buf ( R_139d7_132fda68 , n285810 );
buf ( R_ec64_11ce6248 , n285823 );
buf ( R_12d32_115454f8 , n285834 );
buf ( R_82bb_1204a678 , n285841 );
buf ( R_1472c_13a139c8 , n285846 );
buf ( R_144f7_10565e58 , n285850 );
buf ( R_10dad_12082f98 , n285860 );
buf ( R_b05c_1330b4e8 , n285872 );
buf ( R_13ef1_105714d8 , n285882 );
buf ( R_14635_12b3b038 , n285887 );
buf ( R_117b5_1056fdb8 , n285900 );
buf ( R_14692_11cdf128 , n285904 );
buf ( R_13f_1203dd78 , n285905 );
buf ( R_1055c_105672f8 , n285918 );
buf ( R_1d0_12040258 , n285919 );
buf ( R_13aba_1265cde8 , n285926 );
buf ( R_131e1_102f2ec8 , n285937 );
buf ( R_eb07_1153ef18 , n285950 );
buf ( R_9c9a_1056c578 , n285961 );
buf ( R_10605_11545d18 , n285970 );
buf ( R_13a97_12079218 , n285976 );
buf ( R_1331b_102efc28 , n285987 );
buf ( R_14879_11ce58e8 , n285991 );
buf ( R_14996_102eb3a8 , n285995 );
buf ( R_1405c_11ce34a8 , n285998 );
buf ( R_14945_1056e238 , n286002 );
buf ( R_b65f_11cdba28 , n286011 );
buf ( R_13f3e_13a1e508 , n286020 );
buf ( R_dbc0_132fb9e8 , n286031 );
buf ( R_1351c_13797068 , n286042 );
buf ( R_14804_120788b8 , n286047 );
buf ( R_14a0b_133206c8 , n286051 );
buf ( R_89_126595a8 , n286052 );
buf ( R_13c33_11ce3688 , n286059 );
buf ( R_4f_12b44d18 , n286060 );
buf ( R_cb5a_12b256d8 , n286072 );
buf ( R_13b85_10571258 , n286079 );
buf ( R_138f4_1330a9a8 , n286085 );
buf ( R_ee1a_1264fae8 , n286097 );
buf ( R_10411_102f8828 , n286109 );
buf ( R_14331_1056be98 , n286114 );
buf ( R_14717_1153a378 , n286119 );
buf ( R_94_1330ee68 , n286120 );
buf ( R_e5_1153cfd8 , n286121 );
buf ( R_22a_12b43698 , n286122 );
buf ( R_cba1_13a16e48 , n286141 );
buf ( R_129d1_12047978 , n286151 );
buf ( R_143d8_11cdc2e8 , n286158 );
buf ( R_13070_1264b268 , n286168 );
buf ( R_12915_1056d518 , n286180 );
buf ( R_12942_11cdd0a8 , n286187 );
buf ( R_145a8_12662608 , n286191 );
buf ( R_fda2_1264e328 , n286202 );
buf ( R_ee25_13a16588 , n286213 );
buf ( R_13a1f_11cde2c8 , n286221 );
buf ( R_1432d_11cdddc8 , n286226 );
buf ( R_13be3_12036bb8 , n286232 );
buf ( R_fe10_13a14468 , n286243 );
buf ( R_12610_1204bcf8 , n286253 );
buf ( R_13701_11cdc608 , n286259 );
buf ( R_12597_105711b8 , n286270 );
buf ( R_1441d_12035d58 , n286275 );
buf ( R_1443c_137979c8 , n286281 );
buf ( R_139a7_11ce70a8 , n286287 );
buf ( R_13ad3_1056bdf8 , n286296 );
buf ( R_143e0_102efcc8 , n286301 );
buf ( R_147cc_13315ae8 , n286305 );
buf ( R_1444b_11cdad08 , n286310 );
buf ( R_12631_12036c58 , n286322 );
buf ( R_13dda_102f4fe8 , n286329 );
buf ( R_efd_13a14fa8 , n286332 );
buf ( R_14954_12054358 , n286336 );
buf ( R_1287f_115422f8 , n286346 );
buf ( R_1169f_102f8968 , n286355 );
buf ( R_13a2b_1264b628 , n286367 );
buf ( R_11285_102f9e08 , n286377 );
buf ( R_12548_1056ce38 , n286388 );
buf ( R_1173e_12649fa8 , n286396 );
buf ( R_10b51_13a18a68 , n286403 );
buf ( R_148ca_13a18c48 , n286408 );
buf ( R_12c82_102f0448 , n286419 );
buf ( R_13b79_11543d38 , n286425 );
buf ( R_14057_f8cd618 , n286428 );
buf ( R_a2e4_1056c618 , n286441 );
buf ( R_101e6_1330c7a8 , n286452 );
buf ( R_13a56_f8c0a58 , n286459 );
buf ( R_d6bc_13a1ca28 , n286471 );
buf ( R_4a_1265e648 , n286472 );
buf ( R_115_13316c68 , n286473 );
buf ( R_1224c_12b3d478 , n286484 );
buf ( R_1fa_1265d388 , n286485 );
buf ( R_eeda_11cd81e8 , n286498 );
buf ( R_1455d_11cd9fe8 , n286503 );
buf ( R_1402e_1264dc48 , n286512 );
buf ( R_c753_12039098 , n286523 );
buf ( R_1283c_13a1da68 , n286534 );
buf ( R_aeda_13a1d6a8 , n286545 );
buf ( R_14939_1379f448 , n286549 );
buf ( R_14a20_13a13e28 , n286553 );
buf ( R_13a9d_12081698 , n286560 );
buf ( R_117c0_11ce3e08 , n286569 );
buf ( R_114e1_132f28e8 , n286575 );
buf ( R_1476f_132fb768 , n286580 );
buf ( n25318 , RI19a22f70_2797);
not ( n25319 , n25318 );
not ( n25320 , RI1754a798_67);
nand ( n25321 , n25319 , n25320 );
buf ( n25322 , RI19ad04a8_2209);
buf ( n25323 , RI19a23e70_2789);
buf ( n25324 , n25323 );
nor ( n25325 , n25322 , n25324 );
not ( n25326 , RI1754c610_2);
nand ( n25327 , n25321 , n25325 , n25326 );
buf ( n25328 , n25327 );
not ( n25329 , RI19a23510_2794);
or ( n25330 , n25328 , n25329 );
not ( n25331 , n25325 );
not ( n25332 , n25321 );
or ( n25333 , n25331 , n25332 );
nand ( n25334 , n25333 , n25326 );
buf ( n25335 , n25334 );
buf ( n25336 , n25335 );
not ( n25337 , RI19a859b8_2755);
or ( n25338 , n25336 , n25337 );
nand ( n25339 , n25330 , n25338 );
buf ( n25340 , n25339 );
buf ( n25341 , RI17534808_603);
not ( n25342 , n25341 );
buf ( n25343 , RI173f4d68_1562);
not ( n25344 , n25343 );
not ( n25345 , RI173ac078_1917);
not ( n25346 , n25345 );
or ( n25347 , n25344 , n25346 );
not ( n25348 , RI173f4d68_1562);
buf ( n25349 , RI173ac078_1917);
nand ( n25350 , n25348 , n25349 );
nand ( n25351 , n25347 , n25350 );
not ( n25352 , RI17516358_697);
and ( n25353 , n25351 , n25352 );
not ( n25354 , n25351 );
buf ( n25355 , RI17516358_697);
and ( n25356 , n25354 , n25355 );
nor ( n25357 , n25353 , n25356 );
buf ( n25358 , RI1753aa78_586);
not ( n25359 , n25358 );
nand ( n25360 , n25359 , n25323 );
not ( n25361 , n25360 );
buf ( n25362 , n25361 );
buf ( n25363 , n25362 );
buf ( n25364 , n25363 );
buf ( n25365 , RI19aad828_2471);
nand ( n25366 , n25364 , n25365 );
buf ( n25367 , RI17491398_1028);
and ( n25368 , n25366 , n25367 );
not ( n25369 , n25366 );
not ( n25370 , RI17491398_1028);
and ( n25371 , n25369 , n25370 );
nor ( n25372 , n25368 , n25371 );
xor ( n25373 , n25357 , n25372 );
buf ( n25374 , n25361 );
buf ( n25375 , n25374 );
buf ( n25376 , n25375 );
buf ( n25377 , RI19ac0a40_2326);
nand ( n25378 , n25376 , n25377 );
not ( n25379 , RI1751df18_673);
and ( n25380 , n25378 , n25379 );
not ( n25381 , n25378 );
buf ( n25382 , RI1751df18_673);
and ( n25383 , n25381 , n25382 );
nor ( n25384 , n25380 , n25383 );
xnor ( n25385 , n25373 , n25384 );
not ( n25386 , n25385 );
or ( n25387 , n25342 , n25386 );
or ( n25388 , n25385 , n25341 );
nand ( n25389 , n25387 , n25388 );
buf ( n25390 , RI173c95b0_1774);
not ( n25391 , n25390 );
not ( n25392 , RI17340030_2129);
not ( n25393 , n25392 );
or ( n25394 , n25391 , n25393 );
not ( n25395 , RI173c95b0_1774);
buf ( n25396 , RI17340030_2129);
nand ( n25397 , n25395 , n25396 );
nand ( n25398 , n25394 , n25397 );
not ( n25399 , RI174125e8_1418);
and ( n25400 , n25398 , n25399 );
not ( n25401 , n25398 );
buf ( n25402 , RI174125e8_1418);
and ( n25403 , n25401 , n25402 );
nor ( n25404 , n25400 , n25403 );
buf ( n25405 , n25363 );
buf ( n25406 , RI19a8ffa8_2683);
nand ( n25407 , n25405 , n25406 );
buf ( n25408 , RI17465bf8_1240);
and ( n25409 , n25407 , n25408 );
not ( n25410 , n25407 );
not ( n25411 , RI17465bf8_1240);
and ( n25412 , n25410 , n25411 );
nor ( n25413 , n25409 , n25412 );
xor ( n25414 , n25404 , n25413 );
buf ( n25415 , n25361 );
buf ( n25416 , n25415 );
buf ( n25417 , RI19ac0680_2328);
nand ( n25418 , n25416 , n25417 );
buf ( n25419 , RI174ae8d0_885);
and ( n25420 , n25418 , n25419 );
not ( n25421 , n25418 );
not ( n25422 , RI174ae8d0_885);
and ( n25423 , n25421 , n25422 );
nor ( n25424 , n25420 , n25423 );
xor ( n25425 , n25414 , n25424 );
buf ( n25426 , n25425 );
and ( n25427 , n25389 , n25426 );
not ( n25428 , n25389 );
not ( n25429 , n25426 );
and ( n25430 , n25428 , n25429 );
nor ( n25431 , n25427 , n25430 );
not ( n25432 , n25431 );
not ( n25433 , n25432 );
buf ( n25434 , RI1733be90_2149);
not ( n25435 , n25434 );
buf ( n25436 , RI173c9268_1775);
buf ( n25437 , RI173ff808_1510);
not ( n25438 , n25437 );
not ( n25439 , RI173b67d0_1866);
not ( n25440 , n25439 );
or ( n25441 , n25438 , n25440 );
not ( n25442 , RI173ff808_1510);
buf ( n25443 , RI173b67d0_1866);
nand ( n25444 , n25442 , n25443 );
nand ( n25445 , n25441 , n25444 );
xor ( n25446 , n25436 , n25445 );
buf ( n25447 , RI1752e610_622);
not ( n25448 , RI1749baf0_977);
xor ( n25449 , n25447 , n25448 );
buf ( n25450 , n25361 );
buf ( n25451 , n25450 );
buf ( n25452 , n25451 );
buf ( n25453 , RI19ab9a38_2383);
nand ( n25454 , n25452 , n25453 );
xnor ( n25455 , n25449 , n25454 );
xnor ( n25456 , n25446 , n25455 );
not ( n25457 , n25456 );
not ( n25458 , n25457 );
or ( n25459 , n25435 , n25458 );
not ( n25460 , n25434 );
nand ( n25461 , n25460 , n25456 );
nand ( n25462 , n25459 , n25461 );
buf ( n25463 , RI173d4068_1722);
not ( n25464 , n25463 );
not ( n25465 , RI1738b378_2077);
not ( n25466 , n25465 );
or ( n25467 , n25464 , n25466 );
not ( n25468 , RI173d4068_1722);
buf ( n25469 , RI1738b378_2077);
nand ( n25470 , n25468 , n25469 );
nand ( n25471 , n25467 , n25470 );
buf ( n25472 , RI1744bb40_1367);
and ( n25473 , n25471 , n25472 );
not ( n25474 , n25471 );
not ( n25475 , RI1744bb40_1367);
and ( n25476 , n25474 , n25475 );
nor ( n25477 , n25473 , n25476 );
not ( n25478 , n25477 );
buf ( n25479 , n25415 );
buf ( n25480 , RI19a9c5f0_2595);
nand ( n25481 , n25479 , n25480 );
buf ( n25482 , RI17470350_1189);
and ( n25483 , n25481 , n25482 );
not ( n25484 , n25481 );
not ( n25485 , RI17470350_1189);
and ( n25486 , n25484 , n25485 );
nor ( n25487 , n25483 , n25486 );
xor ( n25488 , n25478 , n25487 );
buf ( n25489 , n25361 );
buf ( n25490 , n25489 );
buf ( n25491 , n25490 );
buf ( n25492 , RI19acb828_2243);
nand ( n25493 , n25491 , n25492 );
buf ( n25494 , RI174b9460_834);
and ( n25495 , n25493 , n25494 );
not ( n25496 , n25493 );
not ( n25497 , RI174b9460_834);
and ( n25498 , n25496 , n25497 );
nor ( n25499 , n25495 , n25498 );
not ( n25500 , n25499 );
xnor ( n25501 , n25488 , n25500 );
not ( n25502 , n25501 );
not ( n25503 , n25502 );
and ( n25504 , n25462 , n25503 );
not ( n25505 , n25462 );
xor ( n25506 , n25477 , n25499 );
not ( n25507 , n25487 );
xnor ( n25508 , n25506 , n25507 );
buf ( n25509 , n25508 );
and ( n25510 , n25505 , n25509 );
nor ( n25511 , n25504 , n25510 );
buf ( n25512 , RI173dd410_1677);
not ( n25513 , n25512 );
buf ( n25514 , RI173cee48_1747);
not ( n25515 , n25514 );
not ( n25516 , RI17345580_2103);
not ( n25517 , n25516 );
or ( n25518 , n25515 , n25517 );
not ( n25519 , RI173cee48_1747);
buf ( n25520 , RI17345580_2103);
nand ( n25521 , n25519 , n25520 );
nand ( n25522 , n25518 , n25521 );
not ( n25523 , RI17446938_1392);
and ( n25524 , n25522 , n25523 );
not ( n25525 , n25522 );
buf ( n25526 , RI17446938_1392);
and ( n25527 , n25525 , n25526 );
nor ( n25528 , n25524 , n25527 );
buf ( n25529 , n25415 );
buf ( n25530 , RI19a8c498_2709);
nand ( n25531 , n25529 , n25530 );
not ( n25532 , RI1746b148_1214);
and ( n25533 , n25531 , n25532 );
not ( n25534 , n25531 );
buf ( n25535 , RI1746b148_1214);
and ( n25536 , n25534 , n25535 );
nor ( n25537 , n25533 , n25536 );
xor ( n25538 , n25528 , n25537 );
buf ( n25539 , n25362 );
buf ( n25540 , n25539 );
buf ( n25541 , RI19abd890_2354);
nand ( n25542 , n25540 , n25541 );
not ( n25543 , RI174b3e20_859);
and ( n25544 , n25542 , n25543 );
not ( n25545 , n25542 );
buf ( n25546 , RI174b3e20_859);
and ( n25547 , n25545 , n25546 );
nor ( n25548 , n25544 , n25547 );
xnor ( n25549 , n25538 , n25548 );
not ( n25550 , n25549 );
not ( n25551 , n25550 );
or ( n25552 , n25513 , n25551 );
not ( n25553 , n25549 );
or ( n25554 , n25553 , n25512 );
nand ( n25555 , n25552 , n25554 );
buf ( n25556 , RI173ec398_1604);
not ( n25557 , n25556 );
not ( n25558 , RI173a36a8_1959);
not ( n25559 , n25558 );
or ( n25560 , n25557 , n25559 );
not ( n25561 , RI173ec398_1604);
buf ( n25562 , RI173a36a8_1959);
nand ( n25563 , n25561 , n25562 );
nand ( n25564 , n25560 , n25563 );
not ( n25565 , RI1747e900_1119);
and ( n25566 , n25564 , n25565 );
not ( n25567 , n25564 );
buf ( n25568 , RI1747e900_1119);
and ( n25569 , n25567 , n25568 );
nor ( n25570 , n25566 , n25569 );
buf ( n25571 , n25489 );
buf ( n25572 , n25571 );
buf ( n25573 , RI19acf1d0_2217);
nand ( n25574 , n25572 , n25573 );
not ( n25575 , RI17510160_716);
and ( n25576 , n25574 , n25575 );
not ( n25577 , n25574 );
buf ( n25578 , RI17510160_716);
and ( n25579 , n25577 , n25578 );
nor ( n25580 , n25576 , n25579 );
xor ( n25581 , n25570 , n25580 );
buf ( n25582 , n25362 );
buf ( n25583 , n25582 );
buf ( n25584 , RI19aa05b0_2566);
nand ( n25585 , n25583 , n25584 );
buf ( n25586 , RI17488680_1071);
and ( n25587 , n25585 , n25586 );
not ( n25588 , n25585 );
not ( n25589 , RI17488680_1071);
and ( n25590 , n25588 , n25589 );
nor ( n25591 , n25587 , n25590 );
xor ( n25592 , n25581 , n25591 );
not ( n25593 , n25592 );
buf ( n25594 , n25593 );
and ( n25595 , n25555 , n25594 );
not ( n25596 , n25555 );
not ( n25597 , n25592 );
not ( n25598 , n25597 );
and ( n25599 , n25596 , n25598 );
nor ( n25600 , n25595 , n25599 );
not ( n25601 , n25600 );
nand ( n25602 , n25511 , n25601 );
not ( n25603 , n25602 );
or ( n25604 , n25433 , n25603 );
or ( n25605 , n25602 , n25432 );
nand ( n25606 , n25604 , n25605 );
not ( n25607 , n25606 );
buf ( n25608 , RI173895f0_2086);
buf ( n25609 , RI1740b9a0_1451);
not ( n25610 , n25609 );
not ( n25611 , RI173c2cb0_1806);
not ( n25612 , n25611 );
or ( n25613 , n25610 , n25612 );
not ( n25614 , RI1740b9a0_1451);
buf ( n25615 , RI173c2cb0_1806);
nand ( n25616 , n25614 , n25615 );
nand ( n25617 , n25613 , n25616 );
xor ( n25618 , n25608 , n25617 );
buf ( n25619 , RI17339730_2161);
buf ( n25620 , RI174a7fd0_917);
xor ( n25621 , n25619 , n25620 );
buf ( n25622 , n25363 );
buf ( n25623 , RI19ab3138_2431);
nand ( n25624 , n25622 , n25623 );
xnor ( n25625 , n25621 , n25624 );
xnor ( n25626 , n25618 , n25625 );
not ( n25627 , n25626 );
buf ( n25628 , n25374 );
buf ( n25629 , RI19a95048_2647);
nand ( n25630 , n25628 , n25629 );
buf ( n25631 , RI1752a308_635);
and ( n25632 , n25630 , n25631 );
not ( n25633 , n25630 );
not ( n25634 , RI1752a308_635);
and ( n25635 , n25633 , n25634 );
nor ( n25636 , n25632 , n25635 );
not ( n25637 , n25636 );
not ( n25638 , n25637 );
not ( n25639 , n25638 );
buf ( n25640 , RI173ee468_1594);
not ( n25641 , n25640 );
not ( n25642 , RI173a5778_1949);
not ( n25643 , n25642 );
or ( n25644 , n25641 , n25643 );
not ( n25645 , RI173ee468_1594);
buf ( n25646 , RI173a5778_1949);
nand ( n25647 , n25645 , n25646 );
nand ( n25648 , n25644 , n25647 );
buf ( n25649 , RI17493120_1019);
and ( n25650 , n25648 , n25649 );
not ( n25651 , n25648 );
not ( n25652 , RI17493120_1019);
and ( n25653 , n25651 , n25652 );
nor ( n25654 , n25650 , n25653 );
buf ( n25655 , n25489 );
buf ( n25656 , n25655 );
buf ( n25657 , RI19a9f548_2574);
nand ( n25658 , n25656 , n25657 );
not ( n25659 , RI1748a750_1061);
and ( n25660 , n25658 , n25659 );
not ( n25661 , n25658 );
buf ( n25662 , RI1748a750_1061);
and ( n25663 , n25661 , n25662 );
nor ( n25664 , n25660 , n25663 );
xor ( n25665 , n25654 , n25664 );
buf ( n25666 , n25451 );
buf ( n25667 , RI19ace168_2224);
nand ( n25668 , n25666 , n25667 );
not ( n25669 , RI17513a18_705);
and ( n25670 , n25668 , n25669 );
not ( n25671 , n25668 );
buf ( n25672 , RI17513a18_705);
and ( n25673 , n25671 , n25672 );
nor ( n25674 , n25670 , n25673 );
xnor ( n25675 , n25665 , n25674 );
not ( n25676 , n25675 );
not ( n25677 , n25676 );
or ( n25678 , n25639 , n25677 );
or ( n25679 , n25676 , n25638 );
nand ( n25680 , n25678 , n25679 );
not ( n25681 , n25680 );
and ( n25682 , n25627 , n25681 );
not ( n25683 , n25626 );
not ( n25684 , n25683 );
and ( n25685 , n25684 , n25680 );
nor ( n25686 , n25682 , n25685 );
buf ( n25687 , RI173cd750_1754);
not ( n25688 , n25687 );
not ( n25689 , RI173441d0_2109);
not ( n25690 , n25689 );
or ( n25691 , n25688 , n25690 );
not ( n25692 , RI173cd750_1754);
buf ( n25693 , RI173441d0_2109);
nand ( n25694 , n25692 , n25693 );
nand ( n25695 , n25691 , n25694 );
not ( n25696 , RI17445588_1398);
and ( n25697 , n25695 , n25696 );
not ( n25698 , n25695 );
buf ( n25699 , RI17445588_1398);
and ( n25700 , n25698 , n25699 );
nor ( n25701 , n25697 , n25700 );
buf ( n25702 , RI19a8dfc8_2697);
nand ( n25703 , n25451 , n25702 );
not ( n25704 , RI17469d98_1220);
and ( n25705 , n25703 , n25704 );
not ( n25706 , n25703 );
buf ( n25707 , RI17469d98_1220);
and ( n25708 , n25706 , n25707 );
nor ( n25709 , n25705 , n25708 );
xor ( n25710 , n25701 , n25709 );
buf ( n25711 , n25582 );
buf ( n25712 , n25711 );
buf ( n25713 , RI19abeda8_2342);
nand ( n25714 , n25712 , n25713 );
not ( n25715 , RI174b2a70_865);
and ( n25716 , n25714 , n25715 );
not ( n25717 , n25714 );
buf ( n25718 , RI174b2a70_865);
and ( n25719 , n25717 , n25718 );
nor ( n25720 , n25716 , n25719 );
xnor ( n25721 , n25710 , n25720 );
not ( n25722 , n25721 );
not ( n25723 , n25722 );
buf ( n25724 , RI173bee58_1825);
not ( n25725 , n25724 );
buf ( n25726 , RI173f9250_1541);
not ( n25727 , n25726 );
not ( n25728 , RI173b0560_1896);
not ( n25729 , n25728 );
or ( n25730 , n25727 , n25729 );
not ( n25731 , RI173f9250_1541);
buf ( n25732 , RI173b0560_1896);
nand ( n25733 , n25731 , n25732 );
nand ( n25734 , n25730 , n25733 );
buf ( n25735 , RI17389938_2085);
and ( n25736 , n25734 , n25735 );
not ( n25737 , n25734 );
not ( n25738 , RI17389938_2085);
and ( n25739 , n25737 , n25738 );
nor ( n25740 , n25736 , n25739 );
buf ( n25741 , n25362 );
buf ( n25742 , RI19aadb70_2470);
nand ( n25743 , n25741 , n25742 );
buf ( n25744 , RI17524b60_652);
and ( n25745 , n25743 , n25744 );
not ( n25746 , n25743 );
not ( n25747 , RI17524b60_652);
and ( n25748 , n25746 , n25747 );
nor ( n25749 , n25745 , n25748 );
xor ( n25750 , n25740 , n25749 );
buf ( n25751 , n25571 );
buf ( n25752 , n25751 );
buf ( n25753 , RI19aab938_2485);
nand ( n25754 , n25752 , n25753 );
buf ( n25755 , RI17495880_1007);
and ( n25756 , n25754 , n25755 );
not ( n25757 , n25754 );
not ( n25758 , RI17495880_1007);
and ( n25759 , n25757 , n25758 );
nor ( n25760 , n25756 , n25759 );
xnor ( n25761 , n25750 , n25760 );
buf ( n25762 , n25761 );
not ( n25763 , n25762 );
or ( n25764 , n25725 , n25763 );
not ( n25765 , n25761 );
not ( n25766 , n25765 );
or ( n25767 , n25766 , n25724 );
nand ( n25768 , n25764 , n25767 );
not ( n25769 , n25768 );
or ( n25770 , n25723 , n25769 );
not ( n25771 , n25721 );
not ( n25772 , n25771 );
not ( n25773 , n25772 );
or ( n25774 , n25768 , n25773 );
nand ( n25775 , n25770 , n25774 );
nand ( n25776 , n25686 , n25775 );
not ( n25777 , n25776 );
buf ( n25778 , RI173e1268_1658);
not ( n25779 , n25778 );
not ( n25780 , RI17398578_2013);
not ( n25781 , n25780 );
or ( n25782 , n25779 , n25781 );
not ( n25783 , RI173e1268_1658);
buf ( n25784 , RI17398578_2013);
nand ( n25785 , n25783 , n25784 );
nand ( n25786 , n25782 , n25785 );
buf ( n25787 , RI17459088_1302);
and ( n25788 , n25786 , n25787 );
not ( n25789 , n25786 );
not ( n25790 , RI17459088_1302);
and ( n25791 , n25789 , n25790 );
nor ( n25792 , n25788 , n25791 );
buf ( n25793 , n25490 );
buf ( n25794 , RI19a93d88_2655);
nand ( n25795 , n25793 , n25794 );
buf ( n25796 , RI1747d898_1124);
and ( n25797 , n25795 , n25796 );
not ( n25798 , n25795 );
not ( n25799 , RI1747d898_1124);
and ( n25800 , n25798 , n25799 );
nor ( n25801 , n25797 , n25800 );
xor ( n25802 , n25792 , n25801 );
buf ( n25803 , n25490 );
buf ( n25804 , RI19ac40a0_2299);
nand ( n25805 , n25803 , n25804 );
buf ( n25806 , RI174ce388_769);
and ( n25807 , n25805 , n25806 );
not ( n25808 , n25805 );
not ( n25809 , RI174ce388_769);
and ( n25810 , n25808 , n25809 );
nor ( n25811 , n25807 , n25810 );
not ( n25812 , n25811 );
xnor ( n25813 , n25802 , n25812 );
not ( n25814 , n25813 );
buf ( n25815 , RI19a9e030_2584);
nand ( n25816 , n25405 , n25815 );
buf ( n25817 , RI1748be48_1054);
and ( n25818 , n25816 , n25817 );
not ( n25819 , n25816 );
not ( n25820 , RI1748be48_1054);
and ( n25821 , n25819 , n25820 );
nor ( n25822 , n25818 , n25821 );
buf ( n25823 , n25822 );
not ( n25824 , n25823 );
and ( n25825 , n25814 , n25824 );
not ( n25826 , n25813 );
not ( n25827 , n25826 );
and ( n25828 , n25827 , n25823 );
nor ( n25829 , n25825 , n25828 );
buf ( n25830 , RI173feae8_1514);
not ( n25831 , n25830 );
not ( n25832 , RI173b5ab0_1870);
not ( n25833 , n25832 );
or ( n25834 , n25831 , n25833 );
not ( n25835 , RI173feae8_1514);
buf ( n25836 , RI173b5ab0_1870);
nand ( n25837 , n25835 , n25836 );
nand ( n25838 , n25834 , n25837 );
not ( n25839 , n25838 );
buf ( n25840 , RI173c0208_1819);
buf ( n25841 , RI19aa7c48_2511);
nand ( n25842 , n25741 , n25841 );
buf ( n25843 , RI1749add0_981);
and ( n25844 , n25842 , n25843 );
not ( n25845 , n25842 );
not ( n25846 , RI1749add0_981);
and ( n25847 , n25845 , n25846 );
nor ( n25848 , n25844 , n25847 );
xor ( n25849 , n25840 , n25848 );
buf ( n25850 , n25415 );
buf ( n25851 , n25850 );
buf ( n25852 , RI19a88e38_2732);
nand ( n25853 , n25851 , n25852 );
not ( n25854 , RI1752d170_626);
and ( n25855 , n25853 , n25854 );
not ( n25856 , n25853 );
buf ( n25857 , RI1752d170_626);
and ( n25858 , n25856 , n25857 );
nor ( n25859 , n25855 , n25858 );
xnor ( n25860 , n25849 , n25859 );
not ( n25861 , n25860 );
not ( n25862 , n25861 );
or ( n25863 , n25839 , n25862 );
not ( n25864 , n25838 );
nand ( n25865 , n25860 , n25864 );
nand ( n25866 , n25863 , n25865 );
buf ( n25867 , n25866 );
not ( n25868 , n25867 );
and ( n25869 , n25829 , n25868 );
not ( n25870 , n25829 );
and ( n25871 , n25870 , n25867 );
nor ( n25872 , n25869 , n25871 );
not ( n25873 , n25872 );
and ( n25874 , n25777 , n25873 );
and ( n25875 , n25872 , n25776 );
nor ( n25876 , n25874 , n25875 );
not ( n25877 , n25876 );
not ( n25878 , n25877 );
buf ( n25879 , n25571 );
buf ( n25880 , n25879 );
buf ( n25881 , RI19a9bfd8_2598);
nand ( n25882 , n25880 , n25881 );
not ( n25883 , RI1746f978_1192);
and ( n25884 , n25882 , n25883 );
not ( n25885 , n25882 );
buf ( n25886 , RI1746f978_1192);
and ( n25887 , n25885 , n25886 );
nor ( n25888 , n25884 , n25887 );
not ( n25889 , n25888 );
buf ( n25890 , RI1733b800_2151);
not ( n25891 , n25890 );
not ( n25892 , RI173c4d80_1796);
not ( n25893 , n25892 );
or ( n25894 , n25891 , n25893 );
not ( n25895 , RI1733b800_2151);
buf ( n25896 , RI173c4d80_1796);
nand ( n25897 , n25895 , n25896 );
nand ( n25898 , n25894 , n25897 );
not ( n25899 , RI1740da70_1441);
and ( n25900 , n25898 , n25899 );
not ( n25901 , n25898 );
buf ( n25902 , RI1740da70_1441);
and ( n25903 , n25901 , n25902 );
nor ( n25904 , n25900 , n25903 );
buf ( n25905 , RI19ac21b0_2313);
nand ( n25906 , n25803 , n25905 );
buf ( n25907 , RI174aa0a0_907);
and ( n25908 , n25906 , n25907 );
not ( n25909 , n25906 );
not ( n25910 , RI174aa0a0_907);
and ( n25911 , n25909 , n25910 );
nor ( n25912 , n25908 , n25911 );
xor ( n25913 , n25904 , n25912 );
buf ( n25914 , n25362 );
buf ( n25915 , n25914 );
buf ( n25916 , n25915 );
buf ( n25917 , RI19a91e98_2669);
nand ( n25918 , n25916 , n25917 );
not ( n25919 , RI174613c8_1262);
and ( n25920 , n25918 , n25919 );
not ( n25921 , n25918 );
buf ( n25922 , RI174613c8_1262);
and ( n25923 , n25921 , n25922 );
nor ( n25924 , n25920 , n25923 );
xnor ( n25925 , n25913 , n25924 );
not ( n25926 , n25925 );
not ( n25927 , n25926 );
not ( n25928 , n25927 );
or ( n25929 , n25889 , n25928 );
not ( n25930 , n25888 );
buf ( n25931 , n25925 );
not ( n25932 , n25931 );
nand ( n25933 , n25930 , n25932 );
nand ( n25934 , n25929 , n25933 );
buf ( n25935 , RI17399298_2009);
not ( n25936 , n25935 );
not ( n25937 , RI173e1f88_1654);
not ( n25938 , n25937 );
or ( n25939 , n25936 , n25938 );
not ( n25940 , RI17399298_2009);
buf ( n25941 , RI173e1f88_1654);
nand ( n25942 , n25940 , n25941 );
nand ( n25943 , n25939 , n25942 );
not ( n25944 , RI17459da8_1298);
and ( n25945 , n25943 , n25944 );
not ( n25946 , n25943 );
buf ( n25947 , RI17459da8_1298);
and ( n25948 , n25946 , n25947 );
nor ( n25949 , n25945 , n25948 );
buf ( n25950 , RI19a86c00_2747);
nand ( n25951 , n25914 , n25950 );
buf ( n25952 , RI174cf828_765);
and ( n25953 , n25951 , n25952 );
not ( n25954 , n25951 );
not ( n25955 , RI174cf828_765);
and ( n25956 , n25954 , n25955 );
nor ( n25957 , n25953 , n25956 );
xor ( n25958 , n25949 , n25957 );
buf ( n25959 , RI19aa5740_2526);
nand ( n25960 , n25741 , n25959 );
not ( n25961 , RI1747e5b8_1120);
xor ( n25962 , n25960 , n25961 );
xnor ( n25963 , n25958 , n25962 );
not ( n25964 , n25963 );
not ( n25965 , n25964 );
and ( n25966 , n25934 , n25965 );
not ( n25967 , n25934 );
not ( n25968 , n25949 );
not ( n25969 , n25957 );
not ( n25970 , n25962 );
or ( n25971 , n25969 , n25970 );
or ( n25972 , n25957 , n25962 );
nand ( n25973 , n25971 , n25972 );
not ( n25974 , n25973 );
or ( n25975 , n25968 , n25974 );
or ( n25976 , n25973 , n25949 );
nand ( n25977 , n25975 , n25976 );
buf ( n25978 , n25977 );
and ( n25979 , n25967 , n25978 );
nor ( n25980 , n25966 , n25979 );
not ( n25981 , n25980 );
not ( n25982 , n25981 );
buf ( n25983 , RI173fda80_1519);
buf ( n25984 , RI173bc068_1839);
not ( n25985 , n25984 );
not ( n25986 , RI17404d58_1484);
not ( n25987 , n25986 );
or ( n25988 , n25985 , n25987 );
not ( n25989 , RI173bc068_1839);
buf ( n25990 , RI17404d58_1484);
nand ( n25991 , n25989 , n25990 );
nand ( n25992 , n25988 , n25991 );
xor ( n25993 , n25983 , n25992 );
buf ( n25994 , RI17332ae8_2194);
not ( n25995 , n25994 );
buf ( n25996 , RI19ab5d48_2410);
nand ( n25997 , n25751 , n25996 );
buf ( n25998 , RI174a1040_951);
and ( n25999 , n25997 , n25998 );
not ( n26000 , n25997 );
not ( n26001 , RI174a1040_951);
and ( n26002 , n26000 , n26001 );
nor ( n26003 , n25999 , n26002 );
not ( n26004 , n26003 );
or ( n26005 , n25995 , n26004 );
or ( n26006 , n26003 , n25994 );
nand ( n26007 , n26005 , n26006 );
xnor ( n26008 , n25993 , n26007 );
buf ( n26009 , n26008 );
not ( n26010 , n26009 );
buf ( n26011 , RI173ad0e0_1912);
not ( n26012 , n26011 );
buf ( n26013 , RI173e7820_1627);
not ( n26014 , n26013 );
not ( n26015 , RI1739e7e8_1983);
not ( n26016 , n26015 );
or ( n26017 , n26014 , n26016 );
not ( n26018 , RI173e7820_1627);
buf ( n26019 , RI1739e7e8_1983);
nand ( n26020 , n26018 , n26019 );
nand ( n26021 , n26017 , n26020 );
buf ( n26022 , RI1745f2f8_1272);
and ( n26023 , n26021 , n26022 );
not ( n26024 , n26021 );
not ( n26025 , RI1745f2f8_1272);
and ( n26026 , n26024 , n26025 );
nor ( n26027 , n26023 , n26026 );
buf ( n26028 , n25655 );
buf ( n26029 , RI19aa1d20_2554);
nand ( n26030 , n26028 , n26029 );
not ( n26031 , RI17483b08_1094);
and ( n26032 , n26030 , n26031 );
not ( n26033 , n26030 );
buf ( n26034 , RI17483b08_1094);
and ( n26035 , n26033 , n26034 );
nor ( n26036 , n26032 , n26035 );
xor ( n26037 , n26027 , n26036 );
buf ( n26038 , RI19a82d30_2774);
nand ( n26039 , n25851 , n26038 );
not ( n26040 , RI17508ac8_739);
and ( n26041 , n26039 , n26040 );
not ( n26042 , n26039 );
buf ( n26043 , RI17508ac8_739);
and ( n26044 , n26042 , n26043 );
nor ( n26045 , n26041 , n26044 );
xnor ( n26046 , n26037 , n26045 );
buf ( n26047 , n26046 );
not ( n26048 , n26047 );
or ( n26049 , n26012 , n26048 );
not ( n26050 , n26046 );
not ( n26051 , n26050 );
or ( n26052 , n26051 , n26011 );
nand ( n26053 , n26049 , n26052 );
not ( n26054 , n26053 );
or ( n26055 , n26010 , n26054 );
or ( n26056 , n26053 , n26009 );
nand ( n26057 , n26055 , n26056 );
buf ( n26058 , n25362 );
buf ( n26059 , n26058 );
buf ( n26060 , RI19a876c8_2742);
nand ( n26061 , n26059 , n26060 );
not ( n26062 , RI174d1208_760);
and ( n26063 , n26061 , n26062 );
not ( n26064 , n26061 );
buf ( n26065 , RI174d1208_760);
and ( n26066 , n26064 , n26065 );
nor ( n26067 , n26063 , n26066 );
not ( n26068 , n26067 );
buf ( n26069 , RI173d46f8_1720);
not ( n26070 , n26069 );
not ( n26071 , RI1738ba08_2075);
not ( n26072 , n26071 );
or ( n26073 , n26070 , n26072 );
not ( n26074 , RI173d46f8_1720);
buf ( n26075 , RI1738ba08_2075);
nand ( n26076 , n26074 , n26075 );
nand ( n26077 , n26073 , n26076 );
not ( n26078 , RI1744c1d0_1365);
and ( n26079 , n26077 , n26078 );
not ( n26080 , n26077 );
buf ( n26081 , RI1744c1d0_1365);
and ( n26082 , n26080 , n26081 );
nor ( n26083 , n26079 , n26082 );
buf ( n26084 , RI19a9ca28_2593);
nand ( n26085 , n25540 , n26084 );
buf ( n26086 , RI174709e0_1187);
and ( n26087 , n26085 , n26086 );
not ( n26088 , n26085 );
not ( n26089 , RI174709e0_1187);
and ( n26090 , n26088 , n26089 );
nor ( n26091 , n26087 , n26090 );
xor ( n26092 , n26083 , n26091 );
buf ( n26093 , RI19acbc60_2241);
nand ( n26094 , n25851 , n26093 );
buf ( n26095 , RI174b9eb0_832);
and ( n26096 , n26094 , n26095 );
not ( n26097 , n26094 );
not ( n26098 , RI174b9eb0_832);
and ( n26099 , n26097 , n26098 );
nor ( n26100 , n26096 , n26099 );
not ( n26101 , n26100 );
xnor ( n26102 , n26092 , n26101 );
not ( n26103 , n26102 );
or ( n26104 , n26068 , n26103 );
not ( n26105 , n26067 );
not ( n26106 , n26083 );
xor ( n26107 , n26106 , n26100 );
xnor ( n26108 , n26107 , n26091 );
not ( n26109 , n26108 );
nand ( n26110 , n26105 , n26109 );
nand ( n26111 , n26104 , n26110 );
buf ( n26112 , RI173a8f40_1932);
not ( n26113 , n26112 );
not ( n26114 , RI173f1c30_1577);
not ( n26115 , n26114 );
or ( n26116 , n26113 , n26115 );
not ( n26117 , RI173a8f40_1932);
buf ( n26118 , RI173f1c30_1577);
nand ( n26119 , n26117 , n26118 );
nand ( n26120 , n26116 , n26119 );
not ( n26121 , RI174b75e8_842);
and ( n26122 , n26120 , n26121 );
not ( n26123 , n26120 );
buf ( n26124 , RI174b75e8_842);
and ( n26125 , n26123 , n26124 );
nor ( n26126 , n26122 , n26125 );
buf ( n26127 , RI19ab0870_2450);
nand ( n26128 , n25405 , n26127 );
buf ( n26129 , RI1748df18_1044);
and ( n26130 , n26128 , n26129 );
not ( n26131 , n26128 );
not ( n26132 , RI1748df18_1044);
and ( n26133 , n26131 , n26132 );
nor ( n26134 , n26130 , n26133 );
xor ( n26135 , n26126 , n26134 );
buf ( n26136 , RI19ac1d78_2315);
nand ( n26137 , n25405 , n26136 );
buf ( n26138 , RI175191c0_688);
and ( n26139 , n26137 , n26138 );
not ( n26140 , n26137 );
not ( n26141 , RI175191c0_688);
and ( n26142 , n26140 , n26141 );
nor ( n26143 , n26139 , n26142 );
not ( n26144 , n26143 );
xnor ( n26145 , n26135 , n26144 );
buf ( n26146 , n26145 );
and ( n26147 , n26111 , n26146 );
not ( n26148 , n26111 );
not ( n26149 , n26146 );
and ( n26150 , n26148 , n26149 );
nor ( n26151 , n26147 , n26150 );
nand ( n26152 , n26057 , n26151 );
not ( n26153 , n26152 );
or ( n26154 , n25982 , n26153 );
or ( n26155 , n26152 , n25981 );
nand ( n26156 , n26154 , n26155 );
not ( n26157 , n26156 );
not ( n26158 , n26157 );
or ( n26159 , n25878 , n26158 );
nand ( n26160 , n25876 , n26156 );
nand ( n26161 , n26159 , n26160 );
buf ( n26162 , n25479 );
buf ( n26163 , RI19abe6a0_2346);
nand ( n26164 , n26162 , n26163 );
not ( n26165 , RI174b1d50_869);
and ( n26166 , n26164 , n26165 );
not ( n26167 , n26164 );
buf ( n26168 , RI174b1d50_869);
and ( n26169 , n26167 , n26168 );
nor ( n26170 , n26166 , n26169 );
buf ( n26171 , RI173db9d0_1685);
not ( n26172 , n26171 );
not ( n26173 , RI17392ce0_2040);
not ( n26174 , n26173 );
or ( n26175 , n26172 , n26174 );
not ( n26176 , RI173db9d0_1685);
buf ( n26177 , RI17392ce0_2040);
nand ( n26178 , n26176 , n26177 );
nand ( n26179 , n26175 , n26178 );
not ( n26180 , RI174534a8_1330);
and ( n26181 , n26179 , n26180 );
not ( n26182 , n26179 );
buf ( n26183 , RI174534a8_1330);
and ( n26184 , n26182 , n26183 );
nor ( n26185 , n26181 , n26184 );
buf ( n26186 , RI19ac7700_2274);
nand ( n26187 , n25405 , n26186 );
buf ( n26188 , RI174c5850_796);
and ( n26189 , n26187 , n26188 );
not ( n26190 , n26187 );
not ( n26191 , RI174c5850_796);
and ( n26192 , n26190 , n26191 );
nor ( n26193 , n26189 , n26192 );
xor ( n26194 , n26185 , n26193 );
buf ( n26195 , RI19a97820_2629);
nand ( n26196 , n25915 , n26195 );
buf ( n26197 , RI17478000_1151);
and ( n26198 , n26196 , n26197 );
not ( n26199 , n26196 );
not ( n26200 , RI17478000_1151);
and ( n26201 , n26199 , n26200 );
nor ( n26202 , n26198 , n26201 );
buf ( n26203 , n26202 );
xnor ( n26204 , n26194 , n26203 );
buf ( n26205 , n26204 );
xor ( n26206 , n26170 , n26205 );
not ( n26207 , RI174146b8_1408);
not ( n26208 , RI17407170_1473);
buf ( n26209 , RI173be480_1828);
nand ( n26210 , n26208 , n26209 );
not ( n26211 , RI173be480_1828);
buf ( n26212 , RI17407170_1473);
nand ( n26213 , n26211 , n26212 );
and ( n26214 , n26210 , n26213 );
xor ( n26215 , n26207 , n26214 );
buf ( n26216 , RI17334f00_2183);
buf ( n26217 , RI174a3458_940);
xor ( n26218 , n26216 , n26217 );
buf ( n26219 , RI19ab4dd0_2417);
nand ( n26220 , n25622 , n26219 );
xnor ( n26221 , n26218 , n26220 );
xnor ( n26222 , n26215 , n26221 );
xnor ( n26223 , n26206 , n26222 );
not ( n26224 , n26223 );
buf ( n26225 , RI1738ca70_2070);
not ( n26226 , n26225 );
buf ( n26227 , RI173c6b08_1787);
not ( n26228 , n26227 );
not ( n26229 , RI1733d588_2142);
not ( n26230 , n26229 );
or ( n26231 , n26228 , n26230 );
not ( n26232 , RI173c6b08_1787);
buf ( n26233 , RI1733d588_2142);
nand ( n26234 , n26232 , n26233 );
nand ( n26235 , n26231 , n26234 );
buf ( n26236 , RI1740f7f8_1432);
and ( n26237 , n26235 , n26236 );
not ( n26238 , n26235 );
not ( n26239 , RI1740f7f8_1432);
and ( n26240 , n26238 , n26239 );
nor ( n26241 , n26237 , n26240 );
buf ( n26242 , n25450 );
buf ( n26243 , RI19a90cc8_2677);
nand ( n26244 , n26242 , n26243 );
not ( n26245 , RI17463150_1253);
and ( n26246 , n26244 , n26245 );
not ( n26247 , n26244 );
buf ( n26248 , RI17463150_1253);
and ( n26249 , n26247 , n26248 );
nor ( n26250 , n26246 , n26249 );
xor ( n26251 , n26241 , n26250 );
buf ( n26252 , RI19ac1148_2322);
nand ( n26253 , n25803 , n26252 );
not ( n26254 , RI174abe28_898);
and ( n26255 , n26253 , n26254 );
not ( n26256 , n26253 );
buf ( n26257 , RI174abe28_898);
and ( n26258 , n26256 , n26257 );
nor ( n26259 , n26255 , n26258 );
xnor ( n26260 , n26251 , n26259 );
buf ( n26261 , n26260 );
not ( n26262 , n26261 );
or ( n26263 , n26226 , n26262 );
or ( n26264 , n26261 , n26225 );
nand ( n26265 , n26263 , n26264 );
buf ( n26266 , n25571 );
buf ( n26267 , RI19aa48b8_2533);
nand ( n26268 , n26266 , n26267 );
buf ( n26269 , RI17480688_1110);
and ( n26270 , n26268 , n26269 );
not ( n26271 , n26268 );
not ( n26272 , RI17480688_1110);
and ( n26273 , n26271 , n26272 );
nor ( n26274 , n26270 , n26273 );
not ( n26275 , n26274 );
buf ( n26276 , n25490 );
buf ( n26277 , RI19a85c10_2754);
nand ( n26278 , n26276 , n26277 );
not ( n26279 , RI175019d0_755);
and ( n26280 , n26278 , n26279 );
not ( n26281 , n26278 );
buf ( n26282 , RI175019d0_755);
and ( n26283 , n26281 , n26282 );
nor ( n26284 , n26280 , n26283 );
not ( n26285 , n26284 );
or ( n26286 , n26275 , n26285 );
or ( n26287 , n26274 , n26284 );
nand ( n26288 , n26286 , n26287 );
buf ( n26289 , RI173e4058_1644);
not ( n26290 , n26289 );
not ( n26291 , RI1739b368_1999);
not ( n26292 , n26291 );
or ( n26293 , n26290 , n26292 );
not ( n26294 , RI173e4058_1644);
buf ( n26295 , RI1739b368_1999);
nand ( n26296 , n26294 , n26295 );
nand ( n26297 , n26293 , n26296 );
not ( n26298 , RI1745be78_1288);
and ( n26299 , n26297 , n26298 );
not ( n26300 , n26297 );
buf ( n26301 , RI1745be78_1288);
and ( n26302 , n26300 , n26301 );
nor ( n26303 , n26299 , n26302 );
and ( n26304 , n26288 , n26303 );
not ( n26305 , n26288 );
not ( n26306 , n26303 );
and ( n26307 , n26305 , n26306 );
nor ( n26308 , n26304 , n26307 );
not ( n26309 , n26308 );
not ( n26310 , n26309 );
buf ( n26311 , n26310 );
and ( n26312 , n26265 , n26311 );
not ( n26313 , n26265 );
not ( n26314 , n26284 );
xor ( n26315 , n26303 , n26314 );
buf ( n26316 , n26274 );
xnor ( n26317 , n26315 , n26316 );
buf ( n26318 , n26317 );
buf ( n26319 , n26318 );
and ( n26320 , n26313 , n26319 );
nor ( n26321 , n26312 , n26320 );
not ( n26322 , n26321 );
nand ( n26323 , n26224 , n26322 );
not ( n26324 , n26323 );
buf ( n26325 , n26028 );
buf ( n26326 , RI19ab5f28_2409);
nand ( n26327 , n26325 , n26326 );
buf ( n26328 , n26327 );
buf ( n26329 , RI174a1388_950);
xor ( n26330 , n26328 , n26329 );
not ( n26331 , n26330 );
buf ( n26332 , RI173f6460_1555);
not ( n26333 , n26332 );
not ( n26334 , RI173ad770_1910);
not ( n26335 , n26334 );
or ( n26336 , n26333 , n26335 );
not ( n26337 , RI173f6460_1555);
buf ( n26338 , RI173ad770_1910);
nand ( n26339 , n26337 , n26338 );
nand ( n26340 , n26336 , n26339 );
not ( n26341 , RI1752f060_620);
and ( n26342 , n26340 , n26341 );
not ( n26343 , n26340 );
buf ( n26344 , RI1752f060_620);
and ( n26345 , n26343 , n26344 );
nor ( n26346 , n26342 , n26345 );
buf ( n26347 , RI19ab3c00_2425);
nand ( n26348 , n25751 , n26347 );
buf ( n26349 , RI17520330_666);
and ( n26350 , n26348 , n26349 );
not ( n26351 , n26348 );
not ( n26352 , RI17520330_666);
and ( n26353 , n26351 , n26352 );
nor ( n26354 , n26350 , n26353 );
xor ( n26355 , n26346 , n26354 );
buf ( n26356 , RI19aac6d0_2480);
nand ( n26357 , n26162 , n26356 );
buf ( n26358 , RI17492a90_1021);
and ( n26359 , n26357 , n26358 );
not ( n26360 , n26357 );
not ( n26361 , RI17492a90_1021);
and ( n26362 , n26360 , n26361 );
nor ( n26363 , n26359 , n26362 );
xnor ( n26364 , n26355 , n26363 );
not ( n26365 , n26364 );
not ( n26366 , n26365 );
not ( n26367 , n26366 );
or ( n26368 , n26331 , n26367 );
not ( n26369 , n26364 );
not ( n26370 , n26369 );
or ( n26371 , n26370 , n26330 );
nand ( n26372 , n26368 , n26371 );
not ( n26373 , n26372 );
buf ( n26374 , RI173caca8_1767);
not ( n26375 , n26374 );
not ( n26376 , RI17341728_2122);
not ( n26377 , n26376 );
or ( n26378 , n26375 , n26377 );
not ( n26379 , RI173caca8_1767);
buf ( n26380 , RI17341728_2122);
nand ( n26381 , n26379 , n26380 );
nand ( n26382 , n26378 , n26381 );
not ( n26383 , RI17413ce0_1411);
and ( n26384 , n26382 , n26383 );
not ( n26385 , n26382 );
buf ( n26386 , RI17413ce0_1411);
and ( n26387 , n26385 , n26386 );
nor ( n26388 , n26384 , n26387 );
buf ( n26389 , RI19abf4b0_2338);
nand ( n26390 , n25405 , n26389 );
buf ( n26391 , RI174affc8_878);
and ( n26392 , n26390 , n26391 );
not ( n26393 , n26390 );
not ( n26394 , RI174affc8_878);
and ( n26395 , n26393 , n26394 );
nor ( n26396 , n26392 , n26395 );
xor ( n26397 , n26388 , n26396 );
buf ( n26398 , n26058 );
buf ( n26399 , RI19a8e8b0_2693);
nand ( n26400 , n26398 , n26399 );
buf ( n26401 , RI174672f0_1233);
and ( n26402 , n26400 , n26401 );
not ( n26403 , n26400 );
not ( n26404 , RI174672f0_1233);
and ( n26405 , n26403 , n26404 );
nor ( n26406 , n26402 , n26405 );
not ( n26407 , n26406 );
xnor ( n26408 , n26397 , n26407 );
buf ( n26409 , n26408 );
not ( n26410 , n26409 );
and ( n26411 , n26373 , n26410 );
and ( n26412 , n26372 , n26409 );
nor ( n26413 , n26411 , n26412 );
not ( n26414 , n26413 );
not ( n26415 , n26414 );
and ( n26416 , n26324 , n26415 );
and ( n26417 , n26323 , n26414 );
nor ( n26418 , n26416 , n26417 );
not ( n26419 , n26418 );
and ( n26420 , n26161 , n26419 );
not ( n26421 , n26161 );
and ( n26422 , n26421 , n26418 );
nor ( n26423 , n26420 , n26422 );
not ( n26424 , n26423 );
not ( n26425 , n25432 );
not ( n26426 , n25511 );
nand ( n26427 , n26425 , n26426 );
not ( n26428 , n26427 );
buf ( n26429 , RI19aac838_2479);
nand ( n26430 , n25741 , n26429 );
buf ( n26431 , RI17492dd8_1020);
and ( n26432 , n26430 , n26431 );
not ( n26433 , n26430 );
not ( n26434 , RI17492dd8_1020);
and ( n26435 , n26433 , n26434 );
nor ( n26436 , n26432 , n26435 );
not ( n26437 , n26436 );
buf ( n26438 , RI173e81f8_1624);
not ( n26439 , n26438 );
not ( n26440 , RI1739f1c0_1980);
not ( n26441 , n26440 );
or ( n26442 , n26439 , n26441 );
not ( n26443 , RI173e81f8_1624);
buf ( n26444 , RI1739f1c0_1980);
nand ( n26445 , n26443 , n26444 );
nand ( n26446 , n26442 , n26445 );
not ( n26447 , RI1745fcd0_1269);
and ( n26448 , n26446 , n26447 );
not ( n26449 , n26446 );
buf ( n26450 , RI1745fcd0_1269);
and ( n26451 , n26449 , n26450 );
nor ( n26452 , n26448 , n26451 );
buf ( n26453 , n25362 );
buf ( n26454 , RI19aa2248_2551);
nand ( n26455 , n26453 , n26454 );
not ( n26456 , RI174844e0_1091);
and ( n26457 , n26455 , n26456 );
not ( n26458 , n26455 );
buf ( n26459 , RI174844e0_1091);
and ( n26460 , n26458 , n26459 );
nor ( n26461 , n26457 , n26460 );
xor ( n26462 , n26452 , n26461 );
buf ( n26463 , n25741 );
buf ( n26464 , RI19a83438_2771);
nand ( n26465 , n26463 , n26464 );
not ( n26466 , RI17509a40_736);
and ( n26467 , n26465 , n26466 );
not ( n26468 , n26465 );
buf ( n26469 , RI17509a40_736);
and ( n26470 , n26468 , n26469 );
nor ( n26471 , n26467 , n26470 );
xnor ( n26472 , n26462 , n26471 );
not ( n26473 , n26472 );
or ( n26474 , n26437 , n26473 );
buf ( n26475 , n26472 );
or ( n26476 , n26475 , n26436 );
nand ( n26477 , n26474 , n26476 );
not ( n26478 , n26477 );
buf ( n26479 , RI174046c8_1486);
buf ( n26480 , RI17405730_1481);
not ( n26481 , n26480 );
not ( n26482 , RI173bca40_1836);
not ( n26483 , n26482 );
or ( n26484 , n26481 , n26483 );
not ( n26485 , RI17405730_1481);
buf ( n26486 , RI173bca40_1836);
nand ( n26487 , n26485 , n26486 );
nand ( n26488 , n26484 , n26487 );
xor ( n26489 , n26479 , n26488 );
buf ( n26490 , RI173334c0_2191);
not ( n204252 , RI174a1a18_948);
xor ( n204253 , n26490 , n204252 );
buf ( n204254 , RI19ab63d8_2407);
nand ( n204255 , n25416 , n204254 );
xnor ( n204256 , n204253 , n204255 );
xnor ( n204257 , n26489 , n204256 );
buf ( n204258 , n204257 );
not ( n204259 , n204258 );
not ( n204260 , n204259 );
or ( n204261 , n26478 , n204260 );
or ( n204262 , n204259 , n26477 );
nand ( n204263 , n204261 , n204262 );
not ( n204264 , n204263 );
and ( n204265 , n26428 , n204264 );
and ( n204266 , n26427 , n204263 );
nor ( n204267 , n204265 , n204266 );
not ( n204268 , n204267 );
not ( n204269 , RI173a2cd0_1962);
not ( n204270 , n204269 );
buf ( n204271 , RI173dcd80_1679);
not ( n204272 , n204271 );
not ( n204273 , RI17394090_2034);
not ( n204274 , n204273 );
or ( n204275 , n204272 , n204274 );
not ( n204276 , RI173dcd80_1679);
buf ( n204277 , RI17394090_2034);
nand ( n204278 , n204276 , n204277 );
nand ( n204279 , n204275 , n204278 );
not ( n204280 , n204279 );
or ( n204281 , n204270 , n204280 );
or ( n204282 , n204279 , n204269 );
nand ( n204283 , n204281 , n204282 );
not ( n204284 , n204283 );
not ( n204285 , RI17454858_1324);
buf ( n204286 , RI19ac5e28_2285);
nand ( n204287 , n25529 , n204286 );
not ( n204288 , n204287 );
buf ( n204289 , RI174c7740_790);
not ( n204290 , n204289 );
and ( n204291 , n204288 , n204290 );
nand ( n204292 , n25628 , n204286 );
and ( n204293 , n204292 , n204289 );
nor ( n204294 , n204291 , n204293 );
xor ( n204295 , n204285 , n204294 );
buf ( n204296 , RI19a96038_2640);
nand ( n204297 , n25583 , n204296 );
not ( n204298 , n204297 );
buf ( n204299 , RI174793b0_1145);
not ( n204300 , n204299 );
and ( n204301 , n204298 , n204300 );
nand ( n204302 , n25376 , n204296 );
and ( n204303 , n204302 , n204299 );
nor ( n204304 , n204301 , n204303 );
xnor ( n204305 , n204295 , n204304 );
not ( n204306 , n204305 );
not ( n204307 , n204306 );
or ( n204308 , n204284 , n204307 );
or ( n204309 , n204306 , n204283 );
nand ( n204310 , n204308 , n204309 );
not ( n204311 , n204310 );
buf ( n204312 , RI173fa2b8_1536);
not ( n204313 , n204312 );
not ( n204314 , RI173b15c8_1891);
not ( n204315 , n204314 );
or ( n204316 , n204313 , n204315 );
not ( n204317 , RI173fa2b8_1536);
buf ( n204318 , RI173b15c8_1891);
nand ( n204319 , n204317 , n204318 );
nand ( n204320 , n204316 , n204319 );
buf ( n204321 , RI17394db0_2030);
and ( n204322 , n204320 , n204321 );
not ( n204323 , n204320 );
not ( n204324 , RI17394db0_2030);
and ( n204325 , n204323 , n204324 );
nor ( n204326 , n204322 , n204325 );
buf ( n204327 , RI19aa9d90_2497);
nand ( n204328 , n26266 , n204327 );
buf ( n204329 , RI174968e8_1002);
and ( n204330 , n204328 , n204329 );
not ( n204331 , n204328 );
not ( n204332 , RI174968e8_1002);
and ( n204333 , n204331 , n204332 );
nor ( n204334 , n204330 , n204333 );
xor ( n204335 , n204326 , n204334 );
buf ( n204336 , n25363 );
buf ( n204337 , RI19a9cc08_2592);
nand ( n204338 , n204336 , n204337 );
buf ( n204339 , RI17526528_647);
and ( n204340 , n204338 , n204339 );
not ( n204341 , n204338 );
not ( n204342 , RI17526528_647);
and ( n204343 , n204341 , n204342 );
nor ( n204344 , n204340 , n204343 );
not ( n204345 , n204344 );
xnor ( n204346 , n204335 , n204345 );
not ( n204347 , n204346 );
not ( n204348 , n204347 );
or ( n204349 , n204311 , n204348 );
buf ( n204350 , n204347 );
or ( n204351 , n204350 , n204310 );
nand ( n204352 , n204349 , n204351 );
not ( n204353 , n204352 );
buf ( n204354 , RI19aa0358_2567);
nand ( n204355 , n26453 , n204354 );
buf ( n204356 , RI17488338_1072);
and ( n204357 , n204355 , n204356 );
not ( n204358 , n204355 );
not ( n204359 , RI17488338_1072);
and ( n204360 , n204358 , n204359 );
nor ( n204361 , n204357 , n204360 );
not ( n204362 , n204361 );
buf ( n204363 , RI19acef78_2218);
nand ( n204364 , n26398 , n204363 );
not ( n204365 , RI1750fc38_717);
and ( n204366 , n204364 , n204365 );
not ( n204367 , n204364 );
buf ( n204368 , RI1750fc38_717);
and ( n204369 , n204367 , n204368 );
nor ( n204370 , n204366 , n204369 );
not ( n204371 , n204370 );
or ( n204372 , n204362 , n204371 );
or ( n204373 , n204361 , n204370 );
nand ( n204374 , n204372 , n204373 );
buf ( n204375 , RI173a3360_1960);
not ( n204376 , n204375 );
not ( n204377 , RI173ec050_1605);
not ( n204378 , n204377 );
or ( n204379 , n204376 , n204378 );
not ( n204380 , RI173a3360_1960);
buf ( n204381 , RI173ec050_1605);
nand ( n204382 , n204380 , n204381 );
nand ( n204383 , n204379 , n204382 );
not ( n204384 , RI1747c4e8_1130);
and ( n204385 , n204383 , n204384 );
not ( n204386 , n204383 );
buf ( n204387 , RI1747c4e8_1130);
and ( n204388 , n204386 , n204387 );
nor ( n204389 , n204385 , n204388 );
xnor ( n204390 , n204374 , n204389 );
buf ( n204391 , n204390 );
not ( n204392 , n204391 );
buf ( n204393 , n25582 );
buf ( n204394 , RI19ac6080_2284);
nand ( n204395 , n204393 , n204394 );
not ( n204396 , RI174c7c68_789);
and ( n204397 , n204395 , n204396 );
not ( n204398 , n204395 );
buf ( n204399 , RI174c7c68_789);
and ( n204400 , n204398 , n204399 );
nor ( n204401 , n204397 , n204400 );
buf ( n204402 , RI173ceb00_1748);
not ( n204403 , n204402 );
not ( n204404 , RI17345238_2104);
not ( n204405 , n204404 );
or ( n204406 , n204403 , n204405 );
not ( n204407 , RI173ceb00_1748);
buf ( n204408 , RI17345238_2104);
nand ( n204409 , n204407 , n204408 );
nand ( n204410 , n204406 , n204409 );
buf ( n204411 , RI174465f0_1393);
and ( n204412 , n204410 , n204411 );
not ( n204413 , n204410 );
not ( n204414 , RI174465f0_1393);
and ( n204415 , n204413 , n204414 );
nor ( n204416 , n204412 , n204415 );
buf ( n204417 , RI19abd6b0_2355);
nand ( n204418 , n25915 , n204417 );
buf ( n204419 , RI174b3ad8_860);
and ( n204420 , n204418 , n204419 );
not ( n204421 , n204418 );
not ( n204422 , RI174b3ad8_860);
and ( n204423 , n204421 , n204422 );
nor ( n204424 , n204420 , n204423 );
xor ( n204425 , n204416 , n204424 );
buf ( n204426 , n26276 );
buf ( n204427 , RI19a8c240_2710);
nand ( n204428 , n204426 , n204427 );
not ( n204429 , RI1746ae00_1215);
and ( n204430 , n204428 , n204429 );
not ( n204431 , n204428 );
buf ( n204432 , RI1746ae00_1215);
and ( n204433 , n204431 , n204432 );
nor ( n204434 , n204430 , n204433 );
xnor ( n204435 , n204425 , n204434 );
not ( n204436 , n204435 );
and ( n204437 , n204401 , n204436 );
not ( n204438 , n204401 );
buf ( n204439 , n204435 );
and ( n204440 , n204438 , n204439 );
nor ( n204441 , n204437 , n204440 );
not ( n204442 , n204441 );
or ( n204443 , n204392 , n204442 );
or ( n204444 , n204441 , n204391 );
nand ( n204445 , n204443 , n204444 );
not ( n204446 , n204445 );
not ( n204447 , n204446 );
nor ( n204448 , n204353 , n204447 );
not ( n204449 , n204448 );
buf ( n204450 , RI19a8a2d8_2723);
nand ( n204451 , n25529 , n204450 );
buf ( n204452 , RI1746f630_1193);
xor ( n204453 , n204451 , n204452 );
buf ( n204454 , n204453 );
not ( n204455 , n204454 );
buf ( n204456 , RI175361d0_598);
buf ( n204457 , RI1740d3e0_1443);
not ( n204458 , n204457 );
not ( n204459 , RI173c46f0_1798);
not ( n204460 , n204459 );
or ( n204461 , n204458 , n204460 );
not ( n204462 , RI1740d3e0_1443);
buf ( n204463 , RI173c46f0_1798);
nand ( n204464 , n204462 , n204463 );
nand ( n204465 , n204461 , n204464 );
xor ( n204466 , n204456 , n204465 );
buf ( n204467 , RI1733b170_2153);
buf ( n204468 , RI174a9a10_909);
xor ( n204469 , n204467 , n204468 );
buf ( n204470 , RI19ab1ef0_2440);
nand ( n204471 , n25793 , n204470 );
xnor ( n204472 , n204469 , n204471 );
xor ( n204473 , n204466 , n204472 );
not ( n204474 , n204473 );
or ( n204475 , n204455 , n204474 );
or ( n204476 , n204473 , n204454 );
nand ( n204477 , n204475 , n204476 );
buf ( n204478 , RI173d3690_1725);
not ( n204479 , n204478 );
not ( n204480 , RI1738a9a0_2080);
not ( n204481 , n204480 );
or ( n204482 , n204479 , n204481 );
not ( n204483 , RI173d3690_1725);
buf ( n204484 , RI1738a9a0_2080);
nand ( n204485 , n204483 , n204484 );
nand ( n204486 , n204482 , n204485 );
not ( n204487 , RI1744b168_1370);
and ( n204488 , n204486 , n204487 );
not ( n204489 , n204486 );
buf ( n204490 , RI1744b168_1370);
and ( n204491 , n204489 , n204490 );
nor ( n204492 , n204488 , n204491 );
buf ( n204493 , n25655 );
buf ( n204494 , RI19acb300_2246);
nand ( n204495 , n204493 , n204494 );
buf ( n204496 , RI174b8650_837);
and ( n204497 , n204495 , n204496 );
not ( n204498 , n204495 );
not ( n204499 , RI174b8650_837);
and ( n204500 , n204498 , n204499 );
nor ( n204501 , n204497 , n204500 );
xor ( n204502 , n204492 , n204501 );
xnor ( n204503 , n204502 , n25888 );
buf ( n204504 , n204503 );
buf ( n204505 , n204504 );
and ( n204506 , n204477 , n204505 );
not ( n204507 , n204477 );
not ( n204508 , n204504 );
and ( n204509 , n204507 , n204508 );
nor ( n204510 , n204506 , n204509 );
not ( n204511 , n204510 );
buf ( n204512 , n25655 );
buf ( n204513 , n204512 );
buf ( n204514 , n204513 );
not ( n204515 , n204514 );
not ( n204516 , RI175385e8_592);
not ( n204517 , RI17539218_590);
not ( n204518 , RI17539e48_588);
and ( n204519 , n204516 , n204517 , n204518 );
buf ( n204520 , RI17537fd0_593);
buf ( n204521 , RI17536770_597);
nor ( n204522 , n204520 , n204521 );
not ( n204523 , RI175379b8_594);
and ( n204524 , n204522 , n204523 );
not ( n204525 , RI17539830_589);
nand ( n204526 , n204515 , n204519 , n204524 , n204525 );
not ( n204527 , n204526 );
and ( n204528 , n204511 , n204527 );
not ( n204529 , n204511 );
and ( n204530 , n204529 , n204526 );
nor ( n204531 , n204528 , n204530 );
not ( n204532 , n204531 );
or ( n204533 , n204449 , n204532 );
or ( n204534 , n204531 , n204448 );
nand ( n204535 , n204533 , n204534 );
not ( n204536 , n204535 );
and ( n204537 , n204268 , n204536 );
and ( n204538 , n204267 , n204535 );
nor ( n204539 , n204537 , n204538 );
not ( n204540 , n204539 );
and ( n204541 , n26424 , n204540 );
not ( n204542 , n26424 );
and ( n204543 , n204542 , n204539 );
nor ( n204544 , n204541 , n204543 );
not ( n204545 , n204544 );
or ( n204546 , n25607 , n204545 );
not ( n204547 , n25606 );
not ( n204548 , n204539 );
not ( n204549 , n26423 );
or ( n204550 , n204548 , n204549 );
not ( n204551 , n26423 );
nand ( n204552 , n204551 , n204540 );
nand ( n204553 , n204550 , n204552 );
nand ( n204554 , n204547 , n204553 );
nand ( n204555 , n204546 , n204554 );
buf ( n204556 , RI174118c8_1422);
not ( n204557 , n204556 );
not ( n204558 , RI173eda90_1597);
buf ( n204559 , RI17403318_1492);
not ( n204560 , n204559 );
not ( n204561 , RI173ba628_1847);
not ( n204562 , n204561 );
or ( n204563 , n204560 , n204562 );
not ( n204564 , RI17403318_1492);
buf ( n204565 , RI173ba628_1847);
nand ( n204566 , n204564 , n204565 );
nand ( n204567 , n204563 , n204566 );
not ( n204568 , n204567 );
xor ( n204569 , n204558 , n204568 );
buf ( n204570 , RI175342e0_604);
not ( n204571 , n204570 );
buf ( n204572 , n25490 );
buf ( n204573 , RI19ab73c8_2400);
nand ( n204574 , n204572 , n204573 );
buf ( n204575 , RI1749f600_959);
and ( n204576 , n204574 , n204575 );
not ( n204577 , n204574 );
not ( n204578 , RI1749f600_959);
and ( n204579 , n204577 , n204578 );
nor ( n204580 , n204576 , n204579 );
not ( n204581 , n204580 );
or ( n204582 , n204571 , n204581 );
or ( n204583 , n204580 , n204570 );
nand ( n204584 , n204582 , n204583 );
xnor ( n204585 , n204569 , n204584 );
buf ( n204586 , n204585 );
not ( n204587 , n204586 );
or ( n204588 , n204557 , n204587 );
or ( n204589 , n204586 , n204556 );
nand ( n204590 , n204588 , n204589 );
buf ( n204591 , RI1744f650_1349);
buf ( n204592 , RI19a99f80_2612);
nand ( n204593 , n25479 , n204592 );
buf ( n204594 , RI17473e60_1171);
and ( n204595 , n204593 , n204594 );
not ( n204596 , n204593 );
not ( n204597 , RI17473e60_1171);
and ( n204598 , n204596 , n204597 );
nor ( n204599 , n204595 , n204598 );
xor ( n204600 , n204591 , n204599 );
buf ( n204601 , RI19ac96e0_2259);
nand ( n204602 , n25666 , n204601 );
not ( n204603 , RI174bf658_815);
and ( n204604 , n204602 , n204603 );
not ( n204605 , n204602 );
buf ( n204606 , RI174bf658_815);
and ( n204607 , n204605 , n204606 );
nor ( n204608 , n204604 , n204607 );
xnor ( n204609 , n204600 , n204608 );
not ( n204610 , n204609 );
not ( n204611 , RI173d7b78_1704);
buf ( n204612 , RI1738ee88_2059);
and ( n204613 , n204611 , n204612 );
not ( n204614 , n204611 );
not ( n204615 , RI1738ee88_2059);
and ( n204616 , n204614 , n204615 );
nor ( n204617 , n204613 , n204616 );
not ( n204618 , n204617 );
and ( n204619 , n204610 , n204618 );
and ( n204620 , n204609 , n204617 );
nor ( n204621 , n204619 , n204620 );
buf ( n204622 , n204621 );
and ( n204623 , n204590 , n204622 );
not ( n204624 , n204590 );
not ( n204625 , n204617 );
not ( n204626 , n204625 );
not ( n204627 , n204609 );
not ( n204628 , n204627 );
or ( n204629 , n204626 , n204628 );
nand ( n204630 , n204609 , n204617 );
nand ( n204631 , n204629 , n204630 );
buf ( n204632 , n204631 );
and ( n204633 , n204624 , n204632 );
nor ( n204634 , n204623 , n204633 );
not ( n204635 , n204634 );
buf ( n204636 , RI17400f00_1503);
not ( n204637 , n204636 );
buf ( n204638 , RI173f2608_1574);
not ( n204639 , n204638 );
not ( n204640 , RI173a9918_1929);
not ( n204641 , n204640 );
or ( n204642 , n204639 , n204641 );
not ( n204643 , RI173f2608_1574);
buf ( n204644 , RI173a9918_1929);
nand ( n204645 , n204643 , n204644 );
nand ( n204646 , n204642 , n204645 );
not ( n204647 , RI174be1b8_819);
and ( n204648 , n204646 , n204647 );
not ( n204649 , n204646 );
buf ( n204650 , RI174be1b8_819);
and ( n204651 , n204649 , n204650 );
nor ( n204652 , n204648 , n204651 );
buf ( n204653 , RI19aae7a0_2465);
nand ( n204654 , n25803 , n204653 );
buf ( n204655 , RI1748ec38_1040);
and ( n204656 , n204654 , n204655 );
not ( n204657 , n204654 );
not ( n204658 , RI1748ec38_1040);
and ( n204659 , n204657 , n204658 );
nor ( n204660 , n204656 , n204659 );
xor ( n204661 , n204652 , n204660 );
buf ( n204662 , RI19a23330_2795);
nand ( n204663 , n204426 , n204662 );
not ( n204664 , RI1751a138_685);
and ( n204665 , n204663 , n204664 );
not ( n204666 , n204663 );
buf ( n204667 , RI1751a138_685);
and ( n204668 , n204666 , n204667 );
nor ( n204669 , n204665 , n204668 );
xnor ( n204670 , n204661 , n204669 );
buf ( n204671 , n204670 );
buf ( n204672 , n204671 );
not ( n204673 , n204672 );
or ( n204674 , n204637 , n204673 );
not ( n204675 , n204670 );
not ( n204676 , n204675 );
not ( n204677 , n204676 );
not ( n204678 , RI17400f00_1503);
nand ( n204679 , n204677 , n204678 );
nand ( n204680 , n204674 , n204679 );
not ( n204681 , n26261 );
and ( n204682 , n204680 , n204681 );
not ( n204683 , n204680 );
and ( n204684 , n204683 , n26261 );
nor ( n204685 , n204682 , n204684 );
not ( n204686 , n204685 );
nand ( n204687 , n204635 , n204686 );
not ( n204688 , n204687 );
buf ( n204689 , RI173ad428_1911);
not ( n204690 , n204689 );
buf ( n204691 , RI173e7b68_1626);
not ( n204692 , n204691 );
not ( n204693 , RI1739eb30_1982);
not ( n204694 , n204693 );
or ( n204695 , n204692 , n204694 );
not ( n204696 , RI173e7b68_1626);
buf ( n204697 , RI1739eb30_1982);
nand ( n204698 , n204696 , n204697 );
nand ( n204699 , n204695 , n204698 );
not ( n204700 , RI1745f640_1271);
and ( n204701 , n204699 , n204700 );
not ( n204702 , n204699 );
buf ( n204703 , RI1745f640_1271);
and ( n204704 , n204702 , n204703 );
nor ( n204705 , n204701 , n204704 );
buf ( n204706 , RI19a82f88_2773);
nand ( n204707 , n26242 , n204706 );
buf ( n204708 , RI17508ff0_738);
and ( n204709 , n204707 , n204708 );
not ( n204710 , n204707 );
not ( n204711 , RI17508ff0_738);
and ( n204712 , n204710 , n204711 );
nor ( n204713 , n204709 , n204712 );
xor ( n204714 , n204705 , n204713 );
buf ( n204715 , RI19aa1f00_2553);
nand ( n204716 , n25622 , n204715 );
buf ( n204717 , RI17483e50_1093);
and ( n204718 , n204716 , n204717 );
not ( n204719 , n204716 );
not ( n204720 , RI17483e50_1093);
and ( n204721 , n204719 , n204720 );
nor ( n204722 , n204718 , n204721 );
xor ( n204723 , n204714 , n204722 );
not ( n204724 , n204723 );
or ( n204725 , n204690 , n204724 );
not ( n204726 , n204723 );
not ( n204727 , n204726 );
not ( n204728 , n204727 );
not ( n204729 , RI173ad428_1911);
nand ( n204730 , n204728 , n204729 );
nand ( n204731 , n204725 , n204730 );
buf ( n204732 , RI173ffe98_1508);
not ( n204733 , RI174050a0_1483);
buf ( n204734 , RI173bc3b0_1838);
nand ( n204735 , n204733 , n204734 );
not ( n204736 , RI173bc3b0_1838);
buf ( n204737 , RI174050a0_1483);
nand ( n204738 , n204736 , n204737 );
and ( n204739 , n204735 , n204738 );
xor ( n204740 , n204732 , n204739 );
buf ( n204741 , RI17332e30_2193);
xor ( n204742 , n204741 , n26329 );
xnor ( n204743 , n204742 , n26327 );
xnor ( n204744 , n204740 , n204743 );
not ( n204745 , n204744 );
not ( n204746 , n204745 );
and ( n204747 , n204731 , n204746 );
not ( n204748 , n204731 );
and ( n204749 , n204748 , n204745 );
nor ( n204750 , n204747 , n204749 );
not ( n204751 , n204750 );
and ( n204752 , n204688 , n204751 );
and ( n204753 , n204687 , n204750 );
nor ( n204754 , n204752 , n204753 );
not ( n204755 , n204754 );
not ( n204756 , n204755 );
buf ( n204757 , RI173e5750_1637);
buf ( n204758 , RI173f4048_1566);
not ( n204759 , n204758 );
not ( n204760 , RI173ab358_1921);
not ( n204761 , n204760 );
or ( n204762 , n204759 , n204761 );
not ( n204763 , RI173f4048_1566);
buf ( n204764 , RI173ab358_1921);
nand ( n204765 , n204763 , n204764 );
nand ( n204766 , n204762 , n204765 );
not ( n204767 , RI1750b408_731);
and ( n204768 , n204766 , n204767 );
not ( n204769 , n204766 );
buf ( n204770 , RI1750b408_731);
and ( n204771 , n204769 , n204770 );
nor ( n204772 , n204768 , n204771 );
buf ( n204773 , RI19abcfa8_2359);
nand ( n204774 , n25479 , n204773 );
buf ( n204775 , RI1751ca78_677);
and ( n204776 , n204774 , n204775 );
not ( n204777 , n204774 );
not ( n204778 , RI1751ca78_677);
and ( n204779 , n204777 , n204778 );
nor ( n204780 , n204776 , n204779 );
xor ( n204781 , n204772 , n204780 );
buf ( n204782 , RI19aad300_2474);
nand ( n204783 , n26059 , n204782 );
not ( n204784 , RI17490678_1032);
and ( n204785 , n204783 , n204784 );
not ( n204786 , n204783 );
buf ( n204787 , RI17490678_1032);
and ( n204788 , n204786 , n204787 );
nor ( n204789 , n204785 , n204788 );
xnor ( n204790 , n204781 , n204789 );
not ( n204791 , n204790 );
not ( n204792 , n204791 );
xor ( n204793 , n204757 , n204792 );
buf ( n204794 , RI1744e5e8_1354);
buf ( n204795 , RI19acb120_2247);
nand ( n204796 , n25628 , n204795 );
buf ( n204797 , RI174bd768_821);
and ( n204798 , n204796 , n204797 );
not ( n204799 , n204796 );
not ( n204800 , RI174bd768_821);
and ( n204801 , n204799 , n204800 );
nor ( n204802 , n204798 , n204801 );
xor ( n204803 , n204794 , n204802 );
buf ( n204804 , RI19a9bd80_2599);
nand ( n204805 , n26059 , n204804 );
not ( n204806 , RI17472df8_1176);
and ( n204807 , n204805 , n204806 );
not ( n204808 , n204805 );
buf ( n204809 , RI17472df8_1176);
and ( n204810 , n204808 , n204809 );
nor ( n204811 , n204807 , n204810 );
xnor ( n204812 , n204803 , n204811 );
not ( n204813 , n204812 );
not ( n204814 , RI173d6b10_1709);
buf ( n204815 , RI1738de20_2064);
and ( n204816 , n204814 , n204815 );
not ( n204817 , n204814 );
not ( n204818 , RI1738de20_2064);
and ( n204819 , n204817 , n204818 );
nor ( n204820 , n204816 , n204819 );
not ( n204821 , n204820 );
and ( n204822 , n204813 , n204821 );
and ( n204823 , n204812 , n204820 );
nor ( n204824 , n204822 , n204823 );
buf ( n204825 , n204824 );
xor ( n204826 , n204793 , n204825 );
not ( n204827 , n204826 );
buf ( n204828 , RI17497950_997);
not ( n204829 , RI173eeaf8_1592);
buf ( n204830 , RI173a5e08_1947);
nand ( n204831 , n204829 , n204830 );
not ( n204832 , RI173a5e08_1947);
buf ( n204833 , RI173eeaf8_1592);
nand ( n204834 , n204832 , n204833 );
and ( n204835 , n204831 , n204834 );
xor ( n204836 , n204828 , n204835 );
buf ( n204837 , RI19acc200_2238);
nand ( n204838 , n25539 , n204837 );
buf ( n204839 , RI17514468_703);
and ( n204840 , n204838 , n204839 );
not ( n204841 , n204838 );
not ( n204842 , RI17514468_703);
and ( n204843 , n204841 , n204842 );
nor ( n204844 , n204840 , n204843 );
not ( n204845 , n204844 );
buf ( n204846 , RI19a9d400_2589);
nand ( n204847 , n25529 , n204846 );
not ( n204848 , RI1748ade0_1059);
and ( n204849 , n204847 , n204848 );
not ( n204850 , n204847 );
buf ( n204851 , RI1748ade0_1059);
and ( n204852 , n204850 , n204851 );
nor ( n204853 , n204849 , n204852 );
not ( n204854 , n204853 );
or ( n204855 , n204845 , n204854 );
or ( n204856 , n204844 , n204853 );
nand ( n204857 , n204855 , n204856 );
xnor ( n204858 , n204836 , n204857 );
buf ( n204859 , n204858 );
not ( n204860 , n204859 );
not ( n204861 , n204860 );
buf ( n204862 , RI173b2630_1886);
not ( n204863 , n204862 );
and ( n204864 , n204861 , n204863 );
and ( n204865 , n204860 , n204862 );
nor ( n204866 , n204864 , n204865 );
buf ( n204867 , RI173b6e60_1864);
not ( n204868 , RI1740c030_1449);
buf ( n204869 , RI173c3340_1804);
and ( n204870 , n204868 , n204869 );
not ( n204871 , n204868 );
not ( n204872 , RI173c3340_1804);
and ( n204873 , n204871 , n204872 );
nor ( n204874 , n204870 , n204873 );
xor ( n204875 , n204867 , n204874 );
buf ( n204876 , RI17339dc0_2159);
not ( n204877 , n204876 );
buf ( n204878 , RI19ab0ff0_2446);
nand ( n204879 , n25491 , n204878 );
buf ( n204880 , RI174a8660_915);
and ( n204881 , n204879 , n204880 );
not ( n204882 , n204879 );
not ( n204883 , RI174a8660_915);
and ( n204884 , n204882 , n204883 );
nor ( n204885 , n204881 , n204884 );
not ( n204886 , n204885 );
or ( n204887 , n204877 , n204886 );
or ( n204888 , n204885 , n204876 );
nand ( n204889 , n204887 , n204888 );
xnor ( n204890 , n204875 , n204889 );
not ( n204891 , n204890 );
buf ( n204892 , n204891 );
and ( n204893 , n204866 , n204892 );
not ( n204894 , n204866 );
not ( n204895 , n204892 );
and ( n204896 , n204894 , n204895 );
nor ( n204897 , n204893 , n204896 );
nand ( n204898 , n204827 , n204897 );
buf ( n204899 , RI1738cdb8_2069);
not ( n204900 , n204899 );
buf ( n204901 , RI173c7198_1785);
not ( n204902 , n204901 );
not ( n204903 , RI1733dc18_2140);
not ( n204904 , n204903 );
or ( n204905 , n204902 , n204904 );
not ( n204906 , RI173c7198_1785);
buf ( n204907 , RI1733dc18_2140);
nand ( n204908 , n204906 , n204907 );
nand ( n204909 , n204905 , n204908 );
buf ( n204910 , RI1740fe88_1430);
and ( n204911 , n204909 , n204910 );
not ( n204912 , n204909 );
not ( n204913 , RI1740fe88_1430);
and ( n204914 , n204912 , n204913 );
nor ( n204915 , n204911 , n204914 );
buf ( n204916 , n26058 );
buf ( n204917 , RI19a90f20_2676);
nand ( n204918 , n204916 , n204917 );
not ( n204919 , RI174637e0_1251);
and ( n204920 , n204918 , n204919 );
not ( n204921 , n204918 );
buf ( n204922 , RI174637e0_1251);
and ( n204923 , n204921 , n204922 );
nor ( n204924 , n204920 , n204923 );
xor ( n204925 , n204915 , n204924 );
buf ( n204926 , n25656 );
buf ( n204927 , RI19ac12b0_2321);
nand ( n204928 , n204926 , n204927 );
not ( n204929 , RI174ac4b8_896);
and ( n204930 , n204928 , n204929 );
not ( n204931 , n204928 );
buf ( n204932 , RI174ac4b8_896);
and ( n204933 , n204931 , n204932 );
nor ( n204934 , n204930 , n204933 );
xnor ( n204935 , n204925 , n204934 );
buf ( n204936 , n204935 );
not ( n204937 , n204936 );
or ( n204938 , n204900 , n204937 );
not ( n204939 , n204936 );
not ( n204940 , RI1738cdb8_2069);
nand ( n204941 , n204939 , n204940 );
nand ( n204942 , n204938 , n204941 );
buf ( n204943 , RI173e43a0_1643);
not ( n204944 , n204943 );
not ( n204945 , RI1739b6b0_1998);
not ( n204946 , n204945 );
or ( n204947 , n204944 , n204946 );
not ( n204948 , RI173e43a0_1643);
buf ( n204949 , RI1739b6b0_1998);
nand ( n204950 , n204948 , n204949 );
nand ( n204951 , n204947 , n204950 );
buf ( n204952 , RI1745c1c0_1287);
and ( n204953 , n204951 , n204952 );
not ( n204954 , n204951 );
not ( n204955 , RI1745c1c0_1287);
and ( n204956 , n204954 , n204955 );
nor ( n204957 , n204953 , n204956 );
buf ( n204958 , RI19a85e68_2753);
nand ( n204959 , n25572 , n204958 );
buf ( n204960 , RI17501ef8_754);
and ( n204961 , n204959 , n204960 );
not ( n204962 , n204959 );
not ( n204963 , RI17501ef8_754);
and ( n204964 , n204962 , n204963 );
nor ( n204965 , n204961 , n204964 );
xor ( n204966 , n204957 , n204965 );
buf ( n204967 , RI19aa4a98_2532);
nand ( n204968 , n204393 , n204967 );
not ( n204969 , RI174809d0_1109);
and ( n204970 , n204968 , n204969 );
not ( n204971 , n204968 );
buf ( n204972 , RI174809d0_1109);
and ( n204973 , n204971 , n204972 );
nor ( n204974 , n204970 , n204973 );
xnor ( n204975 , n204966 , n204974 );
buf ( n204976 , n204975 );
not ( n204977 , n204976 );
not ( n204978 , n204977 );
and ( n204979 , n204942 , n204978 );
not ( n204980 , n204942 );
not ( n204981 , n204976 );
and ( n204982 , n204980 , n204981 );
nor ( n204983 , n204979 , n204982 );
buf ( n204984 , n204983 );
xnor ( n204985 , n204898 , n204984 );
not ( n204986 , n204985 );
not ( n204987 , n204986 );
or ( n204988 , n204756 , n204987 );
nand ( n204989 , n204985 , n204754 );
nand ( n204990 , n204988 , n204989 );
not ( n204991 , n204990 );
not ( n204992 , n204991 );
buf ( n204993 , RI173e4a30_1641);
not ( n204994 , n204993 );
buf ( n204995 , RI173f39b8_1568);
not ( n204996 , n204995 );
not ( n204997 , RI173aacc8_1923);
not ( n204998 , n204997 );
or ( n204999 , n204996 , n204998 );
not ( n205000 , RI173f39b8_1568);
buf ( n205001 , RI173aacc8_1923);
nand ( n205002 , n205000 , n205001 );
nand ( n205003 , n204999 , n205002 );
not ( n205004 , RI17502420_753);
and ( n205005 , n205003 , n205004 );
not ( n205006 , n205003 );
buf ( n205007 , RI17502420_753);
and ( n205008 , n205006 , n205007 );
nor ( n205009 , n205005 , n205008 );
buf ( n205010 , RI19a23150_2796);
nand ( n205011 , n204493 , n205010 );
buf ( n205012 , RI1751c028_679);
and ( n205013 , n205011 , n205012 );
not ( n205014 , n205011 );
not ( n205015 , RI1751c028_679);
and ( n205016 , n205014 , n205015 );
nor ( n205017 , n205013 , n205016 );
xor ( n205018 , n205009 , n205017 );
buf ( n205019 , n25490 );
buf ( n205020 , n205019 );
buf ( n205021 , RI19aaf628_2458);
nand ( n205022 , n205020 , n205021 );
not ( n205023 , RI1748ffe8_1034);
and ( n205024 , n205022 , n205023 );
not ( n205025 , n205022 );
buf ( n205026 , RI1748ffe8_1034);
and ( n205027 , n205025 , n205026 );
nor ( n205028 , n205024 , n205027 );
xnor ( n205029 , n205018 , n205028 );
not ( n205030 , n205029 );
or ( n205031 , n204994 , n205030 );
not ( n205032 , n204993 );
not ( n205033 , n205029 );
nand ( n205034 , n205032 , n205033 );
nand ( n205035 , n205031 , n205034 );
buf ( n205036 , RI173c8200_1780);
not ( n205037 , n205036 );
not ( n205038 , RI1733ec80_2135);
not ( n205039 , n205038 );
or ( n205040 , n205037 , n205039 );
not ( n205041 , RI173c8200_1780);
buf ( n205042 , RI1733ec80_2135);
nand ( n205043 , n205041 , n205042 );
nand ( n205044 , n205040 , n205043 );
buf ( n205045 , RI17410ef0_1425);
and ( n205046 , n205044 , n205045 );
not ( n205047 , n205044 );
not ( n205048 , RI17410ef0_1425);
and ( n205049 , n205047 , n205048 );
nor ( n205050 , n205046 , n205049 );
buf ( n205051 , RI19ac1b98_2316);
nand ( n205052 , n25479 , n205051 );
buf ( n205053 , RI174ad520_891);
and ( n205054 , n205052 , n205053 );
not ( n205055 , n205052 );
not ( n205056 , RI174ad520_891);
and ( n205057 , n205055 , n205056 );
nor ( n205058 , n205054 , n205057 );
xor ( n205059 , n205050 , n205058 );
buf ( n205060 , RI19a919e8_2671);
nand ( n205061 , n25803 , n205060 );
buf ( n205062 , RI17464848_1246);
and ( n205063 , n205061 , n205062 );
not ( n205064 , n205061 );
not ( n205065 , RI17464848_1246);
and ( n205066 , n205064 , n205065 );
nor ( n205067 , n205063 , n205066 );
xnor ( n205068 , n205059 , n205067 );
and ( n205069 , n205035 , n205068 );
not ( n205070 , n205035 );
xor ( n205071 , n205050 , n205067 );
xor ( n205072 , n205071 , n205058 );
not ( n205073 , n205072 );
not ( n205074 , n205073 );
and ( n205075 , n205070 , n205074 );
nor ( n205076 , n205069 , n205075 );
not ( n205077 , n205076 );
buf ( n205078 , RI173f6af0_1553);
buf ( n205079 , RI17404038_1488);
not ( n205080 , n205079 );
not ( n205081 , RI173bb348_1843);
not ( n205082 , n205081 );
or ( n205083 , n205080 , n205082 );
not ( n205084 , RI17404038_1488);
buf ( n205085 , RI173bb348_1843);
nand ( n205086 , n205084 , n205085 );
nand ( n205087 , n205083 , n205086 );
xor ( n205088 , n205078 , n205087 );
buf ( n205089 , RI17535780_600);
not ( n205090 , RI174a0320_955);
xor ( n205091 , n205089 , n205090 );
buf ( n205092 , RI19ab7da0_2396);
nand ( n205093 , n25666 , n205092 );
xnor ( n205094 , n205091 , n205093 );
xnor ( n205095 , n205088 , n205094 );
not ( n205096 , n205095 );
not ( n205097 , n205096 );
buf ( n205098 , RI173f53f8_1560);
not ( n205099 , n205098 );
buf ( n205100 , RI173e6b00_1631);
not ( n205101 , n205100 );
not ( n205102 , RI1739dac8_1987);
not ( n205103 , n205102 );
or ( n205104 , n205101 , n205103 );
not ( n205105 , RI173e6b00_1631);
buf ( n205106 , RI1739dac8_1987);
nand ( n205107 , n205105 , n205106 );
nand ( n205108 , n205104 , n205107 );
buf ( n205109 , RI1745e5d8_1276);
and ( n205110 , n205108 , n205109 );
not ( n205111 , n205108 );
not ( n205112 , RI1745e5d8_1276);
and ( n205113 , n205111 , n205112 );
nor ( n205114 , n205110 , n205113 );
buf ( n205115 , RI19a84e00_2760);
nand ( n205116 , n204493 , n205115 );
buf ( n205117 , RI17507628_743);
and ( n205118 , n205116 , n205117 );
not ( n205119 , n205116 );
not ( n205120 , RI17507628_743);
and ( n205121 , n205119 , n205120 );
nor ( n205122 , n205118 , n205121 );
xor ( n205123 , n205114 , n205122 );
buf ( n205124 , n25914 );
buf ( n205125 , RI19aa3aa8_2540);
nand ( n205126 , n205124 , n205125 );
buf ( n205127 , RI17482de8_1098);
and ( n205128 , n205126 , n205127 );
not ( n205129 , n205126 );
not ( n205130 , RI17482de8_1098);
and ( n205131 , n205129 , n205130 );
nor ( n205132 , n205128 , n205131 );
buf ( n205133 , n205132 );
xnor ( n205134 , n205123 , n205133 );
not ( n205135 , n205134 );
or ( n205136 , n205099 , n205135 );
or ( n205137 , n205134 , n205098 );
nand ( n205138 , n205136 , n205137 );
not ( n205139 , n205138 );
or ( n205140 , n205097 , n205139 );
not ( n205141 , n205138 );
not ( n205142 , n205095 );
not ( n205143 , n205142 );
nand ( n205144 , n205141 , n205143 );
nand ( n205145 , n205140 , n205144 );
not ( n205146 , n205145 );
nand ( n205147 , n205077 , n205146 );
not ( n205148 , n205147 );
not ( n205149 , RI173a3018_1961);
not ( n205150 , n205149 );
buf ( n205151 , RI173dd0c8_1678);
not ( n205152 , n205151 );
not ( n205153 , RI173943d8_2033);
not ( n205154 , n205153 );
or ( n205155 , n205152 , n205154 );
not ( n205156 , RI173dd0c8_1678);
buf ( n205157 , RI173943d8_2033);
nand ( n205158 , n205156 , n205157 );
nand ( n205159 , n205155 , n205158 );
not ( n205160 , n205159 );
or ( n205161 , n205150 , n205160 );
or ( n205162 , n205159 , n205149 );
nand ( n205163 , n205161 , n205162 );
not ( n205164 , n205163 );
buf ( n205165 , RI17454ba0_1323);
buf ( n205166 , RI19a96290_2639);
nand ( n205167 , n25451 , n205166 );
buf ( n205168 , RI174796f8_1144);
and ( n205169 , n205167 , n205168 );
not ( n205170 , n205167 );
not ( n205171 , RI174796f8_1144);
and ( n205172 , n205170 , n205171 );
nor ( n205173 , n205169 , n205172 );
xor ( n205174 , n205165 , n205173 );
xnor ( n205175 , n205174 , n204401 );
not ( n205176 , n205175 );
not ( n205177 , n205176 );
or ( n205178 , n205164 , n205177 );
or ( n205179 , n205176 , n205163 );
nand ( n205180 , n205178 , n205179 );
buf ( n205181 , RI173b1910_1890);
not ( n205182 , n205181 );
not ( n205183 , RI173fa600_1535);
not ( n205184 , n205183 );
or ( n205185 , n205182 , n205184 );
not ( n205186 , RI173b1910_1890);
buf ( n205187 , RI173fa600_1535);
nand ( n205188 , n205186 , n205187 );
nand ( n205189 , n205185 , n205188 );
not ( n205190 , RI173971c8_2019);
and ( n205191 , n205189 , n205190 );
not ( n205192 , n205189 );
buf ( n205193 , RI173971c8_2019);
and ( n205194 , n205192 , n205193 );
nor ( n205195 , n205191 , n205194 );
buf ( n205196 , RI19a9e6c0_2581);
nand ( n205197 , n25583 , n205196 );
buf ( n205198 , RI17526a50_646);
and ( n205199 , n205197 , n205198 );
not ( n205200 , n205197 );
not ( n205201 , RI17526a50_646);
and ( n205202 , n205200 , n205201 );
nor ( n205203 , n205199 , n205202 );
xor ( n205204 , n205195 , n205203 );
buf ( n205205 , RI19aa9f70_2496);
nand ( n205206 , n25752 , n205205 );
not ( n205207 , RI17496c30_1001);
and ( n205208 , n205206 , n205207 );
not ( n205209 , n205206 );
buf ( n205210 , RI17496c30_1001);
and ( n205211 , n205209 , n205210 );
nor ( n205212 , n205208 , n205211 );
xnor ( n205213 , n205204 , n205212 );
not ( n205214 , n205213 );
buf ( n205215 , n205214 );
not ( n205216 , n205215 );
and ( n205217 , n205180 , n205216 );
not ( n205218 , n205180 );
buf ( n205219 , n205213 );
not ( n205220 , n205219 );
buf ( n205221 , n205220 );
and ( n205222 , n205218 , n205221 );
or ( n205223 , n205217 , n205222 );
buf ( n205224 , n205223 );
not ( n205225 , n205224 );
and ( n205226 , n205148 , n205225 );
and ( n205227 , n205147 , n205224 );
nor ( n205228 , n205226 , n205227 );
not ( n205229 , n205228 );
not ( n205230 , n25866 );
not ( n205231 , n205230 );
buf ( n205232 , RI174a2dc8_942);
not ( n205233 , n205232 );
xor ( n205234 , n25792 , n25811 );
not ( n205235 , n25801 );
xor ( n205236 , n205234 , n205235 );
not ( n205237 , n205236 );
or ( n205238 , n205233 , n205237 );
not ( n205239 , n205232 );
nand ( n205240 , n205239 , n25813 );
nand ( n205241 , n205238 , n205240 );
not ( n205242 , n205241 );
and ( n205243 , n205231 , n205242 );
and ( n205244 , n205230 , n205241 );
nor ( n205245 , n205243 , n205244 );
not ( n205246 , n205245 );
buf ( n205247 , RI173cf190_1746);
not ( n205248 , n205247 );
not ( n205249 , RI173458c8_2102);
not ( n205250 , n205249 );
or ( n205251 , n205248 , n205250 );
not ( n205252 , RI173cf190_1746);
buf ( n205253 , RI173458c8_2102);
nand ( n205254 , n205252 , n205253 );
nand ( n205255 , n205251 , n205254 );
buf ( n205256 , RI17446c80_1391);
and ( n205257 , n205255 , n205256 );
not ( n205258 , n205255 );
not ( n205259 , RI17446c80_1391);
and ( n205260 , n205258 , n205259 );
nor ( n205261 , n205257 , n205260 );
buf ( n205262 , RI19a8c6f0_2708);
nand ( n205263 , n204916 , n205262 );
not ( n205264 , RI1746b490_1213);
and ( n205265 , n205263 , n205264 );
not ( n205266 , n205263 );
buf ( n205267 , RI1746b490_1213);
and ( n205268 , n205266 , n205267 );
nor ( n205269 , n205265 , n205268 );
xor ( n205270 , n205261 , n205269 );
buf ( n205271 , n26453 );
buf ( n205272 , RI19abd9f8_2353);
nand ( n205273 , n205271 , n205272 );
not ( n205274 , RI174b4168_858);
and ( n205275 , n205273 , n205274 );
not ( n205276 , n205273 );
buf ( n205277 , RI174b4168_858);
and ( n205278 , n205276 , n205277 );
nor ( n205279 , n205275 , n205278 );
xnor ( n205280 , n205270 , n205279 );
not ( n205281 , n205280 );
not ( n205282 , n205281 );
not ( n205283 , n205282 );
buf ( n205284 , RI173dd758_1676);
not ( n205285 , n205284 );
and ( n205286 , n205283 , n205285 );
and ( n205287 , n205282 , n205284 );
nor ( n205288 , n205286 , n205287 );
buf ( n205289 , RI173a39f0_1958);
not ( n205290 , n205289 );
not ( n205291 , RI173ec6e0_1603);
not ( n205292 , n205291 );
or ( n205293 , n205290 , n205292 );
not ( n205294 , RI173a39f0_1958);
buf ( n205295 , RI173ec6e0_1603);
nand ( n205296 , n205294 , n205295 );
nand ( n205297 , n205293 , n205296 );
buf ( n205298 , RI17480d18_1108);
and ( n205299 , n205297 , n205298 );
not ( n205300 , n205297 );
not ( n205301 , RI17480d18_1108);
and ( n205302 , n205300 , n205301 );
nor ( n205303 , n205299 , n205302 );
buf ( n205304 , RI19acf428_2216);
nand ( n205305 , n26242 , n205304 );
buf ( n205306 , RI17510688_715);
and ( n205307 , n205305 , n205306 );
not ( n205308 , n205305 );
not ( n205309 , RI17510688_715);
and ( n205310 , n205308 , n205309 );
nor ( n205311 , n205307 , n205310 );
xor ( n205312 , n205303 , n205311 );
buf ( n205313 , RI19aa0790_2565);
nand ( n205314 , n204426 , n205313 );
not ( n205315 , RI174889c8_1070);
and ( n205316 , n205314 , n205315 );
not ( n205317 , n205314 );
buf ( n205318 , RI174889c8_1070);
and ( n205319 , n205317 , n205318 );
nor ( n205320 , n205316 , n205319 );
xor ( n205321 , n205312 , n205320 );
buf ( n205322 , n205321 );
and ( n205323 , n205288 , n205322 );
not ( n205324 , n205288 );
not ( n205325 , n205322 );
and ( n205326 , n205324 , n205325 );
nor ( n205327 , n205323 , n205326 );
not ( n205328 , n205327 );
nand ( n205329 , n205246 , n205328 );
buf ( n205330 , RI1733c1d8_2148);
not ( n205331 , n205330 );
not ( n205332 , RI173cb680_1764);
buf ( n205333 , RI173b6b18_1865);
not ( n205334 , n205333 );
not ( n205335 , RI173ffb50_1509);
not ( n205336 , n205335 );
or ( n205337 , n205334 , n205336 );
not ( n205338 , RI173b6b18_1865);
buf ( n205339 , RI173ffb50_1509);
nand ( n205340 , n205338 , n205339 );
nand ( n205341 , n205337 , n205340 );
not ( n205342 , n205341 );
xor ( n205343 , n205332 , n205342 );
buf ( n205344 , RI1752eb38_621);
buf ( n205345 , RI1749be38_976);
xor ( n205346 , n205344 , n205345 );
buf ( n205347 , RI19ab9c18_2382);
nand ( n205348 , n205271 , n205347 );
xnor ( n205349 , n205346 , n205348 );
xnor ( n205350 , n205343 , n205349 );
not ( n205351 , n205350 );
or ( n205352 , n205331 , n205351 );
or ( n205353 , n205350 , n205330 );
nand ( n205354 , n205352 , n205353 );
buf ( n205355 , RI173d43b0_1721);
not ( n205356 , n205355 );
not ( n205357 , RI1738b6c0_2076);
not ( n205358 , n205357 );
or ( n205359 , n205356 , n205358 );
not ( n205360 , RI173d43b0_1721);
buf ( n205361 , RI1738b6c0_2076);
nand ( n205362 , n205360 , n205361 );
nand ( n205363 , n205359 , n205362 );
not ( n205364 , RI1744be88_1366);
and ( n205365 , n205363 , n205364 );
not ( n205366 , n205363 );
buf ( n205367 , RI1744be88_1366);
and ( n205368 , n205366 , n205367 );
nor ( n205369 , n205365 , n205368 );
buf ( n205370 , RI19a9c848_2594);
nand ( n205371 , n26242 , n205370 );
buf ( n205372 , RI17470698_1188);
xor ( n205373 , n205371 , n205372 );
xor ( n205374 , n205369 , n205373 );
buf ( n205375 , RI19acba08_2242);
nand ( n205376 , n205020 , n205375 );
not ( n205377 , RI174b9988_833);
and ( n205378 , n205376 , n205377 );
not ( n205379 , n205376 );
buf ( n205380 , RI174b9988_833);
and ( n205381 , n205379 , n205380 );
nor ( n205382 , n205378 , n205381 );
xnor ( n205383 , n205374 , n205382 );
not ( n205384 , n205383 );
buf ( n205385 , n205384 );
not ( n205386 , n205385 );
and ( n205387 , n205354 , n205386 );
not ( n205388 , n205354 );
not ( n205389 , n205383 );
and ( n205390 , n205388 , n205389 );
nor ( n205391 , n205387 , n205390 );
not ( n205392 , n205391 );
not ( n205393 , n205392 );
and ( n205394 , n205329 , n205393 );
not ( n205395 , n205329 );
and ( n205396 , n205395 , n205392 );
nor ( n205397 , n205394 , n205396 );
not ( n205398 , n205397 );
or ( n205399 , n205229 , n205398 );
or ( n205400 , n205397 , n205228 );
nand ( n205401 , n205399 , n205400 );
buf ( n205402 , RI17450d48_1342);
buf ( n205403 , RI17408520_1467);
not ( n205404 , n205403 );
not ( n205405 , RI173bf830_1822);
not ( n205406 , n205405 );
or ( n205407 , n205404 , n205406 );
not ( n205408 , RI17408520_1467);
buf ( n205409 , RI173bf830_1822);
nand ( n205410 , n205408 , n205409 );
nand ( n205411 , n205407 , n205410 );
xor ( n205412 , n205402 , n205411 );
not ( n205413 , RI173362b0_2177);
buf ( n205414 , RI174a4808_934);
xor ( n205415 , n205413 , n205414 );
buf ( n205416 , RI19ab34f8_2429);
nand ( n205417 , n25793 , n205416 );
xnor ( n205418 , n205415 , n205417 );
xnor ( n205419 , n205412 , n205418 );
buf ( n205420 , n205419 );
not ( n205421 , n205420 );
not ( n205422 , n205421 );
buf ( n205423 , RI173ce470_1750);
not ( n205424 , n205423 );
and ( n205425 , n205422 , n205424 );
not ( n205426 , n205420 );
and ( n205427 , n205426 , n205423 );
nor ( n27667 , n205425 , n205427 );
not ( n27668 , n204279 );
not ( n27669 , n204306 );
or ( n27670 , n27668 , n27669 );
not ( n205432 , n204279 );
nand ( n205433 , n205432 , n204305 );
nand ( n205434 , n27670 , n205433 );
buf ( n205435 , n205434 );
not ( n205436 , n205435 );
and ( n27676 , n27667 , n205436 );
not ( n27677 , n27667 );
and ( n27678 , n27677 , n205435 );
nor ( n27679 , n27676 , n27678 );
not ( n27680 , n27679 );
buf ( n27681 , RI1744b7f8_1368);
not ( n27682 , n27681 );
buf ( n27683 , RI173c5410_1794);
not ( n205445 , n27683 );
not ( n205446 , RI1733be90_2149);
not ( n27686 , n205446 );
or ( n27687 , n205445 , n27686 );
not ( n27688 , RI173c5410_1794);
nand ( n27689 , n27688 , n25434 );
nand ( n205451 , n27687 , n27689 );
not ( n27691 , RI1740e100_1439);
and ( n205453 , n205451 , n27691 );
not ( n27693 , n205451 );
buf ( n27694 , RI1740e100_1439);
and ( n27695 , n27693 , n27694 );
nor ( n27696 , n205453 , n27695 );
buf ( n27697 , RI19a922d0_2667);
nand ( n27698 , n25711 , n27697 );
buf ( n27699 , RI17461a58_1260);
and ( n27700 , n27698 , n27699 );
not ( n27701 , n27698 );
not ( n27702 , RI17461a58_1260);
and ( n205464 , n27701 , n27702 );
nor ( n27704 , n27700 , n205464 );
xor ( n205466 , n27696 , n27704 );
buf ( n27706 , n204336 );
buf ( n27707 , RI19ac25e8_2311);
nand ( n27708 , n27706 , n27707 );
not ( n27709 , RI174aa730_905);
and ( n27710 , n27708 , n27709 );
not ( n27711 , n27708 );
buf ( n27712 , RI174aa730_905);
and ( n27713 , n27711 , n27712 );
nor ( n27714 , n27710 , n27713 );
xnor ( n205476 , n205466 , n27714 );
buf ( n27716 , n205476 );
not ( n205478 , n27716 );
or ( n27718 , n27682 , n205478 );
not ( n205480 , n27704 );
xor ( n27720 , n27696 , n205480 );
xnor ( n27721 , n27720 , n27714 );
not ( n27722 , RI1744b7f8_1368);
nand ( n27723 , n27721 , n27722 );
nand ( n27724 , n27718 , n27723 );
buf ( n27725 , RI173e2960_1651);
not ( n27726 , n27725 );
not ( n27727 , RI17399c70_2006);
not ( n27728 , n27727 );
or ( n205490 , n27726 , n27728 );
not ( n27730 , RI173e2960_1651);
buf ( n205492 , RI17399c70_2006);
nand ( n27732 , n27730 , n205492 );
nand ( n27733 , n205490 , n27732 );
not ( n27734 , RI1745a780_1295);
and ( n27735 , n27733 , n27734 );
not ( n27736 , n27733 );
buf ( n27737 , RI1745a780_1295);
and ( n27738 , n27736 , n27737 );
nor ( n27739 , n27735 , n27738 );
buf ( n27740 , RI19a87218_2744);
nand ( n27741 , n25741 , n27740 );
buf ( n27742 , RI174d07a0_762);
and ( n205504 , n27741 , n27742 );
not ( n27744 , n27741 );
not ( n205506 , RI174d07a0_762);
and ( n27746 , n27744 , n205506 );
nor ( n27747 , n205504 , n27746 );
xor ( n27748 , n27739 , n27747 );
buf ( n27749 , n25741 );
buf ( n27750 , RI19aa5fb0_2523);
nand ( n27751 , n27749 , n27750 );
buf ( n27752 , RI1747ef90_1117);
and ( n27753 , n27751 , n27752 );
not ( n27754 , n27751 );
not ( n205516 , RI1747ef90_1117);
and ( n27756 , n27754 , n205516 );
nor ( n205518 , n27753 , n27756 );
xnor ( n27758 , n27748 , n205518 );
not ( n27759 , n27758 );
and ( n27760 , n27724 , n27759 );
not ( n27761 , n27724 );
not ( n27762 , n27758 );
not ( n27763 , n27762 );
and ( n27764 , n27761 , n27763 );
nor ( n27765 , n27760 , n27764 );
not ( n27766 , n27765 );
nand ( n27767 , n27680 , n27766 );
not ( n27768 , n27767 );
buf ( n27769 , RI173ce128_1751);
not ( n205531 , n27769 );
not ( n27771 , RI17344860_2107);
not ( n205533 , n27771 );
or ( n27773 , n205531 , n205533 );
not ( n27774 , RI173ce128_1751);
buf ( n27775 , RI17344860_2107);
nand ( n27776 , n27774 , n27775 );
nand ( n27777 , n27773 , n27776 );
not ( n27778 , RI17445c18_1396);
and ( n27779 , n27777 , n27778 );
not ( n27780 , n27777 );
buf ( n27781 , RI17445c18_1396);
and ( n205543 , n27780 , n27781 );
nor ( n27783 , n27779 , n205543 );
buf ( n205545 , RI19a8bbb0_2713);
nand ( n27785 , n26242 , n205545 );
buf ( n27786 , RI1746a428_1218);
and ( n27787 , n27785 , n27786 );
not ( n27788 , n27785 );
not ( n27789 , RI1746a428_1218);
and ( n27790 , n27788 , n27789 );
nor ( n27791 , n27787 , n27790 );
xor ( n27792 , n27783 , n27791 );
buf ( n27793 , RI19abd188_2358);
nand ( n27794 , n25416 , n27793 );
not ( n27795 , RI174b3100_863);
and ( n27796 , n27794 , n27795 );
not ( n27797 , n27794 );
buf ( n205559 , RI174b3100_863);
and ( n27799 , n27797 , n205559 );
nor ( n205561 , n27796 , n27799 );
xor ( n27801 , n27792 , n205561 );
not ( n27802 , n27801 );
not ( n27803 , n27802 );
buf ( n27804 , RI173bf1a0_1824);
not ( n27805 , n27804 );
buf ( n27806 , RI19aabb90_2484);
nand ( n27807 , n204572 , n27806 );
buf ( n27808 , RI17495bc8_1006);
and ( n27809 , n27807 , n27808 );
not ( n205571 , n27807 );
not ( n27811 , RI17495bc8_1006);
and ( n205573 , n205571 , n27811 );
nor ( n27813 , n27809 , n205573 );
not ( n27814 , n27813 );
buf ( n27815 , RI19aaf448_2459);
nand ( n27816 , n25915 , n27815 );
not ( n27817 , RI17525088_651);
and ( n27818 , n27816 , n27817 );
not ( n27819 , n27816 );
buf ( n27820 , RI17525088_651);
and ( n27821 , n27819 , n27820 );
nor ( n205583 , n27818 , n27821 );
not ( n27823 , n205583 );
or ( n205585 , n27814 , n27823 );
or ( n27825 , n27813 , n205583 );
nand ( n205587 , n205585 , n27825 );
buf ( n27827 , RI173f9598_1540);
not ( n27828 , n27827 );
not ( n27829 , RI173b08a8_1895);
not ( n27830 , n27829 );
or ( n27831 , n27828 , n27830 );
not ( n27832 , RI173f9598_1540);
buf ( n27833 , RI173b08a8_1895);
nand ( n27834 , n27832 , n27833 );
nand ( n27835 , n27831 , n27834 );
not ( n205597 , RI1738bd50_2074);
and ( n27837 , n27835 , n205597 );
not ( n27838 , n27835 );
buf ( n27839 , RI1738bd50_2074);
and ( n27840 , n27838 , n27839 );
nor ( n27841 , n27837 , n27840 );
xor ( n27842 , n205587 , n27841 );
not ( n27843 , n27842 );
or ( n27844 , n27805 , n27843 );
not ( n27845 , n205583 );
xor ( n27846 , n27841 , n27845 );
buf ( n27847 , n27813 );
xnor ( n27848 , n27846 , n27847 );
not ( n205610 , RI173bf1a0_1824);
nand ( n27850 , n27848 , n205610 );
nand ( n205612 , n27844 , n27850 );
not ( n27852 , n205612 );
or ( n27853 , n27803 , n27852 );
or ( n27854 , n205612 , n27802 );
nand ( n27855 , n27853 , n27854 );
not ( n27856 , n27855 );
and ( n27857 , n27768 , n27856 );
and ( n27858 , n27767 , n27855 );
nor ( n27859 , n27857 , n27858 );
and ( n27860 , n205401 , n27859 );
not ( n205622 , n205401 );
not ( n27862 , n27859 );
and ( n205624 , n205622 , n27862 );
nor ( n27864 , n27860 , n205624 );
not ( n27865 , n27864 );
not ( n27866 , n27865 );
or ( n27867 , n204992 , n27866 );
nand ( n27868 , n27864 , n204990 );
nand ( n27869 , n27867 , n27868 );
buf ( n27870 , n27869 );
and ( n27871 , n204555 , n27870 );
not ( n27872 , n204555 );
and ( n27873 , n27864 , n204990 );
not ( n27874 , n27864 );
and ( n27875 , n27874 , n204991 );
nor ( n27876 , n27873 , n27875 );
not ( n205638 , n27876 );
not ( n27878 , n205638 );
and ( n27879 , n27872 , n27878 );
nor ( n27880 , n27871 , n27879 );
buf ( n27881 , n25358 );
nor ( n27882 , n204514 , n27881 );
not ( n27883 , RI1754c610_2);
not ( n27884 , n27883 );
or ( n27885 , n27882 , n27884 );
buf ( n27886 , n27885 );
not ( n27887 , n27886 );
buf ( n205649 , n27887 );
not ( n27889 , n205649 );
nor ( n205651 , n27880 , n27889 );
buf ( n27891 , RI173fee30_1513);
not ( n27892 , n27891 );
not ( n27893 , RI173b5df8_1869);
not ( n27894 , n27893 );
or ( n27895 , n27892 , n27894 );
not ( n27896 , RI173fee30_1513);
buf ( n27897 , RI173b5df8_1869);
nand ( n27898 , n27896 , n27897 );
nand ( n27899 , n27895 , n27898 );
not ( n205661 , n27899 );
not ( n27901 , n205661 );
buf ( n205663 , RI173c2620_1808);
buf ( n27903 , RI1749b118_980);
not ( n27904 , n27903 );
buf ( n27905 , RI19aa7e28_2510);
nand ( n27906 , n25416 , n27905 );
not ( n27907 , n27906 );
or ( n27908 , n27904 , n27907 );
not ( n27909 , RI1749b118_980);
nand ( n27910 , n25479 , n27909 , n27905 );
nand ( n27911 , n27908 , n27910 );
xor ( n205673 , n205663 , n27911 );
buf ( n27913 , RI19a89e28_2725);
nand ( n205675 , n25405 , n27913 );
not ( n27915 , RI1752d698_625);
and ( n27916 , n205675 , n27915 );
not ( n27917 , n205675 );
buf ( n27918 , RI1752d698_625);
and ( n27919 , n27917 , n27918 );
nor ( n27920 , n27916 , n27919 );
xnor ( n27921 , n205673 , n27920 );
not ( n27922 , n27921 );
not ( n27923 , n27922 );
or ( n27924 , n27901 , n27923 );
nand ( n205686 , n27921 , n27899 );
nand ( n27926 , n27924 , n205686 );
not ( n205688 , n27926 );
not ( n27928 , n205688 );
buf ( n205690 , RI173a7500_1940);
not ( n27930 , n205690 );
buf ( n27931 , RI173988c0_2012);
not ( n27932 , n27931 );
not ( n27933 , RI173e15b0_1657);
not ( n27934 , n27933 );
or ( n27935 , n27932 , n27934 );
not ( n27936 , RI173988c0_2012);
buf ( n27937 , RI173e15b0_1657);
nand ( n27938 , n27936 , n27937 );
nand ( n205700 , n27935 , n27938 );
not ( n27940 , RI174593d0_1301);
and ( n205702 , n205700 , n27940 );
not ( n27942 , n205700 );
buf ( n27943 , RI174593d0_1301);
and ( n27944 , n27942 , n27943 );
nor ( n27945 , n205702 , n27944 );
buf ( n27946 , n25363 );
buf ( n27947 , RI19a93fe0_2654);
nand ( n27948 , n27946 , n27947 );
buf ( n27949 , RI1747dbe0_1123);
xor ( n27950 , n27948 , n27949 );
xor ( n27951 , n27945 , n27950 );
buf ( n27952 , RI19ac4280_2298);
nand ( n27953 , n27706 , n27952 );
not ( n27954 , RI174ce8b0_768);
and ( n205716 , n27953 , n27954 );
not ( n27956 , n27953 );
buf ( n205718 , RI174ce8b0_768);
and ( n27958 , n27956 , n205718 );
nor ( n27959 , n205716 , n27958 );
xnor ( n27960 , n27951 , n27959 );
buf ( n27961 , n27960 );
not ( n27962 , n27961 );
or ( n27963 , n27930 , n27962 );
or ( n27964 , n27961 , n205690 );
nand ( n27965 , n27963 , n27964 );
not ( n27966 , n27965 );
and ( n205728 , n27928 , n27966 );
buf ( n27968 , n205688 );
and ( n27969 , n27968 , n27965 );
nor ( n27970 , n205728 , n27969 );
not ( n27971 , n27970 );
buf ( n27972 , RI17459a60_1299);
buf ( n27973 , RI17398f50_2010);
not ( n27974 , n27973 );
not ( n27975 , RI173e1c40_1655);
not ( n27976 , n27975 );
or ( n27977 , n27974 , n27976 );
not ( n205739 , RI17398f50_2010);
buf ( n27979 , RI173e1c40_1655);
nand ( n205741 , n205739 , n27979 );
nand ( n27981 , n27977 , n205741 );
xor ( n205743 , n27972 , n27981 );
buf ( n27983 , RI19a869a8_2748);
nand ( n27984 , n25539 , n27983 );
buf ( n27985 , RI174cf300_766);
and ( n27986 , n27984 , n27985 );
not ( n27987 , n27984 );
not ( n27988 , RI174cf300_766);
and ( n27989 , n27987 , n27988 );
nor ( n27990 , n27986 , n27989 );
not ( n27991 , n27990 );
buf ( n205753 , RI19aa5560_2527);
nand ( n27993 , n25529 , n205753 );
not ( n205755 , RI1747e270_1121);
and ( n27995 , n27993 , n205755 );
not ( n27996 , n27993 );
buf ( n27997 , RI1747e270_1121);
and ( n27998 , n27996 , n27997 );
nor ( n27999 , n27995 , n27998 );
not ( n28000 , n27999 );
or ( n28001 , n27991 , n28000 );
or ( n28002 , n27990 , n27999 );
nand ( n28003 , n28001 , n28002 );
xnor ( n28004 , n205743 , n28003 );
not ( n205766 , n28004 );
buf ( n28006 , RI173d3348_1726);
not ( n205768 , n28006 );
not ( n28008 , RI1738a658_2081);
not ( n28009 , n28008 );
or ( n28010 , n205768 , n28009 );
not ( n28011 , RI173d3348_1726);
buf ( n28012 , RI1738a658_2081);
nand ( n28013 , n28011 , n28012 );
nand ( n28014 , n28010 , n28013 );
buf ( n28015 , RI1744ae20_1371);
and ( n28016 , n28014 , n28015 );
not ( n28017 , n28014 );
not ( n205779 , RI1744ae20_1371);
and ( n28019 , n28017 , n205779 );
nor ( n205781 , n28016 , n28019 );
xor ( n28021 , n205781 , n204453 );
buf ( n28022 , RI19abbe50_2368);
nand ( n28023 , n25452 , n28022 );
not ( n28024 , RI174b8308_838);
and ( n28025 , n28023 , n28024 );
not ( n28026 , n28023 );
buf ( n28027 , RI174b8308_838);
and ( n28028 , n28026 , n28027 );
nor ( n28029 , n28025 , n28028 );
xnor ( n28030 , n28021 , n28029 );
not ( n28031 , n28030 );
buf ( n28032 , RI19ac4460_2297);
nand ( n28033 , n26453 , n28032 );
buf ( n205795 , RI174cedd8_767);
and ( n28035 , n28033 , n205795 );
not ( n205797 , n28033 );
not ( n28037 , RI174cedd8_767);
and ( n28038 , n205797 , n28037 );
nor ( n28039 , n28035 , n28038 );
buf ( n28040 , n28039 );
not ( n28041 , n28040 );
and ( n28042 , n28031 , n28041 );
not ( n28043 , n28030 );
not ( n28044 , n28043 );
and ( n28045 , n28044 , n28040 );
nor ( n205807 , n28042 , n28045 );
not ( n28047 , n205807 );
and ( n205809 , n205766 , n28047 );
not ( n28049 , n205766 );
and ( n28050 , n28049 , n205807 );
nor ( n28051 , n205809 , n28050 );
not ( n28052 , n28051 );
nand ( n28053 , n27971 , n28052 );
buf ( n28054 , RI173efea8_1586);
buf ( n28055 , RI17403660_1491);
not ( n28056 , n28055 );
not ( n28057 , RI173ba970_1846);
not ( n205819 , n28057 );
or ( n28059 , n28056 , n205819 );
not ( n205821 , RI17403660_1491);
buf ( n28061 , RI173ba970_1846);
nand ( n205823 , n205821 , n28061 );
nand ( n28063 , n28059 , n205823 );
xor ( n28064 , n28054 , n28063 );
not ( n28065 , RI1749f948_958);
xor ( n28066 , n25341 , n28065 );
buf ( n28067 , RI19ab7530_2399);
nand ( n28068 , n204426 , n28067 );
xnor ( n28069 , n28066 , n28068 );
xnor ( n28070 , n28064 , n28069 );
not ( n28071 , n28070 );
not ( n205833 , n28071 );
not ( n28073 , n205833 );
buf ( n205835 , RI19a8fd50_2684);
nand ( n28075 , n204926 , n205835 );
buf ( n28076 , RI17465568_1242);
and ( n28077 , n28075 , n28076 );
not ( n28078 , n28075 );
not ( n28079 , RI17465568_1242);
and ( n28080 , n28078 , n28079 );
nor ( n28081 , n28077 , n28080 );
buf ( n28082 , n28081 );
not ( n28083 , n28082 );
and ( n28084 , n28073 , n28083 );
not ( n205846 , n28071 );
and ( n28086 , n205846 , n28082 );
nor ( n205848 , n28084 , n28086 );
buf ( n28088 , RI1744f998_1348);
buf ( n205850 , RI19a9a160_2611);
nand ( n28090 , n25628 , n205850 );
buf ( n28091 , RI174741a8_1170);
and ( n28092 , n28090 , n28091 );
not ( n28093 , n28090 );
not ( n28094 , RI174741a8_1170);
and ( n28095 , n28093 , n28094 );
nor ( n28096 , n28092 , n28095 );
xor ( n28097 , n28088 , n28096 );
buf ( n28098 , RI19ac9938_2258);
nand ( n205860 , n25851 , n28098 );
not ( n28100 , RI174bfb80_814);
and ( n28101 , n205860 , n28100 );
not ( n28102 , n205860 );
buf ( n28103 , RI174bfb80_814);
and ( n28104 , n28102 , n28103 );
nor ( n28105 , n28101 , n28104 );
xnor ( n28106 , n28097 , n28105 );
not ( n28107 , n28106 );
buf ( n28108 , RI173d7ec0_1703);
not ( n28109 , n28108 );
not ( n28110 , RI1738f1d0_2058);
not ( n28111 , n28110 );
or ( n28112 , n28109 , n28111 );
not ( n28113 , RI173d7ec0_1703);
buf ( n205875 , RI1738f1d0_2058);
nand ( n28115 , n28113 , n205875 );
nand ( n205877 , n28112 , n28115 );
not ( n28117 , n205877 );
not ( n205879 , n28117 );
and ( n28119 , n28107 , n205879 );
and ( n28120 , n28106 , n28117 );
nor ( n28121 , n28119 , n28120 );
buf ( n28122 , n28121 );
and ( n28123 , n205848 , n28122 );
not ( n28124 , n205848 );
not ( n28125 , n28122 );
and ( n28126 , n28124 , n28125 );
nor ( n28127 , n28123 , n28126 );
buf ( n205889 , n28127 );
xnor ( n28129 , n28053 , n205889 );
not ( n205891 , n28129 );
not ( n28131 , RI17460d38_1264);
not ( n28132 , RI17409f60_1459);
buf ( n28133 , RI173c1270_1814);
nand ( n28134 , n28132 , n28133 );
not ( n28135 , RI173c1270_1814);
buf ( n28136 , RI17409f60_1459);
nand ( n28137 , n28135 , n28136 );
and ( n28138 , n28134 , n28137 );
xor ( n28139 , n28131 , n28138 );
buf ( n28140 , RI17337cf0_2169);
buf ( n205902 , RI174a6590_925);
xor ( n28142 , n28140 , n205902 );
buf ( n28143 , RI19ab2148_2439);
nand ( n28144 , n25712 , n28143 );
xnor ( n28145 , n28142 , n28144 );
xnor ( n28146 , n28139 , n28145 );
not ( n28147 , n28146 );
buf ( n28148 , n25490 );
buf ( n28149 , RI19aaa510_2493);
nand ( n28150 , n28148 , n28149 );
buf ( n205912 , RI17497608_998);
and ( n28152 , n28150 , n205912 );
not ( n205914 , n28150 );
not ( n28154 , RI17497608_998);
and ( n28155 , n205914 , n28154 );
nor ( n28156 , n28152 , n28155 );
buf ( n28157 , n28156 );
not ( n28158 , n28157 );
buf ( n28159 , RI173eca28_1602);
not ( n28160 , n28159 );
not ( n28161 , RI173a3d38_1957);
not ( n28162 , n28161 );
or ( n28163 , n28160 , n28162 );
not ( n28164 , RI173eca28_1602);
buf ( n205926 , RI173a3d38_1957);
nand ( n28166 , n28164 , n205926 );
nand ( n205928 , n28163 , n28166 );
buf ( n28168 , RI17483130_1097);
and ( n28169 , n205928 , n28168 );
not ( n28170 , n205928 );
not ( n28171 , RI17483130_1097);
and ( n28172 , n28170 , n28171 );
nor ( n28173 , n28169 , n28172 );
buf ( n28174 , RI19acf680_2215);
nand ( n28175 , n25479 , n28174 );
buf ( n28176 , RI17510bb0_714);
xor ( n205938 , n28175 , n28176 );
xor ( n28178 , n28173 , n205938 );
buf ( n28179 , RI19aa0970_2564);
nand ( n28180 , n25452 , n28179 );
buf ( n28181 , RI17488d10_1069);
and ( n28182 , n28180 , n28181 );
not ( n28183 , n28180 );
not ( n28184 , RI17488d10_1069);
and ( n28185 , n28183 , n28184 );
nor ( n28186 , n28182 , n28185 );
not ( n28187 , n28186 );
xnor ( n28188 , n28178 , n28187 );
not ( n28189 , n28188 );
or ( n28190 , n28158 , n28189 );
or ( n205952 , n28188 , n28157 );
nand ( n28192 , n28190 , n205952 );
not ( n205954 , n28192 );
and ( n28194 , n28147 , n205954 );
and ( n28195 , n28146 , n28192 );
nor ( n28196 , n28194 , n28195 );
not ( n28197 , n27802 );
buf ( n28198 , RI17335c20_2179);
not ( n28199 , n28198 );
not ( n28200 , n27842 );
or ( n28201 , n28199 , n28200 );
not ( n28202 , RI17335c20_2179);
nand ( n205964 , n27848 , n28202 );
nand ( n28204 , n28201 , n205964 );
not ( n205966 , n28204 );
or ( n28206 , n28197 , n205966 );
or ( n28207 , n28204 , n27802 );
nand ( n28208 , n28206 , n28207 );
nand ( n28209 , n28196 , n28208 );
not ( n28210 , n28209 );
buf ( n28211 , RI1745d570_1281);
not ( n28212 , n28211 );
buf ( n28213 , RI173d71a0_1707);
not ( n28214 , n28213 );
not ( n28215 , RI1738e4b0_2062);
not ( n205977 , n28215 );
or ( n28217 , n28214 , n205977 );
not ( n28218 , RI173d71a0_1707);
buf ( n28219 , RI1738e4b0_2062);
nand ( n28220 , n28218 , n28219 );
nand ( n28221 , n28217 , n28220 );
buf ( n28222 , RI1744ec78_1352);
and ( n28223 , n28221 , n28222 );
not ( n28224 , n28221 );
not ( n28225 , RI1744ec78_1352);
and ( n28226 , n28224 , n28225 );
nor ( n205988 , n28223 , n28226 );
not ( n28228 , n205988 );
buf ( n205990 , RI19a99698_2616);
nand ( n28230 , n25850 , n205990 );
buf ( n28231 , RI17473488_1174);
and ( n28232 , n28230 , n28231 );
not ( n28233 , n28230 );
not ( n28234 , RI17473488_1174);
and ( n28235 , n28233 , n28234 );
nor ( n28236 , n28232 , n28235 );
xor ( n28237 , n28228 , n28236 );
buf ( n28238 , n25529 );
buf ( n28239 , RI19ac90c8_2262);
nand ( n28240 , n28238 , n28239 );
not ( n206002 , RI174be6e0_818);
and ( n28242 , n28240 , n206002 );
not ( n206004 , n28240 );
buf ( n28244 , RI174be6e0_818);
and ( n28245 , n206004 , n28244 );
nor ( n28246 , n28242 , n28245 );
xnor ( n28247 , n28237 , n28246 );
not ( n28248 , n28247 );
or ( n28249 , n28212 , n28248 );
xor ( n28250 , n205988 , n28236 );
xnor ( n28251 , n28250 , n28246 );
not ( n28252 , RI1745d570_1281);
nand ( n206014 , n28251 , n28252 );
nand ( n28254 , n28249 , n206014 );
not ( n206016 , n28254 );
buf ( n28256 , RI173f4390_1565);
not ( n28257 , n28256 );
not ( n28258 , RI173ab6a0_1920);
not ( n28259 , n28258 );
or ( n28260 , n28257 , n28259 );
not ( n28261 , RI173f4390_1565);
buf ( n28262 , RI173ab6a0_1920);
nand ( n28263 , n28261 , n28262 );
nand ( n28264 , n28260 , n28263 );
buf ( n28265 , RI1750ecc0_720);
and ( n28266 , n28264 , n28265 );
not ( n28267 , n28264 );
not ( n206029 , RI1750ecc0_720);
and ( n28269 , n28267 , n206029 );
nor ( n206031 , n28266 , n28269 );
buf ( n28271 , RI19abe2e0_2348);
nand ( n206033 , n25583 , n28271 );
buf ( n28273 , RI1751cfa0_676);
and ( n28274 , n206033 , n28273 );
not ( n28275 , n206033 );
not ( n28276 , RI1751cfa0_676);
and ( n28277 , n28275 , n28276 );
nor ( n28278 , n28274 , n28277 );
xor ( n28279 , n206031 , n28278 );
buf ( n28280 , RI19aad468_2473);
nand ( n28281 , n25540 , n28280 );
buf ( n206043 , RI174909c0_1031);
and ( n28283 , n28281 , n206043 );
not ( n206045 , n28281 );
not ( n28285 , RI174909c0_1031);
and ( n28286 , n206045 , n28285 );
nor ( n28287 , n28283 , n28286 );
xnor ( n28288 , n28279 , n28287 );
not ( n28289 , n28288 );
and ( n28290 , n206016 , n28289 );
and ( n28291 , n28254 , n28288 );
nor ( n28292 , n28290 , n28291 );
not ( n28293 , n28292 );
not ( n28294 , n28293 );
and ( n206056 , n28210 , n28294 );
and ( n28296 , n28209 , n28293 );
nor ( n206058 , n206056 , n28296 );
buf ( n28298 , RI19aa3238_2544);
nand ( n28299 , n25376 , n28298 );
not ( n28300 , RI174820c8_1102);
and ( n28301 , n28299 , n28300 );
not ( n28302 , n28299 );
buf ( n28303 , RI174820c8_1102);
and ( n28304 , n28302 , n28303 );
nor ( n28305 , n28301 , n28304 );
not ( n28306 , n28305 );
buf ( n28307 , RI173d74e8_1706);
not ( n28308 , n28307 );
not ( n28309 , RI1738e7f8_2061);
not ( n28310 , n28309 );
or ( n28311 , n28308 , n28310 );
not ( n28312 , RI173d74e8_1706);
buf ( n28313 , RI1738e7f8_2061);
nand ( n28314 , n28312 , n28313 );
nand ( n28315 , n28311 , n28314 );
not ( n28316 , RI1744efc0_1351);
and ( n28317 , n28315 , n28316 );
not ( n206079 , n28315 );
buf ( n28319 , RI1744efc0_1351);
and ( n206081 , n206079 , n28319 );
nor ( n28321 , n28317 , n206081 );
buf ( n28322 , RI19ac92a8_2261);
nand ( n28323 , n25915 , n28322 );
buf ( n28324 , RI174bec08_817);
and ( n28325 , n28323 , n28324 );
not ( n28326 , n28323 );
not ( n28327 , RI174bec08_817);
and ( n28328 , n28326 , n28327 );
nor ( n28329 , n28325 , n28328 );
xor ( n206091 , n28321 , n28329 );
buf ( n28331 , RI19a998f0_2615);
nand ( n206093 , n26276 , n28331 );
buf ( n28333 , RI174737d0_1173);
and ( n28334 , n206093 , n28333 );
not ( n28335 , n206093 );
not ( n28336 , RI174737d0_1173);
and ( n28337 , n28335 , n28336 );
nor ( n28338 , n28334 , n28337 );
xor ( n28339 , n206091 , n28338 );
buf ( n28340 , n28339 );
not ( n28341 , n28340 );
or ( n28342 , n28306 , n28341 );
not ( n28343 , n28305 );
not ( n28344 , n28339 );
nand ( n206106 , n28343 , n28344 );
nand ( n28346 , n28342 , n206106 );
not ( n206108 , n28346 );
buf ( n28348 , RI173f4a20_1563);
not ( n28349 , n28348 );
not ( n28350 , RI173abd30_1918);
not ( n28351 , n28350 );
or ( n28352 , n28349 , n28351 );
not ( n28353 , RI173f4a20_1563);
buf ( n28354 , RI173abd30_1918);
nand ( n28355 , n28353 , n28354 );
nand ( n28356 , n28352 , n28355 );
buf ( n28357 , RI17512aa0_708);
and ( n206119 , n28356 , n28357 );
not ( n28359 , n28356 );
not ( n206121 , RI17512aa0_708);
and ( n28361 , n28359 , n206121 );
nor ( n28362 , n206119 , n28361 );
buf ( n28363 , RI19abf690_2337);
nand ( n28364 , n26242 , n28363 );
buf ( n28365 , RI1751d9f0_674);
and ( n28366 , n28364 , n28365 );
not ( n28367 , n28364 );
not ( n28368 , RI1751d9f0_674);
and ( n28369 , n28367 , n28368 );
nor ( n28370 , n28366 , n28369 );
xor ( n206132 , n28362 , n28370 );
buf ( n28372 , RI19aad648_2472);
nand ( n206134 , n204393 , n28372 );
buf ( n28374 , RI17491050_1029);
and ( n28375 , n206134 , n28374 );
not ( n28376 , n206134 );
not ( n28377 , RI17491050_1029);
and ( n28378 , n28376 , n28377 );
nor ( n28379 , n28375 , n28378 );
xnor ( n28380 , n206132 , n28379 );
not ( n28381 , n28380 );
not ( n28382 , n28381 );
not ( n206144 , n28382 );
and ( n28384 , n206108 , n206144 );
and ( n206146 , n28346 , n28382 );
nor ( n28386 , n28384 , n206146 );
buf ( n28387 , RI173ddaa0_1675);
buf ( n28388 , RI174018d8_1500);
not ( n28389 , n28388 );
not ( n28390 , RI173b8be8_1855);
not ( n28391 , n28390 );
or ( n28392 , n28389 , n28391 );
not ( n28393 , RI174018d8_1500);
buf ( n28394 , RI173b8be8_1855);
nand ( n28395 , n28393 , n28394 );
nand ( n28396 , n28392 , n28395 );
xor ( n206158 , n28387 , n28396 );
buf ( n28398 , RI175319a0_612);
buf ( n206160 , RI1749dbc0_967);
xor ( n28400 , n28398 , n206160 );
buf ( n28401 , RI19ab8b38_2390);
nand ( n28402 , n25916 , n28401 );
xnor ( n28403 , n28400 , n28402 );
xnor ( n28404 , n206158 , n28403 );
buf ( n28405 , n28404 );
not ( n28406 , n28405 );
buf ( n28407 , RI19a23678_2793);
nand ( n28408 , n205271 , n28407 );
not ( n206170 , RI1751ab88_683);
and ( n28410 , n28408 , n206170 );
not ( n206172 , n28408 );
buf ( n28412 , RI1751ab88_683);
and ( n28413 , n206172 , n28412 );
nor ( n28414 , n28410 , n28413 );
not ( n28415 , n28414 );
not ( n28416 , n26308 );
or ( n28417 , n28415 , n28416 );
not ( n28418 , n28414 );
nand ( n28419 , n28418 , n26317 );
nand ( n28420 , n28417 , n28419 );
not ( n28421 , n28420 );
and ( n28422 , n28406 , n28421 );
and ( n28423 , n28405 , n28420 );
nor ( n206185 , n28422 , n28423 );
not ( n28425 , n206185 );
nand ( n28426 , n28386 , n28425 );
buf ( n28427 , RI1744fce0_1347);
not ( n28428 , n28427 );
buf ( n206190 , RI173c98f8_1773);
not ( n28430 , n206190 );
not ( n206192 , RI17340378_2128);
not ( n28432 , n206192 );
or ( n28433 , n28430 , n28432 );
not ( n28434 , RI173c98f8_1773);
buf ( n28435 , RI17340378_2128);
nand ( n28436 , n28434 , n28435 );
nand ( n28437 , n28433 , n28436 );
buf ( n28438 , RI17412930_1417);
and ( n28439 , n28437 , n28438 );
not ( n28440 , n28437 );
not ( n206202 , RI17412930_1417);
and ( n28442 , n28440 , n206202 );
nor ( n206204 , n28439 , n28442 );
buf ( n28444 , RI19a90188_2682);
nand ( n28445 , n25451 , n28444 );
buf ( n28446 , RI17465f40_1239);
and ( n28447 , n28445 , n28446 );
not ( n28448 , n28445 );
not ( n28449 , RI17465f40_1239);
and ( n28450 , n28448 , n28449 );
nor ( n28451 , n28447 , n28450 );
xor ( n28452 , n206204 , n28451 );
buf ( n28453 , RI19ac0860_2327);
nand ( n28454 , n25540 , n28453 );
not ( n206216 , RI174aec18_884);
and ( n28456 , n28454 , n206216 );
not ( n28457 , n28454 );
buf ( n28458 , RI174aec18_884);
and ( n28459 , n28457 , n28458 );
nor ( n28460 , n28456 , n28459 );
xnor ( n28461 , n28452 , n28460 );
not ( n28462 , n28461 );
buf ( n28463 , n28462 );
not ( n28464 , n28463 );
or ( n28465 , n28428 , n28464 );
buf ( n28466 , n28461 );
not ( n28467 , RI1744fce0_1347);
nand ( n28468 , n28466 , n28467 );
nand ( n28469 , n28465 , n28468 );
buf ( n28470 , RI173e7190_1629);
not ( n206232 , n28470 );
not ( n28472 , RI1739e158_1985);
not ( n206234 , n28472 );
or ( n28474 , n206232 , n206234 );
not ( n28475 , RI173e7190_1629);
buf ( n28476 , RI1739e158_1985);
nand ( n28477 , n28475 , n28476 );
nand ( n28478 , n28474 , n28477 );
not ( n28479 , RI1745ec68_1274);
and ( n28480 , n28478 , n28479 );
not ( n28481 , n28478 );
buf ( n28482 , RI1745ec68_1274);
and ( n28483 , n28481 , n28482 );
nor ( n28484 , n28480 , n28483 );
buf ( n206246 , RI19aa3c88_2539);
nand ( n28486 , n26058 , n206246 );
buf ( n28487 , RI17483478_1096);
and ( n28488 , n28486 , n28487 );
not ( n28489 , n28486 );
not ( n28490 , RI17483478_1096);
and ( n28491 , n28489 , n28490 );
nor ( n28492 , n28488 , n28491 );
xor ( n28493 , n28484 , n28492 );
buf ( n28494 , RI19a85058_2759);
nand ( n28495 , n26325 , n28494 );
not ( n206257 , RI17508078_741);
and ( n28497 , n28495 , n206257 );
not ( n206259 , n28495 );
buf ( n28499 , RI17508078_741);
and ( n28500 , n206259 , n28499 );
nor ( n28501 , n28497 , n28500 );
xnor ( n28502 , n28493 , n28501 );
buf ( n28503 , n28502 );
and ( n28504 , n28469 , n28503 );
not ( n28505 , n28469 );
not ( n28506 , n28484 );
xor ( n28507 , n28506 , n28492 );
xnor ( n28508 , n28507 , n28501 );
not ( n28509 , n28508 );
not ( n206271 , n28509 );
buf ( n28511 , n206271 );
and ( n206273 , n28505 , n28511 );
nor ( n28513 , n28504 , n206273 );
and ( n28514 , n28426 , n28513 );
not ( n28515 , n28426 );
not ( n28516 , n28513 );
and ( n28517 , n28515 , n28516 );
nor ( n28518 , n28514 , n28517 );
xor ( n28519 , n206058 , n28518 );
not ( n28520 , n28127 );
nand ( n28521 , n28520 , n28051 );
buf ( n28522 , RI173cc6e8_1759);
not ( n28523 , n28522 );
not ( n28524 , RI17343168_2114);
not ( n206286 , n28524 );
or ( n28526 , n28523 , n206286 );
not ( n28527 , RI173cc6e8_1759);
buf ( n28528 , RI17343168_2114);
nand ( n28529 , n28527 , n28528 );
nand ( n28530 , n28526 , n28529 );
buf ( n28531 , RI17415720_1403);
and ( n28532 , n28530 , n28531 );
not ( n28533 , n28530 );
not ( n28534 , RI17415720_1403);
and ( n28535 , n28533 , n28534 );
nor ( n206297 , n28532 , n28535 );
buf ( n28537 , RI19a8d410_2702);
nand ( n28538 , n204336 , n28537 );
buf ( n28539 , RI17468d30_1225);
and ( n28540 , n28538 , n28539 );
not ( n28541 , n28538 );
not ( n28542 , RI17468d30_1225);
and ( n28543 , n28541 , n28542 );
nor ( n28544 , n28540 , n28543 );
not ( n28545 , n28544 );
xor ( n206307 , n206297 , n28545 );
buf ( n28547 , RI19abe4c0_2347);
nand ( n206309 , n25916 , n28547 );
not ( n28549 , RI174b1a08_870);
and ( n206311 , n206309 , n28549 );
not ( n28551 , n206309 );
buf ( n28552 , RI174b1a08_870);
and ( n28553 , n28551 , n28552 );
nor ( n28554 , n206311 , n28553 );
xnor ( n28555 , n206307 , n28554 );
not ( n28556 , n28555 );
not ( n28557 , n28556 );
not ( n28558 , n28557 );
buf ( n28559 , RI1740fb40_1431);
not ( n206321 , n28559 );
buf ( n28561 , RI173f7ea0_1547);
not ( n206323 , n28561 );
not ( n28563 , RI173af1b0_1902);
not ( n28564 , n28563 );
or ( n28565 , n206323 , n28564 );
not ( n28566 , RI173f7ea0_1547);
buf ( n28567 , RI173af1b0_1902);
nand ( n28568 , n28566 , n28567 );
nand ( n28569 , n28565 , n28568 );
not ( n28570 , RI1733d8d0_2141);
and ( n28571 , n28569 , n28570 );
not ( n28572 , n28569 );
buf ( n28573 , RI1733d8d0_2141);
and ( n206335 , n28572 , n28573 );
nor ( n28575 , n28571 , n206335 );
buf ( n206337 , RI19aa5a88_2525);
nand ( n28577 , n204512 , n206337 );
buf ( n28578 , RI17522c70_658);
and ( n28579 , n28577 , n28578 );
not ( n28580 , n28577 );
not ( n28581 , RI17522c70_658);
and ( n28582 , n28580 , n28581 );
nor ( n28583 , n28579 , n28582 );
xor ( n28584 , n28575 , n28583 );
buf ( n28585 , RI19aaac18_2490);
nand ( n206347 , n204926 , n28585 );
buf ( n28587 , RI174944d0_1013);
and ( n206349 , n206347 , n28587 );
not ( n28589 , n206347 );
not ( n28590 , RI174944d0_1013);
and ( n28591 , n28589 , n28590 );
nor ( n28592 , n206349 , n28591 );
xnor ( n28593 , n28584 , n28592 );
not ( n28594 , n28593 );
not ( n28595 , n28594 );
or ( n28596 , n206321 , n28595 );
not ( n28597 , n28594 );
not ( n28598 , RI1740fb40_1431);
nand ( n28599 , n28597 , n28598 );
nand ( n28600 , n28596 , n28599 );
not ( n28601 , n28600 );
or ( n28602 , n28558 , n28601 );
buf ( n28603 , n28555 );
or ( n28604 , n28600 , n28603 );
nand ( n28605 , n28602 , n28604 );
and ( n28606 , n28521 , n28605 );
not ( n28607 , n28521 );
not ( n206369 , n28605 );
and ( n28609 , n28607 , n206369 );
or ( n206371 , n28606 , n28609 );
xnor ( n28611 , n28519 , n206371 );
buf ( n28612 , RI17444ef8_1400);
buf ( n28613 , RI173dc060_1683);
not ( n28614 , n28613 );
not ( n28615 , RI17393370_2038);
not ( n28616 , n28615 );
or ( n28617 , n28614 , n28616 );
not ( n28618 , RI173dc060_1683);
buf ( n28619 , RI17393370_2038);
nand ( n206381 , n28618 , n28619 );
nand ( n28621 , n28617 , n206381 );
buf ( n28622 , RI17453b38_1328);
and ( n28623 , n28621 , n28622 );
not ( n28624 , n28621 );
not ( n28625 , RI17453b38_1328);
and ( n28626 , n28624 , n28625 );
nor ( n28627 , n28623 , n28626 );
buf ( n28628 , RI19ac7b38_2272);
nand ( n28629 , n26453 , n28628 );
buf ( n28630 , RI174c62a0_794);
and ( n28631 , n28629 , n28630 );
not ( n28632 , n28629 );
not ( n28633 , RI174c62a0_794);
and ( n28634 , n28632 , n28633 );
nor ( n28635 , n28631 , n28634 );
xor ( n206397 , n28627 , n28635 );
buf ( n28637 , n26242 );
buf ( n206399 , RI19a97dc0_2627);
nand ( n28639 , n28637 , n206399 );
buf ( n206401 , RI17478690_1149);
and ( n28641 , n28639 , n206401 );
not ( n28642 , n28639 );
not ( n28643 , RI17478690_1149);
and ( n28644 , n28642 , n28643 );
nor ( n28645 , n28641 , n28644 );
xnor ( n28646 , n206397 , n28645 );
buf ( n28647 , n28646 );
xor ( n28648 , n28612 , n28647 );
not ( n28649 , RI17447ce8_1386);
not ( n206411 , RI17407800_1471);
buf ( n28651 , RI173beb10_1826);
and ( n206413 , n206411 , n28651 );
not ( n28653 , n206411 );
not ( n28654 , RI173beb10_1826);
and ( n28655 , n28653 , n28654 );
nor ( n28656 , n206413 , n28655 );
xor ( n28657 , n28649 , n28656 );
buf ( n28658 , RI17335590_2181);
buf ( n28659 , RI174a3ae8_938);
xor ( n28660 , n28658 , n28659 );
buf ( n28661 , RI19ab52f8_2415);
nand ( n28662 , n204926 , n28661 );
xnor ( n28663 , n28660 , n28662 );
xnor ( n206425 , n28657 , n28663 );
buf ( n28665 , n206425 );
xnor ( n206427 , n28648 , n28665 );
not ( n28667 , n206427 );
not ( n28668 , n28096 );
not ( n28669 , n28668 );
not ( n28670 , n25426 );
or ( n28671 , n28669 , n28670 );
not ( n28672 , n28668 );
nand ( n28673 , n28672 , n25429 );
nand ( n28674 , n28671 , n28673 );
xor ( n28675 , n205114 , n205132 );
xnor ( n206437 , n28675 , n205122 );
not ( n28677 , n206437 );
and ( n28678 , n28674 , n28677 );
not ( n28679 , n28674 );
buf ( n28680 , n206437 );
and ( n28681 , n28679 , n28680 );
nor ( n28682 , n28678 , n28681 );
buf ( n28683 , n204713 );
not ( n28684 , n28683 );
buf ( n28685 , RI173d8f28_1698);
not ( n28686 , n28685 );
not ( n28687 , RI17390238_2053);
not ( n28688 , n28687 );
or ( n28689 , n28686 , n28688 );
not ( n206451 , RI173d8f28_1698);
buf ( n28691 , RI17390238_2053);
nand ( n28692 , n206451 , n28691 );
nand ( n206454 , n28689 , n28692 );
not ( n28694 , RI17450a00_1343);
and ( n206456 , n206454 , n28694 );
not ( n28696 , n206454 );
buf ( n28697 , RI17450a00_1343);
and ( n28698 , n28696 , n28697 );
nor ( n28699 , n206456 , n28698 );
buf ( n28700 , RI19a98630_2623);
nand ( n28701 , n25479 , n28700 );
buf ( n28702 , RI17475210_1165);
and ( n28703 , n28701 , n28702 );
not ( n28704 , n28701 );
not ( n206466 , RI17475210_1165);
and ( n28706 , n28704 , n206466 );
nor ( n206468 , n28703 , n28706 );
xor ( n28708 , n28699 , n206468 );
buf ( n28709 , RI19ac81c8_2269);
nand ( n28710 , n27749 , n28709 );
not ( n28711 , RI174c1548_809);
and ( n28712 , n28710 , n28711 );
not ( n28713 , n28710 );
buf ( n28714 , RI174c1548_809);
and ( n28715 , n28713 , n28714 );
nor ( n28716 , n28712 , n28715 );
xnor ( n28717 , n28708 , n28716 );
not ( n206479 , n28717 );
not ( n28719 , n206479 );
or ( n206481 , n28684 , n28719 );
buf ( n28721 , n28717 );
not ( n28722 , n28721 );
or ( n28723 , n28722 , n28683 );
nand ( n28724 , n206481 , n28723 );
not ( n28725 , n26366 );
xor ( n28726 , n28724 , n28725 );
nor ( n28727 , n28682 , n28726 );
not ( n28728 , n28727 );
and ( n28729 , n28667 , n28728 );
and ( n28730 , n206427 , n28727 );
nor ( n28731 , n28729 , n28730 );
not ( n206493 , n28731 );
buf ( n28733 , RI19ab4380_2422);
nand ( n206495 , n25583 , n28733 );
not ( n28735 , RI174a5f00_927);
and ( n28736 , n206495 , n28735 );
not ( n28737 , n206495 );
buf ( n28738 , RI174a5f00_927);
and ( n28739 , n28737 , n28738 );
nor ( n28740 , n28736 , n28739 );
not ( n28741 , n28740 );
not ( n28742 , n28741 );
buf ( n28743 , RI173fac90_1533);
not ( n28744 , n28743 );
not ( n28745 , RI173b1fa0_1888);
not ( n28746 , n28745 );
or ( n28747 , n28744 , n28746 );
not ( n206509 , RI173fac90_1533);
buf ( n28749 , RI173b1fa0_1888);
nand ( n206511 , n206509 , n28749 );
nand ( n28751 , n28747 , n206511 );
buf ( n206513 , RI1739b9f8_1997);
and ( n28753 , n28751 , n206513 );
not ( n28754 , n28751 );
not ( n28755 , RI1739b9f8_1997);
and ( n28756 , n28754 , n28755 );
nor ( n28757 , n28753 , n28756 );
buf ( n28758 , RI19aa12d0_2559);
nand ( n28759 , n25793 , n28758 );
buf ( n28760 , RI175274a0_644);
and ( n28761 , n28759 , n28760 );
not ( n206523 , n28759 );
not ( n28763 , RI175274a0_644);
and ( n206525 , n206523 , n28763 );
nor ( n28765 , n28761 , n206525 );
xor ( n28766 , n28757 , n28765 );
buf ( n28767 , RI19aaa330_2494);
nand ( n28768 , n27749 , n28767 );
buf ( n28769 , RI174972c0_999);
and ( n28770 , n28768 , n28769 );
not ( n28771 , n28768 );
not ( n28772 , RI174972c0_999);
and ( n28773 , n28771 , n28772 );
nor ( n206535 , n28770 , n28773 );
buf ( n28775 , n206535 );
xor ( n206537 , n28766 , n28775 );
not ( n28777 , n206537 );
or ( n206539 , n28742 , n28777 );
not ( n28779 , n206537 );
not ( n28780 , n28779 );
or ( n28781 , n28780 , n28741 );
nand ( n28782 , n206539 , n28781 );
buf ( n28783 , RI173cf820_1744);
not ( n28784 , n28783 );
not ( n28785 , RI17345f58_2100);
not ( n28786 , n28785 );
or ( n28787 , n28784 , n28786 );
not ( n28788 , RI173cf820_1744);
buf ( n28789 , RI17345f58_2100);
nand ( n28790 , n28788 , n28789 );
nand ( n206552 , n28787 , n28790 );
not ( n28792 , RI17447310_1389);
and ( n206554 , n206552 , n28792 );
not ( n28794 , n206552 );
buf ( n28795 , RI17447310_1389);
and ( n28796 , n28794 , n28795 );
nor ( n28797 , n206554 , n28796 );
buf ( n28798 , RI19abddb8_2351);
nand ( n28799 , n26242 , n28798 );
not ( n28800 , RI174b47f8_856);
and ( n28801 , n28799 , n28800 );
not ( n28802 , n28799 );
buf ( n206564 , RI174b47f8_856);
and ( n28804 , n28802 , n206564 );
nor ( n206566 , n28801 , n28804 );
not ( n28806 , n206566 );
xor ( n28807 , n28797 , n28806 );
buf ( n28808 , RI19a8cb28_2706);
nand ( n28809 , n205124 , n28808 );
buf ( n28810 , RI1746bb20_1211);
and ( n28811 , n28809 , n28810 );
not ( n28812 , n28809 );
not ( n28813 , RI1746bb20_1211);
and ( n28814 , n28812 , n28813 );
nor ( n28815 , n28811 , n28814 );
xnor ( n28816 , n28807 , n28815 );
buf ( n28817 , n28816 );
and ( n28818 , n28782 , n28817 );
not ( n28819 , n28782 );
not ( n206581 , n28815 );
not ( n28821 , n206566 );
or ( n28822 , n206581 , n28821 );
or ( n28823 , n28815 , n206566 );
nand ( n28824 , n28822 , n28823 );
and ( n28825 , n28824 , n28797 );
not ( n28826 , n28824 );
not ( n28827 , n28797 );
and ( n28828 , n28826 , n28827 );
nor ( n28829 , n28825 , n28828 );
buf ( n206591 , n28829 );
and ( n28831 , n28819 , n206591 );
nor ( n206593 , n28818 , n28831 );
not ( n28833 , n206593 );
buf ( n28834 , RI19abcdc8_2360);
nand ( n28835 , n25751 , n28834 );
buf ( n28836 , RI174b6580_847);
and ( n28837 , n28835 , n28836 );
not ( n28838 , n28835 );
not ( n28839 , RI174b6580_847);
and ( n28840 , n28838 , n28839 );
nor ( n28841 , n28837 , n28840 );
buf ( n28842 , n28841 );
buf ( n28843 , RI173e0200_1663);
not ( n206605 , n28843 );
not ( n28845 , RI17397510_2018);
not ( n28846 , n28845 );
or ( n28847 , n206605 , n28846 );
not ( n28848 , RI173e0200_1663);
buf ( n28849 , RI17397510_2018);
nand ( n28850 , n28848 , n28849 );
nand ( n28851 , n28847 , n28850 );
buf ( n28852 , RI17458020_1307);
and ( n28853 , n28851 , n28852 );
not ( n28854 , n28851 );
not ( n28855 , RI17458020_1307);
and ( n28856 , n28854 , n28855 );
nor ( n206618 , n28853 , n28856 );
buf ( n28858 , RI19ac3290_2305);
nand ( n206620 , n25851 , n28858 );
buf ( n28860 , RI174cc9c0_774);
and ( n28861 , n206620 , n28860 );
not ( n28862 , n206620 );
not ( n28863 , RI174cc9c0_774);
and ( n28864 , n28862 , n28863 );
nor ( n28865 , n28861 , n28864 );
xor ( n28866 , n206618 , n28865 );
buf ( n28867 , RI19a93068_2661);
nand ( n28868 , n204916 , n28867 );
buf ( n206630 , RI1747c830_1129);
and ( n28870 , n28868 , n206630 );
not ( n206632 , n28868 );
not ( n28872 , RI1747c830_1129);
and ( n28873 , n206632 , n28872 );
nor ( n28874 , n28870 , n28873 );
not ( n28875 , n28874 );
xnor ( n28876 , n28866 , n28875 );
buf ( n28877 , n28876 );
not ( n28878 , n28877 );
xor ( n28879 , n28842 , n28878 );
xnor ( n28880 , n28879 , n25683 );
not ( n28881 , n28880 );
nand ( n28882 , n28833 , n28881 );
buf ( n28883 , RI174c8be0_786);
and ( n206645 , n28883 , n204976 );
not ( n28885 , n28883 );
and ( n28886 , n28885 , n204977 );
nor ( n28887 , n206645 , n28886 );
buf ( n28888 , RI173dfeb8_1664);
buf ( n28889 , RI17401c20_1499);
not ( n28890 , n28889 );
not ( n28891 , RI173b8f30_1854);
not ( n28892 , n28891 );
or ( n28893 , n28890 , n28892 );
not ( n28894 , RI17401c20_1499);
buf ( n206656 , RI173b8f30_1854);
nand ( n28896 , n28894 , n206656 );
nand ( n206658 , n28893 , n28896 );
xor ( n28898 , n28888 , n206658 );
buf ( n28899 , RI17531ec8_611);
buf ( n28900 , RI1749df08_966);
xor ( n28901 , n28899 , n28900 );
buf ( n28902 , n25491 );
buf ( n28903 , RI19ab8d90_2389);
nand ( n28904 , n28902 , n28903 );
xnor ( n28905 , n28901 , n28904 );
xnor ( n28906 , n28898 , n28905 );
not ( n28907 , n28906 );
not ( n206669 , n28907 );
not ( n28909 , n206669 );
and ( n206671 , n28887 , n28909 );
not ( n28911 , n28887 );
and ( n28912 , n28911 , n206669 );
nor ( n28913 , n206671 , n28912 );
not ( n28914 , n28913 );
and ( n28915 , n28882 , n28914 );
not ( n28916 , n28882 );
and ( n28917 , n28916 , n28913 );
nor ( n28918 , n28915 , n28917 );
not ( n28919 , n28918 );
or ( n206681 , n206493 , n28919 );
not ( n28921 , n28918 );
not ( n206683 , n28731 );
nand ( n28923 , n28921 , n206683 );
nand ( n28924 , n206681 , n28923 );
not ( n28925 , n28924 );
and ( n28926 , n28611 , n28925 );
not ( n28927 , n28611 );
and ( n28928 , n28927 , n28924 );
nor ( n28929 , n28926 , n28928 );
not ( n28930 , n28929 );
or ( n28931 , n205891 , n28930 );
not ( n28932 , n28129 );
and ( n28933 , n28611 , n28924 );
not ( n28934 , n28611 );
and ( n28935 , n28934 , n28925 );
nor ( n28936 , n28933 , n28935 );
nand ( n28937 , n28932 , n28936 );
nand ( n28938 , n28931 , n28937 );
not ( n28939 , n204501 );
not ( n206701 , n25926 );
or ( n28941 , n28939 , n206701 );
not ( n28942 , n204501 );
nand ( n28943 , n28942 , n25931 );
nand ( n28944 , n28941 , n28943 );
and ( n28945 , n28944 , n25965 );
not ( n28946 , n28944 );
and ( n28947 , n28946 , n25978 );
nor ( n28948 , n28945 , n28947 );
not ( n28949 , n28948 );
not ( n28950 , n28949 );
buf ( n28951 , RI17453160_1331);
buf ( n28952 , RI17408868_1466);
not ( n28953 , n28952 );
not ( n28954 , RI173bfb78_1821);
not ( n28955 , n28954 );
or ( n28956 , n28953 , n28955 );
not ( n28957 , RI17408868_1466);
buf ( n28958 , RI173bfb78_1821);
nand ( n28959 , n28957 , n28958 );
nand ( n206721 , n28956 , n28959 );
xor ( n28961 , n28951 , n206721 );
buf ( n206723 , RI173365f8_2176);
not ( n28963 , RI174a4b50_933);
xor ( n28964 , n206723 , n28963 );
buf ( n28965 , RI19ab36d8_2428);
nand ( n28966 , n205271 , n28965 );
xnor ( n28967 , n28964 , n28966 );
xnor ( n28968 , n28961 , n28967 );
not ( n28969 , n28968 );
not ( n28970 , n28969 );
buf ( n28971 , RI173f9c28_1538);
not ( n28972 , n28971 );
buf ( n28973 , RI173eb330_1609);
not ( n28974 , n28973 );
not ( n206736 , RI173a2640_1964);
not ( n28976 , n206736 );
or ( n28977 , n28974 , n28976 );
not ( n28978 , RI173eb330_1609);
buf ( n28979 , RI173a2640_1964);
nand ( n28980 , n28978 , n28979 );
nand ( n28981 , n28977 , n28980 );
buf ( n28982 , RI17475558_1164);
and ( n28983 , n28981 , n28982 );
not ( n28984 , n28981 );
not ( n28985 , RI17475558_1164);
and ( n206747 , n28984 , n28985 );
nor ( n28987 , n28983 , n206747 );
buf ( n206749 , RI19a9fae8_2571);
nand ( n28989 , n25628 , n206749 );
buf ( n28990 , RI17487618_1076);
and ( n28991 , n28989 , n28990 );
not ( n28992 , n28989 );
not ( n28993 , RI17487618_1076);
and ( n28994 , n28992 , n28993 );
nor ( n28995 , n28991 , n28994 );
xor ( n28996 , n28987 , n28995 );
buf ( n28997 , n25879 );
buf ( n28998 , RI19ace870_2221);
nand ( n28999 , n28997 , n28998 );
not ( n29000 , RI1750e798_721);
and ( n29001 , n28999 , n29000 );
not ( n206763 , n28999 );
buf ( n29003 , RI1750e798_721);
and ( n206765 , n206763 , n29003 );
nor ( n29005 , n29001 , n206765 );
xnor ( n29006 , n28996 , n29005 );
not ( n29007 , n29006 );
not ( n29008 , n29007 );
or ( n29009 , n28972 , n29008 );
not ( n29010 , RI173f9c28_1538);
nand ( n29011 , n29006 , n29010 );
nand ( n29012 , n29009 , n29011 );
not ( n29013 , n29012 );
and ( n29014 , n28970 , n29013 );
buf ( n29015 , n28968 );
not ( n206777 , n29015 );
and ( n29017 , n206777 , n29012 );
nor ( n206779 , n29014 , n29017 );
not ( n29019 , n206779 );
buf ( n29020 , RI173a7848_1939);
not ( n29021 , n29020 );
buf ( n29022 , RI17398c08_2011);
not ( n29023 , n29022 );
not ( n29024 , RI173e18f8_1656);
not ( n29025 , n29024 );
or ( n29026 , n29023 , n29025 );
not ( n29027 , RI17398c08_2011);
buf ( n206789 , RI173e18f8_1656);
nand ( n29029 , n29027 , n206789 );
nand ( n206791 , n29026 , n29029 );
not ( n29031 , RI17459718_1300);
and ( n29032 , n206791 , n29031 );
not ( n29033 , n206791 );
buf ( n29034 , RI17459718_1300);
and ( n29035 , n29033 , n29034 );
nor ( n29036 , n29032 , n29035 );
xor ( n29037 , n29036 , n28039 );
buf ( n29038 , RI19a94238_2653);
nand ( n29039 , n28997 , n29038 );
not ( n29040 , RI1747df28_1122);
and ( n29041 , n29039 , n29040 );
not ( n206803 , n29039 );
buf ( n29043 , RI1747df28_1122);
and ( n206805 , n206803 , n29043 );
nor ( n29045 , n29041 , n206805 );
xnor ( n29046 , n29037 , n29045 );
not ( n29047 , n29046 );
or ( n29048 , n29021 , n29047 );
or ( n29049 , n29046 , n29020 );
nand ( n29050 , n29048 , n29049 );
not ( n29051 , n29050 );
buf ( n29052 , RI174a9d58_908);
buf ( n29053 , RI173f0880_1583);
not ( n206815 , n29053 );
not ( n29055 , RI173a7b90_1938);
not ( n29056 , n29055 );
or ( n29057 , n206815 , n29056 );
not ( n29058 , RI173f0880_1583);
buf ( n29059 , RI173a7b90_1938);
nand ( n29060 , n29058 , n29059 );
nand ( n29061 , n29057 , n29060 );
xor ( n29062 , n29052 , n29061 );
buf ( n29063 , RI19aafad8_2456);
nand ( n29064 , n25741 , n29063 );
not ( n29065 , n29064 );
buf ( n29066 , RI1748cb68_1050);
not ( n29067 , n29066 );
and ( n29068 , n29065 , n29067 );
nand ( n29069 , n25656 , n29063 );
and ( n29070 , n29069 , n29066 );
nor ( n206832 , n29068 , n29070 );
not ( n29072 , n206832 );
buf ( n29073 , RI19a85508_2757);
nand ( n29074 , n25751 , n29073 );
not ( n29075 , RI175172d0_694);
and ( n29076 , n29074 , n29075 );
not ( n29077 , n29074 );
buf ( n29078 , RI175172d0_694);
and ( n29079 , n29077 , n29078 );
nor ( n29080 , n29076 , n29079 );
not ( n29081 , n29080 );
or ( n29082 , n29072 , n29081 );
not ( n29083 , n29080 );
not ( n29084 , n206832 );
nand ( n206846 , n29083 , n29084 );
nand ( n29086 , n29082 , n206846 );
xnor ( n206848 , n29062 , n29086 );
buf ( n29088 , n206848 );
not ( n29089 , n29088 );
or ( n29090 , n29051 , n29089 );
or ( n29091 , n29088 , n29050 );
nand ( n29092 , n29090 , n29091 );
not ( n29093 , n29092 );
nand ( n29094 , n29019 , n29093 );
not ( n29095 , n29094 );
or ( n206857 , n28950 , n29095 );
or ( n29097 , n29094 , n28949 );
nand ( n206859 , n206857 , n29097 );
not ( n29099 , n206859 );
buf ( n29100 , RI17340a08_2126);
not ( n29101 , n29100 );
not ( n29102 , RI173f8f08_1542);
not ( n29103 , RI17404380_1487);
buf ( n29104 , RI173bb690_1842);
nand ( n29105 , n29103 , n29104 );
not ( n29106 , RI173bb690_1842);
buf ( n29107 , RI17404380_1487);
nand ( n29108 , n29106 , n29107 );
and ( n29109 , n29105 , n29108 );
xor ( n29110 , n29102 , n29109 );
buf ( n29111 , RI17535ca8_599);
buf ( n29112 , RI174a0668_954);
xor ( n29113 , n29111 , n29112 );
buf ( n206875 , RI19ab7f80_2395);
nand ( n29115 , n28637 , n206875 );
xnor ( n206877 , n29113 , n29115 );
xnor ( n29117 , n29110 , n206877 );
not ( n29118 , n29117 );
or ( n29119 , n29101 , n29118 );
not ( n29120 , n29100 );
buf ( n29121 , RI173f8f08_1542);
xor ( n29122 , n29121 , n29109 );
xnor ( n29123 , n29122 , n206877 );
nand ( n29124 , n29120 , n29123 );
nand ( n29125 , n29119 , n29124 );
buf ( n206887 , RI173d8be0_1699);
not ( n29127 , n206887 );
not ( n29128 , RI1738fef0_2054);
not ( n29129 , n29128 );
or ( n29130 , n29127 , n29129 );
not ( n29131 , RI173d8be0_1699);
buf ( n29132 , RI1738fef0_2054);
nand ( n29133 , n29131 , n29132 );
nand ( n29134 , n29130 , n29133 );
buf ( n29135 , RI174506b8_1344);
and ( n29136 , n29134 , n29135 );
not ( n29137 , n29134 );
not ( n29138 , RI174506b8_1344);
and ( n206900 , n29137 , n29138 );
nor ( n29140 , n29136 , n206900 );
buf ( n206902 , n25415 );
buf ( n29142 , RI19a983d8_2624);
nand ( n29143 , n206902 , n29142 );
buf ( n29144 , RI17474ec8_1166);
and ( n29145 , n29143 , n29144 );
not ( n29146 , n29143 );
not ( n29147 , RI17474ec8_1166);
and ( n29148 , n29146 , n29147 );
nor ( n29149 , n29145 , n29148 );
xor ( n29150 , n29140 , n29149 );
buf ( n29151 , n25571 );
buf ( n29152 , RI19ac7f70_2270);
nand ( n206914 , n29151 , n29152 );
not ( n29154 , RI174c1020_810);
and ( n29155 , n206914 , n29154 );
not ( n29156 , n206914 );
buf ( n29157 , RI174c1020_810);
and ( n29158 , n29156 , n29157 );
nor ( n29159 , n29155 , n29158 );
buf ( n29160 , n29159 );
xnor ( n29161 , n29150 , n29160 );
buf ( n29162 , n29161 );
and ( n29163 , n29125 , n29162 );
not ( n29164 , n29125 );
not ( n29165 , n29149 );
not ( n29166 , n29159 );
or ( n206928 , n29165 , n29166 );
or ( n29168 , n29149 , n29159 );
nand ( n206930 , n206928 , n29168 );
not ( n29170 , n29140 );
and ( n29171 , n206930 , n29170 );
not ( n29172 , n206930 );
and ( n29173 , n29172 , n29140 );
nor ( n29174 , n29171 , n29173 );
buf ( n29175 , n29174 );
and ( n29176 , n29164 , n29175 );
nor ( n29177 , n29163 , n29176 );
not ( n29178 , n29177 );
buf ( n206940 , RI173e2618_1652);
not ( n29180 , n206940 );
not ( n206942 , RI17399928_2007);
not ( n29182 , n206942 );
or ( n29183 , n29180 , n29182 );
not ( n29184 , RI173e2618_1652);
buf ( n29185 , RI17399928_2007);
nand ( n29186 , n29184 , n29185 );
nand ( n29187 , n29183 , n29186 );
buf ( n29188 , RI1745a438_1296);
and ( n29189 , n29187 , n29188 );
not ( n206951 , n29187 );
not ( n29191 , RI1745a438_1296);
and ( n206953 , n206951 , n29191 );
nor ( n29193 , n29189 , n206953 );
buf ( n29194 , RI19a86fc0_2745);
nand ( n29195 , n25451 , n29194 );
buf ( n29196 , RI174d0278_763);
and ( n29197 , n29195 , n29196 );
not ( n29198 , n29195 );
not ( n29199 , RI174d0278_763);
and ( n29200 , n29198 , n29199 );
nor ( n29201 , n29197 , n29200 );
xor ( n206963 , n29193 , n29201 );
buf ( n29203 , n26453 );
buf ( n206965 , RI19aa5dd0_2524);
nand ( n29205 , n29203 , n206965 );
not ( n29206 , RI1747ec48_1118);
and ( n29207 , n29205 , n29206 );
not ( n29208 , n29205 );
buf ( n29209 , RI1747ec48_1118);
and ( n29210 , n29208 , n29209 );
nor ( n29211 , n29207 , n29210 );
xnor ( n29212 , n206963 , n29211 );
not ( n29213 , n29212 );
not ( n29214 , n29213 );
not ( n206976 , n29214 );
not ( n29216 , n206976 );
buf ( n206978 , RI173d39d8_1724);
not ( n29218 , n206978 );
buf ( n29219 , RI173c50c8_1795);
not ( n29220 , n29219 );
not ( n29221 , RI1733bb48_2150);
not ( n29222 , n29221 );
or ( n29223 , n29220 , n29222 );
not ( n29224 , RI173c50c8_1795);
buf ( n29225 , RI1733bb48_2150);
nand ( n29226 , n29224 , n29225 );
nand ( n206988 , n29223 , n29226 );
buf ( n29228 , RI1740ddb8_1440);
and ( n29229 , n206988 , n29228 );
not ( n29230 , n206988 );
not ( n29231 , RI1740ddb8_1440);
and ( n29232 , n29230 , n29231 );
nor ( n29233 , n29229 , n29232 );
buf ( n29234 , RI19ac2390_2312);
nand ( n29235 , n204493 , n29234 );
buf ( n29236 , RI174aa3e8_906);
and ( n29237 , n29235 , n29236 );
not ( n29238 , n29235 );
not ( n29239 , RI174aa3e8_906);
and ( n29240 , n29238 , n29239 );
nor ( n207002 , n29237 , n29240 );
xor ( n29242 , n29233 , n207002 );
buf ( n29243 , RI19a920f0_2668);
nand ( n29244 , n25741 , n29243 );
buf ( n29245 , RI17461710_1261);
and ( n29246 , n29244 , n29245 );
not ( n29247 , n29244 );
not ( n29248 , RI17461710_1261);
and ( n29249 , n29247 , n29248 );
nor ( n29250 , n29246 , n29249 );
xnor ( n207012 , n29242 , n29250 );
not ( n29252 , n207012 );
or ( n29253 , n29218 , n29252 );
or ( n29254 , n207012 , n206978 );
nand ( n29255 , n29253 , n29254 );
not ( n29256 , n29255 );
or ( n29257 , n29216 , n29256 );
not ( n29258 , n29214 );
or ( n29259 , n29255 , n29258 );
nand ( n29260 , n29257 , n29259 );
nand ( n29261 , n29178 , n29260 );
not ( n207023 , n29261 );
buf ( n29263 , RI17335f68_2178);
not ( n207025 , n29263 );
buf ( n29265 , RI173b0bf0_1894);
not ( n29266 , n29265 );
not ( n29267 , RI173f98e0_1539);
not ( n29268 , n29267 );
or ( n29269 , n29266 , n29268 );
not ( n29270 , RI173b0bf0_1894);
buf ( n29271 , RI173f98e0_1539);
nand ( n29272 , n29270 , n29271 );
nand ( n29273 , n29269 , n29272 );
not ( n29274 , RI1738e168_2063);
and ( n29275 , n29273 , n29274 );
not ( n29276 , n29273 );
buf ( n29277 , RI1738e168_2063);
and ( n29278 , n29276 , n29277 );
nor ( n207040 , n29275 , n29278 );
not ( n29280 , n207040 );
buf ( n29281 , RI19a981f8_2625);
nand ( n207043 , n25751 , n29281 );
buf ( n29283 , RI175255b0_650);
and ( n207045 , n207043 , n29283 );
not ( n29285 , n207043 );
not ( n29286 , RI175255b0_650);
and ( n29287 , n29285 , n29286 );
nor ( n29288 , n207045 , n29287 );
xor ( n29289 , n29280 , n29288 );
buf ( n29290 , RI19aa9688_2500);
nand ( n29291 , n204426 , n29290 );
buf ( n29292 , RI17495f10_1005);
and ( n29293 , n29291 , n29292 );
not ( n29294 , n29291 );
not ( n29295 , RI17495f10_1005);
and ( n29296 , n29294 , n29295 );
nor ( n29297 , n29293 , n29296 );
xnor ( n207059 , n29289 , n29297 );
not ( n29299 , n207059 );
or ( n29300 , n207025 , n29299 );
or ( n29301 , n207059 , n29263 );
nand ( n29302 , n29300 , n29301 );
not ( n29303 , n205423 );
not ( n29304 , RI17344ba8_2106);
not ( n29305 , n29304 );
or ( n29306 , n29303 , n29305 );
not ( n29307 , RI173ce470_1750);
buf ( n29308 , RI17344ba8_2106);
nand ( n29309 , n29307 , n29308 );
nand ( n29310 , n29306 , n29309 );
not ( n207072 , RI17445f60_1395);
and ( n29312 , n29310 , n207072 );
not ( n207074 , n29310 );
buf ( n29314 , RI17445f60_1395);
and ( n29315 , n207074 , n29314 );
nor ( n29316 , n29312 , n29315 );
buf ( n29317 , RI19abd2f0_2357);
nand ( n29318 , n204512 , n29317 );
buf ( n29319 , RI174b3448_862);
and ( n29320 , n29318 , n29319 );
not ( n29321 , n29318 );
not ( n29322 , RI174b3448_862);
and ( n207084 , n29321 , n29322 );
nor ( n29324 , n29320 , n207084 );
xor ( n207086 , n29316 , n29324 );
buf ( n29326 , RI19a8be08_2712);
nand ( n29327 , n26325 , n29326 );
buf ( n29328 , RI1746a770_1217);
and ( n29329 , n29327 , n29328 );
not ( n29330 , n29327 );
not ( n29331 , RI1746a770_1217);
and ( n29332 , n29330 , n29331 );
nor ( n29333 , n29329 , n29332 );
xor ( n29334 , n207086 , n29333 );
not ( n29335 , n29334 );
not ( n29336 , n29335 );
and ( n207098 , n29302 , n29336 );
not ( n29338 , n29302 );
not ( n207100 , n29336 );
and ( n29340 , n29338 , n207100 );
nor ( n29341 , n207098 , n29340 );
not ( n29342 , n29341 );
not ( n29343 , n29342 );
and ( n29344 , n207023 , n29343 );
and ( n29345 , n29261 , n29342 );
nor ( n29346 , n29344 , n29345 );
not ( n29347 , n29346 );
or ( n29348 , n29099 , n29347 );
or ( n29349 , n29346 , n206859 );
nand ( n29350 , n29348 , n29349 );
buf ( n29351 , RI173d2cb8_1728);
buf ( n29352 , n27961 );
xor ( n207114 , n29351 , n29352 );
buf ( n29354 , RI17411f58_1420);
buf ( n207116 , RI173c4060_1800);
not ( n29356 , n207116 );
not ( n207118 , RI1740cd50_1445);
not ( n29358 , n207118 );
or ( n29359 , n29356 , n29358 );
not ( n29360 , RI173c4060_1800);
buf ( n29361 , RI1740cd50_1445);
nand ( n29362 , n29360 , n29361 );
nand ( n29363 , n29359 , n29362 );
xor ( n29364 , n29354 , n29363 );
buf ( n29365 , RI1733aae0_2155);
buf ( n29366 , RI174a9380_911);
xor ( n207128 , n29365 , n29366 );
buf ( n29368 , RI19ab1860_2442);
nand ( n29369 , n25666 , n29368 );
xnor ( n29370 , n207128 , n29369 );
xnor ( n29371 , n29364 , n29370 );
buf ( n29372 , n29371 );
xnor ( n29373 , n207114 , n29372 );
not ( n29374 , n29373 );
buf ( n29375 , RI173c39d0_1802);
not ( n29376 , n29375 );
buf ( n29377 , RI173fe110_1517);
not ( n207139 , n29377 );
not ( n29379 , RI173b50d8_1873);
not ( n207141 , n29379 );
or ( n29381 , n207139 , n207141 );
not ( n29382 , RI173fe110_1517);
buf ( n29383 , RI173b50d8_1873);
nand ( n29384 , n29382 , n29383 );
nand ( n29385 , n29381 , n29384 );
buf ( n29386 , RI173b95c0_1852);
and ( n29387 , n29385 , n29386 );
not ( n29388 , n29385 );
not ( n29389 , RI173b95c0_1852);
and ( n207151 , n29388 , n29389 );
nor ( n29391 , n29387 , n207151 );
buf ( n207153 , RI19a88460_2736);
nand ( n29393 , n25572 , n207153 );
buf ( n29394 , RI1752c1f8_629);
and ( n29395 , n29393 , n29394 );
not ( n29396 , n29393 );
not ( n29397 , RI1752c1f8_629);
and ( n29398 , n29396 , n29397 );
nor ( n29399 , n29395 , n29398 );
xor ( n29400 , n29391 , n29399 );
buf ( n29401 , RI19aa71f8_2515);
nand ( n29402 , n25583 , n29401 );
buf ( n207164 , RI1749a3f8_984);
and ( n29404 , n29402 , n207164 );
not ( n29405 , n29402 );
not ( n29406 , RI1749a3f8_984);
and ( n29407 , n29405 , n29406 );
nor ( n29408 , n29404 , n29407 );
xnor ( n29409 , n29400 , n29408 );
not ( n29410 , n29409 );
buf ( n29411 , n29410 );
not ( n207173 , n29411 );
not ( n29413 , n207173 );
or ( n207175 , n29376 , n29413 );
not ( n29415 , n29410 );
not ( n29416 , n29415 );
not ( n29417 , RI173c39d0_1802);
nand ( n29418 , n29416 , n29417 );
nand ( n29419 , n207175 , n29418 );
buf ( n29420 , RI173d2970_1729);
not ( n29421 , n29420 );
not ( n29422 , RI17389c80_2084);
not ( n29423 , n29422 );
or ( n29424 , n29421 , n29423 );
not ( n29425 , RI173d2970_1729);
buf ( n29426 , RI17389c80_2084);
nand ( n29427 , n29425 , n29426 );
nand ( n29428 , n29424 , n29427 );
buf ( n207190 , RI1744a448_1374);
and ( n29430 , n29428 , n207190 );
not ( n207192 , n29428 );
not ( n29432 , RI1744a448_1374);
and ( n29433 , n207192 , n29432 );
nor ( n29434 , n29430 , n29433 );
buf ( n29435 , n25490 );
buf ( n29436 , RI19a89888_2727);
nand ( n29437 , n29435 , n29436 );
not ( n29438 , RI1746ec58_1196);
and ( n29439 , n29437 , n29438 );
not ( n29440 , n29437 );
buf ( n207202 , RI1746ec58_1196);
and ( n29442 , n29440 , n207202 );
nor ( n29443 , n29439 , n29442 );
xor ( n29444 , n29434 , n29443 );
buf ( n29445 , RI19abb5e0_2372);
nand ( n29446 , n26059 , n29445 );
not ( n29447 , RI174b7930_841);
and ( n29448 , n29446 , n29447 );
not ( n29449 , n29446 );
buf ( n29450 , RI174b7930_841);
and ( n29451 , n29449 , n29450 );
nor ( n29452 , n29448 , n29451 );
xnor ( n207214 , n29444 , n29452 );
buf ( n29454 , n207214 );
buf ( n207216 , n29454 );
not ( n29456 , n207216 );
not ( n29457 , n29456 );
and ( n29458 , n29419 , n29457 );
not ( n29459 , n29419 );
not ( n29460 , n207216 );
and ( n29461 , n29459 , n29460 );
nor ( n29462 , n29458 , n29461 );
nand ( n29463 , n29374 , n29462 );
buf ( n29464 , RI19a23858_2792);
nand ( n207226 , n25751 , n29464 );
buf ( n29466 , RI1751b0b0_682);
xor ( n207228 , n207226 , n29466 );
buf ( n29468 , n207228 );
nor ( n29469 , n204976 , n29468 );
not ( n29470 , n29469 );
nand ( n29471 , n29468 , n204976 );
nand ( n29472 , n29470 , n29471 );
xnor ( n29473 , n29472 , n206669 );
not ( n29474 , n29473 );
and ( n29475 , n29463 , n29474 );
not ( n29476 , n29463 );
and ( n29477 , n29476 , n29473 );
nor ( n29478 , n29475 , n29477 );
and ( n29479 , n29350 , n29478 );
not ( n29480 , n29350 );
not ( n207242 , n29478 );
and ( n29482 , n29480 , n207242 );
nor ( n207244 , n29479 , n29482 );
buf ( n29484 , RI173915e8_2047);
not ( n29485 , n29484 );
buf ( n29486 , RI173cb9c8_1763);
not ( n29487 , n29486 );
not ( n29488 , RI17342448_2118);
not ( n29489 , n29488 );
or ( n29490 , n29487 , n29489 );
not ( n29491 , RI173cb9c8_1763);
buf ( n29492 , RI17342448_2118);
nand ( n207254 , n29491 , n29492 );
nand ( n29494 , n29490 , n207254 );
not ( n207256 , RI17414a00_1407);
and ( n29496 , n29494 , n207256 );
not ( n29497 , n29494 );
buf ( n29498 , RI17414a00_1407);
and ( n29499 , n29497 , n29498 );
nor ( n29500 , n29496 , n29499 );
buf ( n29501 , RI19a8f210_2689);
nand ( n29502 , n27946 , n29501 );
buf ( n29503 , RI17468010_1229);
and ( n29504 , n29502 , n29503 );
not ( n29505 , n29502 );
not ( n29506 , RI17468010_1229);
and ( n29507 , n29505 , n29506 );
nor ( n29508 , n29504 , n29507 );
xor ( n29509 , n29500 , n29508 );
buf ( n207271 , RI19abfc30_2334);
nand ( n29511 , n205020 , n207271 );
not ( n207273 , RI174b0ce8_874);
and ( n29513 , n29511 , n207273 );
not ( n29514 , n29511 );
buf ( n29515 , RI174b0ce8_874);
and ( n29516 , n29514 , n29515 );
nor ( n29517 , n29513 , n29516 );
xnor ( n29518 , n29509 , n29517 );
buf ( n29519 , n29518 );
not ( n29520 , n29519 );
or ( n29521 , n29485 , n29520 );
not ( n29522 , n29508 );
xor ( n29523 , n29500 , n29522 );
xnor ( n207285 , n29523 , n29517 );
buf ( n29525 , n207285 );
not ( n29526 , RI173915e8_2047);
nand ( n29527 , n29525 , n29526 );
nand ( n29528 , n29521 , n29527 );
buf ( n29529 , RI173e8f18_1620);
not ( n29530 , n29529 );
not ( n29531 , RI1739fee0_1976);
not ( n29532 , n29531 );
or ( n29533 , n29530 , n29532 );
not ( n29534 , RI173e8f18_1620);
buf ( n207296 , RI1739fee0_1976);
nand ( n29536 , n29534 , n207296 );
nand ( n207298 , n29533 , n29536 );
buf ( n29538 , RI174609f0_1265);
and ( n29539 , n207298 , n29538 );
not ( n29540 , n207298 );
not ( n29541 , RI174609f0_1265);
and ( n29542 , n29540 , n29541 );
nor ( n29543 , n29539 , n29542 );
buf ( n29544 , RI19aa2e78_2546);
nand ( n29545 , n26276 , n29544 );
buf ( n29546 , RI17485200_1087);
and ( n29547 , n29545 , n29546 );
not ( n29548 , n29545 );
not ( n29549 , RI17485200_1087);
and ( n29550 , n29548 , n29549 );
nor ( n29551 , n29547 , n29550 );
xor ( n207313 , n29543 , n29551 );
buf ( n29553 , RI19a83f78_2766);
nand ( n207315 , n25803 , n29553 );
not ( n29555 , RI1750aee0_732);
and ( n29556 , n207315 , n29555 );
not ( n29557 , n207315 );
buf ( n29558 , RI1750aee0_732);
and ( n29559 , n29557 , n29558 );
nor ( n29560 , n29556 , n29559 );
xnor ( n29561 , n207313 , n29560 );
buf ( n29562 , n29561 );
not ( n29563 , n29562 );
not ( n207325 , n29563 );
and ( n29565 , n29528 , n207325 );
not ( n207327 , n29528 );
buf ( n29567 , n29563 );
and ( n29568 , n207327 , n29567 );
nor ( n29569 , n29565 , n29568 );
not ( n29570 , n29569 );
buf ( n29571 , RI173e9f80_1615);
not ( n29572 , n29571 );
buf ( n29573 , RI173db340_1687);
not ( n29574 , n29573 );
not ( n29575 , RI17392650_2042);
not ( n29576 , n29575 );
or ( n207338 , n29574 , n29576 );
not ( n29578 , RI173db340_1687);
buf ( n207340 , RI17392650_2042);
nand ( n29580 , n29578 , n207340 );
nand ( n29581 , n207338 , n29580 );
buf ( n29582 , RI17452e18_1332);
and ( n29583 , n29581 , n29582 );
not ( n29584 , n29581 );
not ( n29585 , RI17452e18_1332);
and ( n29586 , n29584 , n29585 );
nor ( n29587 , n29583 , n29586 );
buf ( n29588 , RI19ac74a8_2275);
nand ( n29589 , n204916 , n29588 );
buf ( n29590 , RI174c4e00_798);
and ( n29591 , n29589 , n29590 );
not ( n29592 , n29589 );
not ( n29593 , RI174c4e00_798);
and ( n207355 , n29592 , n29593 );
nor ( n29595 , n29591 , n207355 );
xor ( n29596 , n29587 , n29595 );
buf ( n29597 , n28148 );
buf ( n29598 , RI19a976b8_2630);
nand ( n29599 , n29597 , n29598 );
buf ( n29600 , RI17477628_1154);
and ( n29601 , n29599 , n29600 );
not ( n29602 , n29599 );
not ( n29603 , RI17477628_1154);
and ( n29604 , n29602 , n29603 );
nor ( n29605 , n29601 , n29604 );
xnor ( n29606 , n29596 , n29605 );
buf ( n29607 , n29606 );
buf ( n29608 , n29607 );
not ( n29609 , n29608 );
or ( n29610 , n29572 , n29609 );
or ( n29611 , n29608 , n29571 );
nand ( n29612 , n29610 , n29611 );
buf ( n29613 , RI173f8878_1544);
not ( n29614 , n29613 );
not ( n207376 , RI173afb88_1899);
not ( n207377 , n207376 );
or ( n29617 , n29614 , n207377 );
not ( n29618 , RI173f8878_1544);
buf ( n207380 , RI173afb88_1899);
nand ( n29620 , n29618 , n207380 );
nand ( n207382 , n29617 , n29620 );
buf ( n29622 , RI17344518_2108);
and ( n29623 , n207382 , n29622 );
not ( n29624 , n207382 );
not ( n29625 , RI17344518_2108);
and ( n29626 , n29624 , n29625 );
nor ( n29627 , n29623 , n29626 );
buf ( n29628 , RI19aaa858_2492);
nand ( n29629 , n205019 , n29628 );
buf ( n29630 , RI17523be8_655);
and ( n207392 , n29629 , n29630 );
not ( n29632 , n29629 );
not ( n207394 , RI17523be8_655);
and ( n29634 , n29632 , n207394 );
nor ( n29635 , n207392 , n29634 );
xor ( n29636 , n29627 , n29635 );
buf ( n29637 , RI19aab410_2487);
nand ( n29638 , n25628 , n29637 );
buf ( n29639 , RI17494ea8_1010);
and ( n29640 , n29638 , n29639 );
not ( n29641 , n29638 );
not ( n29642 , RI17494ea8_1010);
and ( n29643 , n29641 , n29642 );
nor ( n29644 , n29640 , n29643 );
xor ( n29645 , n29636 , n29644 );
not ( n207407 , n29645 );
not ( n29647 , n207407 );
not ( n207409 , n29647 );
and ( n29649 , n29612 , n207409 );
not ( n29650 , n29612 );
and ( n29651 , n29650 , n29647 );
nor ( n29652 , n29649 , n29651 );
not ( n29653 , n29652 );
nand ( n29654 , n29570 , n29653 );
not ( n29655 , n29654 );
buf ( n29656 , RI19abaa28_2376);
nand ( n29657 , n206902 , n29656 );
buf ( n29658 , RI174b68c8_846);
and ( n29659 , n29657 , n29658 );
not ( n29660 , n29657 );
not ( n207422 , RI174b68c8_846);
and ( n29662 , n29660 , n207422 );
nor ( n29663 , n29659 , n29662 );
buf ( n29664 , n29663 );
not ( n29665 , n29664 );
buf ( n29666 , RI173a0228_1975);
buf ( n29667 , RI1740bce8_1450);
not ( n29668 , n29667 );
not ( n207430 , RI173c2ff8_1805);
not ( n29670 , n207430 );
or ( n29671 , n29668 , n29670 );
not ( n29672 , RI1740bce8_1450);
buf ( n29673 , RI173c2ff8_1805);
nand ( n29674 , n29672 , n29673 );
nand ( n29675 , n29671 , n29674 );
xor ( n29676 , n29666 , n29675 );
not ( n29677 , RI17339a78_2160);
not ( n29678 , n29677 );
buf ( n29679 , RI19ab0e10_2447);
nand ( n29680 , n25656 , n29679 );
buf ( n29681 , RI174a8318_916);
and ( n29682 , n29680 , n29681 );
not ( n29683 , n29680 );
not ( n29684 , RI174a8318_916);
and ( n207446 , n29683 , n29684 );
nor ( n29686 , n29682 , n207446 );
not ( n207448 , n29686 );
not ( n29688 , n207448 );
or ( n29689 , n29678 , n29688 );
buf ( n29690 , RI17339a78_2160);
nand ( n29691 , n29686 , n29690 );
nand ( n29692 , n29689 , n29691 );
xor ( n29693 , n29676 , n29692 );
buf ( n29694 , n29693 );
not ( n29695 , n29694 );
or ( n29696 , n29665 , n29695 );
or ( n29697 , n29694 , n29664 );
nand ( n29698 , n29696 , n29697 );
buf ( n29699 , RI173e0548_1662);
not ( n29700 , n29699 );
not ( n29701 , RI17397858_2017);
not ( n29702 , n29701 );
or ( n207464 , n29700 , n29702 );
not ( n29704 , RI173e0548_1662);
buf ( n207466 , RI17397858_2017);
nand ( n29706 , n29704 , n207466 );
nand ( n29707 , n207464 , n29706 );
not ( n29708 , RI17458368_1306);
and ( n29709 , n29707 , n29708 );
not ( n29710 , n29707 );
buf ( n29711 , RI17458368_1306);
and ( n29712 , n29710 , n29711 );
nor ( n29713 , n29709 , n29712 );
buf ( n29714 , RI19ac34e8_2304);
nand ( n29715 , n26453 , n29714 );
buf ( n207477 , RI174ccee8_773);
and ( n29717 , n29715 , n207477 );
not ( n29718 , n29715 );
not ( n29719 , RI174ccee8_773);
and ( n29720 , n29718 , n29719 );
nor ( n29721 , n29717 , n29720 );
xor ( n29722 , n29713 , n29721 );
buf ( n29723 , RI19a932c0_2660);
nand ( n29724 , n25793 , n29723 );
buf ( n29725 , RI1747cb78_1128);
and ( n29726 , n29724 , n29725 );
not ( n29727 , n29724 );
not ( n29728 , RI1747cb78_1128);
and ( n29729 , n29727 , n29728 );
nor ( n207491 , n29726 , n29729 );
xnor ( n29731 , n29722 , n207491 );
buf ( n207493 , n29731 );
not ( n29733 , n207493 );
and ( n207495 , n29698 , n29733 );
not ( n29735 , n29698 );
and ( n29736 , n29735 , n207493 );
nor ( n29737 , n207495 , n29736 );
not ( n29738 , n29737 );
not ( n29739 , n29738 );
and ( n29740 , n29655 , n29739 );
and ( n29741 , n29654 , n29738 );
nor ( n29742 , n29740 , n29741 );
not ( n207504 , n29742 );
buf ( n29744 , RI173b1c58_1889);
buf ( n207506 , n25597 );
and ( n29746 , n29744 , n207506 );
not ( n29747 , n29744 );
not ( n29748 , n25594 );
and ( n29749 , n29747 , n29748 );
nor ( n29750 , n29746 , n29749 );
not ( n29751 , n29750 );
not ( n29752 , n29751 );
buf ( n29753 , RI174098d0_1461);
not ( n29754 , n29753 );
not ( n207516 , RI173c0be0_1816);
not ( n29756 , n207516 );
or ( n29757 , n29754 , n29756 );
not ( n207519 , RI174098d0_1461);
buf ( n29759 , RI173c0be0_1816);
nand ( n207521 , n207519 , n29759 );
nand ( n29761 , n29757 , n207521 );
buf ( n29762 , n29761 );
not ( n29763 , n29762 );
buf ( n29764 , RI17337660_2171);
not ( n29765 , RI1745c508_1286);
xor ( n29766 , n29764 , n29765 );
xnor ( n29767 , n29766 , n28740 );
not ( n29768 , n29767 );
not ( n29769 , n29768 );
or ( n29770 , n29763 , n29769 );
not ( n29771 , n29762 );
nand ( n207533 , n29771 , n29767 );
nand ( n29773 , n29770 , n207533 );
buf ( n207535 , n29773 );
not ( n29775 , n207535 );
not ( n29776 , n29775 );
or ( n29777 , n29752 , n29776 );
nand ( n29778 , n207535 , n29750 );
nand ( n29779 , n29777 , n29778 );
not ( n29780 , n29779 );
not ( n29781 , n26480 );
buf ( n29782 , RI173f6e38_1552);
not ( n29783 , n29782 );
not ( n207545 , RI173ae148_1907);
not ( n29785 , n207545 );
or ( n207547 , n29783 , n29785 );
not ( n29787 , RI173f6e38_1552);
buf ( n29788 , RI173ae148_1907);
nand ( n29789 , n29787 , n29788 );
nand ( n29790 , n207547 , n29789 );
buf ( n29791 , RI17332458_2196);
and ( n29792 , n29790 , n29791 );
not ( n29793 , n29790 );
not ( n29794 , RI17332458_2196);
and ( n29795 , n29793 , n29794 );
nor ( n29796 , n29792 , n29795 );
buf ( n29797 , RI19aaca18_2478);
nand ( n29798 , n25656 , n29797 );
not ( n207560 , RI17493468_1018);
and ( n29800 , n29798 , n207560 );
not ( n29801 , n29798 );
buf ( n29802 , RI17493468_1018);
and ( n207564 , n29801 , n29802 );
nor ( n29804 , n29800 , n207564 );
xor ( n29805 , n29796 , n29804 );
buf ( n207567 , RI19ab6cc0_2403);
nand ( n29807 , n205271 , n207567 );
not ( n29808 , RI175212a8_663);
and ( n29809 , n29807 , n29808 );
not ( n29810 , n29807 );
buf ( n29811 , RI175212a8_663);
and ( n29812 , n29810 , n29811 );
nor ( n29813 , n29809 , n29812 );
xnor ( n29814 , n29805 , n29813 );
buf ( n29815 , n29814 );
not ( n29816 , n29815 );
or ( n29817 , n29781 , n29816 );
or ( n207579 , n29815 , n26480 );
nand ( n29819 , n29817 , n207579 );
not ( n207581 , n29819 );
buf ( n29821 , RI173cb338_1765);
not ( n29822 , n29821 );
not ( n29823 , RI17341db8_2120);
not ( n29824 , n29823 );
or ( n29825 , n29822 , n29824 );
not ( n29826 , RI173cb338_1765);
buf ( n29827 , RI17341db8_2120);
nand ( n29828 , n29826 , n29827 );
nand ( n29829 , n29825 , n29828 );
buf ( n207591 , RI17414370_1409);
and ( n29831 , n29829 , n207591 );
not ( n207593 , n29829 );
not ( n29833 , RI17414370_1409);
and ( n29834 , n207593 , n29833 );
nor ( n29835 , n29831 , n29834 );
buf ( n29836 , RI19a8efb8_2690);
nand ( n29837 , n29435 , n29836 );
not ( n29838 , RI17467980_1231);
and ( n29839 , n29837 , n29838 );
not ( n29840 , n29837 );
buf ( n29841 , RI17467980_1231);
and ( n29842 , n29840 , n29841 );
nor ( n29843 , n29839 , n29842 );
xor ( n29844 , n29835 , n29843 );
buf ( n29845 , RI19abfa50_2335);
nand ( n207607 , n28902 , n29845 );
not ( n29847 , RI174b0658_876);
and ( n207609 , n207607 , n29847 );
not ( n29849 , n207607 );
buf ( n29850 , RI174b0658_876);
and ( n29851 , n29849 , n29850 );
nor ( n29852 , n207609 , n29851 );
xnor ( n29853 , n29844 , n29852 );
buf ( n29854 , n29853 );
not ( n29855 , n29854 );
not ( n29856 , n29855 );
not ( n29857 , n29856 );
and ( n29858 , n207581 , n29857 );
not ( n29859 , n29853 );
not ( n29860 , n29859 );
and ( n29861 , n29819 , n29860 );
nor ( n29862 , n29858 , n29861 );
not ( n29863 , n29862 );
nand ( n207625 , n29780 , n29863 );
buf ( n29865 , RI19a831e0_2772);
nand ( n207627 , n25850 , n29865 );
buf ( n29867 , RI17509518_737);
and ( n29868 , n207627 , n29867 );
not ( n29869 , n207627 );
not ( n29870 , RI17509518_737);
and ( n29871 , n29869 , n29870 );
nor ( n29872 , n29868 , n29871 );
not ( n29873 , n29872 );
not ( n29874 , n29873 );
buf ( n29875 , RI173d95b8_1696);
not ( n29876 , n29875 );
not ( n29877 , RI173908c8_2051);
not ( n29878 , n29877 );
or ( n29879 , n29876 , n29878 );
not ( n29880 , RI173d95b8_1696);
buf ( n29881 , RI173908c8_2051);
nand ( n29882 , n29880 , n29881 );
nand ( n29883 , n29879 , n29882 );
not ( n29884 , RI17451090_1341);
and ( n29885 , n29883 , n29884 );
not ( n29886 , n29883 );
buf ( n29887 , RI17451090_1341);
and ( n29888 , n29886 , n29887 );
nor ( n29889 , n29885 , n29888 );
buf ( n29890 , n25571 );
buf ( n29891 , RI19ac8330_2268);
nand ( n29892 , n29890 , n29891 );
buf ( n29893 , RI174c1f98_807);
and ( n29894 , n29892 , n29893 );
not ( n29895 , n29892 );
not ( n29896 , RI174c1f98_807);
and ( n29897 , n29895 , n29896 );
nor ( n29898 , n29894 , n29897 );
xor ( n29899 , n29889 , n29898 );
buf ( n29900 , RI19a98888_2622);
nand ( n207662 , n26463 , n29900 );
not ( n29902 , RI174758a0_1163);
and ( n207664 , n207662 , n29902 );
not ( n29904 , n207662 );
buf ( n29905 , RI174758a0_1163);
and ( n29906 , n29904 , n29905 );
nor ( n29907 , n207664 , n29906 );
xor ( n29908 , n29899 , n29907 );
buf ( n29909 , n29908 );
not ( n29910 , n29909 );
not ( n29911 , n29910 );
or ( n29912 , n29874 , n29911 );
not ( n29913 , n29910 );
nand ( n207675 , n29913 , n29872 );
nand ( n29915 , n29912 , n207675 );
not ( n207677 , n26436 );
buf ( n29917 , RI19ab54d8_2414);
nand ( n29918 , n25751 , n29917 );
not ( n29919 , RI17520858_665);
and ( n29920 , n29918 , n29919 );
not ( n29921 , n29918 );
buf ( n29922 , RI17520858_665);
and ( n29923 , n29921 , n29922 );
nor ( n29924 , n29920 , n29923 );
not ( n29925 , n29924 );
or ( n207687 , n207677 , n29925 );
or ( n29927 , n26436 , n29924 );
nand ( n207689 , n207687 , n29927 );
buf ( n29929 , RI173f67a8_1554);
not ( n29930 , n29929 );
not ( n29931 , RI173adab8_1909);
not ( n29932 , n29931 );
or ( n29933 , n29930 , n29932 );
not ( n29934 , RI173f67a8_1554);
buf ( n29935 , RI173adab8_1909);
nand ( n29936 , n29934 , n29935 );
nand ( n29937 , n29933 , n29936 );
not ( n29938 , RI17532918_609);
and ( n29939 , n29937 , n29938 );
not ( n29940 , n29937 );
buf ( n29941 , RI17532918_609);
and ( n29942 , n29940 , n29941 );
nor ( n207704 , n29939 , n29942 );
xor ( n29944 , n207689 , n207704 );
buf ( n207706 , n29944 );
and ( n29946 , n29915 , n207706 );
not ( n29947 , n29915 );
not ( n29948 , n207706 );
and ( n29949 , n29947 , n29948 );
nor ( n29950 , n29946 , n29949 );
buf ( n29951 , n29950 );
xor ( n29952 , n207625 , n29951 );
not ( n29953 , n29952 );
or ( n29954 , n207504 , n29953 );
or ( n207716 , n29952 , n29742 );
nand ( n29956 , n29954 , n207716 );
not ( n207718 , n29956 );
and ( n29958 , n207244 , n207718 );
not ( n29959 , n207244 );
and ( n29960 , n29959 , n29956 );
nor ( n29961 , n29958 , n29960 );
buf ( n29962 , n29961 );
and ( n29963 , n28938 , n29962 );
not ( n29964 , n28938 );
not ( n29965 , n29962 );
and ( n29966 , n29964 , n29965 );
nor ( n207728 , n29963 , n29966 );
not ( n29968 , n207728 );
buf ( n29969 , RI17411238_1424);
buf ( n29970 , n28344 );
xor ( n29971 , n29969 , n29970 );
buf ( n29972 , RI173e9260_1619);
buf ( n29973 , RI17402c88_1494);
not ( n29974 , n29973 );
not ( n29975 , RI173b9f98_1849);
not ( n29976 , n29975 );
or ( n29977 , n29974 , n29976 );
not ( n29978 , RI17402c88_1494);
buf ( n29979 , RI173b9f98_1849);
nand ( n29980 , n29978 , n29979 );
nand ( n29981 , n29977 , n29980 );
xor ( n29982 , n29972 , n29981 );
buf ( n29983 , RI17533890_606);
buf ( n29984 , RI1749ef70_961);
xor ( n29985 , n29983 , n29984 );
buf ( n207747 , RI19ab7008_2402);
nand ( n29987 , n29597 , n207747 );
xnor ( n207749 , n29985 , n29987 );
xnor ( n29989 , n29982 , n207749 );
buf ( n29990 , n29989 );
buf ( n29991 , n29990 );
xor ( n29992 , n29971 , n29991 );
not ( n29993 , n29992 );
buf ( n29994 , RI17400870_1505);
not ( n29995 , n29994 );
not ( n29996 , n26146 );
or ( n29997 , n29995 , n29996 );
or ( n207759 , n26146 , n29994 );
nand ( n29999 , n29997 , n207759 );
buf ( n207761 , RI173c6478_1789);
not ( n30001 , n207761 );
not ( n30002 , RI1733cef8_2144);
not ( n30003 , n30002 );
or ( n30004 , n30001 , n30003 );
not ( n30005 , RI173c6478_1789);
buf ( n30006 , RI1733cef8_2144);
nand ( n30007 , n30005 , n30006 );
nand ( n30008 , n30004 , n30007 );
not ( n30009 , RI1740f168_1434);
and ( n207771 , n30008 , n30009 );
not ( n30011 , n30008 );
buf ( n30012 , RI1740f168_1434);
and ( n30013 , n30011 , n30012 );
nor ( n30014 , n207771 , n30013 );
buf ( n30015 , RI19ac30b0_2306);
nand ( n30016 , n25405 , n30015 );
buf ( n30017 , RI174ab798_900);
and ( n30018 , n30016 , n30017 );
not ( n30019 , n30016 );
not ( n30020 , RI174ab798_900);
and ( n30021 , n30019 , n30020 );
nor ( n207783 , n30018 , n30021 );
xor ( n30023 , n30014 , n207783 );
buf ( n207785 , n25529 );
buf ( n30025 , RI19a92e10_2662);
nand ( n30026 , n207785 , n30025 );
not ( n30027 , RI17462ac0_1255);
and ( n30028 , n30026 , n30027 );
not ( n30029 , n30026 );
buf ( n30030 , RI17462ac0_1255);
and ( n30031 , n30029 , n30030 );
nor ( n30032 , n30028 , n30031 );
xnor ( n30033 , n30023 , n30032 );
buf ( n30034 , n30033 );
not ( n207796 , n30034 );
and ( n30036 , n29999 , n207796 );
not ( n207798 , n29999 );
buf ( n30038 , n30034 );
and ( n30039 , n207798 , n30038 );
nor ( n30040 , n30036 , n30039 );
not ( n30041 , n30040 );
nand ( n30042 , n29993 , n30041 );
buf ( n30043 , RI173acd98_1913);
not ( n30044 , n30043 );
buf ( n30045 , RI173e74d8_1628);
not ( n207807 , n30045 );
not ( n30047 , RI1739e4a0_1984);
not ( n30048 , n30047 );
or ( n30049 , n207807 , n30048 );
not ( n30050 , RI173e74d8_1628);
buf ( n30051 , RI1739e4a0_1984);
nand ( n30052 , n30050 , n30051 );
nand ( n30053 , n30049 , n30052 );
buf ( n30054 , RI1745efb0_1273);
and ( n30055 , n30053 , n30054 );
not ( n30056 , n30053 );
not ( n207818 , RI1745efb0_1273);
and ( n30058 , n30056 , n207818 );
nor ( n207820 , n30055 , n30058 );
buf ( n30060 , RI19aa3ee0_2538);
nand ( n30061 , n25451 , n30060 );
buf ( n30062 , RI174837c0_1095);
and ( n30063 , n30061 , n30062 );
not ( n30064 , n30061 );
not ( n30065 , RI174837c0_1095);
and ( n30066 , n30064 , n30065 );
nor ( n30067 , n30063 , n30066 );
not ( n30068 , n30067 );
xor ( n30069 , n207820 , n30068 );
buf ( n30070 , RI19a852b0_2758);
nand ( n30071 , n207785 , n30070 );
not ( n30072 , RI175085a0_740);
and ( n30073 , n30071 , n30072 );
not ( n30074 , n30071 );
buf ( n30075 , RI175085a0_740);
and ( n30076 , n30074 , n30075 );
nor ( n30077 , n30073 , n30076 );
xnor ( n30078 , n30069 , n30077 );
not ( n30079 , n30078 );
or ( n30080 , n30044 , n30079 );
or ( n207842 , n30078 , n30043 );
nand ( n30082 , n30080 , n207842 );
not ( n207844 , n30082 );
not ( n30084 , RI173fb668_1530);
not ( n30085 , RI17404a10_1485);
buf ( n30086 , RI173bbd20_1840);
and ( n30087 , n30085 , n30086 );
not ( n30088 , n30085 );
not ( n30089 , RI173bbd20_1840);
and ( n30090 , n30088 , n30089 );
nor ( n30091 , n30087 , n30090 );
xor ( n207853 , n30084 , n30091 );
buf ( n30093 , RI173327a0_2195);
buf ( n207855 , RI174a0cf8_952);
xor ( n30095 , n30093 , n207855 );
buf ( n30096 , RI19ab5a00_2411);
nand ( n30097 , n29597 , n30096 );
xnor ( n30098 , n30095 , n30097 );
xnor ( n30099 , n207853 , n30098 );
buf ( n30100 , n30099 );
not ( n30101 , n30100 );
or ( n30102 , n207844 , n30101 );
or ( n30103 , n30100 , n30082 );
nand ( n30104 , n30102 , n30103 );
not ( n207866 , n30104 );
and ( n30106 , n30042 , n207866 );
not ( n207868 , n30042 );
and ( n30108 , n207868 , n30104 );
nor ( n30109 , n30106 , n30108 );
not ( n30110 , n30109 );
not ( n30111 , n204570 );
not ( n30112 , n28380 );
or ( n30113 , n30111 , n30112 );
or ( n30114 , n28380 , n204570 );
nand ( n30115 , n30113 , n30114 );
buf ( n30116 , RI1733f9a0_2131);
not ( n207878 , n30116 );
not ( n30118 , RI173c8f20_1776);
not ( n30119 , n30118 );
or ( n30120 , n207878 , n30119 );
not ( n30121 , RI1733f9a0_2131);
buf ( n30122 , RI173c8f20_1776);
nand ( n30123 , n30121 , n30122 );
nand ( n30124 , n30120 , n30123 );
buf ( n30125 , RI17411c10_1421);
and ( n30126 , n30124 , n30125 );
not ( n30127 , n30124 );
not ( n30128 , RI17411c10_1421);
and ( n30129 , n30127 , n30128 );
nor ( n207891 , n30126 , n30129 );
buf ( n30131 , RI19ac04a0_2329);
nand ( n207893 , n26242 , n30131 );
buf ( n30133 , RI174ae240_887);
xor ( n30134 , n207893 , n30133 );
xor ( n30135 , n207891 , n30134 );
xnor ( n30136 , n30135 , n28081 );
buf ( n30137 , n30136 );
and ( n30138 , n30115 , n30137 );
not ( n30139 , n30115 );
not ( n30140 , n30137 );
and ( n30141 , n30139 , n30140 );
nor ( n207903 , n30138 , n30141 );
not ( n30143 , n207903 );
not ( n207905 , n30143 );
not ( n30145 , n29225 );
buf ( n30146 , RI173c6e50_1786);
buf ( n30147 , RI173b6488_1867);
not ( n30148 , n30147 );
not ( n30149 , RI173ff4c0_1511);
not ( n30150 , n30149 );
or ( n30151 , n30148 , n30150 );
not ( n30152 , RI173b6488_1867);
buf ( n30153 , RI173ff4c0_1511);
nand ( n30154 , n30152 , n30153 );
nand ( n30155 , n30151 , n30154 );
xor ( n30156 , n30146 , n30155 );
buf ( n207918 , RI1752e0e8_623);
not ( n30158 , RI1749b7a8_978);
xor ( n30159 , n207918 , n30158 );
buf ( n30160 , RI19ab98d0_2384);
nand ( n30161 , n29203 , n30160 );
xnor ( n30162 , n30159 , n30161 );
xnor ( n30163 , n30156 , n30162 );
not ( n30164 , n30163 );
not ( n30165 , n30164 );
or ( n30166 , n30145 , n30165 );
or ( n30167 , n30164 , n29225 );
nand ( n30168 , n30166 , n30167 );
buf ( n207930 , RI173d3d20_1723);
not ( n30170 , n207930 );
not ( n207932 , RI1738b030_2078);
not ( n30172 , n207932 );
or ( n30173 , n30170 , n30172 );
not ( n30174 , RI173d3d20_1723);
buf ( n30175 , RI1738b030_2078);
nand ( n30176 , n30174 , n30175 );
nand ( n30177 , n30173 , n30176 );
and ( n30178 , n30177 , n27681 );
not ( n30179 , n30177 );
and ( n30180 , n30179 , n27722 );
nor ( n207942 , n30178 , n30180 );
buf ( n30182 , RI19acb648_2244);
nand ( n207944 , n25803 , n30182 );
buf ( n30184 , RI174b8f38_835);
and ( n30185 , n207944 , n30184 );
not ( n30186 , n207944 );
not ( n30187 , RI174b8f38_835);
and ( n30188 , n30186 , n30187 );
nor ( n30189 , n30185 , n30188 );
xor ( n30190 , n207942 , n30189 );
buf ( n30191 , RI19a9c398_2596);
nand ( n30192 , n28148 , n30191 );
buf ( n30193 , RI17470008_1190);
and ( n30194 , n30192 , n30193 );
not ( n30195 , n30192 );
not ( n30196 , RI17470008_1190);
and ( n30197 , n30195 , n30196 );
nor ( n30198 , n30194 , n30197 );
xnor ( n207960 , n30190 , n30198 );
buf ( n30200 , n207960 );
and ( n207962 , n30168 , n30200 );
not ( n30202 , n30168 );
xor ( n30203 , n207942 , n30198 );
not ( n30204 , n30189 );
xnor ( n30205 , n30203 , n30204 );
not ( n30206 , n30205 );
not ( n30207 , n30206 );
and ( n30208 , n30202 , n30207 );
nor ( n30209 , n207962 , n30208 );
not ( n207971 , n205151 );
not ( n30211 , n204436 );
or ( n30212 , n207971 , n30211 );
not ( n30213 , n205151 );
nand ( n30214 , n30213 , n204439 );
nand ( n30215 , n30212 , n30214 );
and ( n30216 , n30215 , n204391 );
not ( n30217 , n30215 );
xor ( n30218 , n204389 , n204361 );
buf ( n30219 , n204370 );
xnor ( n30220 , n30218 , n30219 );
and ( n30221 , n30217 , n30220 );
nor ( n30222 , n30216 , n30221 );
nand ( n30223 , n30209 , n30222 );
not ( n30224 , n30223 );
or ( n207986 , n207905 , n30224 );
or ( n30226 , n30223 , n30143 );
nand ( n30227 , n207986 , n30226 );
not ( n30228 , n30227 );
buf ( n30229 , RI173f22c0_1575);
buf ( n30230 , RI174039a8_1490);
not ( n30231 , n30230 );
not ( n30232 , RI173bacb8_1845);
not ( n30233 , n30232 );
or ( n30234 , n30231 , n30233 );
not ( n30235 , RI174039a8_1490);
buf ( n207997 , RI173bacb8_1845);
nand ( n30237 , n30235 , n207997 );
nand ( n207999 , n30234 , n30237 );
xor ( n30239 , n30229 , n207999 );
buf ( n30240 , RI17534d30_602);
buf ( n30241 , RI1749fc90_957);
xor ( n30242 , n30240 , n30241 );
buf ( n30243 , RI19ab7878_2398);
nand ( n30244 , n25880 , n30243 );
xnor ( n30245 , n30242 , n30244 );
xnor ( n30246 , n30239 , n30245 );
not ( n30247 , n30246 );
not ( n30248 , n25343 );
buf ( n30249 , RI173e6470_1633);
not ( n30250 , n30249 );
not ( n30251 , RI1739d438_1989);
not ( n30252 , n30251 );
or ( n30253 , n30250 , n30252 );
not ( n30254 , RI173e6470_1633);
buf ( n30255 , RI1739d438_1989);
nand ( n208017 , n30254 , n30255 );
nand ( n30257 , n30253 , n208017 );
buf ( n30258 , RI1745df48_1278);
and ( n30259 , n30257 , n30258 );
not ( n30260 , n30257 );
not ( n30261 , RI1745df48_1278);
and ( n208023 , n30260 , n30261 );
nor ( n30263 , n30259 , n208023 );
buf ( n208025 , RI19a84950_2762);
nand ( n30265 , n25364 , n208025 );
buf ( n30266 , RI17506bd8_745);
and ( n30267 , n30265 , n30266 );
not ( n30268 , n30265 );
not ( n30269 , RI17506bd8_745);
and ( n30270 , n30268 , n30269 );
nor ( n30271 , n30267 , n30270 );
xor ( n30272 , n30263 , n30271 );
buf ( n30273 , RI19aa3580_2542);
nand ( n208035 , n207785 , n30273 );
buf ( n30275 , RI17482758_1100);
and ( n208037 , n208035 , n30275 );
not ( n30277 , n208035 );
not ( n30278 , RI17482758_1100);
and ( n30279 , n30277 , n30278 );
nor ( n30280 , n208037 , n30279 );
xnor ( n30281 , n30272 , n30280 );
buf ( n30282 , n30281 );
not ( n30283 , n30282 );
or ( n30284 , n30248 , n30283 );
or ( n30285 , n30282 , n25343 );
nand ( n208047 , n30284 , n30285 );
xor ( n30287 , n30247 , n208047 );
buf ( n208049 , RI173f9f70_1537);
not ( n30289 , n208049 );
not ( n30290 , RI173b1280_1892);
not ( n30291 , n30290 );
or ( n30292 , n30289 , n30291 );
not ( n30293 , RI173f9f70_1537);
buf ( n30294 , RI173b1280_1892);
nand ( n30295 , n30293 , n30294 );
nand ( n30296 , n30292 , n30295 );
not ( n208058 , RI17392998_2041);
and ( n30298 , n30296 , n208058 );
not ( n208060 , n30296 );
buf ( n30300 , RI17392998_2041);
and ( n30301 , n208060 , n30300 );
nor ( n30302 , n30298 , n30301 );
buf ( n30303 , RI19a9b420_2603);
nand ( n30304 , n25451 , n30303 );
buf ( n30305 , RI17526000_648);
and ( n30306 , n30304 , n30305 );
not ( n30307 , n30304 );
not ( n30308 , RI17526000_648);
and ( n30309 , n30307 , n30308 );
nor ( n208071 , n30306 , n30309 );
xor ( n30311 , n30302 , n208071 );
buf ( n208073 , RI19aa9bb0_2498);
nand ( n30313 , n26463 , n208073 );
not ( n208075 , RI174965a0_1003);
and ( n30315 , n30313 , n208075 );
not ( n30316 , n30313 );
buf ( n30317 , RI174965a0_1003);
and ( n30318 , n30316 , n30317 );
nor ( n30319 , n30315 , n30318 );
xnor ( n30320 , n30311 , n30319 );
buf ( n30321 , n30320 );
not ( n30322 , n30321 );
not ( n30323 , n28979 );
buf ( n208085 , RI173dca38_1680);
not ( n30325 , n208085 );
not ( n30326 , RI17393d48_2035);
not ( n30327 , n30326 );
or ( n30328 , n30325 , n30327 );
not ( n30329 , RI173dca38_1680);
buf ( n30330 , RI17393d48_2035);
nand ( n30331 , n30329 , n30330 );
nand ( n30332 , n30328 , n30331 );
not ( n30333 , n30332 );
not ( n30334 , n30333 );
or ( n30335 , n30323 , n30334 );
or ( n30336 , n30333 , n28979 );
nand ( n30337 , n30335 , n30336 );
not ( n30338 , n30337 );
buf ( n208100 , RI17454510_1325);
buf ( n30340 , RI19a95de0_2641);
nand ( n208102 , n25375 , n30340 );
not ( n30342 , n208102 );
buf ( n30343 , RI17479068_1146);
not ( n30344 , n30343 );
and ( n30345 , n30342 , n30344 );
nand ( n30346 , n26058 , n30340 );
and ( n30347 , n30346 , n30343 );
nor ( n30348 , n30345 , n30347 );
xor ( n30349 , n208100 , n30348 );
buf ( n30350 , RI174c7218_791);
not ( n30351 , n30350 );
buf ( n30352 , RI19ac5bd0_2286);
nand ( n30353 , n25416 , n30352 );
not ( n30354 , n30353 );
or ( n208116 , n30351 , n30354 );
buf ( n30356 , n25375 );
nand ( n208118 , n30356 , n30352 );
or ( n30358 , n208118 , n30350 );
nand ( n30359 , n208116 , n30358 );
xnor ( n30360 , n30349 , n30359 );
not ( n30361 , n30360 );
not ( n30362 , n30361 );
or ( n30363 , n30338 , n30362 );
or ( n30364 , n30361 , n30337 );
nand ( n30365 , n30363 , n30364 );
not ( n30366 , n30365 );
and ( n208128 , n30322 , n30366 );
and ( n30368 , n30321 , n30365 );
nor ( n30369 , n208128 , n30368 );
nand ( n30370 , n30287 , n30369 );
not ( n30371 , n30370 );
buf ( n30372 , RI173ebd08_1606);
not ( n30373 , n30372 );
not ( n30374 , n205149 );
or ( n30375 , n30373 , n30374 );
not ( n30376 , RI173ebd08_1606);
buf ( n30377 , RI173a3018_1961);
nand ( n30378 , n30376 , n30377 );
nand ( n30379 , n30375 , n30378 );
buf ( n208141 , RI1747a0d0_1141);
and ( n30381 , n30379 , n208141 );
not ( n208143 , n30379 );
not ( n30383 , RI1747a0d0_1141);
and ( n30384 , n208143 , n30383 );
nor ( n30385 , n30381 , n30384 );
buf ( n30386 , RI19aa0100_2568);
nand ( n30387 , n29890 , n30386 );
buf ( n30388 , RI17487ff0_1073);
and ( n30389 , n30387 , n30388 );
not ( n30390 , n30387 );
not ( n30391 , RI17487ff0_1073);
and ( n30392 , n30390 , n30391 );
nor ( n208154 , n30389 , n30392 );
xor ( n30394 , n30385 , n208154 );
buf ( n30395 , RI19aced20_2219);
nand ( n30396 , n204336 , n30395 );
buf ( n30397 , RI1750f710_718);
and ( n30398 , n30396 , n30397 );
not ( n30399 , n30396 );
not ( n30400 , RI1750f710_718);
and ( n30401 , n30399 , n30400 );
nor ( n30402 , n30398 , n30401 );
not ( n30403 , n30402 );
xor ( n208165 , n30394 , n30403 );
buf ( n30405 , n208165 );
not ( n208167 , n30405 );
buf ( n30407 , n204294 );
not ( n208169 , n30407 );
buf ( n30409 , RI173ce7b8_1749);
not ( n30410 , n30409 );
not ( n30411 , RI17344ef0_2105);
not ( n30412 , n30411 );
or ( n30413 , n30410 , n30412 );
not ( n30414 , RI173ce7b8_1749);
buf ( n30415 , RI17344ef0_2105);
nand ( n30416 , n30414 , n30415 );
nand ( n30417 , n30413 , n30416 );
buf ( n208179 , RI174462a8_1394);
and ( n30419 , n30417 , n208179 );
not ( n208181 , n30417 );
not ( n30421 , RI174462a8_1394);
and ( n30422 , n208181 , n30421 );
nor ( n30423 , n30419 , n30422 );
buf ( n30424 , RI19a8bfe8_2711);
nand ( n30425 , n205124 , n30424 );
buf ( n30426 , RI1746aab8_1216);
and ( n30427 , n30425 , n30426 );
not ( n30428 , n30425 );
not ( n30429 , RI1746aab8_1216);
and ( n30430 , n30428 , n30429 );
nor ( n30431 , n30427 , n30430 );
xor ( n30432 , n30423 , n30431 );
buf ( n30433 , RI19abd4d0_2356);
nand ( n30434 , n25540 , n30433 );
buf ( n208196 , RI174b3790_861);
and ( n30436 , n30434 , n208196 );
not ( n208198 , n30434 );
not ( n30438 , RI174b3790_861);
and ( n30439 , n208198 , n30438 );
nor ( n30440 , n30436 , n30439 );
not ( n30441 , n30440 );
xnor ( n30442 , n30432 , n30441 );
not ( n30443 , n30442 );
or ( n30444 , n208169 , n30443 );
or ( n30445 , n30442 , n30407 );
nand ( n30446 , n30444 , n30445 );
not ( n30447 , n30446 );
or ( n30448 , n208167 , n30447 );
buf ( n208210 , n208165 );
or ( n30450 , n30446 , n208210 );
nand ( n208212 , n30448 , n30450 );
buf ( n30452 , n208212 );
not ( n30453 , n30452 );
and ( n30454 , n30371 , n30453 );
and ( n30455 , n30370 , n30452 );
nor ( n30456 , n30454 , n30455 );
not ( n30457 , n30456 );
or ( n30458 , n30228 , n30457 );
or ( n30459 , n30456 , n30227 );
nand ( n30460 , n30458 , n30459 );
not ( n30461 , n30460 );
buf ( n30462 , RI173cd408_1755);
not ( n30463 , n30462 );
not ( n30464 , RI17343e88_2110);
not ( n30465 , n30464 );
or ( n208227 , n30463 , n30465 );
not ( n30467 , RI173cd408_1755);
buf ( n208229 , RI17343e88_2110);
nand ( n30469 , n30467 , n208229 );
nand ( n30470 , n208227 , n30469 );
not ( n30471 , RI17445240_1399);
and ( n30472 , n30470 , n30471 );
not ( n30473 , n30470 );
buf ( n30474 , RI17445240_1399);
and ( n30475 , n30473 , n30474 );
nor ( n30476 , n30472 , n30475 );
buf ( n30477 , RI19a8dd70_2698);
nand ( n208239 , n25793 , n30477 );
not ( n30479 , RI17469a50_1221);
and ( n208241 , n208239 , n30479 );
not ( n30481 , n208239 );
buf ( n30482 , RI17469a50_1221);
and ( n30483 , n30481 , n30482 );
nor ( n30484 , n208241 , n30483 );
xor ( n30485 , n30476 , n30484 );
buf ( n30486 , RI19abebc8_2343);
nand ( n30487 , n27706 , n30486 );
not ( n30488 , RI174b2728_866);
and ( n30489 , n30487 , n30488 );
not ( n30490 , n30487 );
buf ( n30491 , RI174b2728_866);
and ( n30492 , n30490 , n30491 );
nor ( n30493 , n30489 , n30492 );
xnor ( n30494 , n30485 , n30493 );
not ( n30495 , n30494 );
not ( n30496 , n30495 );
not ( n30497 , n30496 );
not ( n30498 , n30497 );
not ( n30499 , n28651 );
buf ( n30500 , RI173f8bc0_1543);
not ( n30501 , n30500 );
not ( n208263 , RI173afed0_1898);
not ( n30503 , n208263 );
or ( n208265 , n30501 , n30503 );
not ( n30505 , RI173f8bc0_1543);
buf ( n30506 , RI173afed0_1898);
nand ( n30507 , n30505 , n30506 );
nand ( n30508 , n208265 , n30507 );
not ( n30509 , RI17346930_2097);
and ( n30510 , n30508 , n30509 );
not ( n30511 , n30508 );
buf ( n30512 , RI17346930_2097);
and ( n208274 , n30511 , n30512 );
nor ( n30514 , n30510 , n208274 );
buf ( n208276 , RI19aac388_2481);
nand ( n30516 , n25915 , n208276 );
buf ( n30517 , RI17524110_654);
and ( n30518 , n30516 , n30517 );
not ( n30519 , n30516 );
not ( n30520 , RI17524110_654);
and ( n30521 , n30519 , n30520 );
nor ( n30522 , n30518 , n30521 );
xor ( n30523 , n30514 , n30522 );
buf ( n30524 , RI19aab5f0_2486);
nand ( n30525 , n29203 , n30524 );
buf ( n30526 , RI174951f0_1009);
and ( n30527 , n30525 , n30526 );
not ( n208289 , n30525 );
not ( n30529 , RI174951f0_1009);
and ( n208291 , n208289 , n30529 );
nor ( n30531 , n30527 , n208291 );
xor ( n30532 , n30523 , n30531 );
not ( n30533 , n30532 );
not ( n30534 , n30533 );
not ( n30535 , n30534 );
or ( n30536 , n30499 , n30535 );
not ( n30537 , n30533 );
or ( n30538 , n30537 , n28651 );
nand ( n30539 , n30536 , n30538 );
not ( n208301 , n30539 );
or ( n30541 , n30498 , n208301 );
buf ( n208303 , n30494 );
not ( n30543 , n208303 );
or ( n30544 , n30539 , n30543 );
nand ( n30545 , n30541 , n30544 );
not ( n30546 , n30545 );
buf ( n30547 , RI173dc6f0_1681);
not ( n30548 , n30547 );
not ( n30549 , RI17393a00_2036);
not ( n30550 , n30549 );
or ( n30551 , n30548 , n30550 );
not ( n30552 , RI173dc6f0_1681);
buf ( n30553 , RI17393a00_2036);
nand ( n30554 , n30552 , n30553 );
nand ( n30555 , n30551 , n30554 );
not ( n30556 , RI174541c8_1326);
and ( n30557 , n30555 , n30556 );
not ( n30558 , n30555 );
buf ( n208320 , RI174541c8_1326);
and ( n30560 , n30558 , n208320 );
nor ( n30561 , n30557 , n30560 );
buf ( n30562 , RI19a95b88_2642);
nand ( n30563 , n26028 , n30562 );
buf ( n30564 , RI17478d20_1147);
and ( n30565 , n30563 , n30564 );
not ( n30566 , n30563 );
not ( n30567 , RI17478d20_1147);
and ( n30568 , n30566 , n30567 );
nor ( n30569 , n30565 , n30568 );
xor ( n30570 , n30561 , n30569 );
buf ( n30571 , RI19ac5978_2287);
nand ( n30572 , n25376 , n30571 );
not ( n30573 , RI174c6cf0_792);
and ( n30574 , n30572 , n30573 );
not ( n30575 , n30572 );
buf ( n30576 , RI174c6cf0_792);
and ( n30577 , n30575 , n30576 );
nor ( n30578 , n30574 , n30577 );
xnor ( n30579 , n30570 , n30578 );
buf ( n30580 , n30579 );
not ( n30581 , n30580 );
not ( n30582 , n30581 );
xor ( n30583 , n25687 , n30582 );
not ( n30584 , RI17407e90_1469);
and ( n30585 , n30584 , n27804 );
not ( n30586 , n30584 );
and ( n30587 , n30586 , n205610 );
nor ( n208349 , n30585 , n30587 );
not ( n30589 , n208349 );
not ( n30590 , n30589 );
not ( n30591 , RI1744c518_1364);
xor ( n30592 , n28198 , n30591 );
buf ( n30593 , RI19ab5820_2412);
nand ( n30594 , n25491 , n30593 );
not ( n30595 , RI174a4178_936);
and ( n30596 , n30594 , n30595 );
not ( n30597 , n30594 );
buf ( n30598 , RI174a4178_936);
and ( n30599 , n30597 , n30598 );
nor ( n30600 , n30596 , n30599 );
xnor ( n30601 , n30592 , n30600 );
not ( n30602 , n30601 );
not ( n30603 , n30602 );
or ( n30604 , n30590 , n30603 );
nand ( n30605 , n30601 , n208349 );
nand ( n30606 , n30604 , n30605 );
not ( n30607 , n30606 );
not ( n30608 , n30607 );
xnor ( n208370 , n30583 , n30608 );
nand ( n30610 , n30546 , n208370 );
not ( n30611 , n30610 );
buf ( n30612 , RI17332110_2197);
buf ( n30613 , RI1740b658_1452);
not ( n30614 , n30613 );
not ( n30615 , RI173c2968_1807);
not ( n30616 , n30615 );
or ( n30617 , n30614 , n30616 );
not ( n30618 , RI1740b658_1452);
buf ( n208380 , RI173c2968_1807);
nand ( n30620 , n30618 , n208380 );
nand ( n208382 , n30617 , n30620 );
xor ( n30622 , n30612 , n208382 );
buf ( n30623 , RI19ab2f58_2432);
nand ( n30624 , n204512 , n30623 );
buf ( n30625 , RI174a7c88_918);
and ( n30626 , n30624 , n30625 );
not ( n30627 , n30624 );
not ( n30628 , RI174a7c88_918);
and ( n30629 , n30627 , n30628 );
nor ( n30630 , n30626 , n30629 );
not ( n30631 , n30630 );
buf ( n30632 , RI173393e8_2162);
not ( n30633 , n30632 );
and ( n30634 , n30631 , n30633 );
and ( n208396 , n30630 , n30632 );
nor ( n30636 , n30634 , n208396 );
xnor ( n208398 , n30622 , n30636 );
not ( n30638 , n208398 );
not ( n30639 , n30638 );
buf ( n30640 , n25655 );
buf ( n30641 , n30640 );
buf ( n30642 , RI19a93518_2659);
nand ( n30643 , n30641 , n30642 );
not ( n30644 , RI17529de0_636);
and ( n30645 , n30643 , n30644 );
not ( n208407 , n30643 );
buf ( n30647 , RI17529de0_636);
and ( n208409 , n208407 , n30647 );
nor ( n30649 , n30645 , n208409 );
buf ( n30650 , n30649 );
not ( n30651 , n30650 );
buf ( n30652 , RI173a5430_1950);
not ( n30653 , n30652 );
not ( n30654 , RI173ee120_1595);
not ( n30655 , n30654 );
or ( n30656 , n30653 , n30655 );
not ( n30657 , RI173a5430_1950);
buf ( n208419 , RI173ee120_1595);
nand ( n30659 , n30657 , n208419 );
nand ( n30660 , n30656 , n30659 );
buf ( n30661 , RI17490d08_1030);
and ( n30662 , n30660 , n30661 );
not ( n30663 , n30660 );
not ( n30664 , RI17490d08_1030);
and ( n30665 , n30663 , n30664 );
nor ( n30666 , n30662 , n30665 );
buf ( n30667 , RI19a9f368_2575);
nand ( n30668 , n25364 , n30667 );
buf ( n30669 , RI1748a408_1062);
and ( n30670 , n30668 , n30669 );
not ( n30671 , n30668 );
not ( n30672 , RI1748a408_1062);
and ( n30673 , n30671 , n30672 );
nor ( n30674 , n30670 , n30673 );
xor ( n30675 , n30666 , n30674 );
buf ( n30676 , RI19acdf10_2225);
nand ( n30677 , n26325 , n30676 );
not ( n30678 , RI175134f0_706);
and ( n30679 , n30677 , n30678 );
not ( n208441 , n30677 );
buf ( n30681 , RI175134f0_706);
and ( n208443 , n208441 , n30681 );
nor ( n30683 , n30679 , n208443 );
xnor ( n208445 , n30675 , n30683 );
not ( n30685 , n208445 );
not ( n30686 , n30685 );
or ( n30687 , n30651 , n30686 );
not ( n30688 , n30650 );
buf ( n30689 , n208445 );
nand ( n30690 , n30688 , n30689 );
nand ( n30691 , n30687 , n30690 );
not ( n30692 , n30691 );
and ( n30693 , n30639 , n30692 );
not ( n30694 , n208398 );
and ( n30695 , n30694 , n30691 );
nor ( n30696 , n30693 , n30695 );
not ( n30697 , n30696 );
not ( n208459 , n30697 );
and ( n30699 , n30611 , n208459 );
not ( n208461 , n30545 );
nand ( n30701 , n208461 , n208370 );
and ( n30702 , n30701 , n30697 );
nor ( n30703 , n30699 , n30702 );
not ( n30704 , n30703 );
or ( n30705 , n30461 , n30704 );
or ( n30706 , n30703 , n30460 );
nand ( n30707 , n30705 , n30706 );
nand ( n30708 , n30040 , n207866 );
not ( n208470 , n30708 );
buf ( n30710 , RI19a87470_2743);
nand ( n30711 , n204513 , n30710 );
not ( n30712 , RI174d0cc8_761);
and ( n30713 , n30711 , n30712 );
not ( n30714 , n30711 );
buf ( n30715 , RI174d0cc8_761);
and ( n30716 , n30714 , n30715 );
nor ( n30717 , n30713 , n30716 );
not ( n30718 , n30717 );
not ( n30719 , n205383 );
or ( n208481 , n30718 , n30719 );
not ( n30721 , n30717 );
nand ( n30722 , n30721 , n205389 );
nand ( n30723 , n208481 , n30722 );
buf ( n30724 , RI173f18e8_1578);
not ( n30725 , n30724 );
not ( n30726 , RI173a8bf8_1933);
not ( n30727 , n30726 );
or ( n30728 , n30725 , n30727 );
not ( n30729 , RI173f18e8_1578);
buf ( n30730 , RI173a8bf8_1933);
nand ( n30731 , n30729 , n30730 );
nand ( n30732 , n30728 , n30731 );
not ( n30733 , RI174b51d0_853);
and ( n30734 , n30732 , n30733 );
not ( n30735 , n30732 );
buf ( n208497 , RI174b51d0_853);
and ( n30737 , n30735 , n208497 );
nor ( n30738 , n30734 , n30737 );
buf ( n30739 , RI19ab0528_2451);
nand ( n30740 , n204493 , n30739 );
buf ( n30741 , RI1748dbd0_1045);
and ( n30742 , n30740 , n30741 );
not ( n30743 , n30740 );
not ( n30744 , RI1748dbd0_1045);
and ( n208506 , n30743 , n30744 );
nor ( n208507 , n30742 , n208506 );
xor ( n30747 , n30738 , n208507 );
buf ( n30748 , RI19ab3a20_2426);
nand ( n30749 , n204393 , n30748 );
not ( n208511 , RI17518c98_689);
and ( n30751 , n30749 , n208511 );
not ( n208513 , n30749 );
buf ( n30753 , RI17518c98_689);
and ( n30754 , n208513 , n30753 );
nor ( n30755 , n30751 , n30754 );
xnor ( n30756 , n30747 , n30755 );
buf ( n30757 , n30756 );
and ( n30758 , n30723 , n30757 );
not ( n30759 , n30723 );
not ( n30760 , n208507 );
not ( n30761 , n30755 );
or ( n30762 , n30760 , n30761 );
or ( n30763 , n208507 , n30755 );
nand ( n30764 , n30762 , n30763 );
not ( n30765 , n30738 );
and ( n30766 , n30764 , n30765 );
not ( n30767 , n30764 );
and ( n30768 , n30767 , n30738 );
nor ( n30769 , n30766 , n30768 );
not ( n30770 , n30769 );
not ( n30771 , n30770 );
and ( n208533 , n30759 , n30771 );
nor ( n30773 , n30758 , n208533 );
not ( n208535 , n30773 );
not ( n30775 , n208535 );
and ( n30776 , n208470 , n30775 );
and ( n30777 , n30708 , n208535 );
nor ( n30778 , n30776 , n30777 );
not ( n30779 , n30778 );
buf ( n30780 , n28554 );
not ( n30781 , n29607 );
xor ( n30782 , n30780 , n30781 );
not ( n30783 , RI174122a0_1419);
buf ( n208545 , RI173be138_1829);
not ( n30785 , n208545 );
not ( n30786 , RI17406e28_1474);
not ( n30787 , n30786 );
or ( n30788 , n30785 , n30787 );
not ( n30789 , RI173be138_1829);
buf ( n30790 , RI17406e28_1474);
nand ( n30791 , n30789 , n30790 );
nand ( n208553 , n30788 , n30791 );
xor ( n30793 , n30783 , n208553 );
not ( n30794 , RI17334bb8_2184);
not ( n30795 , n30794 );
buf ( n30796 , RI19ab4bf0_2418);
nand ( n30797 , n29890 , n30796 );
not ( n30798 , RI174a3110_941);
and ( n30799 , n30797 , n30798 );
not ( n30800 , n30797 );
buf ( n30801 , RI174a3110_941);
and ( n30802 , n30800 , n30801 );
nor ( n30803 , n30799 , n30802 );
not ( n208565 , n30803 );
or ( n30805 , n30795 , n208565 );
or ( n208567 , n30803 , n30794 );
nand ( n30807 , n30805 , n208567 );
xnor ( n30808 , n30793 , n30807 );
buf ( n30809 , n30808 );
not ( n30810 , n30809 );
xnor ( n30811 , n30782 , n30810 );
not ( n30812 , n30811 );
not ( n30813 , RI1738c728_2071);
not ( n30814 , n30813 );
not ( n30815 , n30814 );
buf ( n208577 , RI173c67c0_1788);
not ( n30817 , n208577 );
not ( n208579 , RI1733d240_2143);
not ( n30819 , n208579 );
or ( n30820 , n30817 , n30819 );
not ( n30821 , RI173c67c0_1788);
buf ( n30822 , RI1733d240_2143);
nand ( n30823 , n30821 , n30822 );
nand ( n30824 , n30820 , n30823 );
buf ( n30825 , RI1740f4b0_1433);
and ( n30826 , n30824 , n30825 );
not ( n30827 , n30824 );
not ( n30828 , RI1740f4b0_1433);
and ( n30829 , n30827 , n30828 );
nor ( n30830 , n30826 , n30829 );
buf ( n30831 , RI19a90a70_2678);
nand ( n30832 , n204572 , n30831 );
not ( n30833 , RI17462e08_1254);
and ( n30834 , n30832 , n30833 );
not ( n208596 , n30832 );
buf ( n30836 , RI17462e08_1254);
and ( n30837 , n208596 , n30836 );
nor ( n30838 , n30834 , n30837 );
xor ( n30839 , n30830 , n30838 );
buf ( n30840 , RI19ac0f68_2323);
nand ( n30841 , n25916 , n30840 );
not ( n30842 , RI174abae0_899);
and ( n30843 , n30841 , n30842 );
not ( n30844 , n30841 );
buf ( n30845 , RI174abae0_899);
and ( n30846 , n30844 , n30845 );
nor ( n30847 , n30843 , n30846 );
xnor ( n30848 , n30839 , n30847 );
not ( n208610 , n30848 );
not ( n30850 , n208610 );
not ( n208612 , n30850 );
or ( n30852 , n30815 , n208612 );
not ( n30853 , n208610 );
or ( n30854 , n30853 , n30814 );
nand ( n30855 , n30852 , n30854 );
buf ( n30856 , RI173e3d10_1645);
not ( n30857 , n30856 );
not ( n30858 , RI1739b020_2000);
not ( n30859 , n30858 );
or ( n208621 , n30857 , n30859 );
not ( n30861 , RI173e3d10_1645);
buf ( n208623 , RI1739b020_2000);
nand ( n30863 , n30861 , n208623 );
nand ( n30864 , n208621 , n30863 );
buf ( n30865 , RI1745bb30_1289);
and ( n30866 , n30864 , n30865 );
not ( n30867 , n30864 );
not ( n30868 , RI1745bb30_1289);
and ( n30869 , n30867 , n30868 );
nor ( n30870 , n30866 , n30869 );
buf ( n30871 , RI19a859b8_2755);
nand ( n30872 , n25529 , n30871 );
not ( n30873 , RI175014a8_756);
and ( n30874 , n30872 , n30873 );
not ( n208636 , n30872 );
buf ( n30876 , RI175014a8_756);
and ( n30877 , n208636 , n30876 );
nor ( n30878 , n30874 , n30877 );
xor ( n30879 , n30870 , n30878 );
buf ( n208641 , RI19aa46d8_2534);
nand ( n30881 , n204916 , n208641 );
buf ( n208643 , RI17480340_1111);
and ( n30883 , n30881 , n208643 );
not ( n30884 , n30881 );
not ( n30885 , RI17480340_1111);
and ( n30886 , n30884 , n30885 );
nor ( n30887 , n30883 , n30886 );
xor ( n30888 , n30879 , n30887 );
not ( n30889 , n30888 );
not ( n30890 , n30889 );
and ( n30891 , n30855 , n30890 );
not ( n208653 , n30855 );
not ( n30893 , n30890 );
and ( n208655 , n208653 , n30893 );
nor ( n30895 , n30891 , n208655 );
buf ( n30896 , n205033 );
not ( n30897 , n30896 );
buf ( n30898 , n30897 );
not ( n30899 , n30898 );
buf ( n30900 , RI173e50c0_1639);
not ( n30901 , n30900 );
buf ( n30902 , RI173d6480_1711);
not ( n30903 , n30902 );
not ( n30904 , RI1738d790_2066);
not ( n30905 , n30904 );
or ( n30906 , n30903 , n30905 );
not ( n30907 , RI173d6480_1711);
buf ( n30908 , RI1738d790_2066);
nand ( n30909 , n30907 , n30908 );
nand ( n30910 , n30906 , n30909 );
buf ( n208672 , RI1744df58_1356);
and ( n30912 , n30910 , n208672 );
not ( n30913 , n30910 );
not ( n30914 , RI1744df58_1356);
and ( n30915 , n30913 , n30914 );
nor ( n30916 , n30912 , n30915 );
not ( n30917 , n30916 );
buf ( n30918 , RI19acadd8_2249);
nand ( n30919 , n25622 , n30918 );
buf ( n30920 , RI174bcd18_823);
and ( n30921 , n30919 , n30920 );
not ( n30922 , n30919 );
not ( n30923 , RI174bcd18_823);
and ( n30924 , n30922 , n30923 );
nor ( n30925 , n30921 , n30924 );
xor ( n208687 , n30917 , n30925 );
buf ( n30927 , RI19a9b8d0_2601);
nand ( n208689 , n25793 , n30927 );
buf ( n30929 , RI17472768_1178);
and ( n30930 , n208689 , n30929 );
not ( n30931 , n208689 );
not ( n30932 , RI17472768_1178);
and ( n30933 , n30931 , n30932 );
nor ( n30934 , n30930 , n30933 );
not ( n30935 , n30934 );
xnor ( n30936 , n208687 , n30935 );
not ( n30937 , n30936 );
or ( n208699 , n30901 , n30937 );
not ( n30939 , n30900 );
xor ( n208701 , n30916 , n30934 );
not ( n30941 , n30925 );
xnor ( n30942 , n208701 , n30941 );
buf ( n30943 , n30942 );
nand ( n30944 , n30939 , n30943 );
nand ( n30945 , n208699 , n30944 );
not ( n30946 , n30945 );
or ( n30947 , n30899 , n30946 );
or ( n30948 , n30945 , n30898 );
nand ( n208710 , n30947 , n30948 );
nand ( n30950 , n30895 , n208710 );
not ( n30951 , n30950 );
or ( n30952 , n30812 , n30951 );
or ( n30953 , n30950 , n30811 );
nand ( n30954 , n30952 , n30953 );
not ( n30955 , n30954 );
or ( n30956 , n30779 , n30955 );
or ( n30957 , n30954 , n30778 );
nand ( n30958 , n30956 , n30957 );
not ( n30959 , n30958 );
and ( n30960 , n30707 , n30959 );
not ( n30961 , n30707 );
and ( n30962 , n30961 , n30958 );
nor ( n30963 , n30960 , n30962 );
buf ( n208725 , n30963 );
not ( n30965 , n208725 );
or ( n208727 , n30110 , n30965 );
not ( n30967 , n30109 );
not ( n30968 , n30963 );
nand ( n30969 , n30967 , n30968 );
nand ( n30970 , n208727 , n30969 );
buf ( n30971 , n208610 );
not ( n30972 , n30971 );
not ( n30973 , n30972 );
buf ( n30974 , RI17400bb8_1504);
not ( n30975 , n30974 );
buf ( n30976 , RI173f1f78_1576);
not ( n30977 , n30976 );
not ( n30978 , RI173a9288_1931);
not ( n30979 , n30978 );
or ( n30980 , n30977 , n30979 );
not ( n30981 , RI173f1f78_1576);
buf ( n30982 , RI173a9288_1931);
nand ( n30983 , n30981 , n30982 );
nand ( n30984 , n30980 , n30983 );
buf ( n30985 , RI174ba3d8_831);
and ( n30986 , n30984 , n30985 );
not ( n30987 , n30984 );
not ( n30988 , RI174ba3d8_831);
and ( n30989 , n30987 , n30988 );
nor ( n30990 , n30986 , n30989 );
buf ( n30991 , RI19ab0a50_2449);
nand ( n208753 , n206902 , n30991 );
buf ( n30993 , RI1748e260_1043);
and ( n208755 , n208753 , n30993 );
not ( n30995 , n208753 );
not ( n30996 , RI1748e260_1043);
and ( n30997 , n30995 , n30996 );
nor ( n30998 , n208755 , n30997 );
xor ( n30999 , n30990 , n30998 );
buf ( n31000 , RI19ad0238_2210);
nand ( n31001 , n25416 , n31000 );
not ( n31002 , RI175196e8_687);
and ( n31003 , n31001 , n31002 );
not ( n31004 , n31001 );
buf ( n31005 , RI175196e8_687);
and ( n31006 , n31004 , n31005 );
nor ( n31007 , n31003 , n31006 );
xor ( n31008 , n30999 , n31007 );
not ( n31009 , n31008 );
or ( n31010 , n30975 , n31009 );
or ( n31011 , n31008 , n30974 );
nand ( n31012 , n31010 , n31011 );
not ( n31013 , n31012 );
or ( n31014 , n30973 , n31013 );
not ( n208776 , n30971 );
or ( n31016 , n31012 , n208776 );
nand ( n208778 , n31014 , n31016 );
not ( n31018 , n208778 );
buf ( n31019 , RI173eb678_1608);
buf ( n31020 , RI173ba2e0_1848);
not ( n31021 , n31020 );
not ( n31022 , RI17402fd0_1493);
not ( n31023 , n31022 );
or ( n31024 , n31021 , n31023 );
not ( n31025 , RI173ba2e0_1848);
buf ( n31026 , RI17402fd0_1493);
nand ( n31027 , n31025 , n31026 );
nand ( n31028 , n31024 , n31027 );
xor ( n208790 , n31019 , n31028 );
buf ( n31030 , RI17533db8_605);
not ( n208792 , RI1749f2b8_960);
xor ( n31032 , n31030 , n208792 );
buf ( n31033 , RI19ab71e8_2401);
nand ( n31034 , n30641 , n31033 );
xnor ( n31035 , n31032 , n31034 );
xnor ( n31036 , n208790 , n31035 );
not ( n31037 , n31036 );
not ( n31038 , n31037 );
buf ( n31039 , RI17411580_1423);
not ( n31040 , n31039 );
and ( n31041 , n31038 , n31040 );
and ( n31042 , n31037 , n31039 );
nor ( n31043 , n31041 , n31042 );
buf ( n31044 , RI173d7830_1705);
not ( n31045 , n31044 );
not ( n31046 , RI1738eb40_2060);
not ( n31047 , n31046 );
or ( n31048 , n31045 , n31047 );
not ( n31049 , RI173d7830_1705);
buf ( n31050 , RI1738eb40_2060);
nand ( n31051 , n31049 , n31050 );
nand ( n31052 , n31048 , n31051 );
not ( n31053 , n31052 );
buf ( n31054 , RI1744f308_1350);
buf ( n31055 , RI19ac9500_2260);
nand ( n208817 , n25741 , n31055 );
buf ( n31057 , RI174bf130_816);
and ( n208819 , n208817 , n31057 );
not ( n31059 , n208817 );
not ( n31060 , RI174bf130_816);
and ( n31061 , n31059 , n31060 );
nor ( n31062 , n208819 , n31061 );
xor ( n31063 , n31054 , n31062 );
buf ( n31064 , RI19a99d28_2613);
nand ( n31065 , n29203 , n31064 );
not ( n31066 , RI17473b18_1172);
and ( n31067 , n31065 , n31066 );
not ( n208829 , n31065 );
buf ( n31069 , RI17473b18_1172);
and ( n31070 , n208829 , n31069 );
nor ( n31071 , n31067 , n31070 );
xnor ( n31072 , n31063 , n31071 );
and ( n31073 , n31053 , n31072 );
not ( n31074 , n31053 );
not ( n31075 , n31072 );
and ( n31076 , n31074 , n31075 );
nor ( n31077 , n31073 , n31076 );
buf ( n31078 , n31077 );
and ( n31079 , n31043 , n31078 );
not ( n31080 , n31043 );
not ( n31081 , n31078 );
and ( n208843 , n31080 , n31081 );
nor ( n31083 , n31079 , n208843 );
not ( n31084 , n31083 );
nand ( n31085 , n31084 , n25981 );
not ( n31086 , n31085 );
or ( n31087 , n31018 , n31086 );
or ( n31088 , n31085 , n208778 );
nand ( n31089 , n31087 , n31088 );
not ( n31090 , n31089 );
buf ( n31091 , RI173b0218_1897);
not ( n208853 , n31091 );
buf ( n31093 , RI173ee7b0_1593);
not ( n208855 , n31093 );
not ( n31095 , RI173a5ac0_1948);
not ( n31096 , n31095 );
or ( n31097 , n208855 , n31096 );
not ( n31098 , RI173ee7b0_1593);
buf ( n31099 , RI173a5ac0_1948);
nand ( n31100 , n31098 , n31099 );
nand ( n31101 , n31097 , n31100 );
not ( n31102 , RI17495538_1008);
and ( n31103 , n31101 , n31102 );
not ( n31104 , n31101 );
buf ( n31105 , RI17495538_1008);
and ( n208867 , n31104 , n31105 );
nor ( n31107 , n31103 , n208867 );
buf ( n208869 , RI19ace3c0_2223);
nand ( n31109 , n29890 , n208869 );
buf ( n31110 , RI17513f40_704);
and ( n31111 , n31109 , n31110 );
not ( n31112 , n31109 );
not ( n31113 , RI17513f40_704);
and ( n31114 , n31112 , n31113 );
nor ( n31115 , n31111 , n31114 );
xor ( n31116 , n31107 , n31115 );
buf ( n31117 , RI19a9f728_2573);
nand ( n31118 , n26463 , n31117 );
not ( n31119 , RI1748aa98_1060);
and ( n31120 , n31118 , n31119 );
not ( n31121 , n31118 );
buf ( n208883 , RI1748aa98_1060);
and ( n31123 , n31121 , n208883 );
nor ( n208885 , n31120 , n31123 );
xnor ( n31125 , n31116 , n208885 );
not ( n31126 , n31125 );
not ( n31127 , n31126 );
not ( n31128 , n31127 );
or ( n31129 , n208853 , n31128 );
or ( n31130 , n31127 , n31091 );
nand ( n31131 , n31129 , n31130 );
and ( n31132 , n31131 , n29694 );
not ( n31133 , n31131 );
xor ( n31134 , n29666 , n29675 );
xnor ( n31135 , n31134 , n29692 );
buf ( n31136 , n31135 );
buf ( n31137 , n31136 );
and ( n31138 , n31133 , n31137 );
nor ( n31139 , n31132 , n31138 );
not ( n31140 , n31139 );
nand ( n31141 , n31140 , n26414 );
not ( n31142 , n31141 );
buf ( n208904 , RI173e5408_1638);
buf ( n31144 , RI173f3d00_1567);
not ( n208906 , n31144 );
not ( n31146 , RI173ab010_1922);
not ( n31147 , n31146 );
or ( n31148 , n208906 , n31147 );
not ( n31149 , RI173f3d00_1567);
buf ( n31150 , RI173ab010_1922);
nand ( n31151 , n31149 , n31150 );
nand ( n31152 , n31148 , n31151 );
not ( n31153 , RI17507b50_742);
and ( n31154 , n31152 , n31153 );
not ( n208916 , n31152 );
buf ( n31156 , RI17507b50_742);
and ( n31157 , n208916 , n31156 );
nor ( n31158 , n31154 , n31157 );
buf ( n31159 , RI19aaf790_2457);
nand ( n31160 , n204916 , n31159 );
buf ( n31161 , RI17490330_1033);
and ( n31162 , n31160 , n31161 );
not ( n31163 , n31160 );
not ( n31164 , RI17490330_1033);
and ( n31165 , n31163 , n31164 );
nor ( n31166 , n31162 , n31165 );
xor ( n31167 , n31158 , n31166 );
buf ( n31168 , RI19a83b40_2768);
nand ( n31169 , n26266 , n31168 );
buf ( n31170 , RI1751c550_678);
and ( n31171 , n31169 , n31170 );
not ( n31172 , n31169 );
not ( n208934 , RI1751c550_678);
and ( n31174 , n31172 , n208934 );
nor ( n208936 , n31171 , n31174 );
xor ( n31176 , n31167 , n208936 );
buf ( n31177 , n31176 );
xor ( n31178 , n208904 , n31177 );
buf ( n31179 , RI1744e2a0_1355);
buf ( n31180 , RI173d67c8_1710);
not ( n31181 , n31180 );
not ( n31182 , RI1738dad8_2065);
not ( n208944 , n31182 );
or ( n31184 , n31181 , n208944 );
not ( n208946 , RI173d67c8_1710);
buf ( n31186 , RI1738dad8_2065);
nand ( n31187 , n208946 , n31186 );
nand ( n31188 , n31184 , n31187 );
xor ( n31189 , n31179 , n31188 );
buf ( n31190 , RI19acaf40_2248);
nand ( n31191 , n25628 , n31190 );
buf ( n31192 , RI174bd240_822);
and ( n31193 , n31191 , n31192 );
not ( n31194 , n31191 );
not ( n31195 , RI174bd240_822);
and ( n31196 , n31194 , n31195 );
nor ( n31197 , n31193 , n31196 );
not ( n31198 , n31197 );
buf ( n31199 , RI19a9bb28_2600);
nand ( n31200 , n25529 , n31199 );
buf ( n31201 , RI17472ab0_1177);
and ( n31202 , n31200 , n31201 );
not ( n31203 , n31200 );
not ( n31204 , RI17472ab0_1177);
and ( n31205 , n31203 , n31204 );
nor ( n31206 , n31202 , n31205 );
not ( n31207 , n31206 );
not ( n31208 , n31207 );
or ( n31209 , n31198 , n31208 );
not ( n31210 , n31197 );
nand ( n31211 , n31206 , n31210 );
nand ( n31212 , n31209 , n31211 );
xnor ( n31213 , n31189 , n31212 );
xnor ( n31214 , n31178 , n31213 );
not ( n31215 , n31214 );
not ( n31216 , n31215 );
and ( n31217 , n31142 , n31216 );
and ( n31218 , n31141 , n31215 );
nor ( n208980 , n31217 , n31218 );
not ( n31220 , n208980 );
and ( n208982 , n31090 , n31220 );
and ( n31222 , n31089 , n208980 );
nor ( n31223 , n208982 , n31222 );
not ( n31224 , n31223 );
buf ( n31225 , RI1744b4b0_1369);
not ( n31226 , n31225 );
buf ( n31227 , n207012 );
not ( n31228 , n31227 );
or ( n31229 , n31226 , n31228 );
or ( n208991 , n31227 , n31225 );
nand ( n31231 , n31229 , n208991 );
and ( n31232 , n31231 , n29258 );
not ( n31233 , n31231 );
and ( n31234 , n31233 , n29214 );
nor ( n31235 , n31232 , n31234 );
nand ( n31236 , n25872 , n31235 );
not ( n31237 , n31236 );
not ( n208999 , n27769 );
buf ( n31239 , RI1744e930_1353);
not ( n209001 , RI174081d8_1468);
buf ( n31241 , RI173bf4e8_1823);
nand ( n31242 , n209001 , n31241 );
not ( n31243 , RI173bf4e8_1823);
buf ( n31244 , RI174081d8_1468);
nand ( n31245 , n31243 , n31244 );
and ( n31246 , n31242 , n31245 );
xor ( n31247 , n31239 , n31246 );
buf ( n31248 , RI174a44c0_935);
xor ( n31249 , n29263 , n31248 );
buf ( n31250 , RI19ab3318_2430);
nand ( n31251 , n207785 , n31250 );
xnor ( n31252 , n31249 , n31251 );
xnor ( n31253 , n31247 , n31252 );
not ( n31254 , n31253 );
not ( n31255 , n31254 );
or ( n31256 , n208999 , n31255 );
or ( n31257 , n31254 , n27769 );
nand ( n31258 , n31256 , n31257 );
not ( n31259 , n30360 );
not ( n31260 , n30333 );
and ( n31261 , n31259 , n31260 );
and ( n31262 , n30360 , n30333 );
nor ( n31263 , n31261 , n31262 );
buf ( n31264 , n31263 );
and ( n31265 , n31258 , n31264 );
not ( n31266 , n31258 );
not ( n31267 , n30332 );
not ( n31268 , n30360 );
not ( n31269 , n31268 );
or ( n209031 , n31267 , n31269 );
nand ( n31271 , n30360 , n30333 );
nand ( n209033 , n209031 , n31271 );
buf ( n31273 , n209033 );
and ( n31274 , n31266 , n31273 );
nor ( n31275 , n31265 , n31274 );
not ( n31276 , n31275 );
not ( n31277 , n31276 );
and ( n31278 , n31237 , n31277 );
and ( n31279 , n31236 , n31276 );
nor ( n31280 , n31278 , n31279 );
not ( n31281 , n31280 );
buf ( n31282 , RI173f50b0_1561);
not ( n31283 , n31282 );
buf ( n209045 , RI173e67b8_1632);
not ( n31285 , n209045 );
not ( n209047 , RI1739d780_1988);
not ( n31287 , n209047 );
or ( n31288 , n31285 , n31287 );
not ( n31289 , RI173e67b8_1632);
buf ( n31290 , RI1739d780_1988);
nand ( n31291 , n31289 , n31290 );
nand ( n31292 , n31288 , n31291 );
buf ( n31293 , RI1745e290_1277);
and ( n31294 , n31292 , n31293 );
not ( n31295 , n31292 );
not ( n31296 , RI1745e290_1277);
and ( n31297 , n31295 , n31296 );
nor ( n31298 , n31294 , n31297 );
buf ( n31299 , RI19a84ba8_2761);
nand ( n209061 , n25803 , n31299 );
buf ( n31301 , RI17507100_744);
and ( n209063 , n209061 , n31301 );
not ( n31303 , n209061 );
not ( n31304 , RI17507100_744);
and ( n31305 , n31303 , n31304 );
nor ( n31306 , n209063 , n31305 );
xor ( n31307 , n31298 , n31306 );
buf ( n31308 , RI19aa38c8_2541);
nand ( n31309 , n25491 , n31308 );
buf ( n31310 , RI17482aa0_1099);
and ( n31311 , n31309 , n31310 );
not ( n31312 , n31309 );
not ( n31313 , RI17482aa0_1099);
and ( n31314 , n31312 , n31313 );
nor ( n31315 , n31311 , n31314 );
not ( n31316 , n31315 );
xor ( n31317 , n31307 , n31316 );
not ( n31318 , n31317 );
or ( n31319 , n31283 , n31318 );
not ( n31320 , n31282 );
xor ( n31321 , n31298 , n31315 );
not ( n31322 , n31306 );
xnor ( n31323 , n31321 , n31322 );
nand ( n31324 , n31320 , n31323 );
nand ( n31325 , n31319 , n31324 );
buf ( n31326 , RI173f46d8_1564);
buf ( n31327 , RI17403cf0_1489);
not ( n31328 , n31327 );
not ( n31329 , RI173bb000_1844);
not ( n31330 , n31329 );
or ( n31331 , n31328 , n31330 );
not ( n31332 , RI17403cf0_1489);
buf ( n31333 , RI173bb000_1844);
nand ( n31334 , n31332 , n31333 );
nand ( n31335 , n31331 , n31334 );
xor ( n31336 , n31326 , n31335 );
buf ( n31337 , RI17535258_601);
not ( n31338 , RI1749ffd8_956);
xor ( n31339 , n31337 , n31338 );
buf ( n31340 , RI19ab7a58_2397);
nand ( n31341 , n25879 , n31340 );
xnor ( n31342 , n31339 , n31341 );
xnor ( n31343 , n31336 , n31342 );
not ( n31344 , n31343 );
and ( n31345 , n31325 , n31344 );
not ( n31346 , n31325 );
and ( n31347 , n31346 , n31343 );
nor ( n31348 , n31345 , n31347 );
not ( n31349 , n31348 );
not ( n31350 , n31349 );
buf ( n31351 , RI173e22d0_1653);
not ( n31352 , n31351 );
buf ( n209114 , RI173f3670_1569);
not ( n31354 , n209114 );
not ( n31355 , RI173aa980_1924);
not ( n31356 , n31355 );
or ( n31357 , n31354 , n31356 );
not ( n209119 , RI173f3670_1569);
buf ( n31359 , RI173aa980_1924);
nand ( n209121 , n209119 , n31359 );
nand ( n31361 , n31357 , n209121 );
not ( n31362 , RI174cfd50_764);
and ( n31363 , n31361 , n31362 );
not ( n31364 , n31361 );
buf ( n31365 , RI174cfd50_764);
and ( n31366 , n31364 , n31365 );
nor ( n31367 , n31363 , n31366 );
buf ( n31368 , RI19a23c18_2790);
nand ( n31369 , n29151 , n31368 );
buf ( n31370 , RI1751bb00_680);
and ( n31371 , n31369 , n31370 );
not ( n31372 , n31369 );
not ( n31373 , RI1751bb00_680);
and ( n31374 , n31372 , n31373 );
nor ( n31375 , n31371 , n31374 );
xor ( n31376 , n31367 , n31375 );
buf ( n31377 , RI19aaf268_2460);
nand ( n31378 , n26463 , n31377 );
buf ( n31379 , RI1748fca0_1035);
and ( n31380 , n31378 , n31379 );
not ( n31381 , n31378 );
not ( n31382 , RI1748fca0_1035);
and ( n31383 , n31381 , n31382 );
nor ( n209145 , n31380 , n31383 );
xnor ( n209146 , n31376 , n209145 );
not ( n31386 , n209146 );
not ( n31387 , n31386 );
or ( n31388 , n31352 , n31387 );
not ( n31389 , n209146 );
or ( n31390 , n31389 , n31351 );
nand ( n31391 , n31388 , n31390 );
buf ( n209153 , RI173c7eb8_1781);
not ( n31393 , n209153 );
not ( n31394 , RI1733e938_2136);
not ( n31395 , n31394 );
or ( n31396 , n31393 , n31395 );
not ( n31397 , RI173c7eb8_1781);
buf ( n31398 , RI1733e938_2136);
nand ( n31399 , n31397 , n31398 );
nand ( n31400 , n31396 , n31399 );
not ( n31401 , RI17410ba8_1426);
and ( n31402 , n31400 , n31401 );
not ( n31403 , n31400 );
buf ( n31404 , RI17410ba8_1426);
and ( n31405 , n31403 , n31404 );
nor ( n31406 , n31402 , n31405 );
buf ( n31407 , RI19a91808_2672);
nand ( n31408 , n25803 , n31407 );
not ( n31409 , RI17464500_1247);
and ( n31410 , n31408 , n31409 );
not ( n31411 , n31408 );
buf ( n31412 , RI17464500_1247);
and ( n31413 , n31411 , n31412 );
nor ( n31414 , n31410 , n31413 );
xor ( n209176 , n31406 , n31414 );
buf ( n31416 , RI19ac1a30_2317);
nand ( n31417 , n25416 , n31416 );
not ( n31418 , RI174ad1d8_892);
and ( n31419 , n31417 , n31418 );
not ( n31420 , n31417 );
buf ( n31421 , RI174ad1d8_892);
and ( n31422 , n31420 , n31421 );
nor ( n31423 , n31419 , n31422 );
xnor ( n31424 , n209176 , n31423 );
buf ( n31425 , n31424 );
and ( n31426 , n31391 , n31425 );
not ( n31427 , n31391 );
not ( n31428 , n31424 );
and ( n31429 , n31427 , n31428 );
nor ( n31430 , n31426 , n31429 );
not ( n31431 , n31430 );
nand ( n31432 , n31431 , n204511 );
not ( n31433 , n31432 );
or ( n31434 , n31350 , n31433 );
nand ( n31435 , n31431 , n204511 );
or ( n31436 , n31435 , n31349 );
nand ( n31437 , n31434 , n31436 );
not ( n31438 , n31437 );
not ( n31439 , n31438 );
buf ( n31440 , RI173e0f20_1659);
not ( n31441 , n31440 );
not ( n31442 , RI17398230_2014);
not ( n31443 , n31442 );
or ( n31444 , n31441 , n31443 );
not ( n31445 , RI173e0f20_1659);
buf ( n209207 , RI17398230_2014);
nand ( n31447 , n31445 , n209207 );
nand ( n209209 , n31444 , n31447 );
not ( n31449 , RI17458d40_1303);
and ( n31450 , n209209 , n31449 );
not ( n31451 , n209209 );
buf ( n31452 , RI17458d40_1303);
and ( n31453 , n31451 , n31452 );
nor ( n31454 , n31450 , n31453 );
buf ( n31455 , RI19ac3d58_2300);
nand ( n209217 , n25583 , n31455 );
buf ( n31457 , RI174cde60_770);
and ( n31458 , n209217 , n31457 );
not ( n31459 , n209217 );
not ( n31460 , RI174cde60_770);
and ( n31461 , n31459 , n31460 );
nor ( n31462 , n31458 , n31461 );
xor ( n31463 , n31454 , n31462 );
buf ( n31464 , RI19a93ba8_2656);
nand ( n31465 , n205020 , n31464 );
buf ( n31466 , RI1747d550_1125);
and ( n209228 , n31465 , n31466 );
not ( n31468 , n31465 );
not ( n31469 , RI1747d550_1125);
and ( n31470 , n31468 , n31469 );
nor ( n31471 , n209228 , n31470 );
xnor ( n31472 , n31463 , n31471 );
not ( n31473 , n31472 );
not ( n31474 , n31473 );
buf ( n31475 , RI174a09b0_953);
not ( n31476 , n31475 );
and ( n31477 , n31474 , n31476 );
and ( n31478 , n31473 , n31475 );
nor ( n31479 , n31477 , n31478 );
buf ( n31480 , RI173fe7a0_1515);
not ( n209242 , n31480 );
not ( n31482 , RI173b5768_1871);
not ( n31483 , n31482 );
or ( n31484 , n209242 , n31483 );
not ( n31485 , RI173fe7a0_1515);
buf ( n31486 , RI173b5768_1871);
nand ( n31487 , n31485 , n31486 );
nand ( n31488 , n31484 , n31487 );
buf ( n31489 , RI173bddf0_1830);
and ( n209251 , n31488 , n31489 );
not ( n31491 , n31488 );
not ( n31492 , RI173bddf0_1830);
and ( n31493 , n31491 , n31492 );
nor ( n31494 , n209251 , n31493 );
buf ( n31495 , RI19a88be0_2733);
nand ( n31496 , n25376 , n31495 );
not ( n31497 , RI1752cc48_627);
and ( n31498 , n31496 , n31497 );
not ( n31499 , n31496 );
buf ( n31500 , RI1752cc48_627);
and ( n31501 , n31499 , n31500 );
nor ( n31502 , n31498 , n31501 );
not ( n31503 , n31502 );
xor ( n31504 , n31494 , n31503 );
buf ( n31505 , RI19aa7a68_2512);
nand ( n31506 , n28997 , n31505 );
buf ( n31507 , RI1749aa88_982);
and ( n31508 , n31506 , n31507 );
not ( n209270 , n31506 );
not ( n31510 , RI1749aa88_982);
and ( n31511 , n209270 , n31510 );
nor ( n31512 , n31508 , n31511 );
buf ( n31513 , n31512 );
xnor ( n31514 , n31504 , n31513 );
buf ( n31515 , n31514 );
and ( n31516 , n31479 , n31515 );
not ( n31517 , n31479 );
not ( n31518 , n31512 );
not ( n209280 , n31502 );
or ( n31520 , n31518 , n209280 );
or ( n209282 , n31512 , n31502 );
nand ( n31522 , n31520 , n209282 );
and ( n31523 , n31522 , n31494 );
not ( n31524 , n31522 );
not ( n31525 , n31494 );
and ( n31526 , n31524 , n31525 );
nor ( n31527 , n31523 , n31526 );
buf ( n31528 , n31527 );
and ( n31529 , n31517 , n31528 );
nor ( n31530 , n31516 , n31529 );
not ( n31531 , n31530 );
nand ( n31532 , n31531 , n204263 );
and ( n31533 , n31532 , n25601 );
not ( n31534 , n31532 );
and ( n31535 , n31534 , n25600 );
nor ( n31536 , n31533 , n31535 );
not ( n31537 , n31536 );
not ( n31538 , n31537 );
or ( n31539 , n31439 , n31538 );
nand ( n31540 , n31437 , n31536 );
nand ( n209302 , n31539 , n31540 );
not ( n31542 , n209302 );
or ( n31543 , n31281 , n31542 );
or ( n31544 , n209302 , n31280 );
nand ( n31545 , n31543 , n31544 );
not ( n31546 , n31545 );
or ( n31547 , n31224 , n31546 );
not ( n31548 , n31545 );
not ( n31549 , n31223 );
nand ( n31550 , n31548 , n31549 );
nand ( n209312 , n31547 , n31550 );
buf ( n31552 , n209312 );
and ( n31553 , n30970 , n31552 );
not ( n31554 , n30970 );
not ( n31555 , n31545 );
not ( n31556 , n31555 );
not ( n31557 , n31549 );
and ( n31558 , n31556 , n31557 );
and ( n31559 , n31555 , n31549 );
nor ( n31560 , n31558 , n31559 );
buf ( n31561 , n31560 );
and ( n31562 , n31554 , n31561 );
nor ( n31563 , n31553 , n31562 );
not ( n31564 , n31563 );
nor ( n31565 , n29968 , n31564 );
nand ( n31566 , n205651 , n31565 );
not ( n31567 , n31563 );
not ( n31568 , n27880 );
not ( n31569 , n31568 );
or ( n31570 , n31567 , n31569 );
buf ( n31571 , n27886 );
buf ( n31572 , n31571 );
nor ( n31573 , n207728 , n31572 );
nand ( n209335 , n31570 , n31573 );
and ( n31575 , n27882 , n27883 );
buf ( n31576 , n31575 );
buf ( n31577 , n31576 );
nand ( n31578 , n31577 , n28076 );
nand ( n31579 , n31566 , n209335 , n31578 );
buf ( n31580 , n31579 );
not ( n31581 , n205098 );
not ( n31582 , RI173ac708_1915);
not ( n31583 , n31582 );
or ( n31584 , n31581 , n31583 );
not ( n31585 , RI173f53f8_1560);
buf ( n209347 , RI173ac708_1915);
nand ( n31587 , n31585 , n209347 );
nand ( n209349 , n31584 , n31587 );
not ( n31589 , RI1751d4c8_675);
and ( n31590 , n209349 , n31589 );
not ( n31591 , n209349 );
buf ( n31592 , RI1751d4c8_675);
and ( n31593 , n31591 , n31592 );
nor ( n31594 , n31590 , n31593 );
buf ( n31595 , RI19ac36c8_2303);
nand ( n31596 , n25803 , n31595 );
buf ( n31597 , RI1751e968_671);
and ( n31598 , n31596 , n31597 );
not ( n31599 , n31596 );
not ( n31600 , RI1751e968_671);
and ( n31601 , n31599 , n31600 );
nor ( n209363 , n31598 , n31601 );
xor ( n31603 , n31594 , n209363 );
buf ( n209365 , RI19aadfa8_2468);
nand ( n31605 , n204572 , n209365 );
buf ( n209367 , RI17491a28_1026);
and ( n31607 , n31605 , n209367 );
not ( n31608 , n31605 );
not ( n31609 , RI17491a28_1026);
and ( n31610 , n31608 , n31609 );
nor ( n31611 , n31607 , n31610 );
not ( n31612 , n31611 );
xor ( n31613 , n31603 , n31612 );
xor ( n31614 , n31293 , n31613 );
xnor ( n31615 , n31614 , n28121 );
buf ( n31616 , RI173e2ff0_1649);
not ( n31617 , n31616 );
not ( n31618 , RI1739a300_2004);
not ( n31619 , n31618 );
or ( n31620 , n31617 , n31619 );
not ( n31621 , RI173e2ff0_1649);
buf ( n31622 , RI1739a300_2004);
nand ( n31623 , n31621 , n31622 );
nand ( n209385 , n31620 , n31623 );
buf ( n31625 , RI1745ae10_1293);
and ( n31626 , n209385 , n31625 );
not ( n209388 , n209385 );
not ( n31628 , RI1745ae10_1293);
and ( n209390 , n209388 , n31628 );
nor ( n31630 , n31626 , n209390 );
buf ( n31631 , RI19aa62f8_2521);
nand ( n31632 , n25364 , n31631 );
buf ( n31633 , RI1747f620_1115);
xor ( n31634 , n31632 , n31633 );
xor ( n31635 , n31630 , n31634 );
xor ( n31636 , n31635 , n26067 );
buf ( n31637 , n31636 );
not ( n31638 , n31637 );
not ( n31639 , n205355 );
buf ( n31640 , RI173c5aa0_1792);
not ( n31641 , n31640 );
not ( n31642 , RI1733c520_2147);
not ( n31643 , n31642 );
or ( n31644 , n31641 , n31643 );
not ( n31645 , RI173c5aa0_1792);
buf ( n31646 , RI1733c520_2147);
nand ( n31647 , n31645 , n31646 );
nand ( n31648 , n31644 , n31647 );
not ( n31649 , RI1740e790_1437);
and ( n31650 , n31648 , n31649 );
not ( n31651 , n31648 );
buf ( n31652 , RI1740e790_1437);
and ( n31653 , n31651 , n31652 );
nor ( n31654 , n31650 , n31653 );
buf ( n31655 , RI19a92708_2665);
nand ( n31656 , n25751 , n31655 );
buf ( n31657 , RI174620e8_1258);
and ( n31658 , n31656 , n31657 );
not ( n31659 , n31656 );
not ( n31660 , RI174620e8_1258);
and ( n31661 , n31659 , n31660 );
nor ( n31662 , n31658 , n31661 );
xor ( n31663 , n31654 , n31662 );
buf ( n31664 , RI19ac2a98_2309);
nand ( n31665 , n25583 , n31664 );
not ( n31666 , RI174aadc0_903);
and ( n31667 , n31665 , n31666 );
not ( n31668 , n31665 );
buf ( n31669 , RI174aadc0_903);
and ( n31670 , n31668 , n31669 );
nor ( n31671 , n31667 , n31670 );
xor ( n31672 , n31663 , n31671 );
not ( n31673 , n31672 );
not ( n209435 , n31673 );
or ( n31675 , n31639 , n209435 );
not ( n209437 , n31672 );
or ( n31677 , n209437 , n205355 );
nand ( n31678 , n31675 , n31677 );
not ( n31679 , n31678 );
or ( n31680 , n31638 , n31679 );
or ( n31681 , n31678 , n31637 );
nand ( n31682 , n31680 , n31681 );
not ( n31683 , n31682 );
nand ( n31684 , n31615 , n31683 );
not ( n31685 , n31684 );
buf ( n31686 , RI173d9900_1695);
not ( n31687 , n31686 );
not ( n31688 , RI17390c10_2050);
not ( n31689 , n31688 );
or ( n31690 , n31687 , n31689 );
not ( n31691 , RI173d9900_1695);
buf ( n31692 , RI17390c10_2050);
nand ( n31693 , n31691 , n31692 );
nand ( n31694 , n31690 , n31693 );
not ( n31695 , n31694 );
buf ( n31696 , RI19ac8510_2267);
nand ( n31697 , n25540 , n31696 );
buf ( n31698 , RI174c24c0_806);
and ( n31699 , n31697 , n31698 );
not ( n31700 , n31697 );
not ( n31701 , RI174c24c0_806);
and ( n31702 , n31700 , n31701 );
nor ( n31703 , n31699 , n31702 );
not ( n31704 , n31703 );
buf ( n209466 , RI19a98ae0_2621);
nand ( n31706 , n25851 , n209466 );
buf ( n209468 , RI17475be8_1162);
and ( n31708 , n31706 , n209468 );
not ( n31709 , n31706 );
not ( n31710 , RI17475be8_1162);
and ( n31711 , n31709 , n31710 );
nor ( n31712 , n31708 , n31711 );
not ( n31713 , n31712 );
not ( n31714 , n31713 );
or ( n31715 , n31704 , n31714 );
not ( n31716 , n31703 );
nand ( n31717 , n31712 , n31716 );
nand ( n31718 , n31715 , n31717 );
buf ( n31719 , RI174513d8_1340);
and ( n31720 , n31718 , n31719 );
not ( n31721 , n31718 );
not ( n31722 , RI174513d8_1340);
and ( n31723 , n31721 , n31722 );
nor ( n31724 , n31720 , n31723 );
and ( n31725 , n31695 , n31724 );
not ( n31726 , n31695 );
not ( n31727 , n31724 );
and ( n31728 , n31726 , n31727 );
nor ( n209490 , n31725 , n31728 );
not ( n31730 , n209490 );
not ( n31731 , n31730 );
buf ( n31732 , RI173413e0_2123);
xor ( n31733 , n204732 , n204739 );
xnor ( n31734 , n31733 , n204743 );
not ( n31735 , n31734 );
and ( n31736 , n31732 , n31735 );
not ( n31737 , n31732 );
and ( n31738 , n31737 , n31734 );
nor ( n31739 , n31736 , n31738 );
not ( n31740 , n31739 );
and ( n209502 , n31731 , n31740 );
and ( n31742 , n31730 , n31739 );
nor ( n209504 , n209502 , n31742 );
not ( n31744 , n209504 );
not ( n31745 , n31744 );
and ( n31746 , n31685 , n31745 );
and ( n31747 , n31684 , n31744 );
nor ( n31748 , n31746 , n31747 );
not ( n31749 , n31748 );
buf ( n31750 , RI17337318_2172);
not ( n31751 , RI1745a0f0_1297);
xor ( n31752 , n31750 , n31751 );
buf ( n31753 , RI174a5bb8_928);
not ( n31754 , n31753 );
buf ( n209516 , RI19ab4038_2423);
nand ( n31756 , n205019 , n209516 );
not ( n209518 , n31756 );
or ( n31758 , n31754 , n209518 );
nand ( n31759 , n29151 , n209516 );
or ( n31760 , n31759 , n31753 );
nand ( n31761 , n31758 , n31760 );
xnor ( n31762 , n31752 , n31761 );
not ( n31763 , n31762 );
not ( n31764 , n31763 );
buf ( n31765 , RI173c0898_1817);
not ( n31766 , n31765 );
not ( n209528 , RI17409588_1462);
not ( n31768 , n209528 );
or ( n31769 , n31766 , n31768 );
not ( n31770 , RI173c0898_1817);
buf ( n31771 , RI17409588_1462);
nand ( n31772 , n31770 , n31771 );
nand ( n31773 , n31769 , n31772 );
not ( n31774 , n31773 );
and ( n31775 , n31764 , n31774 );
and ( n31776 , n31763 , n31773 );
nor ( n31777 , n31775 , n31776 );
buf ( n31778 , n31777 );
not ( n31779 , n31778 );
not ( n31780 , n205187 );
not ( n31781 , n30220 );
or ( n31782 , n31780 , n31781 );
nand ( n31783 , n204390 , n205183 );
nand ( n31784 , n31782 , n31783 );
not ( n209546 , n31784 );
and ( n31786 , n31779 , n209546 );
and ( n209548 , n31778 , n31784 );
nor ( n31788 , n31786 , n209548 );
not ( n31789 , n31788 );
not ( n31790 , n29185 );
not ( n31791 , n207960 );
or ( n31792 , n31790 , n31791 );
not ( n31793 , n29185 );
nand ( n31794 , n31793 , n30205 );
nand ( n31795 , n31792 , n31794 );
buf ( n31796 , RI173f1258_1580);
not ( n31797 , n31796 );
not ( n31798 , RI173a8568_1935);
not ( n31799 , n31798 );
or ( n209561 , n31797 , n31799 );
not ( n31801 , RI173f1258_1580);
buf ( n31802 , RI173a8568_1935);
nand ( n31803 , n31801 , n31802 );
nand ( n31804 , n209561 , n31803 );
not ( n31805 , RI174b09a0_875);
and ( n31806 , n31804 , n31805 );
not ( n31807 , n31804 );
buf ( n31808 , RI174b09a0_875);
and ( n31809 , n31807 , n31808 );
nor ( n31810 , n31806 , n31809 );
buf ( n31811 , RI19a94df0_2648);
nand ( n31812 , n25583 , n31811 );
buf ( n31813 , RI17518248_691);
and ( n31814 , n31812 , n31813 );
not ( n31815 , n31812 );
not ( n31816 , RI17518248_691);
and ( n31817 , n31815 , n31816 );
nor ( n209579 , n31814 , n31817 );
xor ( n31819 , n31810 , n209579 );
buf ( n31820 , RI19ab01e0_2453);
nand ( n31821 , n205271 , n31820 );
buf ( n31822 , RI1748d540_1047);
and ( n31823 , n31821 , n31822 );
not ( n31824 , n31821 );
not ( n31825 , RI1748d540_1047);
and ( n31826 , n31824 , n31825 );
nor ( n31827 , n31823 , n31826 );
xnor ( n31828 , n31819 , n31827 );
not ( n31829 , n31828 );
and ( n31830 , n31795 , n31829 );
not ( n31831 , n31795 );
buf ( n31832 , n31828 );
and ( n31833 , n31831 , n31832 );
nor ( n31834 , n31830 , n31833 );
nand ( n31835 , n31789 , n31834 );
not ( n209597 , n25500 );
not ( n31837 , n209597 );
buf ( n31838 , RI173c5758_1793);
not ( n31839 , n31838 );
not ( n31840 , RI1733c1d8_2148);
not ( n31841 , n31840 );
or ( n31842 , n31839 , n31841 );
not ( n31843 , RI173c5758_1793);
nand ( n31844 , n31843 , n205330 );
nand ( n31845 , n31842 , n31844 );
buf ( n31846 , RI1740e448_1438);
and ( n31847 , n31845 , n31846 );
not ( n31848 , n31845 );
not ( n31849 , RI1740e448_1438);
and ( n31850 , n31848 , n31849 );
nor ( n31851 , n31847 , n31850 );
buf ( n31852 , RI19a92528_2666);
nand ( n31853 , n29435 , n31852 );
not ( n31854 , RI17461da0_1259);
and ( n31855 , n31853 , n31854 );
not ( n31856 , n31853 );
buf ( n31857 , RI17461da0_1259);
and ( n31858 , n31856 , n31857 );
nor ( n31859 , n31855 , n31858 );
xor ( n31860 , n31851 , n31859 );
buf ( n31861 , RI19ac2840_2310);
nand ( n31862 , n25712 , n31861 );
not ( n209624 , RI174aaa78_904);
and ( n31864 , n31862 , n209624 );
not ( n209626 , n31862 );
buf ( n31866 , RI174aaa78_904);
and ( n209628 , n209626 , n31866 );
nor ( n31868 , n31864 , n209628 );
xnor ( n31869 , n31860 , n31868 );
not ( n31870 , n31869 );
not ( n31871 , n31870 );
or ( n31872 , n31837 , n31871 );
or ( n31873 , n31870 , n209597 );
nand ( n31874 , n31872 , n31873 );
buf ( n31875 , RI173e2ca8_1650);
not ( n31876 , n31875 );
not ( n31877 , RI17399fb8_2005);
not ( n31878 , n31877 );
or ( n31879 , n31876 , n31878 );
not ( n31880 , RI173e2ca8_1650);
buf ( n31881 , RI17399fb8_2005);
nand ( n31882 , n31880 , n31881 );
nand ( n31883 , n31879 , n31882 );
buf ( n31884 , RI1745aac8_1294);
and ( n31885 , n31883 , n31884 );
not ( n31886 , n31883 );
not ( n31887 , RI1745aac8_1294);
and ( n31888 , n31886 , n31887 );
nor ( n31889 , n31885 , n31888 );
buf ( n31890 , RI19aa6190_2522);
nand ( n31891 , n29151 , n31890 );
not ( n31892 , RI1747f2d8_1116);
and ( n31893 , n31891 , n31892 );
not ( n31894 , n31891 );
buf ( n31895 , RI1747f2d8_1116);
and ( n31896 , n31894 , n31895 );
nor ( n31897 , n31893 , n31896 );
xor ( n31898 , n31889 , n31897 );
xnor ( n31899 , n31898 , n30717 );
buf ( n31900 , n31899 );
and ( n209662 , n31874 , n31900 );
not ( n31902 , n31874 );
not ( n31903 , n31897 );
xor ( n31904 , n31889 , n31903 );
xnor ( n31905 , n31904 , n30717 );
not ( n31906 , n31905 );
not ( n31907 , n31906 );
and ( n31908 , n31902 , n31907 );
nor ( n31909 , n209662 , n31908 );
buf ( n31910 , n31909 );
and ( n31911 , n31835 , n31910 );
not ( n209673 , n31835 );
not ( n31913 , n31910 );
and ( n209675 , n209673 , n31913 );
nor ( n31915 , n31911 , n209675 );
not ( n31916 , n31915 );
not ( n31917 , n31916 );
nand ( n31918 , n209504 , n31682 );
buf ( n31919 , RI17336940_2175);
not ( n31920 , n31919 );
not ( n31921 , n204347 );
or ( n31922 , n31920 , n31921 );
not ( n31923 , n31919 );
not ( n31924 , n204326 );
xor ( n31925 , n31924 , n204344 );
xnor ( n31926 , n31925 , n204334 );
nand ( n31927 , n31923 , n31926 );
nand ( n31928 , n31922 , n31927 );
not ( n209690 , n25550 );
and ( n209691 , n31928 , n209690 );
not ( n31931 , n31928 );
buf ( n31932 , n25553 );
and ( n31933 , n31931 , n31932 );
nor ( n31934 , n209691 , n31933 );
and ( n31935 , n31918 , n31934 );
not ( n31936 , n31918 );
not ( n31937 , n31934 );
and ( n31938 , n31936 , n31937 );
nor ( n31939 , n31935 , n31938 );
not ( n31940 , n31939 );
not ( n31941 , n31940 );
or ( n209703 , n31917 , n31941 );
nand ( n31943 , n31939 , n31915 );
nand ( n209705 , n209703 , n31943 );
buf ( n31945 , RI173c43a8_1799);
xor ( n31946 , n31945 , n28044 );
xnor ( n31947 , n31946 , n205230 );
not ( n31948 , n31947 );
not ( n31949 , n25896 );
not ( n31950 , RI173c4a38_1797);
buf ( n31951 , RI173ff178_1512);
not ( n31952 , n31951 );
not ( n31953 , RI173b6140_1868);
not ( n31954 , n31953 );
or ( n31955 , n31952 , n31954 );
not ( n31956 , RI173ff178_1512);
buf ( n31957 , RI173b6140_1868);
nand ( n31958 , n31956 , n31957 );
nand ( n31959 , n31955 , n31958 );
xor ( n31960 , n31950 , n31959 );
buf ( n209722 , RI1752dbc0_624);
buf ( n31962 , RI1749b460_979);
xor ( n209724 , n209722 , n31962 );
buf ( n31964 , RI19ab96f0_2385);
nand ( n31965 , n205019 , n31964 );
xnor ( n31966 , n209724 , n31965 );
xor ( n31967 , n31960 , n31966 );
not ( n31968 , n31967 );
or ( n31969 , n31949 , n31968 );
buf ( n31970 , RI173c4a38_1797);
xor ( n31971 , n31970 , n31959 );
xor ( n209733 , n31971 , n31966 );
nand ( n31973 , n209733 , n25892 );
nand ( n209735 , n31969 , n31973 );
not ( n31975 , n209735 );
not ( n31976 , n206978 );
not ( n31977 , RI1738ace8_2079);
not ( n31978 , n31977 );
or ( n31979 , n31976 , n31978 );
not ( n31980 , RI173d39d8_1724);
buf ( n31981 , RI1738ace8_2079);
nand ( n209743 , n31980 , n31981 );
nand ( n31983 , n31979 , n209743 );
and ( n31984 , n31983 , n31225 );
not ( n31985 , n31983 );
not ( n31986 , RI1744b4b0_1369);
and ( n31987 , n31985 , n31986 );
nor ( n31988 , n31984 , n31987 );
buf ( n31989 , RI19acb4e0_2245);
nand ( n31990 , n25491 , n31989 );
buf ( n31991 , RI174b8a10_836);
and ( n31992 , n31990 , n31991 );
not ( n31993 , n31990 );
not ( n31994 , RI174b8a10_836);
and ( n31995 , n31993 , n31994 );
nor ( n31996 , n31992 , n31995 );
xor ( n31997 , n31988 , n31996 );
buf ( n31998 , RI19a9c1b8_2597);
nand ( n31999 , n25479 , n31998 );
buf ( n32000 , RI1746fcc0_1191);
and ( n32001 , n31999 , n32000 );
not ( n32002 , n31999 );
not ( n32003 , RI1746fcc0_1191);
and ( n32004 , n32002 , n32003 );
nor ( n32005 , n32001 , n32004 );
xnor ( n32006 , n31997 , n32005 );
buf ( n32007 , n32006 );
not ( n32008 , n32007 );
and ( n32009 , n31975 , n32008 );
not ( n32010 , n32006 );
not ( n32011 , n32010 );
and ( n32012 , n209735 , n32011 );
nor ( n32013 , n32009 , n32012 );
not ( n32014 , n32013 );
nand ( n32015 , n31948 , n32014 );
not ( n32016 , n32015 );
buf ( n32017 , n205017 );
not ( n32018 , n208904 );
not ( n32019 , RI1739c3d0_1994);
not ( n32020 , n32019 );
or ( n32021 , n32018 , n32020 );
not ( n32022 , RI173e5408_1638);
buf ( n32023 , RI1739c3d0_1994);
nand ( n209785 , n32022 , n32023 );
nand ( n32025 , n32021 , n209785 );
not ( n32026 , RI1745cee0_1283);
and ( n32027 , n32025 , n32026 );
not ( n32028 , n32025 );
buf ( n32029 , RI1745cee0_1283);
and ( n32030 , n32028 , n32029 );
nor ( n32031 , n32027 , n32030 );
buf ( n32032 , RI19a864f8_2750);
nand ( n32033 , n25479 , n32032 );
not ( n32034 , RI17503398_750);
and ( n209796 , n32033 , n32034 );
not ( n32036 , n32033 );
buf ( n209798 , RI17503398_750);
and ( n32038 , n32036 , n209798 );
nor ( n32039 , n209796 , n32038 );
xor ( n32040 , n32031 , n32039 );
buf ( n32041 , RI19aa5218_2529);
nand ( n32042 , n25451 , n32041 );
buf ( n32043 , RI174816f0_1105);
and ( n32044 , n32042 , n32043 );
not ( n32045 , n32042 );
not ( n32046 , RI174816f0_1105);
and ( n32047 , n32045 , n32046 );
nor ( n32048 , n32044 , n32047 );
xor ( n32049 , n32040 , n32048 );
buf ( n32050 , n32049 );
and ( n32051 , n32017 , n32050 );
not ( n32052 , n32017 );
not ( n32053 , n32049 );
and ( n32054 , n32052 , n32053 );
nor ( n32055 , n32051 , n32054 );
not ( n32056 , n32055 );
not ( n32057 , n32056 );
not ( n32058 , RI17402940_1495);
buf ( n32059 , RI173b9c50_1850);
and ( n32060 , n32058 , n32059 );
not ( n32061 , n32058 );
not ( n32062 , RI173b9c50_1850);
and ( n32063 , n32061 , n32062 );
nor ( n32064 , n32060 , n32063 );
not ( n32065 , n32064 );
buf ( n32066 , RI17533368_607);
not ( n32067 , RI173e6e48_1630);
xor ( n32068 , n32066 , n32067 );
buf ( n32069 , RI19ab9498_2386);
nand ( n32070 , n28238 , n32069 );
not ( n32071 , RI1749ec28_962);
and ( n32072 , n32070 , n32071 );
not ( n32073 , n32070 );
buf ( n32074 , RI1749ec28_962);
and ( n32075 , n32073 , n32074 );
nor ( n32076 , n32072 , n32075 );
xnor ( n32077 , n32068 , n32076 );
not ( n32078 , n32077 );
or ( n32079 , n32065 , n32078 );
or ( n32080 , n32077 , n32064 );
nand ( n32081 , n32079 , n32080 );
buf ( n32082 , n32081 );
not ( n209844 , n32082 );
not ( n32084 , n209844 );
or ( n209846 , n32057 , n32084 );
nand ( n32086 , n32082 , n32055 );
nand ( n32087 , n209846 , n32086 );
not ( n32088 , n32087 );
and ( n32089 , n32016 , n32088 );
and ( n32090 , n32015 , n32087 );
nor ( n32091 , n32089 , n32090 );
not ( n32092 , n32091 );
and ( n32093 , n209705 , n32092 );
not ( n32094 , n209705 );
and ( n32095 , n32094 , n32091 );
nor ( n32096 , n32093 , n32095 );
not ( n32097 , n32096 );
buf ( n32098 , RI19a838e8_2769);
nand ( n32099 , n204512 , n32098 );
buf ( n32100 , RI1750a490_734);
and ( n32101 , n32099 , n32100 );
not ( n32102 , n32099 );
not ( n32103 , RI1750a490_734);
and ( n32104 , n32102 , n32103 );
nor ( n32105 , n32101 , n32104 );
not ( n32106 , n32105 );
buf ( n32107 , RI173d9f90_1693);
not ( n32108 , n32107 );
not ( n32109 , RI173912a0_2048);
not ( n32110 , n32109 );
or ( n32111 , n32108 , n32110 );
not ( n209873 , RI173d9f90_1693);
buf ( n32113 , RI173912a0_2048);
nand ( n209875 , n209873 , n32113 );
nand ( n32115 , n32111 , n209875 );
not ( n32116 , RI17451a68_1338);
and ( n32117 , n32115 , n32116 );
not ( n32118 , n32115 );
buf ( n32119 , RI17451a68_1338);
and ( n32120 , n32118 , n32119 );
nor ( n32121 , n32117 , n32120 );
buf ( n32122 , RI19a98f90_2619);
nand ( n209884 , n26453 , n32122 );
buf ( n32124 , RI17476278_1160);
xor ( n209886 , n209884 , n32124 );
xor ( n32126 , n32121 , n209886 );
buf ( n32127 , RI19ac89c0_2265);
nand ( n32128 , n26162 , n32127 );
not ( n32129 , RI174c2f10_804);
and ( n32130 , n32128 , n32129 );
not ( n32131 , n32128 );
buf ( n32132 , RI174c2f10_804);
and ( n209894 , n32131 , n32132 );
nor ( n32134 , n32130 , n209894 );
xnor ( n32135 , n32126 , n32134 );
buf ( n32136 , n32135 );
and ( n32137 , n32106 , n32136 );
not ( n32138 , n32106 );
not ( n32139 , n32135 );
and ( n32140 , n32138 , n32139 );
or ( n32141 , n32137 , n32140 );
buf ( n32142 , RI173f74c8_1550);
not ( n32143 , n32142 );
not ( n32144 , RI173ae7d8_1905);
not ( n32145 , n32144 );
or ( n32146 , n32143 , n32145 );
not ( n32147 , RI173f74c8_1550);
buf ( n32148 , RI173ae7d8_1905);
nand ( n32149 , n32147 , n32148 );
nand ( n32150 , n32146 , n32149 );
buf ( n32151 , RI17336c88_2174);
and ( n32152 , n32150 , n32151 );
not ( n32153 , n32150 );
not ( n32154 , RI17336c88_2174);
and ( n32155 , n32153 , n32154 );
nor ( n32156 , n32152 , n32155 );
buf ( n32157 , RI19aacdd8_2476);
nand ( n32158 , n30640 , n32157 );
not ( n32159 , RI17493af8_1016);
and ( n209921 , n32158 , n32159 );
not ( n32161 , n32158 );
buf ( n32162 , RI17493af8_1016);
and ( n32163 , n32161 , n32162 );
nor ( n32164 , n209921 , n32163 );
xor ( n32165 , n32156 , n32164 );
buf ( n32166 , RI19ab9df8_2381);
nand ( n32167 , n25851 , n32166 );
not ( n32168 , RI17521cf8_661);
and ( n32169 , n32167 , n32168 );
not ( n32170 , n32167 );
buf ( n32171 , RI17521cf8_661);
and ( n32172 , n32170 , n32171 );
nor ( n32173 , n32169 , n32172 );
xnor ( n32174 , n32165 , n32173 );
buf ( n32175 , n32174 );
not ( n32176 , n32175 );
buf ( n32177 , n32176 );
and ( n32178 , n32141 , n32177 );
not ( n32179 , n32141 );
not ( n32180 , n32174 );
not ( n209942 , n32180 );
not ( n32182 , n209942 );
not ( n32183 , n32182 );
and ( n32184 , n32179 , n32183 );
nor ( n32185 , n32178 , n32184 );
not ( n32186 , n32185 );
not ( n32187 , RI173b2978_1885);
buf ( n32188 , RI17485548_1086);
buf ( n32189 , RI19a9e8a0_2580);
nand ( n209951 , n25490 , n32189 );
buf ( n32191 , RI17489058_1068);
and ( n209953 , n209951 , n32191 );
not ( n32193 , n209951 );
not ( n32194 , RI17489058_1068);
and ( n32195 , n32193 , n32194 );
nor ( n32196 , n209953 , n32195 );
xor ( n32197 , n32188 , n32196 );
buf ( n32198 , RI19acd358_2230);
nand ( n32199 , n25656 , n32198 );
not ( n32200 , RI175110d8_713);
and ( n32201 , n32199 , n32200 );
not ( n32202 , n32199 );
buf ( n32203 , RI175110d8_713);
and ( n209965 , n32202 , n32203 );
nor ( n32205 , n32201 , n209965 );
xnor ( n32206 , n32197 , n32205 );
not ( n32207 , n32206 );
not ( n32208 , RI173ecd70_1601);
buf ( n32209 , RI173a4080_1956);
and ( n32210 , n32208 , n32209 );
not ( n32211 , n32208 );
not ( n32212 , RI173a4080_1956);
and ( n32213 , n32211 , n32212 );
nor ( n32214 , n32210 , n32213 );
not ( n32215 , n32214 );
and ( n32216 , n32207 , n32215 );
and ( n32217 , n32206 , n32214 );
nor ( n32218 , n32216 , n32217 );
buf ( n32219 , n32218 );
xor ( n32220 , n32187 , n32219 );
buf ( n32221 , RI17477970_1153);
not ( n32222 , RI1740a2a8_1458);
buf ( n32223 , RI173c15b8_1813);
nand ( n32224 , n32222 , n32223 );
not ( n32225 , RI173c15b8_1813);
buf ( n32226 , RI1740a2a8_1458);
nand ( n32227 , n32225 , n32226 );
and ( n32228 , n32224 , n32227 );
xor ( n32229 , n32221 , n32228 );
buf ( n32230 , RI17338038_2168);
buf ( n32231 , RI174a68d8_924);
xor ( n32232 , n32230 , n32231 );
buf ( n32233 , RI19ab2328_2438);
nand ( n32234 , n205271 , n32233 );
xnor ( n32235 , n32232 , n32234 );
xor ( n32236 , n32229 , n32235 );
and ( n32237 , n32220 , n32236 );
not ( n32238 , n32220 );
xor ( n210000 , n32221 , n32228 );
xnor ( n32240 , n210000 , n32235 );
buf ( n210002 , n32240 );
and ( n32242 , n32238 , n210002 );
nor ( n32243 , n32237 , n32242 );
buf ( n32244 , RI17406108_1478);
not ( n32245 , n32244 );
buf ( n32246 , RI173aeb20_1904);
not ( n32247 , n32246 );
not ( n32248 , RI173f7810_1549);
not ( n32249 , n32248 );
or ( n210011 , n32247 , n32249 );
not ( n32251 , RI173aeb20_1904);
buf ( n32252 , RI173f7810_1549);
nand ( n32253 , n32251 , n32252 );
nand ( n32254 , n210011 , n32253 );
not ( n32255 , RI173390a0_2163);
and ( n32256 , n32254 , n32255 );
not ( n32257 , n32254 );
buf ( n32258 , RI173390a0_2163);
and ( n32259 , n32257 , n32258 );
nor ( n32260 , n32256 , n32259 );
buf ( n32261 , RI19aad120_2475);
nand ( n32262 , n29890 , n32261 );
not ( n32263 , RI17493e40_1015);
and ( n32264 , n32262 , n32263 );
not ( n32265 , n32262 );
buf ( n32266 , RI17493e40_1015);
and ( n32267 , n32265 , n32266 );
nor ( n210029 , n32264 , n32267 );
xor ( n32269 , n32260 , n210029 );
buf ( n32270 , RI19abba90_2370);
nand ( n32271 , n29203 , n32270 );
buf ( n32272 , RI17522220_660);
and ( n32273 , n32271 , n32272 );
not ( n32274 , n32271 );
not ( n32275 , RI17522220_660);
and ( n32276 , n32274 , n32275 );
nor ( n32277 , n32273 , n32276 );
xor ( n32278 , n32269 , n32277 );
not ( n32279 , n32278 );
buf ( n32280 , n32279 );
not ( n32281 , n32280 );
or ( n32282 , n32245 , n32281 );
buf ( n210044 , n32278 );
not ( n32284 , n210044 );
not ( n210046 , n32284 );
not ( n32286 , RI17406108_1478);
nand ( n32287 , n210046 , n32286 );
nand ( n32288 , n32282 , n32287 );
buf ( n32289 , RI173cc058_1761);
not ( n32290 , n32289 );
not ( n32291 , RI17342ad8_2116);
not ( n32292 , n32291 );
or ( n32293 , n32290 , n32292 );
not ( n32294 , RI173cc058_1761);
buf ( n32295 , RI17342ad8_2116);
nand ( n32296 , n32294 , n32295 );
nand ( n32297 , n32293 , n32296 );
buf ( n32298 , RI17415090_1405);
and ( n32299 , n32297 , n32298 );
not ( n32300 , n32297 );
not ( n32301 , RI17415090_1405);
and ( n32302 , n32300 , n32301 );
nor ( n32303 , n32299 , n32302 );
buf ( n32304 , RI19a8cd80_2705);
nand ( n32305 , n26463 , n32304 );
buf ( n32306 , RI174686a0_1227);
and ( n32307 , n32305 , n32306 );
not ( n32308 , n32305 );
not ( n32309 , RI174686a0_1227);
and ( n32310 , n32308 , n32309 );
nor ( n32311 , n32307 , n32310 );
xor ( n32312 , n32303 , n32311 );
buf ( n32313 , RI19abdf98_2350);
nand ( n32314 , n25405 , n32313 );
buf ( n210076 , RI174b1378_872);
and ( n32316 , n32314 , n210076 );
not ( n210078 , n32314 );
not ( n32318 , RI174b1378_872);
and ( n32319 , n210078 , n32318 );
nor ( n32320 , n32316 , n32319 );
xor ( n32321 , n32312 , n32320 );
not ( n32322 , n32321 );
buf ( n32323 , n32322 );
and ( n32324 , n32288 , n32323 );
not ( n32325 , n32288 );
buf ( n32326 , n32321 );
and ( n32327 , n32325 , n32326 );
nor ( n32328 , n32324 , n32327 );
not ( n32329 , n32328 );
nand ( n32330 , n32243 , n32329 );
not ( n32331 , n32330 );
or ( n32332 , n32186 , n32331 );
not ( n32333 , n32328 );
nand ( n32334 , n32333 , n32243 );
or ( n32335 , n32334 , n32185 );
nand ( n32336 , n32332 , n32335 );
not ( n32337 , n32336 );
buf ( n32338 , n206902 );
buf ( n32339 , RI19abb298_2373);
nand ( n32340 , n32338 , n32339 );
not ( n32341 , RI174b72a0_843);
and ( n32342 , n32340 , n32341 );
not ( n32343 , n32340 );
buf ( n32344 , RI174b72a0_843);
and ( n32345 , n32343 , n32344 );
nor ( n32346 , n32342 , n32345 );
not ( n32347 , n31473 );
xor ( n32348 , n32346 , n32347 );
not ( n32349 , RI173e46e8_1642);
not ( n32350 , RI1740c6c0_1447);
and ( n32351 , n32350 , n29375 );
not ( n32352 , n32350 );
and ( n32353 , n32352 , n29417 );
nor ( n32354 , n32351 , n32353 );
xor ( n32355 , n32349 , n32354 );
buf ( n32356 , RI1733a450_2157);
buf ( n210118 , RI174a8cf0_913);
xor ( n32358 , n32356 , n210118 );
buf ( n210120 , RI19ab1518_2444);
nand ( n32360 , n28902 , n210120 );
xnor ( n32361 , n32358 , n32360 );
xnor ( n32362 , n32355 , n32361 );
buf ( n32363 , n32362 );
xor ( n32364 , n32348 , n32363 );
not ( n32365 , n32364 );
not ( n32366 , n32365 );
buf ( n32367 , RI17391fc0_2044);
not ( n32368 , n32367 );
buf ( n32369 , RI173cc3a0_1760);
not ( n32370 , n32369 );
not ( n32371 , RI17342e20_2115);
not ( n32372 , n32371 );
or ( n32373 , n32370 , n32372 );
not ( n210135 , RI173cc3a0_1760);
buf ( n32375 , RI17342e20_2115);
nand ( n210137 , n210135 , n32375 );
nand ( n32377 , n32373 , n210137 );
buf ( n32378 , RI174153d8_1404);
and ( n32379 , n32377 , n32378 );
not ( n32380 , n32377 );
not ( n32381 , RI174153d8_1404);
and ( n32382 , n32380 , n32381 );
nor ( n32383 , n32379 , n32382 );
buf ( n32384 , RI19a8cfd8_2704);
nand ( n32385 , n28148 , n32384 );
buf ( n32386 , RI174689e8_1226);
and ( n32387 , n32385 , n32386 );
not ( n32388 , n32385 );
not ( n32389 , RI174689e8_1226);
and ( n32390 , n32388 , n32389 );
nor ( n32391 , n32387 , n32390 );
xor ( n32392 , n32383 , n32391 );
buf ( n210154 , RI19abe100_2349);
nand ( n32394 , n204926 , n210154 );
not ( n32395 , RI174b16c0_871);
and ( n32396 , n32394 , n32395 );
not ( n32397 , n32394 );
buf ( n32398 , RI174b16c0_871);
and ( n32399 , n32397 , n32398 );
nor ( n32400 , n32396 , n32399 );
xnor ( n32401 , n32392 , n32400 );
not ( n32402 , n32401 );
not ( n32403 , n32402 );
or ( n32404 , n32368 , n32403 );
buf ( n32405 , n32401 );
not ( n32406 , n32405 );
or ( n32407 , n32406 , n32367 );
nand ( n32408 , n32404 , n32407 );
buf ( n32409 , RI173a0f48_1971);
not ( n32410 , n32409 );
not ( n32411 , RI173e9c38_1616);
not ( n32412 , n32411 );
or ( n32413 , n32410 , n32412 );
not ( n32414 , RI173a0f48_1971);
buf ( n32415 , RI173e9c38_1616);
nand ( n32416 , n32414 , n32415 );
nand ( n210178 , n32413 , n32416 );
buf ( n32418 , RI174658b0_1241);
and ( n210180 , n210178 , n32418 );
not ( n32420 , n210178 );
not ( n32421 , RI174658b0_1241);
and ( n32422 , n32420 , n32421 );
nor ( n32423 , n210180 , n32422 );
buf ( n32424 , RI19acfd88_2212);
nand ( n32425 , n26058 , n32424 );
buf ( n32426 , RI1750c380_728);
and ( n32427 , n32425 , n32426 );
not ( n32428 , n32425 );
not ( n32429 , RI1750c380_728);
and ( n32430 , n32428 , n32429 );
nor ( n32431 , n32427 , n32430 );
xor ( n32432 , n32423 , n32431 );
buf ( n32433 , RI19aa0f10_2561);
nand ( n32434 , n25376 , n32433 );
not ( n32435 , RI17485f20_1083);
and ( n32436 , n32434 , n32435 );
not ( n32437 , n32434 );
buf ( n32438 , RI17485f20_1083);
and ( n32439 , n32437 , n32438 );
nor ( n32440 , n32436 , n32439 );
xnor ( n32441 , n32432 , n32440 );
buf ( n32442 , n32441 );
not ( n32443 , n32442 );
and ( n32444 , n32408 , n32443 );
not ( n32445 , n32408 );
and ( n32446 , n32445 , n32442 );
nor ( n32447 , n32444 , n32446 );
buf ( n32448 , RI173ea958_1612);
not ( n32449 , n32448 );
not ( n32450 , n28647 );
or ( n210212 , n32449 , n32450 );
or ( n32452 , n28647 , n32448 );
nand ( n210214 , n210212 , n32452 );
buf ( n32454 , n27848 );
and ( n32455 , n210214 , n32454 );
not ( n32456 , n210214 );
buf ( n32457 , n27842 );
and ( n32458 , n32456 , n32457 );
nor ( n32459 , n32455 , n32458 );
nand ( n32460 , n32447 , n32459 );
not ( n32461 , n32460 );
and ( n32462 , n32366 , n32461 );
and ( n32463 , n32365 , n32460 );
nor ( n32464 , n32462 , n32463 );
not ( n32465 , n32464 );
and ( n32466 , n32337 , n32465 );
and ( n32467 , n32336 , n32464 );
nor ( n32468 , n32466 , n32467 );
not ( n32469 , n32468 );
and ( n32470 , n32097 , n32469 );
and ( n32471 , n32468 , n32096 );
nor ( n32472 , n32470 , n32471 );
not ( n32473 , n32472 );
not ( n32474 , n32473 );
or ( n32475 , n31749 , n32474 );
or ( n32476 , n32473 , n31748 );
nand ( n32477 , n32475 , n32476 );
not ( n32478 , n32477 );
not ( n32479 , n29762 );
not ( n32480 , n29768 );
or ( n32481 , n32479 , n32480 );
or ( n32482 , n29768 , n29762 );
nand ( n32483 , n32481 , n32482 );
not ( n32484 , n32483 );
not ( n210246 , n25593 );
buf ( n210247 , RI173fa948_1534);
buf ( n32487 , n210247 );
not ( n210249 , n32487 );
and ( n210250 , n210246 , n210249 );
and ( n32490 , n25593 , n32487 );
nor ( n210252 , n210250 , n32490 );
not ( n210253 , n210252 );
and ( n32493 , n32484 , n210253 );
and ( n32494 , n29773 , n210252 );
nor ( n32495 , n32493 , n32494 );
not ( n32496 , n32495 );
not ( n32497 , n32496 );
not ( n32498 , n25761 );
buf ( n32499 , RI1744a100_1375);
not ( n32500 , n32499 );
and ( n210262 , n32498 , n32500 );
and ( n32502 , n25761 , n32499 );
nor ( n210264 , n210262 , n32502 );
and ( n32504 , n210264 , n25722 );
not ( n32505 , n210264 );
and ( n32506 , n32505 , n25772 );
nor ( n32507 , n32504 , n32506 );
not ( n32508 , n32507 );
buf ( n32509 , RI19a8e220_2696);
nand ( n32510 , n204572 , n32509 );
not ( n32511 , RI17466918_1236);
and ( n32512 , n32510 , n32511 );
not ( n32513 , n32510 );
buf ( n32514 , RI17466918_1236);
and ( n32515 , n32513 , n32514 );
nor ( n32516 , n32512 , n32515 );
buf ( n32517 , n32516 );
not ( n32518 , n32517 );
not ( n32519 , n30099 );
or ( n32520 , n32518 , n32519 );
not ( n32521 , n32517 );
buf ( n32522 , RI173fb668_1530);
xor ( n32523 , n32522 , n30091 );
xnor ( n32524 , n32523 , n30098 );
nand ( n32525 , n32521 , n32524 );
nand ( n32526 , n32520 , n32525 );
and ( n32527 , n32526 , n28722 );
not ( n32528 , n32526 );
and ( n32529 , n32528 , n28721 );
nor ( n32530 , n32527 , n32529 );
nand ( n32531 , n32508 , n32530 );
not ( n32532 , n32531 );
or ( n32533 , n32497 , n32532 );
not ( n32534 , n32507 );
nand ( n32535 , n32534 , n32530 );
or ( n32536 , n32535 , n32496 );
nand ( n32537 , n32533 , n32536 );
not ( n32538 , n32537 );
buf ( n32539 , RI173d8208_1702);
not ( n32540 , n32539 );
not ( n32541 , RI1738f518_2057);
not ( n32542 , n32541 );
or ( n32543 , n32540 , n32542 );
not ( n32544 , RI173d8208_1702);
buf ( n32545 , RI1738f518_2057);
nand ( n32546 , n32544 , n32545 );
nand ( n32547 , n32543 , n32546 );
not ( n32548 , n32547 );
buf ( n32549 , RI19ac9b90_2257);
nand ( n32550 , n25539 , n32549 );
buf ( n32551 , RI174c00a8_813);
and ( n32552 , n32550 , n32551 );
not ( n32553 , n32550 );
not ( n32554 , RI174c00a8_813);
and ( n32555 , n32553 , n32554 );
nor ( n32556 , n32552 , n32555 );
xor ( n32557 , n28467 , n32556 );
buf ( n32558 , RI19a9a3b8_2610);
nand ( n32559 , n29435 , n32558 );
buf ( n32560 , RI174744f0_1169);
and ( n32561 , n32559 , n32560 );
not ( n32562 , n32559 );
not ( n32563 , RI174744f0_1169);
and ( n32564 , n32562 , n32563 );
nor ( n32565 , n32561 , n32564 );
xnor ( n32566 , n32557 , n32565 );
not ( n32567 , n32566 );
not ( n32568 , n32567 );
or ( n32569 , n32548 , n32568 );
not ( n32570 , n32547 );
nand ( n32571 , n32566 , n32570 );
nand ( n32572 , n32569 , n32571 );
xor ( n32573 , n205109 , n32572 );
buf ( n32574 , RI173f5740_1559);
not ( n32575 , n32574 );
not ( n32576 , RI173aca50_1914);
not ( n32577 , n32576 );
or ( n32578 , n32575 , n32577 );
not ( n32579 , RI173f5740_1559);
buf ( n32580 , RI173aca50_1914);
nand ( n32581 , n32579 , n32580 );
nand ( n32582 , n32578 , n32581 );
not ( n32583 , RI17520d80_664);
and ( n32584 , n32582 , n32583 );
not ( n32585 , n32582 );
buf ( n32586 , RI17520d80_664);
and ( n32587 , n32585 , n32586 );
nor ( n32588 , n32584 , n32587 );
buf ( n32589 , RI19aae110_2467);
nand ( n32590 , n25751 , n32589 );
buf ( n32591 , RI17491d70_1025);
and ( n32592 , n32590 , n32591 );
not ( n32593 , n32590 );
not ( n32594 , RI17491d70_1025);
and ( n32595 , n32593 , n32594 );
nor ( n32596 , n32592 , n32595 );
xor ( n32597 , n32588 , n32596 );
buf ( n32598 , RI19ac4f28_2292);
nand ( n32599 , n26266 , n32598 );
buf ( n32600 , RI1751ee90_670);
and ( n32601 , n32599 , n32600 );
not ( n32602 , n32599 );
not ( n210364 , RI1751ee90_670);
and ( n32604 , n32602 , n210364 );
nor ( n210366 , n32601 , n32604 );
not ( n32606 , n210366 );
xnor ( n32607 , n32597 , n32606 );
buf ( n32608 , n32607 );
xor ( n32609 , n32573 , n32608 );
buf ( n32610 , RI19aa8bc0_2505);
nand ( n32611 , n204926 , n32610 );
not ( n32612 , RI174989b8_992);
and ( n32613 , n32611 , n32612 );
not ( n32614 , n32611 );
buf ( n32615 , RI174989b8_992);
and ( n32616 , n32614 , n32615 );
nor ( n32617 , n32613 , n32616 );
not ( n32618 , n32617 );
buf ( n32619 , RI173a50e8_1951);
not ( n32620 , n32619 );
not ( n32621 , RI173eddd8_1596);
not ( n32622 , n32621 );
or ( n32623 , n32620 , n32622 );
not ( n32624 , RI173a50e8_1951);
buf ( n32625 , RI173eddd8_1596);
nand ( n32626 , n32624 , n32625 );
nand ( n32627 , n32623 , n32626 );
buf ( n32628 , RI1748e8f0_1041);
and ( n32629 , n32627 , n32628 );
not ( n32630 , n32627 );
not ( n32631 , RI1748e8f0_1041);
and ( n32632 , n32630 , n32631 );
nor ( n32633 , n32629 , n32632 );
buf ( n32634 , RI19acdcb8_2226);
nand ( n32635 , n26242 , n32634 );
buf ( n32636 , RI17512fc8_707);
and ( n32637 , n32635 , n32636 );
not ( n32638 , n32635 );
not ( n32639 , RI17512fc8_707);
and ( n32640 , n32638 , n32639 );
nor ( n32641 , n32637 , n32640 );
xor ( n32642 , n32633 , n32641 );
buf ( n32643 , RI19a9f188_2576);
nand ( n32644 , n32338 , n32643 );
not ( n32645 , RI1748a0c0_1063);
and ( n32646 , n32644 , n32645 );
not ( n32647 , n32644 );
buf ( n32648 , RI1748a0c0_1063);
and ( n32649 , n32647 , n32648 );
nor ( n32650 , n32646 , n32649 );
xnor ( n32651 , n32642 , n32650 );
not ( n32652 , n32651 );
not ( n32653 , n32652 );
or ( n32654 , n32618 , n32653 );
buf ( n32655 , n32651 );
not ( n32656 , n32617 );
nand ( n32657 , n32655 , n32656 );
nand ( n32658 , n32654 , n32657 );
not ( n32659 , n32658 );
buf ( n32660 , RI17512578_709);
buf ( n32661 , RI1740afc8_1454);
not ( n32662 , n32661 );
not ( n32663 , RI173c22d8_1809);
not ( n32664 , n32663 );
or ( n32665 , n32662 , n32664 );
not ( n32666 , RI1740afc8_1454);
buf ( n32667 , RI173c22d8_1809);
nand ( n210429 , n32666 , n32667 );
nand ( n32669 , n32665 , n210429 );
xor ( n32670 , n32660 , n32669 );
buf ( n32671 , RI17338d58_2164);
not ( n32672 , n32671 );
buf ( n32673 , RI19ab2d78_2433);
nand ( n32674 , n204336 , n32673 );
buf ( n32675 , RI174a75f8_920);
and ( n32676 , n32674 , n32675 );
not ( n32677 , n32674 );
not ( n32678 , RI174a75f8_920);
and ( n32679 , n32677 , n32678 );
nor ( n32680 , n32676 , n32679 );
not ( n32681 , n32680 );
or ( n32682 , n32672 , n32681 );
or ( n32683 , n32680 , n32671 );
nand ( n32684 , n32682 , n32683 );
xnor ( n32685 , n32670 , n32684 );
not ( n32686 , n32685 );
and ( n32687 , n32659 , n32686 );
not ( n32688 , n32685 );
not ( n32689 , n32688 );
and ( n32690 , n32689 , n32658 );
nor ( n32691 , n32687 , n32690 );
not ( n32692 , n32691 );
nand ( n32693 , n32609 , n32692 );
not ( n32694 , n32693 );
not ( n32695 , n26069 );
buf ( n32696 , RI173c5de8_1791);
not ( n32697 , n32696 );
not ( n32698 , RI1733c868_2146);
not ( n32699 , n32698 );
or ( n32700 , n32697 , n32699 );
not ( n32701 , RI173c5de8_1791);
buf ( n32702 , RI1733c868_2146);
nand ( n32703 , n32701 , n32702 );
nand ( n32704 , n32700 , n32703 );
not ( n32705 , RI1740ead8_1436);
and ( n32706 , n32704 , n32705 );
not ( n32707 , n32704 );
buf ( n32708 , RI1740ead8_1436);
and ( n32709 , n32707 , n32708 );
nor ( n32710 , n32706 , n32709 );
buf ( n32711 , RI19ac2cf0_2308);
nand ( n32712 , n27946 , n32711 );
buf ( n32713 , RI174ab108_902);
and ( n32714 , n32712 , n32713 );
not ( n32715 , n32712 );
not ( n32716 , RI174ab108_902);
and ( n32717 , n32715 , n32716 );
nor ( n32718 , n32714 , n32717 );
xor ( n210480 , n32710 , n32718 );
buf ( n32720 , RI19a92960_2664);
nand ( n32721 , n25666 , n32720 );
buf ( n32722 , RI17462430_1257);
and ( n32723 , n32721 , n32722 );
not ( n32724 , n32721 );
not ( n32725 , RI17462430_1257);
and ( n32726 , n32724 , n32725 );
nor ( n32727 , n32723 , n32726 );
xnor ( n210489 , n210480 , n32727 );
not ( n32729 , n210489 );
not ( n32730 , n32729 );
or ( n32731 , n32695 , n32730 );
or ( n32732 , n32729 , n26069 );
nand ( n32733 , n32731 , n32732 );
buf ( n32734 , RI173e3338_1648);
not ( n32735 , n32734 );
not ( n32736 , RI1739a648_2003);
not ( n210498 , n32736 );
or ( n32738 , n32735 , n210498 );
not ( n32739 , RI173e3338_1648);
buf ( n32740 , RI1739a648_2003);
nand ( n32741 , n32739 , n32740 );
nand ( n32742 , n32738 , n32741 );
not ( n32743 , RI1745b158_1292);
and ( n32744 , n32742 , n32743 );
not ( n32745 , n32742 );
buf ( n32746 , RI1745b158_1292);
and ( n32747 , n32745 , n32746 );
nor ( n32748 , n32744 , n32747 );
buf ( n32749 , RI19a87920_2741);
nand ( n32750 , n30640 , n32749 );
buf ( n32751 , RI17500530_759);
and ( n32752 , n32750 , n32751 );
not ( n32753 , n32750 );
not ( n32754 , RI17500530_759);
and ( n32755 , n32753 , n32754 );
nor ( n32756 , n32752 , n32755 );
xor ( n32757 , n32748 , n32756 );
buf ( n32758 , RI19aa6640_2520);
nand ( n32759 , n25405 , n32758 );
not ( n32760 , RI1747f968_1114);
and ( n32761 , n32759 , n32760 );
not ( n32762 , n32759 );
buf ( n32763 , RI1747f968_1114);
and ( n32764 , n32762 , n32763 );
nor ( n32765 , n32761 , n32764 );
xnor ( n32766 , n32757 , n32765 );
not ( n32767 , n32766 );
buf ( n32768 , n32767 );
not ( n32769 , n32768 );
and ( n32770 , n32733 , n32769 );
not ( n32771 , n32733 );
not ( n210533 , n32756 );
not ( n32773 , n32765 );
or ( n32774 , n210533 , n32773 );
or ( n32775 , n32756 , n32765 );
nand ( n32776 , n32774 , n32775 );
not ( n32777 , n32748 );
and ( n32778 , n32776 , n32777 );
not ( n32779 , n32776 );
and ( n32780 , n32779 , n32748 );
nor ( n32781 , n32778 , n32780 );
not ( n32782 , n32781 );
not ( n32783 , n32782 );
and ( n32784 , n32771 , n32783 );
nor ( n32785 , n32770 , n32784 );
not ( n32786 , n32785 );
not ( n32787 , n32786 );
and ( n32788 , n32694 , n32787 );
and ( n32789 , n32693 , n32786 );
nor ( n32790 , n32788 , n32789 );
not ( n32791 , n32790 );
or ( n32792 , n32538 , n32791 );
or ( n32793 , n32537 , n32790 );
nand ( n210555 , n32792 , n32793 );
buf ( n32795 , RI173f5a88_1558);
not ( n32796 , n32795 );
not ( n32797 , RI173acd98_1913);
not ( n32798 , n32797 );
or ( n32799 , n32796 , n32798 );
not ( n32800 , RI173f5a88_1558);
nand ( n32801 , n32800 , n30043 );
nand ( n32802 , n32799 , n32801 );
buf ( n210564 , RI17524638_653);
and ( n32804 , n32802 , n210564 );
not ( n32805 , n32802 );
not ( n32806 , RI17524638_653);
and ( n32807 , n32805 , n32806 );
nor ( n32808 , n32804 , n32807 );
buf ( n32809 , RI19aae458_2466);
nand ( n32810 , n25803 , n32809 );
buf ( n32811 , RI174920b8_1024);
and ( n32812 , n32810 , n32811 );
not ( n32813 , n32810 );
not ( n32814 , RI174920b8_1024);
and ( n32815 , n32813 , n32814 );
nor ( n32816 , n32812 , n32815 );
xor ( n32817 , n32808 , n32816 );
buf ( n32818 , RI19ac6878_2281);
nand ( n32819 , n26398 , n32818 );
buf ( n32820 , RI1751f3b8_669);
and ( n32821 , n32819 , n32820 );
not ( n32822 , n32819 );
not ( n32823 , RI1751f3b8_669);
and ( n32824 , n32822 , n32823 );
nor ( n32825 , n32821 , n32824 );
xor ( n210587 , n32817 , n32825 );
buf ( n32827 , n210587 );
xor ( n210589 , n28492 , n32827 );
not ( n32829 , RI17450028_1346);
buf ( n32830 , RI19ac9de8_2256);
nand ( n32831 , n25375 , n32830 );
buf ( n32832 , RI174c05d0_812);
and ( n32833 , n32831 , n32832 );
not ( n32834 , n32831 );
not ( n32835 , RI174c05d0_812);
and ( n32836 , n32834 , n32835 );
nor ( n32837 , n32833 , n32836 );
xor ( n32838 , n32829 , n32837 );
buf ( n32839 , RI19a9a610_2609);
nand ( n32840 , n26266 , n32839 );
buf ( n32841 , RI17474838_1168);
and ( n32842 , n32840 , n32841 );
not ( n32843 , n32840 );
not ( n32844 , RI17474838_1168);
and ( n32845 , n32843 , n32844 );
nor ( n32846 , n32842 , n32845 );
xnor ( n32847 , n32838 , n32846 );
not ( n32848 , n32847 );
buf ( n32849 , RI173d8550_1701);
not ( n32850 , n32849 );
not ( n32851 , RI1738f860_2056);
not ( n32852 , n32851 );
or ( n32853 , n32850 , n32852 );
not ( n32854 , RI173d8550_1701);
buf ( n32855 , RI1738f860_2056);
nand ( n32856 , n32854 , n32855 );
nand ( n32857 , n32853 , n32856 );
not ( n32858 , n32857 );
not ( n32859 , n32858 );
and ( n32860 , n32848 , n32859 );
and ( n32861 , n32847 , n32858 );
nor ( n32862 , n32860 , n32861 );
buf ( n32863 , n32862 );
xnor ( n32864 , n210589 , n32863 );
not ( n32865 , n32864 );
not ( n32866 , n29887 );
buf ( n210628 , RI173ca960_1768);
not ( n210629 , n210628 );
not ( n32869 , RI173413e0_2123);
not ( n210631 , n32869 );
or ( n210632 , n210629 , n210631 );
not ( n32872 , RI173ca960_1768);
nand ( n32873 , n32872 , n31732 );
nand ( n32874 , n210632 , n32873 );
buf ( n32875 , RI17413998_1412);
and ( n32876 , n32874 , n32875 );
not ( n32877 , n32874 );
not ( n32878 , RI17413998_1412);
and ( n32879 , n32877 , n32878 );
nor ( n32880 , n32876 , n32879 );
buf ( n32881 , RI19abf2d0_2339);
nand ( n32882 , n25751 , n32881 );
buf ( n32883 , RI174afc80_879);
and ( n32884 , n32882 , n32883 );
not ( n32885 , n32882 );
not ( n32886 , RI174afc80_879);
and ( n32887 , n32885 , n32886 );
nor ( n210649 , n32884 , n32887 );
xor ( n32889 , n32880 , n210649 );
buf ( n32890 , RI19a8e6d0_2694);
nand ( n32891 , n32338 , n32890 );
buf ( n32892 , RI17466fa8_1234);
and ( n32893 , n32891 , n32892 );
not ( n32894 , n32891 );
not ( n32895 , RI17466fa8_1234);
and ( n32896 , n32894 , n32895 );
nor ( n32897 , n32893 , n32896 );
xnor ( n32898 , n32889 , n32897 );
not ( n32899 , n32898 );
not ( n32900 , n32899 );
not ( n32901 , n32900 );
or ( n32902 , n32866 , n32901 );
not ( n32903 , n32898 );
nand ( n32904 , n32903 , n29884 );
nand ( n32905 , n32902 , n32904 );
not ( n32906 , n26475 );
and ( n32907 , n32905 , n32906 );
not ( n32908 , n32905 );
not ( n32909 , n26472 );
not ( n32910 , n32909 );
and ( n32911 , n32908 , n32910 );
nor ( n32912 , n32907 , n32911 );
nand ( n32913 , n32865 , n32912 );
xor ( n32914 , n29219 , n30207 );
buf ( n32915 , n30163 );
not ( n32916 , n32915 );
xnor ( n32917 , n32914 , n32916 );
not ( n32918 , n32917 );
and ( n32919 , n32913 , n32918 );
not ( n32920 , n32913 );
and ( n32921 , n32920 , n32917 );
nor ( n32922 , n32919 , n32921 );
and ( n32923 , n210555 , n32922 );
not ( n32924 , n210555 );
not ( n32925 , n32922 );
and ( n32926 , n32924 , n32925 );
nor ( n32927 , n32923 , n32926 );
buf ( n32928 , n206468 );
buf ( n32929 , RI173ca618_1769);
not ( n32930 , n32929 );
not ( n32931 , RI17341098_2124);
not ( n32932 , n32931 );
or ( n32933 , n32930 , n32932 );
not ( n32934 , RI173ca618_1769);
buf ( n32935 , RI17341098_2124);
nand ( n32936 , n32934 , n32935 );
nand ( n32937 , n32933 , n32936 );
buf ( n32938 , RI17413650_1413);
and ( n32939 , n32937 , n32938 );
not ( n32940 , n32937 );
not ( n32941 , RI17413650_1413);
and ( n32942 , n32940 , n32941 );
nor ( n32943 , n32939 , n32942 );
buf ( n32944 , RI19abf0f0_2340);
nand ( n32945 , n29151 , n32944 );
buf ( n32946 , RI174af938_880);
and ( n32947 , n32945 , n32946 );
not ( n32948 , n32945 );
not ( n32949 , RI174af938_880);
and ( n32950 , n32948 , n32949 );
nor ( n32951 , n32947 , n32950 );
xor ( n32952 , n32943 , n32951 );
buf ( n32953 , RI19a8e478_2695);
nand ( n32954 , n30641 , n32953 );
buf ( n32955 , RI17466c60_1235);
and ( n32956 , n32954 , n32955 );
not ( n32957 , n32954 );
not ( n32958 , RI17466c60_1235);
and ( n32959 , n32957 , n32958 );
nor ( n32960 , n32956 , n32959 );
xnor ( n32961 , n32952 , n32960 );
buf ( n32962 , n32961 );
xor ( n32963 , n32928 , n32962 );
buf ( n32964 , RI173e7eb0_1625);
not ( n32965 , n32964 );
not ( n32966 , RI1739ee78_1981);
not ( n32967 , n32966 );
or ( n32968 , n32965 , n32967 );
not ( n32969 , RI173e7eb0_1625);
buf ( n32970 , RI1739ee78_1981);
nand ( n32971 , n32969 , n32970 );
nand ( n32972 , n32968 , n32971 );
not ( n32973 , RI1745f988_1270);
and ( n32974 , n32972 , n32973 );
not ( n32975 , n32972 );
buf ( n210737 , RI1745f988_1270);
and ( n32977 , n32975 , n210737 );
nor ( n32978 , n32974 , n32977 );
xor ( n32979 , n32978 , n29872 );
buf ( n32980 , RI19aa2068_2552);
nand ( n32981 , n25479 , n32980 );
not ( n32982 , RI17484198_1092);
and ( n32983 , n32981 , n32982 );
not ( n32984 , n32981 );
buf ( n32985 , RI17484198_1092);
and ( n32986 , n32984 , n32985 );
nor ( n32987 , n32983 , n32986 );
xnor ( n32988 , n32979 , n32987 );
buf ( n32989 , n32988 );
xor ( n32990 , n32963 , n32989 );
not ( n32991 , n32990 );
not ( n32992 , n206777 );
not ( n32993 , n208179 );
and ( n32994 , n32992 , n32993 );
and ( n32995 , n206777 , n208179 );
nor ( n32996 , n32994 , n32995 );
not ( n32997 , n205159 );
not ( n32998 , n205176 );
or ( n32999 , n32997 , n32998 );
not ( n33000 , n205159 );
nand ( n33001 , n205175 , n33000 );
nand ( n33002 , n32999 , n33001 );
not ( n33003 , n33002 );
and ( n33004 , n32996 , n33003 );
not ( n33005 , n32996 );
not ( n33006 , n33003 );
and ( n33007 , n33005 , n33006 );
nor ( n33008 , n33004 , n33007 );
not ( n33009 , n33008 );
nand ( n33010 , n32991 , n33009 );
not ( n33011 , n33010 );
buf ( n33012 , RI17406450_1477);
not ( n33013 , n32402 );
xor ( n33014 , n33012 , n33013 );
not ( n33015 , RI173f7b58_1548);
buf ( n33016 , RI173aee68_1903);
and ( n33017 , n33015 , n33016 );
not ( n33018 , n33015 );
not ( n33019 , RI173aee68_1903);
and ( n33020 , n33018 , n33019 );
nor ( n33021 , n33017 , n33020 );
not ( n33022 , n33021 );
buf ( n33023 , RI1733b4b8_2152);
buf ( n33024 , RI19aaaa38_2491);
nand ( n33025 , n26453 , n33024 );
buf ( n33026 , RI17494188_1014);
and ( n33027 , n33025 , n33026 );
not ( n33028 , n33025 );
not ( n33029 , RI17494188_1014);
and ( n33030 , n33028 , n33029 );
nor ( n33031 , n33027 , n33030 );
xor ( n33032 , n33023 , n33031 );
buf ( n33033 , RI19aa4318_2536);
nand ( n33034 , n25803 , n33033 );
not ( n33035 , RI17522748_659);
and ( n33036 , n33034 , n33035 );
not ( n33037 , n33034 );
buf ( n33038 , RI17522748_659);
and ( n33039 , n33037 , n33038 );
nor ( n33040 , n33036 , n33039 );
xnor ( n33041 , n33032 , n33040 );
not ( n33042 , n33041 );
or ( n33043 , n33022 , n33042 );
or ( n33044 , n33041 , n33021 );
nand ( n33045 , n33043 , n33044 );
buf ( n33046 , n33045 );
not ( n33047 , n33046 );
xor ( n33048 , n33014 , n33047 );
not ( n33049 , n33048 );
not ( n33050 , n33049 );
and ( n33051 , n33011 , n33050 );
and ( n33052 , n33010 , n33049 );
nor ( n33053 , n33051 , n33052 );
not ( n33054 , n33053 );
buf ( n33055 , RI19ab29b8_2435);
nand ( n33056 , n25851 , n33055 );
buf ( n33057 , RI174a6f68_922);
and ( n33058 , n33056 , n33057 );
not ( n33059 , n33056 );
not ( n33060 , RI174a6f68_922);
and ( n33061 , n33059 , n33060 );
nor ( n33062 , n33058 , n33061 );
buf ( n33063 , RI173fc388_1526);
not ( n33064 , n33063 );
not ( n33065 , RI173b3350_1882);
not ( n33066 , n33065 );
or ( n33067 , n33064 , n33066 );
not ( n33068 , RI173fc388_1526);
buf ( n33069 , RI173b3350_1882);
nand ( n33070 , n33068 , n33069 );
nand ( n33071 , n33067 , n33070 );
buf ( n33072 , RI173a71b8_1941);
and ( n33073 , n33071 , n33072 );
not ( n33074 , n33071 );
not ( n33075 , RI173a71b8_1941);
and ( n33076 , n33074 , n33075 );
nor ( n33077 , n33073 , n33076 );
buf ( n33078 , RI19a90368_2681);
nand ( n33079 , n25879 , n33078 );
buf ( n33080 , RI17529390_638);
and ( n33081 , n33079 , n33080 );
not ( n33082 , n33079 );
not ( n33083 , RI17529390_638);
and ( n33084 , n33082 , n33083 );
nor ( n33085 , n33081 , n33084 );
xor ( n33086 , n33077 , n33085 );
buf ( n33087 , RI19aa8878_2506);
nand ( n33088 , n26463 , n33087 );
buf ( n33089 , RI17498670_993);
and ( n33090 , n33088 , n33089 );
not ( n33091 , n33088 );
not ( n33092 , RI17498670_993);
and ( n33093 , n33091 , n33092 );
nor ( n33094 , n33090 , n33093 );
xnor ( n33095 , n33086 , n33094 );
buf ( n33096 , n33095 );
and ( n33097 , n33062 , n33096 );
not ( n33098 , n33062 );
not ( n33099 , n33096 );
and ( n33100 , n33098 , n33099 );
nor ( n33101 , n33097 , n33100 );
buf ( n33102 , RI173d0bd0_1738);
not ( n33103 , n33102 );
not ( n33104 , RI17347308_2094);
not ( n33105 , n33104 );
or ( n33106 , n33103 , n33105 );
not ( n33107 , RI173d0bd0_1738);
buf ( n33108 , RI17347308_2094);
nand ( n33109 , n33107 , n33108 );
nand ( n33110 , n33106 , n33109 );
not ( n33111 , RI174486c0_1383);
and ( n33112 , n33110 , n33111 );
not ( n33113 , n33110 );
buf ( n33114 , RI174486c0_1383);
and ( n33115 , n33113 , n33114 );
nor ( n33116 , n33112 , n33115 );
buf ( n33117 , RI19a8af08_2718);
nand ( n33118 , n205019 , n33117 );
buf ( n33119 , RI1746ced0_1205);
and ( n33120 , n33118 , n33119 );
not ( n33121 , n33118 );
not ( n33122 , RI1746ced0_1205);
and ( n33123 , n33121 , n33122 );
nor ( n33124 , n33120 , n33123 );
xor ( n33125 , n33116 , n33124 );
buf ( n33126 , RI19abc8a0_2363);
nand ( n33127 , n25666 , n33126 );
not ( n33128 , RI174b5ba8_850);
and ( n33129 , n33127 , n33128 );
not ( n33130 , n33127 );
buf ( n33131 , RI174b5ba8_850);
and ( n33132 , n33130 , n33131 );
nor ( n33133 , n33129 , n33132 );
xnor ( n33134 , n33125 , n33133 );
buf ( n33135 , n33134 );
and ( n33136 , n33101 , n33135 );
not ( n33137 , n33101 );
not ( n33138 , n33124 );
xor ( n33139 , n33116 , n33138 );
xnor ( n33140 , n33139 , n33133 );
buf ( n33141 , n33140 );
buf ( n33142 , n33141 );
and ( n33143 , n33137 , n33142 );
nor ( n33144 , n33136 , n33143 );
not ( n33145 , n33144 );
not ( n33146 , n204770 );
buf ( n33147 , RI1739ca60_1992);
not ( n33148 , n33147 );
not ( n33149 , RI173e5a98_1636);
not ( n33150 , n33149 );
or ( n33151 , n33148 , n33150 );
not ( n33152 , RI1739ca60_1992);
buf ( n33153 , RI173e5a98_1636);
nand ( n33154 , n33152 , n33153 );
nand ( n33155 , n33151 , n33154 );
and ( n33156 , n33155 , n28211 );
not ( n33157 , n33155 );
and ( n33158 , n33157 , n28252 );
nor ( n33159 , n33156 , n33158 );
buf ( n33160 , RI19a841d0_2765);
nand ( n33161 , n29435 , n33160 );
buf ( n33162 , RI17503de8_748);
and ( n33163 , n33161 , n33162 );
not ( n33164 , n33161 );
not ( n33165 , RI17503de8_748);
and ( n33166 , n33164 , n33165 );
nor ( n33167 , n33163 , n33166 );
xor ( n33168 , n33159 , n33167 );
buf ( n33169 , RI19aa3058_2545);
nand ( n33170 , n25416 , n33169 );
buf ( n33171 , RI17481d80_1103);
and ( n33172 , n33170 , n33171 );
not ( n33173 , n33170 );
not ( n33174 , RI17481d80_1103);
and ( n33175 , n33173 , n33174 );
nor ( n33176 , n33172 , n33175 );
xnor ( n33177 , n33168 , n33176 );
not ( n33178 , n33177 );
not ( n210940 , n33178 );
not ( n210941 , n210940 );
or ( n33181 , n33146 , n210941 );
buf ( n33182 , n33177 );
buf ( n33183 , n33182 );
or ( n33184 , n33183 , n204770 );
nand ( n33185 , n33181 , n33184 );
not ( n33186 , n31037 );
not ( n33187 , n33186 );
and ( n33188 , n33185 , n33187 );
not ( n33189 , n33185 );
and ( n33190 , n33189 , n33186 );
nor ( n33191 , n33188 , n33190 );
nand ( n210953 , n33145 , n33191 );
not ( n33193 , n210953 );
buf ( n33194 , RI173eaca0_1611);
buf ( n33195 , n207059 );
xor ( n33196 , n33194 , n33195 );
not ( n33197 , RI173dc3a8_1682);
not ( n33198 , n33197 );
buf ( n33199 , RI173936b8_2037);
not ( n33200 , n33199 );
and ( n33201 , n33198 , n33200 );
and ( n33202 , n33199 , n33197 );
nor ( n33203 , n33201 , n33202 );
not ( n33204 , n33203 );
not ( n33205 , n33204 );
not ( n33206 , RI17453e80_1327);
buf ( n33207 , RI19ac7d90_2271);
nand ( n33208 , n26242 , n33207 );
buf ( n33209 , RI174c67c8_793);
and ( n33210 , n33208 , n33209 );
not ( n33211 , n33208 );
not ( n33212 , RI174c67c8_793);
and ( n33213 , n33211 , n33212 );
nor ( n33214 , n33210 , n33213 );
xor ( n33215 , n33206 , n33214 );
buf ( n33216 , RI19a98018_2626);
nand ( n33217 , n204572 , n33216 );
buf ( n33218 , RI174789d8_1148);
and ( n33219 , n33217 , n33218 );
not ( n33220 , n33217 );
not ( n33221 , RI174789d8_1148);
and ( n33222 , n33220 , n33221 );
nor ( n33223 , n33219 , n33222 );
xnor ( n33224 , n33215 , n33223 );
not ( n33225 , n33224 );
not ( n33226 , n33225 );
or ( n210988 , n33205 , n33226 );
nand ( n33228 , n33224 , n33203 );
nand ( n33229 , n210988 , n33228 );
not ( n33230 , n33229 );
xnor ( n33231 , n33196 , n33230 );
not ( n33232 , n33231 );
not ( n33233 , n33232 );
or ( n33234 , n33193 , n33233 );
or ( n33235 , n33232 , n210953 );
nand ( n33236 , n33234 , n33235 );
not ( n33237 , n33236 );
and ( n33238 , n33054 , n33237 );
and ( n33239 , n33053 , n33236 );
nor ( n33240 , n33238 , n33239 );
not ( n33241 , n33240 );
not ( n33242 , n33241 );
and ( n33243 , n32927 , n33242 );
not ( n33244 , n32927 );
and ( n33245 , n33244 , n33241 );
nor ( n33246 , n33243 , n33245 );
buf ( n33247 , n33246 );
not ( n33248 , n33247 );
and ( n33249 , n32478 , n33248 );
and ( n33250 , n32477 , n33247 );
nor ( n33251 , n33249 , n33250 );
buf ( n33252 , n27885 );
buf ( n33253 , n33252 );
buf ( n33254 , n33253 );
not ( n33255 , n33254 );
nand ( n33256 , n33251 , n33255 );
buf ( n33257 , RI173406c0_2127);
not ( n33258 , n33257 );
not ( n33259 , n205142 );
or ( n33260 , n33258 , n33259 );
buf ( n33261 , n205095 );
not ( n33262 , n33261 );
or ( n33263 , n33262 , n33257 );
nand ( n33264 , n33260 , n33263 );
not ( n33265 , n33264 );
not ( n33266 , RI17450370_1345);
buf ( n33267 , RI19aca040_2255);
nand ( n33268 , n25582 , n33267 );
buf ( n33269 , RI174c0af8_811);
and ( n33270 , n33268 , n33269 );
not ( n33271 , n33268 );
not ( n33272 , RI174c0af8_811);
and ( n33273 , n33271 , n33272 );
nor ( n33274 , n33270 , n33273 );
xor ( n33275 , n33266 , n33274 );
buf ( n33276 , RI19a9a868_2608);
nand ( n33277 , n25803 , n33276 );
buf ( n33278 , RI17474b80_1167);
and ( n33279 , n33277 , n33278 );
not ( n33280 , n33277 );
not ( n33281 , RI17474b80_1167);
and ( n33282 , n33280 , n33281 );
nor ( n33283 , n33279 , n33282 );
xnor ( n33284 , n33275 , n33283 );
not ( n33285 , n33284 );
buf ( n33286 , RI173d8898_1700);
not ( n33287 , n33286 );
not ( n33288 , RI1738fba8_2055);
not ( n33289 , n33288 );
or ( n33290 , n33287 , n33289 );
not ( n33291 , RI173d8898_1700);
buf ( n33292 , RI1738fba8_2055);
nand ( n33293 , n33291 , n33292 );
nand ( n33294 , n33290 , n33293 );
not ( n33295 , n33294 );
not ( n33296 , n33295 );
and ( n33297 , n33285 , n33296 );
and ( n33298 , n33284 , n33295 );
nor ( n33299 , n33297 , n33298 );
buf ( n33300 , n33299 );
not ( n33301 , n33300 );
and ( n33302 , n33265 , n33301 );
buf ( n33303 , n33299 );
and ( n33304 , n33264 , n33303 );
nor ( n33305 , n33302 , n33304 );
not ( n33306 , n33305 );
not ( n33307 , n33306 );
not ( n33308 , n204478 );
not ( n33309 , n25931 );
or ( n33310 , n33308 , n33309 );
not ( n33311 , n204478 );
nand ( n33312 , n33311 , n25926 );
nand ( n33313 , n33310 , n33312 );
and ( n33314 , n33313 , n25965 );
not ( n33315 , n33313 );
and ( n33316 , n33315 , n25978 );
nor ( n33317 , n33314 , n33316 );
nand ( n33318 , n28293 , n33317 );
not ( n33319 , n33318 );
and ( n33320 , n33307 , n33319 );
and ( n33321 , n33306 , n33318 );
nor ( n33322 , n33320 , n33321 );
not ( n33323 , n33322 );
not ( n33324 , n33323 );
not ( n33325 , n27971 );
not ( n33326 , n205426 );
not ( n33327 , n29271 );
buf ( n33328 , RI173a22f8_1965);
not ( n33329 , n33328 );
not ( n33330 , RI173eafe8_1610);
not ( n33331 , n33330 );
or ( n33332 , n33329 , n33331 );
not ( n33333 , RI173a22f8_1965);
buf ( n33334 , RI173eafe8_1610);
nand ( n33335 , n33333 , n33334 );
nand ( n33336 , n33332 , n33335 );
buf ( n33337 , RI17473140_1175);
and ( n33338 , n33336 , n33337 );
not ( n33339 , n33336 );
not ( n33340 , RI17473140_1175);
and ( n33341 , n33339 , n33340 );
nor ( n33342 , n33338 , n33341 );
not ( n33343 , n33342 );
buf ( n33344 , RI19a9f908_2572);
nand ( n33345 , n25376 , n33344 );
buf ( n33346 , RI174872d0_1077);
and ( n33347 , n33345 , n33346 );
not ( n33348 , n33345 );
not ( n33349 , RI174872d0_1077);
and ( n33350 , n33348 , n33349 );
nor ( n33351 , n33347 , n33350 );
buf ( n33352 , n33351 );
xor ( n33353 , n33343 , n33352 );
buf ( n33354 , RI19ace618_2222);
nand ( n33355 , n25752 , n33354 );
not ( n33356 , RI1750e270_722);
and ( n33357 , n33355 , n33356 );
not ( n33358 , n33355 );
buf ( n33359 , RI1750e270_722);
and ( n33360 , n33358 , n33359 );
nor ( n33361 , n33357 , n33360 );
xnor ( n33362 , n33353 , n33361 );
not ( n33363 , n33362 );
or ( n33364 , n33327 , n33363 );
xor ( n33365 , n33342 , n33351 );
xnor ( n33366 , n33365 , n33361 );
nand ( n33367 , n33366 , n29267 );
nand ( n33368 , n33364 , n33367 );
not ( n33369 , n33368 );
and ( n33370 , n33326 , n33369 );
and ( n33371 , n205426 , n33368 );
nor ( n33372 , n33370 , n33371 );
nand ( n33373 , n33372 , n28605 );
not ( n33374 , n33373 );
or ( n33375 , n33325 , n33374 );
or ( n33376 , n33373 , n27971 );
nand ( n33377 , n33375 , n33376 );
not ( n33378 , n33377 );
not ( n33379 , n33378 );
or ( n33380 , n33324 , n33379 );
nand ( n33381 , n33377 , n33322 );
nand ( n33382 , n33380 , n33381 );
not ( n211144 , n33382 );
not ( n33384 , n25826 );
xor ( n33385 , n29420 , n33384 );
buf ( n33386 , RI173fb320_1531);
buf ( n33387 , RI1740ca08_1446);
not ( n33388 , n33387 );
not ( n33389 , RI173c3d18_1801);
not ( n33390 , n33389 );
or ( n33391 , n33388 , n33390 );
not ( n33392 , RI1740ca08_1446);
buf ( n33393 , RI173c3d18_1801);
nand ( n33394 , n33392 , n33393 );
nand ( n33395 , n33391 , n33394 );
xor ( n33396 , n33386 , n33395 );
buf ( n33397 , RI1733a798_2156);
not ( n33398 , RI174a9038_912);
xor ( n33399 , n33397 , n33398 );
buf ( n33400 , RI19ab16f8_2443);
nand ( n33401 , n205124 , n33400 );
xnor ( n33402 , n33399 , n33401 );
xnor ( n33403 , n33396 , n33402 );
not ( n33404 , n33403 );
xnor ( n33405 , n33385 , n33404 );
not ( n33406 , n33405 );
nand ( n33407 , n33406 , n28516 );
not ( n33408 , n33407 );
buf ( n33409 , RI173c3688_1803);
not ( n33410 , n33409 );
buf ( n33411 , RI173fddc8_1518);
not ( n33412 , n33411 );
not ( n33413 , RI173b4d90_1874);
not ( n33414 , n33413 );
or ( n33415 , n33412 , n33414 );
not ( n33416 , RI173fddc8_1518);
buf ( n33417 , RI173b4d90_1874);
nand ( n33418 , n33416 , n33417 );
nand ( n33419 , n33415 , n33418 );
not ( n33420 , RI173b71a8_1863);
and ( n33421 , n33419 , n33420 );
not ( n33422 , n33419 );
buf ( n33423 , RI173b71a8_1863);
and ( n33424 , n33422 , n33423 );
nor ( n33425 , n33421 , n33424 );
buf ( n33426 , RI19a88208_2737);
nand ( n33427 , n30640 , n33426 );
buf ( n33428 , RI1752bcd0_630);
and ( n33429 , n33427 , n33428 );
not ( n33430 , n33427 );
not ( n33431 , RI1752bcd0_630);
and ( n33432 , n33430 , n33431 );
nor ( n33433 , n33429 , n33432 );
xor ( n33434 , n33425 , n33433 );
buf ( n33435 , RI19aa7090_2516);
nand ( n33436 , n204336 , n33435 );
buf ( n33437 , RI1749a0b0_985);
and ( n33438 , n33436 , n33437 );
not ( n33439 , n33436 );
not ( n33440 , RI1749a0b0_985);
and ( n33441 , n33439 , n33440 );
nor ( n33442 , n33438 , n33441 );
xor ( n33443 , n33434 , n33442 );
buf ( n33444 , n33443 );
not ( n33445 , n33444 );
or ( n33446 , n33410 , n33445 );
or ( n33447 , n33444 , n33409 );
nand ( n33448 , n33446 , n33447 );
buf ( n33449 , RI173d22e0_1731);
not ( n33450 , n33449 );
not ( n33451 , RI173892a8_2087);
not ( n33452 , n33451 );
or ( n33453 , n33450 , n33452 );
not ( n33454 , RI173d22e0_1731);
buf ( n33455 , RI173892a8_2087);
nand ( n33456 , n33454 , n33455 );
nand ( n33457 , n33453 , n33456 );
buf ( n211219 , RI17449db8_1376);
and ( n33459 , n33457 , n211219 );
not ( n33460 , n33457 );
not ( n33461 , RI17449db8_1376);
and ( n33462 , n33460 , n33461 );
nor ( n33463 , n33459 , n33462 );
buf ( n33464 , RI19a89720_2728);
nand ( n33465 , n206902 , n33464 );
buf ( n33466 , RI1746e5c8_1198);
and ( n33467 , n33465 , n33466 );
not ( n33468 , n33465 );
not ( n33469 , RI1746e5c8_1198);
and ( n33470 , n33468 , n33469 );
nor ( n33471 , n33467 , n33470 );
xor ( n33472 , n33463 , n33471 );
xnor ( n33473 , n33472 , n32346 );
not ( n33474 , n33473 );
not ( n33475 , n33474 );
and ( n33476 , n33448 , n33475 );
not ( n33477 , n33448 );
and ( n33478 , n33477 , n33474 );
nor ( n33479 , n33476 , n33478 );
not ( n33480 , n33479 );
not ( n33481 , n33480 );
not ( n33482 , n33481 );
and ( n33483 , n33408 , n33482 );
and ( n33484 , n33407 , n33481 );
nor ( n33485 , n33483 , n33484 );
not ( n33486 , n33485 );
and ( n33487 , n211144 , n33486 );
and ( n33488 , n33382 , n33485 );
nor ( n33489 , n33487 , n33488 );
not ( n33490 , n32415 );
buf ( n33491 , RI173daff8_1688);
not ( n33492 , n33491 );
not ( n33493 , RI17392308_2043);
not ( n33494 , n33493 );
or ( n33495 , n33492 , n33494 );
not ( n33496 , RI173daff8_1688);
buf ( n33497 , RI17392308_2043);
nand ( n33498 , n33496 , n33497 );
nand ( n33499 , n33495 , n33498 );
buf ( n33500 , RI17452ad0_1333);
and ( n33501 , n33499 , n33500 );
not ( n33502 , n33499 );
not ( n33503 , RI17452ad0_1333);
and ( n33504 , n33502 , n33503 );
nor ( n33505 , n33501 , n33504 );
buf ( n33506 , RI19ac7250_2276);
nand ( n33507 , n25803 , n33506 );
buf ( n33508 , RI174c48d8_799);
and ( n211270 , n33507 , n33508 );
not ( n211271 , n33507 );
not ( n33511 , RI174c48d8_799);
and ( n33512 , n211271 , n33511 );
nor ( n33513 , n211270 , n33512 );
xor ( n33514 , n33505 , n33513 );
buf ( n33515 , RI19a97460_2631);
nand ( n33516 , n26266 , n33515 );
buf ( n33517 , RI174772e0_1155);
and ( n33518 , n33516 , n33517 );
not ( n33519 , n33516 );
not ( n33520 , RI174772e0_1155);
and ( n33521 , n33519 , n33520 );
nor ( n33522 , n33518 , n33521 );
not ( n33523 , n33522 );
xnor ( n33524 , n33514 , n33523 );
not ( n33525 , n33524 );
not ( n33526 , n33525 );
or ( n33527 , n33490 , n33526 );
not ( n33528 , n33525 );
nand ( n33529 , n33528 , n32411 );
nand ( n33530 , n33527 , n33529 );
buf ( n33531 , RI173f8530_1545);
not ( n33532 , n33531 );
not ( n33533 , RI173af840_1900);
not ( n33534 , n33533 );
or ( n33535 , n33532 , n33534 );
not ( n33536 , RI173f8530_1545);
buf ( n33537 , RI173af840_1900);
nand ( n33538 , n33536 , n33537 );
nand ( n33539 , n33535 , n33538 );
not ( n33540 , RI17342100_2119);
and ( n211302 , n33539 , n33540 );
not ( n33542 , n33539 );
buf ( n33543 , RI17342100_2119);
and ( n33544 , n33542 , n33543 );
nor ( n33545 , n211302 , n33544 );
buf ( n33546 , RI19aa8f80_2503);
nand ( n33547 , n25711 , n33546 );
buf ( n33548 , RI175236c0_656);
and ( n33549 , n33547 , n33548 );
not ( n33550 , n33547 );
not ( n33551 , RI175236c0_656);
and ( n33552 , n33550 , n33551 );
nor ( n33553 , n33549 , n33552 );
xor ( n33554 , n33545 , n33553 );
buf ( n33555 , RI19aab0c8_2488);
nand ( n33556 , n204426 , n33555 );
buf ( n33557 , RI17494b60_1011);
and ( n33558 , n33556 , n33557 );
not ( n33559 , n33556 );
not ( n33560 , RI17494b60_1011);
and ( n33561 , n33559 , n33560 );
nor ( n33562 , n33558 , n33561 );
xnor ( n33563 , n33554 , n33562 );
buf ( n33564 , n33563 );
not ( n33565 , n33564 );
buf ( n33566 , n33565 );
not ( n33567 , n33566 );
and ( n33568 , n33530 , n33567 );
not ( n33569 , n33530 );
and ( n33570 , n33569 , n33566 );
nor ( n33571 , n33568 , n33570 );
not ( n33572 , n33571 );
nand ( n33573 , n28913 , n33572 );
not ( n33574 , n32113 );
not ( n33575 , n29860 );
or ( n33576 , n33574 , n33575 );
not ( n33577 , n29854 );
nand ( n33578 , n33577 , n32109 );
nand ( n33579 , n33576 , n33578 );
buf ( n33580 , RI173e8bd0_1621);
not ( n33581 , n33580 );
not ( n33582 , RI1739fb98_1977);
not ( n33583 , n33582 );
or ( n33584 , n33581 , n33583 );
not ( n33585 , RI173e8bd0_1621);
buf ( n33586 , RI1739fb98_1977);
nand ( n33587 , n33585 , n33586 );
nand ( n33588 , n33584 , n33587 );
not ( n33589 , RI174606a8_1266);
and ( n33590 , n33588 , n33589 );
not ( n33591 , n33588 );
buf ( n33592 , RI174606a8_1266);
and ( n33593 , n33591 , n33592 );
nor ( n33594 , n33590 , n33593 );
buf ( n33595 , RI19aa2c20_2547);
nand ( n33596 , n29890 , n33595 );
buf ( n33597 , RI17484eb8_1088);
and ( n33598 , n33596 , n33597 );
not ( n33599 , n33596 );
not ( n33600 , RI17484eb8_1088);
and ( n33601 , n33599 , n33600 );
nor ( n33602 , n33598 , n33601 );
xor ( n33603 , n33594 , n33602 );
buf ( n33604 , RI19a83d20_2767);
nand ( n33605 , n25711 , n33604 );
buf ( n33606 , RI1750a9b8_733);
and ( n33607 , n33605 , n33606 );
not ( n33608 , n33605 );
not ( n33609 , RI1750a9b8_733);
and ( n33610 , n33608 , n33609 );
nor ( n33611 , n33607 , n33610 );
not ( n33612 , n33611 );
xnor ( n33613 , n33603 , n33612 );
buf ( n33614 , n33613 );
and ( n33615 , n33579 , n33614 );
not ( n33616 , n33579 );
xor ( n33617 , n33594 , n33611 );
xnor ( n33618 , n33617 , n33602 );
buf ( n33619 , n33618 );
and ( n33620 , n33616 , n33619 );
nor ( n33621 , n33615 , n33620 );
xnor ( n33622 , n33573 , n33621 );
not ( n33623 , n33622 );
buf ( n33624 , RI173caff0_1766);
not ( n33625 , n33624 );
not ( n33626 , RI17341a70_2121);
not ( n33627 , n33626 );
or ( n33628 , n33625 , n33627 );
not ( n33629 , RI173caff0_1766);
buf ( n33630 , RI17341a70_2121);
nand ( n33631 , n33629 , n33630 );
nand ( n33632 , n33628 , n33631 );
buf ( n33633 , RI17414028_1410);
and ( n33634 , n33632 , n33633 );
not ( n33635 , n33632 );
not ( n33636 , RI17414028_1410);
and ( n33637 , n33635 , n33636 );
nor ( n33638 , n33634 , n33637 );
buf ( n33639 , RI19a8ed60_2691);
nand ( n33640 , n25741 , n33639 );
buf ( n33641 , RI17467638_1232);
and ( n33642 , n33640 , n33641 );
not ( n33643 , n33640 );
not ( n33644 , RI17467638_1232);
and ( n33645 , n33643 , n33644 );
nor ( n33646 , n33642 , n33645 );
not ( n33647 , n33646 );
xor ( n33648 , n33638 , n33647 );
buf ( n33649 , RI19abf870_2336);
nand ( n33650 , n26463 , n33649 );
not ( n33651 , RI174b0310_877);
and ( n33652 , n33650 , n33651 );
not ( n33653 , n33650 );
buf ( n33654 , RI174b0310_877);
and ( n33655 , n33653 , n33654 );
nor ( n33656 , n33652 , n33655 );
xnor ( n33657 , n33648 , n33656 );
buf ( n211419 , n33657 );
not ( n33659 , n211419 );
buf ( n33660 , RI174053e8_1482);
not ( n33661 , n33660 );
not ( n33662 , n207706 );
or ( n33663 , n33661 , n33662 );
or ( n33664 , n207706 , n33660 );
nand ( n33665 , n33663 , n33664 );
not ( n33666 , n33665 );
or ( n33667 , n33659 , n33666 );
or ( n33668 , n33665 , n211419 );
nand ( n33669 , n33667 , n33668 );
not ( n33670 , n33669 );
not ( n33671 , n206427 );
nand ( n33672 , n33670 , n33671 );
not ( n33673 , n33672 );
nand ( n33674 , n30220 , n205181 );
not ( n33675 , n33674 );
nor ( n33676 , n30220 , n205181 );
nor ( n33677 , n33675 , n33676 );
not ( n33678 , n33677 );
not ( n33679 , n31773 );
not ( n33680 , n33679 );
not ( n33681 , n31762 );
or ( n33682 , n33680 , n33681 );
or ( n33683 , n31762 , n33679 );
nand ( n33684 , n33682 , n33683 );
buf ( n33685 , n33684 );
not ( n33686 , n33685 );
or ( n33687 , n33678 , n33686 );
or ( n33688 , n33685 , n33677 );
nand ( n33689 , n33687 , n33688 );
not ( n33690 , n33689 );
not ( n33691 , n33690 );
not ( n33692 , n33691 );
and ( n33693 , n33673 , n33692 );
not ( n33694 , n33669 );
nand ( n33695 , n33694 , n33671 );
and ( n33696 , n33695 , n33691 );
nor ( n33697 , n33693 , n33696 );
not ( n33698 , n33697 );
not ( n33699 , n33698 );
or ( n33700 , n33623 , n33699 );
not ( n33701 , n33622 );
nand ( n33702 , n33701 , n33697 );
nand ( n33703 , n33700 , n33702 );
and ( n33704 , n33489 , n33703 );
not ( n33705 , n33489 );
not ( n33706 , n33703 );
and ( n33707 , n33705 , n33706 );
nor ( n33708 , n33704 , n33707 );
buf ( n33709 , n33708 );
not ( n33710 , n33709 );
not ( n33711 , n205230 );
buf ( n33712 , RI173a6e70_1942);
not ( n33713 , n33712 );
not ( n33714 , n205236 );
or ( n33715 , n33713 , n33714 );
or ( n33716 , n205236 , n33712 );
nand ( n33717 , n33715 , n33716 );
not ( n33718 , n33717 );
and ( n33719 , n33711 , n33718 );
and ( n33720 , n25868 , n33717 );
nor ( n33721 , n33719 , n33720 );
not ( n33722 , n27827 );
not ( n33723 , n33194 );
not ( n33724 , RI173a1fb0_1966);
not ( n33725 , n33724 );
or ( n33726 , n33723 , n33725 );
not ( n33727 , RI173eaca0_1611);
buf ( n33728 , RI173a1fb0_1966);
nand ( n33729 , n33727 , n33728 );
nand ( n33730 , n33726 , n33729 );
buf ( n33731 , RI17470d28_1186);
and ( n33732 , n33730 , n33731 );
not ( n33733 , n33730 );
not ( n33734 , RI17470d28_1186);
and ( n33735 , n33733 , n33734 );
nor ( n33736 , n33732 , n33735 );
buf ( n33737 , RI19aa19d8_2555);
nand ( n33738 , n25793 , n33737 );
not ( n33739 , RI17486f88_1078);
and ( n33740 , n33738 , n33739 );
not ( n33741 , n33738 );
buf ( n33742 , RI17486f88_1078);
and ( n33743 , n33741 , n33742 );
nor ( n33744 , n33740 , n33743 );
xor ( n33745 , n33736 , n33744 );
buf ( n33746 , RI19a82b50_2775);
nand ( n33747 , n25880 , n33746 );
not ( n33748 , RI1750dd48_723);
and ( n33749 , n33747 , n33748 );
not ( n33750 , n33747 );
buf ( n33751 , RI1750dd48_723);
and ( n33752 , n33750 , n33751 );
nor ( n33753 , n33749 , n33752 );
xnor ( n33754 , n33745 , n33753 );
not ( n33755 , n33754 );
not ( n33756 , n33755 );
not ( n33757 , n33756 );
or ( n33758 , n33722 , n33757 );
not ( n33759 , n33754 );
not ( n33760 , n33759 );
or ( n33761 , n33760 , n27827 );
nand ( n33762 , n33758 , n33761 );
not ( n33763 , n33762 );
not ( n33764 , n31253 );
not ( n33765 , n33764 );
or ( n33766 , n33763 , n33765 );
not ( n33767 , n31254 );
not ( n33768 , n33767 );
or ( n33769 , n33768 , n33762 );
nand ( n33770 , n33766 , n33769 );
nand ( n33771 , n33721 , n33770 );
not ( n33772 , RI173f0538_1584);
and ( n33773 , n33772 , n29020 );
not ( n33774 , n33772 );
not ( n33775 , RI173a7848_1939);
and ( n33776 , n33774 , n33775 );
nor ( n33777 , n33773 , n33776 );
buf ( n33778 , RI19acd100_2231);
nand ( n33779 , n30640 , n33778 );
buf ( n33780 , RI17516da8_695);
and ( n33781 , n33779 , n33780 );
not ( n211543 , n33779 );
not ( n211544 , RI17516da8_695);
and ( n33784 , n211543 , n211544 );
nor ( n33785 , n33781 , n33784 );
not ( n33786 , n33785 );
buf ( n33787 , n25914 );
buf ( n33788 , RI19a9e468_2582);
nand ( n33789 , n33787 , n33788 );
not ( n33790 , RI1748c820_1051);
and ( n33791 , n33789 , n33790 );
not ( n33792 , n33789 );
buf ( n33793 , RI1748c820_1051);
and ( n33794 , n33792 , n33793 );
nor ( n33795 , n33791 , n33794 );
not ( n33796 , n33795 );
or ( n33797 , n33786 , n33796 );
not ( n33798 , n33795 );
not ( n33799 , n33785 );
nand ( n33800 , n33798 , n33799 );
nand ( n33801 , n33797 , n33800 );
not ( n33802 , RI174a7940_919);
and ( n33803 , n33801 , n33802 );
not ( n33804 , n33801 );
buf ( n33805 , RI174a7940_919);
and ( n33806 , n33804 , n33805 );
nor ( n33807 , n33803 , n33806 );
not ( n33808 , n33807 );
and ( n33809 , n33777 , n33808 );
not ( n33810 , n33777 );
and ( n33811 , n33810 , n33807 );
nor ( n33812 , n33809 , n33811 );
not ( n33813 , n33812 );
buf ( n33814 , n27959 );
not ( n33815 , n33814 );
buf ( n33816 , RI173d3000_1727);
not ( n33817 , n33816 );
not ( n33818 , RI1738a310_2082);
not ( n33819 , n33818 );
or ( n33820 , n33817 , n33819 );
not ( n33821 , RI173d3000_1727);
buf ( n33822 , RI1738a310_2082);
nand ( n33823 , n33821 , n33822 );
nand ( n33824 , n33820 , n33823 );
not ( n33825 , RI1744aad8_1372);
and ( n33826 , n33824 , n33825 );
not ( n33827 , n33824 );
buf ( n33828 , RI1744aad8_1372);
and ( n33829 , n33827 , n33828 );
nor ( n33830 , n33826 , n33829 );
buf ( n33831 , RI19abbc70_2369);
nand ( n33832 , n25479 , n33831 );
buf ( n33833 , RI174b7fc0_839);
and ( n33834 , n33832 , n33833 );
not ( n33835 , n33832 );
not ( n33836 , RI174b7fc0_839);
and ( n33837 , n33835 , n33836 );
nor ( n33838 , n33834 , n33837 );
xor ( n33839 , n33830 , n33838 );
buf ( n33840 , RI19a8a080_2724);
nand ( n33841 , n26059 , n33840 );
not ( n33842 , RI1746f2e8_1194);
and ( n33843 , n33841 , n33842 );
not ( n33844 , n33841 );
buf ( n33845 , RI1746f2e8_1194);
and ( n33846 , n33844 , n33845 );
nor ( n33847 , n33843 , n33846 );
xnor ( n33848 , n33839 , n33847 );
buf ( n33849 , n33848 );
not ( n33850 , n33849 );
or ( n33851 , n33815 , n33850 );
not ( n33852 , n33814 );
not ( n33853 , n33848 );
nand ( n33854 , n33852 , n33853 );
nand ( n33855 , n33851 , n33854 );
not ( n33856 , n33855 );
and ( n33857 , n33813 , n33856 );
not ( n33858 , n33812 );
not ( n33859 , n33858 );
and ( n33860 , n33859 , n33855 );
nor ( n33861 , n33857 , n33860 );
and ( n33862 , n33771 , n33861 );
not ( n33863 , n33771 );
not ( n33864 , n33861 );
and ( n33865 , n33863 , n33864 );
nor ( n33866 , n33862 , n33865 );
not ( n33867 , n33866 );
buf ( n33868 , RI17457cd8_1308);
buf ( n33869 , RI17409240_1463);
not ( n33870 , n33869 );
not ( n33871 , RI173c0550_1818);
not ( n33872 , n33871 );
or ( n33873 , n33870 , n33872 );
not ( n33874 , RI17409240_1463);
buf ( n33875 , RI173c0550_1818);
nand ( n33876 , n33874 , n33875 );
nand ( n33877 , n33873 , n33876 );
xor ( n33878 , n33868 , n33877 );
buf ( n33879 , RI17336fd0_2173);
buf ( n33880 , RI174a5870_929);
xor ( n33881 , n33879 , n33880 );
buf ( n33882 , RI19ab3de0_2424);
nand ( n33883 , n27749 , n33882 );
xnor ( n33884 , n33881 , n33883 );
xnor ( n33885 , n33878 , n33884 );
buf ( n33886 , n33885 );
not ( n33887 , n33886 );
not ( n33888 , n204318 );
not ( n33889 , n30405 );
or ( n33890 , n33888 , n33889 );
not ( n33891 , n208165 );
nand ( n33892 , n33891 , n204314 );
nand ( n33893 , n33890 , n33892 );
not ( n33894 , n33893 );
or ( n33895 , n33887 , n33894 );
or ( n33896 , n33886 , n33893 );
nand ( n33897 , n33895 , n33896 );
not ( n33898 , n26045 );
not ( n33899 , n29174 );
or ( n33900 , n33898 , n33899 );
not ( n33901 , n26045 );
nand ( n33902 , n33901 , n29161 );
nand ( n33903 , n33900 , n33902 );
buf ( n33904 , RI173f6118_1556);
not ( n33905 , n33904 );
not ( n33906 , n204729 );
or ( n33907 , n33905 , n33906 );
not ( n33908 , RI173f6118_1556);
nand ( n33909 , n33908 , n204689 );
nand ( n33910 , n33907 , n33909 );
not ( n33911 , RI1752b7a8_631);
and ( n33912 , n33910 , n33911 );
not ( n33913 , n33910 );
buf ( n33914 , RI1752b7a8_631);
and ( n33915 , n33913 , n33914 );
nor ( n33916 , n33912 , n33915 );
not ( n33917 , n33916 );
buf ( n33918 , RI19ab2508_2437);
nand ( n33919 , n25405 , n33918 );
buf ( n33920 , RI1751fe08_667);
and ( n33921 , n33919 , n33920 );
not ( n33922 , n33919 );
not ( n33923 , RI1751fe08_667);
and ( n33924 , n33922 , n33923 );
nor ( n33925 , n33921 , n33924 );
xor ( n33926 , n33917 , n33925 );
buf ( n33927 , RI19aac040_2482);
nand ( n33928 , n30356 , n33927 );
buf ( n33929 , RI17492748_1022);
and ( n33930 , n33928 , n33929 );
not ( n33931 , n33928 );
not ( n33932 , RI17492748_1022);
and ( n33933 , n33931 , n33932 );
nor ( n33934 , n33930 , n33933 );
xnor ( n33935 , n33926 , n33934 );
buf ( n33936 , n33935 );
not ( n33937 , n33936 );
and ( n33938 , n33903 , n33937 );
not ( n33939 , n33903 );
and ( n33940 , n33939 , n33936 );
nor ( n33941 , n33938 , n33940 );
not ( n33942 , n33941 );
nand ( n33943 , n33897 , n33942 );
buf ( n33944 , n204599 );
not ( n33945 , n33944 );
xor ( n33946 , n207891 , n30134 );
xnor ( n33947 , n33946 , n28081 );
not ( n33948 , n33947 );
not ( n33949 , n33948 );
or ( n33950 , n33945 , n33949 );
or ( n33951 , n33948 , n33944 );
nand ( n33952 , n33950 , n33951 );
not ( n33953 , n31323 );
not ( n33954 , n33953 );
and ( n33955 , n33952 , n33954 );
not ( n33956 , n33952 );
buf ( n33957 , n31317 );
and ( n33958 , n33956 , n33957 );
nor ( n33959 , n33955 , n33958 );
buf ( n33960 , n33959 );
not ( n33961 , n33960 );
and ( n33962 , n33943 , n33961 );
not ( n33963 , n33943 );
and ( n33964 , n33963 , n33960 );
nor ( n33965 , n33962 , n33964 );
not ( n33966 , n33965 );
not ( n33967 , n33966 );
buf ( n33968 , RI173db688_1686);
buf ( n33969 , RI173b88a0_1856);
not ( n33970 , n33969 );
not ( n33971 , RI17401590_1501);
not ( n33972 , n33971 );
or ( n33973 , n33970 , n33972 );
not ( n33974 , RI173b88a0_1856);
buf ( n33975 , RI17401590_1501);
nand ( n33976 , n33974 , n33975 );
nand ( n33977 , n33973 , n33976 );
xor ( n33978 , n33968 , n33977 );
buf ( n33979 , RI17531478_613);
not ( n33980 , RI1749d878_968);
xor ( n33981 , n33979 , n33980 );
buf ( n33982 , RI19ab8958_2391);
nand ( n33983 , n25376 , n33982 );
xnor ( n33984 , n33981 , n33983 );
xnor ( n33985 , n33978 , n33984 );
not ( n33986 , n33985 );
not ( n33987 , n33986 );
buf ( n33988 , RI19a23510_2794);
nand ( n33989 , n205271 , n33988 );
not ( n33990 , RI1751a660_684);
and ( n33991 , n33989 , n33990 );
not ( n33992 , n33989 );
buf ( n33993 , RI1751a660_684);
and ( n33994 , n33992 , n33993 );
nor ( n33995 , n33991 , n33994 );
not ( n33996 , n33995 );
not ( n33997 , n30888 );
or ( n33998 , n33996 , n33997 );
not ( n33999 , n33995 );
nand ( n34000 , n33999 , n30889 );
nand ( n34001 , n33998 , n34000 );
not ( n34002 , n34001 );
and ( n34003 , n33987 , n34002 );
buf ( n34004 , n33986 );
and ( n34005 , n34004 , n34001 );
nor ( n34006 , n34003 , n34005 );
not ( n34007 , n204869 );
buf ( n34008 , RI19a88028_2738);
nand ( n34009 , n25879 , n34008 );
buf ( n34010 , RI1752b280_632);
and ( n34011 , n34009 , n34010 );
not ( n34012 , n34009 );
not ( n34013 , RI1752b280_632);
and ( n34014 , n34012 , n34013 );
nor ( n34015 , n34011 , n34014 );
not ( n34016 , n34015 );
buf ( n34017 , RI19aa6d48_2517);
nand ( n34018 , n30356 , n34017 );
not ( n34019 , RI17499a20_987);
and ( n34020 , n34018 , n34019 );
not ( n34021 , n34018 );
buf ( n34022 , RI17499a20_987);
and ( n34023 , n34021 , n34022 );
nor ( n34024 , n34020 , n34023 );
not ( n34025 , n34024 );
or ( n34026 , n34016 , n34025 );
or ( n34027 , n34015 , n34024 );
nand ( n34028 , n34026 , n34027 );
buf ( n34029 , RI173fd738_1520);
not ( n34030 , n34029 );
not ( n34031 , RI173b4700_1876);
not ( n34032 , n34031 );
or ( n34033 , n34030 , n34032 );
not ( n34034 , RI173fd738_1520);
buf ( n34035 , RI173b4700_1876);
nand ( n34036 , n34034 , n34035 );
nand ( n34037 , n34033 , n34036 );
buf ( n34038 , RI173b4a48_1875);
and ( n34039 , n34037 , n34038 );
not ( n34040 , n34037 );
not ( n34041 , RI173b4a48_1875);
and ( n34042 , n34040 , n34041 );
nor ( n34043 , n34039 , n34042 );
not ( n34044 , n34043 );
xor ( n211806 , n34028 , n34044 );
buf ( n211807 , n211806 );
not ( n34047 , n211807 );
or ( n34048 , n34007 , n34047 );
not ( n34049 , n204869 );
xor ( n34050 , n34043 , n34015 );
xnor ( n34051 , n34050 , n34024 );
nand ( n34052 , n34049 , n34051 );
nand ( n34053 , n34048 , n34052 );
buf ( n34054 , RI173d1f98_1732);
not ( n34055 , n34054 );
not ( n34056 , RI173599e0_2088);
not ( n34057 , n34056 );
or ( n34058 , n34055 , n34057 );
not ( n34059 , RI173d1f98_1732);
buf ( n34060 , RI173599e0_2088);
nand ( n34061 , n34059 , n34060 );
nand ( n34062 , n34058 , n34061 );
not ( n34063 , RI17449a70_1377);
and ( n34064 , n34062 , n34063 );
not ( n34065 , n34062 );
buf ( n34066 , RI17449a70_1377);
and ( n34067 , n34065 , n34066 );
nor ( n34068 , n34064 , n34067 );
buf ( n34069 , RI19a894c8_2729);
nand ( n34070 , n25793 , n34069 );
buf ( n34071 , RI1746e280_1199);
and ( n34072 , n34070 , n34071 );
not ( n34073 , n34070 );
not ( n34074 , RI1746e280_1199);
and ( n34075 , n34073 , n34074 );
nor ( n34076 , n34072 , n34075 );
not ( n34077 , n34076 );
xor ( n34078 , n34068 , n34077 );
buf ( n34079 , RI19abaf50_2374);
nand ( n34080 , n28997 , n34079 );
not ( n34081 , RI174b6f58_844);
and ( n34082 , n34080 , n34081 );
not ( n34083 , n34080 );
buf ( n34084 , RI174b6f58_844);
and ( n34085 , n34083 , n34084 );
nor ( n34086 , n34082 , n34085 );
buf ( n34087 , n34086 );
xnor ( n34088 , n34078 , n34087 );
buf ( n34089 , n34088 );
buf ( n34090 , n34089 );
and ( n34091 , n34053 , n34090 );
not ( n34092 , n34053 );
not ( n34093 , n34076 );
not ( n34094 , n34086 );
or ( n34095 , n34093 , n34094 );
or ( n34096 , n34076 , n34086 );
nand ( n34097 , n34095 , n34096 );
and ( n34098 , n34097 , n34068 );
not ( n34099 , n34097 );
not ( n34100 , n34068 );
and ( n34101 , n34099 , n34100 );
nor ( n34102 , n34098 , n34101 );
buf ( n34103 , n34102 );
buf ( n34104 , n34103 );
and ( n34105 , n34092 , n34104 );
nor ( n34106 , n34091 , n34105 );
nand ( n34107 , n34006 , n34106 );
not ( n34108 , n34107 );
not ( n34109 , n33176 );
not ( n34110 , n28251 );
or ( n34111 , n34109 , n34110 );
or ( n34112 , n28251 , n33176 );
nand ( n34113 , n34111 , n34112 );
not ( n34114 , n34113 );
buf ( n34115 , n28288 );
not ( n34116 , n34115 );
and ( n34117 , n34114 , n34116 );
and ( n34118 , n34113 , n34115 );
nor ( n34119 , n34117 , n34118 );
not ( n34120 , n34119 );
not ( n34121 , n34120 );
and ( n34122 , n34108 , n34121 );
and ( n34123 , n34107 , n34120 );
nor ( n34124 , n34122 , n34123 );
not ( n34125 , n34124 );
not ( n34126 , n34125 );
or ( n34127 , n33967 , n34126 );
nand ( n34128 , n34124 , n33965 );
nand ( n34129 , n34127 , n34128 );
buf ( n34130 , RI19abcbe8_2361);
nand ( n34131 , n25451 , n34130 );
buf ( n34132 , RI174b6238_848);
and ( n34133 , n34131 , n34132 );
not ( n34134 , n34131 );
not ( n34135 , RI174b6238_848);
and ( n34136 , n34134 , n34135 );
nor ( n34137 , n34133 , n34136 );
buf ( n34138 , n34137 );
buf ( n34139 , n208398 );
or ( n34140 , n34138 , n34139 );
not ( n34141 , n30638 );
nand ( n34142 , n34141 , n34138 );
nand ( n34143 , n34140 , n34142 );
not ( n34144 , n34143 );
buf ( n34145 , RI173dfb70_1665);
not ( n34146 , n34145 );
not ( n34147 , RI17396e80_2020);
not ( n34148 , n34147 );
or ( n34149 , n34146 , n34148 );
not ( n34150 , RI173dfb70_1665);
buf ( n34151 , RI17396e80_2020);
nand ( n34152 , n34150 , n34151 );
nand ( n34153 , n34149 , n34152 );
buf ( n34154 , RI17457648_1310);
and ( n34155 , n34153 , n34154 );
not ( n34156 , n34153 );
not ( n34157 , RI17457648_1310);
and ( n34158 , n34156 , n34157 );
nor ( n34159 , n34155 , n34158 );
buf ( n34160 , RI19a95930_2643);
nand ( n34161 , n25479 , n34160 );
buf ( n34162 , RI1747c1a0_1131);
and ( n34163 , n34161 , n34162 );
not ( n34164 , n34161 );
not ( n34165 , RI1747c1a0_1131);
and ( n34166 , n34164 , n34165 );
nor ( n34167 , n34163 , n34166 );
xor ( n34168 , n34159 , n34167 );
buf ( n34169 , RI19ac5720_2288);
nand ( n34170 , n25880 , n34169 );
not ( n34171 , RI174cbf70_776);
and ( n34172 , n34170 , n34171 );
not ( n34173 , n34170 );
buf ( n34174 , RI174cbf70_776);
and ( n34175 , n34173 , n34174 );
nor ( n34176 , n34172 , n34175 );
xor ( n34177 , n34168 , n34176 );
not ( n34178 , n34177 );
not ( n34179 , n34178 );
buf ( n34180 , n34179 );
not ( n34181 , n34180 );
and ( n34182 , n34144 , n34181 );
and ( n34183 , n34143 , n34180 );
nor ( n34184 , n34182 , n34183 );
buf ( n34185 , RI17390f58_2049);
not ( n34186 , n34185 );
not ( n34187 , n33657 );
or ( n34188 , n34186 , n34187 );
not ( n34189 , n34185 );
xor ( n34190 , n33638 , n33646 );
xnor ( n34191 , n34190 , n33656 );
nand ( n34192 , n34189 , n34191 );
nand ( n34193 , n34188 , n34192 );
buf ( n34194 , RI173e8888_1622);
not ( n34195 , n34194 );
not ( n34196 , RI1739f850_1978);
not ( n34197 , n34196 );
or ( n34198 , n34195 , n34197 );
not ( n34199 , RI173e8888_1622);
buf ( n34200 , RI1739f850_1978);
nand ( n34201 , n34199 , n34200 );
and ( n34202 , n34198 , n34201 );
buf ( n34203 , RI17460360_1267);
and ( n34204 , n34202 , n34203 );
not ( n34205 , n34202 );
not ( n34206 , RI17460360_1267);
and ( n34207 , n34205 , n34206 );
nor ( n34208 , n34204 , n34207 );
buf ( n34209 , RI19aa27e8_2549);
nand ( n34210 , n204512 , n34209 );
buf ( n34211 , RI17484b70_1089);
and ( n34212 , n34210 , n34211 );
not ( n34213 , n34210 );
not ( n34214 , RI17484b70_1089);
and ( n34215 , n34213 , n34214 );
nor ( n34216 , n34212 , n34215 );
or ( n34217 , n34208 , n34216 );
xnor ( n34218 , n34217 , n32106 );
not ( n34219 , n34218 );
not ( n34220 , n34219 );
and ( n34221 , n34193 , n34220 );
not ( n34222 , n34193 );
xor ( n34223 , n34208 , n32105 );
not ( n34224 , n34216 );
xor ( n34225 , n34223 , n34224 );
not ( n34226 , n34225 );
not ( n34227 , n34226 );
and ( n34228 , n34222 , n34227 );
nor ( n34229 , n34221 , n34228 );
nand ( n34230 , n34184 , n34229 );
buf ( n34231 , RI173cf4d8_1745);
not ( n34232 , n34231 );
not ( n34233 , RI17345c10_2101);
not ( n34234 , n34233 );
or ( n34235 , n34232 , n34234 );
not ( n34236 , RI173cf4d8_1745);
buf ( n34237 , RI17345c10_2101);
nand ( n34238 , n34236 , n34237 );
nand ( n34239 , n34235 , n34238 );
buf ( n34240 , RI17446fc8_1390);
and ( n34241 , n34239 , n34240 );
not ( n34242 , n34239 );
not ( n34243 , RI17446fc8_1390);
and ( n34244 , n34242 , n34243 );
nor ( n34245 , n34241 , n34244 );
buf ( n34246 , RI19a8c948_2707);
nand ( n34247 , n25751 , n34246 );
not ( n34248 , RI1746b7d8_1212);
and ( n34249 , n34247 , n34248 );
not ( n34250 , n34247 );
buf ( n34251 , RI1746b7d8_1212);
and ( n34252 , n34250 , n34251 );
nor ( n34253 , n34249 , n34252 );
or ( n34254 , n34245 , n34253 );
buf ( n212016 , RI19abdbd8_2352);
nand ( n212017 , n204393 , n212016 );
not ( n34257 , RI174b44b0_857);
and ( n212019 , n212017 , n34257 );
not ( n212020 , n212017 );
buf ( n34260 , RI174b44b0_857);
and ( n34261 , n212020 , n34260 );
nor ( n34262 , n212019 , n34261 );
or ( n34263 , n34254 , n34262 );
buf ( n34264 , n34263 );
not ( n34265 , n34264 );
not ( n34266 , n34265 );
buf ( n34267 , n31761 );
not ( n34268 , n34267 );
not ( n34269 , n210247 );
not ( n34270 , RI173b1c58_1889);
not ( n34271 , n34270 );
or ( n34272 , n34269 , n34271 );
not ( n34273 , RI173fa948_1534);
nand ( n34274 , n34273 , n29744 );
nand ( n34275 , n34272 , n34274 );
buf ( n34276 , RI173995e0_2008);
and ( n34277 , n34275 , n34276 );
not ( n34278 , n34275 );
not ( n34279 , RI173995e0_2008);
and ( n34280 , n34278 , n34279 );
nor ( n34281 , n34277 , n34280 );
buf ( n34282 , RI19a9fcc8_2570);
nand ( n34283 , n25656 , n34282 );
buf ( n34284 , RI17526f78_645);
and ( n34285 , n34283 , n34284 );
not ( n34286 , n34283 );
not ( n34287 , RI17526f78_645);
and ( n34288 , n34286 , n34287 );
nor ( n34289 , n34285 , n34288 );
xor ( n34290 , n34281 , n34289 );
buf ( n34291 , RI19aaa150_2495);
nand ( n34292 , n25405 , n34291 );
buf ( n34293 , RI17496f78_1000);
and ( n34294 , n34292 , n34293 );
not ( n34295 , n34292 );
not ( n34296 , RI17496f78_1000);
and ( n34297 , n34295 , n34296 );
nor ( n34298 , n34294 , n34297 );
xnor ( n34299 , n34290 , n34298 );
not ( n34300 , n34299 );
or ( n34301 , n34268 , n34300 );
not ( n34302 , n34267 );
not ( n34303 , n34299 );
nand ( n34304 , n34302 , n34303 );
nand ( n34305 , n34301 , n34304 );
not ( n34306 , n34305 );
or ( n34307 , n34266 , n34306 );
not ( n34308 , n34264 );
or ( n34309 , n34305 , n34308 );
nand ( n34310 , n34307 , n34309 );
not ( n34311 , n34310 );
and ( n34312 , n34230 , n34311 );
not ( n34313 , n34230 );
and ( n34314 , n34313 , n34310 );
nor ( n34315 , n34312 , n34314 );
not ( n34316 , n34315 );
and ( n34317 , n34129 , n34316 );
not ( n34318 , n34129 );
and ( n34319 , n34318 , n34315 );
nor ( n34320 , n34317 , n34319 );
buf ( n34321 , RI173358d8_2180);
not ( n34322 , n34321 );
not ( n34323 , n25762 );
or ( n34324 , n34322 , n34323 );
not ( n34325 , n34321 );
and ( n34326 , n34325 , n25765 );
nand ( n34327 , n34324 , n34326 );
not ( n34328 , n25722 );
nand ( n34329 , n34327 , n34328 );
not ( n34330 , n34327 );
buf ( n34331 , n25771 );
nand ( n34332 , n34330 , n34331 );
nor ( n34333 , n34329 , n34332 );
not ( n34334 , n34333 );
not ( n34335 , n32863 );
not ( n34336 , n34335 );
xor ( n34337 , n31326 , n31335 );
xnor ( n34338 , n34337 , n31342 );
not ( n34339 , n34338 );
not ( n34340 , n34339 );
not ( n34341 , n28435 );
and ( n34342 , n34340 , n34341 );
and ( n34343 , n31344 , n28435 );
nor ( n34344 , n34342 , n34343 );
not ( n34345 , n34344 );
and ( n34346 , n34336 , n34345 );
and ( n34347 , n34335 , n34344 );
nor ( n34348 , n34346 , n34347 );
not ( n34349 , n34348 );
nand ( n34350 , n34334 , n34349 );
not ( n34351 , n34350 );
buf ( n34352 , RI17409c18_1460);
not ( n34353 , n34352 );
not ( n34354 , RI173c0f28_1815);
not ( n34355 , n34354 );
or ( n34356 , n34353 , n34355 );
not ( n34357 , RI17409c18_1460);
buf ( n34358 , RI173c0f28_1815);
nand ( n34359 , n34357 , n34358 );
nand ( n34360 , n34356 , n34359 );
not ( n34361 , n34360 );
buf ( n34362 , RI173379a8_2170);
not ( n34363 , RI1745e920_1275);
xor ( n34364 , n34362 , n34363 );
buf ( n34365 , RI174a6248_926);
not ( n34366 , n34365 );
buf ( n34367 , RI19ab4560_2421);
nand ( n34368 , n25751 , n34367 );
not ( n34369 , n34368 );
or ( n34370 , n34366 , n34369 );
nand ( n34371 , n30356 , n34367 );
or ( n34372 , n34371 , n34365 );
nand ( n34373 , n34370 , n34372 );
xnor ( n34374 , n34364 , n34373 );
not ( n34375 , n34374 );
not ( n34376 , n34375 );
or ( n34377 , n34361 , n34376 );
not ( n34378 , n34360 );
nand ( n34379 , n34374 , n34378 );
nand ( n34380 , n34377 , n34379 );
buf ( n34381 , n34380 );
not ( n34382 , n34381 );
not ( n34383 , n34382 );
not ( n34384 , n205321 );
nor ( n34385 , n34384 , n28775 );
not ( n34386 , n34385 );
nand ( n34387 , n28775 , n34384 );
nand ( n34388 , n34386 , n34387 );
not ( n34389 , n34388 );
or ( n34390 , n34383 , n34389 );
not ( n34391 , n34381 );
or ( n34392 , n34388 , n34391 );
nand ( n34393 , n34390 , n34392 );
not ( n34394 , n34393 );
and ( n34395 , n34351 , n34394 );
and ( n34396 , n34350 , n34393 );
nor ( n34397 , n34395 , n34396 );
not ( n34398 , n34397 );
not ( n34399 , n34398 );
not ( n34400 , n33721 );
nand ( n34401 , n33861 , n34400 );
buf ( n34402 , RI19a8faf8_2685);
nand ( n34403 , n204426 , n34402 );
buf ( n34404 , RI17465220_1243);
and ( n34405 , n34403 , n34404 );
not ( n34406 , n34403 );
not ( n34407 , RI17465220_1243);
and ( n34408 , n34406 , n34407 );
nor ( n34409 , n34405 , n34408 );
buf ( n34410 , n34409 );
not ( n34411 , n34410 );
buf ( n34412 , RI173eda90_1597);
xor ( n34413 , n34412 , n204567 );
not ( n34414 , n204584 );
xnor ( n34415 , n34413 , n34414 );
buf ( n34416 , n34415 );
not ( n34417 , n34416 );
or ( n34418 , n34411 , n34417 );
or ( n34419 , n34416 , n34410 );
nand ( n34420 , n34418 , n34419 );
and ( n34421 , n34420 , n204632 );
not ( n34422 , n34420 );
and ( n34423 , n34422 , n204622 );
nor ( n34424 , n34421 , n34423 );
not ( n34425 , n34424 );
and ( n34426 , n34401 , n34425 );
not ( n34427 , n34401 );
and ( n34428 , n34427 , n34424 );
nor ( n34429 , n34426 , n34428 );
not ( n34430 , n34429 );
not ( n34431 , n34430 );
or ( n34432 , n34399 , n34431 );
nand ( n34433 , n34429 , n34397 );
nand ( n34434 , n34432 , n34433 );
and ( n34435 , n34320 , n34434 );
not ( n34436 , n34320 );
not ( n34437 , n34434 );
and ( n34438 , n34436 , n34437 );
nor ( n34439 , n34435 , n34438 );
not ( n34440 , n34439 );
or ( n34441 , n33867 , n34440 );
not ( n34442 , n33866 );
not ( n34443 , n34437 );
not ( n34444 , n34320 );
not ( n34445 , n34444 );
or ( n34446 , n34443 , n34445 );
nand ( n34447 , n34320 , n34434 );
nand ( n34448 , n34446 , n34447 );
nand ( n34449 , n34442 , n34448 );
nand ( n34450 , n34441 , n34449 );
not ( n34451 , n34450 );
or ( n34452 , n33710 , n34451 );
or ( n34453 , n34450 , n33709 );
nand ( n34454 , n34452 , n34453 );
not ( n34455 , n34454 );
not ( n34456 , n207190 );
not ( n34457 , n33404 );
or ( n34458 , n34456 , n34457 );
or ( n34459 , n33404 , n207190 );
nand ( n34460 , n34458 , n34459 );
buf ( n34461 , n205236 );
and ( n34462 , n34460 , n34461 );
not ( n34463 , n34460 );
not ( n34464 , n25826 );
and ( n34465 , n34463 , n34464 );
nor ( n34466 , n34462 , n34465 );
not ( n34467 , n30220 );
not ( n34468 , n205173 );
not ( n34469 , n34468 );
not ( n34470 , n204436 );
or ( n34471 , n34469 , n34470 );
nand ( n34472 , n204439 , n205173 );
nand ( n34473 , n34471 , n34472 );
not ( n34474 , n34473 );
or ( n34475 , n34467 , n34474 );
not ( n34476 , n30220 );
not ( n34477 , n34476 );
or ( n34478 , n34473 , n34477 );
nand ( n212240 , n34475 , n34478 );
nand ( n212241 , n34466 , n212240 );
not ( n34481 , n212241 );
buf ( n34482 , RI1740a5f0_1457);
not ( n34483 , n34482 );
buf ( n34484 , RI173fc040_1527);
not ( n34485 , n34484 );
not ( n34486 , RI173b3008_1883);
not ( n34487 , n34486 );
or ( n34488 , n34485 , n34487 );
not ( n34489 , RI173fc040_1527);
buf ( n34490 , RI173b3008_1883);
nand ( n34491 , n34489 , n34490 );
nand ( n34492 , n34488 , n34491 );
not ( n34493 , RI173a4da0_1952);
and ( n34494 , n34492 , n34493 );
not ( n34495 , n34492 );
buf ( n34496 , RI173a4da0_1952);
and ( n34497 , n34495 , n34496 );
nor ( n34498 , n34494 , n34497 );
buf ( n34499 , RI19aa8530_2507);
nand ( n34500 , n33787 , n34499 );
buf ( n34501 , RI17498328_994);
and ( n34502 , n34500 , n34501 );
not ( n34503 , n34500 );
not ( n34504 , RI17498328_994);
and ( n34505 , n34503 , n34504 );
nor ( n34506 , n34502 , n34505 );
xor ( n34507 , n34498 , n34506 );
buf ( n34508 , RI19a8eb08_2692);
nand ( n34509 , n204513 , n34508 );
not ( n34510 , RI17528e68_639);
and ( n34511 , n34509 , n34510 );
not ( n34512 , n34509 );
buf ( n34513 , RI17528e68_639);
and ( n34514 , n34512 , n34513 );
nor ( n34515 , n34511 , n34514 );
xnor ( n34516 , n34507 , n34515 );
not ( n34517 , n34516 );
or ( n34518 , n34483 , n34517 );
not ( n34519 , n34482 );
xor ( n34520 , n34498 , n34506 );
xnor ( n34521 , n34520 , n34515 );
not ( n34522 , n34521 );
and ( n34523 , n34519 , n34522 );
and ( n34524 , n34518 , n34523 );
buf ( n34525 , RI173d0888_1739);
not ( n34526 , n34525 );
not ( n34527 , RI17346fc0_2095);
not ( n34528 , n34527 );
or ( n34529 , n34526 , n34528 );
not ( n34530 , RI173d0888_1739);
buf ( n34531 , RI17346fc0_2095);
and ( n34532 , n34530 , n34531 );
and ( n34533 , n34529 , n34532 );
buf ( n34534 , RI17448378_1384);
and ( n34535 , n34533 , n34534 );
not ( n34536 , n34533 );
not ( n34537 , RI17448378_1384);
and ( n34538 , n34536 , n34537 );
nor ( n34539 , n34535 , n34538 );
buf ( n34540 , RI19a8acb0_2719);
nand ( n34541 , n205019 , n34540 );
buf ( n34542 , RI1746cb88_1206);
and ( n34543 , n34541 , n34542 );
not ( n34544 , n34541 );
not ( n34545 , RI1746cb88_1206);
and ( n34546 , n34544 , n34545 );
nor ( n34547 , n34543 , n34546 );
xor ( n34548 , n34539 , n34547 );
buf ( n34549 , RI19abc6c0_2364);
nand ( n34550 , n205271 , n34549 );
not ( n34551 , RI174b5860_851);
and ( n34552 , n34550 , n34551 );
not ( n34553 , n34550 );
buf ( n34554 , RI174b5860_851);
and ( n34555 , n34553 , n34554 );
nor ( n34556 , n34552 , n34555 );
xnor ( n34557 , n34548 , n34556 );
buf ( n34558 , n34557 );
and ( n34559 , n34524 , n34558 );
not ( n34560 , n34524 );
not ( n34561 , n34547 );
xor ( n34562 , n34539 , n34561 );
xnor ( n34563 , n34562 , n34556 );
buf ( n34564 , n34563 );
and ( n34565 , n34560 , n34564 );
nor ( n34566 , n34559 , n34565 );
not ( n34567 , n34566 );
and ( n34568 , n34481 , n34567 );
and ( n34569 , n212241 , n34566 );
nor ( n34570 , n34568 , n34569 );
not ( n34571 , n34570 );
not ( n34572 , n34571 );
buf ( n34573 , RI1733fce8_2130);
not ( n34574 , n34573 );
not ( n34575 , n32441 );
not ( n34576 , n34575 );
or ( n34577 , n34574 , n34576 );
not ( n34578 , n34573 );
nand ( n34579 , n34578 , n32441 );
nand ( n34580 , n34577 , n34579 );
not ( n34581 , n34580 );
not ( n34582 , n26222 );
and ( n34583 , n34581 , n34582 );
and ( n34584 , n26222 , n34580 );
nor ( n34585 , n34583 , n34584 );
not ( n34586 , n34585 );
buf ( n34587 , RI173eee40_1591);
not ( n34588 , n34587 );
not ( n34589 , n207493 );
not ( n34590 , n34589 );
or ( n34591 , n34588 , n34590 );
or ( n34592 , n29733 , n34587 );
nand ( n34593 , n34591 , n34592 );
not ( n34594 , n33444 );
and ( n34595 , n34593 , n34594 );
not ( n34596 , n34593 );
not ( n34597 , n33444 );
not ( n34598 , n34597 );
and ( n34599 , n34596 , n34598 );
nor ( n34600 , n34595 , n34599 );
not ( n34601 , n34600 );
nand ( n34602 , n34586 , n34601 );
not ( n34603 , n30689 );
not ( n34604 , n34603 );
buf ( n34605 , RI173964a8_2023);
not ( n34606 , n34605 );
not ( n34607 , n33134 );
or ( n34608 , n34606 , n34607 );
or ( n34609 , n33134 , n34605 );
nand ( n34610 , n34608 , n34609 );
not ( n34611 , n34610 );
or ( n34612 , n34604 , n34611 );
buf ( n34613 , n30685 );
or ( n34614 , n34610 , n34613 );
nand ( n34615 , n34612 , n34614 );
buf ( n34616 , n34615 );
not ( n34617 , n34616 );
and ( n34618 , n34602 , n34617 );
not ( n34619 , n34602 );
and ( n34620 , n34619 , n34616 );
nor ( n34621 , n34618 , n34620 );
not ( n34622 , n34621 );
not ( n34623 , n34622 );
not ( n34624 , n34566 );
not ( n34625 , n34466 );
nand ( n34626 , n34624 , n34625 );
not ( n34627 , n34626 );
not ( n34628 , RI173cdde0_1752);
not ( n34629 , RI174001e0_1507);
buf ( n34630 , RI173b74f0_1862);
and ( n34631 , n34629 , n34630 );
not ( n34632 , n34629 );
not ( n34633 , RI173b74f0_1862);
and ( n34634 , n34632 , n34633 );
nor ( n34635 , n34631 , n34634 );
xor ( n34636 , n34628 , n34635 );
buf ( n34637 , RI1752f588_619);
buf ( n34638 , RI1749c4c8_974);
xor ( n34639 , n34637 , n34638 );
buf ( n34640 , RI19aba050_2380);
nand ( n34641 , n26325 , n34640 );
xnor ( n34642 , n34639 , n34641 );
xnor ( n34643 , n34636 , n34642 );
not ( n34644 , n34643 );
not ( n34645 , n34644 );
not ( n34646 , n34645 );
not ( n34647 , n31802 );
not ( n212409 , n27759 );
or ( n212410 , n34647 , n212409 );
nand ( n34650 , n27758 , n31798 );
nand ( n34651 , n212410 , n34650 );
not ( n34652 , n34651 );
and ( n34653 , n34646 , n34652 );
buf ( n34654 , n34643 );
and ( n34655 , n34654 , n34651 );
nor ( n34656 , n34653 , n34655 );
not ( n34657 , n34656 );
not ( n34658 , n34657 );
and ( n34659 , n34627 , n34658 );
and ( n34660 , n34626 , n34657 );
nor ( n34661 , n34659 , n34660 );
not ( n34662 , n34661 );
not ( n34663 , n34662 );
or ( n34664 , n34623 , n34663 );
nand ( n34665 , n34661 , n34621 );
nand ( n34666 , n34664 , n34665 );
buf ( n34667 , RI173d1c50_1733);
not ( n34668 , n34667 );
not ( n34669 , RI17359698_2089);
not ( n34670 , n34669 );
or ( n34671 , n34668 , n34670 );
not ( n34672 , RI173d1c50_1733);
buf ( n34673 , RI17359698_2089);
nand ( n34674 , n34672 , n34673 );
nand ( n34675 , n34671 , n34674 );
not ( n34676 , RI17449728_1378);
and ( n34677 , n34675 , n34676 );
not ( n34678 , n34675 );
buf ( n34679 , RI17449728_1378);
and ( n34680 , n34678 , n34679 );
nor ( n34681 , n34677 , n34680 );
buf ( n34682 , RI19a89270_2730);
nand ( n34683 , n33787 , n34682 );
buf ( n34684 , RI1746df38_1200);
and ( n34685 , n34683 , n34684 );
not ( n34686 , n34683 );
not ( n34687 , RI1746df38_1200);
and ( n34688 , n34686 , n34687 );
nor ( n34689 , n34685 , n34688 );
xor ( n34690 , n34681 , n34689 );
buf ( n34691 , RI19abad70_2375);
nand ( n34692 , n204426 , n34691 );
not ( n34693 , RI174b6c10_845);
and ( n34694 , n34692 , n34693 );
not ( n34695 , n34692 );
buf ( n34696 , RI174b6c10_845);
and ( n34697 , n34695 , n34696 );
nor ( n34698 , n34694 , n34697 );
xnor ( n34699 , n34690 , n34698 );
buf ( n34700 , n34699 );
xor ( n34701 , n29666 , n34700 );
buf ( n34702 , RI173fd3f0_1521);
not ( n34703 , n34702 );
not ( n34704 , RI173b43b8_1877);
not ( n34705 , n34704 );
or ( n34706 , n34703 , n34705 );
not ( n34707 , RI173fd3f0_1521);
buf ( n34708 , RI173b43b8_1877);
nand ( n34709 , n34707 , n34708 );
nand ( n34710 , n34706 , n34709 );
not ( n34711 , n34710 );
buf ( n34712 , RI19a87dd0_2739);
nand ( n34713 , n25529 , n34712 );
buf ( n34714 , RI1752ad58_633);
and ( n34715 , n34713 , n34714 );
not ( n34716 , n34713 );
not ( n34717 , RI1752ad58_633);
and ( n34718 , n34716 , n34717 );
nor ( n34719 , n34715 , n34718 );
xor ( n34720 , n204862 , n34719 );
buf ( n34721 , RI19aa6b68_2518);
nand ( n34722 , n25583 , n34721 );
buf ( n34723 , RI174996d8_988);
and ( n34724 , n34722 , n34723 );
not ( n34725 , n34722 );
not ( n34726 , RI174996d8_988);
and ( n34727 , n34725 , n34726 );
nor ( n34728 , n34724 , n34727 );
xnor ( n34729 , n34720 , n34728 );
not ( n34730 , n34729 );
or ( n34731 , n34711 , n34730 );
not ( n34732 , n34729 );
not ( n34733 , n34710 );
nand ( n34734 , n34732 , n34733 );
nand ( n34735 , n34731 , n34734 );
not ( n34736 , n34735 );
xnor ( n34737 , n34701 , n34736 );
not ( n34738 , n27891 );
not ( n34739 , n33777 );
or ( n34740 , n34738 , n34739 );
or ( n34741 , n33777 , n27891 );
nand ( n34742 , n34740 , n34741 );
xor ( n34743 , n34742 , n33807 );
xnor ( n34744 , n34743 , n209733 );
buf ( n34745 , n34744 );
or ( n34746 , n34737 , n34745 );
not ( n34747 , n205106 );
not ( n34748 , n32570 );
or ( n34749 , n34747 , n34748 );
nand ( n34750 , n32547 , n205102 );
nand ( n34751 , n34749 , n34750 );
not ( n34752 , n34751 );
not ( n34753 , n32566 );
not ( n34754 , n34753 );
or ( n34755 , n34752 , n34754 );
or ( n34756 , n34753 , n34751 );
nand ( n34757 , n34755 , n34756 );
not ( n34758 , n32607 );
not ( n34759 , n34758 );
and ( n34760 , n34757 , n34759 );
not ( n34761 , n34757 );
xor ( n34762 , n32588 , n210366 );
xnor ( n34763 , n34762 , n32596 );
and ( n34764 , n34761 , n34763 );
nor ( n34765 , n34760 , n34764 );
and ( n34766 , n34746 , n34765 );
not ( n34767 , n34746 );
not ( n34768 , n34765 );
and ( n34769 , n34767 , n34768 );
nor ( n34770 , n34766 , n34769 );
and ( n34771 , n34666 , n34770 );
not ( n34772 , n34666 );
not ( n34773 , n34770 );
and ( n34774 , n34772 , n34773 );
nor ( n34775 , n34771 , n34774 );
buf ( n34776 , RI173c9f88_1771);
not ( n34777 , n34776 );
not ( n34778 , RI17340a08_2126);
not ( n34779 , n34778 );
or ( n34780 , n34777 , n34779 );
not ( n34781 , RI173c9f88_1771);
nand ( n34782 , n34781 , n29100 );
nand ( n34783 , n34780 , n34782 );
not ( n34784 , RI17412fc0_1415);
and ( n34785 , n34783 , n34784 );
not ( n34786 , n34783 );
buf ( n34787 , RI17412fc0_1415);
and ( n34788 , n34786 , n34787 );
nor ( n34789 , n34785 , n34788 );
buf ( n34790 , RI19ac0d88_2324);
nand ( n34791 , n25539 , n34790 );
buf ( n34792 , RI174af2a8_882);
and ( n34793 , n34791 , n34792 );
not ( n34794 , n34791 );
not ( n34795 , RI174af2a8_882);
and ( n34796 , n34794 , n34795 );
nor ( n34797 , n34793 , n34796 );
xor ( n34798 , n34789 , n34797 );
buf ( n34799 , RI19a90818_2679);
nand ( n34800 , n25793 , n34799 );
not ( n34801 , RI174665d0_1237);
and ( n34802 , n34800 , n34801 );
not ( n34803 , n34800 );
buf ( n34804 , RI174665d0_1237);
and ( n34805 , n34803 , n34804 );
nor ( n34806 , n34802 , n34805 );
xnor ( n34807 , n34798 , n34806 );
not ( n34808 , n34807 );
not ( n34809 , n33286 );
and ( n34810 , n34808 , n34809 );
and ( n34811 , n34807 , n33286 );
nor ( n34812 , n34810 , n34811 );
and ( n34813 , n34812 , n26051 );
not ( n34814 , n34812 );
and ( n34815 , n34814 , n26050 );
nor ( n34816 , n34813 , n34815 );
buf ( n34817 , n34816 );
not ( n34818 , n34817 );
xor ( n34819 , n207040 , n29288 );
xnor ( n34820 , n34819 , n29297 );
xor ( n34821 , n33731 , n34820 );
not ( n34822 , n33204 );
not ( n34823 , n33225 );
or ( n34824 , n34822 , n34823 );
nand ( n34825 , n34824 , n33228 );
xnor ( n34826 , n34821 , n34825 );
not ( n34827 , n34826 );
nand ( n34828 , n34818 , n34827 );
not ( n34829 , n34828 );
and ( n34830 , n31773 , n205249 );
not ( n34831 , n31773 );
and ( n34832 , n34831 , n205253 );
nor ( n34833 , n34830 , n34832 );
not ( n34834 , n34833 );
not ( n34835 , n34834 );
not ( n34836 , n31763 );
or ( n34837 , n34835 , n34836 );
nand ( n34838 , n31762 , n34833 );
nand ( n34839 , n34837 , n34838 );
buf ( n34840 , RI173ddde8_1674);
not ( n212602 , n34840 );
not ( n212603 , RI173950f8_2029);
not ( n34843 , n212603 );
or ( n34844 , n212602 , n34843 );
not ( n34845 , RI173ddde8_1674);
buf ( n34846 , RI173950f8_2029);
nand ( n34847 , n34845 , n34846 );
nand ( n34848 , n34844 , n34847 );
buf ( n34849 , RI174558c0_1319);
and ( n34850 , n34848 , n34849 );
not ( n34851 , n34848 );
not ( n34852 , RI174558c0_1319);
and ( n34853 , n34851 , n34852 );
nor ( n34854 , n34850 , n34853 );
buf ( n34855 , RI19a96bf0_2635);
nand ( n34856 , n26028 , n34855 );
buf ( n34857 , RI1747a418_1140);
and ( n34858 , n34856 , n34857 );
not ( n34859 , n34856 );
not ( n212621 , RI1747a418_1140);
and ( n212622 , n34859 , n212621 );
nor ( n212623 , n34858 , n212622 );
xor ( n212624 , n34854 , n212623 );
buf ( n34864 , RI19ac69e0_2280);
nand ( n34865 , n28238 , n34864 );
not ( n34866 , RI174c9108_785);
and ( n34867 , n34865 , n34866 );
not ( n34868 , n34865 );
buf ( n34869 , RI174c9108_785);
and ( n34870 , n34868 , n34869 );
nor ( n34871 , n34867 , n34870 );
xnor ( n34872 , n212624 , n34871 );
not ( n34873 , n34872 );
and ( n34874 , n34839 , n34873 );
not ( n34875 , n34839 );
not ( n34876 , n34873 );
and ( n34877 , n34875 , n34876 );
nor ( n34878 , n34874 , n34877 );
not ( n34879 , n34878 );
not ( n34880 , n34879 );
and ( n34881 , n34829 , n34880 );
and ( n34882 , n34828 , n34879 );
nor ( n34883 , n34881 , n34882 );
not ( n34884 , n34883 );
not ( n34885 , n31020 );
not ( n34886 , n28288 );
or ( n34887 , n34885 , n34886 );
or ( n34888 , n28288 , n31020 );
nand ( n34889 , n34887 , n34888 );
buf ( n34890 , RI173c8bd8_1777);
not ( n34891 , n34890 );
not ( n34892 , RI1733f658_2132);
not ( n34893 , n34892 );
or ( n34894 , n34891 , n34893 );
not ( n34895 , RI173c8bd8_1777);
buf ( n34896 , RI1733f658_2132);
nand ( n34897 , n34895 , n34896 );
nand ( n34898 , n34894 , n34897 );
and ( n34899 , n34898 , n204556 );
not ( n34900 , n34898 );
not ( n34901 , RI174118c8_1422);
and ( n34902 , n34900 , n34901 );
nor ( n34903 , n34899 , n34902 );
buf ( n34904 , RI19ac0338_2330);
nand ( n34905 , n25405 , n34904 );
buf ( n34906 , RI174adef8_888);
and ( n34907 , n34905 , n34906 );
not ( n34908 , n34905 );
not ( n34909 , RI174adef8_888);
and ( n34910 , n34908 , n34909 );
nor ( n34911 , n34907 , n34910 );
xor ( n34912 , n34903 , n34911 );
xnor ( n34913 , n34912 , n34409 );
buf ( n34914 , n34913 );
and ( n34915 , n34889 , n34914 );
not ( n34916 , n34889 );
not ( n34917 , n34914 );
and ( n34918 , n34916 , n34917 );
nor ( n34919 , n34915 , n34918 );
not ( n34920 , n34919 );
not ( n34921 , n34920 );
not ( n34922 , n28121 );
not ( n34923 , n30118 );
not ( n34924 , n28070 );
xor ( n34925 , n34923 , n34924 );
nand ( n34926 , n28071 , n30122 );
nand ( n34927 , n34925 , n34926 );
not ( n34928 , n34927 );
or ( n34929 , n34922 , n34928 );
or ( n34930 , n34927 , n28122 );
nand ( n34931 , n34929 , n34930 );
not ( n34932 , n34931 );
buf ( n34933 , RI17454ee8_1322);
not ( n34934 , n34933 );
not ( n34935 , n25550 );
or ( n34936 , n34934 , n34935 );
not ( n34937 , RI17454ee8_1322);
nand ( n34938 , n209690 , n34937 );
nand ( n34939 , n34936 , n34938 );
not ( n34940 , n207506 );
xnor ( n34941 , n34939 , n34940 );
not ( n34942 , n34941 );
nand ( n34943 , n34932 , n34942 );
not ( n34944 , n34943 );
or ( n34945 , n34921 , n34944 );
or ( n34946 , n34943 , n34920 );
nand ( n34947 , n34945 , n34946 );
not ( n34948 , n34947 );
and ( n34949 , n34884 , n34948 );
and ( n34950 , n34883 , n34947 );
nor ( n34951 , n34949 , n34950 );
and ( n34952 , n34775 , n34951 );
not ( n34953 , n34775 );
not ( n34954 , n34951 );
and ( n34955 , n34953 , n34954 );
nor ( n34956 , n34952 , n34955 );
not ( n34957 , n34956 );
or ( n34958 , n34572 , n34957 );
not ( n34959 , n34571 );
not ( n34960 , n34951 );
not ( n34961 , n34775 );
or ( n34962 , n34960 , n34961 );
and ( n34963 , n34666 , n34773 );
not ( n34964 , n34666 );
and ( n34965 , n34964 , n34770 );
nor ( n34966 , n34963 , n34965 );
nand ( n34967 , n34966 , n34954 );
nand ( n34968 , n34962 , n34967 );
nand ( n34969 , n34959 , n34968 );
nand ( n34970 , n34958 , n34969 );
buf ( n34971 , RI17455578_1320);
not ( n34972 , RI17408bb0_1465);
buf ( n34973 , RI173bfec0_1820);
nand ( n34974 , n34972 , n34973 );
not ( n34975 , RI173bfec0_1820);
buf ( n34976 , RI17408bb0_1465);
nand ( n34977 , n34975 , n34976 );
and ( n34978 , n34974 , n34977 );
xor ( n34979 , n34971 , n34978 );
buf ( n34980 , RI174a4e98_932);
xor ( n34981 , n31919 , n34980 );
buf ( n34982 , RI19ab3840_2427);
nand ( n34983 , n205020 , n34982 );
xnor ( n34984 , n34981 , n34983 );
xnor ( n34985 , n34979 , n34984 );
xor ( n34986 , n204434 , n34985 );
not ( n34987 , n25512 );
not ( n34988 , RI17394720_2032);
not ( n34989 , n34988 );
or ( n34990 , n34987 , n34989 );
not ( n34991 , RI173dd410_1677);
buf ( n34992 , RI17394720_2032);
nand ( n34993 , n34991 , n34992 );
nand ( n34994 , n34990 , n34993 );
and ( n34995 , n34994 , n34937 );
not ( n34996 , n34994 );
and ( n34997 , n34996 , n34933 );
nor ( n34998 , n34995 , n34997 );
buf ( n34999 , RI19a964e8_2638);
nand ( n35000 , n204393 , n34999 );
buf ( n35001 , RI17479a40_1143);
and ( n35002 , n35000 , n35001 );
not ( n35003 , n35000 );
not ( n35004 , RI17479a40_1143);
and ( n35005 , n35003 , n35004 );
nor ( n35006 , n35002 , n35005 );
xor ( n35007 , n34998 , n35006 );
buf ( n35008 , RI19ac63c8_2283);
nand ( n35009 , n25851 , n35008 );
buf ( n35010 , RI174c8190_788);
and ( n35011 , n35009 , n35010 );
not ( n35012 , n35009 );
not ( n35013 , RI174c8190_788);
and ( n35014 , n35012 , n35013 );
nor ( n35015 , n35011 , n35014 );
not ( n35016 , n35015 );
xnor ( n35017 , n35007 , n35016 );
xnor ( n35018 , n34986 , n35017 );
not ( n35019 , n35018 );
not ( n35020 , n33274 );
not ( n35021 , n34807 );
not ( n35022 , n35021 );
or ( n35023 , n35020 , n35022 );
or ( n35024 , n35021 , n33274 );
nand ( n35025 , n35023 , n35024 );
and ( n35026 , n35025 , n26047 );
not ( n35027 , n35025 );
not ( n35028 , n26047 );
and ( n35029 , n35027 , n35028 );
nor ( n35030 , n35026 , n35029 );
not ( n35031 , n35030 );
nand ( n35032 , n35019 , n35031 );
not ( n35033 , n204867 );
not ( n35034 , n211806 );
or ( n35035 , n35033 , n35034 );
or ( n35036 , n211806 , n204867 );
nand ( n35037 , n35035 , n35036 );
not ( n35038 , n35037 );
not ( n35039 , n34102 );
and ( n35040 , n35038 , n35039 );
and ( n35041 , n35037 , n34103 );
nor ( n35042 , n35040 , n35041 );
not ( n35043 , n35042 );
xnor ( n35044 , n35032 , n35043 );
not ( n35045 , n35044 );
not ( n35046 , n35045 );
buf ( n35047 , RI173d6e58_1708);
buf ( n35048 , RI173b8210_1858);
not ( n35049 , n35048 );
not ( n35050 , n204678 );
or ( n35051 , n35049 , n35050 );
not ( n35052 , RI173b8210_1858);
nand ( n35053 , n35052 , n204636 );
nand ( n35054 , n35051 , n35053 );
xor ( n35055 , n35047 , n35054 );
buf ( n35056 , RI17530a28_615);
buf ( n35057 , RI1749d1e8_970);
xor ( n35058 , n35056 , n35057 );
buf ( n35059 , RI19ab82c8_2394);
nand ( n35060 , n204426 , n35059 );
xnor ( n35061 , n35058 , n35060 );
not ( n35062 , n35061 );
xnor ( n35063 , n35055 , n35062 );
not ( n35064 , n35063 );
buf ( n35065 , RI1739a990_2002);
not ( n35066 , n35065 );
not ( n35067 , RI173e3680_1647);
not ( n35068 , n35067 );
or ( n35069 , n35066 , n35068 );
not ( n35070 , RI1739a990_2002);
buf ( n35071 , RI173e3680_1647);
nand ( n35072 , n35070 , n35071 );
nand ( n212834 , n35069 , n35072 );
not ( n212835 , RI1745b4a0_1291);
and ( n35075 , n212834 , n212835 );
not ( n35076 , n212834 );
buf ( n35077 , RI1745b4a0_1291);
and ( n35078 , n35076 , n35077 );
nor ( n35079 , n35075 , n35078 );
buf ( n35080 , RI19a87b78_2740);
nand ( n35081 , n25879 , n35080 );
buf ( n35082 , RI17500a58_758);
and ( n35083 , n35081 , n35082 );
not ( n35084 , n35081 );
not ( n35085 , RI17500a58_758);
and ( n35086 , n35084 , n35085 );
nor ( n35087 , n35083 , n35086 );
xor ( n35088 , n35079 , n35087 );
buf ( n35089 , RI19aa6988_2519);
nand ( n35090 , n25583 , n35089 );
not ( n35091 , RI1747fcb0_1113);
and ( n35092 , n35090 , n35091 );
not ( n35093 , n35090 );
buf ( n35094 , RI1747fcb0_1113);
and ( n35095 , n35093 , n35094 );
nor ( n35096 , n35092 , n35095 );
xnor ( n35097 , n35088 , n35096 );
not ( n35098 , n35097 );
not ( n35099 , n35098 );
buf ( n35100 , n30998 );
not ( n35101 , n35100 );
and ( n35102 , n35099 , n35101 );
and ( n35103 , n35098 , n35100 );
nor ( n35104 , n35102 , n35103 );
not ( n35105 , n35104 );
or ( n35106 , n35064 , n35105 );
buf ( n35107 , n35063 );
or ( n35108 , n35107 , n35104 );
nand ( n35109 , n35106 , n35108 );
not ( n35110 , n35109 );
and ( n35111 , n27899 , n204467 );
not ( n35112 , n27899 );
not ( n35113 , RI1733b170_2153);
and ( n35114 , n35112 , n35113 );
nor ( n35115 , n35111 , n35114 );
not ( n35116 , n27921 );
xor ( n35117 , n35115 , n35116 );
xnor ( n35118 , n35117 , n25926 );
not ( n35119 , n35118 );
nand ( n35120 , n35110 , n35119 );
not ( n35121 , n33337 );
not ( n35122 , n30579 );
or ( n35123 , n35121 , n35122 );
or ( n35124 , n30579 , n33337 );
nand ( n35125 , n35123 , n35124 );
buf ( n35126 , RI173b0f38_1893);
not ( n35127 , n35126 );
not ( n35128 , n29010 );
or ( n35129 , n35127 , n35128 );
not ( n35130 , RI173b0f38_1893);
nand ( n35131 , n35130 , n28971 );
nand ( n35132 , n35129 , n35131 );
buf ( n35133 , RI17390580_2052);
and ( n35134 , n35132 , n35133 );
not ( n35135 , n35132 );
not ( n35136 , RI17390580_2052);
and ( n35137 , n35135 , n35136 );
nor ( n35138 , n35134 , n35137 );
buf ( n35139 , RI19a99ad0_2614);
nand ( n35140 , n25741 , n35139 );
buf ( n35141 , RI17525ad8_649);
and ( n35142 , n35140 , n35141 );
not ( n35143 , n35140 );
not ( n35144 , RI17525ad8_649);
and ( n35145 , n35143 , n35144 );
nor ( n35146 , n35142 , n35145 );
xor ( n35147 , n35138 , n35146 );
buf ( n35148 , RI19aa9868_2499);
nand ( n35149 , n26059 , n35148 );
buf ( n35150 , RI17496258_1004);
and ( n35151 , n35149 , n35150 );
not ( n35152 , n35149 );
not ( n35153 , RI17496258_1004);
and ( n35154 , n35152 , n35153 );
nor ( n35155 , n35151 , n35154 );
xnor ( n35156 , n35147 , n35155 );
xor ( n35157 , n35125 , n35156 );
not ( n35158 , n35157 );
and ( n35159 , n35120 , n35158 );
not ( n35160 , n35120 );
and ( n35161 , n35160 , n35157 );
nor ( n35162 , n35159 , n35161 );
not ( n35163 , n35162 );
not ( n35164 , n35163 );
or ( n35165 , n35046 , n35164 );
nand ( n35166 , n35162 , n35044 );
nand ( n35167 , n35165 , n35166 );
xor ( n35168 , n28995 , n209033 );
not ( n35169 , n30321 );
xnor ( n35170 , n35168 , n35169 );
not ( n35171 , n35170 );
buf ( n35172 , RI19aa7540_2514);
nand ( n35173 , n29151 , n35172 );
buf ( n35174 , RI17523198_657);
and ( n35175 , n35173 , n35174 );
not ( n35176 , n35173 );
not ( n35177 , RI17523198_657);
and ( n35178 , n35176 , n35177 );
nor ( n35179 , n35175 , n35178 );
buf ( n35180 , n35179 );
not ( n35181 , n35180 );
not ( n35182 , n35181 );
not ( n35183 , n32443 );
or ( n35184 , n35182 , n35183 );
nand ( n35185 , n32442 , n35180 );
nand ( n35186 , n35184 , n35185 );
not ( n35187 , n35186 );
buf ( n35188 , n26222 );
not ( n35189 , n35188 );
and ( n35190 , n35187 , n35189 );
and ( n35191 , n35188 , n35186 );
nor ( n35192 , n35190 , n35191 );
not ( n35193 , n35192 );
nand ( n35194 , n35171 , n35193 );
buf ( n35195 , RI17455230_1321);
not ( n35196 , n35195 );
not ( n35197 , n205280 );
or ( n35198 , n35196 , n35197 );
not ( n35199 , n205280 );
not ( n35200 , n35199 );
or ( n35201 , n35200 , n35195 );
nand ( n35202 , n35198 , n35201 );
and ( n35203 , n35202 , n205322 );
not ( n35204 , n35202 );
and ( n35205 , n35204 , n205325 );
nor ( n35206 , n35203 , n35205 );
and ( n35207 , n35194 , n35206 );
not ( n35208 , n35194 );
not ( n35209 , n35206 );
and ( n35210 , n35208 , n35209 );
nor ( n35211 , n35207 , n35210 );
and ( n35212 , n35167 , n35211 );
not ( n35213 , n35167 );
not ( n35214 , n35211 );
and ( n35215 , n35213 , n35214 );
nor ( n35216 , n35212 , n35215 );
not ( n35217 , n35216 );
not ( n35218 , n35217 );
not ( n35219 , n35006 );
not ( n35220 , n35219 );
not ( n35221 , n25553 );
or ( n35222 , n35220 , n35221 );
not ( n35223 , n35219 );
not ( n35224 , n25553 );
nand ( n35225 , n35223 , n35224 );
nand ( n35226 , n35222 , n35225 );
and ( n35227 , n35226 , n34940 );
not ( n35228 , n35226 );
not ( n35229 , n29748 );
and ( n35230 , n35228 , n35229 );
nor ( n35231 , n35227 , n35230 );
not ( n35232 , n35231 );
buf ( n35233 , RI19acd5b0_2229);
nand ( n35234 , n30641 , n35233 );
not ( n35235 , RI17511600_712);
and ( n35236 , n35234 , n35235 );
not ( n35237 , n35234 );
buf ( n35238 , RI17511600_712);
and ( n35239 , n35237 , n35238 );
nor ( n35240 , n35236 , n35239 );
not ( n35241 , n35240 );
buf ( n35242 , RI17395ad0_2026);
not ( n35243 , n35242 );
not ( n35244 , RI173de7c0_1671);
not ( n35245 , n35244 );
or ( n35246 , n35243 , n35245 );
not ( n35247 , RI17395ad0_2026);
buf ( n35248 , RI173de7c0_1671);
nand ( n35249 , n35247 , n35248 );
nand ( n35250 , n35246 , n35249 );
buf ( n35251 , RI17456298_1316);
and ( n35252 , n35250 , n35251 );
not ( n35253 , n35250 );
not ( n35254 , RI17456298_1316);
and ( n35255 , n35253 , n35254 );
nor ( n35256 , n35252 , n35255 );
buf ( n35257 , RI19a946e8_2651);
nand ( n35258 , n25479 , n35257 );
buf ( n35259 , RI1747adf0_1137);
and ( n35260 , n35258 , n35259 );
not ( n35261 , n35258 );
not ( n35262 , RI1747adf0_1137);
and ( n35263 , n35261 , n35262 );
nor ( n35264 , n35260 , n35263 );
xor ( n35265 , n35256 , n35264 );
buf ( n35266 , RI19ac4910_2295);
nand ( n35267 , n205124 , n35266 );
not ( n35268 , RI174ca080_782);
and ( n35269 , n35267 , n35268 );
not ( n35270 , n35267 );
buf ( n35271 , RI174ca080_782);
and ( n35272 , n35270 , n35271 );
nor ( n35273 , n35269 , n35272 );
xor ( n35274 , n35265 , n35273 );
buf ( n35275 , n35274 );
not ( n35276 , n35275 );
or ( n213038 , n35241 , n35276 );
or ( n213039 , n35240 , n35275 );
nand ( n35279 , n213038 , n213039 );
buf ( n213041 , n34516 );
buf ( n213042 , n213041 );
and ( n35282 , n35279 , n213042 );
not ( n35283 , n35279 );
not ( n35284 , n213042 );
and ( n35285 , n35283 , n35284 );
nor ( n35286 , n35282 , n35285 );
not ( n35287 , n35286 );
nand ( n35288 , n35232 , n35287 );
not ( n35289 , n35288 );
buf ( n35290 , RI1744a790_1373);
not ( n35291 , n27961 );
xor ( n35292 , n35290 , n35291 );
xor ( n35293 , n35292 , n29372 );
not ( n35294 , n35293 );
not ( n35295 , n35294 );
or ( n35296 , n35289 , n35295 );
or ( n35297 , n35294 , n35288 );
nand ( n35298 , n35296 , n35297 );
not ( n35299 , n35298 );
not ( n35300 , n35299 );
xor ( n35301 , n205058 , n28247 );
xnor ( n35302 , n35301 , n32082 );
not ( n35303 , n35302 );
buf ( n35304 , RI1749cb58_972);
not ( n35305 , n35304 );
buf ( n35306 , RI19aba578_2378);
nand ( n35307 , n28637 , n35306 );
not ( n35308 , n35307 );
or ( n35309 , n35305 , n35308 );
or ( n35310 , n35307 , n35304 );
nand ( n35311 , n35309 , n35310 );
not ( n35312 , n35311 );
not ( n35313 , n26146 );
or ( n35314 , n35312 , n35313 );
or ( n35315 , n35311 , n26145 );
nand ( n35316 , n35314 , n35315 );
and ( n35317 , n35316 , n207796 );
not ( n35318 , n35316 );
and ( n35319 , n35318 , n30038 );
nor ( n35320 , n35317 , n35319 );
not ( n35321 , n35320 );
nand ( n35322 , n35303 , n35321 );
not ( n35323 , n35322 );
not ( n35324 , n33543 );
not ( n35325 , n29571 );
not ( n35326 , RI173a1290_1970);
not ( n35327 , n35326 );
or ( n35328 , n35325 , n35327 );
not ( n35329 , RI173e9f80_1615);
buf ( n35330 , RI173a1290_1970);
nand ( n35331 , n35329 , n35330 );
nand ( n35332 , n35328 , n35331 );
not ( n35333 , RI17467cc8_1230);
and ( n35334 , n35332 , n35333 );
not ( n35335 , n35332 );
buf ( n35336 , RI17467cc8_1230);
and ( n35337 , n35335 , n35336 );
nor ( n35338 , n35334 , n35337 );
buf ( n35339 , RI19aa10f0_2560);
nand ( n35340 , n28148 , n35339 );
buf ( n35341 , RI17486268_1082);
and ( n35342 , n35340 , n35341 );
not ( n35343 , n35340 );
not ( n35344 , RI17486268_1082);
and ( n35345 , n35343 , n35344 );
nor ( n35346 , n35342 , n35345 );
xor ( n35347 , n35338 , n35346 );
buf ( n35348 , RI19acffe0_2211);
nand ( n35349 , n25491 , n35348 );
buf ( n35350 , RI1750c8a8_727);
and ( n35351 , n35349 , n35350 );
not ( n35352 , n35349 );
not ( n35353 , RI1750c8a8_727);
and ( n35354 , n35352 , n35353 );
nor ( n35355 , n35351 , n35354 );
not ( n35356 , n35355 );
xnor ( n35357 , n35347 , n35356 );
buf ( n35358 , n35357 );
not ( n35359 , n35358 );
or ( n35360 , n35324 , n35359 );
or ( n35361 , n35358 , n33543 );
nand ( n35362 , n35360 , n35361 );
not ( n35363 , n35362 );
not ( n35364 , RI174458d0_1397);
buf ( n35365 , RI174074b8_1472);
not ( n35366 , n35365 );
not ( n35367 , RI173be7c8_1827);
not ( n35368 , n35367 );
or ( n35369 , n35366 , n35368 );
not ( n35370 , RI174074b8_1472);
buf ( n35371 , RI173be7c8_1827);
nand ( n35372 , n35370 , n35371 );
nand ( n35373 , n35369 , n35372 );
xor ( n35374 , n35364 , n35373 );
buf ( n35375 , RI19ab5118_2416);
nand ( n35376 , n28148 , n35375 );
buf ( n35377 , RI174a37a0_939);
and ( n35378 , n35376 , n35377 );
not ( n35379 , n35376 );
not ( n35380 , RI174a37a0_939);
and ( n35381 , n35379 , n35380 );
nor ( n35382 , n35378 , n35381 );
not ( n35383 , n35382 );
buf ( n35384 , RI17335248_2182);
not ( n35385 , n35384 );
and ( n35386 , n35383 , n35385 );
and ( n35387 , n35382 , n35384 );
nor ( n35388 , n35386 , n35387 );
xor ( n35389 , n35374 , n35388 );
not ( n35390 , n35389 );
not ( n35391 , n35390 );
and ( n35392 , n35363 , n35391 );
buf ( n35393 , n35390 );
and ( n35394 , n35362 , n35393 );
nor ( n35395 , n35392 , n35394 );
not ( n35396 , n35395 );
not ( n35397 , n35396 );
and ( n35398 , n35323 , n35397 );
and ( n35399 , n35322 , n35396 );
nor ( n35400 , n35398 , n35399 );
not ( n35401 , n35400 );
not ( n35402 , n35401 );
or ( n35403 , n35300 , n35402 );
nand ( n35404 , n35400 , n35298 );
nand ( n35405 , n35403 , n35404 );
not ( n35406 , n35405 );
and ( n35407 , n35218 , n35406 );
and ( n35408 , n35217 , n35405 );
nor ( n35409 , n35407 , n35408 );
buf ( n35410 , n35409 );
and ( n35411 , n34970 , n35410 );
not ( n35412 , n34970 );
and ( n35413 , n35216 , n35405 );
not ( n35414 , n35216 );
not ( n35415 , n35405 );
and ( n35416 , n35414 , n35415 );
nor ( n35417 , n35413 , n35416 );
buf ( n35418 , n35417 );
and ( n35419 , n35412 , n35418 );
nor ( n35420 , n35411 , n35419 );
not ( n35421 , n35420 );
nand ( n35422 , n34455 , n35421 );
or ( n35423 , n33256 , n35422 );
not ( n35424 , n35421 );
not ( n35425 , n33251 );
or ( n35426 , n35424 , n35425 );
buf ( n35427 , n27885 );
buf ( n35428 , n35427 );
nor ( n35429 , n34455 , n35428 );
nand ( n35430 , n35426 , n35429 );
buf ( n35431 , n31575 );
buf ( n35432 , RI1733f310_2133);
nand ( n35433 , n35431 , n35432 );
nand ( n35434 , n35423 , n35430 , n35433 );
buf ( n35435 , n35434 );
nor ( n35436 , n204263 , n25431 );
not ( n35437 , n35436 );
not ( n35438 , n31531 );
and ( n35439 , n35437 , n35438 );
and ( n35440 , n35436 , n31531 );
nor ( n35441 , n35439 , n35440 );
not ( n35442 , n35441 );
not ( n35443 , n35442 );
not ( n35444 , n31560 );
or ( n35445 , n35443 , n35444 );
not ( n35446 , n35442 );
nand ( n35447 , n35446 , n209312 );
nand ( n35448 , n35445 , n35447 );
not ( n35449 , n27968 );
buf ( n35450 , RI19a9e288_2583);
nand ( n35451 , n26325 , n35450 );
not ( n35452 , RI1748c4d8_1052);
and ( n35453 , n35451 , n35452 );
not ( n35454 , n35451 );
buf ( n35455 , RI1748c4d8_1052);
and ( n35456 , n35454 , n35455 );
nor ( n35457 , n35453 , n35456 );
not ( n35458 , n35457 );
not ( n35459 , n27961 );
or ( n35460 , n35458 , n35459 );
or ( n35461 , n35457 , n27960 );
nand ( n213223 , n35460 , n35461 );
not ( n213224 , n213223 );
and ( n35464 , n35449 , n213224 );
and ( n35465 , n27968 , n213223 );
nor ( n35466 , n35464 , n35465 );
not ( n35467 , n35466 );
not ( n35468 , n35467 );
buf ( n35469 , RI19a96998_2636);
nand ( n35470 , n25416 , n35469 );
buf ( n35471 , RI1752a830_634);
and ( n35472 , n35470 , n35471 );
not ( n35473 , n35470 );
not ( n35474 , RI1752a830_634);
and ( n35475 , n35473 , n35474 );
nor ( n35476 , n35472 , n35475 );
buf ( n35477 , n35476 );
not ( n35478 , n35477 );
not ( n35479 , n31126 );
or ( n35480 , n35478 , n35479 );
buf ( n35481 , n31125 );
not ( n35482 , n35481 );
or ( n35483 , n35482 , n35477 );
nand ( n35484 , n35480 , n35483 );
not ( n35485 , n35484 );
not ( n35486 , n31136 );
and ( n35487 , n35485 , n35486 );
and ( n35488 , n35484 , n31137 );
nor ( n35489 , n35487 , n35488 );
nand ( n35490 , n35489 , n27855 );
not ( n35491 , n35490 );
or ( n35492 , n35468 , n35491 );
or ( n35493 , n35467 , n35490 );
nand ( n35494 , n35492 , n35493 );
not ( n35495 , n35494 );
not ( n35496 , n31282 );
not ( n35497 , RI173ac3c0_1916);
not ( n35498 , n35497 );
or ( n35499 , n35496 , n35498 );
not ( n35500 , RI173f50b0_1561);
buf ( n35501 , RI173ac3c0_1916);
nand ( n35502 , n35500 , n35501 );
nand ( n35503 , n35499 , n35502 );
buf ( n35504 , RI17519c10_686);
and ( n35505 , n35503 , n35504 );
not ( n35506 , n35503 );
not ( n35507 , RI17519c10_686);
and ( n35508 , n35506 , n35507 );
nor ( n35509 , n35505 , n35508 );
buf ( n35510 , RI19aadd50_2469);
nand ( n35511 , n26453 , n35510 );
buf ( n35512 , RI174916e0_1027);
and ( n35513 , n35511 , n35512 );
not ( n35514 , n35511 );
not ( n35515 , RI174916e0_1027);
and ( n35516 , n35514 , n35515 );
nor ( n35517 , n35513 , n35516 );
xor ( n35518 , n35509 , n35517 );
buf ( n35519 , RI19ac1f58_2314);
nand ( n35520 , n205020 , n35519 );
not ( n35521 , RI1751e440_672);
and ( n35522 , n35520 , n35521 );
not ( n35523 , n35520 );
buf ( n35524 , RI1751e440_672);
and ( n35525 , n35523 , n35524 );
nor ( n35526 , n35522 , n35525 );
xnor ( n35527 , n35518 , n35526 );
xor ( n35528 , n30240 , n35527 );
xnor ( n35529 , n35528 , n28462 );
not ( n35530 , n35529 );
nand ( n35531 , n205392 , n35530 );
not ( n35532 , n35531 );
not ( n35533 , RI17406ae0_1475);
not ( n35534 , RI17405a78_1480);
buf ( n35535 , RI173bcd88_1835);
and ( n35536 , n35534 , n35535 );
not ( n35537 , n35534 );
not ( n35538 , RI173bcd88_1835);
and ( n35539 , n35537 , n35538 );
nor ( n35540 , n35536 , n35539 );
xor ( n35541 , n35533 , n35540 );
buf ( n35542 , RI17333808_2190);
buf ( n35543 , RI174a1d60_947);
xor ( n35544 , n35542 , n35543 );
buf ( n35545 , RI19ab65b8_2406);
nand ( n35546 , n25803 , n35545 );
xnor ( n35547 , n35544 , n35546 );
xnor ( n35548 , n35541 , n35547 );
not ( n35549 , n35548 );
buf ( n35550 , n29804 );
buf ( n35551 , RI173e8540_1623);
not ( n35552 , n35551 );
not ( n35553 , RI1739f508_1979);
not ( n35554 , n35553 );
or ( n35555 , n35552 , n35554 );
not ( n35556 , RI173e8540_1623);
buf ( n35557 , RI1739f508_1979);
nand ( n35558 , n35556 , n35557 );
nand ( n35559 , n35555 , n35558 );
not ( n35560 , RI17460018_1268);
and ( n35561 , n35559 , n35560 );
not ( n35562 , n35559 );
buf ( n35563 , RI17460018_1268);
and ( n35564 , n35562 , n35563 );
nor ( n35565 , n35561 , n35564 );
buf ( n35566 , RI19aa24a0_2550);
nand ( n35567 , n25364 , n35566 );
buf ( n35568 , RI17484828_1090);
and ( n35569 , n35567 , n35568 );
not ( n35570 , n35567 );
not ( n35571 , RI17484828_1090);
and ( n35572 , n35570 , n35571 );
nor ( n35573 , n35569 , n35572 );
xor ( n35574 , n35565 , n35573 );
buf ( n35575 , RI19a83690_2770);
nand ( n35576 , n26242 , n35575 );
buf ( n35577 , RI17509f68_735);
and ( n35578 , n35576 , n35577 );
not ( n35579 , n35576 );
not ( n35580 , RI17509f68_735);
and ( n35581 , n35579 , n35580 );
nor ( n35582 , n35578 , n35581 );
not ( n35583 , n35582 );
xnor ( n35584 , n35574 , n35583 );
and ( n35585 , n35550 , n35584 );
not ( n35586 , n35550 );
not ( n35587 , n35565 );
xor ( n35588 , n35587 , n35582 );
not ( n35589 , n35573 );
xnor ( n35590 , n35588 , n35589 );
and ( n35591 , n35586 , n35590 );
nor ( n35592 , n35585 , n35591 );
not ( n35593 , n35592 );
not ( n35594 , n35593 );
or ( n35595 , n35549 , n35594 );
not ( n35596 , n35548 );
nand ( n35597 , n35592 , n35596 );
nand ( n35598 , n35595 , n35597 );
not ( n35599 , n35598 );
not ( n35600 , n35599 );
not ( n213362 , n35600 );
and ( n213363 , n35532 , n213362 );
not ( n35603 , n35529 );
nand ( n35604 , n35603 , n205392 );
and ( n35605 , n35604 , n35600 );
nor ( n35606 , n213363 , n35605 );
not ( n35607 , n35606 );
or ( n35608 , n35495 , n35607 );
or ( n35609 , n35606 , n35494 );
nand ( n35610 , n35608 , n35609 );
buf ( n35611 , n25924 );
not ( n35612 , n35611 );
not ( n35613 , n31967 );
or ( n35614 , n35612 , n35613 );
not ( n35615 , n35611 );
nand ( n35616 , n35615 , n209733 );
nand ( n35617 , n35614 , n35616 );
and ( n35618 , n35617 , n32011 );
not ( n35619 , n35617 );
xor ( n35620 , n31988 , n32005 );
not ( n35621 , n31996 );
xnor ( n35622 , n35620 , n35621 );
not ( n35623 , n35622 );
not ( n35624 , n35623 );
and ( n35625 , n35619 , n35624 );
nor ( n35626 , n35618 , n35625 );
not ( n35627 , RI175373a0_595);
not ( n35628 , n35627 );
not ( n35629 , RI1753a460_587);
not ( n35630 , RI17536770_597);
nand ( n35631 , n35629 , n35630 );
nand ( n35632 , n204517 , n204523 );
nor ( n35633 , n35628 , n35631 , n35632 );
xor ( n35634 , n35626 , n35633 );
not ( n35635 , n25597 );
not ( n35636 , n35635 );
not ( n35637 , n25549 );
not ( n35638 , n35016 );
not ( n35639 , n35638 );
and ( n35640 , n35637 , n35639 );
and ( n35641 , n25549 , n35638 );
nor ( n35642 , n35640 , n35641 );
not ( n35643 , n35642 );
or ( n213405 , n35636 , n35643 );
or ( n213406 , n35642 , n25598 );
nand ( n35646 , n213405 , n213406 );
buf ( n35647 , n35646 );
not ( n35648 , n35647 );
nand ( n35649 , n35648 , n205224 );
and ( n35650 , n35634 , n35649 );
not ( n35651 , n35634 );
not ( n35652 , n35649 );
and ( n35653 , n35651 , n35652 );
nor ( n35654 , n35650 , n35653 );
and ( n35655 , n35610 , n35654 );
not ( n35656 , n35610 );
not ( n35657 , n35654 );
and ( n35658 , n35656 , n35657 );
nor ( n35659 , n35655 , n35658 );
buf ( n35660 , RI19abe808_2345);
nand ( n35661 , n27749 , n35660 );
buf ( n35662 , RI174b2098_868);
and ( n35663 , n35661 , n35662 );
not ( n35664 , n35661 );
not ( n35665 , RI174b2098_868);
and ( n35666 , n35664 , n35665 );
nor ( n35667 , n35663 , n35666 );
not ( n35668 , n35667 );
not ( n35669 , n35668 );
not ( n35670 , n35390 );
or ( n35671 , n35669 , n35670 );
not ( n35672 , n35668 );
nand ( n35673 , n35672 , n35389 );
nand ( n35674 , n35671 , n35673 );
buf ( n35675 , RI173dbd18_1684);
not ( n35676 , n35675 );
not ( n35677 , RI17393028_2039);
not ( n35678 , n35677 );
or ( n35679 , n35676 , n35678 );
not ( n35680 , RI173dbd18_1684);
buf ( n35681 , RI17393028_2039);
nand ( n35682 , n35680 , n35681 );
nand ( n35683 , n35679 , n35682 );
buf ( n35684 , RI174537f0_1329);
and ( n35685 , n35683 , n35684 );
not ( n35686 , n35683 );
not ( n35687 , RI174537f0_1329);
and ( n35688 , n35686 , n35687 );
nor ( n35689 , n35685 , n35688 );
buf ( n35690 , RI19a97b68_2628);
nand ( n35691 , n26276 , n35690 );
buf ( n35692 , RI17478348_1150);
xor ( n35693 , n35691 , n35692 );
xor ( n35694 , n35689 , n35693 );
buf ( n35695 , RI19ac7958_2273);
nand ( n35696 , n28637 , n35695 );
not ( n35697 , RI174c5d78_795);
and ( n35698 , n35696 , n35697 );
not ( n35699 , n35696 );
buf ( n35700 , RI174c5d78_795);
and ( n35701 , n35699 , n35700 );
nor ( n35702 , n35698 , n35701 );
xor ( n35703 , n35694 , n35702 );
buf ( n35704 , n35703 );
buf ( n35705 , n35704 );
xnor ( n35706 , n35674 , n35705 );
not ( n35707 , n35706 );
nand ( n35708 , n35707 , n204983 );
not ( n35709 , n35708 );
buf ( n35710 , RI19ab6090_2408);
nand ( n35711 , n205271 , n35710 );
not ( n35712 , n35711 );
buf ( n35713 , RI174a16d0_949);
not ( n35714 , n35713 );
and ( n35715 , n35712 , n35714 );
and ( n35716 , n35711 , n35713 );
nor ( n35717 , n35715 , n35716 );
not ( n35718 , n35717 );
not ( n35719 , n35718 );
not ( n35720 , n207706 );
or ( n35721 , n35719 , n35720 );
not ( n35722 , n29944 );
nand ( n35723 , n35722 , n35717 );
nand ( n35724 , n35721 , n35723 );
not ( n35725 , n35724 );
not ( n35726 , n211419 );
and ( n35727 , n35725 , n35726 );
and ( n35728 , n35724 , n211419 );
nor ( n35729 , n35727 , n35728 );
not ( n35730 , n35729 );
not ( n35731 , n35730 );
and ( n35732 , n35709 , n35731 );
and ( n35733 , n35708 , n35730 );
nor ( n35734 , n35732 , n35733 );
not ( n35735 , n35734 );
not ( n35736 , n35735 );
not ( n35737 , n32005 );
xor ( n35738 , n29233 , n29250 );
not ( n35739 , n207002 );
xnor ( n35740 , n35738 , n35739 );
not ( n35741 , n35740 );
or ( n35742 , n35737 , n35741 );
or ( n35743 , n35740 , n32005 );
nand ( n35744 , n35742 , n35743 );
and ( n35745 , n35744 , n29258 );
not ( n35746 , n35744 );
and ( n35747 , n35746 , n29214 );
nor ( n35748 , n35745 , n35747 );
not ( n35749 , n35748 );
not ( n35750 , n35749 );
buf ( n35751 , n32756 );
xor ( n35752 , n30990 , n30998 );
xnor ( n35753 , n35752 , n31007 );
buf ( n35754 , n35753 );
xor ( n35755 , n35751 , n35754 );
buf ( n35756 , RI1744c860_1363);
buf ( n35757 , RI19acbe40_2240);
nand ( n35758 , n25879 , n35757 );
buf ( n35759 , RI174ba900_830);
and ( n35760 , n35758 , n35759 );
not ( n35761 , n35758 );
not ( n35762 , RI174ba900_830);
and ( n35763 , n35761 , n35762 );
nor ( n35764 , n35760 , n35763 );
xor ( n35765 , n35756 , n35764 );
buf ( n35766 , RI19a9ce60_2591);
nand ( n35767 , n25711 , n35766 );
not ( n35768 , RI17471070_1185);
and ( n35769 , n35767 , n35768 );
not ( n35770 , n35767 );
buf ( n35771 , RI17471070_1185);
and ( n35772 , n35770 , n35771 );
nor ( n35773 , n35769 , n35772 );
xnor ( n35774 , n35765 , n35773 );
not ( n35775 , n35774 );
not ( n35776 , RI173d4d88_1718);
buf ( n35777 , RI1738c098_2073);
and ( n35778 , n35776 , n35777 );
not ( n35779 , n35776 );
not ( n35780 , RI1738c098_2073);
and ( n35781 , n35779 , n35780 );
nor ( n35782 , n35778 , n35781 );
not ( n35783 , n35782 );
and ( n35784 , n35775 , n35783 );
and ( n35785 , n35774 , n35782 );
nor ( n35786 , n35784 , n35785 );
not ( n35787 , n35786 );
xnor ( n35788 , n35755 , n35787 );
not ( n35789 , n35788 );
nand ( n35790 , n35789 , n204750 );
not ( n35791 , n35790 );
or ( n35792 , n35750 , n35791 );
or ( n35793 , n35790 , n35749 );
nand ( n35794 , n35792 , n35793 );
not ( n35795 , n35794 );
not ( n35796 , n35795 );
or ( n35797 , n35736 , n35796 );
nand ( n35798 , n35794 , n35734 );
nand ( n35799 , n35797 , n35798 );
and ( n35800 , n35659 , n35799 );
not ( n35801 , n35659 );
not ( n35802 , n35799 );
and ( n35803 , n35801 , n35802 );
nor ( n35804 , n35800 , n35803 );
buf ( n35805 , n35804 );
and ( n35806 , n35448 , n35805 );
not ( n35807 , n35448 );
and ( n35808 , n35659 , n35802 );
not ( n35809 , n35659 );
and ( n35810 , n35809 , n35799 );
nor ( n35811 , n35808 , n35810 );
not ( n35812 , n35811 );
not ( n35813 , n35812 );
and ( n35814 , n35807 , n35813 );
nor ( n35815 , n35806 , n35814 );
not ( n35816 , n205649 );
nor ( n35817 , n35815 , n35816 );
not ( n35818 , n31326 );
xor ( n35819 , n31594 , n31611 );
not ( n35820 , n209363 );
xnor ( n35821 , n35819 , n35820 );
not ( n35822 , n35821 );
or ( n35823 , n35818 , n35822 );
or ( n35824 , n35821 , n31326 );
nand ( n35825 , n35823 , n35824 );
not ( n35826 , n33257 );
not ( n35827 , RI173c9c40_1772);
not ( n35828 , n35827 );
or ( n35829 , n35826 , n35828 );
not ( n35830 , RI173406c0_2127);
buf ( n35831 , RI173c9c40_1772);
nand ( n35832 , n35830 , n35831 );
nand ( n35833 , n35829 , n35832 );
not ( n35834 , RI17412c78_1416);
and ( n35835 , n35833 , n35834 );
not ( n35836 , n35833 );
buf ( n35837 , RI17412c78_1416);
and ( n35838 , n35836 , n35837 );
nor ( n35839 , n35835 , n35838 );
buf ( n35840 , RI19ac0ba8_2325);
nand ( n35841 , n29151 , n35840 );
buf ( n35842 , RI174aef60_883);
and ( n35843 , n35841 , n35842 );
not ( n35844 , n35841 );
not ( n35845 , RI174aef60_883);
and ( n213607 , n35844 , n35845 );
nor ( n213608 , n35843 , n213607 );
xor ( n35848 , n35839 , n213608 );
buf ( n35849 , RI19a905c0_2680);
nand ( n35850 , n26059 , n35849 );
buf ( n35851 , RI17466288_1238);
and ( n35852 , n35850 , n35851 );
not ( n35853 , n35850 );
not ( n35854 , RI17466288_1238);
and ( n35855 , n35853 , n35854 );
nor ( n35856 , n35852 , n35855 );
xnor ( n35857 , n35848 , n35856 );
buf ( n35858 , n35857 );
and ( n213620 , n35825 , n35858 );
not ( n213621 , n35825 );
not ( n35861 , n35858 );
and ( n35862 , n213621 , n35861 );
nor ( n35863 , n213620 , n35862 );
not ( n35864 , n35863 );
not ( n35865 , n30032 );
buf ( n35866 , RI173d4a40_1719);
not ( n35867 , n30974 );
not ( n35868 , RI173b7ec8_1859);
not ( n35869 , n35868 );
or ( n35870 , n35867 , n35869 );
not ( n35871 , RI17400bb8_1504);
buf ( n35872 , RI173b7ec8_1859);
nand ( n35873 , n35871 , n35872 );
nand ( n35874 , n35870 , n35873 );
xor ( n35875 , n35866 , n35874 );
buf ( n35876 , RI17530500_616);
buf ( n35877 , RI1749cea0_971);
xor ( n35878 , n35876 , n35877 );
buf ( n35879 , RI19aba8c0_2377);
nand ( n35880 , n28902 , n35879 );
xnor ( n35881 , n35878 , n35880 );
xnor ( n35882 , n35875 , n35881 );
not ( n35883 , n35882 );
or ( n35884 , n35865 , n35883 );
not ( n35885 , n30032 );
not ( n35886 , n35874 );
xor ( n35887 , n35866 , n35886 );
xnor ( n35888 , n35887 , n35881 );
nand ( n35889 , n35885 , n35888 );
nand ( n35890 , n35884 , n35889 );
buf ( n35891 , RI173d5418_1716);
not ( n35892 , n35891 );
not ( n35893 , n30813 );
or ( n35894 , n35892 , n35893 );
not ( n35895 , RI173d5418_1716);
buf ( n35896 , RI1738c728_2071);
nand ( n35897 , n35895 , n35896 );
nand ( n35898 , n35894 , n35897 );
buf ( n35899 , RI1744cef0_1361);
and ( n35900 , n35898 , n35899 );
not ( n35901 , n35898 );
not ( n35902 , RI1744cef0_1361);
and ( n35903 , n35901 , n35902 );
nor ( n35904 , n35900 , n35903 );
buf ( n35905 , RI19a9aac0_2607);
nand ( n35906 , n25582 , n35905 );
buf ( n35907 , RI17471700_1183);
and ( n35908 , n35906 , n35907 );
not ( n35909 , n35906 );
not ( n35910 , RI17471700_1183);
and ( n35911 , n35909 , n35910 );
nor ( n35912 , n35908 , n35911 );
xor ( n35913 , n35904 , n35912 );
buf ( n35914 , RI19aca298_2254);
nand ( n35915 , n204916 , n35914 );
not ( n35916 , RI174bb350_828);
and ( n35917 , n35915 , n35916 );
not ( n35918 , n35915 );
buf ( n35919 , RI174bb350_828);
and ( n35920 , n35918 , n35919 );
nor ( n35921 , n35917 , n35920 );
xnor ( n35922 , n35913 , n35921 );
not ( n35923 , n35922 );
and ( n35924 , n35890 , n35923 );
not ( n35925 , n35890 );
buf ( n35926 , n35922 );
and ( n35927 , n35925 , n35926 );
nor ( n35928 , n35924 , n35927 );
not ( n35929 , n35928 );
nand ( n35930 , n35864 , n35929 );
not ( n35931 , n35548 );
not ( n35932 , n29782 );
not ( n35933 , n35584 );
or ( n35934 , n35932 , n35933 );
not ( n35935 , n29782 );
nand ( n35936 , n35935 , n35590 );
nand ( n35937 , n35934 , n35936 );
not ( n35938 , n35937 );
or ( n35939 , n35931 , n35938 );
not ( n35940 , n35596 );
or ( n35941 , n35940 , n35937 );
nand ( n35942 , n35939 , n35941 );
buf ( n35943 , n35942 );
xnor ( n35944 , n35930 , n35943 );
buf ( n35945 , n35944 );
not ( n35946 , n35945 );
buf ( n35947 , RI173df198_1668);
not ( n35948 , n35947 );
not ( n35949 , n33134 );
or ( n35950 , n35948 , n35949 );
not ( n35951 , n35947 );
nand ( n35952 , n35951 , n33140 );
nand ( n35953 , n35950 , n35952 );
and ( n35954 , n35953 , n34603 );
not ( n35955 , n35953 );
and ( n35956 , n35955 , n30689 );
nor ( n35957 , n35954 , n35956 );
not ( n35958 , n31884 );
xor ( n35959 , n205369 , n205373 );
xnor ( n35960 , n35959 , n205382 );
not ( n35961 , n35960 );
or ( n35962 , n35958 , n35961 );
or ( n35963 , n35960 , n31884 );
nand ( n35964 , n35962 , n35963 );
and ( n35965 , n35964 , n30756 );
not ( n35966 , n35964 );
and ( n35967 , n35966 , n30771 );
nor ( n35968 , n35965 , n35967 );
not ( n35969 , n35968 );
nand ( n35970 , n35957 , n35969 );
not ( n35971 , n204907 );
not ( n35972 , n33986 );
or ( n35973 , n35971 , n35972 );
or ( n35974 , n33986 , n204907 );
nand ( n35975 , n35973 , n35974 );
buf ( n35976 , RI19a9b1c8_2604);
nand ( n35977 , n25915 , n35976 );
buf ( n35978 , RI174720d8_1180);
and ( n35979 , n35977 , n35978 );
not ( n35980 , n35977 );
not ( n35981 , RI174720d8_1180);
and ( n35982 , n35980 , n35981 );
nor ( n35983 , n35979 , n35982 );
not ( n35984 , n35983 );
buf ( n35985 , RI19aca9a0_2251);
nand ( n35986 , n204572 , n35985 );
not ( n35987 , RI174bc2c8_825);
and ( n35988 , n35986 , n35987 );
not ( n35989 , n35986 );
buf ( n35990 , RI174bc2c8_825);
and ( n35991 , n35989 , n35990 );
nor ( n35992 , n35988 , n35991 );
not ( n35993 , n35992 );
or ( n35994 , n35984 , n35993 );
or ( n35995 , n35983 , n35992 );
nand ( n35996 , n35994 , n35995 );
buf ( n35997 , RI173d5df0_1713);
not ( n35998 , n35997 );
not ( n35999 , RI1738d100_2068);
not ( n36000 , n35999 );
or ( n36001 , n35998 , n36000 );
not ( n36002 , RI173d5df0_1713);
buf ( n36003 , RI1738d100_2068);
nand ( n36004 , n36002 , n36003 );
nand ( n36005 , n36001 , n36004 );
buf ( n36006 , RI1744d8c8_1358);
and ( n213768 , n36005 , n36006 );
not ( n213769 , n36005 );
not ( n36009 , RI1744d8c8_1358);
and ( n36010 , n213769 , n36009 );
nor ( n36011 , n213768 , n36010 );
not ( n213773 , n36011 );
and ( n213774 , n35996 , n213773 );
not ( n36014 , n35996 );
and ( n213776 , n36014 , n36011 );
nor ( n213777 , n213774 , n213776 );
not ( n36017 , n213777 );
not ( n36018 , n36017 );
and ( n36019 , n35975 , n36018 );
not ( n36020 , n35975 );
buf ( n36021 , n35983 );
xor ( n36022 , n36011 , n36021 );
buf ( n36023 , n35992 );
xnor ( n36024 , n36022 , n36023 );
buf ( n36025 , n36024 );
and ( n36026 , n36020 , n36025 );
nor ( n36027 , n36019 , n36026 );
not ( n36028 , n36027 );
xnor ( n36029 , n35970 , n36028 );
not ( n36030 , n36029 );
not ( n36031 , n36030 );
not ( n36032 , n35942 );
nand ( n36033 , n36032 , n35863 );
not ( n36034 , n36033 );
not ( n36035 , RI173a4710_1954);
not ( n36036 , n36035 );
not ( n36037 , n36036 );
buf ( n36038 , RI173deb08_1670);
not ( n36039 , n36038 );
not ( n36040 , RI17395e18_2025);
not ( n36041 , n36040 );
or ( n36042 , n36039 , n36041 );
not ( n36043 , RI173deb08_1670);
buf ( n36044 , RI17395e18_2025);
nand ( n36045 , n36043 , n36044 );
nand ( n36046 , n36042 , n36045 );
not ( n36047 , RI174565e0_1315);
and ( n36048 , n36046 , n36047 );
not ( n36049 , n36046 );
buf ( n36050 , RI174565e0_1315);
and ( n36051 , n36049 , n36050 );
nor ( n36052 , n36048 , n36051 );
buf ( n36053 , RI19ac4b68_2294);
nand ( n36054 , n25416 , n36053 );
buf ( n36055 , RI174ca5a8_781);
and ( n36056 , n36054 , n36055 );
not ( n36057 , n36054 );
not ( n36058 , RI174ca5a8_781);
and ( n36059 , n36057 , n36058 );
nor ( n36060 , n36056 , n36059 );
xor ( n36061 , n36052 , n36060 );
buf ( n36062 , RI19a94940_2650);
nand ( n36063 , n25416 , n36062 );
buf ( n36064 , RI1747b138_1136);
and ( n36065 , n36063 , n36064 );
not ( n36066 , n36063 );
not ( n36067 , RI1747b138_1136);
and ( n36068 , n36066 , n36067 );
nor ( n36069 , n36065 , n36068 );
xnor ( n36070 , n36061 , n36069 );
not ( n36071 , n36070 );
not ( n36072 , n36071 );
or ( n36073 , n36037 , n36072 );
not ( n36074 , n36070 );
or ( n36075 , n36074 , n36036 );
nand ( n36076 , n36073 , n36075 );
and ( n36077 , n36076 , n33096 );
not ( n36078 , n36076 );
and ( n36079 , n36078 , n33099 );
nor ( n36080 , n36077 , n36079 );
not ( n36081 , n36080 );
not ( n36082 , n36081 );
and ( n36083 , n36034 , n36082 );
and ( n36084 , n36033 , n36081 );
nor ( n36085 , n36083 , n36084 );
not ( n36086 , n36085 );
not ( n36087 , n36086 );
or ( n36088 , n36031 , n36087 );
nand ( n36089 , n36085 , n36029 );
nand ( n36090 , n36088 , n36089 );
buf ( n36091 , RI173cfb68_1743);
xor ( n36092 , n36091 , n35275 );
buf ( n36093 , n28146 );
xnor ( n36094 , n36092 , n36093 );
buf ( n36095 , RI1744d238_1360);
not ( n36096 , n36095 );
not ( n36097 , n26261 );
or ( n36098 , n36096 , n36097 );
or ( n36099 , n26261 , n36095 );
nand ( n36100 , n36098 , n36099 );
and ( n36101 , n36100 , n26319 );
not ( n36102 , n36100 );
and ( n36103 , n36102 , n26311 );
nor ( n36104 , n36101 , n36103 );
nand ( n36105 , n36094 , n36104 );
not ( n213867 , n36105 );
not ( n213868 , n29759 );
not ( n36108 , n28779 );
or ( n36109 , n213868 , n36108 );
or ( n36110 , n28779 , n29759 );
nand ( n36111 , n36109 , n36110 );
and ( n36112 , n36111 , n206591 );
not ( n36113 , n36111 );
and ( n36114 , n36113 , n28817 );
nor ( n36115 , n36112 , n36114 );
not ( n36116 , n36115 );
not ( n36117 , n36116 );
and ( n36118 , n213867 , n36117 );
and ( n36119 , n36105 , n36116 );
nor ( n36120 , n36118 , n36119 );
and ( n36121 , n36090 , n36120 );
not ( n36122 , n36090 );
not ( n36123 , n36120 );
and ( n36124 , n36122 , n36123 );
nor ( n36125 , n36121 , n36124 );
not ( n36126 , n36125 );
not ( n36127 , n33016 );
buf ( n36128 , RI17461080_1263);
buf ( n36129 , RI173a08b8_1973);
not ( n36130 , n36129 );
not ( n36131 , RI173e95a8_1618);
not ( n36132 , n36131 );
or ( n36133 , n36130 , n36132 );
not ( n36134 , RI173a08b8_1973);
buf ( n36135 , RI173e95a8_1618);
nand ( n36136 , n36134 , n36135 );
nand ( n36137 , n36133 , n36136 );
buf ( n36138 , n36137 );
xor ( n36139 , n36128 , n36138 );
buf ( n36140 , RI19acf8d8_2214);
nand ( n36141 , n27946 , n36140 );
not ( n36142 , RI1750b930_730);
and ( n36143 , n36141 , n36142 );
not ( n36144 , n36141 );
buf ( n36145 , RI1750b930_730);
and ( n36146 , n36144 , n36145 );
nor ( n36147 , n36143 , n36146 );
not ( n36148 , n36147 );
not ( n36149 , n36148 );
buf ( n36150 , RI19aa0b50_2563);
nand ( n36151 , n27946 , n36150 );
buf ( n36152 , RI17485890_1085);
and ( n36153 , n36151 , n36152 );
not ( n36154 , n36151 );
not ( n36155 , RI17485890_1085);
and ( n36156 , n36154 , n36155 );
nor ( n36157 , n36153 , n36156 );
not ( n36158 , n36157 );
not ( n36159 , n36158 );
or ( n36160 , n36149 , n36159 );
nand ( n36161 , n36157 , n36147 );
nand ( n36162 , n36160 , n36161 );
xnor ( n213924 , n36139 , n36162 );
not ( n213925 , n213924 );
or ( n36165 , n36127 , n213925 );
not ( n213927 , RI17461080_1263);
xor ( n213928 , n213927 , n36137 );
xor ( n36168 , n213928 , n36162 );
or ( n36169 , n36168 , n33016 );
nand ( n36170 , n36165 , n36169 );
buf ( n36171 , RI173bdaa8_1831);
not ( n36172 , n36171 );
not ( n36173 , RI17406798_1476);
not ( n213935 , n36173 );
or ( n213936 , n36172 , n213935 );
not ( n36176 , RI173bdaa8_1831);
buf ( n36177 , RI17406798_1476);
nand ( n36178 , n36176 , n36177 );
nand ( n36179 , n213936 , n36178 );
xor ( n36180 , n28559 , n36179 );
buf ( n36181 , RI17334528_2186);
buf ( n36182 , RI174a2a80_943);
xor ( n36183 , n36181 , n36182 );
buf ( n36184 , RI19ab48a8_2419);
nand ( n36185 , n28637 , n36184 );
xnor ( n36186 , n36183 , n36185 );
xnor ( n36187 , n36180 , n36186 );
not ( n36188 , n36187 );
not ( n36189 , n36188 );
not ( n36190 , n36189 );
and ( n36191 , n36170 , n36190 );
not ( n36192 , n36170 );
and ( n36193 , n36192 , n36189 );
nor ( n36194 , n36191 , n36193 );
not ( n36195 , n36194 );
xor ( n36196 , n32938 , n29910 );
xnor ( n36197 , n36196 , n26009 );
not ( n36198 , n36197 );
buf ( n36199 , RI17402940_1495);
not ( n36200 , n36199 );
not ( n36201 , n31177 );
or ( n36202 , n36200 , n36201 );
or ( n36203 , n31177 , n36199 );
nand ( n36204 , n36202 , n36203 );
buf ( n36205 , RI173c8548_1779);
not ( n36206 , n36205 );
not ( n36207 , RI1733efc8_2134);
not ( n36208 , n36207 );
or ( n36209 , n36206 , n36208 );
not ( n36210 , RI173c8548_1779);
buf ( n36211 , RI1733efc8_2134);
nand ( n36212 , n36210 , n36211 );
nand ( n36213 , n36209 , n36212 );
and ( n36214 , n36213 , n29969 );
not ( n36215 , n36213 );
not ( n36216 , RI17411238_1424);
and ( n36217 , n36215 , n36216 );
nor ( n36218 , n36214 , n36217 );
buf ( n36219 , RI19a8f648_2687);
nand ( n36220 , n25622 , n36219 );
buf ( n36221 , RI17464b90_1245);
and ( n36222 , n36220 , n36221 );
not ( n36223 , n36220 );
not ( n36224 , RI17464b90_1245);
and ( n36225 , n36223 , n36224 );
nor ( n36226 , n36222 , n36225 );
not ( n36227 , n36226 );
xor ( n36228 , n36218 , n36227 );
buf ( n36229 , RI19abff78_2332);
nand ( n36230 , n204513 , n36229 );
not ( n36231 , RI174ad868_890);
and ( n36232 , n36230 , n36231 );
not ( n36233 , n36230 );
buf ( n36234 , RI174ad868_890);
and ( n36235 , n36233 , n36234 );
nor ( n36236 , n36232 , n36235 );
xnor ( n36237 , n36228 , n36236 );
buf ( n36238 , n36237 );
and ( n36239 , n36204 , n36238 );
not ( n36240 , n36204 );
xor ( n36241 , n36218 , n36226 );
xnor ( n36242 , n36241 , n36236 );
buf ( n36243 , n36242 );
and ( n36244 , n36240 , n36243 );
nor ( n36245 , n36239 , n36244 );
nand ( n36246 , n36198 , n36245 );
not ( n36247 , n36246 );
or ( n36248 , n36195 , n36247 );
not ( n36249 , n36245 );
not ( n36250 , n36249 );
nand ( n36251 , n36250 , n36198 );
or ( n36252 , n36251 , n36194 );
nand ( n36253 , n36248 , n36252 );
not ( n36254 , n36253 );
buf ( n36255 , n209733 );
xor ( n214017 , n205663 , n36255 );
xor ( n214018 , n33802 , n33777 );
xnor ( n36258 , n214018 , n33801 );
xnor ( n36259 , n214017 , n36258 );
xor ( n36260 , n32808 , n32825 );
buf ( n36261 , n32816 );
xnor ( n36262 , n36260 , n36261 );
not ( n36263 , n36262 );
not ( n36264 , n36263 );
xor ( n36265 , n28470 , n36264 );
xnor ( n36266 , n36265 , n32863 );
nand ( n36267 , n36259 , n36266 );
not ( n36268 , n36267 );
not ( n36269 , n28313 );
buf ( n36270 , RI19a8f8a0_2686);
nand ( n36271 , n25364 , n36270 );
buf ( n36272 , RI17464ed8_1244);
and ( n36273 , n36271 , n36272 );
not ( n36274 , n36271 );
not ( n36275 , RI17464ed8_1244);
and ( n36276 , n36274 , n36275 );
nor ( n36277 , n36273 , n36276 );
not ( n36278 , n36277 );
buf ( n36279 , RI19ac0158_2331);
nand ( n36280 , n25451 , n36279 );
not ( n36281 , RI174adbb0_889);
and ( n36282 , n36280 , n36281 );
not ( n36283 , n36280 );
buf ( n36284 , RI174adbb0_889);
and ( n36285 , n36283 , n36284 );
nor ( n36286 , n36282 , n36285 );
not ( n36287 , n36286 );
or ( n36288 , n36278 , n36287 );
or ( n36289 , n36277 , n36286 );
nand ( n36290 , n36288 , n36289 );
buf ( n36291 , RI173c8890_1778);
not ( n36292 , n36291 );
not ( n36293 , RI1733f310_2133);
not ( n36294 , n36293 );
or ( n36295 , n36292 , n36294 );
not ( n36296 , RI173c8890_1778);
nand ( n214058 , n36296 , n35432 );
nand ( n214059 , n36295 , n214058 );
not ( n36299 , RI17411580_1423);
and ( n36300 , n214059 , n36299 );
not ( n36301 , n214059 );
and ( n36302 , n36301 , n31039 );
nor ( n36303 , n36300 , n36302 );
not ( n36304 , n36303 );
and ( n36305 , n36290 , n36304 );
not ( n36306 , n36290 );
and ( n36307 , n36306 , n36303 );
nor ( n36308 , n36305 , n36307 );
not ( n36309 , n36308 );
not ( n36310 , n36309 );
or ( n36311 , n36269 , n36310 );
not ( n36312 , n36309 );
nand ( n36313 , n36312 , n28309 );
nand ( n36314 , n36311 , n36313 );
buf ( n36315 , RI173e6128_1634);
not ( n36316 , n36315 );
not ( n36317 , RI1739d0f0_1990);
not ( n36318 , n36317 );
or ( n36319 , n36316 , n36318 );
not ( n36320 , RI173e6128_1634);
buf ( n36321 , RI1739d0f0_1990);
nand ( n36322 , n36320 , n36321 );
nand ( n36323 , n36319 , n36322 );
buf ( n36324 , RI1745dc00_1279);
and ( n36325 , n36323 , n36324 );
not ( n36326 , n36323 );
not ( n36327 , RI1745dc00_1279);
and ( n36328 , n36326 , n36327 );
nor ( n36329 , n36325 , n36328 );
buf ( n36330 , RI19aa3418_2543);
nand ( n36331 , n26242 , n36330 );
not ( n36332 , RI17482410_1101);
and ( n36333 , n36331 , n36332 );
not ( n36334 , n36331 );
buf ( n36335 , RI17482410_1101);
and ( n36336 , n36334 , n36335 );
nor ( n36337 , n36333 , n36336 );
xor ( n36338 , n36329 , n36337 );
buf ( n36339 , RI19a846f8_2763);
nand ( n36340 , n25880 , n36339 );
not ( n36341 , RI175066b0_746);
and ( n36342 , n36340 , n36341 );
not ( n36343 , n36340 );
buf ( n36344 , RI175066b0_746);
and ( n36345 , n36343 , n36344 );
nor ( n36346 , n36342 , n36345 );
xnor ( n36347 , n36338 , n36346 );
not ( n36348 , n36347 );
buf ( n36349 , n36348 );
not ( n36350 , n36349 );
and ( n36351 , n36314 , n36350 );
not ( n36352 , n36314 );
and ( n36353 , n36352 , n36349 );
nor ( n36354 , n36351 , n36353 );
not ( n36355 , n36354 );
not ( n36356 , n36355 );
and ( n36357 , n36268 , n36356 );
and ( n36358 , n36267 , n36355 );
nor ( n36359 , n36357 , n36358 );
not ( n36360 , n36359 );
or ( n36361 , n36254 , n36360 );
or ( n36362 , n36253 , n36359 );
nand ( n36363 , n36361 , n36362 );
not ( n36364 , n36363 );
or ( n36365 , n36126 , n36364 );
or ( n36366 , n36363 , n36125 );
nand ( n36367 , n36365 , n36366 );
not ( n36368 , n36367 );
not ( n36369 , n36368 );
or ( n36370 , n35946 , n36369 );
not ( n36371 , n35945 );
buf ( n36372 , n36367 );
nand ( n36373 , n36371 , n36372 );
nand ( n36374 , n36370 , n36373 );
not ( n36375 , n36374 );
xor ( n36376 , n32765 , n35754 );
buf ( n36377 , n35786 );
xnor ( n36378 , n36376 , n36377 );
not ( n36379 , n36378 );
buf ( n36380 , n31967 );
xor ( n36381 , n27920 , n36380 );
xnor ( n36382 , n36381 , n36258 );
not ( n36383 , n36382 );
nand ( n36384 , n36379 , n36383 );
not ( n36385 , n36384 );
buf ( n36386 , RI1744d580_1359);
not ( n36387 , n36386 );
not ( n36388 , n204936 );
or ( n36389 , n36387 , n36388 );
not ( n36390 , RI1744d580_1359);
nand ( n36391 , n204939 , n36390 );
nand ( n36392 , n36389 , n36391 );
and ( n36393 , n36392 , n204978 );
not ( n36394 , n36392 );
and ( n36395 , n36394 , n204981 );
nor ( n36396 , n36393 , n36395 );
not ( n36397 , n36396 );
and ( n36398 , n36385 , n36397 );
not ( n36399 , n36396 );
not ( n36400 , n36399 );
and ( n36401 , n36384 , n36400 );
nor ( n36402 , n36398 , n36401 );
not ( n36403 , n36402 );
not ( n36404 , n36403 );
not ( n214166 , n205078 );
not ( n214167 , n32607 );
or ( n36407 , n214166 , n214167 );
not ( n36408 , n205078 );
nand ( n36409 , n36408 , n34763 );
nand ( n36410 , n36407 , n36409 );
not ( n36411 , n35021 );
and ( n36412 , n36410 , n36411 );
not ( n36413 , n36410 );
buf ( n36414 , n34807 );
not ( n36415 , n36414 );
and ( n36416 , n36413 , n36415 );
nor ( n36417 , n36412 , n36416 );
not ( n36418 , n36417 );
not ( n36419 , n36418 );
buf ( n36420 , n30838 );
not ( n36421 , n35054 );
xor ( n36422 , n35047 , n36421 );
xnor ( n36423 , n36422 , n35061 );
xor ( n36424 , n36420 , n36423 );
buf ( n36425 , RI173d5760_1715);
not ( n36426 , n36425 );
not ( n36427 , RI1738ca70_2070);
not ( n36428 , n36427 );
or ( n36429 , n36426 , n36428 );
not ( n36430 , RI173d5760_1715);
nand ( n36431 , n36430 , n26225 );
nand ( n36432 , n36429 , n36431 );
not ( n36433 , RI1744d238_1360);
and ( n36434 , n36432 , n36433 );
not ( n36435 , n36432 );
and ( n36436 , n36435 , n36095 );
nor ( n36437 , n36434 , n36436 );
buf ( n36438 , RI19aca4f0_2253);
nand ( n36439 , n25628 , n36438 );
buf ( n36440 , RI174bb878_827);
and ( n36441 , n36439 , n36440 );
not ( n36442 , n36439 );
not ( n36443 , RI174bb878_827);
and ( n36444 , n36442 , n36443 );
nor ( n36445 , n36441 , n36444 );
xor ( n36446 , n36437 , n36445 );
buf ( n36447 , RI19a9ad18_2606);
nand ( n36448 , n204916 , n36447 );
not ( n36449 , RI17471a48_1182);
and ( n36450 , n36448 , n36449 );
not ( n36451 , n36448 );
buf ( n36452 , RI17471a48_1182);
and ( n36453 , n36451 , n36452 );
nor ( n36454 , n36450 , n36453 );
xnor ( n36455 , n36446 , n36454 );
not ( n36456 , n36455 );
not ( n36457 , n36456 );
xnor ( n36458 , n36424 , n36457 );
not ( n36459 , n36458 );
buf ( n36460 , RI19ac5108_2291);
nand ( n36461 , n26242 , n36460 );
buf ( n36462 , RI174caff8_779);
and ( n36463 , n36461 , n36462 );
not ( n36464 , n36461 );
not ( n36465 , RI174caff8_779);
and ( n36466 , n36464 , n36465 );
nor ( n36467 , n36463 , n36466 );
buf ( n214229 , n36467 );
not ( n214230 , n214229 );
not ( n36470 , n33140 );
or ( n214232 , n214230 , n36470 );
or ( n214233 , n33140 , n214229 );
nand ( n36473 , n214232 , n214233 );
not ( n214235 , n30689 );
and ( n214236 , n36473 , n214235 );
not ( n36476 , n36473 );
and ( n36477 , n36476 , n30689 );
nor ( n36478 , n214236 , n36477 );
not ( n36479 , n36478 );
nand ( n36480 , n36459 , n36479 );
not ( n36481 , n36480 );
or ( n36482 , n36419 , n36481 );
nand ( n36483 , n36459 , n36479 );
or ( n36484 , n36483 , n36418 );
nand ( n36485 , n36482 , n36484 );
not ( n36486 , n36485 );
not ( n36487 , n29644 );
buf ( n36488 , RI173ea2c8_1614);
not ( n36489 , n36488 );
not ( n36490 , RI173a15d8_1969);
not ( n36491 , n36490 );
or ( n36492 , n36489 , n36491 );
not ( n36493 , RI173ea2c8_1614);
buf ( n36494 , RI173a15d8_1969);
nand ( n36495 , n36493 , n36494 );
nand ( n36496 , n36492 , n36495 );
not ( n36497 , RI1746a0e0_1219);
and ( n36498 , n36496 , n36497 );
not ( n36499 , n36496 );
buf ( n36500 , RI1746a0e0_1219);
and ( n36501 , n36499 , n36500 );
nor ( n36502 , n36498 , n36501 );
buf ( n36503 , RI19aa1438_2558);
nand ( n36504 , n26028 , n36503 );
not ( n36505 , RI174865b0_1081);
and ( n36506 , n36504 , n36505 );
not ( n36507 , n36504 );
buf ( n36508 , RI174865b0_1081);
and ( n36509 , n36507 , n36508 );
nor ( n36510 , n36506 , n36509 );
xor ( n36511 , n36502 , n36510 );
buf ( n36512 , RI19a82538_2778);
nand ( n36513 , n25711 , n36512 );
buf ( n36514 , RI1750cdd0_726);
and ( n36515 , n36513 , n36514 );
not ( n36516 , n36513 );
not ( n36517 , RI1750cdd0_726);
and ( n36518 , n36516 , n36517 );
nor ( n36519 , n36515 , n36518 );
xor ( n36520 , n36511 , n36519 );
not ( n36521 , n36520 );
or ( n36522 , n36487 , n36521 );
or ( n36523 , n36520 , n29644 );
nand ( n36524 , n36522 , n36523 );
nor ( n36525 , n36524 , n206425 );
not ( n36526 , n36525 );
nand ( n36527 , n28665 , n36524 );
nand ( n36528 , n36526 , n36527 );
not ( n36529 , n36528 );
not ( n36530 , n26490 );
not ( n36531 , n29814 );
or ( n36532 , n36530 , n36531 );
not ( n36533 , n26490 );
not ( n36534 , n29814 );
nand ( n36535 , n36533 , n36534 );
nand ( n36536 , n36532 , n36535 );
and ( n36537 , n36536 , n33577 );
not ( n36538 , n36536 );
and ( n36539 , n36538 , n29860 );
nor ( n36540 , n36537 , n36539 );
nand ( n36541 , n36529 , n36540 );
not ( n36542 , n36541 );
not ( n36543 , n31625 );
not ( n36544 , n26108 );
or ( n36545 , n36543 , n36544 );
or ( n36546 , n26108 , n31625 );
nand ( n36547 , n36545 , n36546 );
and ( n36548 , n36547 , n26149 );
not ( n36549 , n36547 );
and ( n36550 , n36549 , n26146 );
nor ( n36551 , n36548 , n36550 );
not ( n36552 , n36551 );
not ( n36553 , n36552 );
not ( n36554 , n36553 );
and ( n36555 , n36542 , n36554 );
and ( n36556 , n36541 , n36553 );
nor ( n36557 , n36555 , n36556 );
not ( n36558 , n36557 );
or ( n36559 , n36486 , n36558 );
or ( n36560 , n36557 , n36485 );
nand ( n36561 , n36559 , n36560 );
not ( n36562 , n36561 );
not ( n36563 , n36562 );
or ( n36564 , n36404 , n36563 );
nand ( n36565 , n36402 , n36561 );
nand ( n36566 , n36564 , n36565 );
not ( n36567 , n29052 );
not ( n36568 , n205766 );
not ( n36569 , n36568 );
or ( n36570 , n36567 , n36569 );
not ( n36571 , n29052 );
buf ( n36572 , n28004 );
not ( n36573 , n36572 );
nand ( n36574 , n36571 , n36573 );
nand ( n36575 , n36570 , n36574 );
and ( n36576 , n36575 , n32915 );
not ( n36577 , n36575 );
and ( n36578 , n36577 , n32916 );
nor ( n36579 , n36576 , n36578 );
not ( n36580 , n36579 );
not ( n36581 , n36580 );
not ( n36582 , n36581 );
not ( n36583 , RI174a3458_940);
and ( n36584 , n26220 , n36583 );
not ( n36585 , n26220 );
and ( n36586 , n36585 , n26217 );
nor ( n36587 , n36584 , n36586 );
not ( n36588 , n36587 );
not ( n36589 , n33565 );
or ( n36590 , n36588 , n36589 );
or ( n36591 , n33565 , n36587 );
nand ( n36592 , n36590 , n36591 );
buf ( n36593 , RI173ccd78_1757);
not ( n36594 , n36593 );
not ( n36595 , RI173437f8_2112);
not ( n36596 , n36595 );
or ( n36597 , n36594 , n36596 );
not ( n36598 , RI173ccd78_1757);
buf ( n36599 , RI173437f8_2112);
nand ( n36600 , n36598 , n36599 );
nand ( n36601 , n36597 , n36600 );
buf ( n36602 , RI17444bb0_1401);
and ( n36603 , n36601 , n36602 );
not ( n36604 , n36601 );
not ( n36605 , RI17444bb0_1401);
and ( n36606 , n36604 , n36605 );
nor ( n36607 , n36603 , n36606 );
not ( n36608 , n36607 );
buf ( n36609 , RI19a8d8c0_2700);
nand ( n36610 , n26325 , n36609 );
not ( n36611 , RI174693c0_1223);
and ( n36612 , n36610 , n36611 );
not ( n36613 , n36610 );
buf ( n36614 , RI174693c0_1223);
and ( n36615 , n36613 , n36614 );
nor ( n36616 , n36612 , n36615 );
xor ( n36617 , n36608 , n36616 );
xnor ( n36618 , n36617 , n35668 );
not ( n36619 , n36618 );
not ( n36620 , n36619 );
and ( n36621 , n36592 , n36620 );
not ( n36622 , n36592 );
xor ( n36623 , n36607 , n35667 );
not ( n36624 , n36616 );
xnor ( n36625 , n36623 , n36624 );
buf ( n36626 , n36625 );
and ( n36627 , n36622 , n36626 );
nor ( n36628 , n36621 , n36627 );
not ( n36629 , n36628 );
not ( n36630 , n205284 );
not ( n36631 , RI17394a68_2031);
not ( n36632 , n36631 );
or ( n36633 , n36630 , n36632 );
not ( n36634 , RI173dd758_1676);
buf ( n36635 , RI17394a68_2031);
nand ( n36636 , n36634 , n36635 );
nand ( n36637 , n36633 , n36636 );
and ( n36638 , n36637 , n35195 );
not ( n36639 , n36637 );
not ( n36640 , RI17455230_1321);
and ( n36641 , n36639 , n36640 );
nor ( n36642 , n36638 , n36641 );
not ( n36643 , n36642 );
buf ( n36644 , RI19ac6620_2282);
nand ( n36645 , n25711 , n36644 );
buf ( n36646 , RI174c86b8_787);
and ( n36647 , n36645 , n36646 );
not ( n36648 , n36645 );
not ( n36649 , RI174c86b8_787);
and ( n36650 , n36648 , n36649 );
nor ( n36651 , n36647 , n36650 );
xor ( n36652 , n36643 , n36651 );
buf ( n36653 , RI19a96740_2637);
nand ( n36654 , n25405 , n36653 );
buf ( n36655 , RI17479d88_1142);
and ( n36656 , n36654 , n36655 );
not ( n36657 , n36654 );
not ( n214419 , RI17479d88_1142);
and ( n214420 , n36657 , n214419 );
nor ( n36660 , n36656 , n214420 );
buf ( n214422 , n36660 );
xnor ( n36662 , n36652 , n214422 );
not ( n36663 , n36662 );
buf ( n36664 , n36663 );
xor ( n36665 , n25548 , n36664 );
xnor ( n36666 , n36665 , n33886 );
not ( n36667 , n36666 );
nand ( n36668 , n36629 , n36667 );
not ( n36669 , n36668 );
or ( n36670 , n36582 , n36669 );
or ( n36671 , n36668 , n36581 );
nand ( n36672 , n36670 , n36671 );
not ( n36673 , n36672 );
buf ( n36674 , n32039 );
not ( n36675 , n36674 );
not ( n36676 , n31213 );
or ( n36677 , n36675 , n36676 );
or ( n36678 , n31213 , n36674 );
nand ( n36679 , n36677 , n36678 );
and ( n36680 , n36679 , n31177 );
not ( n36681 , n36679 );
xor ( n36682 , n31158 , n208936 );
buf ( n36683 , n31166 );
xnor ( n36684 , n36682 , n36683 );
buf ( n36685 , n36684 );
and ( n36686 , n36681 , n36685 );
nor ( n36687 , n36680 , n36686 );
not ( n36688 , n36687 );
not ( n36689 , n36454 );
not ( n36690 , n26261 );
or ( n36691 , n36689 , n36690 );
not ( n36692 , n36454 );
nand ( n36693 , n36692 , n204681 );
nand ( n36694 , n36691 , n36693 );
and ( n36695 , n36694 , n26311 );
not ( n36696 , n36694 );
and ( n36697 , n36696 , n26319 );
nor ( n36698 , n36695 , n36697 );
nand ( n36699 , n36688 , n36698 );
not ( n36700 , n36699 );
not ( n36701 , n32875 );
not ( n36702 , n204744 );
not ( n36703 , n36702 );
or ( n36704 , n36701 , n36703 );
not ( n36705 , n204744 );
or ( n214467 , n36705 , n32875 );
nand ( n214468 , n36704 , n214467 );
not ( n36708 , n214468 );
xor ( n36709 , n31722 , n31695 );
xnor ( n36710 , n36709 , n31718 );
buf ( n214472 , n36710 );
not ( n214473 , n214472 );
and ( n36713 , n36708 , n214473 );
and ( n36714 , n214468 , n214472 );
nor ( n36715 , n36713 , n36714 );
not ( n36716 , n36715 );
not ( n36717 , n36716 );
and ( n36718 , n36700 , n36717 );
and ( n36719 , n36699 , n36716 );
nor ( n36720 , n36718 , n36719 );
not ( n36721 , n36720 );
and ( n36722 , n36673 , n36721 );
and ( n36723 , n36672 , n36720 );
nor ( n36724 , n36722 , n36723 );
and ( n36725 , n36566 , n36724 );
not ( n36726 , n36566 );
not ( n36727 , n36724 );
and ( n36728 , n36726 , n36727 );
nor ( n36729 , n36725 , n36728 );
buf ( n36730 , n36729 );
not ( n36731 , n36730 );
and ( n36732 , n36375 , n36731 );
and ( n36733 , n36374 , n36730 );
nor ( n36734 , n36732 , n36733 );
not ( n36735 , n31036 );
not ( n36736 , n36735 );
not ( n36737 , n36291 );
and ( n36738 , n36736 , n36737 );
and ( n36739 , n36735 , n36291 );
nor ( n36740 , n36738 , n36739 );
and ( n36741 , n36740 , n31078 );
not ( n36742 , n36740 );
and ( n36743 , n36742 , n31081 );
nor ( n36744 , n36741 , n36743 );
not ( n36745 , n36744 );
buf ( n36746 , RI17454858_1324);
not ( n36747 , n36746 );
xor ( n36748 , n30423 , n30440 );
buf ( n36749 , n30431 );
xnor ( n36750 , n36748 , n36749 );
buf ( n36751 , n36750 );
not ( n36752 , n36751 );
or ( n36753 , n36747 , n36752 );
or ( n36754 , n36751 , n36746 );
nand ( n36755 , n36753 , n36754 );
and ( n36756 , n36755 , n208210 );
not ( n36757 , n36755 );
not ( n36758 , n208210 );
and ( n36759 , n36757 , n36758 );
nor ( n36760 , n36756 , n36759 );
not ( n36761 , n36760 );
nand ( n36762 , n36745 , n36761 );
not ( n36763 , n36238 );
not ( n36764 , n32059 );
not ( n36765 , n31176 );
or ( n36766 , n36764 , n36765 );
or ( n36767 , n31176 , n32059 );
nand ( n36768 , n36766 , n36767 );
not ( n36769 , n36768 );
or ( n36770 , n36763 , n36769 );
or ( n36771 , n36768 , n36238 );
nand ( n36772 , n36770 , n36771 );
and ( n36773 , n36762 , n36772 );
not ( n36774 , n36762 );
not ( n36775 , n36772 );
and ( n36776 , n36774 , n36775 );
nor ( n36777 , n36773 , n36776 );
not ( n36778 , n36777 );
buf ( n36779 , RI173a4a58_1953);
not ( n36780 , n36779 );
not ( n36781 , RI173ed748_1598);
not ( n36782 , n36781 );
or ( n36783 , n36780 , n36782 );
not ( n36784 , RI173a4a58_1953);
buf ( n36785 , RI173ed748_1598);
nand ( n36786 , n36784 , n36785 );
nand ( n36787 , n36783 , n36786 );
not ( n36788 , RI1748c190_1053);
and ( n36789 , n36787 , n36788 );
not ( n36790 , n36787 );
buf ( n36791 , RI1748c190_1053);
and ( n36792 , n36790 , n36791 );
nor ( n36793 , n36789 , n36792 );
buf ( n36794 , RI19a9efa8_2577);
nand ( n36795 , n25479 , n36794 );
buf ( n36796 , RI17489a30_1065);
and ( n36797 , n36795 , n36796 );
not ( n36798 , n36795 );
not ( n36799 , RI17489a30_1065);
and ( n36800 , n36798 , n36799 );
nor ( n36801 , n36797 , n36800 );
xor ( n36802 , n36793 , n36801 );
buf ( n36803 , RI19acda60_2227);
nand ( n36804 , n27946 , n36803 );
buf ( n36805 , RI17512050_710);
and ( n36806 , n36804 , n36805 );
not ( n36807 , n36804 );
not ( n36808 , RI17512050_710);
and ( n36809 , n36807 , n36808 );
nor ( n36810 , n36806 , n36809 );
not ( n36811 , n36810 );
xnor ( n36812 , n36802 , n36811 );
buf ( n36813 , n36812 );
not ( n36814 , n36813 );
not ( n36815 , n36044 );
buf ( n36816 , RI173d0540_1740);
not ( n36817 , n36816 );
not ( n36818 , RI17346c78_2096);
not ( n36819 , n36818 );
or ( n36820 , n36817 , n36819 );
not ( n36821 , RI173d0540_1740);
buf ( n36822 , RI17346c78_2096);
nand ( n36823 , n36821 , n36822 );
nand ( n36824 , n36820 , n36823 );
buf ( n36825 , RI17448030_1385);
and ( n36826 , n36824 , n36825 );
not ( n36827 , n36824 );
not ( n36828 , RI17448030_1385);
and ( n36829 , n36827 , n36828 );
nor ( n36830 , n36826 , n36829 );
buf ( n36831 , RI19a8aad0_2720);
nand ( n36832 , n26242 , n36831 );
not ( n36833 , RI1746c840_1207);
and ( n36834 , n36832 , n36833 );
not ( n36835 , n36832 );
buf ( n36836 , RI1746c840_1207);
and ( n36837 , n36835 , n36836 );
nor ( n36838 , n36834 , n36837 );
xor ( n36839 , n36830 , n36838 );
buf ( n36840 , RI19abc4e0_2365);
nand ( n36841 , n27749 , n36840 );
not ( n36842 , RI174b5518_852);
and ( n36843 , n36841 , n36842 );
not ( n36844 , n36841 );
buf ( n36845 , RI174b5518_852);
and ( n36846 , n36844 , n36845 );
nor ( n36847 , n36843 , n36846 );
xnor ( n36848 , n36839 , n36847 );
buf ( n36849 , n36848 );
not ( n36850 , n36849 );
or ( n36851 , n36815 , n36850 );
or ( n36852 , n36849 , n36044 );
nand ( n36853 , n36851 , n36852 );
not ( n36854 , n36853 );
or ( n36855 , n36814 , n36854 );
or ( n36856 , n36853 , n36813 );
nand ( n36857 , n36855 , n36856 );
not ( n36858 , n36857 );
not ( n36859 , n34736 );
not ( n36860 , n36859 );
not ( n36861 , n36860 );
not ( n36862 , n31093 );
not ( n36863 , n34177 );
or ( n36864 , n36862 , n36863 );
or ( n36865 , n34179 , n31093 );
nand ( n36866 , n36864 , n36865 );
not ( n36867 , n36866 );
and ( n36868 , n36861 , n36867 );
and ( n36869 , n36860 , n36866 );
nor ( n36870 , n36868 , n36869 );
not ( n36871 , n36870 );
nand ( n36872 , n36858 , n36871 );
not ( n36873 , n36872 );
buf ( n36874 , RI19ac1670_2319);
nand ( n36875 , n32338 , n36874 );
not ( n36876 , RI174acb48_894);
and ( n36877 , n36875 , n36876 );
not ( n214639 , n36875 );
buf ( n214640 , RI174acb48_894);
and ( n36880 , n214639 , n214640 );
nor ( n36881 , n36877 , n36880 );
not ( n36882 , n36881 );
not ( n36883 , n28907 );
not ( n36884 , n36883 );
or ( n36885 , n36882 , n36884 );
not ( n36886 , n36881 );
not ( n36887 , n28906 );
nand ( n36888 , n36886 , n36887 );
nand ( n36889 , n36885 , n36888 );
buf ( n36890 , n30936 );
and ( n36891 , n36889 , n36890 );
not ( n36892 , n36889 );
and ( n36893 , n36892 , n30943 );
nor ( n36894 , n36891 , n36893 );
not ( n36895 , n36894 );
not ( n36896 , n36895 );
and ( n36897 , n36873 , n36896 );
and ( n36898 , n36872 , n36895 );
nor ( n36899 , n36897 , n36898 );
not ( n36900 , n36899 );
buf ( n36901 , RI173cfeb0_1742);
not ( n36902 , n36901 );
not ( n36903 , RI173465e8_2098);
not ( n36904 , n36903 );
or ( n36905 , n36902 , n36904 );
not ( n36906 , RI173cfeb0_1742);
buf ( n36907 , RI173465e8_2098);
nand ( n36908 , n36906 , n36907 );
nand ( n36909 , n36905 , n36908 );
not ( n36910 , RI174479a0_1387);
and ( n36911 , n36909 , n36910 );
not ( n36912 , n36909 );
buf ( n36913 , RI174479a0_1387);
and ( n36914 , n36912 , n36913 );
nor ( n36915 , n36911 , n36914 );
buf ( n36916 , RI19a8a878_2721);
nand ( n36917 , n28238 , n36916 );
buf ( n36918 , RI1746c1b0_1209);
and ( n36919 , n36917 , n36918 );
not ( n36920 , n36917 );
not ( n36921 , RI1746c1b0_1209);
and ( n36922 , n36920 , n36921 );
nor ( n36923 , n36919 , n36922 );
xor ( n36924 , n36915 , n36923 );
buf ( n36925 , RI19abc378_2366);
nand ( n36926 , n25803 , n36925 );
buf ( n36927 , RI174b4e88_854);
and ( n36928 , n36926 , n36927 );
not ( n36929 , n36926 );
not ( n36930 , RI174b4e88_854);
and ( n36931 , n36929 , n36930 );
nor ( n36932 , n36928 , n36931 );
not ( n36933 , n36932 );
xnor ( n36934 , n36924 , n36933 );
xor ( n36935 , n28136 , n36934 );
buf ( n36936 , RI173fb9b0_1529);
not ( n36937 , n36936 );
not ( n36938 , n32187 );
or ( n36939 , n36937 , n36938 );
not ( n36940 , RI173fb9b0_1529);
buf ( n36941 , RI173b2978_1885);
nand ( n36942 , n36940 , n36941 );
nand ( n36943 , n36939 , n36942 );
not ( n36944 , n36943 );
not ( n36945 , RI173a0570_1974);
buf ( n36946 , RI19a8b958_2714);
nand ( n36947 , n25751 , n36946 );
buf ( n36948 , RI17528418_641);
and ( n36949 , n36947 , n36948 );
not ( n36950 , n36947 );
not ( n214712 , RI17528418_641);
and ( n214713 , n36950 , n214712 );
nor ( n36953 , n36949 , n214713 );
xor ( n214715 , n36945 , n36953 );
buf ( n214716 , RI19aa8080_2509);
nand ( n36956 , n25666 , n214716 );
not ( n36957 , RI17497c98_996);
and ( n36958 , n36956 , n36957 );
not ( n36959 , n36956 );
buf ( n36960 , RI17497c98_996);
and ( n36961 , n36959 , n36960 );
nor ( n36962 , n36958 , n36961 );
xnor ( n36963 , n214715 , n36962 );
not ( n36964 , n36963 );
or ( n36965 , n36944 , n36964 );
not ( n36966 , n36963 );
not ( n36967 , n36943 );
nand ( n36968 , n36966 , n36967 );
nand ( n36969 , n36965 , n36968 );
not ( n36970 , n36969 );
xnor ( n36971 , n36935 , n36970 );
not ( n36972 , n36971 );
buf ( n36973 , RI173a7ed8_1937);
not ( n36974 , n36973 );
not ( n36975 , n25963 );
or ( n36976 , n36974 , n36975 );
or ( n36977 , n25963 , n36973 );
nand ( n36978 , n36976 , n36977 );
not ( n36979 , n36978 );
not ( n36980 , n25457 );
or ( n36981 , n36979 , n36980 );
buf ( n36982 , n25456 );
not ( n36983 , n36982 );
or ( n36984 , n36983 , n36978 );
nand ( n36985 , n36981 , n36984 );
not ( n36986 , n36985 );
nand ( n36987 , n36972 , n36986 );
not ( n36988 , n205311 );
xor ( n36989 , n34854 , n212623 );
xnor ( n36990 , n36989 , n34871 );
not ( n36991 , n36990 );
or ( n36992 , n36988 , n36991 );
or ( n36993 , n36990 , n205311 );
nand ( n36994 , n36992 , n36993 );
buf ( n36995 , RI173fafd8_1532);
not ( n36996 , n36995 );
not ( n36997 , RI173b22e8_1887);
not ( n36998 , n36997 );
or ( n36999 , n36996 , n36998 );
not ( n37000 , RI173fafd8_1532);
buf ( n37001 , RI173b22e8_1887);
nand ( n37002 , n37000 , n37001 );
nand ( n37003 , n36999 , n37002 );
buf ( n37004 , RI1739de10_1986);
and ( n37005 , n37003 , n37004 );
not ( n37006 , n37003 );
not ( n37007 , RI1739de10_1986);
and ( n37008 , n37006 , n37007 );
nor ( n37009 , n37005 , n37008 );
xor ( n37010 , n37009 , n28156 );
buf ( n37011 , RI19aa29c8_2548);
nand ( n37012 , n28238 , n37011 );
not ( n37013 , RI175279c8_643);
and ( n37014 , n37012 , n37013 );
not ( n37015 , n37012 );
buf ( n37016 , RI175279c8_643);
and ( n37017 , n37015 , n37016 );
nor ( n37018 , n37014 , n37017 );
xnor ( n37019 , n37010 , n37018 );
not ( n37020 , n37019 );
and ( n37021 , n36994 , n37020 );
not ( n37022 , n36994 );
not ( n37023 , n37020 );
and ( n37024 , n37022 , n37023 );
nor ( n37025 , n37021 , n37024 );
and ( n37026 , n36987 , n37025 );
not ( n37027 , n36987 );
not ( n37028 , n37025 );
and ( n37029 , n37027 , n37028 );
nor ( n37030 , n37026 , n37029 );
not ( n37031 , n37030 );
or ( n37032 , n36900 , n37031 );
or ( n37033 , n37030 , n36899 );
nand ( n37034 , n37032 , n37033 );
not ( n37035 , n33397 );
buf ( n37036 , RI173fe458_1516);
not ( n37037 , n37036 );
not ( n37038 , RI173b5420_1872);
not ( n37039 , n37038 );
or ( n37040 , n37037 , n37039 );
not ( n37041 , RI173fe458_1516);
buf ( n37042 , RI173b5420_1872);
nand ( n37043 , n37041 , n37042 );
nand ( n37044 , n37040 , n37043 );
not ( n37045 , n37044 );
not ( n37046 , n37045 );
or ( n37047 , n37035 , n37046 );
not ( n37048 , RI1733a798_2156);
nand ( n37049 , n37044 , n37048 );
nand ( n37050 , n37047 , n37049 );
not ( n37051 , RI173bb9d8_1841);
buf ( n37052 , RI19a88a00_2734);
nand ( n37053 , n25656 , n37052 );
buf ( n37054 , RI1752c720_628);
and ( n37055 , n37053 , n37054 );
not ( n37056 , n37053 );
not ( n37057 , RI1752c720_628);
and ( n37058 , n37056 , n37057 );
nor ( n37059 , n37055 , n37058 );
xor ( n37060 , n37051 , n37059 );
buf ( n37061 , RI19aa7888_2513);
nand ( n37062 , n25628 , n37061 );
buf ( n37063 , RI1749a740_983);
and ( n37064 , n37062 , n37063 );
not ( n37065 , n37062 );
not ( n37066 , RI1749a740_983);
and ( n37067 , n37065 , n37066 );
nor ( n37068 , n37064 , n37067 );
xnor ( n37069 , n37060 , n37068 );
not ( n37070 , n37069 );
and ( n37071 , n37050 , n37070 );
not ( n37072 , n37050 );
and ( n37073 , n37072 , n37069 );
or ( n37074 , n37071 , n37073 );
not ( n37075 , n29351 );
not ( n37076 , RI17389fc8_2083);
not ( n37077 , n37076 );
or ( n37078 , n37075 , n37077 );
not ( n37079 , RI173d2cb8_1728);
buf ( n37080 , RI17389fc8_2083);
nand ( n37081 , n37079 , n37080 );
nand ( n37082 , n37078 , n37081 );
not ( n37083 , RI1744a790_1373);
and ( n37084 , n37082 , n37083 );
not ( n37085 , n37082 );
and ( n37086 , n37085 , n35290 );
nor ( n37087 , n37084 , n37086 );
buf ( n37088 , RI19abb748_2371);
nand ( n37089 , n27946 , n37088 );
buf ( n37090 , RI174b7c78_840);
and ( n37091 , n37089 , n37090 );
not ( n37092 , n37089 );
not ( n37093 , RI174b7c78_840);
and ( n37094 , n37092 , n37093 );
nor ( n37095 , n37091 , n37094 );
xor ( n37096 , n37087 , n37095 );
buf ( n37097 , RI19a89bd0_2726);
nand ( n37098 , n26162 , n37097 );
buf ( n37099 , RI1746efa0_1195);
and ( n37100 , n37098 , n37099 );
not ( n37101 , n37098 );
not ( n37102 , RI1746efa0_1195);
and ( n37103 , n37101 , n37102 );
nor ( n37104 , n37100 , n37103 );
xnor ( n37105 , n37096 , n37104 );
buf ( n37106 , n37105 );
and ( n37107 , n37074 , n37106 );
not ( n214869 , n37074 );
not ( n214870 , n37106 );
and ( n37110 , n214869 , n214870 );
nor ( n37111 , n37107 , n37110 );
buf ( n37112 , n37111 );
not ( n37113 , n37112 );
not ( n37114 , n204404 );
xor ( n37115 , n34971 , n34978 );
xnor ( n37116 , n37115 , n34984 );
not ( n37117 , n37116 );
or ( n37118 , n37114 , n37117 );
not ( n37119 , n204404 );
not ( n37120 , n37116 );
nand ( n37121 , n37119 , n37120 );
nand ( n37122 , n37118 , n37121 );
buf ( n37123 , n35017 );
and ( n37124 , n37122 , n37123 );
not ( n37125 , n37122 );
xor ( n37126 , n34998 , n35015 );
xor ( n37127 , n37126 , n35219 );
buf ( n37128 , n37127 );
and ( n37129 , n37125 , n37128 );
nor ( n37130 , n37124 , n37129 );
not ( n37131 , n32539 );
not ( n37132 , n28462 );
or ( n37133 , n37131 , n37132 );
or ( n37134 , n28462 , n32539 );
nand ( n37135 , n37133 , n37134 );
and ( n37136 , n37135 , n28502 );
not ( n37137 , n37135 );
and ( n37138 , n37137 , n206271 );
nor ( n37139 , n37136 , n37138 );
not ( n37140 , n37139 );
nand ( n37141 , n37130 , n37140 );
not ( n37142 , n37141 );
or ( n37143 , n37113 , n37142 );
or ( n37144 , n37141 , n37112 );
nand ( n37145 , n37143 , n37144 );
not ( n37146 , n37145 );
not ( n37147 , n31480 );
buf ( n37148 , RI173efb60_1587);
not ( n37149 , n37148 );
not ( n37150 , RI173a6e70_1942);
not ( n37151 , n37150 );
or ( n37152 , n37149 , n37151 );
not ( n37153 , RI173efb60_1587);
nand ( n37154 , n37153 , n33712 );
nand ( n37155 , n37152 , n37154 );
and ( n37156 , n37155 , n205232 );
not ( n37157 , n37155 );
not ( n37158 , RI174a2dc8_942);
and ( n37159 , n37157 , n37158 );
nor ( n37160 , n37156 , n37159 );
not ( n37161 , n37160 );
buf ( n37162 , RI19accc50_2233);
nand ( n37163 , n204336 , n37162 );
buf ( n37164 , RI17515e30_698);
and ( n37165 , n37163 , n37164 );
not ( n37166 , n37163 );
not ( n37167 , RI17515e30_698);
and ( n37168 , n37166 , n37167 );
nor ( n37169 , n37165 , n37168 );
xor ( n37170 , n37161 , n37169 );
xnor ( n37171 , n37170 , n25822 );
not ( n37172 , n37171 );
not ( n37173 , n37172 );
or ( n37174 , n37147 , n37173 );
not ( n37175 , n31480 );
nand ( n37176 , n37175 , n37171 );
nand ( n37177 , n37174 , n37176 );
buf ( n37178 , RI17457990_1309);
not ( n37179 , RI1740d098_1444);
and ( n37180 , n37179 , n31945 );
not ( n37181 , n37179 );
not ( n37182 , RI173c43a8_1799);
and ( n37183 , n37181 , n37182 );
nor ( n37184 , n37180 , n37183 );
xor ( n37185 , n37178 , n37184 );
buf ( n37186 , RI1733ae28_2154);
buf ( n37187 , RI174a96c8_910);
xor ( n37188 , n37186 , n37187 );
buf ( n37189 , RI19ab1ba8_2441);
nand ( n37190 , n25622 , n37189 );
xnor ( n37191 , n37188 , n37190 );
xnor ( n37192 , n37185 , n37191 );
buf ( n37193 , n37192 );
and ( n37194 , n37177 , n37193 );
not ( n37195 , n37177 );
not ( n37196 , n37193 );
and ( n37197 , n37195 , n37196 );
nor ( n37198 , n37194 , n37197 );
not ( n37199 , n204609 );
not ( n37200 , n204617 );
not ( n37201 , n30255 );
and ( n37202 , n37200 , n37201 );
and ( n37203 , n204617 , n30255 );
nor ( n37204 , n37202 , n37203 );
not ( n37205 , n37204 );
and ( n37206 , n37199 , n37205 );
and ( n37207 , n204609 , n37204 );
nor ( n37208 , n37206 , n37207 );
not ( n37209 , n37208 );
xor ( n37210 , n35509 , n35517 );
xnor ( n37211 , n37210 , n35526 );
buf ( n37212 , n37211 );
not ( n214974 , n37212 );
and ( n214975 , n37209 , n214974 );
and ( n37215 , n37208 , n37212 );
nor ( n37216 , n214975 , n37215 );
nand ( n37217 , n37198 , n37216 );
not ( n37218 , n37217 );
not ( n37219 , n28105 );
xor ( n37220 , n25404 , n25424 );
not ( n37221 , n25413 );
xnor ( n37222 , n37220 , n37221 );
not ( n37223 , n37222 );
or ( n37224 , n37219 , n37223 );
or ( n37225 , n28105 , n37222 );
nand ( n37226 , n37224 , n37225 );
and ( n37227 , n37226 , n28680 );
not ( n37228 , n37226 );
not ( n37229 , n206437 );
and ( n37230 , n37228 , n37229 );
nor ( n37231 , n37227 , n37230 );
not ( n37232 , n37231 );
not ( n37233 , n37232 );
and ( n37234 , n37218 , n37233 );
nand ( n37235 , n37216 , n37198 );
and ( n37236 , n37235 , n37232 );
nor ( n37237 , n37234 , n37236 );
not ( n37238 , n37237 );
or ( n37239 , n37146 , n37238 );
or ( n37240 , n37145 , n37237 );
nand ( n37241 , n37239 , n37240 );
nand ( n37242 , n36744 , n36775 );
not ( n37243 , n37242 );
buf ( n37244 , RI1740d728_1442);
not ( n37245 , n33012 );
not ( n37246 , RI173bd760_1832);
not ( n37247 , n37246 );
or ( n37248 , n37245 , n37247 );
not ( n37249 , RI17406450_1477);
buf ( n37250 , RI173bd760_1832);
nand ( n37251 , n37249 , n37250 );
nand ( n37252 , n37248 , n37251 );
xor ( n37253 , n37244 , n37252 );
buf ( n37254 , RI173341e0_2187);
not ( n37255 , RI174a2738_944);
xor ( n37256 , n37254 , n37255 );
buf ( n37257 , RI19ab4740_2420);
nand ( n37258 , n204426 , n37257 );
xnor ( n37259 , n37256 , n37258 );
xnor ( n37260 , n37253 , n37259 );
not ( n37261 , n37260 );
not ( n37262 , n37261 );
not ( n37263 , n32277 );
not ( n37264 , n29561 );
or ( n37265 , n37263 , n37264 );
or ( n37266 , n29561 , n32277 );
nand ( n37267 , n37265 , n37266 );
not ( n37268 , n37267 );
and ( n37269 , n37262 , n37268 );
not ( n215031 , n37261 );
not ( n215032 , n215031 );
and ( n37272 , n215032 , n37267 );
nor ( n37273 , n37269 , n37272 );
not ( n37274 , n37273 );
not ( n37275 , n37274 );
and ( n37276 , n37243 , n37275 );
and ( n37277 , n37242 , n37274 );
nor ( n37278 , n37276 , n37277 );
and ( n37279 , n37241 , n37278 );
not ( n37280 , n37241 );
not ( n37281 , n37278 );
and ( n37282 , n37280 , n37281 );
nor ( n37283 , n37279 , n37282 );
not ( n37284 , n37283 );
and ( n37285 , n37034 , n37284 );
not ( n37286 , n37034 );
and ( n37287 , n37286 , n37283 );
nor ( n37288 , n37285 , n37287 );
not ( n37289 , n37288 );
not ( n37290 , n37289 );
not ( n37291 , n37290 );
or ( n37292 , n36778 , n37291 );
not ( n37293 , n36777 );
nand ( n37294 , n37289 , n37293 );
nand ( n37295 , n37292 , n37294 );
buf ( n37296 , n31472 );
not ( n37297 , n37296 );
xor ( n37298 , n211219 , n37297 );
xnor ( n37299 , n37298 , n32363 );
buf ( n37300 , n204304 );
not ( n37301 , n37300 );
not ( n37302 , n30442 );
not ( n37303 , n37302 );
not ( n37304 , n37303 );
or ( n37305 , n37301 , n37304 );
or ( n37306 , n30442 , n37300 );
nand ( n37307 , n37305 , n37306 );
and ( n37308 , n37307 , n36758 );
not ( n37309 , n37307 );
and ( n37310 , n37309 , n208210 );
nor ( n37311 , n37308 , n37310 );
nand ( n37312 , n37299 , n37311 );
not ( n37313 , n32226 );
buf ( n37314 , RI173fbcf8_1528);
not ( n37315 , n37314 );
not ( n37316 , RI173b2cc0_1884);
not ( n37317 , n37316 );
or ( n37318 , n37315 , n37317 );
not ( n37319 , RI173fbcf8_1528);
buf ( n37320 , RI173b2cc0_1884);
nand ( n37321 , n37319 , n37320 );
nand ( n37322 , n37318 , n37321 );
not ( n37323 , RI173a2988_1963);
and ( n37324 , n37322 , n37323 );
not ( n37325 , n37322 );
buf ( n37326 , RI173a2988_1963);
and ( n37327 , n37325 , n37326 );
nor ( n37328 , n37324 , n37327 );
buf ( n37329 , RI19aa81e8_2508);
nand ( n37330 , n204572 , n37329 );
buf ( n37331 , RI17497fe0_995);
and ( n37332 , n37330 , n37331 );
not ( n37333 , n37330 );
not ( n37334 , RI17497fe0_995);
and ( n37335 , n37333 , n37334 );
nor ( n37336 , n37332 , n37335 );
xor ( n37337 , n37328 , n37336 );
buf ( n37338 , RI19a8d230_2703);
nand ( n37339 , n25803 , n37338 );
buf ( n37340 , RI17528940_640);
and ( n37341 , n37339 , n37340 );
not ( n37342 , n37339 );
not ( n37343 , RI17528940_640);
and ( n215105 , n37342 , n37343 );
nor ( n215106 , n37341 , n215105 );
xor ( n37346 , n37337 , n215106 );
buf ( n37347 , n37346 );
not ( n37348 , n37347 );
or ( n37349 , n37313 , n37348 );
or ( n37350 , n37347 , n32226 );
nand ( n37351 , n37349 , n37350 );
not ( n37352 , n36848 );
not ( n37353 , n37352 );
and ( n37354 , n37351 , n37353 );
not ( n37355 , n37351 );
not ( n37356 , n36849 );
and ( n37357 , n37355 , n37356 );
nor ( n37358 , n37354 , n37357 );
and ( n37359 , n37312 , n37358 );
not ( n37360 , n37312 );
not ( n37361 , n37358 );
and ( n37362 , n37360 , n37361 );
nor ( n37363 , n37359 , n37362 );
not ( n37364 , n28573 );
buf ( n37365 , RI173e98f0_1617);
not ( n37366 , n37365 );
not ( n37367 , RI173a0c00_1972);
not ( n37368 , n37367 );
or ( n37369 , n37366 , n37368 );
not ( n37370 , RI173e98f0_1617);
buf ( n37371 , RI173a0c00_1972);
nand ( n37372 , n37370 , n37371 );
nand ( n37373 , n37369 , n37372 );
not ( n37374 , RI17463498_1252);
and ( n37375 , n37373 , n37374 );
not ( n37376 , n37373 );
buf ( n37377 , RI17463498_1252);
and ( n215139 , n37376 , n37377 );
nor ( n215140 , n37375 , n215139 );
buf ( n37380 , RI19acfb30_2213);
nand ( n215142 , n26453 , n37380 );
buf ( n215143 , RI1750be58_729);
and ( n37383 , n215142 , n215143 );
not ( n37384 , n215142 );
not ( n37385 , RI1750be58_729);
and ( n37386 , n37384 , n37385 );
nor ( n37387 , n37383 , n37386 );
xor ( n37388 , n215140 , n37387 );
buf ( n37389 , RI19aa0d30_2562);
nand ( n37390 , n29203 , n37389 );
not ( n37391 , RI17485bd8_1084);
and ( n37392 , n37390 , n37391 );
not ( n37393 , n37390 );
buf ( n37394 , RI17485bd8_1084);
and ( n37395 , n37393 , n37394 );
nor ( n37396 , n37392 , n37395 );
xnor ( n37397 , n37388 , n37396 );
buf ( n37398 , n37397 );
not ( n37399 , n37398 );
or ( n37400 , n37364 , n37399 );
or ( n37401 , n37398 , n28573 );
nand ( n37402 , n37400 , n37401 );
not ( n37403 , n37402 );
not ( n37404 , n30810 );
and ( n37405 , n37403 , n37404 );
not ( n37406 , n30808 );
buf ( n37407 , n37406 );
and ( n37408 , n37402 , n37407 );
nor ( n37409 , n37405 , n37408 );
buf ( n37410 , n34641 );
not ( n37411 , RI1749c4c8_974);
and ( n37412 , n37410 , n37411 );
not ( n37413 , n37410 );
and ( n37414 , n37413 , n34638 );
or ( n37415 , n37412 , n37414 );
not ( n37416 , n37415 );
buf ( n37417 , RI173f15a0_1579);
not ( n37418 , n37417 );
not ( n37419 , RI173a88b0_1934);
not ( n37420 , n37419 );
or ( n37421 , n37418 , n37420 );
not ( n37422 , RI173f15a0_1579);
buf ( n37423 , RI173a88b0_1934);
nand ( n37424 , n37422 , n37423 );
nand ( n37425 , n37421 , n37424 );
not ( n37426 , RI174b2db8_864);
and ( n37427 , n37425 , n37426 );
not ( n37428 , n37425 );
buf ( n37429 , RI174b2db8_864);
and ( n37430 , n37428 , n37429 );
nor ( n37431 , n37427 , n37430 );
buf ( n37432 , RI19aa40c0_2537);
nand ( n37433 , n25451 , n37432 );
buf ( n37434 , RI17518770_690);
and ( n37435 , n37433 , n37434 );
not ( n37436 , n37433 );
not ( n37437 , RI17518770_690);
and ( n37438 , n37436 , n37437 );
nor ( n37439 , n37435 , n37438 );
xor ( n37440 , n37431 , n37439 );
buf ( n37441 , RI19ab03c0_2452);
nand ( n37442 , n25628 , n37441 );
not ( n37443 , RI1748d888_1046);
and ( n37444 , n37442 , n37443 );
not ( n37445 , n37442 );
buf ( n37446 , RI1748d888_1046);
and ( n37447 , n37445 , n37446 );
nor ( n37448 , n37444 , n37447 );
xnor ( n37449 , n37440 , n37448 );
not ( n37450 , n37449 );
not ( n37451 , n37450 );
or ( n37452 , n37416 , n37451 );
or ( n37453 , n37450 , n37415 );
nand ( n37454 , n37452 , n37453 );
buf ( n37455 , n210489 );
and ( n37456 , n37454 , n37455 );
not ( n37457 , n37454 );
not ( n37458 , n37455 );
and ( n37459 , n37457 , n37458 );
nor ( n37460 , n37456 , n37459 );
nand ( n37461 , n37409 , n37460 );
not ( n37462 , n37461 );
not ( n37463 , n204833 );
not ( n37464 , n28876 );
not ( n37465 , n37464 );
or ( n37466 , n37463 , n37465 );
or ( n37467 , n37464 , n204833 );
nand ( n37468 , n37466 , n37467 );
buf ( n37469 , n211807 );
and ( n37470 , n37468 , n37469 );
not ( n37471 , n37468 );
buf ( n37472 , n34051 );
and ( n37473 , n37471 , n37472 );
nor ( n37474 , n37470 , n37473 );
not ( n37475 , n37474 );
not ( n37476 , n37475 );
and ( n37477 , n37462 , n37476 );
and ( n37478 , n37461 , n37475 );
nor ( n37479 , n37477 , n37478 );
nand ( n37480 , n37363 , n37479 );
not ( n37481 , n37480 );
nor ( n37482 , n37363 , n37479 );
nor ( n37483 , n37481 , n37482 );
not ( n37484 , n37483 );
buf ( n37485 , n208507 );
not ( n37486 , n37485 );
xor ( n37487 , n31630 , n31634 );
xnor ( n37488 , n37487 , n26067 );
not ( n37489 , n37488 );
or ( n37490 , n37486 , n37489 );
or ( n37491 , n37488 , n37485 );
nand ( n37492 , n37490 , n37491 );
not ( n37493 , n37492 );
buf ( n215255 , RI173d2628_1730);
not ( n215256 , RI17400870_1505);
buf ( n37496 , RI173b7b80_1860);
and ( n37497 , n215256 , n37496 );
not ( n37498 , n215256 );
not ( n37499 , RI173b7b80_1860);
and ( n37500 , n37498 , n37499 );
nor ( n37501 , n37497 , n37500 );
xor ( n37502 , n215255 , n37501 );
buf ( n37503 , RI1752ffd8_617);
xor ( n37504 , n37503 , n35304 );
xnor ( n37505 , n37504 , n35307 );
xnor ( n37506 , n37502 , n37505 );
not ( n37507 , n37506 );
not ( n37508 , n37507 );
or ( n37509 , n37493 , n37508 );
not ( n37510 , n37506 );
or ( n37511 , n37510 , n37492 );
nand ( n37512 , n37509 , n37511 );
buf ( n37513 , RI1746e910_1197);
not ( n37514 , n37513 );
not ( n37515 , n28646 );
or ( n37516 , n37514 , n37515 );
or ( n37517 , n28646 , n37513 );
nand ( n37518 , n37516 , n37517 );
and ( n37519 , n37518 , n32457 );
not ( n37520 , n37518 );
and ( n37521 , n37520 , n32454 );
nor ( n37522 , n37519 , n37521 );
nand ( n37523 , n37512 , n37522 );
not ( n37524 , n37523 );
not ( n37525 , n32849 );
not ( n37526 , n35857 );
not ( n37527 , n37526 );
or ( n37528 , n37525 , n37527 );
not ( n37529 , n35857 );
or ( n37530 , n37529 , n32849 );
nand ( n37531 , n37528 , n37530 );
not ( n37532 , n30078 );
not ( n37533 , n37532 );
and ( n37534 , n37531 , n37533 );
not ( n37535 , n37531 );
xor ( n37536 , n207820 , n30067 );
xnor ( n37537 , n37536 , n30077 );
not ( n37538 , n37537 );
not ( n37539 , n37538 );
and ( n37540 , n37535 , n37539 );
nor ( n37541 , n37534 , n37540 );
not ( n37542 , n37541 );
not ( n37543 , n37542 );
and ( n37544 , n37524 , n37543 );
not ( n37545 , n37541 );
and ( n37546 , n37523 , n37545 );
nor ( n37547 , n37544 , n37546 );
not ( n37548 , n37547 );
buf ( n37549 , RI174a5528_930);
buf ( n37550 , RI19accea8_2232);
nand ( n37551 , n30640 , n37550 );
buf ( n37552 , RI17516880_696);
and ( n37553 , n37551 , n37552 );
not ( n37554 , n37551 );
not ( n37555 , RI17516880_696);
and ( n37556 , n37554 , n37555 );
nor ( n37557 , n37553 , n37556 );
xor ( n37558 , n37549 , n37557 );
xnor ( n37559 , n37558 , n35457 );
buf ( n37560 , n37559 );
not ( n37561 , n37560 );
not ( n37562 , RI173f01f0_1585);
not ( n37563 , n37562 );
not ( n37564 , n205690 );
and ( n37565 , n37563 , n37564 );
and ( n37566 , n205690 , n37562 );
nor ( n37567 , n37565 , n37566 );
not ( n37568 , n37567 );
not ( n37569 , n25830 );
and ( n37570 , n37568 , n37569 );
and ( n37571 , n37567 , n25830 );
nor ( n37572 , n37570 , n37571 );
not ( n37573 , n37572 );
and ( n37574 , n37561 , n37573 );
and ( n37575 , n37560 , n37572 );
nor ( n37576 , n37574 , n37575 );
not ( n37577 , n204465 );
xor ( n37578 , n204456 , n37577 );
xnor ( n37579 , n37578 , n204472 );
not ( n37580 , n37579 );
not ( n37581 , n37580 );
and ( n37582 , n37576 , n37581 );
not ( n37583 , n37576 );
and ( n37584 , n37583 , n37580 );
nor ( n37585 , n37582 , n37584 );
not ( n37586 , n37585 );
not ( n37587 , n37586 );
buf ( n37588 , n29333 );
not ( n37589 , n37588 );
not ( n37590 , n205419 );
or ( n37591 , n37589 , n37590 );
or ( n37592 , n205419 , n37588 );
nand ( n37593 , n37591 , n37592 );
xor ( n37594 , n37593 , n205434 );
not ( n37595 , n25608 );
buf ( n37596 , RI173fd0a8_1522);
not ( n37597 , n37596 );
not ( n37598 , RI173b4070_1878);
not ( n37599 , n37598 );
or ( n37600 , n37597 , n37599 );
not ( n37601 , RI173fd0a8_1522);
buf ( n37602 , RI173b4070_1878);
nand ( n37603 , n37601 , n37602 );
nand ( n37604 , n37600 , n37603 );
not ( n37605 , RI173b0218_1897);
and ( n37606 , n37604 , n37605 );
not ( n37607 , n37604 );
and ( n37608 , n37607 , n31091 );
nor ( n37609 , n37606 , n37608 );
xor ( n37610 , n37609 , n35476 );
buf ( n37611 , RI19aa9430_2501);
nand ( n37612 , n27749 , n37611 );
buf ( n37613 , RI17499390_989);
and ( n37614 , n37612 , n37613 );
not ( n37615 , n37612 );
not ( n37616 , RI17499390_989);
and ( n37617 , n37615 , n37616 );
nor ( n37618 , n37614 , n37617 );
xor ( n37619 , n37610 , n37618 );
not ( n37620 , n37619 );
or ( n37621 , n37595 , n37620 );
or ( n37622 , n37619 , n25608 );
nand ( n37623 , n37621 , n37622 );
buf ( n37624 , RI173d1908_1734);
not ( n37625 , n37624 );
not ( n37626 , RI17359350_2090);
not ( n37627 , n37626 );
or ( n37628 , n37625 , n37627 );
not ( n37629 , RI173d1908_1734);
buf ( n37630 , RI17359350_2090);
nand ( n37631 , n37629 , n37630 );
nand ( n37632 , n37628 , n37631 );
not ( n37633 , RI174493e0_1379);
and ( n37634 , n37632 , n37633 );
not ( n37635 , n37632 );
buf ( n37636 , RI174493e0_1379);
and ( n37637 , n37635 , n37636 );
nor ( n37638 , n37634 , n37637 );
xor ( n37639 , n37638 , n29663 );
buf ( n37640 , RI19a89018_2731);
nand ( n37641 , n28238 , n37640 );
buf ( n37642 , RI1746dbf0_1201);
and ( n37643 , n37641 , n37642 );
not ( n37644 , n37641 );
not ( n37645 , RI1746dbf0_1201);
and ( n37646 , n37644 , n37645 );
nor ( n37647 , n37643 , n37646 );
xnor ( n37648 , n37639 , n37647 );
buf ( n37649 , n37648 );
and ( n37650 , n37623 , n37649 );
not ( n37651 , n37623 );
not ( n37652 , n37648 );
and ( n37653 , n37651 , n37652 );
nor ( n37654 , n37650 , n37653 );
not ( n215416 , n37654 );
nand ( n215417 , n37594 , n215416 );
not ( n37657 , n215417 );
or ( n37658 , n37587 , n37657 );
nand ( n37659 , n37594 , n215416 );
or ( n37660 , n37659 , n37586 );
nand ( n37661 , n37658 , n37660 );
not ( n37662 , n37661 );
or ( n37663 , n37548 , n37662 );
or ( n37664 , n37661 , n37547 );
nand ( n37665 , n37663 , n37664 );
not ( n37666 , n37665 );
buf ( n37667 , n33744 );
buf ( n37668 , n34820 );
xor ( n37669 , n37667 , n37668 );
xnor ( n37670 , n37669 , n33230 );
not ( n37671 , n205165 );
not ( n37672 , n204436 );
or ( n37673 , n37671 , n37672 );
not ( n37674 , n204439 );
or ( n37675 , n37674 , n205165 );
nand ( n37676 , n37673 , n37675 );
not ( n37677 , n37676 );
not ( n37678 , n34477 );
and ( n37679 , n37677 , n37678 );
and ( n37680 , n37676 , n34477 );
nor ( n37681 , n37679 , n37680 );
nand ( n37682 , n37670 , n37681 );
not ( n37683 , n37682 );
not ( n37684 , n34890 );
not ( n37685 , n204586 );
or ( n37686 , n37684 , n37685 );
or ( n37687 , n204586 , n34890 );
nand ( n37688 , n37686 , n37687 );
and ( n37689 , n37688 , n204622 );
not ( n37690 , n37688 );
and ( n37691 , n37690 , n204632 );
nor ( n37692 , n37689 , n37691 );
not ( n37693 , n37692 );
not ( n37694 , n37693 );
and ( n37695 , n37683 , n37694 );
nand ( n37696 , n37681 , n37670 );
and ( n37697 , n37696 , n37693 );
nor ( n37698 , n37695 , n37697 );
not ( n37699 , n37698 );
or ( n37700 , n37666 , n37699 );
or ( n37701 , n37698 , n37665 );
nand ( n37702 , n37700 , n37701 );
not ( n37703 , n37702 );
or ( n37704 , n37484 , n37703 );
not ( n37705 , n37483 );
not ( n37706 , n37702 );
nand ( n37707 , n37705 , n37706 );
nand ( n37708 , n37704 , n37707 );
buf ( n37709 , n37708 );
and ( n37710 , n37295 , n37709 );
not ( n37711 , n37295 );
buf ( n37712 , n37702 );
buf ( n37713 , n37483 );
xor ( n37714 , n37712 , n37713 );
buf ( n37715 , n37714 );
and ( n37716 , n37711 , n37715 );
nor ( n37717 , n37710 , n37716 );
not ( n37718 , n37717 );
nand ( n37719 , n35817 , n36734 , n37718 );
not ( n37720 , n35815 );
not ( n37721 , n37720 );
not ( n37722 , n36734 );
or ( n37723 , n37721 , n37722 );
buf ( n37724 , n33252 );
buf ( n37725 , n37724 );
nor ( n37726 , n37718 , n37725 );
nand ( n37727 , n37723 , n37726 );
buf ( n37728 , n35431 );
nand ( n37729 , n37728 , n31919 );
nand ( n37730 , n37719 , n37727 , n37729 );
buf ( n37731 , n37730 );
buf ( n37732 , RI17514990_702);
buf ( n37733 , n37732 );
not ( n37734 , n33096 );
buf ( n37735 , RI19a9ed50_2578);
nand ( n37736 , n25451 , n37735 );
buf ( n37737 , RI174896e8_1066);
and ( n37738 , n37736 , n37737 );
not ( n37739 , n37736 );
not ( n37740 , RI174896e8_1066);
and ( n37741 , n37739 , n37740 );
nor ( n37742 , n37738 , n37741 );
buf ( n37743 , n37742 );
not ( n37744 , n37743 );
not ( n37745 , n37744 );
not ( n37746 , n36070 );
not ( n37747 , n37746 );
or ( n37748 , n37745 , n37747 );
not ( n37749 , n36071 );
nand ( n37750 , n37749 , n37743 );
nand ( n37751 , n37748 , n37750 );
not ( n37752 , n37751 );
or ( n37753 , n37734 , n37752 );
or ( n37754 , n37751 , n33096 );
nand ( n37755 , n37753 , n37754 );
not ( n37756 , n37755 );
not ( n37757 , n204345 );
not ( n37758 , n208165 );
or ( n37759 , n37757 , n37758 );
xor ( n37760 , n30385 , n30402 );
not ( n37761 , n208154 );
xnor ( n37762 , n37760 , n37761 );
nand ( n37763 , n37762 , n204344 );
nand ( n37764 , n37759 , n37763 );
not ( n37765 , n37764 );
not ( n37766 , n33886 );
and ( n37767 , n37765 , n37766 );
and ( n37768 , n37764 , n33886 );
nor ( n37769 , n37767 , n37768 );
buf ( n37770 , RI173bc6f8_1837);
not ( n37771 , n37770 );
not ( n37772 , n29944 );
or ( n37773 , n37771 , n37772 );
xor ( n37774 , n207704 , n26436 );
buf ( n37775 , n29924 );
xnor ( n37776 , n37774 , n37775 );
or ( n37777 , n37770 , n37776 );
nand ( n37778 , n37773 , n37777 );
and ( n37779 , n37778 , n34191 );
not ( n37780 , n37778 );
and ( n37781 , n37780 , n211419 );
nor ( n37782 , n37779 , n37781 );
nand ( n37783 , n37769 , n37782 );
not ( n37784 , n37783 );
or ( n37785 , n37756 , n37784 );
or ( n37786 , n37783 , n37755 );
nand ( n37787 , n37785 , n37786 );
not ( n37788 , n37787 );
not ( n37789 , n204789 );
not ( n37790 , n210940 );
or ( n37791 , n37789 , n37790 );
not ( n37792 , n204789 );
nand ( n37793 , n37792 , n33178 );
nand ( n37794 , n37791 , n37793 );
not ( n37795 , n31036 );
and ( n37796 , n37794 , n37795 );
not ( n37797 , n37794 );
and ( n37798 , n37797 , n33186 );
nor ( n37799 , n37796 , n37798 );
not ( n37800 , n35056 );
not ( n37801 , n204675 );
not ( n37802 , n37801 );
or ( n37803 , n37800 , n37802 );
not ( n37804 , n35056 );
nand ( n37805 , n37804 , n204675 );
nand ( n37806 , n37803 , n37805 );
and ( n37807 , n37806 , n204681 );
not ( n37808 , n37806 );
and ( n37809 , n37808 , n26261 );
nor ( n37810 , n37807 , n37809 );
nand ( n37811 , n37799 , n37810 );
not ( n37812 , n37811 );
buf ( n37813 , RI17487960_1075);
not ( n37814 , n37813 );
not ( n37815 , n35274 );
or ( n37816 , n37814 , n37815 );
or ( n37817 , n35274 , n37813 );
nand ( n215579 , n37816 , n37817 );
not ( n215580 , n34516 );
not ( n37820 , n215580 );
and ( n37821 , n215579 , n37820 );
not ( n37822 , n215579 );
and ( n37823 , n37822 , n215580 );
nor ( n37824 , n37821 , n37823 );
not ( n37825 , n37824 );
not ( n215587 , n37825 );
and ( n215588 , n37812 , n215587 );
and ( n215589 , n37811 , n37825 );
nor ( n215590 , n215588 , n215589 );
not ( n37830 , n215590 );
buf ( n37831 , RI173df4e0_1667);
not ( n37832 , n37831 );
not ( n37833 , RI173967f0_2022);
not ( n37834 , n37833 );
or ( n37835 , n37832 , n37834 );
not ( n37836 , RI173df4e0_1667);
buf ( n37837 , RI173967f0_2022);
nand ( n37838 , n37836 , n37837 );
nand ( n37839 , n37835 , n37838 );
not ( n37840 , RI17456fb8_1312);
and ( n37841 , n37839 , n37840 );
not ( n37842 , n37839 );
buf ( n37843 , RI17456fb8_1312);
and ( n37844 , n37842 , n37843 );
nor ( n37845 , n37841 , n37844 );
buf ( n37846 , RI19a954f8_2645);
nand ( n37847 , n30640 , n37846 );
not ( n37848 , RI1747bb10_1133);
and ( n37849 , n37847 , n37848 );
not ( n37850 , n37847 );
buf ( n37851 , RI1747bb10_1133);
and ( n37852 , n37850 , n37851 );
nor ( n37853 , n37849 , n37852 );
xor ( n37854 , n37845 , n37853 );
buf ( n37855 , RI19ac52e8_2290);
nand ( n37856 , n25711 , n37855 );
not ( n37857 , RI174cb520_778);
and ( n37858 , n37856 , n37857 );
not ( n37859 , n37856 );
buf ( n37860 , RI174cb520_778);
and ( n37861 , n37859 , n37860 );
nor ( n37862 , n37858 , n37861 );
xnor ( n37863 , n37854 , n37862 );
not ( n37864 , n37863 );
not ( n37865 , n37864 );
xor ( n37866 , n33138 , n37865 );
buf ( n37867 , RI174bdc90_820);
not ( n37868 , RI1740ac80_1455);
buf ( n37869 , RI173c1f90_1810);
and ( n37870 , n37868 , n37869 );
not ( n37871 , n37868 );
not ( n37872 , RI173c1f90_1810);
and ( n37873 , n37871 , n37872 );
nor ( n37874 , n37870 , n37873 );
xor ( n37875 , n37867 , n37874 );
buf ( n37876 , RI17338a10_2165);
buf ( n37877 , RI174a72b0_921);
xor ( n37878 , n37876 , n37877 );
buf ( n37879 , RI19ab2b98_2434);
nand ( n37880 , n204513 , n37879 );
xnor ( n37881 , n37878 , n37880 );
xnor ( n37882 , n37875 , n37881 );
xnor ( n37883 , n37866 , n37882 );
not ( n37884 , n37398 );
buf ( n37885 , RI19ac6e18_2278);
nand ( n37886 , n205019 , n37885 );
not ( n37887 , RI174c3e88_801);
and ( n37888 , n37886 , n37887 );
not ( n37889 , n37886 );
buf ( n37890 , RI174c3e88_801);
and ( n37891 , n37889 , n37890 );
nor ( n37892 , n37888 , n37891 );
buf ( n37893 , n37892 );
not ( n37894 , n37893 );
not ( n37895 , n32322 );
or ( n37896 , n37894 , n37895 );
not ( n37897 , n37893 );
xor ( n37898 , n32303 , n32320 );
not ( n37899 , n32311 );
xnor ( n37900 , n37898 , n37899 );
nand ( n37901 , n37897 , n37900 );
nand ( n37902 , n37896 , n37901 );
not ( n37903 , n37902 );
or ( n37904 , n37884 , n37903 );
or ( n37905 , n37902 , n37398 );
nand ( n37906 , n37904 , n37905 );
nand ( n37907 , n37883 , n37906 );
buf ( n37908 , RI173a8220_1936);
not ( n37909 , n37908 );
not ( n37910 , RI173f0f10_1581);
not ( n37911 , n37910 );
or ( n37912 , n37909 , n37911 );
not ( n37913 , RI173a8220_1936);
buf ( n37914 , RI173f0f10_1581);
nand ( n37915 , n37913 , n37914 );
nand ( n37916 , n37912 , n37915 );
not ( n37917 , RI174ae588_886);
and ( n37918 , n37916 , n37917 );
not ( n215680 , n37916 );
buf ( n215681 , RI174ae588_886);
and ( n37921 , n215680 , n215681 );
nor ( n37922 , n37918 , n37921 );
buf ( n37923 , RI19a887a8_2735);
nand ( n37924 , n26276 , n37923 );
buf ( n37925 , RI17517d20_692);
and ( n37926 , n37924 , n37925 );
not ( n37927 , n37924 );
not ( n37928 , RI17517d20_692);
and ( n37929 , n37927 , n37928 );
nor ( n37930 , n37926 , n37929 );
xor ( n37931 , n37922 , n37930 );
buf ( n37932 , RI19ab0000_2454);
nand ( n37933 , n25851 , n37932 );
not ( n37934 , RI1748d1f8_1048);
and ( n37935 , n37933 , n37934 );
not ( n37936 , n37933 );
buf ( n37937 , RI1748d1f8_1048);
and ( n37938 , n37936 , n37937 );
nor ( n37939 , n37935 , n37938 );
xnor ( n37940 , n37931 , n37939 );
not ( n37941 , n37940 );
not ( n37942 , n25436 );
and ( n37943 , n37941 , n37942 );
and ( n37944 , n37940 , n25436 );
nor ( n37945 , n37943 , n37944 );
buf ( n37946 , n31869 );
xor ( n37947 , n37945 , n37946 );
not ( n37948 , n37947 );
and ( n37949 , n37907 , n37948 );
not ( n37950 , n37907 );
and ( n37951 , n37950 , n37947 );
nor ( n37952 , n37949 , n37951 );
not ( n37953 , n37952 );
or ( n37954 , n37830 , n37953 );
or ( n37955 , n37952 , n215590 );
nand ( n37956 , n37954 , n37955 );
not ( n37957 , n37755 );
not ( n37958 , n37769 );
nand ( n37959 , n37957 , n37958 );
not ( n37960 , n37959 );
buf ( n37961 , RI17457300_1311);
not ( n37962 , n37961 );
not ( n37963 , n34137 );
buf ( n37964 , RI19a8b4a8_2716);
nand ( n37965 , n29435 , n37964 );
not ( n37966 , RI1746d560_1203);
and ( n37967 , n37965 , n37966 );
not ( n37968 , n37965 );
buf ( n37969 , RI1746d560_1203);
and ( n37970 , n37968 , n37969 );
nor ( n37971 , n37967 , n37970 );
not ( n37972 , n37971 );
or ( n37973 , n37963 , n37972 );
or ( n37974 , n34137 , n37971 );
nand ( n37975 , n37973 , n37974 );
buf ( n37976 , RI173d1278_1736);
not ( n37977 , n37976 );
not ( n37978 , RI17358cc0_2092);
not ( n37979 , n37978 );
or ( n37980 , n37977 , n37979 );
not ( n37981 , RI173d1278_1736);
buf ( n37982 , RI17358cc0_2092);
nand ( n37983 , n37981 , n37982 );
nand ( n37984 , n37980 , n37983 );
buf ( n37985 , RI17448d50_1381);
and ( n37986 , n37984 , n37985 );
not ( n37987 , n37984 );
not ( n37988 , RI17448d50_1381);
and ( n37989 , n37987 , n37988 );
nor ( n37990 , n37986 , n37989 );
xnor ( n37991 , n37975 , n37990 );
not ( n37992 , n37991 );
or ( n37993 , n37962 , n37992 );
xor ( n37994 , n37990 , n34137 );
buf ( n37995 , n37971 );
xnor ( n37996 , n37994 , n37995 );
not ( n37997 , RI17457300_1311);
nand ( n37998 , n37996 , n37997 );
nand ( n37999 , n37993 , n37998 );
buf ( n38000 , n35481 );
not ( n38001 , n38000 );
and ( n38002 , n37999 , n38001 );
not ( n38003 , n37999 );
and ( n38004 , n38003 , n38000 );
nor ( n38005 , n38002 , n38004 );
not ( n38006 , n38005 );
and ( n38007 , n37960 , n38006 );
and ( n38008 , n37959 , n38005 );
nor ( n38009 , n38007 , n38008 );
not ( n38010 , n38009 );
and ( n38011 , n37956 , n38010 );
not ( n38012 , n37956 );
and ( n38013 , n38012 , n38009 );
nor ( n38014 , n38011 , n38013 );
not ( n38015 , n38014 );
not ( n38016 , n205193 );
not ( n38017 , n30220 );
or ( n38018 , n38016 , n38017 );
nand ( n38019 , n204391 , n205190 );
nand ( n38020 , n38018 , n38019 );
and ( n38021 , n38020 , n31778 );
not ( n38022 , n38020 );
and ( n38023 , n38022 , n33685 );
nor ( n38024 , n38021 , n38023 );
not ( n38025 , n38024 );
not ( n38026 , n38025 );
buf ( n38027 , RI19abef88_2341);
nand ( n38028 , n25491 , n38027 );
buf ( n38029 , RI174af5f0_881);
and ( n38030 , n38028 , n38029 );
not ( n38031 , n38028 );
not ( n38032 , RI174af5f0_881);
and ( n38033 , n38031 , n38032 );
nor ( n38034 , n38030 , n38033 );
buf ( n38035 , n38034 );
xor ( n38036 , n38035 , n28722 );
buf ( n38037 , n32524 );
xnor ( n38038 , n38036 , n38037 );
not ( n38039 , n32076 );
not ( n38040 , n38039 );
not ( n215802 , n36685 );
or ( n215803 , n38040 , n215802 );
or ( n38043 , n36685 , n38039 );
nand ( n38044 , n215803 , n38043 );
and ( n38045 , n38044 , n36238 );
not ( n38046 , n38044 );
and ( n38047 , n38046 , n36243 );
nor ( n38048 , n38045 , n38047 );
nand ( n38049 , n38038 , n38048 );
not ( n38050 , n38049 );
or ( n38051 , n38026 , n38050 );
or ( n38052 , n38049 , n38025 );
nand ( n38053 , n38051 , n38052 );
not ( n38054 , n38053 );
buf ( n38055 , RI1740ee20_1435);
buf ( n38056 , RI173d50d0_1717);
not ( n38057 , n38056 );
not ( n38058 , RI1738c3e0_2072);
not ( n38059 , n38058 );
or ( n38060 , n38057 , n38059 );
not ( n38061 , RI173d50d0_1717);
buf ( n38062 , RI1738c3e0_2072);
nand ( n38063 , n38061 , n38062 );
nand ( n38064 , n38060 , n38063 );
not ( n38065 , RI1744cba8_1362);
and ( n38066 , n38064 , n38065 );
not ( n38067 , n38064 );
buf ( n38068 , RI1744cba8_1362);
and ( n38069 , n38067 , n38068 );
nor ( n38070 , n38066 , n38069 );
buf ( n38071 , RI19acc020_2239);
nand ( n38072 , n205019 , n38071 );
buf ( n38073 , RI174bae28_829);
and ( n38074 , n38072 , n38073 );
not ( n38075 , n38072 );
not ( n38076 , RI174bae28_829);
and ( n38077 , n38075 , n38076 );
nor ( n38078 , n38074 , n38077 );
xor ( n38079 , n38070 , n38078 );
buf ( n38080 , RI19a9d1a8_2590);
nand ( n38081 , n29203 , n38080 );
not ( n38082 , RI174713b8_1184);
and ( n38083 , n38081 , n38082 );
not ( n38084 , n38081 );
buf ( n38085 , RI174713b8_1184);
and ( n38086 , n38084 , n38085 );
nor ( n38087 , n38083 , n38086 );
xnor ( n38088 , n38079 , n38087 );
buf ( n38089 , n38088 );
not ( n38090 , n38089 );
xor ( n38091 , n38055 , n38090 );
xnor ( n38092 , n38091 , n37510 );
not ( n38093 , n38092 );
not ( n38094 , n38093 );
buf ( n38095 , n37853 );
not ( n38096 , n38095 );
buf ( n38097 , RI173d0f18_1737);
not ( n38098 , n38097 );
not ( n38099 , RI17347650_2093);
not ( n38100 , n38099 );
or ( n38101 , n38098 , n38100 );
not ( n38102 , RI173d0f18_1737);
buf ( n38103 , RI17347650_2093);
nand ( n38104 , n38102 , n38103 );
nand ( n38105 , n38101 , n38104 );
not ( n38106 , RI17448a08_1382);
and ( n38107 , n38105 , n38106 );
not ( n38108 , n38105 );
buf ( n38109 , RI17448a08_1382);
and ( n38110 , n38108 , n38109 );
nor ( n38111 , n38107 , n38110 );
buf ( n38112 , RI19abca80_2362);
nand ( n38113 , n25451 , n38112 );
buf ( n38114 , RI174b5ef0_849);
and ( n38115 , n38113 , n38114 );
not ( n38116 , n38113 );
not ( n38117 , RI174b5ef0_849);
and ( n38118 , n38116 , n38117 );
nor ( n38119 , n38115 , n38118 );
xor ( n38120 , n38111 , n38119 );
buf ( n38121 , RI19a8b250_2717);
nand ( n38122 , n25622 , n38121 );
not ( n38123 , RI1746d218_1204);
and ( n38124 , n38122 , n38123 );
not ( n38125 , n38122 );
buf ( n38126 , RI1746d218_1204);
and ( n38127 , n38125 , n38126 );
nor ( n38128 , n38124 , n38127 );
xor ( n38129 , n38120 , n38128 );
not ( n38130 , n38129 );
not ( n38131 , n38130 );
or ( n38132 , n38096 , n38131 );
not ( n38133 , n38095 );
nand ( n38134 , n38133 , n38129 );
nand ( n38135 , n38132 , n38134 );
not ( n38136 , n25675 );
buf ( n38137 , n38136 );
and ( n38138 , n38135 , n38137 );
not ( n38139 , n38135 );
not ( n38140 , n38136 );
buf ( n38141 , n38140 );
and ( n38142 , n38139 , n38141 );
nor ( n38143 , n38138 , n38142 );
buf ( n38144 , RI19acc5c0_2236);
nand ( n38145 , n204426 , n38144 );
not ( n38146 , RI17514eb8_701);
and ( n38147 , n38145 , n38146 );
not ( n38148 , n38145 );
buf ( n38149 , RI17514eb8_701);
and ( n38150 , n38148 , n38149 );
nor ( n38151 , n38147 , n38150 );
buf ( n38152 , n38151 );
not ( n38153 , n38152 );
buf ( n38154 , RI173e0890_1661);
not ( n38155 , n38154 );
not ( n38156 , RI17397ba0_2016);
not ( n38157 , n38156 );
or ( n38158 , n38155 , n38157 );
not ( n38159 , RI173e0890_1661);
buf ( n38160 , RI17397ba0_2016);
nand ( n38161 , n38159 , n38160 );
nand ( n38162 , n38158 , n38161 );
not ( n38163 , RI174586b0_1305);
and ( n38164 , n38162 , n38163 );
not ( n38165 , n38162 );
buf ( n38166 , RI174586b0_1305);
and ( n38167 , n38165 , n38166 );
nor ( n38168 , n38164 , n38167 );
buf ( n38169 , RI19ac3920_2302);
nand ( n38170 , n204512 , n38169 );
buf ( n38171 , RI174cd410_772);
and ( n38172 , n38170 , n38171 );
not ( n38173 , n38170 );
not ( n38174 , RI174cd410_772);
and ( n38175 , n38173 , n38174 );
nor ( n38176 , n38172 , n38175 );
buf ( n38177 , n38176 );
xor ( n38178 , n38168 , n38177 );
buf ( n38179 , RI19a936f8_2658);
nand ( n38180 , n26266 , n38179 );
not ( n38181 , RI1747cec0_1127);
and ( n38182 , n38180 , n38181 );
not ( n38183 , n38180 );
buf ( n38184 , RI1747cec0_1127);
and ( n38185 , n38183 , n38184 );
nor ( n38186 , n38182 , n38185 );
buf ( n38187 , n38186 );
xnor ( n38188 , n38178 , n38187 );
not ( n38189 , n38188 );
or ( n38190 , n38153 , n38189 );
not ( n38191 , n38152 );
not ( n38192 , n38176 );
not ( n215954 , n38186 );
or ( n215955 , n38192 , n215954 );
or ( n38195 , n38176 , n38186 );
nand ( n38196 , n215955 , n38195 );
not ( n38197 , n38168 );
and ( n38198 , n38196 , n38197 );
not ( n38199 , n38196 );
and ( n38200 , n38199 , n38168 );
nor ( n38201 , n38198 , n38200 );
nand ( n38202 , n38191 , n38201 );
nand ( n38203 , n38190 , n38202 );
not ( n38204 , n29409 );
not ( n38205 , n38204 );
and ( n38206 , n38203 , n38205 );
not ( n38207 , n38203 );
and ( n38208 , n38207 , n29411 );
nor ( n38209 , n38206 , n38208 );
nor ( n38210 , n38143 , n38209 );
not ( n38211 , n38210 );
and ( n38212 , n38094 , n38211 );
and ( n38213 , n38093 , n38210 );
nor ( n38214 , n38212 , n38213 );
not ( n38215 , n38214 );
and ( n38216 , n38054 , n38215 );
and ( n38217 , n38053 , n38214 );
nor ( n38218 , n38216 , n38217 );
not ( n38219 , n38218 );
and ( n38220 , n38015 , n38219 );
and ( n38221 , n38014 , n38218 );
nor ( n38222 , n38220 , n38221 );
not ( n38223 , n38222 );
or ( n38224 , n37788 , n38223 );
not ( n38225 , n37787 );
not ( n38226 , n38218 );
not ( n38227 , n38014 );
or ( n38228 , n38226 , n38227 );
not ( n38229 , n38014 );
not ( n38230 , n38218 );
nand ( n38231 , n38229 , n38230 );
nand ( n38232 , n38228 , n38231 );
nand ( n38233 , n38225 , n38232 );
nand ( n38234 , n38224 , n38233 );
not ( n38235 , n37626 );
not ( n38236 , n29693 );
or ( n38237 , n38235 , n38236 );
not ( n38238 , n37626 );
nand ( n38239 , n38238 , n31135 );
nand ( n38240 , n38237 , n38239 );
and ( n38241 , n38240 , n29733 );
not ( n38242 , n38240 );
and ( n38243 , n38242 , n207493 );
nor ( n38244 , n38241 , n38243 );
not ( n38245 , n33491 );
not ( n38246 , n28555 );
or ( n38247 , n38245 , n38246 );
not ( n38248 , n33491 );
xor ( n38249 , n206297 , n28544 );
xnor ( n38250 , n38249 , n28554 );
nand ( n38251 , n38248 , n38250 );
nand ( n38252 , n38247 , n38251 );
xor ( n38253 , n35338 , n35355 );
not ( n38254 , n35346 );
xor ( n38255 , n38253 , n38254 );
not ( n38256 , n38255 );
not ( n38257 , n38256 );
and ( n38258 , n38252 , n38257 );
not ( n38259 , n38252 );
and ( n38260 , n38259 , n35358 );
nor ( n38261 , n38258 , n38260 );
nand ( n38262 , n38244 , n38261 );
not ( n38263 , n38262 );
not ( n38264 , n204936 );
buf ( n38265 , RI17530f50_614);
not ( n38266 , n38265 );
buf ( n38267 , RI173f2950_1573);
not ( n38268 , n38267 );
not ( n38269 , RI173a9c60_1928);
not ( n38270 , n38269 );
or ( n38271 , n38268 , n38270 );
not ( n38272 , RI173f2950_1573);
buf ( n38273 , RI173a9c60_1928);
nand ( n38274 , n38272 , n38273 );
nand ( n38275 , n38271 , n38274 );
not ( n38276 , RI174c1a70_808);
and ( n38277 , n38275 , n38276 );
not ( n38278 , n38275 );
buf ( n38279 , RI174c1a70_808);
and ( n38280 , n38278 , n38279 );
nor ( n38281 , n38277 , n38280 );
buf ( n38282 , RI19aae980_2464);
nand ( n38283 , n25539 , n38282 );
buf ( n38284 , RI1748ef80_1039);
and ( n38285 , n38283 , n38284 );
not ( n38286 , n38283 );
not ( n38287 , RI1748ef80_1039);
and ( n216049 , n38286 , n38287 );
nor ( n216050 , n38285 , n216049 );
xor ( n38290 , n38281 , n216050 );
xnor ( n216052 , n38290 , n33995 );
not ( n216053 , n216052 );
or ( n38293 , n38266 , n216053 );
or ( n38294 , n216052 , n38265 );
nand ( n38295 , n38293 , n38294 );
not ( n38296 , n38295 );
or ( n38297 , n38264 , n38296 );
or ( n38298 , n38295 , n204936 );
nand ( n38299 , n38297 , n38298 );
not ( n38300 , n38299 );
and ( n38301 , n38263 , n38300 );
and ( n38302 , n38262 , n38299 );
nor ( n38303 , n38301 , n38302 );
not ( n38304 , n38303 );
not ( n38305 , n28404 );
buf ( n38306 , RI173f2c98_1572);
not ( n38307 , n38306 );
not ( n38308 , n26308 );
or ( n38309 , n38307 , n38308 );
not ( n38310 , n38306 );
nand ( n38311 , n38310 , n26317 );
nand ( n38312 , n38309 , n38311 );
xor ( n38313 , n38305 , n38312 );
not ( n38314 , n36129 );
buf ( n38315 , RI19a97028_2633);
nand ( n38316 , n25656 , n38315 );
buf ( n38317 , RI17476c50_1157);
and ( n38318 , n38316 , n38317 );
not ( n38319 , n38316 );
not ( n38320 , RI17476c50_1157);
and ( n38321 , n38319 , n38320 );
nor ( n38322 , n38318 , n38321 );
not ( n38323 , n38322 );
not ( n38324 , n37892 );
or ( n38325 , n38323 , n38324 );
or ( n38326 , n38322 , n37892 );
nand ( n38327 , n38325 , n38326 );
buf ( n38328 , RI173da968_1690);
not ( n38329 , n38328 );
not ( n38330 , RI17391c78_2045);
not ( n38331 , n38330 );
or ( n38332 , n38329 , n38331 );
not ( n38333 , RI173da968_1690);
buf ( n38334 , RI17391c78_2045);
nand ( n38335 , n38333 , n38334 );
nand ( n38336 , n38332 , n38335 );
not ( n38337 , RI17452440_1335);
and ( n38338 , n38336 , n38337 );
not ( n38339 , n38336 );
buf ( n38340 , RI17452440_1335);
and ( n38341 , n38339 , n38340 );
nor ( n38342 , n38338 , n38341 );
and ( n38343 , n38327 , n38342 );
not ( n38344 , n38327 );
not ( n38345 , n38342 );
and ( n38346 , n38344 , n38345 );
nor ( n38347 , n38343 , n38346 );
not ( n38348 , n38347 );
or ( n38349 , n38314 , n38348 );
or ( n38350 , n38347 , n36129 );
nand ( n38351 , n38349 , n38350 );
not ( n38352 , n38351 );
not ( n38353 , n28597 );
not ( n38354 , n38353 );
and ( n38355 , n38352 , n38354 );
buf ( n38356 , n28594 );
and ( n38357 , n38351 , n38356 );
nor ( n38358 , n38355 , n38357 );
nand ( n38359 , n38313 , n38358 );
buf ( n38360 , RI19ac6ff8_2277);
nand ( n38361 , n25416 , n38360 );
not ( n38362 , RI174c43b0_800);
and ( n38363 , n38361 , n38362 );
not ( n38364 , n38361 );
buf ( n38365 , RI174c43b0_800);
and ( n38366 , n38364 , n38365 );
nor ( n38367 , n38363 , n38366 );
not ( n38368 , n38367 );
not ( n38369 , n32406 );
or ( n38370 , n38368 , n38369 );
not ( n38371 , n38367 );
not ( n38372 , n32402 );
nand ( n38373 , n38371 , n38372 );
nand ( n38374 , n38370 , n38373 );
and ( n38375 , n38374 , n32443 );
not ( n216137 , n38374 );
and ( n216138 , n216137 , n32442 );
nor ( n38378 , n38375 , n216138 );
xor ( n38379 , n38359 , n38378 );
not ( n38380 , n38379 );
or ( n38381 , n38304 , n38380 );
or ( n38382 , n38379 , n38303 );
nand ( n38383 , n38381 , n38382 );
not ( n38384 , n38383 );
not ( n38385 , n38384 );
not ( n38386 , n29860 );
not ( n38387 , n38386 );
not ( n38388 , n36534 );
not ( n38389 , n38388 );
not ( n38390 , n26486 );
and ( n38391 , n38389 , n38390 );
and ( n38392 , n29815 , n26486 );
nor ( n38393 , n38391 , n38392 );
not ( n38394 , n38393 );
or ( n38395 , n38387 , n38394 );
buf ( n38396 , n29854 );
not ( n38397 , n38396 );
or ( n38398 , n38393 , n38397 );
nand ( n38399 , n38395 , n38398 );
buf ( n38400 , n38399 );
not ( n38401 , n38400 );
buf ( n38402 , RI173da620_1691);
not ( n38403 , n38402 );
not ( n38404 , RI17391930_2046);
not ( n38405 , n38404 );
or ( n38406 , n38403 , n38405 );
not ( n38407 , RI173da620_1691);
buf ( n38408 , RI17391930_2046);
nand ( n38409 , n38407 , n38408 );
nand ( n38410 , n38406 , n38409 );
buf ( n38411 , RI174520f8_1336);
and ( n38412 , n38410 , n38411 );
not ( n38413 , n38410 );
not ( n38414 , RI174520f8_1336);
and ( n38415 , n38413 , n38414 );
nor ( n38416 , n38412 , n38415 );
buf ( n38417 , RI19ac8e70_2263);
nand ( n38418 , n205124 , n38417 );
buf ( n38419 , RI174c3960_802);
and ( n38420 , n38418 , n38419 );
not ( n38421 , n38418 );
not ( n38422 , RI174c3960_802);
and ( n38423 , n38421 , n38422 );
nor ( n38424 , n38420 , n38423 );
xor ( n38425 , n38416 , n38424 );
buf ( n38426 , RI19a99440_2617);
nand ( n38427 , n204426 , n38426 );
buf ( n38428 , RI17476908_1158);
and ( n38429 , n38427 , n38428 );
not ( n38430 , n38427 );
not ( n38431 , RI17476908_1158);
and ( n38432 , n38430 , n38431 );
nor ( n38433 , n38429 , n38432 );
xnor ( n38434 , n38425 , n38433 );
buf ( n38435 , n38434 );
buf ( n38436 , n38435 );
xor ( n38437 , n29486 , n38436 );
buf ( n38438 , RI17405dc0_1479);
not ( n38439 , n38438 );
not ( n38440 , RI173bd0d0_1834);
not ( n38441 , n38440 );
or ( n38442 , n38439 , n38441 );
not ( n38443 , RI17405dc0_1479);
buf ( n38444 , RI173bd0d0_1834);
nand ( n38445 , n38443 , n38444 );
nand ( n38446 , n38442 , n38445 );
not ( n38447 , n38446 );
not ( n38448 , n38447 );
buf ( n38449 , RI17333b50_2189);
not ( n38450 , RI17408ef8_1464);
xor ( n38451 , n38449 , n38450 );
buf ( n216213 , RI19ab6900_2405);
nand ( n216214 , n25583 , n216213 );
not ( n38454 , RI174a20a8_946);
and ( n216216 , n216214 , n38454 );
not ( n216217 , n216214 );
buf ( n38457 , RI174a20a8_946);
and ( n38458 , n216217 , n38457 );
nor ( n38459 , n216216 , n38458 );
xnor ( n38460 , n38451 , n38459 );
not ( n38461 , n38460 );
or ( n38462 , n38448 , n38461 );
or ( n216224 , n38460 , n38447 );
nand ( n216225 , n38462 , n216224 );
xnor ( n216226 , n38437 , n216225 );
nand ( n216227 , n38401 , n216226 );
not ( n38467 , n216227 );
not ( n38468 , n33685 );
not ( n38469 , n204390 );
buf ( n38470 , n205203 );
not ( n38471 , n38470 );
and ( n38472 , n38469 , n38471 );
and ( n38473 , n204390 , n38470 );
nor ( n38474 , n38472 , n38473 );
not ( n38475 , n38474 );
and ( n38476 , n38468 , n38475 );
and ( n38477 , n33685 , n38474 );
nor ( n38478 , n38476 , n38477 );
not ( n38479 , n38478 );
not ( n38480 , n38479 );
and ( n38481 , n38467 , n38480 );
not ( n38482 , n38400 );
nand ( n38483 , n38482 , n216226 );
and ( n38484 , n38483 , n38479 );
nor ( n38485 , n38481 , n38484 );
not ( n38486 , n38485 );
not ( n38487 , n38486 );
or ( n38488 , n38385 , n38487 );
nand ( n38489 , n38485 , n38383 );
nand ( n38490 , n38488 , n38489 );
not ( n38491 , n29361 );
not ( n38492 , n31515 );
or ( n38493 , n38491 , n38492 );
nand ( n38494 , n31528 , n207118 );
nand ( n38495 , n38493 , n38494 );
and ( n38496 , n38495 , n33853 );
not ( n38497 , n38495 );
not ( n38498 , n33853 );
and ( n38499 , n38497 , n38498 );
nor ( n216261 , n38496 , n38499 );
not ( n216262 , n32049 );
nand ( n38502 , n216262 , n205001 );
not ( n38503 , n38502 );
nor ( n38504 , n32053 , n205001 );
nor ( n38505 , n38503 , n38504 );
not ( n38506 , n38505 );
not ( n38507 , n32082 );
or ( n38508 , n38506 , n38507 );
or ( n38509 , n32082 , n38505 );
nand ( n38510 , n38508 , n38509 );
not ( n38511 , n38510 );
nand ( n38512 , n216261 , n38511 );
not ( n38513 , n38512 );
xor ( n38514 , n37045 , n37069 );
not ( n38515 , n38514 );
buf ( n38516 , RI19acc818_2235);
nand ( n38517 , n25741 , n38516 );
buf ( n38518 , RI175153e0_700);
and ( n38519 , n38517 , n38518 );
not ( n38520 , n38517 );
not ( n38521 , RI175153e0_700);
and ( n38522 , n38520 , n38521 );
nor ( n38523 , n38519 , n38522 );
buf ( n38524 , n38523 );
not ( n38525 , n38524 );
buf ( n38526 , RI17397ee8_2015);
not ( n38527 , n38526 );
not ( n38528 , RI173e0bd8_1660);
not ( n38529 , n38528 );
or ( n38530 , n38527 , n38529 );
not ( n38531 , RI17397ee8_2015);
buf ( n38532 , RI173e0bd8_1660);
nand ( n38533 , n38531 , n38532 );
nand ( n38534 , n38530 , n38533 );
not ( n38535 , RI174589f8_1304);
and ( n38536 , n38534 , n38535 );
not ( n38537 , n38534 );
buf ( n38538 , RI174589f8_1304);
and ( n38539 , n38537 , n38538 );
nor ( n38540 , n38536 , n38539 );
buf ( n38541 , RI19ac3b00_2301);
nand ( n38542 , n25751 , n38541 );
buf ( n38543 , RI174cd938_771);
and ( n38544 , n38542 , n38543 );
not ( n38545 , n38542 );
not ( n38546 , RI174cd938_771);
and ( n38547 , n38545 , n38546 );
nor ( n38548 , n38544 , n38547 );
xor ( n38549 , n38540 , n38548 );
buf ( n38550 , RI19a93950_2657);
nand ( n38551 , n25451 , n38550 );
buf ( n38552 , RI1747d208_1126);
and ( n38553 , n38551 , n38552 );
not ( n38554 , n38551 );
not ( n38555 , RI1747d208_1126);
and ( n38556 , n38554 , n38555 );
nor ( n38557 , n38553 , n38556 );
xnor ( n38558 , n38549 , n38557 );
not ( n38559 , n38558 );
or ( n38560 , n38525 , n38559 );
or ( n38561 , n38558 , n38524 );
nand ( n38562 , n38560 , n38561 );
not ( n38563 , n38562 );
and ( n38564 , n38515 , n38563 );
not ( n38565 , n37044 );
not ( n38566 , n37070 );
or ( n38567 , n38565 , n38566 );
nand ( n38568 , n37069 , n37045 );
nand ( n38569 , n38567 , n38568 );
not ( n38570 , n38569 );
and ( n38571 , n38570 , n38562 );
nor ( n38572 , n38564 , n38571 );
not ( n38573 , n38572 );
not ( n38574 , n38573 );
and ( n38575 , n38513 , n38574 );
and ( n38576 , n38512 , n38573 );
nor ( n38577 , n38575 , n38576 );
not ( n38578 , n38577 );
not ( n38579 , n38578 );
buf ( n38580 , n32951 );
buf ( n38581 , n29909 );
xor ( n38582 , n38580 , n38581 );
not ( n38583 , RI173fda80_1519);
xor ( n38584 , n38583 , n25992 );
xnor ( n38585 , n38584 , n26007 );
buf ( n38586 , n38585 );
buf ( n38587 , n38586 );
xnor ( n38588 , n38582 , n38587 );
not ( n38589 , n38588 );
not ( n38590 , n29022 );
not ( n38591 , n28043 );
or ( n38592 , n38590 , n38591 );
or ( n38593 , n28043 , n29022 );
nand ( n38594 , n38592 , n38593 );
and ( n38595 , n38594 , n36572 );
not ( n38596 , n38594 );
and ( n38597 , n38596 , n36573 );
nor ( n216359 , n38595 , n38597 );
not ( n216360 , n31875 );
not ( n38600 , n205383 );
or ( n38601 , n216360 , n38600 );
not ( n38602 , n205384 );
or ( n38603 , n38602 , n31875 );
nand ( n38604 , n38601 , n38603 );
not ( n38605 , n38604 );
not ( n38606 , n30757 );
and ( n38607 , n38605 , n38606 );
and ( n38608 , n38604 , n30757 );
nor ( n38609 , n38607 , n38608 );
not ( n38610 , n38609 );
nand ( n38611 , n216359 , n38610 );
not ( n38612 , n38611 );
or ( n38613 , n38589 , n38612 );
or ( n38614 , n38611 , n38588 );
nand ( n38615 , n38613 , n38614 );
not ( n38616 , n38615 );
not ( n38617 , n38616 );
or ( n38618 , n38579 , n38617 );
nand ( n38619 , n38615 , n38577 );
nand ( n38620 , n38618 , n38619 );
and ( n38621 , n38490 , n38620 );
not ( n38622 , n38490 );
not ( n38623 , n38620 );
and ( n38624 , n38622 , n38623 );
nor ( n38625 , n38621 , n38624 );
not ( n38626 , n38625 );
not ( n38627 , n38626 );
and ( n38628 , n38234 , n38627 );
not ( n38629 , n38234 );
and ( n38630 , n38490 , n38623 );
not ( n38631 , n38490 );
and ( n38632 , n38631 , n38620 );
nor ( n38633 , n38630 , n38632 );
buf ( n38634 , n38633 );
and ( n38635 , n38629 , n38634 );
nor ( n38636 , n38628 , n38635 );
buf ( n38637 , n35427 );
not ( n38638 , n38637 );
nand ( n38639 , n38636 , n38638 );
buf ( n38640 , RI17410860_1427);
not ( n38641 , n38640 );
not ( n38642 , RI17401f68_1498);
buf ( n38643 , RI173b9278_1853);
nand ( n38644 , n38642 , n38643 );
not ( n38645 , RI173b9278_1853);
buf ( n38646 , RI17401f68_1498);
nand ( n38647 , n38645 , n38646 );
and ( n38648 , n38644 , n38647 );
xor ( n38649 , n31351 , n38648 );
buf ( n38650 , RI175323f0_610);
not ( n38651 , RI1749e250_965);
xor ( n216413 , n38650 , n38651 );
buf ( n216414 , RI19ab8f70_2388);
nand ( n38654 , n26059 , n216414 );
xnor ( n216416 , n216413 , n38654 );
xnor ( n216417 , n38649 , n216416 );
buf ( n38657 , n216417 );
not ( n38658 , n38657 );
or ( n38659 , n38641 , n38658 );
or ( n38660 , n38657 , n38640 );
nand ( n38661 , n38659 , n38660 );
buf ( n38662 , n31213 );
and ( n38663 , n38661 , n38662 );
not ( n38664 , n38661 );
not ( n38665 , n31188 );
and ( n38666 , n31212 , n31179 );
not ( n38667 , n31212 );
not ( n38668 , RI1744e2a0_1355);
and ( n38669 , n38667 , n38668 );
nor ( n38670 , n38666 , n38669 );
not ( n38671 , n38670 );
not ( n38672 , n38671 );
or ( n38673 , n38665 , n38672 );
not ( n38674 , n31188 );
nand ( n38675 , n38670 , n38674 );
nand ( n38676 , n38673 , n38675 );
buf ( n38677 , n38676 );
and ( n38678 , n38664 , n38677 );
nor ( n38679 , n38663 , n38678 );
buf ( n38680 , n31471 );
not ( n38681 , n38680 );
not ( n38682 , n207214 );
not ( n38683 , n38682 );
or ( n38684 , n38681 , n38683 );
or ( n38685 , n38682 , n38680 );
nand ( n38686 , n38684 , n38685 );
xor ( n38687 , n37160 , n25822 );
not ( n38688 , n37169 );
xnor ( n38689 , n38687 , n38688 );
not ( n38690 , n38689 );
not ( n38691 , n38690 );
and ( n38692 , n38686 , n38691 );
not ( n38693 , n38686 );
not ( n38694 , n38691 );
and ( n38695 , n38693 , n38694 );
nor ( n38696 , n38692 , n38695 );
nand ( n38697 , n38679 , n38696 );
not ( n38698 , n205339 );
not ( n38699 , n31832 );
not ( n38700 , n38699 );
or ( n38701 , n38698 , n38700 );
nand ( n38702 , n31832 , n205335 );
nand ( n38703 , n38701 , n38702 );
buf ( n38704 , n31673 );
not ( n38705 , n38704 );
and ( n38706 , n38703 , n38705 );
not ( n38707 , n38703 );
buf ( n38708 , n31672 );
not ( n38709 , n38708 );
and ( n38710 , n38707 , n38709 );
nor ( n38711 , n38706 , n38710 );
not ( n38712 , n38711 );
and ( n38713 , n38697 , n38712 );
not ( n38714 , n38697 );
and ( n38715 , n38714 , n38711 );
nor ( n38716 , n38713 , n38715 );
not ( n38717 , n38716 );
and ( n38718 , n204758 , n33182 );
not ( n38719 , n204758 );
not ( n38720 , n33182 );
and ( n38721 , n38719 , n38720 );
nor ( n38722 , n38718 , n38721 );
and ( n38723 , n38722 , n33186 );
not ( n38724 , n38722 );
and ( n38725 , n38724 , n37795 );
nor ( n38726 , n38723 , n38725 );
not ( n38727 , n216052 );
buf ( n38728 , RI173d9270_1697);
not ( n216490 , n38728 );
and ( n216491 , n38727 , n216490 );
xor ( n38731 , n38281 , n216050 );
xnor ( n216493 , n38731 , n33995 );
and ( n216494 , n216493 , n38728 );
nor ( n38734 , n216491 , n216494 );
and ( n216496 , n38734 , n204936 );
not ( n216497 , n38734 );
and ( n38737 , n216497 , n204939 );
nor ( n38738 , n216496 , n38737 );
nand ( n38739 , n38726 , n38738 );
not ( n38740 , n38739 );
buf ( n38741 , RI173a1c68_1967);
not ( n38742 , n38741 );
not ( n38743 , n28646 );
or ( n38744 , n38742 , n38743 );
not ( n38745 , n28627 );
xor ( n38746 , n38745 , n28635 );
xnor ( n38747 , n38746 , n28645 );
not ( n38748 , RI173a1c68_1967);
nand ( n38749 , n38747 , n38748 );
nand ( n38750 , n38744 , n38749 );
not ( n38751 , n38750 );
not ( n38752 , n32457 );
and ( n38753 , n38751 , n38752 );
and ( n38754 , n38750 , n32457 );
nor ( n38755 , n38753 , n38754 );
not ( n38756 , n38755 );
not ( n38757 , n38756 );
and ( n38758 , n38740 , n38757 );
and ( n38759 , n38739 , n38756 );
nor ( n38760 , n38758 , n38759 );
not ( n38761 , n30547 );
xor ( n38762 , n27783 , n27791 );
xor ( n38763 , n38762 , n205561 );
not ( n38764 , n38763 );
not ( n38765 , n38764 );
or ( n38766 , n38761 , n38765 );
not ( n38767 , n30547 );
nand ( n38768 , n38767 , n38763 );
nand ( n38769 , n38766 , n38768 );
buf ( n38770 , n29007 );
not ( n38771 , n38770 );
and ( n38772 , n38769 , n38771 );
not ( n38773 , n38769 );
buf ( n38774 , n29006 );
not ( n38775 , n38774 );
and ( n38776 , n38773 , n38775 );
nor ( n38777 , n38772 , n38776 );
not ( n38778 , n38777 );
not ( n38779 , n211807 );
not ( n38780 , n204828 );
xor ( n38781 , n206618 , n28874 );
not ( n38782 , n28865 );
xor ( n38783 , n38781 , n38782 );
not ( n38784 , n38783 );
or ( n38785 , n38780 , n38784 );
or ( n38786 , n38783 , n204828 );
nand ( n38787 , n38785 , n38786 );
not ( n38788 , n38787 );
or ( n38789 , n38779 , n38788 );
or ( n38790 , n38787 , n211807 );
nand ( n38791 , n38789 , n38790 );
buf ( n38792 , n38791 );
nand ( n38793 , n38778 , n38792 );
not ( n38794 , n33822 );
not ( n38795 , n37192 );
not ( n38796 , n38795 );
or ( n38797 , n38794 , n38796 );
not ( n38798 , n33822 );
nand ( n38799 , n38798 , n37192 );
nand ( n38800 , n38797 , n38799 );
buf ( n38801 , n29046 );
not ( n38802 , n38801 );
and ( n38803 , n38800 , n38802 );
not ( n38804 , n38800 );
not ( n38805 , n29046 );
buf ( n38806 , n38805 );
not ( n38807 , n38806 );
and ( n38808 , n38804 , n38807 );
nor ( n38809 , n38803 , n38808 );
not ( n38810 , n38809 );
and ( n38811 , n38793 , n38810 );
not ( n38812 , n38793 );
and ( n38813 , n38812 , n38809 );
nor ( n38814 , n38811 , n38813 );
xor ( n38815 , n38760 , n38814 );
not ( n38816 , n36593 );
not ( n38817 , n35389 );
not ( n38818 , n38817 );
or ( n38819 , n38816 , n38818 );
not ( n38820 , n36593 );
buf ( n38821 , RI174458d0_1397);
xor ( n38822 , n38821 , n35373 );
xnor ( n38823 , n38822 , n35388 );
nand ( n216585 , n38820 , n38823 );
nand ( n216586 , n38819 , n216585 );
not ( n38826 , n35704 );
and ( n38827 , n216586 , n38826 );
not ( n38828 , n216586 );
not ( n38829 , n35703 );
not ( n38830 , n38829 );
and ( n38831 , n38828 , n38830 );
nor ( n38832 , n38827 , n38831 );
not ( n38833 , n38832 );
not ( n38834 , n37559 );
not ( n38835 , n37567 );
and ( n38836 , n38834 , n38835 );
and ( n38837 , n37559 , n37567 );
nor ( n38838 , n38836 , n38837 );
buf ( n38839 , n38838 );
not ( n38840 , n38839 );
not ( n216602 , n25787 );
not ( n216603 , n214870 );
or ( n38843 , n216602 , n216603 );
not ( n38844 , n37106 );
or ( n38845 , n38844 , n25787 );
nand ( n38846 , n38843 , n38845 );
not ( n38847 , n38846 );
and ( n38848 , n38840 , n38847 );
and ( n38849 , n38839 , n38846 );
nor ( n38850 , n38848 , n38849 );
not ( n38851 , n38850 );
nand ( n38852 , n38833 , n38851 );
not ( n38853 , n208545 );
buf ( n38854 , RI173f81e8_1546);
not ( n38855 , n38854 );
not ( n38856 , RI173af4f8_1901);
not ( n38857 , n38856 );
or ( n38858 , n38855 , n38857 );
not ( n38859 , RI173f81e8_1546);
buf ( n38860 , RI173af4f8_1901);
nand ( n38861 , n38859 , n38860 );
nand ( n38862 , n38858 , n38861 );
not ( n38863 , RI1733fce8_2130);
and ( n38864 , n38862 , n38863 );
not ( n38865 , n38862 );
and ( n38866 , n38865 , n34573 );
nor ( n38867 , n38864 , n38866 );
xor ( n38868 , n38867 , n35179 );
buf ( n38869 , RI19aaad80_2489);
nand ( n38870 , n26059 , n38869 );
buf ( n38871 , RI17494818_1012);
and ( n38872 , n38870 , n38871 );
not ( n38873 , n38870 );
not ( n38874 , RI17494818_1012);
and ( n38875 , n38873 , n38874 );
nor ( n38876 , n38872 , n38875 );
xnor ( n38877 , n38868 , n38876 );
not ( n38878 , n38877 );
not ( n38879 , n38878 );
or ( n38880 , n38853 , n38879 );
or ( n38881 , n38878 , n208545 );
nand ( n38882 , n38880 , n38881 );
buf ( n38883 , RI173cca30_1758);
not ( n38884 , n38883 );
not ( n38885 , RI173434b0_2113);
not ( n38886 , n38885 );
or ( n38887 , n38884 , n38886 );
not ( n38888 , RI173cca30_1758);
buf ( n38889 , RI173434b0_2113);
nand ( n38890 , n38888 , n38889 );
nand ( n38891 , n38887 , n38890 );
buf ( n38892 , RI17415a68_1402);
and ( n216654 , n38891 , n38892 );
not ( n216655 , n38891 );
not ( n38895 , RI17415a68_1402);
and ( n38896 , n216655 , n38895 );
nor ( n38897 , n216654 , n38896 );
buf ( n38898 , RI19a8d668_2701);
nand ( n38899 , n204493 , n38898 );
not ( n38900 , RI17469078_1224);
and ( n38901 , n38899 , n38900 );
not ( n38902 , n38899 );
buf ( n38903 , RI17469078_1224);
and ( n38904 , n38902 , n38903 );
nor ( n38905 , n38901 , n38904 );
xor ( n38906 , n38897 , n38905 );
xnor ( n38907 , n38906 , n26170 );
buf ( n38908 , n38907 );
and ( n38909 , n38882 , n38908 );
not ( n38910 , n38882 );
not ( n38911 , n38907 );
buf ( n38912 , n38911 );
and ( n38913 , n38910 , n38912 );
nor ( n38914 , n38909 , n38913 );
buf ( n38915 , n38914 );
and ( n38916 , n38852 , n38915 );
not ( n38917 , n38852 );
not ( n38918 , n38915 );
and ( n38919 , n38917 , n38918 );
nor ( n38920 , n38916 , n38919 );
xor ( n38921 , n38815 , n38920 );
not ( n38922 , n38711 );
not ( n38923 , n38679 );
nand ( n38924 , n38922 , n38923 );
not ( n38925 , n38924 );
not ( n38926 , n31344 );
not ( n38927 , n35501 );
not ( n38928 , n31317 );
or ( n38929 , n38927 , n38928 );
or ( n38930 , n31317 , n35501 );
nand ( n38931 , n38929 , n38930 );
not ( n38932 , n38931 );
or ( n38933 , n38926 , n38932 );
or ( n38934 , n38931 , n31344 );
nand ( n38935 , n38933 , n38934 );
buf ( n38936 , n38935 );
not ( n38937 , n38936 );
and ( n38938 , n38925 , n38937 );
and ( n38939 , n38924 , n38936 );
nor ( n38940 , n38938 , n38939 );
not ( n38941 , n38940 );
not ( n38942 , n26289 );
buf ( n38943 , RI173d5aa8_1714);
not ( n38944 , n38943 );
not ( n38945 , n204940 );
or ( n38946 , n38944 , n38945 );
not ( n38947 , RI173d5aa8_1714);
nand ( n38948 , n38947 , n204899 );
nand ( n38949 , n38946 , n38948 );
and ( n38950 , n38949 , n36386 );
not ( n38951 , n38949 );
and ( n38952 , n38951 , n36390 );
nor ( n38953 , n38950 , n38952 );
buf ( n38954 , RI19aca748_2252);
nand ( n216716 , n30640 , n38954 );
buf ( n216717 , RI174bbda0_826);
and ( n38957 , n216716 , n216717 );
not ( n38958 , n216716 );
not ( n38959 , RI174bbda0_826);
and ( n38960 , n38958 , n38959 );
nor ( n38961 , n38957 , n38960 );
xor ( n38962 , n38953 , n38961 );
buf ( n38963 , RI19a9af70_2605);
nand ( n38964 , n205124 , n38963 );
not ( n38965 , RI17471d90_1181);
and ( n38966 , n38964 , n38965 );
not ( n38967 , n38964 );
buf ( n38968 , RI17471d90_1181);
and ( n38969 , n38967 , n38968 );
nor ( n38970 , n38966 , n38969 );
xor ( n38971 , n38962 , n38970 );
not ( n38972 , n38971 );
not ( n38973 , n38972 );
not ( n38974 , n38973 );
or ( n38975 , n38942 , n38974 );
or ( n38976 , n38973 , n26289 );
nand ( n38977 , n38975 , n38976 );
buf ( n38978 , RI173f2fe0_1571);
not ( n38979 , n38978 );
not ( n38980 , RI173aa2f0_1926);
not ( n38981 , n38980 );
or ( n38982 , n38979 , n38981 );
not ( n38983 , RI173f2fe0_1571);
buf ( n38984 , RI173aa2f0_1926);
nand ( n38985 , n38983 , n38984 );
nand ( n38986 , n38982 , n38985 );
and ( n38987 , n38986 , n28883 );
not ( n38988 , n38986 );
not ( n38989 , RI174c8be0_786);
and ( n38990 , n38988 , n38989 );
nor ( n38991 , n38987 , n38990 );
xor ( n38992 , n38991 , n207228 );
buf ( n38993 , RI19aaeea8_2462);
nand ( n38994 , n28637 , n38993 );
buf ( n38995 , RI1748f610_1037);
and ( n38996 , n38994 , n38995 );
not ( n38997 , n38994 );
not ( n38998 , RI1748f610_1037);
and ( n38999 , n38997 , n38998 );
nor ( n39000 , n38996 , n38999 );
xor ( n39001 , n38992 , n39000 );
buf ( n39002 , n39001 );
and ( n39003 , n38977 , n39002 );
not ( n39004 , n38977 );
xor ( n39005 , n38991 , n207228 );
xnor ( n39006 , n39005 , n39000 );
buf ( n39007 , n39006 );
not ( n39008 , n39007 );
not ( n39009 , n39008 );
and ( n39010 , n39004 , n39009 );
nor ( n39011 , n39003 , n39010 );
not ( n39012 , n39011 );
nor ( n39013 , n36812 , n33072 );
not ( n39014 , n39013 );
nand ( n39015 , n36813 , n33072 );
nand ( n39016 , n39014 , n39015 );
not ( n39017 , RI174bdc90_820);
xor ( n39018 , n39017 , n37874 );
xnor ( n39019 , n39018 , n37881 );
buf ( n39020 , n39019 );
and ( n39021 , n39016 , n39020 );
not ( n39022 , n39016 );
buf ( n39023 , n37882 );
and ( n39024 , n39022 , n39023 );
nor ( n39025 , n39021 , n39024 );
not ( n39026 , n39025 );
nand ( n39027 , n39012 , n39026 );
not ( n39028 , n26075 );
not ( n39029 , n32729 );
or ( n39030 , n39028 , n39029 );
not ( n39031 , n26075 );
nand ( n39032 , n39031 , n37455 );
nand ( n39033 , n39030 , n39032 );
and ( n39034 , n39033 , n32783 );
not ( n39035 , n39033 );
not ( n39036 , n32768 );
and ( n39037 , n39035 , n39036 );
nor ( n39038 , n39034 , n39037 );
not ( n39039 , n39038 );
and ( n39040 , n39027 , n39039 );
not ( n39041 , n39027 );
and ( n39042 , n39041 , n39038 );
nor ( n39043 , n39040 , n39042 );
not ( n39044 , n39043 );
and ( n39045 , n38941 , n39044 );
and ( n39046 , n38940 , n39043 );
nor ( n39047 , n39045 , n39046 );
not ( n39048 , n39047 );
and ( n39049 , n38921 , n39048 );
not ( n39050 , n38921 );
and ( n39051 , n39050 , n39047 );
nor ( n39052 , n39049 , n39051 );
not ( n39053 , n39052 );
or ( n39054 , n38717 , n39053 );
not ( n39055 , n38716 );
and ( n39056 , n38921 , n39047 );
not ( n39057 , n38921 );
and ( n39058 , n39057 , n39048 );
nor ( n39059 , n39056 , n39058 );
nand ( n39060 , n39055 , n39059 );
nand ( n39061 , n39054 , n39060 );
buf ( n39062 , n33085 );
not ( n39063 , n39062 );
xor ( n39064 , n36793 , n36810 );
xnor ( n39065 , n39064 , n36801 );
not ( n39066 , n39065 );
or ( n39067 , n39063 , n39066 );
or ( n39068 , n39065 , n39062 );
nand ( n216830 , n39067 , n39068 );
not ( n216831 , n216830 );
not ( n39071 , n216831 );
not ( n39072 , n39023 );
or ( n39073 , n39071 , n39072 );
nand ( n39074 , n39020 , n216830 );
nand ( n39075 , n39073 , n39074 );
buf ( n39076 , RI19a9d9a0_2587);
nand ( n39077 , n206902 , n39076 );
buf ( n39078 , RI1748b470_1057);
xor ( n39079 , n39077 , n39078 );
not ( n39080 , n39079 );
not ( n39081 , n38201 );
or ( n39082 , n39080 , n39081 );
or ( n39083 , n38201 , n39079 );
nand ( n39084 , n39082 , n39083 );
and ( n39085 , n39084 , n38205 );
not ( n39086 , n39084 );
and ( n39087 , n39086 , n38204 );
nor ( n39088 , n39085 , n39087 );
nand ( n39089 , n39075 , n39088 );
not ( n39090 , n39089 );
not ( n39091 , n27943 );
not ( n39092 , n33848 );
or ( n39093 , n39091 , n39092 );
or ( n39094 , n33849 , n27943 );
nand ( n39095 , n39093 , n39094 );
not ( n39096 , n39095 );
not ( n39097 , n39096 );
not ( n39098 , n33858 );
or ( n39099 , n39097 , n39098 );
nand ( n39100 , n36258 , n39095 );
nand ( n39101 , n39099 , n39100 );
not ( n39102 , n39101 );
or ( n39103 , n39090 , n39102 );
or ( n39104 , n39101 , n39089 );
nand ( n39105 , n39103 , n39104 );
not ( n216867 , n39105 );
buf ( n216868 , RI17499d68_986);
not ( n39108 , n207493 );
and ( n39109 , n216868 , n39108 );
not ( n39110 , n216868 );
and ( n39111 , n39110 , n207493 );
or ( n39112 , n39109 , n39111 );
and ( n39113 , n39112 , n33444 );
not ( n39114 , n39112 );
and ( n39115 , n39114 , n34594 );
nor ( n39116 , n39113 , n39115 );
not ( n39117 , n39116 );
buf ( n39118 , RI19aabcf8_2483);
nand ( n39119 , n29203 , n39118 );
buf ( n39120 , RI17492400_1023);
and ( n39121 , n39119 , n39120 );
not ( n39122 , n39119 );
not ( n39123 , RI17492400_1023);
and ( n39124 , n39122 , n39123 );
nor ( n39125 , n39121 , n39124 );
not ( n39126 , n39125 );
not ( n39127 , n26050 );
or ( n39128 , n39126 , n39127 );
or ( n39129 , n26050 , n39125 );
nand ( n39130 , n39128 , n39129 );
not ( n39131 , n39130 );
not ( n39132 , n39131 );
not ( n39133 , n38586 );
or ( n39134 , n39132 , n39133 );
nand ( n39135 , n26008 , n39130 );
nand ( n39136 , n39134 , n39135 );
not ( n39137 , n29983 );
not ( n39138 , n204792 );
or ( n39139 , n39137 , n39138 );
not ( n39140 , n29983 );
nand ( n39141 , n39140 , n204791 );
nand ( n39142 , n39139 , n39141 );
and ( n39143 , n39142 , n36309 );
not ( n39144 , n39142 );
not ( n39145 , n36309 );
and ( n39146 , n39144 , n39145 );
nor ( n39147 , n39143 , n39146 );
nor ( n39148 , n39136 , n39147 );
not ( n39149 , n39148 );
or ( n39150 , n39117 , n39149 );
or ( n39151 , n39148 , n39116 );
nand ( n39152 , n39150 , n39151 );
not ( n39153 , n39152 );
not ( n39154 , n39153 );
or ( n39155 , n216867 , n39154 );
not ( n39156 , n39105 );
nand ( n39157 , n39156 , n39152 );
nand ( n216919 , n39155 , n39157 );
buf ( n216920 , n29443 );
not ( n39160 , n216920 );
not ( n39161 , n33404 );
or ( n39162 , n39160 , n39161 );
not ( n39163 , n216920 );
nand ( n39164 , n39163 , n33403 );
nand ( n39165 , n39162 , n39164 );
and ( n39166 , n39165 , n34464 );
not ( n39167 , n39165 );
and ( n39168 , n39167 , n34461 );
nor ( n39169 , n39166 , n39168 );
not ( n39170 , n39169 );
not ( n39171 , n30578 );
not ( n39172 , n38764 );
or ( n39173 , n39171 , n39172 );
not ( n39174 , n30578 );
nand ( n39175 , n39174 , n38763 );
nand ( n39176 , n39173 , n39175 );
and ( n39177 , n39176 , n38771 );
not ( n39178 , n39176 );
and ( n39179 , n39178 , n38770 );
nor ( n39180 , n39177 , n39179 );
nand ( n39181 , n39170 , n39180 );
not ( n39182 , n39181 );
not ( n39183 , n38306 );
not ( n39184 , RI173a9fa8_1927);
not ( n39185 , n39184 );
or ( n39186 , n39183 , n39185 );
not ( n216948 , RI173f2c98_1572);
buf ( n216949 , RI173a9fa8_1927);
nand ( n39189 , n216948 , n216949 );
nand ( n216951 , n39186 , n39189 );
buf ( n216952 , RI174c5328_797);
and ( n39192 , n216951 , n216952 );
not ( n39193 , n216951 );
not ( n39194 , RI174c5328_797);
and ( n39195 , n39193 , n39194 );
nor ( n39196 , n39192 , n39195 );
buf ( n39197 , RI19aaeb60_2463);
nand ( n39198 , n204493 , n39197 );
buf ( n39199 , RI1748f2c8_1038);
and ( n39200 , n39198 , n39199 );
not ( n39201 , n39198 );
not ( n39202 , RI1748f2c8_1038);
and ( n39203 , n39201 , n39202 );
nor ( n39204 , n39200 , n39203 );
xor ( n39205 , n39196 , n39204 );
xnor ( n39206 , n39205 , n28414 );
not ( n39207 , n39206 );
not ( n39208 , n39207 );
not ( n39209 , n33968 );
and ( n39210 , n39208 , n39209 );
buf ( n39211 , n39206 );
not ( n39212 , n39211 );
and ( n39213 , n39212 , n33968 );
nor ( n39214 , n39210 , n39213 );
buf ( n39215 , RI173c74e0_1784);
not ( n39216 , n39215 );
not ( n39217 , RI1733df60_2139);
not ( n39218 , n39217 );
or ( n39219 , n39216 , n39218 );
not ( n39220 , RI173c74e0_1784);
buf ( n39221 , RI1733df60_2139);
nand ( n39222 , n39220 , n39221 );
nand ( n39223 , n39219 , n39222 );
not ( n216985 , RI174101d0_1429);
and ( n216986 , n39223 , n216985 );
not ( n39226 , n39223 );
buf ( n39227 , RI174101d0_1429);
and ( n39228 , n39226 , n39227 );
nor ( n39229 , n216986 , n39228 );
not ( n39230 , n39229 );
buf ( n39231 , RI19ac1490_2320);
nand ( n39232 , n26028 , n39231 );
buf ( n39233 , RI174ac800_895);
xor ( n39234 , n39232 , n39233 );
xor ( n39235 , n39230 , n39234 );
buf ( n216997 , RI19a91100_2675);
nand ( n216998 , n28637 , n216997 );
buf ( n216999 , RI17463b28_1250);
and ( n217000 , n216998 , n216999 );
not ( n39240 , n216998 );
not ( n217002 , RI17463b28_1250);
and ( n217003 , n39240 , n217002 );
nor ( n39243 , n217000 , n217003 );
xnor ( n39244 , n39235 , n39243 );
not ( n39245 , n39244 );
not ( n39246 , n39245 );
and ( n39247 , n39214 , n39246 );
not ( n39248 , n39214 );
xor ( n39249 , n39229 , n39234 );
xnor ( n39250 , n39249 , n39243 );
buf ( n39251 , n39250 );
and ( n39252 , n39248 , n39251 );
nor ( n39253 , n39247 , n39252 );
buf ( n39254 , n39253 );
not ( n39255 , n39254 );
and ( n39256 , n39182 , n39255 );
and ( n39257 , n39181 , n39254 );
nor ( n39258 , n39256 , n39257 );
and ( n39259 , n216919 , n39258 );
not ( n39260 , n216919 );
not ( n39261 , n39258 );
and ( n39262 , n39260 , n39261 );
nor ( n39263 , n39259 , n39262 );
not ( n39264 , n39263 );
not ( n39265 , n38839 );
not ( n39266 , n205235 );
not ( n39267 , n37105 );
not ( n39268 , n39267 );
or ( n39269 , n39266 , n39268 );
not ( n39270 , n205235 );
nand ( n39271 , n39270 , n37106 );
nand ( n39272 , n39269 , n39271 );
not ( n39273 , n39272 );
and ( n39274 , n39265 , n39273 );
and ( n39275 , n38839 , n39272 );
nor ( n39276 , n39274 , n39275 );
buf ( n39277 , n29201 );
not ( n39278 , n39277 );
not ( n39279 , n39278 );
not ( n39280 , n207960 );
or ( n39281 , n39279 , n39280 );
nand ( n39282 , n30205 , n39277 );
nand ( n39283 , n39281 , n39282 );
not ( n39284 , n39283 );
not ( n39285 , n31829 );
and ( n39286 , n39284 , n39285 );
and ( n39287 , n39283 , n31829 );
nor ( n39288 , n39286 , n39287 );
not ( n39289 , n39288 );
nand ( n39290 , n39276 , n39289 );
not ( n39291 , n39290 );
not ( n39292 , n31401 );
buf ( n39293 , RI174025f8_1496);
not ( n217055 , n39293 );
not ( n217056 , RI173b9908_1851);
not ( n39296 , n217056 );
or ( n39297 , n217055 , n39296 );
not ( n39298 , RI174025f8_1496);
buf ( n39299 , RI173b9908_1851);
nand ( n39300 , n39298 , n39299 );
nand ( n39301 , n39297 , n39300 );
not ( n39302 , n39301 );
buf ( n39303 , RI17532e40_608);
xor ( n39304 , n39303 , n204993 );
buf ( n39305 , RI19ab92b8_2387);
nand ( n39306 , n25751 , n39305 );
not ( n39307 , RI1749e8e0_963);
and ( n39308 , n39306 , n39307 );
not ( n39309 , n39306 );
buf ( n217071 , RI1749e8e0_963);
and ( n217072 , n39309 , n217071 );
nor ( n39312 , n39308 , n217072 );
xnor ( n39313 , n39304 , n39312 );
not ( n39314 , n39313 );
or ( n39315 , n39302 , n39314 );
not ( n39316 , n39313 );
not ( n39317 , n39301 );
nand ( n39318 , n39316 , n39317 );
nand ( n39319 , n39315 , n39318 );
buf ( n39320 , n39319 );
not ( n39321 , n39320 );
or ( n39322 , n39292 , n39321 );
or ( n39323 , n39320 , n31401 );
nand ( n39324 , n39322 , n39323 );
and ( n39325 , n39324 , n204825 );
not ( n39326 , n39324 );
not ( n39327 , n204825 );
and ( n39328 , n39326 , n39327 );
nor ( n39329 , n39325 , n39328 );
not ( n39330 , n39329 );
not ( n39331 , n39330 );
or ( n39332 , n39291 , n39331 );
or ( n39333 , n39330 , n39290 );
nand ( n39334 , n39332 , n39333 );
not ( n39335 , n39334 );
buf ( n39336 , RI173dacb0_1689);
not ( n39337 , n39336 );
not ( n39338 , RI17391fc0_2044);
not ( n39339 , n39338 );
or ( n39340 , n39337 , n39339 );
not ( n39341 , RI173dacb0_1689);
nand ( n39342 , n39341 , n32367 );
nand ( n39343 , n39340 , n39342 );
buf ( n39344 , RI17452788_1334);
and ( n39345 , n39343 , n39344 );
not ( n39346 , n39343 );
not ( n39347 , RI17452788_1334);
and ( n39348 , n39346 , n39347 );
nor ( n39349 , n39345 , n39348 );
buf ( n39350 , RI19a97208_2632);
nand ( n217112 , n25628 , n39350 );
buf ( n217113 , RI17476f98_1156);
and ( n39353 , n217112 , n217113 );
not ( n217115 , n217112 );
not ( n39355 , RI17476f98_1156);
and ( n217117 , n217115 , n39355 );
nor ( n217118 , n39353 , n217117 );
xor ( n39358 , n39349 , n217118 );
xnor ( n39359 , n39358 , n38367 );
not ( n39360 , n39359 );
not ( n39361 , n39360 );
xor ( n39362 , n32320 , n39361 );
xnor ( n39363 , n39362 , n215031 );
buf ( n39364 , n29115 );
not ( n39365 , n39364 );
not ( n39366 , n29112 );
and ( n39367 , n39365 , n39366 );
and ( n39368 , n39364 , n29112 );
nor ( n39369 , n39367 , n39368 );
not ( n39370 , n39369 );
not ( n39371 , n210587 );
or ( n39372 , n39370 , n39371 );
or ( n39373 , n210587 , n39369 );
nand ( n39374 , n39372 , n39373 );
not ( n39375 , n39374 );
not ( n39376 , n38034 );
not ( n39377 , n32516 );
or ( n39378 , n39376 , n39377 );
or ( n39379 , n38034 , n32516 );
nand ( n39380 , n39378 , n39379 );
buf ( n39381 , RI173ca2d0_1770);
not ( n39382 , n39381 );
not ( n39383 , RI17340d50_2125);
not ( n39384 , n39383 );
or ( n39385 , n39382 , n39384 );
not ( n39386 , RI173ca2d0_1770);
buf ( n39387 , RI17340d50_2125);
nand ( n39388 , n39386 , n39387 );
nand ( n39389 , n39385 , n39388 );
buf ( n39390 , RI17413308_1414);
and ( n39391 , n39389 , n39390 );
not ( n39392 , n39389 );
not ( n39393 , RI17413308_1414);
and ( n39394 , n39392 , n39393 );
nor ( n39395 , n39391 , n39394 );
not ( n39396 , n39395 );
and ( n39397 , n39380 , n39396 );
not ( n39398 , n39380 );
and ( n39399 , n39398 , n39395 );
nor ( n39400 , n39397 , n39399 );
buf ( n39401 , n39400 );
buf ( n39402 , n39401 );
not ( n39403 , n39402 );
and ( n39404 , n39375 , n39403 );
and ( n39405 , n39374 , n39401 );
nor ( n39406 , n39404 , n39405 );
nand ( n39407 , n39363 , n39406 );
not ( n39408 , n39407 );
buf ( n39409 , RI173a95d0_1930);
not ( n39410 , n39409 );
not ( n39411 , n32655 );
not ( n39412 , n39411 );
or ( n39413 , n39410 , n39412 );
not ( n39414 , RI173a95d0_1930);
nand ( n39415 , n32655 , n39414 );
nand ( n39416 , n39413 , n39415 );
buf ( n39417 , n32685 );
buf ( n39418 , n39417 );
xnor ( n39419 , n39416 , n39418 );
not ( n39420 , n39419 );
and ( n39421 , n39408 , n39420 );
not ( n39422 , n39406 );
not ( n39423 , n39422 );
nand ( n39424 , n39423 , n39363 );
and ( n39425 , n39424 , n39419 );
nor ( n39426 , n39421 , n39425 );
not ( n39427 , n39426 );
or ( n39428 , n39335 , n39427 );
or ( n217190 , n39426 , n39334 );
nand ( n217191 , n39428 , n217190 );
not ( n39431 , n217191 );
and ( n39432 , n39264 , n39431 );
and ( n39433 , n39263 , n217191 );
nor ( n39434 , n39432 , n39433 );
buf ( n39435 , n39434 );
and ( n39436 , n39061 , n39435 );
not ( n39437 , n39061 );
not ( n39438 , n39263 );
not ( n39439 , n39438 );
not ( n39440 , n217191 );
not ( n39441 , n39440 );
or ( n39442 , n39439 , n39441 );
nand ( n39443 , n39263 , n217191 );
nand ( n39444 , n39442 , n39443 );
buf ( n39445 , n39444 );
and ( n39446 , n39437 , n39445 );
nor ( n39447 , n39436 , n39446 );
buf ( n39448 , RI173c6130_1790);
not ( n39449 , n39448 );
not ( n39450 , RI1733cbb0_2145);
not ( n39451 , n39450 );
or ( n39452 , n39449 , n39451 );
not ( n39453 , RI173c6130_1790);
buf ( n39454 , RI1733cbb0_2145);
nand ( n39455 , n39453 , n39454 );
nand ( n39456 , n39452 , n39455 );
not ( n39457 , RI1740ee20_1435);
and ( n39458 , n39456 , n39457 );
not ( n39459 , n39456 );
and ( n39460 , n39459 , n38055 );
nor ( n39461 , n39458 , n39460 );
buf ( n39462 , RI19a92bb8_2663);
nand ( n39463 , n25583 , n39462 );
buf ( n39464 , RI17462778_1256);
and ( n39465 , n39463 , n39464 );
not ( n39466 , n39463 );
not ( n39467 , RI17462778_1256);
and ( n39468 , n39466 , n39467 );
nor ( n39469 , n39465 , n39468 );
xor ( n39470 , n39461 , n39469 );
buf ( n39471 , RI19ac2f48_2307);
nand ( n39472 , n25712 , n39471 );
not ( n39473 , RI174ab450_901);
and ( n39474 , n39472 , n39473 );
not ( n39475 , n39472 );
buf ( n39476 , RI174ab450_901);
and ( n39477 , n39475 , n39476 );
nor ( n39478 , n39474 , n39477 );
xnor ( n39479 , n39470 , n39478 );
buf ( n39480 , n39479 );
buf ( n39481 , n39480 );
not ( n217243 , n39481 );
buf ( n217244 , RI19aba398_2379);
nand ( n39484 , n25452 , n217244 );
buf ( n39485 , RI1749c810_973);
and ( n39486 , n39484 , n39485 );
not ( n39487 , n39484 );
not ( n39488 , RI1749c810_973);
and ( n39489 , n39487 , n39488 );
nor ( n39490 , n39486 , n39489 );
nor ( n39491 , n30769 , n39490 );
not ( n39492 , n39491 );
nand ( n39493 , n30769 , n39490 );
nand ( n39494 , n39492 , n39493 );
not ( n39495 , n39494 );
or ( n39496 , n217243 , n39495 );
or ( n39497 , n39494 , n39480 );
nand ( n39498 , n39496 , n39497 );
not ( n39499 , n39498 );
not ( n39500 , n31423 );
not ( n39501 , n39319 );
not ( n39502 , n39501 );
or ( n39503 , n39500 , n39502 );
not ( n39504 , n31423 );
nand ( n39505 , n39504 , n39319 );
nand ( n39506 , n39503 , n39505 );
and ( n39507 , n39506 , n39327 );
not ( n39508 , n39506 );
and ( n39509 , n39508 , n204825 );
nor ( n39510 , n39507 , n39509 );
nand ( n39511 , n39499 , n39510 );
and ( n39512 , n39511 , n34585 );
not ( n39513 , n39511 );
and ( n39514 , n39513 , n34586 );
nor ( n39515 , n39512 , n39514 );
not ( n39516 , n39515 );
nand ( n39517 , n34585 , n39498 );
and ( n39518 , n39517 , n34601 );
not ( n39519 , n39517 );
and ( n39520 , n39519 , n34600 );
nor ( n39521 , n39518 , n39520 );
not ( n39522 , n39521 );
not ( n39523 , n34570 );
or ( n39524 , n39522 , n39523 );
or ( n39525 , n34570 , n39521 );
nand ( n39526 , n39524 , n39525 );
not ( n39527 , n36749 );
not ( n39528 , n28968 );
or ( n39529 , n39527 , n39528 );
or ( n39530 , n28968 , n36749 );
nand ( n39531 , n39529 , n39530 );
xor ( n39532 , n33000 , n205175 );
and ( n39533 , n39531 , n39532 );
not ( n39534 , n39531 );
and ( n39535 , n39534 , n33002 );
nor ( n39536 , n39533 , n39535 );
not ( n39537 , n39536 );
nand ( n39538 , n34737 , n39537 );
not ( n39539 , n39538 );
not ( n39540 , n34745 );
and ( n39541 , n39539 , n39540 );
and ( n39542 , n39538 , n34745 );
nor ( n39543 , n39541 , n39542 );
and ( n39544 , n39526 , n39543 );
not ( n39545 , n39526 );
not ( n39546 , n39543 );
and ( n39547 , n39545 , n39546 );
nor ( n39548 , n39544 , n39547 );
not ( n39549 , n33352 );
not ( n39550 , n39549 );
not ( n39551 , n30580 );
or ( n39552 , n39550 , n39551 );
not ( n39553 , n30579 );
not ( n39554 , n39553 );
not ( n39555 , n39554 );
nand ( n39556 , n39555 , n33352 );
nand ( n39557 , n39552 , n39556 );
buf ( n39558 , n35156 );
not ( n39559 , n39558 );
and ( n39560 , n39557 , n39559 );
not ( n39561 , n39557 );
and ( n39562 , n39561 , n39558 );
nor ( n39563 , n39560 , n39562 );
nand ( n39564 , n39563 , n34941 );
and ( n39565 , n39564 , n34932 );
not ( n39566 , n39564 );
and ( n217328 , n39566 , n34931 );
nor ( n217329 , n39565 , n217328 );
buf ( n39569 , n35888 );
not ( n39570 , n26134 );
and ( n39571 , n39570 , n32766 );
not ( n39572 , n39570 );
and ( n39573 , n39572 , n32781 );
nor ( n39574 , n39571 , n39573 );
not ( n217336 , n39574 );
and ( n217337 , n39569 , n217336 );
not ( n217338 , n39569 );
and ( n217339 , n217338 , n39574 );
nor ( n39579 , n217337 , n217339 );
nand ( n39580 , n34826 , n39579 );
not ( n39581 , n39580 );
not ( n39582 , n34817 );
and ( n39583 , n39581 , n39582 );
and ( n39584 , n39580 , n34817 );
nor ( n39585 , n39583 , n39584 );
and ( n39586 , n217329 , n39585 );
not ( n39587 , n217329 );
not ( n39588 , n39585 );
and ( n39589 , n39587 , n39588 );
nor ( n39590 , n39586 , n39589 );
not ( n39591 , n39590 );
and ( n39592 , n39548 , n39591 );
not ( n39593 , n39548 );
and ( n39594 , n39593 , n39590 );
nor ( n39595 , n39592 , n39594 );
not ( n39596 , n39595 );
or ( n39597 , n39516 , n39596 );
not ( n39598 , n39595 );
not ( n39599 , n39515 );
nand ( n39600 , n39598 , n39599 );
nand ( n39601 , n39597 , n39600 );
buf ( n39602 , n35109 );
not ( n39603 , n39602 );
and ( n39604 , n29761 , n34237 );
not ( n39605 , n29761 );
and ( n39606 , n39605 , n34233 );
nor ( n39607 , n39604 , n39606 );
xor ( n39608 , n39607 , n29768 );
buf ( n39609 , RI173de130_1673);
not ( n39610 , n39609 );
not ( n39611 , RI17395440_2028);
not ( n39612 , n39611 );
or ( n39613 , n39610 , n39612 );
not ( n39614 , RI173de130_1673);
buf ( n39615 , RI17395440_2028);
nand ( n39616 , n39614 , n39615 );
nand ( n39617 , n39613 , n39616 );
not ( n39618 , RI17455c08_1318);
and ( n39619 , n39617 , n39618 );
not ( n39620 , n39617 );
buf ( n39621 , RI17455c08_1318);
and ( n39622 , n39620 , n39621 );
nor ( n39623 , n39619 , n39622 );
buf ( n39624 , RI19ac6bc0_2279);
nand ( n39625 , n25405 , n39624 );
buf ( n39626 , RI174c9630_784);
and ( n39627 , n39625 , n39626 );
not ( n39628 , n39625 );
not ( n39629 , RI174c9630_784);
and ( n39630 , n39628 , n39629 );
nor ( n39631 , n39627 , n39630 );
xor ( n39632 , n39623 , n39631 );
buf ( n39633 , RI19a96e48_2634);
nand ( n39634 , n25666 , n39633 );
buf ( n39635 , RI1747a760_1139);
and ( n39636 , n39634 , n39635 );
not ( n39637 , n39634 );
not ( n39638 , RI1747a760_1139);
and ( n39639 , n39637 , n39638 );
nor ( n39640 , n39636 , n39639 );
xnor ( n39641 , n39632 , n39640 );
not ( n39642 , n39641 );
xor ( n39643 , n39608 , n39642 );
nand ( n39644 , n35118 , n39643 );
not ( n39645 , n39644 );
or ( n39646 , n39603 , n39645 );
or ( n39647 , n39602 , n39644 );
nand ( n39648 , n39646 , n39647 );
not ( n39649 , n39648 );
not ( n39650 , n32857 );
not ( n39651 , n28472 );
and ( n39652 , n39650 , n39651 );
and ( n39653 , n32857 , n28472 );
nor ( n39654 , n39652 , n39653 );
buf ( n39655 , n32847 );
xor ( n39656 , n39654 , n39655 );
xnor ( n39657 , n39656 , n210587 );
nand ( n39658 , n35030 , n39657 );
not ( n39659 , n39658 );
not ( n217421 , n35019 );
not ( n217422 , n217421 );
and ( n39662 , n39659 , n217422 );
and ( n39663 , n39658 , n217421 );
nor ( n39664 , n39662 , n39663 );
not ( n39665 , n39664 );
or ( n39666 , n39649 , n39665 );
or ( n39667 , n39648 , n39664 );
nand ( n39668 , n39666 , n39667 );
not ( n39669 , n30137 );
not ( n39670 , n204565 );
buf ( n39671 , n28380 );
not ( n39672 , n39671 );
or ( n39673 , n39670 , n39672 );
not ( n39674 , n204565 );
nand ( n39675 , n39674 , n28381 );
nand ( n39676 , n39673 , n39675 );
not ( n39677 , n39676 );
or ( n39678 , n39669 , n39677 );
not ( n39679 , n30140 );
or ( n39680 , n39676 , n39679 );
nand ( n39681 , n39678 , n39680 );
nand ( n39682 , n35192 , n39681 );
not ( n39683 , n39682 );
not ( n39684 , n35170 );
and ( n39685 , n39683 , n39684 );
and ( n39686 , n39682 , n35170 );
nor ( n39687 , n39685 , n39686 );
and ( n39688 , n39668 , n39687 );
not ( n39689 , n39668 );
not ( n39690 , n39687 );
and ( n39691 , n39689 , n39690 );
nor ( n39692 , n39688 , n39691 );
not ( n39693 , n39692 );
buf ( n39694 , RI173d01f8_1741);
not ( n39695 , RI17400528_1506);
buf ( n39696 , RI173b7838_1861);
and ( n39697 , n39695 , n39696 );
not ( n39698 , n39695 );
not ( n39699 , RI173b7838_1861);
and ( n39700 , n39698 , n39699 );
nor ( n39701 , n39697 , n39700 );
xor ( n39702 , n39694 , n39701 );
buf ( n39703 , RI1752fab0_618);
xor ( n39704 , n39703 , n39485 );
xnor ( n39705 , n39704 , n39484 );
xnor ( n39706 , n39702 , n39705 );
buf ( n39707 , n39706 );
not ( n39708 , n37423 );
not ( n39709 , n31900 );
or ( n39710 , n39708 , n39709 );
or ( n39711 , n31900 , n37423 );
nand ( n39712 , n39710 , n39711 );
and ( n217474 , n39707 , n39712 );
not ( n217475 , n39707 );
not ( n39715 , n39712 );
and ( n217477 , n217475 , n39715 );
nor ( n217478 , n217474 , n217477 );
nand ( n39718 , n217478 , n35286 );
not ( n39719 , n39718 );
not ( n39720 , n35232 );
not ( n39721 , n39720 );
and ( n39722 , n39719 , n39721 );
and ( n39723 , n39718 , n39720 );
nor ( n39724 , n39722 , n39723 );
not ( n39725 , n39724 );
not ( n39726 , n37837 );
not ( n39727 , n38130 );
or ( n39728 , n39726 , n39727 );
or ( n39729 , n37837 , n38130 );
nand ( n39730 , n39728 , n39729 );
and ( n39731 , n39730 , n38137 );
not ( n39732 , n39730 );
not ( n39733 , n38137 );
and ( n39734 , n39732 , n39733 );
nor ( n39735 , n39731 , n39734 );
nand ( n39736 , n35302 , n39735 );
and ( n39737 , n39736 , n35321 );
not ( n39738 , n39736 );
and ( n39739 , n39738 , n35320 );
nor ( n39740 , n39737 , n39739 );
not ( n39741 , n39740 );
or ( n39742 , n39725 , n39741 );
or ( n39743 , n39740 , n39724 );
nand ( n39744 , n39742 , n39743 );
not ( n39745 , n39744 );
and ( n39746 , n39693 , n39745 );
and ( n39747 , n39744 , n39692 );
nor ( n39748 , n39746 , n39747 );
not ( n39749 , n39748 );
not ( n217511 , n39749 );
and ( n217512 , n39601 , n217511 );
not ( n39752 , n39601 );
not ( n217514 , n39748 );
buf ( n217515 , n217514 );
buf ( n39755 , n217515 );
and ( n39756 , n39752 , n39755 );
nor ( n39757 , n217512 , n39756 );
nand ( n39758 , n39447 , n39757 );
or ( n39759 , n38639 , n39758 );
not ( n39760 , n39757 );
not ( n39761 , n38636 );
or ( n39762 , n39760 , n39761 );
buf ( n39763 , n35427 );
nor ( n39764 , n39447 , n39763 );
nand ( n39765 , n39762 , n39764 );
buf ( n39766 , n31575 );
buf ( n39767 , n39766 );
nand ( n39768 , n39767 , n32409 );
nand ( n39769 , n39759 , n39765 , n39768 );
buf ( n39770 , n39769 );
buf ( n39771 , RI173a0570_1974);
not ( n39772 , n39771 );
not ( n39773 , n32219 );
or ( n39774 , n39772 , n39773 );
or ( n39775 , n32219 , n39771 );
nand ( n39776 , n39774 , n39775 );
and ( n39777 , n39776 , n32236 );
not ( n39778 , n39776 );
and ( n39779 , n39778 , n210002 );
nor ( n39780 , n39777 , n39779 );
not ( n39781 , n39780 );
not ( n39782 , n33656 );
not ( n39783 , n204259 );
or ( n39784 , n39782 , n39783 );
not ( n39785 , n33656 );
nand ( n39786 , n39785 , n204258 );
nand ( n39787 , n39784 , n39786 );
xor ( n39788 , n39787 , n32136 );
not ( n39789 , n25426 );
buf ( n39790 , RI1749f948_958);
not ( n39791 , n39790 );
buf ( n39792 , n28068 );
not ( n39793 , n39792 );
or ( n39794 , n39791 , n39793 );
or ( n39795 , n39792 , n39790 );
nand ( n39796 , n39794 , n39795 );
not ( n39797 , n39796 );
buf ( n39798 , n25385 );
not ( n39799 , n39798 );
or ( n39800 , n39797 , n39799 );
not ( n39801 , n39796 );
not ( n39802 , n25372 );
not ( n39803 , n25384 );
or ( n39804 , n39802 , n39803 );
or ( n39805 , n25372 , n25384 );
nand ( n39806 , n39804 , n39805 );
not ( n39807 , n25357 );
and ( n39808 , n39806 , n39807 );
not ( n39809 , n39806 );
and ( n39810 , n39809 , n25357 );
nor ( n39811 , n39808 , n39810 );
nand ( n39812 , n39801 , n39811 );
nand ( n39813 , n39800 , n39812 );
not ( n39814 , n39813 );
or ( n39815 , n39789 , n39814 );
or ( n39816 , n39813 , n25426 );
nand ( n39817 , n39815 , n39816 );
nor ( n39818 , n39788 , n39817 );
not ( n39819 , n39818 );
and ( n39820 , n39781 , n39819 );
and ( n39821 , n39780 , n39818 );
nor ( n39822 , n39820 , n39821 );
not ( n39823 , n39822 );
not ( n217585 , n39823 );
xor ( n217586 , n204910 , n36018 );
xnor ( n39826 , n217586 , n34004 );
buf ( n217588 , RI173ef188_1590);
not ( n217589 , n217588 );
not ( n39829 , RI173a6498_1945);
not ( n39830 , n39829 );
or ( n39831 , n217589 , n39830 );
not ( n39832 , RI173ef188_1590);
buf ( n39833 , RI173a6498_1945);
nand ( n39834 , n39832 , n39833 );
nand ( n39835 , n39831 , n39834 );
buf ( n39836 , RI1749c180_975);
and ( n39837 , n39835 , n39836 );
not ( n39838 , n39835 );
not ( n39839 , RI1749c180_975);
and ( n39840 , n39838 , n39839 );
nor ( n39841 , n39837 , n39840 );
not ( n39842 , n39841 );
xor ( n39843 , n39842 , n39079 );
xnor ( n39844 , n39843 , n38151 );
buf ( n39845 , n39844 );
not ( n39846 , n39845 );
buf ( n39847 , n207491 );
not ( n39848 , n39847 );
xor ( n39849 , n34681 , n34689 );
xor ( n39850 , n39849 , n34698 );
not ( n39851 , n39850 );
or ( n39852 , n39848 , n39851 );
or ( n39853 , n39850 , n39847 );
nand ( n39854 , n39852 , n39853 );
not ( n39855 , n39854 );
or ( n39856 , n39846 , n39855 );
or ( n39857 , n39854 , n39845 );
nand ( n39858 , n39856 , n39857 );
buf ( n39859 , n39858 );
nand ( n39860 , n39826 , n39859 );
xor ( n39861 , n31951 , n35740 );
xnor ( n39862 , n39861 , n29088 );
not ( n39863 , n39862 );
and ( n39864 , n39860 , n39863 );
not ( n39865 , n39860 );
and ( n39866 , n39865 , n39862 );
nor ( n39867 , n39864 , n39866 );
not ( n39868 , n39867 );
not ( n39869 , n39868 );
nand ( n39870 , n39780 , n39817 );
not ( n39871 , n39870 );
not ( n39872 , n35071 );
not ( n39873 , n38088 );
buf ( n39874 , n39873 );
not ( n39875 , n39874 );
not ( n39876 , n39875 );
or ( n39877 , n39872 , n39876 );
nand ( n39878 , n38090 , n35067 );
nand ( n39879 , n39877 , n39878 );
xnor ( n39880 , n39879 , n204672 );
buf ( n39881 , n39880 );
not ( n39882 , n39881 );
and ( n39883 , n39871 , n39882 );
and ( n39884 , n39870 , n39881 );
nor ( n39885 , n39883 , n39884 );
not ( n39886 , n39885 );
not ( n39887 , n39886 );
or ( n39888 , n39869 , n39887 );
nand ( n39889 , n39885 , n39867 );
nand ( n217651 , n39888 , n39889 );
not ( n217652 , n30661 );
not ( n39892 , n37864 );
or ( n39893 , n217652 , n39892 );
or ( n39894 , n37864 , n30661 );
nand ( n39895 , n39893 , n39894 );
buf ( n39896 , RI173fcd60_1523);
not ( n39897 , n39896 );
not ( n39898 , RI173b3d28_1879);
not ( n39899 , n39898 );
or ( n39900 , n39897 , n39899 );
not ( n39901 , RI173fcd60_1523);
buf ( n39902 , RI173b3d28_1879);
nand ( n39903 , n39901 , n39902 );
nand ( n39904 , n39900 , n39903 );
not ( n39905 , RI173ade00_1908);
and ( n39906 , n39904 , n39905 );
not ( n39907 , n39904 );
buf ( n39908 , RI173ade00_1908);
and ( n39909 , n39907 , n39908 );
nor ( n39910 , n39906 , n39909 );
xor ( n39911 , n39910 , n25636 );
buf ( n39912 , RI19aa90e8_2502);
nand ( n39913 , n25405 , n39912 );
buf ( n39914 , RI17499048_990);
and ( n39915 , n39913 , n39914 );
not ( n39916 , n39913 );
not ( n39917 , RI17499048_990);
and ( n39918 , n39916 , n39917 );
nor ( n39919 , n39915 , n39918 );
not ( n39920 , n39919 );
xor ( n39921 , n39911 , n39920 );
not ( n39922 , n39921 );
xor ( n39923 , n39895 , n39922 );
buf ( n39924 , n35517 );
not ( n39925 , n39924 );
not ( n39926 , n31323 );
or ( n39927 , n39925 , n39926 );
or ( n39928 , n31323 , n39924 );
nand ( n39929 , n39927 , n39928 );
and ( n39930 , n39929 , n31343 );
not ( n39931 , n39929 );
and ( n39932 , n39931 , n31344 );
nor ( n39933 , n39930 , n39932 );
nand ( n39934 , n39923 , n39933 );
not ( n39935 , n39934 );
not ( n39936 , n35675 );
buf ( n39937 , RI173cd0c0_1756);
not ( n39938 , n39937 );
not ( n39939 , RI17343b40_2111);
not ( n39940 , n39939 );
or ( n39941 , n39938 , n39940 );
not ( n39942 , RI173cd0c0_1756);
buf ( n39943 , RI17343b40_2111);
nand ( n39944 , n39942 , n39943 );
nand ( n39945 , n39941 , n39944 );
not ( n39946 , RI17444ef8_1400);
and ( n39947 , n39945 , n39946 );
not ( n39948 , n39945 );
and ( n39949 , n39948 , n28612 );
nor ( n39950 , n39947 , n39949 );
buf ( n39951 , RI19a8db18_2699);
nand ( n39952 , n25622 , n39951 );
buf ( n39953 , RI17469708_1222);
and ( n39954 , n39952 , n39953 );
not ( n39955 , n39952 );
not ( n217717 , RI17469708_1222);
and ( n217718 , n39955 , n217717 );
nor ( n39958 , n39954 , n217718 );
xor ( n39959 , n39950 , n39958 );
buf ( n39960 , RI19abe9e8_2344);
nand ( n39961 , n27706 , n39960 );
not ( n39962 , RI174b23e0_867);
and ( n39963 , n39961 , n39962 );
not ( n39964 , n39961 );
buf ( n39965 , RI174b23e0_867);
and ( n39966 , n39964 , n39965 );
nor ( n39967 , n39963 , n39966 );
xnor ( n39968 , n39959 , n39967 );
not ( n39969 , n39968 );
or ( n39970 , n39936 , n39969 );
not ( n39971 , n35675 );
not ( n39972 , n39958 );
xor ( n39973 , n39950 , n39972 );
xnor ( n39974 , n39973 , n39967 );
nand ( n39975 , n39971 , n39974 );
nand ( n39976 , n39970 , n39975 );
not ( n39977 , n32448 );
not ( n39978 , n38748 );
or ( n39979 , n39977 , n39978 );
not ( n39980 , RI173ea958_1612);
nand ( n39981 , n39980 , n38741 );
nand ( n39982 , n39979 , n39981 );
and ( n39983 , n39982 , n37513 );
not ( n39984 , n39982 );
not ( n39985 , RI1746e910_1197);
and ( n39986 , n39984 , n39985 );
nor ( n39987 , n39983 , n39986 );
buf ( n39988 , RI19a82970_2776);
nand ( n39989 , n25850 , n39988 );
buf ( n39990 , RI1750d820_724);
and ( n39991 , n39989 , n39990 );
not ( n39992 , n39989 );
not ( n39993 , RI1750d820_724);
and ( n39994 , n39992 , n39993 );
nor ( n39995 , n39991 , n39994 );
xor ( n39996 , n39987 , n39995 );
buf ( n39997 , RI19aa17f8_2556);
nand ( n39998 , n27946 , n39997 );
not ( n39999 , RI17486c40_1079);
and ( n40000 , n39998 , n39999 );
not ( n40001 , n39998 );
buf ( n40002 , RI17486c40_1079);
and ( n40003 , n40001 , n40002 );
nor ( n40004 , n40000 , n40003 );
xor ( n40005 , n39996 , n40004 );
not ( n40006 , n40005 );
not ( n40007 , n40006 );
and ( n40008 , n39976 , n40007 );
not ( n40009 , n39976 );
and ( n40010 , n40009 , n40006 );
nor ( n40011 , n40008 , n40010 );
not ( n40012 , n40011 );
not ( n40013 , n40012 );
and ( n40014 , n39935 , n40013 );
and ( n40015 , n39934 , n40012 );
nor ( n40016 , n40014 , n40015 );
not ( n40017 , n40016 );
not ( n40018 , n209114 );
not ( n40019 , n30900 );
not ( n40020 , RI1739c088_1995);
not ( n40021 , n40020 );
or ( n40022 , n40019 , n40021 );
not ( n40023 , RI173e50c0_1639);
buf ( n40024 , RI1739c088_1995);
nand ( n40025 , n40023 , n40024 );
nand ( n40026 , n40022 , n40025 );
buf ( n40027 , RI1745cb98_1284);
and ( n40028 , n40026 , n40027 );
not ( n40029 , n40026 );
not ( n40030 , RI1745cb98_1284);
and ( n40031 , n40029 , n40030 );
nor ( n40032 , n40028 , n40031 );
buf ( n40033 , RI19a86318_2751);
nand ( n40034 , n25851 , n40033 );
not ( n40035 , RI17502e70_751);
and ( n40036 , n40034 , n40035 );
not ( n40037 , n40034 );
buf ( n40038 , RI17502e70_751);
and ( n40039 , n40037 , n40038 );
nor ( n40040 , n40036 , n40039 );
not ( n40041 , n40040 );
xor ( n40042 , n40032 , n40041 );
buf ( n40043 , RI19aa4ed0_2530);
nand ( n40044 , n204336 , n40043 );
buf ( n40045 , RI174813a8_1106);
and ( n40046 , n40044 , n40045 );
not ( n40047 , n40044 );
not ( n40048 , RI174813a8_1106);
and ( n40049 , n40047 , n40048 );
nor ( n40050 , n40046 , n40049 );
buf ( n40051 , n40050 );
xor ( n40052 , n40042 , n40051 );
not ( n40053 , n40052 );
not ( n40054 , n40053 );
or ( n217816 , n40018 , n40054 );
xor ( n217817 , n40032 , n40050 );
xnor ( n40057 , n217817 , n40040 );
not ( n217819 , n40057 );
or ( n217820 , n217819 , n209114 );
nand ( n40060 , n217816 , n217820 );
not ( n40061 , n40060 );
buf ( n40062 , n39501 );
not ( n40063 , n40062 );
or ( n40064 , n40061 , n40063 );
not ( n40065 , n40060 );
not ( n40066 , n39501 );
nand ( n40067 , n40065 , n40066 );
nand ( n40068 , n40064 , n40067 );
not ( n40069 , n40068 );
not ( n40070 , n215255 );
xor ( n40071 , n26126 , n26143 );
xnor ( n40072 , n40071 , n39570 );
not ( n217834 , n40072 );
or ( n217835 , n40070 , n217834 );
or ( n40075 , n40072 , n215255 );
nand ( n40076 , n217835 , n40075 );
and ( n40077 , n40076 , n30038 );
not ( n40078 , n40076 );
and ( n40079 , n40078 , n207796 );
nor ( n40080 , n40077 , n40079 );
buf ( n40081 , n37647 );
not ( n40082 , n40081 );
not ( n40083 , n29693 );
or ( n40084 , n40082 , n40083 );
or ( n40085 , n29693 , n40081 );
nand ( n40086 , n40084 , n40085 );
and ( n40087 , n40086 , n207493 );
not ( n40088 , n40086 );
and ( n40089 , n40088 , n39108 );
nor ( n40090 , n40087 , n40089 );
nand ( n40091 , n40080 , n40090 );
not ( n40092 , n40091 );
or ( n40093 , n40069 , n40092 );
or ( n40094 , n40068 , n40091 );
nand ( n40095 , n40093 , n40094 );
not ( n40096 , n40095 );
or ( n40097 , n40017 , n40096 );
or ( n40098 , n40095 , n40016 );
nand ( n40099 , n40097 , n40098 );
buf ( n40100 , n25664 );
not ( n40101 , n37619 );
xor ( n40102 , n40100 , n40101 );
buf ( n40103 , RI173df828_1666);
not ( n40104 , n40103 );
not ( n40105 , RI17396b38_2021);
not ( n40106 , n40105 );
or ( n40107 , n40104 , n40106 );
not ( n40108 , RI173df828_1666);
buf ( n40109 , RI17396b38_2021);
nand ( n40110 , n40108 , n40109 );
nand ( n40111 , n40107 , n40110 );
not ( n40112 , n40111 );
buf ( n40113 , RI19a95750_2644);
nand ( n40114 , n204512 , n40113 );
buf ( n40115 , RI1747be58_1132);
and ( n40116 , n40114 , n40115 );
not ( n40117 , n40114 );
not ( n40118 , RI1747be58_1132);
and ( n40119 , n40117 , n40118 );
nor ( n40120 , n40116 , n40119 );
xor ( n40121 , n37961 , n40120 );
buf ( n40122 , RI19ac5540_2289);
nand ( n217884 , n205020 , n40122 );
not ( n217885 , RI174cba48_777);
and ( n40125 , n217884 , n217885 );
not ( n40126 , n217884 );
buf ( n40127 , RI174cba48_777);
and ( n40128 , n40126 , n40127 );
nor ( n40129 , n40125 , n40128 );
xnor ( n40130 , n40121 , n40129 );
not ( n40131 , n40130 );
not ( n40132 , n40131 );
or ( n40133 , n40112 , n40132 );
not ( n40134 , n40111 );
nand ( n40135 , n40134 , n40130 );
nand ( n40136 , n40133 , n40135 );
xnor ( n40137 , n40102 , n40136 );
not ( n40138 , n40137 );
not ( n40139 , n38166 );
not ( n40140 , n34103 );
or ( n40141 , n40139 , n40140 );
nand ( n40142 , n34089 , n38163 );
nand ( n40143 , n40141 , n40142 );
buf ( n40144 , RI173ef4d0_1589);
not ( n40145 , n40144 );
not ( n40146 , RI173a67e0_1944);
not ( n40147 , n40146 );
or ( n40148 , n40145 , n40147 );
not ( n40149 , RI173ef4d0_1589);
buf ( n40150 , RI173a67e0_1944);
nand ( n40151 , n40149 , n40150 );
nand ( n40152 , n40148 , n40151 );
not ( n40153 , RI1749e598_964);
and ( n40154 , n40152 , n40153 );
not ( n40155 , n40152 );
buf ( n40156 , RI1749e598_964);
and ( n40157 , n40155 , n40156 );
nor ( n40158 , n40154 , n40157 );
xor ( n40159 , n40158 , n38523 );
buf ( n40160 , RI19a9dbf8_2586);
nand ( n40161 , n25622 , n40160 );
buf ( n40162 , RI1748b7b8_1056);
and ( n40163 , n40161 , n40162 );
not ( n40164 , n40161 );
not ( n40165 , RI1748b7b8_1056);
and ( n40166 , n40164 , n40165 );
nor ( n40167 , n40163 , n40166 );
xnor ( n40168 , n40159 , n40167 );
buf ( n40169 , n40168 );
not ( n40170 , n40169 );
and ( n40171 , n40143 , n40170 );
not ( n40172 , n40143 );
and ( n217934 , n40172 , n40169 );
nor ( n217935 , n40171 , n217934 );
nand ( n40175 , n40138 , n217935 );
not ( n40176 , n40175 );
not ( n40177 , n33524 );
not ( n40178 , n40177 );
xor ( n40179 , n32369 , n40178 );
xnor ( n40180 , n40179 , n36189 );
not ( n40181 , n40180 );
and ( n40182 , n40176 , n40181 );
and ( n40183 , n40175 , n40180 );
nor ( n40184 , n40182 , n40183 );
and ( n40185 , n40099 , n40184 );
not ( n40186 , n40099 );
not ( n40187 , n40184 );
and ( n40188 , n40186 , n40187 );
nor ( n40189 , n40185 , n40188 );
and ( n40190 , n217651 , n40189 );
not ( n40191 , n217651 );
not ( n40192 , n40189 );
and ( n40193 , n40191 , n40192 );
nor ( n40194 , n40190 , n40193 );
not ( n40195 , n40194 );
or ( n40196 , n217585 , n40195 );
not ( n40197 , n39823 );
not ( n40198 , n40192 );
not ( n40199 , n217651 );
not ( n40200 , n40199 );
or ( n40201 , n40198 , n40200 );
nand ( n40202 , n217651 , n40189 );
nand ( n40203 , n40201 , n40202 );
nand ( n40204 , n40197 , n40203 );
nand ( n40205 , n40196 , n40204 );
not ( n40206 , n40205 );
buf ( n40207 , n34689 );
not ( n40208 , n40207 );
xor ( n40209 , n204867 , n204874 );
xnor ( n40210 , n40209 , n204889 );
not ( n40211 , n40210 );
or ( n40212 , n40208 , n40211 );
or ( n40213 , n40210 , n40207 );
nand ( n40214 , n40212 , n40213 );
buf ( n40215 , n38201 );
and ( n40216 , n40214 , n40215 );
not ( n40217 , n40214 );
buf ( n40218 , n38188 );
and ( n40219 , n40217 , n40218 );
nor ( n217981 , n40216 , n40219 );
not ( n217982 , n217981 );
xor ( n40222 , n26185 , n26202 );
not ( n40223 , n26193 );
xnor ( n40224 , n40222 , n40223 );
not ( n40225 , n40224 );
not ( n40226 , n36494 );
and ( n40227 , n40225 , n40226 );
and ( n40228 , n40224 , n36494 );
nor ( n40229 , n40227 , n40228 );
buf ( n40230 , n30532 );
buf ( n40231 , n40230 );
and ( n40232 , n40229 , n40231 );
not ( n40233 , n40229 );
not ( n40234 , n40231 );
and ( n40235 , n40233 , n40234 );
nor ( n40236 , n40232 , n40235 );
not ( n40237 , n35702 );
not ( n40238 , n39968 );
or ( n40239 , n40237 , n40238 );
not ( n40240 , n35702 );
nand ( n40241 , n40240 , n39974 );
nand ( n40242 , n40239 , n40241 );
and ( n40243 , n40242 , n40007 );
not ( n40244 , n40242 );
and ( n40245 , n40244 , n40006 );
nor ( n40246 , n40243 , n40245 );
nand ( n40247 , n40236 , n40246 );
not ( n40248 , n40247 );
or ( n40249 , n217982 , n40248 );
or ( n40250 , n40247 , n217981 );
nand ( n40251 , n40249 , n40250 );
not ( n40252 , n40251 );
not ( n40253 , n29426 );
not ( n40254 , n33404 );
or ( n40255 , n40253 , n40254 );
or ( n40256 , n33404 , n29426 );
nand ( n40257 , n40255 , n40256 );
and ( n40258 , n40257 , n34461 );
not ( n40259 , n40257 );
and ( n40260 , n40259 , n34464 );
nor ( n40261 , n40258 , n40260 );
not ( n40262 , n40261 );
not ( n218024 , n38650 );
not ( n218025 , n209146 );
not ( n40265 , n218025 );
or ( n40266 , n218024 , n40265 );
not ( n40267 , n209146 );
or ( n40268 , n40267 , n38650 );
nand ( n40269 , n40266 , n40268 );
not ( n40270 , n31425 );
and ( n40271 , n40269 , n40270 );
not ( n40272 , n40269 );
not ( n40273 , n31428 );
and ( n40274 , n40272 , n40273 );
nor ( n40275 , n40271 , n40274 );
nand ( n40276 , n40262 , n40275 );
not ( n40277 , n40276 );
not ( n40278 , n31612 );
not ( n40279 , n206437 );
or ( n40280 , n40278 , n40279 );
not ( n40281 , n31612 );
nand ( n40282 , n40281 , n37229 );
nand ( n40283 , n40280 , n40282 );
not ( n40284 , n40283 );
not ( n40285 , n205143 );
not ( n40286 , n40285 );
and ( n40287 , n40284 , n40286 );
and ( n40288 , n205142 , n40283 );
nor ( n40289 , n40287 , n40288 );
not ( n40290 , n40289 );
not ( n40291 , n40290 );
and ( n40292 , n40277 , n40291 );
and ( n40293 , n40276 , n40290 );
nor ( n40294 , n40292 , n40293 );
not ( n40295 , n40294 );
or ( n40296 , n40252 , n40295 );
or ( n40297 , n40294 , n40251 );
nand ( n40298 , n40296 , n40297 );
not ( n40299 , n40298 );
not ( n40300 , n40299 );
buf ( n40301 , n36953 );
not ( n40302 , n40301 );
not ( n40303 , n32219 );
not ( n40304 , n40303 );
or ( n40305 , n40302 , n40304 );
or ( n40306 , n40303 , n40301 );
nand ( n40307 , n40305 , n40306 );
and ( n40308 , n40307 , n32236 );
not ( n40309 , n40307 );
and ( n40310 , n40309 , n210002 );
nor ( n40311 , n40308 , n40310 );
not ( n40312 , n38372 );
xor ( n40313 , n37250 , n40312 );
not ( n40314 , n33045 );
xnor ( n40315 , n40313 , n40314 );
not ( n40316 , n40315 );
nand ( n40317 , n40311 , n40316 );
not ( n40318 , n40317 );
not ( n40319 , n208885 );
not ( n40320 , n34177 );
or ( n40321 , n40319 , n40320 );
not ( n40322 , n208885 );
xor ( n218084 , n34159 , n34167 );
xnor ( n218085 , n218084 , n34176 );
nand ( n40325 , n40322 , n218085 );
nand ( n40326 , n40321 , n40325 );
not ( n40327 , n40326 );
not ( n40328 , n34736 );
or ( n40329 , n40327 , n40328 );
or ( n40330 , n34736 , n40326 );
nand ( n40331 , n40329 , n40330 );
not ( n40332 , n40331 );
and ( n40333 , n40318 , n40332 );
and ( n40334 , n40317 , n40331 );
nor ( n40335 , n40333 , n40334 );
not ( n40336 , n40335 );
not ( n40337 , n40336 );
or ( n40338 , n40300 , n40337 );
nand ( n40339 , n40298 , n40335 );
nand ( n40340 , n40338 , n40339 );
and ( n40341 , n28354 , n36349 );
not ( n40342 , n28354 );
and ( n40343 , n40342 , n36350 );
nor ( n40344 , n40341 , n40343 );
not ( n40345 , n205833 );
and ( n40346 , n40344 , n40345 );
not ( n40347 , n40344 );
and ( n40348 , n40347 , n205846 );
nor ( n40349 , n40346 , n40348 );
not ( n40350 , n40349 );
buf ( n40351 , n33785 );
not ( n40352 , n40351 );
not ( n40353 , n38806 );
or ( n40354 , n40352 , n40353 );
or ( n40355 , n38806 , n40351 );
nand ( n40356 , n40354 , n40355 );
and ( n40357 , n40356 , n29088 );
not ( n40358 , n40356 );
not ( n40359 , n29088 );
and ( n40360 , n40358 , n40359 );
nor ( n40361 , n40357 , n40360 );
nand ( n40362 , n40350 , n40361 );
not ( n40363 , n38187 );
not ( n40364 , n34103 );
or ( n40365 , n40363 , n40364 );
not ( n40366 , n38187 );
nand ( n40367 , n40366 , n34089 );
nand ( n40368 , n40365 , n40367 );
not ( n40369 , n40168 );
not ( n40370 , n40369 );
and ( n40371 , n40368 , n40370 );
not ( n40372 , n40368 );
and ( n40373 , n40372 , n40170 );
nor ( n40374 , n40371 , n40373 );
not ( n40375 , n40374 );
and ( n40376 , n40362 , n40375 );
not ( n40377 , n40362 );
and ( n40378 , n40377 , n40374 );
nor ( n40379 , n40376 , n40378 );
not ( n40380 , n40379 );
not ( n40381 , n40380 );
buf ( n40382 , n29852 );
buf ( n40383 , RI173da2d8_1692);
not ( n40384 , n40383 );
not ( n40385 , n29526 );
or ( n218147 , n40384 , n40385 );
not ( n218148 , RI173da2d8_1692);
nand ( n40388 , n218148 , n29484 );
nand ( n40389 , n218147 , n40388 );
not ( n40390 , RI17451db0_1337);
and ( n40391 , n40389 , n40390 );
not ( n40392 , n40389 );
buf ( n40393 , RI17451db0_1337);
and ( n40394 , n40392 , n40393 );
nor ( n40395 , n40391 , n40394 );
buf ( n40396 , RI19ac8c18_2264);
nand ( n40397 , n25711 , n40396 );
buf ( n40398 , RI174c3438_803);
and ( n40399 , n40397 , n40398 );
not ( n40400 , n40397 );
not ( n40401 , RI174c3438_803);
and ( n40402 , n40400 , n40401 );
nor ( n40403 , n40399 , n40402 );
xor ( n40404 , n40395 , n40403 );
buf ( n40405 , RI19a991e8_2618);
nand ( n40406 , n28637 , n40405 );
not ( n40407 , RI174765c0_1159);
and ( n40408 , n40406 , n40407 );
not ( n40409 , n40406 );
buf ( n40410 , RI174765c0_1159);
and ( n40411 , n40409 , n40410 );
nor ( n40412 , n40408 , n40411 );
xnor ( n40413 , n40404 , n40412 );
buf ( n40414 , n40413 );
xor ( n40415 , n40382 , n40414 );
xnor ( n40416 , n40415 , n35940 );
not ( n40417 , n25469 );
buf ( n40418 , n31869 );
not ( n40419 , n40418 );
or ( n40420 , n40417 , n40419 );
or ( n40421 , n37946 , n25469 );
nand ( n40422 , n40420 , n40421 );
and ( n40423 , n40422 , n31907 );
not ( n40424 , n40422 );
not ( n40425 , n31900 );
not ( n40426 , n40425 );
and ( n40427 , n40424 , n40426 );
nor ( n40428 , n40423 , n40427 );
nand ( n40429 , n40416 , n40428 );
not ( n40430 , n40429 );
buf ( n40431 , n30244 );
not ( n40432 , RI1749fc90_957);
and ( n40433 , n40431 , n40432 );
not ( n40434 , n40431 );
and ( n40435 , n40434 , n30241 );
or ( n40436 , n40433 , n40435 );
not ( n40437 , n40436 );
not ( n40438 , n37212 );
or ( n40439 , n40437 , n40438 );
or ( n40440 , n37212 , n40436 );
nand ( n218202 , n40439 , n40440 );
not ( n218203 , n28466 );
and ( n40443 , n218202 , n218203 );
not ( n40444 , n218202 );
and ( n40445 , n40444 , n28466 );
or ( n40446 , n40443 , n40445 );
not ( n40447 , n40446 );
and ( n40448 , n40430 , n40447 );
and ( n40449 , n40429 , n40446 );
nor ( n40450 , n40448 , n40449 );
not ( n40451 , n40450 );
not ( n40452 , n40451 );
or ( n40453 , n40381 , n40452 );
nand ( n40454 , n40450 , n40379 );
nand ( n40455 , n40453 , n40454 );
not ( n40456 , n40455 );
and ( n40457 , n40340 , n40456 );
not ( n40458 , n40340 );
and ( n40459 , n40458 , n40455 );
nor ( n40460 , n40457 , n40459 );
not ( n40461 , n40460 );
and ( n40462 , n40206 , n40461 );
and ( n40463 , n40205 , n40460 );
nor ( n40464 , n40462 , n40463 );
buf ( n40465 , n31571 );
not ( n40466 , n40465 );
nand ( n40467 , n40464 , n40466 );
not ( n40468 , n32134 );
not ( n40469 , n29854 );
or ( n40470 , n40468 , n40469 );
not ( n40471 , n32134 );
nand ( n40472 , n40471 , n29859 );
nand ( n40473 , n40470 , n40472 );
and ( n40474 , n40473 , n33614 );
not ( n40475 , n40473 );
and ( n40476 , n40475 , n33618 );
nor ( n40477 , n40474 , n40476 );
not ( n40478 , n40477 );
not ( n40479 , n40478 );
buf ( n40480 , n35882 );
not ( n40481 , n40480 );
not ( n40482 , n26118 );
not ( n40483 , n32766 );
or ( n40484 , n40482 , n40483 );
nand ( n40485 , n32781 , n26114 );
nand ( n40486 , n40484 , n40485 );
not ( n40487 , n40486 );
or ( n40488 , n40481 , n40487 );
not ( n40489 , n40486 );
nand ( n40490 , n40489 , n39569 );
nand ( n40491 , n40488 , n40490 );
buf ( n40492 , RI173d9c48_1694);
not ( n40493 , n40492 );
not ( n40494 , RI17390f58_2049);
not ( n40495 , n40494 );
or ( n40496 , n40493 , n40495 );
not ( n40497 , RI173d9c48_1694);
nand ( n40498 , n40497 , n34185 );
nand ( n40499 , n40496 , n40498 );
not ( n40500 , RI17451720_1339);
and ( n40501 , n40499 , n40500 );
not ( n40502 , n40499 );
buf ( n40503 , RI17451720_1339);
and ( n40504 , n40502 , n40503 );
nor ( n40505 , n40501 , n40504 );
buf ( n40506 , RI19ac8768_2266);
nand ( n40507 , n26058 , n40506 );
buf ( n40508 , RI174c29e8_805);
and ( n40509 , n40507 , n40508 );
not ( n40510 , n40507 );
not ( n40511 , RI174c29e8_805);
and ( n40512 , n40510 , n40511 );
nor ( n40513 , n40509 , n40512 );
xor ( n40514 , n40505 , n40513 );
buf ( n40515 , RI19a98d38_2620);
nand ( n40516 , n28148 , n40515 );
not ( n40517 , RI17475f30_1161);
and ( n40518 , n40516 , n40517 );
not ( n40519 , n40516 );
buf ( n218281 , RI17475f30_1161);
and ( n218282 , n40519 , n218281 );
nor ( n40522 , n40518 , n218282 );
xnor ( n40523 , n40514 , n40522 );
not ( n40524 , n40523 );
not ( n40525 , n35557 );
and ( n40526 , n40524 , n40525 );
and ( n40527 , n40523 , n35557 );
nor ( n40528 , n40526 , n40527 );
buf ( n40529 , RI173f7180_1551);
not ( n40530 , n40529 );
not ( n40531 , RI173ae490_1906);
not ( n218293 , n40531 );
or ( n218294 , n40530 , n218293 );
not ( n40534 , RI173f7180_1551);
buf ( n40535 , RI173ae490_1906);
nand ( n218297 , n40534 , n40535 );
nand ( n218298 , n218294 , n218297 );
buf ( n40538 , RI17334870_2185);
and ( n218300 , n218298 , n40538 );
not ( n218301 , n218298 );
not ( n40541 , RI17334870_2185);
and ( n40542 , n218301 , n40541 );
nor ( n40543 , n218300 , n40542 );
not ( n40544 , n40543 );
buf ( n40545 , RI19aacbf8_2477);
nand ( n40546 , n25741 , n40545 );
buf ( n40547 , RI174937b0_1017);
and ( n40548 , n40546 , n40547 );
not ( n40549 , n40546 );
not ( n40550 , RI174937b0_1017);
and ( n40551 , n40549 , n40550 );
nor ( n40552 , n40548 , n40551 );
xor ( n40553 , n40544 , n40552 );
buf ( n40554 , RI19ab8778_2392);
nand ( n40555 , n204926 , n40554 );
not ( n40556 , RI175217d0_662);
and ( n40557 , n40555 , n40556 );
not ( n40558 , n40555 );
buf ( n40559 , RI175217d0_662);
and ( n40560 , n40558 , n40559 );
nor ( n40561 , n40557 , n40560 );
xnor ( n40562 , n40553 , n40561 );
not ( n40563 , n40562 );
not ( n40564 , n40563 );
and ( n40565 , n40528 , n40564 );
not ( n40566 , n40528 );
xor ( n40567 , n40543 , n40552 );
xnor ( n40568 , n40567 , n40561 );
buf ( n40569 , n40568 );
and ( n40570 , n40566 , n40569 );
nor ( n40571 , n40565 , n40570 );
not ( n40572 , n40571 );
nand ( n40573 , n40491 , n40572 );
not ( n40574 , n40573 );
or ( n40575 , n40479 , n40574 );
not ( n40576 , n40571 );
nand ( n40577 , n40576 , n40491 );
or ( n40578 , n40577 , n40478 );
nand ( n40579 , n40575 , n40578 );
not ( n40580 , n40579 );
not ( n40581 , n40580 );
nand ( n40582 , n40477 , n40571 );
not ( n40583 , n40582 );
not ( n40584 , n37746 );
buf ( n40585 , n36923 );
not ( n40586 , n40585 );
not ( n40587 , n40586 );
not ( n40588 , n32236 );
or ( n40589 , n40587 , n40588 );
nand ( n218351 , n32240 , n40585 );
nand ( n218352 , n40589 , n218351 );
not ( n40592 , n218352 );
or ( n40593 , n40584 , n40592 );
or ( n40594 , n218352 , n36071 );
nand ( n40595 , n40593 , n40594 );
not ( n40596 , n40595 );
or ( n40597 , n40583 , n40596 );
or ( n40598 , n40595 , n40582 );
nand ( n40599 , n40597 , n40598 );
not ( n40600 , n40599 );
not ( n40601 , n39703 );
not ( n40602 , n30756 );
or ( n40603 , n40601 , n40602 );
not ( n218365 , n39703 );
nand ( n218366 , n218365 , n30769 );
nand ( n40606 , n40603 , n218366 );
not ( n40607 , n39481 );
and ( n40608 , n40606 , n40607 );
not ( n218370 , n40606 );
and ( n218371 , n218370 , n39480 );
nor ( n40611 , n40608 , n218371 );
not ( n40612 , n40611 );
not ( n40613 , n33104 );
not ( n40614 , n37882 );
or ( n40615 , n40613 , n40614 );
not ( n40616 , n33104 );
nand ( n40617 , n40616 , n39019 );
nand ( n40618 , n40615 , n40617 );
not ( n40619 , n37863 );
not ( n40620 , n40619 );
not ( n40621 , n40620 );
and ( n40622 , n40618 , n40621 );
not ( n40623 , n40618 );
and ( n40624 , n40623 , n40620 );
nor ( n40625 , n40622 , n40624 );
not ( n40626 , n40625 );
nand ( n40627 , n40612 , n40626 );
not ( n40628 , n40627 );
not ( n40629 , n209145 );
not ( n40630 , n40052 );
or ( n40631 , n40629 , n40630 );
or ( n40632 , n40057 , n209145 );
nand ( n40633 , n40631 , n40632 );
and ( n40634 , n40633 , n40062 );
not ( n218396 , n40633 );
and ( n218397 , n218396 , n39320 );
or ( n40637 , n40634 , n218397 );
not ( n40638 , n40637 );
not ( n40639 , n40638 );
not ( n40640 , n40639 );
and ( n40641 , n40628 , n40640 );
and ( n218403 , n40627 , n40639 );
nor ( n218404 , n40641 , n218403 );
not ( n218405 , n218404 );
or ( n218406 , n40600 , n218405 );
or ( n40646 , n218404 , n40599 );
nand ( n40647 , n218406 , n40646 );
buf ( n40648 , n40647 );
not ( n40649 , n40648 );
buf ( n40650 , n31115 );
nor ( n40651 , n218085 , n40650 );
not ( n40652 , n40651 );
nand ( n40653 , n218085 , n40650 );
nand ( n40654 , n40652 , n40653 );
not ( n40655 , n40654 );
not ( n40656 , n34736 );
and ( n40657 , n40655 , n40656 );
and ( n40658 , n34736 , n40654 );
nor ( n40659 , n40657 , n40658 );
not ( n40660 , n28405 );
not ( n40661 , n39184 );
not ( n40662 , n26317 );
or ( n40663 , n40661 , n40662 );
nand ( n40664 , n26308 , n216949 );
nand ( n40665 , n40663 , n40664 );
not ( n40666 , n40665 );
or ( n40667 , n40660 , n40666 );
or ( n40668 , n40665 , n28405 );
nand ( n40669 , n40667 , n40668 );
nand ( n218431 , n40659 , n40669 );
not ( n218432 , n36069 );
not ( n40672 , n37352 );
or ( n40673 , n218432 , n40672 );
or ( n40674 , n37352 , n36069 );
nand ( n40675 , n40673 , n40674 );
and ( n40676 , n40675 , n36813 );
not ( n40677 , n40675 );
buf ( n40678 , n39065 );
and ( n40679 , n40677 , n40678 );
nor ( n40680 , n40676 , n40679 );
and ( n40681 , n218431 , n40680 );
not ( n40682 , n218431 );
not ( n40683 , n40680 );
and ( n40684 , n40682 , n40683 );
nor ( n40685 , n40681 , n40684 );
not ( n40686 , n40685 );
not ( n40687 , n40686 );
not ( n40688 , n205426 );
buf ( n40689 , n29288 );
not ( n40690 , n40689 );
not ( n40691 , n33366 );
or ( n40692 , n40690 , n40691 );
or ( n40693 , n33366 , n40689 );
nand ( n40694 , n40692 , n40693 );
not ( n40695 , n40694 );
and ( n40696 , n40688 , n40695 );
not ( n40697 , n205420 );
and ( n40698 , n40697 , n40694 );
nor ( n40699 , n40696 , n40698 );
not ( n40700 , n32962 );
not ( n40701 , n30089 );
buf ( n40702 , RI173f5dd0_1557);
not ( n40703 , n40702 );
not ( n40704 , RI173ad0e0_1912);
not ( n40705 , n40704 );
or ( n40706 , n40703 , n40705 );
not ( n40707 , RI173f5dd0_1557);
nand ( n40708 , n40707 , n26011 );
nand ( n40709 , n40706 , n40708 );
buf ( n40710 , RI17527ef0_642);
and ( n40711 , n40709 , n40710 );
not ( n40712 , n40709 );
not ( n40713 , RI17527ef0_642);
and ( n40714 , n40712 , n40713 );
nor ( n40715 , n40711 , n40714 );
buf ( n40716 , RI19ab0c30_2448);
nand ( n40717 , n25879 , n40716 );
buf ( n40718 , RI1751f8e0_668);
and ( n40719 , n40717 , n40718 );
not ( n40720 , n40717 );
not ( n40721 , RI1751f8e0_668);
and ( n218483 , n40720 , n40721 );
nor ( n218484 , n40719 , n218483 );
xor ( n40724 , n40715 , n218484 );
xnor ( n40725 , n40724 , n39125 );
not ( n40726 , n40725 );
not ( n40727 , n40726 );
or ( n40728 , n40701 , n40727 );
or ( n40729 , n40726 , n30089 );
nand ( n40730 , n40728 , n40729 );
not ( n40731 , n40730 );
or ( n40732 , n40700 , n40731 );
not ( n40733 , n32961 );
not ( n40734 , n40733 );
or ( n40735 , n40730 , n40734 );
nand ( n40736 , n40732 , n40735 );
nand ( n40737 , n40699 , n40736 );
not ( n40738 , n36970 );
not ( n40739 , n28187 );
not ( n40740 , n39642 );
or ( n40741 , n40739 , n40740 );
not ( n40742 , n28187 );
buf ( n40743 , n39641 );
nand ( n40744 , n40742 , n40743 );
nand ( n40745 , n40741 , n40744 );
not ( n40746 , n40745 );
and ( n40747 , n40738 , n40746 );
and ( n40748 , n36970 , n40745 );
nor ( n40749 , n40747 , n40748 );
not ( n218511 , n40749 );
and ( n218512 , n40737 , n218511 );
not ( n40752 , n40737 );
and ( n40753 , n40752 , n40749 );
nor ( n40754 , n218512 , n40753 );
not ( n40755 , n40754 );
not ( n40756 , n40755 );
or ( n40757 , n40687 , n40756 );
nand ( n40758 , n40754 , n40685 );
nand ( n40759 , n40757 , n40758 );
not ( n40760 , n32863 );
not ( n40761 , n28460 );
nor ( n40762 , n40761 , n31343 );
not ( n40763 , n40762 );
not ( n40764 , n28460 );
nand ( n40765 , n40764 , n31343 );
nand ( n40766 , n40763 , n40765 );
not ( n40767 , n40766 );
and ( n40768 , n40760 , n40767 );
and ( n40769 , n32863 , n40766 );
nor ( n40770 , n40768 , n40769 );
not ( n40771 , n38526 );
buf ( n40772 , n33473 );
not ( n40773 , n40772 );
not ( n40774 , n40773 );
or ( n40775 , n40771 , n40774 );
buf ( n40776 , n33474 );
or ( n40777 , n40776 , n38526 );
nand ( n40778 , n40775 , n40777 );
not ( n40779 , RI174a09b0_953);
buf ( n40780 , RI173ef818_1588);
not ( n218542 , n40780 );
not ( n218543 , RI173a6b28_1943);
not ( n40783 , n218543 );
or ( n218545 , n218542 , n40783 );
not ( n218546 , RI173ef818_1588);
buf ( n40786 , RI173a6b28_1943);
nand ( n40787 , n218546 , n40786 );
nand ( n40788 , n218545 , n40787 );
not ( n40789 , n40788 );
xor ( n40790 , n40779 , n40789 );
buf ( n40791 , RI19acc9f8_2234);
nand ( n40792 , n26453 , n40791 );
buf ( n40793 , RI17515908_699);
and ( n40794 , n40792 , n40793 );
not ( n40795 , n40792 );
not ( n40796 , RI17515908_699);
and ( n40797 , n40795 , n40796 );
nor ( n40798 , n40794 , n40797 );
not ( n40799 , n40798 );
buf ( n40800 , RI19a9de50_2585);
nand ( n40801 , n25572 , n40800 );
not ( n40802 , RI1748bb00_1055);
and ( n40803 , n40801 , n40802 );
not ( n40804 , n40801 );
buf ( n40805 , RI1748bb00_1055);
and ( n40806 , n40804 , n40805 );
nor ( n40807 , n40803 , n40806 );
not ( n40808 , n40807 );
or ( n40809 , n40799 , n40808 );
or ( n40810 , n40798 , n40807 );
nand ( n40811 , n40809 , n40810 );
xnor ( n40812 , n40790 , n40811 );
buf ( n40813 , n40812 );
not ( n40814 , n40813 );
and ( n40815 , n40778 , n40814 );
not ( n40816 , n40778 );
and ( n40817 , n40816 , n40813 );
nor ( n40818 , n40815 , n40817 );
nand ( n40819 , n40770 , n40818 );
not ( n40820 , n40819 );
buf ( n40821 , n28904 );
not ( n40822 , RI1749df08_966);
and ( n40823 , n40821 , n40822 );
not ( n40824 , n40821 );
and ( n40825 , n40824 , n28900 );
or ( n40826 , n40823 , n40825 );
not ( n40827 , n40826 );
buf ( n40828 , RI173f3328_1570);
not ( n40829 , n40828 );
not ( n40830 , RI173aa638_1925);
not ( n40831 , n40830 );
or ( n40832 , n40829 , n40831 );
not ( n40833 , RI173f3328_1570);
buf ( n40834 , RI173aa638_1925);
nand ( n218596 , n40833 , n40834 );
nand ( n218597 , n40832 , n218596 );
buf ( n40837 , RI174cc498_775);
and ( n40838 , n218597 , n40837 );
not ( n40839 , n218597 );
not ( n40840 , RI174cc498_775);
and ( n40841 , n40839 , n40840 );
nor ( n40842 , n40838 , n40841 );
buf ( n40843 , RI19aaf088_2461);
nand ( n40844 , n204393 , n40843 );
buf ( n40845 , RI1748f958_1036);
and ( n40846 , n40844 , n40845 );
not ( n40847 , n40844 );
not ( n40848 , RI1748f958_1036);
and ( n40849 , n40847 , n40848 );
nor ( n40850 , n40846 , n40849 );
xor ( n40851 , n40842 , n40850 );
buf ( n40852 , RI19a23a38_2791);
nand ( n40853 , n25540 , n40852 );
buf ( n40854 , RI1751b5d8_681);
and ( n40855 , n40853 , n40854 );
not ( n40856 , n40853 );
not ( n40857 , RI1751b5d8_681);
and ( n40858 , n40856 , n40857 );
nor ( n40859 , n40855 , n40858 );
not ( n40860 , n40859 );
xnor ( n40861 , n40851 , n40860 );
buf ( n40862 , n40861 );
not ( n218624 , n40862 );
or ( n218625 , n40827 , n218624 );
or ( n40865 , n40862 , n40826 );
nand ( n40866 , n218625 , n40865 );
buf ( n40867 , RI173c7b70_1782);
not ( n40868 , n40867 );
not ( n40869 , RI1733e5f0_2137);
not ( n40870 , n40869 );
or ( n40871 , n40868 , n40870 );
not ( n40872 , RI173c7b70_1782);
buf ( n40873 , RI1733e5f0_2137);
nand ( n40874 , n40872 , n40873 );
nand ( n40875 , n40871 , n40874 );
and ( n40876 , n40875 , n38640 );
not ( n40877 , n40875 );
not ( n40878 , RI17410860_1427);
and ( n40879 , n40877 , n40878 );
nor ( n40880 , n40876 , n40879 );
buf ( n40881 , RI19ac1850_2318);
nand ( n40882 , n204493 , n40881 );
buf ( n40883 , RI174ace90_893);
xor ( n40884 , n40882 , n40883 );
xor ( n40885 , n40880 , n40884 );
buf ( n40886 , RI19a915b0_2673);
nand ( n40887 , n28637 , n40886 );
buf ( n40888 , RI174641b8_1248);
and ( n40889 , n40887 , n40888 );
not ( n40890 , n40887 );
not ( n40891 , RI174641b8_1248);
and ( n40892 , n40890 , n40891 );
nor ( n40893 , n40889 , n40892 );
xnor ( n218655 , n40885 , n40893 );
buf ( n218656 , n218655 );
not ( n40896 , n218656 );
and ( n40897 , n40866 , n40896 );
not ( n40898 , n40866 );
and ( n40899 , n40898 , n218656 );
nor ( n40900 , n40897 , n40899 );
not ( n40901 , n40900 );
and ( n40902 , n40820 , n40901 );
and ( n40903 , n40819 , n40900 );
nor ( n40904 , n40902 , n40903 );
buf ( n40905 , n40904 );
and ( n40906 , n40759 , n40905 );
not ( n40907 , n40759 );
not ( n40908 , n40905 );
and ( n40909 , n40907 , n40908 );
nor ( n40910 , n40906 , n40909 );
not ( n40911 , n40910 );
or ( n40912 , n40649 , n40911 );
or ( n40913 , n40910 , n40648 );
nand ( n40914 , n40912 , n40913 );
not ( n40915 , n40914 );
or ( n40916 , n40581 , n40915 );
xor ( n40917 , n40904 , n40759 );
xnor ( n40918 , n40917 , n40647 );
or ( n218680 , n40918 , n40580 );
nand ( n218681 , n40916 , n218680 );
not ( n40921 , n218681 );
xor ( n40922 , n31970 , n206848 );
xor ( n40923 , n40922 , n35740 );
not ( n40924 , n40923 );
not ( n40925 , n35063 );
not ( n40926 , n30976 );
not ( n40927 , n35097 );
or ( n40928 , n40926 , n40927 );
or ( n40929 , n35097 , n30976 );
nand ( n40930 , n40928 , n40929 );
nor ( n40931 , n40925 , n40930 );
not ( n40932 , n40931 );
not ( n40933 , n40930 );
not ( n40934 , n40933 );
not ( n40935 , n35063 );
nand ( n40936 , n40934 , n40935 );
nand ( n40937 , n40932 , n40936 );
not ( n40938 , n40937 );
nand ( n40939 , n40924 , n40938 );
not ( n40940 , n40939 );
not ( n40941 , n32175 );
not ( n40942 , n34200 );
xor ( n40943 , n32121 , n209886 );
xnor ( n40944 , n40943 , n32134 );
not ( n40945 , n40944 );
or ( n40946 , n40942 , n40945 );
or ( n40947 , n40944 , n34200 );
nand ( n40948 , n40946 , n40947 );
not ( n40949 , n40948 );
or ( n40950 , n40941 , n40949 );
or ( n40951 , n40948 , n209942 );
nand ( n40952 , n40950 , n40951 );
not ( n40953 , n40952 );
and ( n40954 , n40940 , n40953 );
and ( n40955 , n40939 , n40952 );
nor ( n40956 , n40954 , n40955 );
not ( n40957 , n40956 );
not ( n40958 , n40957 );
not ( n40959 , n38103 );
not ( n40960 , RI17512578_709);
not ( n40961 , n32669 );
xor ( n40962 , n40960 , n40961 );
xnor ( n40963 , n40962 , n32684 );
not ( n40964 , n40963 );
or ( n40965 , n40959 , n40964 );
or ( n40966 , n40963 , n38103 );
nand ( n40967 , n40965 , n40966 );
not ( n40968 , n40967 );
not ( n40969 , n40136 );
not ( n40970 , n40969 );
and ( n218732 , n40968 , n40970 );
and ( n218733 , n40967 , n40969 );
nor ( n40973 , n218732 , n218733 );
not ( n40974 , n40973 );
not ( n40975 , n40974 );
not ( n40976 , n36969 );
not ( n40977 , n40976 );
not ( n40978 , n28168 );
not ( n40979 , n39642 );
or ( n40980 , n40978 , n40979 );
or ( n40981 , n39642 , n28168 );
nand ( n40982 , n40980 , n40981 );
not ( n40983 , n40982 );
and ( n218745 , n40977 , n40983 );
and ( n218746 , n40976 , n40982 );
nor ( n40986 , n218745 , n218746 );
not ( n218748 , n40986 );
not ( n218749 , n38402 );
buf ( n40989 , RI173cbd10_1762);
not ( n40990 , n40989 );
not ( n40991 , RI17342790_2117);
not ( n40992 , n40991 );
or ( n40993 , n40990 , n40992 );
not ( n40994 , RI173cbd10_1762);
buf ( n40995 , RI17342790_2117);
nand ( n40996 , n40994 , n40995 );
nand ( n40997 , n40993 , n40996 );
not ( n40998 , RI17414d48_1406);
and ( n40999 , n40997 , n40998 );
not ( n41000 , n40997 );
buf ( n41001 , RI17414d48_1406);
and ( n41002 , n41000 , n41001 );
nor ( n41003 , n40999 , n41002 );
buf ( n41004 , RI19a8f3f0_2688);
nand ( n41005 , n26453 , n41004 );
buf ( n41006 , RI17468358_1228);
xor ( n41007 , n41005 , n41006 );
xor ( n41008 , n41003 , n41007 );
buf ( n41009 , RI19abfd98_2333);
nand ( n41010 , n25752 , n41009 );
not ( n41011 , RI174b1030_873);
and ( n41012 , n41010 , n41011 );
not ( n218774 , n41010 );
buf ( n218775 , RI174b1030_873);
and ( n41015 , n218774 , n218775 );
nor ( n41016 , n41012 , n41015 );
xnor ( n41017 , n41008 , n41016 );
not ( n41018 , n41017 );
or ( n41019 , n218749 , n41018 );
or ( n41020 , n41017 , n38402 );
nand ( n41021 , n41019 , n41020 );
not ( n41022 , n41021 );
not ( n41023 , n41022 );
not ( n41024 , n36168 );
not ( n218786 , n41024 );
or ( n218787 , n41023 , n218786 );
nand ( n41027 , n213924 , n41021 );
nand ( n41028 , n218787 , n41027 );
not ( n41029 , n41028 );
nand ( n41030 , n218748 , n41029 );
not ( n41031 , n41030 );
or ( n41032 , n40975 , n41031 );
or ( n41033 , n41030 , n40974 );
nand ( n41034 , n41032 , n41033 );
not ( n41035 , n41034 );
not ( n41036 , n41035 );
or ( n41037 , n40958 , n41036 );
nand ( n41038 , n41034 , n40956 );
nand ( n41039 , n41037 , n41038 );
not ( n41040 , n40523 );
not ( n41041 , n41040 );
xor ( n41042 , n26374 , n41041 );
not ( n41043 , RI174022b0_1497);
not ( n41044 , RI174053e8_1482);
and ( n41045 , n41044 , n37770 );
not ( n41046 , n41044 );
not ( n41047 , RI173bc6f8_1837);
and ( n41048 , n41046 , n41047 );
nor ( n41049 , n41045 , n41048 );
xor ( n41050 , n41043 , n41049 );
buf ( n41051 , RI17333178_2192);
xor ( n41052 , n41051 , n35713 );
xnor ( n41053 , n41052 , n35711 );
xnor ( n41054 , n41050 , n41053 );
buf ( n41055 , n41054 );
xnor ( n41056 , n41042 , n41055 );
not ( n41057 , n34613 );
buf ( n41058 , RI17456c70_1313);
not ( n41059 , n41058 );
not ( n41060 , n33134 );
or ( n41061 , n41059 , n41060 );
not ( n41062 , n33134 );
not ( n41063 , n41062 );
or ( n41064 , n41063 , n41058 );
nand ( n41065 , n41061 , n41064 );
not ( n41066 , n41065 );
or ( n41067 , n41057 , n41066 );
or ( n41068 , n41065 , n214235 );
nand ( n41069 , n41067 , n41068 );
nand ( n41070 , n41056 , n41069 );
buf ( n41071 , n32900 );
not ( n218833 , n41071 );
not ( n218834 , n25984 );
not ( n41074 , n33936 );
or ( n41075 , n218834 , n41074 );
not ( n41076 , n33935 );
not ( n41077 , n41076 );
or ( n41078 , n41077 , n25984 );
nand ( n41079 , n41075 , n41078 );
not ( n41080 , n41079 );
or ( n41081 , n218833 , n41080 );
not ( n41082 , n32903 );
or ( n41083 , n41079 , n41082 );
nand ( n41084 , n41081 , n41083 );
not ( n41085 , n41084 );
and ( n41086 , n41070 , n41085 );
not ( n41087 , n41070 );
and ( n41088 , n41087 , n41084 );
or ( n41089 , n41086 , n41088 );
not ( n41090 , n41089 );
and ( n41091 , n41039 , n41090 );
not ( n41092 , n41039 );
and ( n41093 , n41092 , n41089 );
nor ( n41094 , n41091 , n41093 );
not ( n41095 , n209207 );
not ( n41096 , n207216 );
or ( n41097 , n41095 , n41096 );
nand ( n41098 , n29456 , n31442 );
nand ( n41099 , n41097 , n41098 );
buf ( n41100 , n38690 );
and ( n41101 , n41099 , n41100 );
not ( n41102 , n41099 );
not ( n218864 , n41100 );
and ( n218865 , n41102 , n218864 );
nor ( n41105 , n41101 , n218865 );
not ( n41106 , n41105 );
not ( n41107 , n41106 );
not ( n41108 , n25941 );
not ( n41109 , n32011 );
or ( n41110 , n41108 , n41109 );
nand ( n41111 , n35622 , n25937 );
nand ( n41112 , n41110 , n41111 );
buf ( n41113 , n37940 );
buf ( n41114 , n41113 );
xor ( n41115 , n41112 , n41114 );
not ( n41116 , n30300 );
buf ( n41117 , RI173eb9c0_1607);
not ( n41118 , n41117 );
not ( n41119 , n204269 );
or ( n41120 , n41118 , n41119 );
not ( n41121 , RI173eb9c0_1607);
buf ( n41122 , RI173a2cd0_1962);
nand ( n41123 , n41121 , n41122 );
nand ( n41124 , n41120 , n41123 );
not ( n41125 , RI17477cb8_1152);
and ( n41126 , n41124 , n41125 );
not ( n41127 , n41124 );
buf ( n41128 , RI17477cb8_1152);
and ( n41129 , n41127 , n41128 );
nor ( n41130 , n41126 , n41129 );
buf ( n41131 , RI19a9ff20_2569);
nand ( n41132 , n206902 , n41131 );
not ( n41133 , RI17487ca8_1074);
and ( n218895 , n41132 , n41133 );
not ( n218896 , n41132 );
buf ( n41136 , RI17487ca8_1074);
and ( n41137 , n218896 , n41136 );
nor ( n41138 , n218895 , n41137 );
xor ( n41139 , n41130 , n41138 );
buf ( n41140 , RI19aceac8_2220);
nand ( n41141 , n28238 , n41140 );
not ( n41142 , RI1750f1e8_719);
and ( n41143 , n41141 , n41142 );
not ( n41144 , n41141 );
buf ( n41145 , RI1750f1e8_719);
and ( n41146 , n41144 , n41145 );
nor ( n41147 , n41143 , n41146 );
xnor ( n41148 , n41139 , n41147 );
buf ( n41149 , n41148 );
not ( n41150 , n41149 );
not ( n41151 , n41150 );
or ( n41152 , n41116 , n41151 );
nand ( n41153 , n41149 , n208058 );
nand ( n41154 , n41152 , n41153 );
not ( n41155 , n41154 );
buf ( n218917 , n37116 );
not ( n218918 , n218917 );
not ( n41158 , n218918 );
and ( n41159 , n41155 , n41158 );
and ( n41160 , n41154 , n218918 );
nor ( n41161 , n41159 , n41160 );
not ( n41162 , n41161 );
nand ( n41163 , n41115 , n41162 );
not ( n41164 , n41163 );
or ( n41165 , n41107 , n41164 );
or ( n41166 , n41163 , n41106 );
nand ( n41167 , n41165 , n41166 );
not ( n41168 , n41167 );
not ( n41169 , n26102 );
xor ( n41170 , n31652 , n41169 );
xor ( n41171 , n41170 , n34645 );
not ( n41172 , n41171 );
buf ( n41173 , RI1740c378_1448);
not ( n218935 , n41173 );
not ( n218936 , n33444 );
or ( n41176 , n218935 , n218936 );
not ( n218938 , RI1740c378_1448);
nand ( n218939 , n34597 , n218938 );
nand ( n41179 , n41176 , n218939 );
and ( n41180 , n41179 , n40773 );
not ( n41181 , n41179 );
and ( n41182 , n41181 , n40772 );
nor ( n41183 , n41180 , n41182 );
nand ( n41184 , n41172 , n41183 );
not ( n41185 , n41184 );
not ( n41186 , n38984 );
not ( n41187 , n204976 );
not ( n41188 , n41187 );
or ( n41189 , n41186 , n41188 );
or ( n41190 , n204981 , n38984 );
nand ( n41191 , n41189 , n41190 );
not ( n41192 , n41191 );
not ( n41193 , n206669 );
and ( n41194 , n41192 , n41193 );
buf ( n41195 , n36883 );
and ( n41196 , n41191 , n41195 );
nor ( n41197 , n41194 , n41196 );
not ( n41198 , n41197 );
not ( n41199 , n41198 );
and ( n41200 , n41185 , n41199 );
not ( n41201 , n41183 );
not ( n41202 , n41201 );
nand ( n41203 , n41202 , n41172 );
and ( n41204 , n41203 , n41198 );
nor ( n41205 , n41200 , n41204 );
not ( n41206 , n41205 );
or ( n41207 , n41168 , n41206 );
not ( n41208 , n41167 );
not ( n41209 , n41205 );
nand ( n41210 , n41208 , n41209 );
nand ( n41211 , n41207 , n41210 );
not ( n41212 , n41211 );
and ( n41213 , n41094 , n41212 );
not ( n41214 , n41094 );
and ( n41215 , n41214 , n41211 );
nor ( n41216 , n41213 , n41215 );
buf ( n41217 , n41216 );
not ( n41218 , n41217 );
and ( n41219 , n40921 , n41218 );
not ( n218981 , n41216 );
not ( n218982 , n218981 );
and ( n41222 , n218681 , n218982 );
nor ( n218984 , n41219 , n41222 );
not ( n218985 , n218984 );
not ( n41225 , n205409 );
xor ( n41226 , n35138 , n35146 );
xnor ( n41227 , n41226 , n35155 );
not ( n41228 , n41227 );
or ( n41229 , n41225 , n41228 );
or ( n41230 , n35156 , n205409 );
nand ( n41231 , n41229 , n41230 );
and ( n41232 , n41231 , n36751 );
not ( n41233 , n41231 );
and ( n41234 , n41233 , n37303 );
nor ( n41235 , n41232 , n41234 );
not ( n41236 , n41235 );
buf ( n41237 , RI173cda98_1753);
nand ( n41238 , n218938 , n33409 );
not ( n41239 , RI173c3688_1803);
nand ( n41240 , n41239 , n41173 );
and ( n41241 , n41238 , n41240 );
xor ( n41242 , n41237 , n41241 );
buf ( n41243 , RI19ab11d0_2445);
nand ( n41244 , n28148 , n41243 );
buf ( n41245 , RI174a89a8_914);
and ( n41246 , n41244 , n41245 );
not ( n41247 , n41244 );
not ( n219009 , RI174a89a8_914);
and ( n219010 , n41247 , n219009 );
nor ( n41250 , n41246 , n219010 );
not ( n41251 , n41250 );
buf ( n41252 , RI1733a108_2158);
not ( n41253 , n41252 );
and ( n41254 , n41251 , n41253 );
and ( n41255 , n41250 , n41252 );
nor ( n41256 , n41254 , n41255 );
xor ( n41257 , n41242 , n41256 );
not ( n41258 , n41257 );
not ( n41259 , n41258 );
not ( n219021 , n34587 );
not ( n219022 , RI173a6150_1946);
not ( n41262 , n219022 );
or ( n41263 , n219021 , n41262 );
not ( n41264 , RI173eee40_1591);
buf ( n41265 , RI173a6150_1946);
nand ( n41266 , n41264 , n41265 );
nand ( n41267 , n41263 , n41266 );
not ( n41268 , RI17499d68_986);
and ( n41269 , n41267 , n41268 );
not ( n41270 , n41267 );
and ( n41271 , n41270 , n216868 );
nor ( n41272 , n41269 , n41271 );
buf ( n41273 , RI19acc3e0_2237);
nand ( n41274 , n26453 , n41273 );
not ( n41275 , RI17514990_702);
and ( n41276 , n41274 , n41275 );
not ( n41277 , n41274 );
and ( n41278 , n41277 , n37732 );
nor ( n41279 , n41276 , n41278 );
not ( n41280 , n41279 );
xor ( n41281 , n41272 , n41280 );
buf ( n41282 , RI19a9d658_2588);
nand ( n41283 , n25656 , n41282 );
buf ( n41284 , RI1748b128_1058);
and ( n41285 , n41283 , n41284 );
not ( n41286 , n41283 );
not ( n41287 , RI1748b128_1058);
and ( n41288 , n41286 , n41287 );
nor ( n41289 , n41285 , n41288 );
buf ( n41290 , n41289 );
xnor ( n219052 , n41281 , n41290 );
and ( n219053 , n34015 , n219052 );
not ( n41293 , n34015 );
not ( n41294 , n41289 );
not ( n41295 , n41279 );
or ( n41296 , n41294 , n41295 );
or ( n41297 , n41289 , n41279 );
nand ( n41298 , n41296 , n41297 );
and ( n41299 , n41298 , n41272 );
not ( n41300 , n41298 );
not ( n41301 , n41272 );
and ( n41302 , n41300 , n41301 );
nor ( n41303 , n41299 , n41302 );
and ( n41304 , n41293 , n41303 );
nor ( n41305 , n219053 , n41304 );
not ( n41306 , n41305 );
not ( n41307 , n41306 );
or ( n41308 , n41259 , n41307 );
nand ( n41309 , n41305 , n41257 );
nand ( n41310 , n41308 , n41309 );
not ( n41311 , n41310 );
nand ( n41312 , n41236 , n41311 );
not ( n41313 , n41312 );
buf ( n41314 , n27999 );
not ( n41315 , n41314 );
not ( n41316 , n204504 );
or ( n41317 , n41315 , n41316 );
not ( n41318 , n41314 );
not ( n41319 , n204503 );
nand ( n41320 , n41318 , n41319 );
nand ( n41321 , n41317 , n41320 );
buf ( n41322 , RI173f0bc8_1582);
not ( n219084 , n41322 );
not ( n219085 , RI173a7ed8_1937);
not ( n41325 , n219085 );
or ( n41326 , n219084 , n41325 );
not ( n41327 , RI173f0bc8_1582);
nand ( n41328 , n41327 , n36973 );
nand ( n41329 , n41326 , n41328 );
not ( n41330 , RI174ac170_897);
and ( n41331 , n41329 , n41330 );
not ( n41332 , n41329 );
buf ( n219094 , RI174ac170_897);
and ( n219095 , n41332 , n219094 );
nor ( n41335 , n41331 , n219095 );
buf ( n41336 , RI19a86de0_2746);
nand ( n41337 , n29890 , n41336 );
buf ( n41338 , RI175177f8_693);
and ( n41339 , n41337 , n41338 );
not ( n41340 , n41337 );
not ( n41341 , RI175177f8_693);
and ( n41342 , n41340 , n41341 );
nor ( n41343 , n41339 , n41342 );
xor ( n41344 , n41335 , n41343 );
buf ( n41345 , RI19aafcb8_2455);
nand ( n41346 , n28238 , n41345 );
not ( n41347 , RI1748ceb0_1049);
and ( n219109 , n41346 , n41347 );
not ( n219110 , n41346 );
buf ( n41350 , RI1748ceb0_1049);
and ( n41351 , n219110 , n41350 );
nor ( n219113 , n219109 , n41351 );
xnor ( n41353 , n41344 , n219113 );
not ( n219115 , n41353 );
not ( n219116 , n219115 );
buf ( n41356 , n219116 );
and ( n41357 , n41321 , n41356 );
not ( n41358 , n41321 );
not ( n41359 , n41353 );
not ( n41360 , n41359 );
not ( n41361 , n41360 );
and ( n41362 , n41358 , n41361 );
nor ( n41363 , n41357 , n41362 );
not ( n41364 , n41363 );
not ( n41365 , n41364 );
and ( n41366 , n41313 , n41365 );
and ( n41367 , n41312 , n41364 );
nor ( n41368 , n41366 , n41367 );
buf ( n41369 , n41368 );
not ( n41370 , n41369 );
not ( n41371 , n25507 );
not ( n41372 , n37946 );
or ( n41373 , n41371 , n41372 );
not ( n41374 , n25507 );
not ( n41375 , n40418 );
nand ( n41376 , n41374 , n41375 );
nand ( n41377 , n41373 , n41376 );
and ( n41378 , n41377 , n40426 );
not ( n41379 , n41377 );
and ( n41380 , n41379 , n31907 );
nor ( n41381 , n41378 , n41380 );
buf ( n41382 , RI19a85760_2756);
nand ( n41383 , n25479 , n41382 );
buf ( n41384 , RI17500f80_757);
and ( n41385 , n41383 , n41384 );
not ( n41386 , n41383 );
not ( n41387 , RI17500f80_757);
and ( n41388 , n41386 , n41387 );
nor ( n41389 , n41385 , n41388 );
not ( n41390 , n41389 );
not ( n41391 , n35922 );
or ( n41392 , n41390 , n41391 );
or ( n41393 , n35922 , n41389 );
nand ( n41394 , n41392 , n41393 );
buf ( n41395 , n216493 );
and ( n219157 , n41394 , n41395 );
not ( n219158 , n41394 );
not ( n41398 , n41395 );
and ( n41399 , n219158 , n41398 );
nor ( n41400 , n219157 , n41399 );
not ( n41401 , n41400 );
nand ( n41402 , n41381 , n41401 );
not ( n41403 , n41402 );
not ( n41404 , n41403 );
buf ( n41405 , n30246 );
not ( n41406 , n41405 );
not ( n41407 , n25402 );
and ( n219169 , n41406 , n41407 );
and ( n219170 , n41405 , n25402 );
nor ( n41410 , n219169 , n219170 );
buf ( n41411 , n32572 );
not ( n41412 , n41411 );
and ( n41413 , n41410 , n41412 );
not ( n41414 , n41410 );
not ( n41415 , n41411 );
not ( n41416 , n41415 );
and ( n41417 , n41414 , n41416 );
nor ( n41418 , n41413 , n41417 );
not ( n41419 , n41418 );
not ( n41420 , n41419 );
or ( n41421 , n41404 , n41420 );
nand ( n41422 , n41418 , n41402 );
nand ( n41423 , n41421 , n41422 );
buf ( n41424 , n30493 );
not ( n41425 , n41424 );
not ( n41426 , RI17407b48_1470);
and ( n41427 , n41426 , n25724 );
not ( n41428 , n41426 );
not ( n41429 , RI173bee58_1825);
and ( n41430 , n41428 , n41429 );
nor ( n41431 , n41427 , n41430 );
xor ( n41432 , n32499 , n41431 );
buf ( n41433 , RI19ab5640_2413);
nand ( n41434 , n25451 , n41433 );
not ( n41435 , n41434 );
buf ( n41436 , RI174a3e30_937);
not ( n41437 , n41436 );
and ( n41438 , n41435 , n41437 );
nand ( n219200 , n204393 , n41433 );
and ( n219201 , n219200 , n41436 );
nor ( n41441 , n41438 , n219201 );
not ( n41442 , n41441 );
not ( n41443 , n34321 );
and ( n41444 , n41442 , n41443 );
and ( n41445 , n41441 , n34321 );
nor ( n41446 , n41444 , n41445 );
xnor ( n41447 , n41432 , n41446 );
not ( n41448 , n41447 );
not ( n41449 , n41448 );
not ( n41450 , n41449 );
or ( n41451 , n41425 , n41450 );
not ( n41452 , n41424 );
nand ( n41453 , n41452 , n41448 );
nand ( n219215 , n41451 , n41453 );
and ( n219216 , n219215 , n33229 );
not ( n41456 , n219215 );
and ( n41457 , n41456 , n33230 );
nor ( n219219 , n219216 , n41457 );
buf ( n219220 , n35546 );
not ( n41460 , n219220 );
not ( n41461 , n35543 );
and ( n41462 , n41460 , n41461 );
and ( n41463 , n219220 , n35543 );
nor ( n41464 , n41462 , n41463 );
not ( n41465 , n41464 );
not ( n41466 , n41465 );
not ( n41467 , n40562 );
or ( n41468 , n41466 , n41467 );
nand ( n41469 , n40569 , n41464 );
nand ( n41470 , n41468 , n41469 );
not ( n41471 , n41470 );
not ( n41472 , n29519 );
and ( n41473 , n41471 , n41472 );
and ( n41474 , n41470 , n29519 );
nor ( n41475 , n41473 , n41474 );
nand ( n41476 , n219219 , n41475 );
not ( n41477 , n33423 );
not ( n41478 , n39845 );
or ( n41479 , n41477 , n41478 );
or ( n41480 , n39845 , n33423 );
nand ( n41481 , n41479 , n41480 );
not ( n41482 , n32363 );
and ( n41483 , n41481 , n41482 );
not ( n41484 , n41481 );
and ( n41485 , n41484 , n32363 );
nor ( n41486 , n41483 , n41485 );
not ( n41487 , n41486 );
and ( n41488 , n41476 , n41487 );
not ( n41489 , n41476 );
and ( n41490 , n41489 , n41486 );
nor ( n41491 , n41488 , n41490 );
xnor ( n41492 , n41423 , n41491 );
not ( n41493 , n41492 );
not ( n41494 , n32244 );
not ( n41495 , RI173bd418_1833);
not ( n41496 , n41495 );
or ( n41497 , n41494 , n41496 );
buf ( n41498 , RI173bd418_1833);
nand ( n41499 , n32286 , n41498 );
nand ( n41500 , n41497 , n41499 );
not ( n41501 , n41500 );
not ( n41502 , n41501 );
buf ( n41503 , RI17333e98_2188);
not ( n41504 , RI1740b310_1453);
xor ( n41505 , n41503 , n41504 );
buf ( n41506 , RI174a23f0_945);
not ( n41507 , n41506 );
buf ( n219269 , RI19ab6ae0_2404);
nand ( n219270 , n25850 , n219269 );
not ( n41510 , n219270 );
or ( n41511 , n41507 , n41510 );
nand ( n41512 , n26028 , n219269 );
or ( n41513 , n41512 , n41506 );
nand ( n41514 , n41511 , n41513 );
xnor ( n41515 , n41505 , n41514 );
not ( n41516 , n41515 );
or ( n41517 , n41502 , n41516 );
or ( n41518 , n41515 , n41501 );
nand ( n41519 , n41517 , n41518 );
buf ( n41520 , n41519 );
not ( n41521 , n41520 );
buf ( n41522 , n32164 );
and ( n41523 , n41522 , n33613 );
not ( n41524 , n41522 );
and ( n41525 , n41524 , n33618 );
nor ( n41526 , n41523 , n41525 );
not ( n41527 , n41526 );
and ( n41528 , n41521 , n41527 );
and ( n41529 , n41520 , n41526 );
nor ( n41530 , n41528 , n41529 );
not ( n41531 , n36411 );
not ( n41532 , n205089 );
not ( n41533 , n32607 );
or ( n41534 , n41532 , n41533 );
or ( n41535 , n32607 , n205089 );
nand ( n41536 , n41534 , n41535 );
not ( n41537 , n41536 );
or ( n41538 , n41531 , n41537 );
or ( n41539 , n41536 , n36411 );
nand ( n41540 , n41538 , n41539 );
nand ( n41541 , n41530 , n41540 );
not ( n41542 , n41541 );
not ( n41543 , n33805 );
not ( n41544 , n29046 );
or ( n41545 , n41543 , n41544 );
or ( n41546 , n29046 , n33805 );
nand ( n41547 , n41545 , n41546 );
not ( n41548 , n41547 );
not ( n41549 , n41548 );
not ( n219311 , n29088 );
not ( n219312 , n219311 );
or ( n41552 , n41549 , n219312 );
nand ( n219314 , n29088 , n41547 );
nand ( n219315 , n41552 , n219314 );
not ( n41555 , n219315 );
and ( n41556 , n41542 , n41555 );
and ( n41557 , n41541 , n219315 );
nor ( n41558 , n41556 , n41557 );
not ( n41559 , n41558 );
nand ( n41560 , n41310 , n41363 );
not ( n41561 , n205367 );
not ( n41562 , n31673 );
or ( n41563 , n41561 , n41562 );
or ( n41564 , n209437 , n205367 );
nand ( n41565 , n41563 , n41564 );
and ( n41566 , n41565 , n31637 );
not ( n219328 , n41565 );
buf ( n219329 , n37488 );
and ( n41569 , n219328 , n219329 );
nor ( n41570 , n41566 , n41569 );
and ( n41571 , n41560 , n41570 );
not ( n41572 , n41560 );
not ( n41573 , n41570 );
and ( n41574 , n41572 , n41573 );
nor ( n41575 , n41571 , n41574 );
not ( n41576 , n41575 );
or ( n41577 , n41559 , n41576 );
or ( n41578 , n41575 , n41558 );
nand ( n41579 , n41577 , n41578 );
not ( n41580 , n205480 );
not ( n41581 , n25457 );
or ( n41582 , n41580 , n41581 );
not ( n41583 , n205480 );
nand ( n41584 , n41583 , n36982 );
nand ( n41585 , n41582 , n41584 );
and ( n41586 , n41585 , n25509 );
not ( n41587 , n41585 );
and ( n41588 , n41587 , n25503 );
nor ( n41589 , n41586 , n41588 );
not ( n41590 , n41589 );
xor ( n41591 , n28173 , n205938 );
xnor ( n41592 , n41591 , n28186 );
buf ( n41593 , n41592 );
buf ( n41594 , n41593 );
not ( n219356 , n41594 );
not ( n219357 , n34871 );
not ( n41597 , n34264 );
not ( n219359 , n41597 );
or ( n219360 , n219357 , n219359 );
not ( n41600 , n34871 );
nand ( n41601 , n41600 , n34264 );
nand ( n41602 , n219360 , n41601 );
not ( n41603 , n41602 );
or ( n41604 , n219356 , n41603 );
or ( n41605 , n41602 , n41594 );
nand ( n41606 , n41604 , n41605 );
nand ( n41607 , n41590 , n41606 );
not ( n41608 , n41607 );
not ( n41609 , n29972 );
not ( n41610 , n204790 );
or ( n41611 , n41609 , n41610 );
or ( n41612 , n204790 , n29972 );
nand ( n41613 , n41611 , n41612 );
and ( n41614 , n41613 , n39145 );
not ( n41615 , n41613 );
and ( n41616 , n41615 , n36309 );
nor ( n41617 , n41614 , n41616 );
not ( n41618 , n41617 );
and ( n41619 , n41608 , n41618 );
and ( n41620 , n41607 , n41617 );
nor ( n41621 , n41619 , n41620 );
not ( n41622 , n41621 );
and ( n41623 , n41579 , n41622 );
not ( n41624 , n41579 );
and ( n41625 , n41624 , n41621 );
nor ( n41626 , n41623 , n41625 );
not ( n41627 , n41626 );
or ( n41628 , n41493 , n41627 );
not ( n41629 , n41626 );
not ( n41630 , n41492 );
nand ( n41631 , n41629 , n41630 );
nand ( n41632 , n41628 , n41631 );
not ( n41633 , n41632 );
or ( n41634 , n41370 , n41633 );
not ( n219396 , n41632 );
not ( n219397 , n219396 );
or ( n41637 , n219397 , n41369 );
nand ( n41638 , n41634 , n41637 );
buf ( n41639 , n39631 );
not ( n41640 , n41639 );
not ( n41641 , n28816 );
or ( n41642 , n41640 , n41641 );
or ( n41643 , n28816 , n41639 );
nand ( n41644 , n41642 , n41643 );
not ( n41645 , n41644 );
not ( n41646 , n32219 );
or ( n41647 , n41645 , n41646 );
or ( n41648 , n32219 , n41644 );
nand ( n41649 , n41647 , n41648 );
not ( n41650 , n41649 );
not ( n41651 , n26008 );
not ( n41652 , n40702 );
not ( n41653 , n26046 );
or ( n41654 , n41652 , n41653 );
or ( n41655 , n26046 , n40702 );
nand ( n41656 , n41654 , n41655 );
not ( n41657 , n41656 );
or ( n41658 , n41651 , n41657 );
not ( n41659 , n41656 );
nand ( n41660 , n41659 , n38586 );
nand ( n41661 , n41658 , n41660 );
not ( n41662 , n205289 );
not ( n41663 , n34873 );
or ( n41664 , n41662 , n41663 );
not ( n41665 , n205289 );
nand ( n41666 , n41665 , n36990 );
nand ( n41667 , n41664 , n41666 );
not ( n41668 , n37019 );
buf ( n219430 , n41668 );
and ( n219431 , n41667 , n219430 );
not ( n41671 , n41667 );
and ( n41672 , n41671 , n37023 );
nor ( n41673 , n219431 , n41672 );
nand ( n41674 , n41661 , n41673 );
not ( n41675 , n41674 );
or ( n41676 , n41650 , n41675 );
or ( n41677 , n41674 , n41649 );
nand ( n41678 , n41676 , n41677 );
not ( n41679 , n41678 );
xor ( n41680 , n215255 , n37501 );
xnor ( n41681 , n41680 , n37505 );
xor ( n41682 , n39454 , n41681 );
xnor ( n41683 , n41682 , n39874 );
buf ( n41684 , RI19a8a530_2722);
nand ( n41685 , n29890 , n41684 );
buf ( n41686 , RI1746be68_1210);
and ( n41687 , n41685 , n41686 );
not ( n41688 , n41685 );
not ( n41689 , RI1746be68_1210);
and ( n41690 , n41688 , n41689 );
nor ( n41691 , n41687 , n41690 );
not ( n41692 , n41691 );
buf ( n41693 , RI19abc198_2367);
nand ( n41694 , n29435 , n41693 );
not ( n41695 , RI174b4b40_855);
and ( n219457 , n41694 , n41695 );
not ( n219458 , n41694 );
buf ( n41698 , RI174b4b40_855);
and ( n41699 , n219458 , n41698 );
nor ( n41700 , n219457 , n41699 );
not ( n41701 , n41700 );
or ( n41702 , n41692 , n41701 );
or ( n41703 , n41691 , n41700 );
nand ( n41704 , n41702 , n41703 );
not ( n41705 , n36091 );
not ( n41706 , RI173462a0_2099);
not ( n41707 , n41706 );
or ( n219469 , n41705 , n41707 );
not ( n219470 , RI173cfb68_1743);
buf ( n41710 , RI173462a0_2099);
nand ( n41711 , n219470 , n41710 );
nand ( n41712 , n219469 , n41711 );
not ( n41713 , RI17447658_1388);
and ( n41714 , n41712 , n41713 );
not ( n41715 , n41712 );
buf ( n41716 , RI17447658_1388);
and ( n41717 , n41715 , n41716 );
nor ( n41718 , n41714 , n41717 );
and ( n41719 , n41704 , n41718 );
not ( n219481 , n41704 );
not ( n219482 , n41718 );
and ( n41722 , n219481 , n219482 );
nor ( n41723 , n41719 , n41722 );
not ( n41724 , n41723 );
buf ( n41725 , RI173de478_1672);
not ( n41726 , n41725 );
and ( n41727 , n41724 , n41726 );
and ( n41728 , n41723 , n41725 );
nor ( n41729 , n41727 , n41728 );
buf ( n41730 , RI173ed0b8_1600);
not ( n41731 , n41730 );
not ( n41732 , RI173a43c8_1955);
not ( n41733 , n41732 );
or ( n41734 , n41731 , n41733 );
not ( n41735 , RI173ed0b8_1600);
buf ( n41736 , RI173a43c8_1955);
nand ( n41737 , n41735 , n41736 );
nand ( n41738 , n41734 , n41737 );
and ( n41739 , n41738 , n37813 );
not ( n41740 , n41738 );
not ( n41741 , RI17487960_1075);
and ( n41742 , n41740 , n41741 );
nor ( n41743 , n41739 , n41742 );
buf ( n41744 , RI19a9eaf8_2579);
nand ( n41745 , n25364 , n41744 );
not ( n41746 , RI174893a0_1067);
and ( n41747 , n41745 , n41746 );
not ( n219509 , n41745 );
buf ( n219510 , RI174893a0_1067);
and ( n41750 , n219509 , n219510 );
nor ( n41751 , n41747 , n41750 );
xor ( n41752 , n41743 , n41751 );
xnor ( n41753 , n41752 , n35240 );
not ( n41754 , n41753 );
buf ( n41755 , n41754 );
not ( n41756 , n41755 );
and ( n41757 , n41729 , n41756 );
not ( n41758 , n41729 );
and ( n41759 , n41758 , n41755 );
nor ( n41760 , n41757 , n41759 );
nand ( n41761 , n41683 , n41760 );
not ( n41762 , n41761 );
and ( n41763 , n29111 , n210587 );
not ( n41764 , n29111 );
and ( n41765 , n41764 , n36262 );
nor ( n41766 , n41763 , n41765 );
xor ( n41767 , n41766 , n39401 );
not ( n41768 , n41767 );
not ( n41769 , n41768 );
and ( n41770 , n41762 , n41769 );
and ( n41771 , n41761 , n41768 );
nor ( n41772 , n41770 , n41771 );
not ( n41773 , n41772 );
or ( n41774 , n41679 , n41773 );
or ( n41775 , n41772 , n41678 );
nand ( n219537 , n41774 , n41775 );
not ( n219538 , n36663 );
xor ( n41778 , n25514 , n219538 );
xnor ( n41779 , n41778 , n33886 );
not ( n41780 , n28958 );
not ( n41781 , n30321 );
or ( n41782 , n41780 , n41781 );
or ( n41783 , n28958 , n30320 );
nand ( n41784 , n41782 , n41783 );
not ( n41785 , n37674 );
and ( n41786 , n41784 , n41785 );
not ( n41787 , n41784 );
and ( n41788 , n41787 , n204436 );
nor ( n41789 , n41786 , n41788 );
not ( n41790 , n41789 );
nand ( n41791 , n41779 , n41790 );
not ( n41792 , n41791 );
not ( n41793 , n32363 );
buf ( n41794 , n33433 );
not ( n41795 , n41794 );
xor ( n41796 , n39841 , n39079 );
xnor ( n41797 , n41796 , n38151 );
not ( n41798 , n41797 );
or ( n41799 , n41795 , n41798 );
or ( n41800 , n41797 , n41794 );
nand ( n41801 , n41799 , n41800 );
not ( n41802 , n41801 );
and ( n41803 , n41793 , n41802 );
and ( n41804 , n32363 , n41801 );
nor ( n41805 , n41803 , n41804 );
not ( n41806 , n41805 );
not ( n41807 , n41806 );
and ( n41808 , n41792 , n41807 );
and ( n41809 , n41791 , n41806 );
nor ( n41810 , n41808 , n41809 );
and ( n41811 , n219537 , n41810 );
not ( n41812 , n219537 );
not ( n41813 , n41810 );
and ( n41814 , n41812 , n41813 );
nor ( n41815 , n41811 , n41814 );
not ( n41816 , n41815 );
not ( n41817 , n41816 );
buf ( n41818 , n30878 );
not ( n41819 , n41818 );
not ( n41820 , n36455 );
or ( n41821 , n41819 , n41820 );
not ( n41822 , n41818 );
nand ( n219584 , n41822 , n36456 );
nand ( n219585 , n41821 , n219584 );
and ( n41825 , n219585 , n39212 );
not ( n41826 , n219585 );
and ( n41827 , n41826 , n39211 );
nor ( n41828 , n41825 , n41827 );
not ( n41829 , n41828 );
not ( n41830 , n41829 );
buf ( n41831 , RI173c7828_1783);
not ( n41832 , n41831 );
not ( n219594 , RI1733e2a8_2138);
not ( n219595 , n219594 );
or ( n41835 , n41832 , n219595 );
not ( n41836 , RI173c7828_1783);
buf ( n41837 , RI1733e2a8_2138);
nand ( n41838 , n41836 , n41837 );
nand ( n41839 , n41835 , n41838 );
buf ( n41840 , RI17410518_1428);
and ( n41841 , n41839 , n41840 );
not ( n41842 , n41839 );
not ( n41843 , RI17410518_1428);
and ( n41844 , n41842 , n41843 );
nor ( n41845 , n41841 , n41844 );
buf ( n41846 , RI19a91358_2674);
nand ( n41847 , n25364 , n41846 );
buf ( n41848 , RI17463e70_1249);
and ( n41849 , n41847 , n41848 );
not ( n41850 , n41847 );
not ( n41851 , RI17463e70_1249);
and ( n41852 , n41850 , n41851 );
nor ( n41853 , n41849 , n41852 );
xor ( n41854 , n41845 , n41853 );
xnor ( n41855 , n41854 , n36881 );
not ( n41856 , n41855 );
buf ( n41857 , n41856 );
not ( n41858 , n41857 );
not ( n41859 , n28388 );
not ( n41860 , n39007 );
or ( n219622 , n41859 , n41860 );
not ( n219623 , n39008 );
or ( n41863 , n219623 , n28388 );
nand ( n219625 , n219622 , n41863 );
not ( n219626 , n219625 );
or ( n41866 , n41858 , n219626 );
or ( n41867 , n219625 , n41857 );
nand ( n41868 , n41866 , n41867 );
not ( n41869 , n35940 );
not ( n41870 , n29788 );
not ( n41871 , n35584 );
or ( n41872 , n41870 , n41871 );
not ( n41873 , n29788 );
nand ( n41874 , n41873 , n35590 );
nand ( n41875 , n41872 , n41874 );
not ( n41876 , n41875 );
or ( n41877 , n41869 , n41876 );
buf ( n41878 , n35548 );
or ( n41879 , n41878 , n41875 );
nand ( n41880 , n41877 , n41879 );
not ( n41881 , n41880 );
nand ( n41882 , n41868 , n41881 );
not ( n41883 , n41882 );
or ( n41884 , n41830 , n41883 );
or ( n41885 , n41882 , n41829 );
nand ( n41886 , n41884 , n41885 );
buf ( n41887 , n41886 );
not ( n41888 , n41887 );
buf ( n219650 , n25720 );
xor ( n219651 , n219650 , n30580 );
buf ( n41891 , n30606 );
xnor ( n41892 , n219651 , n41891 );
not ( n41893 , n41892 );
buf ( n41894 , n39811 );
xor ( n41895 , n36315 , n41894 );
xnor ( n41896 , n41895 , n31081 );
not ( n41897 , n41896 );
not ( n41898 , n30908 );
not ( n41899 , n218656 );
or ( n41900 , n41898 , n41899 );
or ( n219662 , n218656 , n30908 );
nand ( n219663 , n41900 , n219662 );
not ( n41903 , n219663 );
buf ( n41904 , n32053 );
not ( n41905 , n41904 );
and ( n41906 , n41903 , n41905 );
and ( n41907 , n219663 , n41904 );
nor ( n41908 , n41906 , n41907 );
nand ( n41909 , n41897 , n41908 );
not ( n41910 , n41909 );
or ( n41911 , n41893 , n41910 );
not ( n41912 , n41908 );
not ( n219674 , n41912 );
nand ( n219675 , n219674 , n41897 );
or ( n41915 , n219675 , n41892 );
nand ( n41916 , n41911 , n41915 );
not ( n41917 , n41916 );
not ( n41918 , n41917 );
or ( n41919 , n41888 , n41918 );
not ( n41920 , n41886 );
nand ( n41921 , n41920 , n41916 );
nand ( n41922 , n41919 , n41921 );
not ( n41923 , n41922 );
not ( n41924 , n41923 );
or ( n41925 , n41817 , n41924 );
not ( n41926 , n41923 );
not ( n41927 , n41816 );
nand ( n41928 , n41926 , n41927 );
nand ( n41929 , n41925 , n41928 );
buf ( n41930 , n41929 );
and ( n41931 , n41638 , n41930 );
not ( n41932 , n41638 );
xor ( n41933 , n41922 , n41815 );
not ( n41934 , n41933 );
not ( n41935 , n41934 );
and ( n41936 , n41932 , n41935 );
nor ( n41937 , n41931 , n41936 );
not ( n41938 , n41937 );
nand ( n41939 , n218985 , n41938 );
or ( n219701 , n40467 , n41939 );
buf ( n219702 , n33252 );
nor ( n41942 , n40464 , n219702 );
nand ( n41943 , n41942 , n41939 );
buf ( n41944 , n31575 );
buf ( n41945 , n41944 );
nand ( n41946 , n41945 , n36941 );
nand ( n41947 , n219701 , n41943 , n41946 );
buf ( n41948 , n41947 );
not ( n41949 , RI19a97820_2629);
or ( n41950 , n25328 , n41949 );
not ( n41951 , RI19a8d8c0_2700);
or ( n41952 , n25336 , n41951 );
nand ( n41953 , n41950 , n41952 );
buf ( n41954 , n41953 );
not ( n219716 , RI19aadfa8_2468);
or ( n219717 , n25328 , n219716 );
not ( n41957 , RI19aa3aa8_2540);
or ( n41958 , n25335 , n41957 );
nand ( n41959 , n219717 , n41958 );
buf ( n41960 , n41959 );
not ( n41961 , n41767 );
buf ( n41962 , n210029 );
not ( n41963 , n41962 );
not ( n41964 , n29561 );
not ( n41965 , n41964 );
or ( n41966 , n41963 , n41965 );
not ( n219728 , n41962 );
nand ( n219729 , n219728 , n29561 );
nand ( n41969 , n41966 , n219729 );
not ( n41970 , n41969 );
not ( n41971 , n215031 );
not ( n41972 , n41971 );
and ( n41973 , n41970 , n41972 );
and ( n41974 , n37261 , n41969 );
nor ( n41975 , n41973 , n41974 );
nand ( n41976 , n41961 , n41975 );
not ( n41977 , n41976 );
not ( n41978 , n27972 );
not ( n41979 , n204504 );
or ( n41980 , n41978 , n41979 );
not ( n41981 , RI17459a60_1299);
nand ( n41982 , n41319 , n41981 );
nand ( n41983 , n41980 , n41982 );
not ( n41984 , n41983 );
not ( n41985 , n41360 );
and ( n41986 , n41984 , n41985 );
and ( n41987 , n41983 , n41356 );
nor ( n41988 , n41986 , n41987 );
not ( n41989 , n41988 );
not ( n41990 , n41989 );
and ( n41991 , n41977 , n41990 );
and ( n41992 , n41976 , n41989 );
nor ( n41993 , n41991 , n41992 );
not ( n41994 , n41993 );
not ( n41995 , n41994 );
not ( n41996 , n41975 );
nand ( n41997 , n41996 , n41988 );
not ( n219759 , n41997 );
not ( n219760 , n41760 );
not ( n42000 , n219760 );
not ( n42001 , n42000 );
and ( n42002 , n219759 , n42001 );
and ( n42003 , n41997 , n42000 );
nor ( n42004 , n42002 , n42003 );
not ( n42005 , n42004 );
buf ( n42006 , n31859 );
not ( n42007 , n42006 );
not ( n42008 , n205350 );
or ( n42009 , n42007 , n42008 );
or ( n42010 , n205350 , n42006 );
nand ( n42011 , n42009 , n42010 );
and ( n42012 , n42011 , n205386 );
not ( n219774 , n42011 );
and ( n219775 , n219774 , n205389 );
nor ( n42015 , n42012 , n219775 );
not ( n42016 , n42015 );
not ( n42017 , n31019 );
not ( n42018 , n28288 );
or ( n42019 , n42017 , n42018 );
not ( n42020 , n31019 );
xor ( n42021 , n206031 , n28287 );
not ( n42022 , n28278 );
xnor ( n42023 , n42021 , n42022 );
nand ( n42024 , n42020 , n42023 );
nand ( n42025 , n42019 , n42024 );
and ( n42026 , n42025 , n34914 );
not ( n42027 , n42025 );
and ( n42028 , n42027 , n34917 );
nor ( n42029 , n42026 , n42028 );
nand ( n42030 , n42016 , n42029 );
not ( n42031 , n41661 );
and ( n42032 , n42030 , n42031 );
not ( n42033 , n42030 );
and ( n42034 , n42033 , n41661 );
nor ( n42035 , n42032 , n42034 );
not ( n42036 , n42035 );
or ( n42037 , n42005 , n42036 );
or ( n42038 , n42035 , n42004 );
nand ( n42039 , n42037 , n42038 );
not ( n42040 , n41779 );
not ( n42041 , n26081 );
not ( n42042 , n32729 );
or ( n42043 , n42041 , n42042 );
nand ( n42044 , n37455 , n26078 );
nand ( n42045 , n42043 , n42044 );
and ( n42046 , n42045 , n39036 );
not ( n42047 , n42045 );
and ( n42048 , n42047 , n32783 );
nor ( n42049 , n42046 , n42048 );
not ( n42050 , n25962 );
not ( n42051 , n32006 );
or ( n42052 , n42050 , n42051 );
not ( n42053 , n25962 );
nand ( n219815 , n42053 , n35622 );
nand ( n219816 , n42052 , n219815 );
not ( n42056 , n219816 );
not ( n42057 , n37940 );
not ( n42058 , n42057 );
not ( n42059 , n42058 );
and ( n42060 , n42056 , n42059 );
and ( n42061 , n219816 , n42058 );
nor ( n219823 , n42060 , n42061 );
not ( n219824 , n219823 );
nand ( n42064 , n42049 , n219824 );
not ( n42065 , n42064 );
and ( n219827 , n42040 , n42065 );
and ( n219828 , n42064 , n41779 );
nor ( n42068 , n219827 , n219828 );
and ( n42069 , n42039 , n42068 );
not ( n42070 , n42039 );
not ( n42071 , n42068 );
and ( n42072 , n42070 , n42071 );
nor ( n42073 , n42069 , n42072 );
not ( n42074 , n41897 );
not ( n42075 , n29386 );
not ( n42076 , n40369 );
or ( n42077 , n42075 , n42076 );
nand ( n42078 , n40169 , n29389 );
nand ( n219840 , n42077 , n42078 );
buf ( n219841 , n33404 );
xor ( n42081 , n219840 , n219841 );
not ( n42082 , n38459 );
not ( n42083 , n42082 );
not ( n42084 , n32176 );
or ( n42085 , n42083 , n42084 );
or ( n42086 , n32176 , n42082 );
nand ( n42087 , n42085 , n42086 );
xor ( n42088 , n41003 , n41007 );
xnor ( n219850 , n42088 , n41016 );
not ( n219851 , n219850 );
not ( n42091 , n219851 );
not ( n42092 , n42091 );
and ( n42093 , n42087 , n42092 );
not ( n42094 , n42087 );
buf ( n42095 , n219850 );
not ( n42096 , n42095 );
not ( n42097 , n42096 );
and ( n42098 , n42094 , n42097 );
nor ( n42099 , n42093 , n42098 );
nand ( n42100 , n42081 , n42099 );
not ( n42101 , n42100 );
and ( n42102 , n42074 , n42101 );
and ( n219864 , n41897 , n42100 );
nor ( n219865 , n42102 , n219864 );
not ( n42105 , n219865 );
not ( n219867 , n42105 );
not ( n219868 , n31637 );
buf ( n42108 , n205373 );
not ( n42109 , n42108 );
not ( n42110 , n31673 );
not ( n42111 , n42110 );
or ( n42112 , n42109 , n42111 );
not ( n42113 , n31672 );
not ( n42114 , n42113 );
or ( n42115 , n42114 , n42108 );
nand ( n42116 , n42112 , n42115 );
not ( n42117 , n42116 );
or ( n42118 , n219868 , n42117 );
or ( n42119 , n42116 , n31637 );
nand ( n219881 , n42118 , n42119 );
not ( n219882 , n219881 );
not ( n42122 , n219882 );
not ( n42123 , n28438 );
not ( n42124 , n31344 );
or ( n42125 , n42123 , n42124 );
or ( n42126 , n31344 , n28438 );
nand ( n42127 , n42125 , n42126 );
not ( n42128 , n42127 );
not ( n219890 , n32863 );
and ( n219891 , n42128 , n219890 );
and ( n42131 , n42127 , n32863 );
nor ( n42132 , n219891 , n42131 );
nand ( n42133 , n42122 , n42132 );
not ( n42134 , n41868 );
and ( n42135 , n42133 , n42134 );
not ( n42136 , n42133 );
not ( n42137 , n42134 );
and ( n42138 , n42136 , n42137 );
nor ( n42139 , n42135 , n42138 );
not ( n42140 , n42139 );
not ( n219902 , n42140 );
or ( n219903 , n219867 , n219902 );
nand ( n42143 , n219865 , n42139 );
nand ( n219905 , n219903 , n42143 );
and ( n219906 , n42073 , n219905 );
not ( n42146 , n42073 );
not ( n42147 , n219905 );
and ( n42148 , n42146 , n42147 );
nor ( n42149 , n219906 , n42148 );
not ( n42150 , n42149 );
or ( n42151 , n41995 , n42150 );
not ( n219913 , n41994 );
and ( n219914 , n42073 , n42147 );
not ( n42154 , n42073 );
and ( n42155 , n42154 , n219905 );
nor ( n42156 , n219914 , n42155 );
nand ( n42157 , n219913 , n42156 );
nand ( n42158 , n42151 , n42157 );
not ( n42159 , n33404 );
not ( n42160 , n42159 );
buf ( n42161 , n29399 );
and ( n42162 , n42161 , n40168 );
not ( n42163 , n42161 );
and ( n42164 , n42163 , n40369 );
or ( n42165 , n42162 , n42164 );
not ( n219927 , n42165 );
not ( n219928 , n219927 );
or ( n42168 , n42160 , n219928 );
nand ( n42169 , n42165 , n33404 );
nand ( n42170 , n42168 , n42169 );
not ( n42171 , n34973 );
not ( n42172 , n204347 );
or ( n42173 , n42171 , n42172 );
not ( n42174 , n204346 );
or ( n42175 , n42174 , n34973 );
nand ( n42176 , n42173 , n42175 );
and ( n42177 , n42176 , n31932 );
not ( n42178 , n42176 );
and ( n42179 , n42178 , n25549 );
nor ( n42180 , n42177 , n42179 );
nor ( n42181 , n42170 , n42180 );
not ( n42182 , n42181 );
not ( n42183 , n29211 );
not ( n42184 , n207960 );
or ( n42185 , n42183 , n42184 );
not ( n42186 , n29211 );
nand ( n42187 , n42186 , n30205 );
nand ( n42188 , n42185 , n42187 );
not ( n42189 , n31832 );
and ( n42190 , n42188 , n42189 );
not ( n42191 , n42188 );
and ( n42192 , n42191 , n31828 );
nor ( n42193 , n42190 , n42192 );
not ( n42194 , n42193 );
not ( n42195 , n42194 );
not ( n42196 , n42195 );
and ( n219958 , n42182 , n42196 );
and ( n219959 , n42181 , n42195 );
nor ( n42199 , n219958 , n219959 );
not ( n42200 , n42199 );
not ( n42201 , n42200 );
nand ( n42202 , n34225 , n40535 );
not ( n42203 , n42202 );
nor ( n42204 , n34225 , n40535 );
nor ( n42205 , n42203 , n42204 );
not ( n42206 , n42205 );
buf ( n42207 , n216225 );
not ( n42208 , n42207 );
or ( n219970 , n42206 , n42208 );
or ( n219971 , n42207 , n42205 );
nand ( n42211 , n219970 , n219971 );
not ( n219973 , n26314 );
not ( n219974 , n38972 );
or ( n42214 , n219973 , n219974 );
not ( n219976 , n38971 );
or ( n219977 , n219976 , n26314 );
nand ( n42217 , n42214 , n219977 );
and ( n219979 , n42217 , n39007 );
not ( n219980 , n42217 );
and ( n42220 , n219980 , n39002 );
nor ( n219982 , n219979 , n42220 );
nand ( n219983 , n42211 , n219982 );
buf ( n42223 , n26091 );
and ( n42224 , n42223 , n37455 );
not ( n42225 , n42223 );
and ( n42226 , n42225 , n32729 );
nor ( n42227 , n42224 , n42226 );
and ( n42228 , n42227 , n32769 );
not ( n42229 , n42227 );
and ( n42230 , n42229 , n32783 );
nor ( n219992 , n42228 , n42230 );
not ( n219993 , n219992 );
and ( n42233 , n219983 , n219993 );
not ( n42234 , n219983 );
and ( n42235 , n42234 , n219992 );
nor ( n42236 , n42233 , n42235 );
not ( n42237 , n42236 );
not ( n42238 , n42237 );
or ( n42239 , n42201 , n42238 );
nand ( n42240 , n42236 , n42199 );
nand ( n42241 , n42239 , n42240 );
not ( n42242 , n205561 );
not ( n220004 , n31254 );
or ( n220005 , n42242 , n220004 );
not ( n42245 , n205561 );
nand ( n42246 , n42245 , n31253 );
nand ( n42247 , n220005 , n42246 );
and ( n42248 , n42247 , n31273 );
not ( n42249 , n42247 );
and ( n42250 , n42249 , n31264 );
nor ( n42251 , n42248 , n42250 );
not ( n42252 , n42251 );
not ( n42253 , n204757 );
not ( n42254 , RI1739c718_1993);
not ( n42255 , n42254 );
or ( n42256 , n42253 , n42255 );
not ( n42257 , RI173e5750_1637);
buf ( n42258 , RI1739c718_1993);
nand ( n42259 , n42257 , n42258 );
nand ( n42260 , n42256 , n42259 );
buf ( n42261 , RI1745d228_1282);
and ( n42262 , n42260 , n42261 );
not ( n42263 , n42260 );
not ( n42264 , RI1745d228_1282);
and ( n42265 , n42263 , n42264 );
nor ( n42266 , n42262 , n42265 );
buf ( n42267 , RI19aa53f8_2528);
nand ( n42268 , n25539 , n42267 );
not ( n42269 , RI17481a38_1104);
and ( n42270 , n42268 , n42269 );
not ( n42271 , n42268 );
buf ( n42272 , RI17481a38_1104);
and ( n42273 , n42271 , n42272 );
nor ( n220035 , n42270 , n42273 );
xor ( n220036 , n42266 , n220035 );
buf ( n42276 , RI19a86750_2749);
nand ( n42277 , n29435 , n42276 );
not ( n42278 , RI175038c0_749);
and ( n42279 , n42277 , n42278 );
not ( n42280 , n42277 );
buf ( n42281 , RI175038c0_749);
and ( n42282 , n42280 , n42281 );
nor ( n42283 , n42279 , n42282 );
xnor ( n42284 , n220036 , n42283 );
buf ( n42285 , n42284 );
not ( n220047 , n42285 );
not ( n220048 , n31186 );
not ( n42288 , n31428 );
or ( n42289 , n220048 , n42288 );
or ( n42290 , n40270 , n31186 );
nand ( n42291 , n42289 , n42290 );
not ( n42292 , n42291 );
or ( n42293 , n220047 , n42292 );
or ( n42294 , n42291 , n42285 );
nand ( n42295 , n42293 , n42294 );
nand ( n42296 , n42252 , n42295 );
not ( n42297 , n42296 );
buf ( n42298 , n41514 );
not ( n42299 , n42298 );
not ( n42300 , n210044 );
not ( n42301 , n42300 );
or ( n42302 , n42299 , n42301 );
not ( n42303 , n42300 );
not ( n42304 , n42298 );
nand ( n42305 , n42303 , n42304 );
nand ( n42306 , n42302 , n42305 );
and ( n42307 , n42306 , n32323 );
not ( n42308 , n42306 );
and ( n42309 , n42308 , n32326 );
nor ( n42310 , n42307 , n42309 );
not ( n42311 , n42310 );
not ( n42312 , n42311 );
and ( n220074 , n42297 , n42312 );
and ( n220075 , n42296 , n42311 );
nor ( n42315 , n220074 , n220075 );
and ( n42316 , n42241 , n42315 );
not ( n42317 , n42241 );
not ( n42318 , n42315 );
and ( n42319 , n42317 , n42318 );
nor ( n42320 , n42316 , n42319 );
not ( n42321 , n42320 );
not ( n42322 , n42321 );
not ( n42323 , n40976 );
not ( n42324 , n205926 );
not ( n42325 , n40743 );
not ( n42326 , n42325 );
or ( n42327 , n42324 , n42326 );
or ( n220089 , n42325 , n205926 );
nand ( n220090 , n42327 , n220089 );
not ( n42330 , n220090 );
and ( n42331 , n42323 , n42330 );
and ( n42332 , n36970 , n220090 );
nor ( n42333 , n42331 , n42332 );
not ( n42334 , n42333 );
buf ( n42335 , RI19ac46b8_2296);
nand ( n42336 , n25915 , n42335 );
buf ( n42337 , RI174c9b58_783);
and ( n42338 , n42336 , n42337 );
not ( n42339 , n42336 );
not ( n42340 , RI174c9b58_783);
and ( n42341 , n42339 , n42340 );
nor ( n42342 , n42338 , n42341 );
not ( n42343 , n42342 );
not ( n42344 , n42343 );
not ( n42345 , n42344 );
not ( n42346 , n41691 );
xor ( n42347 , n41718 , n42346 );
xnor ( n42348 , n42347 , n41700 );
not ( n42349 , n42348 );
or ( n42350 , n42345 , n42349 );
or ( n42351 , n42348 , n42344 );
nand ( n42352 , n42350 , n42351 );
and ( n220114 , n42352 , n41756 );
not ( n220115 , n42352 );
not ( n42355 , n41754 );
not ( n42356 , n42355 );
and ( n42357 , n220115 , n42356 );
nor ( n42358 , n220114 , n42357 );
buf ( n42359 , n42358 );
nand ( n42360 , n42334 , n42359 );
buf ( n42361 , n31662 );
not ( n42362 , n42361 );
buf ( n42363 , RI173cdde0_1752);
not ( n42364 , n34635 );
xor ( n220126 , n42363 , n42364 );
xnor ( n220127 , n220126 , n34642 );
not ( n42367 , n220127 );
not ( n42368 , n42367 );
or ( n42369 , n42362 , n42368 );
or ( n42370 , n42367 , n42361 );
nand ( n42371 , n42369 , n42370 );
buf ( n42372 , n26102 );
and ( n42373 , n42371 , n42372 );
not ( n42374 , n42371 );
not ( n42375 , n42372 );
and ( n42376 , n42374 , n42375 );
nor ( n42377 , n42373 , n42376 );
and ( n42378 , n42360 , n42377 );
not ( n42379 , n42360 );
not ( n42380 , n42377 );
and ( n42381 , n42379 , n42380 );
nor ( n42382 , n42378 , n42381 );
not ( n42383 , n42382 );
not ( n220145 , n42383 );
not ( n220146 , n30002 );
not ( n42386 , n35888 );
or ( n42387 , n220146 , n42386 );
not ( n42388 , n30002 );
nand ( n42389 , n42388 , n35882 );
nand ( n42390 , n42387 , n42389 );
not ( n42391 , n35926 );
and ( n220153 , n42390 , n42391 );
not ( n220154 , n42390 );
not ( n42394 , n35923 );
and ( n220156 , n220154 , n42394 );
nor ( n220157 , n220153 , n220156 );
buf ( n42397 , n32962 );
not ( n42398 , n42397 );
not ( n42399 , n30093 );
not ( n42400 , n40726 );
not ( n42401 , n42400 );
or ( n42402 , n42399 , n42401 );
not ( n42403 , n30093 );
nand ( n42404 , n42403 , n40726 );
nand ( n220166 , n42402 , n42404 );
not ( n220167 , n220166 );
or ( n42407 , n42398 , n220167 );
or ( n42408 , n220166 , n42397 );
nand ( n42409 , n42407 , n42408 );
nor ( n42410 , n220157 , n42409 );
not ( n42411 , n33031 );
not ( n42412 , n42411 );
not ( n42413 , n213924 );
or ( n42414 , n42412 , n42413 );
or ( n42415 , n36168 , n42411 );
nand ( n42416 , n42414 , n42415 );
and ( n220178 , n42416 , n36189 );
not ( n220179 , n42416 );
and ( n42419 , n220179 , n36190 );
nor ( n42420 , n220178 , n42419 );
not ( n42421 , n42420 );
not ( n42422 , n42421 );
and ( n42423 , n42410 , n42422 );
not ( n42424 , n42410 );
and ( n220186 , n42424 , n42421 );
nor ( n220187 , n42423 , n220186 );
not ( n42427 , n220187 );
not ( n42428 , n42427 );
or ( n42429 , n220145 , n42428 );
nand ( n42430 , n220187 , n42382 );
nand ( n42431 , n42429 , n42430 );
not ( n42432 , n42431 );
not ( n42433 , n42432 );
or ( n42434 , n42322 , n42433 );
nand ( n42435 , n42320 , n42431 );
nand ( n42436 , n42434 , n42435 );
buf ( n220198 , n42436 );
and ( n220199 , n42158 , n220198 );
not ( n42439 , n42158 );
not ( n220201 , n220198 );
and ( n220202 , n42439 , n220201 );
nor ( n42442 , n220199 , n220202 );
not ( n42443 , n205649 );
nor ( n42444 , n42442 , n42443 );
not ( n42445 , n204844 );
not ( n42446 , n28877 );
or ( n42447 , n42445 , n42446 );
or ( n42448 , n28877 , n204844 );
nand ( n42449 , n42447 , n42448 );
and ( n42450 , n42449 , n37472 );
not ( n42451 , n42449 );
and ( n220213 , n42451 , n37469 );
nor ( n220214 , n42450 , n220213 );
not ( n42454 , n220214 );
nand ( n42455 , n41198 , n42454 );
not ( n42456 , n42455 );
buf ( n42457 , RI19a94b98_2649);
nand ( n42458 , n205124 , n42457 );
buf ( n42459 , RI1747b480_1135);
and ( n42460 , n42458 , n42459 );
not ( n42461 , n42458 );
not ( n42462 , RI1747b480_1135);
and ( n42463 , n42461 , n42462 );
nor ( n220225 , n42460 , n42463 );
not ( n220226 , n220225 );
not ( n42466 , n220226 );
not ( n42467 , n34564 );
or ( n42468 , n42466 , n42467 );
not ( n42469 , n220226 );
nand ( n42470 , n42469 , n34558 );
nand ( n42471 , n42468 , n42470 );
buf ( n42472 , n32652 );
not ( n42473 , n42472 );
and ( n42474 , n42471 , n42473 );
not ( n42475 , n42471 );
and ( n220237 , n42475 , n42472 );
nor ( n220238 , n42474 , n220237 );
not ( n42478 , n220238 );
and ( n42479 , n42456 , n42478 );
and ( n42480 , n42455 , n220238 );
nor ( n42481 , n42479 , n42480 );
not ( n42482 , n42481 );
not ( n42483 , n42482 );
not ( n42484 , n41069 );
not ( n42485 , n37347 );
buf ( n42486 , n32196 );
not ( n42487 , n42486 );
not ( n220249 , n42487 );
not ( n220250 , n41725 );
not ( n42490 , RI17395788_2027);
not ( n42491 , n42490 );
or ( n42492 , n220250 , n42491 );
not ( n42493 , RI173de478_1672);
buf ( n42494 , RI17395788_2027);
nand ( n42495 , n42493 , n42494 );
nand ( n42496 , n42492 , n42495 );
not ( n42497 , RI17455f50_1317);
and ( n42498 , n42496 , n42497 );
not ( n42499 , n42496 );
buf ( n42500 , RI17455f50_1317);
and ( n42501 , n42499 , n42500 );
nor ( n42502 , n42498 , n42501 );
buf ( n42503 , RI19a94490_2652);
nand ( n42504 , n26266 , n42503 );
buf ( n42505 , RI1747aaa8_1138);
and ( n42506 , n42504 , n42505 );
not ( n42507 , n42504 );
not ( n42508 , RI1747aaa8_1138);
and ( n42509 , n42507 , n42508 );
nor ( n42510 , n42506 , n42509 );
xor ( n42511 , n42502 , n42510 );
xnor ( n42512 , n42511 , n42343 );
not ( n220274 , n42512 );
or ( n220275 , n220249 , n220274 );
xor ( n42515 , n42502 , n42342 );
buf ( n220277 , n42510 );
xnor ( n220278 , n42515 , n220277 );
nand ( n42518 , n220278 , n42486 );
nand ( n42519 , n220275 , n42518 );
not ( n42520 , n42519 );
or ( n42521 , n42485 , n42520 );
or ( n42522 , n42519 , n37347 );
nand ( n42523 , n42521 , n42522 );
not ( n42524 , n42523 );
not ( n42525 , n29015 );
buf ( n42526 , n35146 );
not ( n42527 , n42526 );
not ( n220289 , n29006 );
or ( n220290 , n42527 , n220289 );
or ( n42530 , n29006 , n42526 );
nand ( n42531 , n220290 , n42530 );
not ( n42532 , n42531 );
not ( n42533 , n42532 );
or ( n42534 , n42525 , n42533 );
nand ( n42535 , n206777 , n42531 );
nand ( n42536 , n42534 , n42535 );
nand ( n42537 , n42524 , n42536 );
not ( n42538 , n42537 );
or ( n42539 , n42484 , n42538 );
not ( n42540 , n42523 );
nand ( n42541 , n42540 , n42536 );
or ( n42542 , n42541 , n41069 );
nand ( n42543 , n42539 , n42542 );
not ( n42544 , n42543 );
not ( n42545 , n32082 );
buf ( n42546 , n205028 );
and ( n42547 , n42546 , n216262 );
not ( n42548 , n42546 );
and ( n42549 , n42548 , n32049 );
nor ( n42550 , n42547 , n42549 );
not ( n42551 , n42550 );
and ( n42552 , n42545 , n42551 );
and ( n42553 , n32082 , n42550 );
nor ( n42554 , n42552 , n42553 );
not ( n42555 , n30034 );
not ( n42556 , n37503 );
not ( n42557 , n40072 );
or ( n42558 , n42556 , n42557 );
or ( n220320 , n26145 , n37503 );
nand ( n220321 , n42558 , n220320 );
not ( n42561 , n220321 );
or ( n42562 , n42555 , n42561 );
or ( n42563 , n220321 , n30038 );
nand ( n42564 , n42562 , n42563 );
nand ( n42565 , n42554 , n42564 );
not ( n42566 , n42565 );
not ( n220328 , n218748 );
and ( n220329 , n42566 , n220328 );
and ( n42569 , n42565 , n218748 );
nor ( n220331 , n220329 , n42569 );
not ( n220332 , n220331 );
or ( n42572 , n42544 , n220332 );
or ( n42573 , n220331 , n42543 );
nand ( n42574 , n42572 , n42573 );
not ( n42575 , n36838 );
buf ( n42576 , RI1748e5a8_1042);
not ( n42577 , n34482 );
not ( n42578 , RI173c1900_1812);
not ( n42579 , n42578 );
or ( n42580 , n42577 , n42579 );
not ( n42581 , RI1740a5f0_1457);
buf ( n220343 , RI173c1900_1812);
nand ( n220344 , n42581 , n220343 );
nand ( n42584 , n42580 , n220344 );
xor ( n220346 , n42576 , n42584 );
buf ( n220347 , RI17338380_2167);
not ( n42587 , RI174a6c20_923);
xor ( n42588 , n220347 , n42587 );
buf ( n42589 , RI19ab2670_2436);
nand ( n42590 , n204926 , n42589 );
xnor ( n42591 , n42588 , n42590 );
xnor ( n42592 , n220346 , n42591 );
not ( n42593 , n42592 );
not ( n42594 , n42593 );
or ( n42595 , n42575 , n42594 );
or ( n42596 , n42593 , n36838 );
nand ( n42597 , n42595 , n42596 );
buf ( n42598 , RI173dee50_1669);
not ( n42599 , n42598 );
not ( n42600 , RI17396160_2024);
not ( n42601 , n42600 );
or ( n42602 , n42599 , n42601 );
not ( n42603 , RI173dee50_1669);
buf ( n42604 , RI17396160_2024);
nand ( n42605 , n42603 , n42604 );
nand ( n42606 , n42602 , n42605 );
not ( n42607 , RI17456928_1314);
and ( n42608 , n42606 , n42607 );
not ( n42609 , n42606 );
buf ( n42610 , RI17456928_1314);
and ( n42611 , n42609 , n42610 );
nor ( n42612 , n42608 , n42611 );
xor ( n42613 , n42612 , n220225 );
buf ( n42614 , RI19ac4dc0_2293);
nand ( n42615 , n26398 , n42614 );
buf ( n42616 , RI174caad0_780);
and ( n42617 , n42615 , n42616 );
not ( n42618 , n42615 );
not ( n42619 , RI174caad0_780);
and ( n42620 , n42618 , n42619 );
nor ( n42621 , n42617 , n42620 );
not ( n42622 , n42621 );
xnor ( n42623 , n42613 , n42622 );
not ( n42624 , n42623 );
and ( n42625 , n42597 , n42624 );
not ( n42626 , n42597 );
buf ( n42627 , n42623 );
and ( n42628 , n42626 , n42627 );
nor ( n42629 , n42625 , n42628 );
not ( n42630 , n42629 );
buf ( n42631 , n40403 );
not ( n42632 , n42631 );
not ( n42633 , n207285 );
or ( n42634 , n42632 , n42633 );
or ( n42635 , n207285 , n42631 );
nand ( n42636 , n42634 , n42635 );
and ( n42637 , n42636 , n29563 );
not ( n42638 , n42636 );
not ( n220400 , n41964 );
and ( n220401 , n42638 , n220400 );
nor ( n42641 , n42637 , n220401 );
not ( n42642 , n42641 );
nand ( n42643 , n42630 , n42642 );
xor ( n42644 , n42643 , n40923 );
xor ( n42645 , n42574 , n42644 );
not ( n42646 , n220214 );
nor ( n42647 , n42646 , n220238 );
and ( n42648 , n42647 , n41171 );
not ( n42649 , n42647 );
and ( n42650 , n42649 , n41172 );
nor ( n220412 , n42648 , n42650 );
not ( n220413 , n220412 );
not ( n42653 , n220413 );
not ( n42654 , n33303 );
not ( n42655 , n205142 );
buf ( n42656 , n213608 );
nor ( n42657 , n42655 , n42656 );
not ( n42658 , n42657 );
nand ( n220420 , n42656 , n205143 );
nand ( n220421 , n42658 , n220420 );
not ( n42661 , n220421 );
or ( n220423 , n42654 , n42661 );
or ( n220424 , n220421 , n33300 );
nand ( n42664 , n220423 , n220424 );
buf ( n42665 , RI1749e250_965);
and ( n42666 , n38654 , n42665 );
not ( n42667 , n38654 );
and ( n42668 , n42667 , n38651 );
nor ( n42669 , n42666 , n42668 );
not ( n42670 , n42669 );
not ( n220432 , n40267 );
not ( n220433 , n220432 );
or ( n220434 , n42670 , n220433 );
buf ( n220435 , n218025 );
not ( n42675 , n220435 );
or ( n42676 , n42675 , n42669 );
nand ( n42677 , n220434 , n42676 );
and ( n42678 , n42677 , n40273 );
not ( n42679 , n42677 );
not ( n42680 , n40270 );
not ( n42681 , n42680 );
and ( n42682 , n42679 , n42681 );
nor ( n42683 , n42678 , n42682 );
not ( n42684 , n42683 );
nand ( n42685 , n42664 , n42684 );
and ( n220447 , n42685 , n41161 );
not ( n220448 , n42685 );
and ( n42688 , n220448 , n41162 );
nor ( n42689 , n220447 , n42688 );
not ( n42690 , n42689 );
not ( n42691 , n42690 );
or ( n42692 , n42653 , n42691 );
nand ( n42693 , n42689 , n220412 );
nand ( n42694 , n42692 , n42693 );
not ( n220456 , n42694 );
and ( n220457 , n42645 , n220456 );
not ( n42697 , n42645 );
and ( n220459 , n42697 , n42694 );
nor ( n220460 , n220457 , n220459 );
not ( n42700 , n220460 );
or ( n42701 , n42483 , n42700 );
not ( n42702 , n42482 );
and ( n42703 , n42645 , n42694 );
not ( n42704 , n42645 );
and ( n42705 , n42704 , n220456 );
nor ( n220467 , n42703 , n42705 );
nand ( n220468 , n42702 , n220467 );
nand ( n42708 , n42701 , n220468 );
buf ( n42709 , n38424 );
not ( n220471 , n42709 );
not ( n220472 , n219851 );
or ( n42712 , n220471 , n220472 );
or ( n42713 , n219851 , n42709 );
nand ( n42714 , n42712 , n42713 );
not ( n42715 , n42714 );
not ( n42716 , n42715 );
not ( n42717 , n41024 );
or ( n42718 , n42716 , n42717 );
nand ( n220480 , n36168 , n42714 );
nand ( n220481 , n42718 , n220480 );
not ( n42721 , n220481 );
not ( n42722 , n33586 );
not ( n42723 , n40414 );
or ( n42724 , n42722 , n42723 );
or ( n42725 , n40414 , n33586 );
nand ( n42726 , n42724 , n42725 );
and ( n42727 , n42726 , n32280 );
not ( n42728 , n42726 );
and ( n42729 , n42728 , n42303 );
nor ( n42730 , n42727 , n42729 );
not ( n220492 , n204638 );
buf ( n220493 , RI1739acd8_2001);
not ( n42733 , n220493 );
not ( n42734 , RI173e39c8_1646);
not ( n42735 , n42734 );
or ( n42736 , n42733 , n42735 );
not ( n42737 , RI1739acd8_2001);
buf ( n42738 , RI173e39c8_1646);
nand ( n42739 , n42737 , n42738 );
nand ( n42740 , n42736 , n42739 );
not ( n42741 , RI1745b7e8_1290);
and ( n42742 , n42740 , n42741 );
not ( n220504 , n42740 );
buf ( n220505 , RI1745b7e8_1290);
and ( n42745 , n220504 , n220505 );
nor ( n42746 , n42742 , n42745 );
xor ( n42747 , n42746 , n41389 );
buf ( n42748 , RI19aa44f8_2535);
nand ( n42749 , n27749 , n42748 );
buf ( n42750 , RI1747fff8_1112);
and ( n42751 , n42749 , n42750 );
not ( n42752 , n42749 );
not ( n42753 , RI1747fff8_1112);
and ( n42754 , n42752 , n42753 );
nor ( n42755 , n42751 , n42754 );
xnor ( n42756 , n42747 , n42755 );
not ( n220518 , n42756 );
not ( n220519 , n220518 );
or ( n42759 , n220492 , n220519 );
not ( n42760 , n42756 );
or ( n42761 , n42760 , n204638 );
nand ( n42762 , n42759 , n42761 );
not ( n42763 , n42762 );
buf ( n42764 , RI173b8558_1857);
not ( n42765 , n42764 );
not ( n42766 , RI17401248_1502);
not ( n220528 , n42766 );
or ( n220529 , n42765 , n220528 );
not ( n42769 , RI173b8558_1857);
buf ( n220531 , RI17401248_1502);
nand ( n220532 , n42769 , n220531 );
nand ( n42772 , n220529 , n220532 );
xor ( n220534 , n38728 , n42772 );
buf ( n220535 , RI1749d530_969);
xor ( n42775 , n38265 , n220535 );
buf ( n42776 , RI19ab8430_2393);
nand ( n42777 , n29597 , n42776 );
xnor ( n42778 , n42775 , n42777 );
xnor ( n42779 , n220534 , n42778 );
not ( n42780 , n42779 );
or ( n220542 , n42763 , n42780 );
buf ( n220543 , n42779 );
or ( n42783 , n220543 , n42762 );
nand ( n220545 , n220542 , n42783 );
nand ( n220546 , n42730 , n220545 );
not ( n42786 , n220546 );
or ( n42787 , n42721 , n42786 );
buf ( n42788 , n220545 );
nand ( n42789 , n42730 , n42788 );
or ( n42790 , n220481 , n42789 );
nand ( n42791 , n42787 , n42790 );
not ( n42792 , n42791 );
and ( n42793 , n37982 , n208398 );
not ( n42794 , n37982 );
not ( n42795 , RI17332110_2197);
xor ( n220557 , n42795 , n208382 );
xnor ( n220558 , n220557 , n30636 );
and ( n42798 , n42794 , n220558 );
nor ( n220560 , n42793 , n42798 );
and ( n220561 , n220560 , n34179 );
not ( n42801 , n220560 );
buf ( n42802 , n218085 );
and ( n42803 , n42801 , n42802 );
nor ( n42804 , n220561 , n42803 );
not ( n42805 , n38328 );
not ( n42806 , n37900 );
not ( n220568 , n42806 );
or ( n220569 , n42805 , n220568 );
or ( n42809 , n42806 , n38328 );
nand ( n42810 , n220569 , n42809 );
and ( n42811 , n42810 , n37397 );
not ( n42812 , n42810 );
not ( n220574 , n37398 );
and ( n220575 , n42812 , n220574 );
nor ( n42815 , n42811 , n220575 );
not ( n220577 , n42815 );
nand ( n220578 , n42804 , n220577 );
not ( n42818 , n30853 );
not ( n42819 , n35876 );
not ( n42820 , n31008 );
or ( n42821 , n42819 , n42820 );
not ( n42822 , n35876 );
nand ( n42823 , n42822 , n35753 );
nand ( n42824 , n42821 , n42823 );
not ( n42825 , n42824 );
or ( n42826 , n42818 , n42825 );
or ( n42827 , n42824 , n30853 );
nand ( n220589 , n42826 , n42827 );
and ( n220590 , n220578 , n220589 );
not ( n42830 , n220578 );
not ( n42831 , n220589 );
and ( n42832 , n42830 , n42831 );
nor ( n42833 , n220590 , n42832 );
not ( n42834 , n42833 );
or ( n42835 , n42792 , n42834 );
not ( n42836 , n42791 );
not ( n42837 , n42833 );
nand ( n42838 , n42836 , n42837 );
nand ( n42839 , n42835 , n42838 );
xor ( n220601 , n33624 , n32139 );
xnor ( n220602 , n220601 , n204259 );
not ( n42842 , n26409 );
not ( n42843 , n204734 );
not ( n42844 , n26364 );
not ( n42845 , n42844 );
or ( n42846 , n42843 , n42845 );
or ( n42847 , n26365 , n204734 );
nand ( n42848 , n42846 , n42847 );
not ( n42849 , n42848 );
or ( n42850 , n42842 , n42849 );
or ( n42851 , n42848 , n26409 );
nand ( n220613 , n42850 , n42851 );
buf ( n220614 , n220613 );
not ( n42854 , n220614 );
nand ( n220616 , n220602 , n42854 );
not ( n220617 , n220616 );
buf ( n42857 , n208071 );
not ( n220619 , n42857 );
not ( n220620 , n41148 );
or ( n42860 , n220619 , n220620 );
or ( n220622 , n41148 , n42857 );
nand ( n220623 , n42860 , n220622 );
and ( n42863 , n220623 , n218917 );
not ( n42864 , n220623 );
and ( n42865 , n42864 , n37120 );
nor ( n42866 , n42863 , n42865 );
buf ( n42867 , n42866 );
not ( n42868 , n42867 );
and ( n220630 , n220617 , n42868 );
and ( n220631 , n220616 , n42867 );
nor ( n42871 , n220630 , n220631 );
buf ( n42872 , n42871 );
xor ( n42873 , n42839 , n42872 );
not ( n42874 , n34797 );
not ( n42875 , n42874 );
not ( n42876 , n29117 );
or ( n42877 , n42875 , n42876 );
nand ( n42878 , n29123 , n34797 );
nand ( n42879 , n42877 , n42878 );
not ( n42880 , n42879 );
not ( n220642 , n29175 );
and ( n220643 , n42880 , n220642 );
and ( n42883 , n42879 , n29175 );
nor ( n42884 , n220643 , n42883 );
not ( n42885 , n42884 );
not ( n42886 , n42885 );
not ( n42887 , n38839 );
nor ( n42888 , n39267 , n25784 );
not ( n42889 , n42888 );
not ( n42890 , n25780 );
nand ( n220652 , n42890 , n214870 );
nand ( n220653 , n42889 , n220652 );
not ( n42893 , n220653 );
and ( n220655 , n42887 , n42893 );
and ( n220656 , n38839 , n220653 );
nor ( n42896 , n220655 , n220656 );
not ( n42897 , n206940 );
not ( n42898 , n30200 );
or ( n42899 , n42897 , n42898 );
not ( n42900 , n206940 );
nand ( n42901 , n42900 , n30205 );
nand ( n42902 , n42899 , n42901 );
and ( n42903 , n42902 , n42189 );
not ( n42904 , n42902 );
and ( n42905 , n42904 , n31832 );
nor ( n220667 , n42903 , n42905 );
not ( n220668 , n220667 );
nand ( n42908 , n42896 , n220668 );
not ( n42909 , n42908 );
or ( n42910 , n42886 , n42909 );
or ( n42911 , n42908 , n42885 );
nand ( n42912 , n42910 , n42911 );
not ( n42913 , n42912 );
not ( n42914 , n40834 );
buf ( n42915 , RI19a860c0_2752);
nand ( n42916 , n25850 , n42915 );
buf ( n42917 , RI17502948_752);
and ( n220679 , n42916 , n42917 );
not ( n220680 , n42916 );
not ( n42920 , RI17502948_752);
and ( n42921 , n220680 , n42920 );
nor ( n42922 , n220679 , n42921 );
not ( n42923 , n42922 );
buf ( n42924 , RI19aa4cf0_2531);
nand ( n42925 , n25479 , n42924 );
not ( n42926 , RI17481060_1107);
and ( n42927 , n42925 , n42926 );
not ( n220689 , n42925 );
buf ( n220690 , RI17481060_1107);
and ( n42930 , n220689 , n220690 );
nor ( n42931 , n42927 , n42930 );
not ( n42932 , n42931 );
or ( n42933 , n42923 , n42932 );
or ( n42934 , n42922 , n42931 );
nand ( n42935 , n42933 , n42934 );
buf ( n42936 , RI173e4d78_1640);
not ( n42937 , n42936 );
not ( n42938 , RI1739bd40_1996);
not ( n42939 , n42938 );
or ( n42940 , n42937 , n42939 );
not ( n42941 , RI173e4d78_1640);
buf ( n42942 , RI1739bd40_1996);
nand ( n42943 , n42941 , n42942 );
nand ( n42944 , n42940 , n42943 );
not ( n42945 , RI1745c850_1285);
and ( n42946 , n42944 , n42945 );
not ( n42947 , n42944 );
buf ( n42948 , RI1745c850_1285);
and ( n42949 , n42947 , n42948 );
nor ( n42950 , n42946 , n42949 );
buf ( n42951 , n42950 );
and ( n42952 , n42935 , n42951 );
not ( n220714 , n42935 );
not ( n220715 , n42951 );
and ( n42955 , n220714 , n220715 );
nor ( n42956 , n42952 , n42955 );
not ( n42957 , n42956 );
or ( n42958 , n42914 , n42957 );
or ( n42959 , n42956 , n40834 );
nand ( n42960 , n42958 , n42959 );
not ( n42961 , n42960 );
not ( n42962 , n42961 );
not ( n42963 , RI173e22d0_1653);
xor ( n220725 , n42963 , n38648 );
xnor ( n220726 , n220725 , n216416 );
buf ( n42966 , n220726 );
not ( n42967 , n42966 );
or ( n42968 , n42962 , n42967 );
nand ( n42969 , n38657 , n42960 );
nand ( n42970 , n42968 , n42969 );
not ( n42971 , n42970 );
buf ( n42972 , RI1740c6c0_1447);
not ( n42973 , n42972 );
not ( n42974 , n29415 );
or ( n42975 , n42973 , n42974 );
not ( n220737 , n42972 );
nand ( n220738 , n220737 , n38204 );
nand ( n42978 , n42975 , n220738 );
and ( n42979 , n42978 , n29456 );
not ( n42980 , n42978 );
and ( n42981 , n42980 , n207216 );
nor ( n42982 , n42979 , n42981 );
nand ( n42983 , n42971 , n42982 );
not ( n42984 , n42983 );
not ( n42985 , n41280 );
not ( n42986 , n207493 );
or ( n42987 , n42985 , n42986 );
or ( n220749 , n207493 , n41280 );
nand ( n220750 , n42987 , n220749 );
xor ( n42990 , n220750 , n33444 );
not ( n42991 , n42990 );
not ( n42992 , n42991 );
and ( n42993 , n42984 , n42992 );
and ( n42994 , n42983 , n42991 );
nor ( n42995 , n42993 , n42994 );
not ( n42996 , n42995 );
and ( n42997 , n42913 , n42996 );
and ( n42998 , n42912 , n42995 );
nor ( n42999 , n42997 , n42998 );
buf ( n220761 , n42999 );
and ( n220762 , n42873 , n220761 );
not ( n43002 , n42873 );
not ( n43003 , n220761 );
and ( n43004 , n43002 , n43003 );
nor ( n43005 , n220762 , n43004 );
buf ( n43006 , n43005 );
and ( n43007 , n42708 , n43006 );
not ( n220769 , n42708 );
xor ( n220770 , n42871 , n42839 );
xnor ( n43010 , n220770 , n42999 );
buf ( n43011 , n43010 );
and ( n43012 , n220769 , n43011 );
nor ( n43013 , n43007 , n43012 );
not ( n43014 , n39211 );
not ( n43015 , n43014 );
not ( n43016 , n30865 );
not ( n43017 , n36455 );
or ( n220779 , n43016 , n43017 );
or ( n220780 , n36455 , n30865 );
nand ( n43020 , n220779 , n220780 );
not ( n43021 , n43020 );
or ( n43022 , n43015 , n43021 );
or ( n43023 , n43020 , n43014 );
nand ( n43024 , n43022 , n43023 );
not ( n43025 , n43024 );
not ( n43026 , n205426 );
buf ( n43027 , n29297 );
not ( n43028 , n43027 );
not ( n43029 , n43028 );
not ( n43030 , n33362 );
or ( n220792 , n43029 , n43030 );
nand ( n220793 , n33366 , n43027 );
nand ( n43033 , n220792 , n220793 );
not ( n43034 , n43033 );
and ( n43035 , n43026 , n43034 );
and ( n43036 , n205426 , n43033 );
nor ( n43037 , n43035 , n43036 );
not ( n43038 , n33021 );
not ( n43039 , n37254 );
and ( n43040 , n43038 , n43039 );
and ( n43041 , n33021 , n37254 );
nor ( n43042 , n43040 , n43041 );
not ( n220804 , n43042 );
not ( n220805 , n33041 );
or ( n43045 , n220804 , n220805 );
or ( n43046 , n33041 , n43042 );
nand ( n43047 , n43045 , n43046 );
and ( n43048 , n43047 , n33013 );
not ( n43049 , n43047 );
and ( n43050 , n43049 , n40312 );
nor ( n43051 , n43048 , n43050 );
nand ( n43052 , n43037 , n43051 );
not ( n220814 , n43052 );
or ( n220815 , n43025 , n220814 );
or ( n43055 , n43052 , n43024 );
nand ( n43056 , n220815 , n43055 );
not ( n43057 , n43056 );
buf ( n43058 , n41853 );
not ( n43059 , n43058 );
not ( n43060 , RI173dfeb8_1664);
not ( n43061 , n206658 );
xor ( n43062 , n43060 , n43061 );
xnor ( n43063 , n43062 , n28905 );
not ( n43064 , n43063 );
not ( n220826 , n43064 );
or ( n220827 , n43059 , n220826 );
or ( n43067 , n43064 , n43058 );
nand ( n43068 , n220827 , n43067 );
and ( n43069 , n43068 , n30936 );
not ( n43070 , n43068 );
and ( n43071 , n43070 , n30943 );
nor ( n43072 , n43069 , n43071 );
buf ( n43073 , n219052 );
not ( n43074 , n43073 );
not ( n220836 , n38782 );
not ( n220837 , n220836 );
not ( n43077 , n37648 );
or ( n43078 , n220837 , n43077 );
or ( n43079 , n37648 , n220836 );
nand ( n43080 , n43078 , n43079 );
not ( n43081 , n43080 );
not ( n43082 , n43081 );
or ( n220844 , n43074 , n43082 );
buf ( n220845 , n41303 );
nand ( n43085 , n43080 , n220845 );
nand ( n43086 , n220844 , n43085 );
nand ( n43087 , n43072 , n43086 );
not ( n43088 , n43087 );
not ( n220850 , n26369 );
not ( n220851 , n204732 );
and ( n43091 , n220850 , n220851 );
and ( n43092 , n26369 , n204732 );
nor ( n43093 , n43091 , n43092 );
and ( n43094 , n43093 , n26409 );
not ( n43095 , n43093 );
not ( n43096 , n26408 );
and ( n43097 , n43095 , n43096 );
nor ( n43098 , n43094 , n43097 );
not ( n43099 , n43098 );
and ( n43100 , n43088 , n43099 );
and ( n43101 , n43087 , n43098 );
nor ( n220863 , n43100 , n43101 );
not ( n220864 , n220863 );
or ( n43104 , n43057 , n220864 );
or ( n43105 , n220863 , n43056 );
nand ( n43106 , n43104 , n43105 );
buf ( n220868 , n209579 );
not ( n220869 , n220868 );
not ( n43109 , n220869 );
not ( n43110 , n27759 );
or ( n43111 , n43109 , n43110 );
not ( n43112 , n27759 );
nand ( n43113 , n43112 , n220868 );
nand ( n43114 , n43111 , n43113 );
and ( n43115 , n43114 , n34644 );
not ( n43116 , n43114 );
not ( n220878 , n34644 );
and ( n220879 , n43116 , n220878 );
nor ( n43119 , n43115 , n220879 );
and ( n43120 , n26316 , n38973 );
not ( n43121 , n26316 );
buf ( n43122 , n38972 );
and ( n43123 , n43121 , n43122 );
nor ( n43124 , n43120 , n43123 );
not ( n220886 , n43124 );
not ( n220887 , n39007 );
and ( n43127 , n220886 , n220887 );
and ( n220889 , n43124 , n39009 );
nor ( n220890 , n43127 , n220889 );
nand ( n43130 , n43119 , n220890 );
nor ( n220892 , n31428 , n31179 );
not ( n220893 , n220892 );
nand ( n43133 , n40270 , n31179 );
nand ( n220895 , n220893 , n43133 );
not ( n220896 , n42285 );
and ( n43136 , n220895 , n220896 );
not ( n43137 , n220895 );
and ( n43138 , n43137 , n42285 );
nor ( n43139 , n43136 , n43138 );
not ( n43140 , n43139 );
xor ( n43141 , n43130 , n43140 );
not ( n43142 , n43141 );
and ( n43143 , n43106 , n43142 );
not ( n220905 , n43106 );
and ( n220906 , n220905 , n43141 );
nor ( n43146 , n43143 , n220906 );
not ( n43147 , n43146 );
buf ( n43148 , n30600 );
not ( n43149 , n43148 );
not ( n43150 , n27842 );
or ( n43151 , n43149 , n43150 );
not ( n43152 , n43148 );
nand ( n43153 , n43152 , n32454 );
nand ( n43154 , n43151 , n43153 );
not ( n43155 , n27802 );
and ( n220917 , n43154 , n43155 );
not ( n220918 , n43154 );
and ( n43158 , n220918 , n27802 );
nor ( n43159 , n220917 , n43158 );
not ( n43160 , n43159 );
xor ( n43161 , n41700 , n35275 );
xor ( n43162 , n43161 , n36093 );
nand ( n43163 , n43160 , n43162 );
not ( n43164 , n43163 );
not ( n43165 , n39707 );
not ( n43166 , n43165 );
not ( n43167 , n37429 );
not ( n220929 , n31900 );
or ( n220930 , n43167 , n220929 );
or ( n43170 , n31900 , n37429 );
nand ( n220932 , n220930 , n43170 );
not ( n220933 , n220932 );
or ( n43173 , n43166 , n220933 );
or ( n43174 , n220932 , n43165 );
nand ( n43175 , n43173 , n43174 );
not ( n43176 , n43175 );
not ( n43177 , n43176 );
not ( n43178 , n43177 );
and ( n43179 , n43164 , n43178 );
not ( n43180 , n43159 );
nand ( n43181 , n43180 , n43162 );
and ( n43182 , n43181 , n43177 );
nor ( n220944 , n43179 , n43182 );
not ( n220945 , n220944 );
buf ( n43185 , n36346 );
xor ( n43186 , n43185 , n41894 );
xnor ( n43187 , n43186 , n31078 );
not ( n43188 , n30935 );
not ( n43189 , n218656 );
or ( n43190 , n43188 , n43189 );
not ( n220952 , n30935 );
not ( n220953 , n218656 );
nand ( n43193 , n220952 , n220953 );
nand ( n43194 , n43190 , n43193 );
and ( n43195 , n43194 , n41904 );
not ( n43196 , n43194 );
not ( n43197 , n41904 );
and ( n43198 , n43196 , n43197 );
nor ( n43199 , n43195 , n43198 );
nand ( n43200 , n43187 , n43199 );
not ( n43201 , n38435 );
xor ( n43202 , n29498 , n43201 );
not ( n220964 , n216225 );
not ( n220965 , n220964 );
xor ( n43205 , n43202 , n220965 );
not ( n43206 , n43205 );
and ( n43207 , n43200 , n43206 );
not ( n43208 , n43200 );
and ( n43209 , n43208 , n43205 );
nor ( n43210 , n43207 , n43209 );
not ( n43211 , n43210 );
or ( n43212 , n220945 , n43211 );
or ( n43213 , n43210 , n220944 );
nand ( n43214 , n43212 , n43213 );
not ( n220976 , n43214 );
or ( n220977 , n43147 , n220976 );
or ( n43217 , n43214 , n43146 );
nand ( n43218 , n220977 , n43217 );
buf ( n43219 , n43218 );
not ( n43220 , n43219 );
not ( n43221 , n43220 );
not ( n43222 , n39243 );
not ( n220984 , n28404 );
not ( n220985 , n220984 );
or ( n43225 , n43222 , n220985 );
or ( n43226 , n220984 , n39243 );
nand ( n43227 , n43225 , n43226 );
buf ( n43228 , RI173d6138_1712);
not ( n43229 , n43228 );
not ( n43230 , RI1738d448_2067);
not ( n43231 , n43230 );
or ( n220993 , n43229 , n43231 );
not ( n220994 , RI173d6138_1712);
buf ( n43234 , RI1738d448_2067);
nand ( n43235 , n220994 , n43234 );
nand ( n43236 , n220993 , n43235 );
not ( n43237 , RI1744dc10_1357);
and ( n43238 , n43236 , n43237 );
not ( n43239 , n43236 );
buf ( n43240 , RI1744dc10_1357);
and ( n43241 , n43239 , n43240 );
nor ( n43242 , n43238 , n43241 );
buf ( n43243 , RI19a9b678_2602);
nand ( n43244 , n25741 , n43243 );
buf ( n221006 , RI17472420_1179);
and ( n221007 , n43244 , n221006 );
not ( n43247 , n43244 );
not ( n43248 , RI17472420_1179);
and ( n43249 , n43247 , n43248 );
nor ( n43250 , n221007 , n43249 );
xor ( n43251 , n43242 , n43250 );
buf ( n43252 , RI19acabf8_2250);
nand ( n221014 , n25540 , n43252 );
not ( n221015 , RI174bc7f0_824);
and ( n43255 , n221014 , n221015 );
not ( n43256 , n221014 );
buf ( n43257 , RI174bc7f0_824);
and ( n43258 , n43256 , n43257 );
nor ( n43259 , n43255 , n43258 );
xnor ( n43260 , n43251 , n43259 );
buf ( n43261 , n43260 );
not ( n43262 , n43261 );
and ( n43263 , n43227 , n43262 );
not ( n43264 , n43227 );
and ( n43265 , n43264 , n43261 );
nor ( n43266 , n43263 , n43265 );
not ( n43267 , n25983 );
xor ( n43268 , n33916 , n33934 );
not ( n43269 , n33925 );
xnor ( n43270 , n43268 , n43269 );
not ( n43271 , n43270 );
or ( n43272 , n43267 , n43271 );
not ( n43273 , n25983 );
not ( n43274 , n43270 );
nand ( n43275 , n43273 , n43274 );
nand ( n43276 , n43272 , n43275 );
and ( n43277 , n43276 , n41082 );
not ( n43278 , n43276 );
not ( n43279 , n32900 );
and ( n43280 , n43278 , n43279 );
nor ( n43281 , n43277 , n43280 );
nand ( n43282 , n43266 , n43281 );
not ( n43283 , n33015 );
not ( n43284 , n36138 );
or ( n43285 , n43283 , n43284 );
or ( n43286 , n36138 , n33015 );
nand ( n43287 , n43285 , n43286 );
and ( n221049 , n36162 , n36128 );
not ( n221050 , n36162 );
and ( n43290 , n221050 , n213927 );
nor ( n43291 , n221049 , n43290 );
xor ( n43292 , n43287 , n43291 );
nor ( n43293 , n36187 , n43292 );
not ( n43294 , n43293 );
nand ( n43295 , n36189 , n43292 );
nand ( n43296 , n43294 , n43295 );
not ( n43297 , n43296 );
and ( n43298 , n43282 , n43297 );
not ( n43299 , n43282 );
and ( n221061 , n43299 , n43296 );
nor ( n221062 , n43298 , n221061 );
not ( n43302 , n221062 );
xor ( n43303 , n33102 , n40621 );
xnor ( n43304 , n43303 , n39020 );
not ( n43305 , n208672 );
not ( n43306 , n218656 );
or ( n43307 , n43305 , n43306 );
or ( n221069 , n218656 , n208672 );
nand ( n221070 , n43307 , n221069 );
not ( n43310 , n221070 );
not ( n43311 , n41904 );
and ( n43312 , n43310 , n43311 );
and ( n43313 , n221070 , n41904 );
nor ( n43314 , n43312 , n43313 );
not ( n43315 , n43314 );
nand ( n43316 , n43304 , n43315 );
not ( n43317 , n43316 );
not ( n43318 , n220343 );
not ( n43319 , n213041 );
or ( n221081 , n43318 , n43319 );
not ( n221082 , n220343 );
nand ( n43322 , n221082 , n215580 );
nand ( n43323 , n221081 , n43322 );
and ( n43324 , n43323 , n34564 );
not ( n43325 , n43323 );
buf ( n43326 , n34558 );
and ( n43327 , n43325 , n43326 );
nor ( n43328 , n43324 , n43327 );
buf ( n43329 , n43328 );
not ( n221091 , n43329 );
not ( n221092 , n221091 );
and ( n43332 , n43317 , n221092 );
and ( n221094 , n43316 , n221091 );
nor ( n221095 , n43332 , n221094 );
not ( n43335 , n221095 );
not ( n43336 , n43335 );
and ( n43337 , n220505 , n35923 );
not ( n43338 , n220505 );
xor ( n43339 , n35904 , n35912 );
xnor ( n43340 , n43339 , n35921 );
and ( n43341 , n43338 , n43340 );
nor ( n43342 , n43337 , n43341 );
and ( n43343 , n43342 , n41395 );
not ( n43344 , n43342 );
and ( n221106 , n43344 , n41398 );
nor ( n221107 , n43343 , n221106 );
not ( n43347 , n28843 );
not ( n43348 , n37652 );
or ( n43349 , n43347 , n43348 );
or ( n43350 , n37652 , n28843 );
nand ( n43351 , n43349 , n43350 );
and ( n43352 , n43351 , n220845 );
not ( n43353 , n43351 );
and ( n221115 , n43353 , n43073 );
nor ( n221116 , n43352 , n221115 );
nand ( n221117 , n221107 , n221116 );
not ( n221118 , n221117 );
not ( n43358 , n204825 );
and ( n221120 , n39301 , n31394 );
not ( n221121 , n39301 );
and ( n43361 , n221121 , n31398 );
or ( n43362 , n221120 , n43361 );
not ( n43363 , n43362 );
buf ( n43364 , n39313 );
not ( n43365 , n43364 );
or ( n43366 , n43363 , n43365 );
or ( n221128 , n43364 , n43362 );
nand ( n221129 , n43366 , n221128 );
not ( n43369 , n221129 );
and ( n43370 , n43358 , n43369 );
and ( n43371 , n204825 , n221129 );
nor ( n43372 , n43370 , n43371 );
not ( n43373 , n43372 );
not ( n43374 , n43373 );
and ( n43375 , n221118 , n43374 );
and ( n43376 , n221117 , n43373 );
nor ( n221138 , n43375 , n43376 );
not ( n221139 , n221138 );
and ( n43379 , n40111 , n25642 );
not ( n43380 , n40111 );
and ( n43381 , n43380 , n25646 );
or ( n43382 , n43379 , n43381 );
and ( n43383 , n43382 , n40131 );
not ( n43384 , n43382 );
and ( n43385 , n43384 , n40130 );
nor ( n43386 , n43383 , n43385 );
not ( n221148 , n43386 );
buf ( n221149 , n40101 );
not ( n43389 , n221149 );
and ( n43390 , n221148 , n43389 );
and ( n43391 , n43386 , n221149 );
nor ( n43392 , n43390 , n43391 );
not ( n221154 , n43392 );
not ( n221155 , n221154 );
not ( n43395 , n43281 );
nand ( n43396 , n43297 , n43395 );
not ( n43397 , n43396 );
or ( n43398 , n221155 , n43397 );
or ( n43399 , n43396 , n221154 );
nand ( n43400 , n43398 , n43399 );
not ( n43401 , n43400 );
or ( n43402 , n221139 , n43401 );
or ( n43403 , n43400 , n221138 );
nand ( n43404 , n43402 , n43403 );
not ( n221166 , n43404 );
not ( n221167 , n221166 );
or ( n43407 , n43336 , n221167 );
nand ( n43408 , n43404 , n221095 );
nand ( n43409 , n43407 , n43408 );
not ( n43410 , n31808 );
not ( n43411 , n27759 );
or ( n43412 , n43410 , n43411 );
nand ( n43413 , n27758 , n31805 );
nand ( n43414 , n43412 , n43413 );
not ( n43415 , n43414 );
not ( n43416 , n220878 );
and ( n221178 , n43415 , n43416 );
and ( n221179 , n220878 , n43414 );
nor ( n43419 , n221178 , n221179 );
not ( n43420 , n43419 );
not ( n43421 , n32964 );
not ( n43422 , n29910 );
or ( n43423 , n43421 , n43422 );
not ( n43424 , n32964 );
nand ( n43425 , n43424 , n29913 );
nand ( n43426 , n43423 , n43425 );
and ( n43427 , n43426 , n207706 );
not ( n43428 , n43426 );
and ( n221190 , n43428 , n29948 );
nor ( n221191 , n43427 , n221190 );
nand ( n43431 , n43420 , n221191 );
not ( n43432 , n32545 );
not ( n43433 , n28463 );
or ( n43434 , n43432 , n43433 );
or ( n221196 , n28463 , n32545 );
nand ( n221197 , n43434 , n221196 );
and ( n43437 , n221197 , n28511 );
not ( n43438 , n221197 );
and ( n43439 , n43438 , n28503 );
nor ( n43440 , n43437 , n43439 );
not ( n43441 , n43440 );
and ( n43442 , n43431 , n43441 );
not ( n221204 , n43431 );
and ( n221205 , n221204 , n43440 );
nor ( n43445 , n43442 , n221205 );
not ( n43446 , n43445 );
not ( n43447 , n43446 );
not ( n43448 , n28055 );
not ( n43449 , n39798 );
or ( n43450 , n43448 , n43449 );
not ( n43451 , n28055 );
nand ( n43452 , n43451 , n41894 );
nand ( n43453 , n43450 , n43452 );
and ( n43454 , n43453 , n25429 );
not ( n43455 , n43453 );
and ( n43456 , n43455 , n25426 );
nor ( n43457 , n43454 , n43456 );
not ( n43458 , n43457 );
not ( n43459 , n40413 );
not ( n43460 , n43459 );
buf ( n43461 , n43460 );
xor ( n43462 , n207591 , n43461 );
xnor ( n43463 , n43462 , n41878 );
not ( n43464 , n43463 );
nand ( n43465 , n43458 , n43464 );
not ( n43466 , n43465 );
not ( n43467 , n28665 );
not ( n43468 , n207380 );
not ( n43469 , n36520 );
not ( n43470 , n43469 );
or ( n221232 , n43468 , n43470 );
not ( n221233 , n36520 );
buf ( n43473 , n221233 );
or ( n43474 , n43473 , n207380 );
nand ( n43475 , n221232 , n43474 );
not ( n43476 , n43475 );
or ( n43477 , n43467 , n43476 );
or ( n43478 , n28665 , n43475 );
nand ( n43479 , n43477 , n43478 );
buf ( n43480 , n43479 );
not ( n43481 , n43480 );
and ( n43482 , n43466 , n43481 );
not ( n43483 , n43457 );
nand ( n43484 , n43483 , n43464 );
and ( n43485 , n43484 , n43480 );
nor ( n43486 , n43482 , n43485 );
not ( n43487 , n43486 );
not ( n43488 , n43487 );
or ( n43489 , n43447 , n43488 );
nand ( n43490 , n43486 , n43445 );
nand ( n43491 , n43489 , n43490 );
and ( n43492 , n43409 , n43491 );
not ( n43493 , n43409 );
not ( n43494 , n43491 );
and ( n43495 , n43493 , n43494 );
nor ( n43496 , n43492 , n43495 );
not ( n43497 , n43496 );
not ( n43498 , n43497 );
or ( n43499 , n43302 , n43498 );
not ( n43500 , n221062 );
and ( n43501 , n43409 , n43491 );
not ( n221263 , n43409 );
and ( n221264 , n221263 , n43494 );
nor ( n43504 , n43501 , n221264 );
nand ( n43505 , n43500 , n43504 );
nand ( n43506 , n43499 , n43505 );
not ( n43507 , n43506 );
or ( n43508 , n43221 , n43507 );
or ( n43509 , n43506 , n43220 );
nand ( n221271 , n43508 , n43509 );
not ( n221272 , n221271 );
nand ( n43512 , n42444 , n43013 , n221272 );
not ( n43513 , n42442 );
not ( n43514 , n43513 );
not ( n43515 , n43013 );
or ( n43516 , n43514 , n43515 );
buf ( n43517 , n27886 );
buf ( n221279 , n43517 );
nor ( n221280 , n221272 , n221279 );
nand ( n221281 , n43516 , n221280 );
nand ( n221282 , n31577 , n206564 );
nand ( n43522 , n43512 , n221281 , n221282 );
buf ( n43523 , n43522 );
not ( n43524 , RI19ac6ff8_2277);
or ( n43525 , n25328 , n43524 );
not ( n43526 , RI19abe100_2349);
or ( n43527 , n25336 , n43526 );
nand ( n43528 , n43525 , n43527 );
buf ( n43529 , n43528 );
buf ( n221291 , n31895 );
nand ( n221292 , n42420 , n42409 );
not ( n43532 , n221292 );
not ( n43533 , n42058 );
not ( n43534 , n25947 );
not ( n43535 , n32006 );
or ( n43536 , n43534 , n43535 );
nand ( n43537 , n35622 , n25944 );
nand ( n43538 , n43536 , n43537 );
not ( n43539 , n43538 );
or ( n43540 , n43533 , n43539 );
or ( n43541 , n43538 , n41114 );
nand ( n221303 , n43540 , n43541 );
not ( n221304 , n221303 );
and ( n43544 , n43532 , n221304 );
and ( n43545 , n221292 , n221303 );
nor ( n43546 , n43544 , n43545 );
not ( n43547 , n43546 );
not ( n43548 , n35756 );
not ( n43549 , n39480 );
or ( n43550 , n43548 , n43549 );
or ( n221312 , n39480 , n35756 );
nand ( n221313 , n43550 , n221312 );
buf ( n43553 , n35097 );
buf ( n43554 , n43553 );
and ( n43555 , n221313 , n43554 );
not ( n43556 , n221313 );
not ( n43557 , n43553 );
and ( n43558 , n43556 , n43557 );
nor ( n221320 , n43555 , n43558 );
nand ( n221321 , n42194 , n221320 );
not ( n43561 , n221321 );
buf ( n221323 , n34872 );
xor ( n221324 , n205247 , n221323 );
xnor ( n43564 , n221324 , n31778 );
not ( n43565 , n43564 );
or ( n43566 , n43561 , n43565 );
or ( n43567 , n43564 , n221321 );
nand ( n43568 , n43566 , n43567 );
not ( n43569 , n43568 );
not ( n43570 , n43569 );
not ( n43571 , n204558 );
not ( n43572 , n28381 );
or ( n43573 , n43571 , n43572 );
not ( n221335 , n204558 );
nand ( n221336 , n221335 , n28380 );
nand ( n43576 , n43573 , n221336 );
not ( n43577 , n30136 );
and ( n221339 , n43576 , n43577 );
not ( n221340 , n43576 );
and ( n43580 , n221340 , n30137 );
nor ( n43581 , n221339 , n43580 );
not ( n43582 , n43581 );
nand ( n43583 , n43582 , n42380 );
not ( n43584 , n43583 );
not ( n43585 , n204744 );
not ( n43586 , n33904 );
not ( n43587 , n204727 );
or ( n43588 , n43586 , n43587 );
not ( n43589 , n204723 );
nand ( n43590 , n43589 , n33908 );
nand ( n43591 , n43588 , n43590 );
not ( n221353 , n43591 );
not ( n221354 , n221353 );
or ( n43594 , n43585 , n221354 );
nand ( n43595 , n36705 , n43591 );
nand ( n43596 , n43594 , n43595 );
not ( n43597 , n43596 );
and ( n43598 , n43584 , n43597 );
not ( n43599 , n43581 );
nand ( n43600 , n43599 , n42380 );
and ( n221362 , n43600 , n43596 );
nor ( n221363 , n43598 , n221362 );
not ( n43603 , n221363 );
not ( n221365 , n43603 );
or ( n221366 , n43570 , n221365 );
nand ( n43606 , n221363 , n43568 );
nand ( n221368 , n221366 , n43606 );
not ( n221369 , n221303 );
nand ( n43609 , n221369 , n42421 );
not ( n43610 , n43609 );
buf ( n43611 , RI173ed400_1599);
not ( n43612 , n43611 );
not ( n43613 , n36035 );
or ( n43614 , n43612 , n43613 );
not ( n43615 , RI173ed400_1599);
buf ( n43616 , RI173a4710_1954);
nand ( n221378 , n43615 , n43616 );
nand ( n221379 , n43614 , n221378 );
not ( n43619 , RI17489d78_1064);
and ( n43620 , n221379 , n43619 );
not ( n43621 , n221379 );
buf ( n43622 , RI17489d78_1064);
and ( n43623 , n43621 , n43622 );
nor ( n43624 , n43620 , n43623 );
xor ( n43625 , n43624 , n37742 );
buf ( n43626 , RI19acd808_2228);
nand ( n43627 , n25656 , n43626 );
buf ( n43628 , RI17511b28_711);
and ( n221390 , n43627 , n43628 );
not ( n221391 , n43627 );
not ( n43631 , RI17511b28_711);
and ( n43632 , n221391 , n43631 );
nor ( n43633 , n221390 , n43632 );
not ( n43634 , n43633 );
xnor ( n43635 , n43625 , n43634 );
buf ( n43636 , n43635 );
not ( n43637 , n43636 );
not ( n43638 , n35248 );
not ( n43639 , n36934 );
or ( n43640 , n43638 , n43639 );
xor ( n221402 , n36915 , n36932 );
xnor ( n221403 , n221402 , n40585 );
nand ( n43643 , n221403 , n35244 );
nand ( n43644 , n43640 , n43643 );
not ( n43645 , n43644 );
or ( n221407 , n43637 , n43645 );
or ( n221408 , n43644 , n43635 );
nand ( n43648 , n221407 , n221408 );
not ( n43649 , n43648 );
and ( n43650 , n43610 , n43649 );
not ( n43651 , n221303 );
nand ( n43652 , n43651 , n42421 );
and ( n43653 , n43652 , n43648 );
nor ( n43654 , n43650 , n43653 );
not ( n43655 , n43654 );
and ( n43656 , n221368 , n43655 );
not ( n43657 , n221368 );
and ( n221419 , n43657 , n43654 );
nor ( n221420 , n43656 , n221419 );
not ( n43660 , n221420 );
not ( n43661 , n35837 );
not ( n43662 , n205142 );
or ( n43663 , n43661 , n43662 );
or ( n43664 , n205096 , n35837 );
nand ( n43665 , n43663 , n43664 );
xor ( n43666 , n43665 , n33300 );
nand ( n43667 , n219992 , n43666 );
not ( n43668 , n43667 );
not ( n43669 , n28889 );
xor ( n221431 , n40842 , n40859 );
buf ( n221432 , n40850 );
xnor ( n43672 , n221431 , n221432 );
buf ( n221434 , n43672 );
not ( n221435 , n221434 );
or ( n43675 , n43669 , n221435 );
or ( n221437 , n221434 , n28889 );
nand ( n221438 , n43675 , n221437 );
and ( n43678 , n221438 , n218656 );
not ( n43679 , n221438 );
and ( n43680 , n43679 , n40896 );
nor ( n43681 , n43678 , n43680 );
not ( n43682 , n43681 );
not ( n43683 , n43682 );
and ( n43684 , n43668 , n43683 );
not ( n43685 , n219993 );
nand ( n221447 , n43685 , n43666 );
and ( n221448 , n221447 , n43682 );
nor ( n43688 , n43684 , n221448 );
not ( n43689 , n43688 );
xor ( n43690 , n30249 , n37212 );
xnor ( n43691 , n43690 , n204621 );
not ( n43692 , n43691 );
buf ( n43693 , RI173bb9d8_1841);
not ( n43694 , n43693 );
not ( n43695 , n40812 );
not ( n43696 , n43695 );
not ( n43697 , n43696 );
or ( n221459 , n43694 , n43697 );
or ( n221460 , n43696 , n43693 );
nand ( n43700 , n221459 , n221460 );
not ( n221462 , n29371 );
not ( n221463 , n221462 );
and ( n43703 , n43700 , n221463 );
not ( n43704 , n43700 );
not ( n43705 , n29372 );
and ( n43706 , n43704 , n43705 );
nor ( n43707 , n43703 , n43706 );
nand ( n43708 , n43707 , n42311 );
not ( n43709 , n43708 );
or ( n43710 , n43692 , n43709 );
or ( n43711 , n43708 , n43691 );
nand ( n43712 , n43710 , n43711 );
not ( n43713 , n43712 );
or ( n43714 , n43689 , n43713 );
or ( n43715 , n43712 , n43688 );
nand ( n43716 , n43714 , n43715 );
not ( n221478 , n43716 );
not ( n221479 , n221478 );
or ( n43719 , n43660 , n221479 );
not ( n43720 , n221420 );
nand ( n43721 , n43720 , n43716 );
nand ( n43722 , n43719 , n43721 );
not ( n43723 , n43722 );
or ( n43724 , n43547 , n43723 );
not ( n43725 , n43722 );
not ( n43726 , n43725 );
or ( n43727 , n43726 , n43546 );
nand ( n43728 , n43724 , n43727 );
and ( n43729 , n37258 , n37255 );
not ( n221491 , n37258 );
buf ( n221492 , RI174a2738_944);
and ( n43732 , n221491 , n221492 );
nor ( n43733 , n43729 , n43732 );
xor ( n43734 , n43733 , n32406 );
not ( n43735 , n33046 );
xnor ( n43736 , n43734 , n43735 );
not ( n43737 , n43736 );
not ( n43738 , n43737 );
not ( n43739 , n205420 );
buf ( n43740 , n29324 );
not ( n221502 , n43740 );
and ( n221503 , n43739 , n221502 );
and ( n43743 , n205420 , n43740 );
nor ( n43744 , n221503 , n43743 );
and ( n43745 , n43744 , n205436 );
not ( n43746 , n43744 );
and ( n43747 , n43746 , n205435 );
nor ( n43748 , n43745 , n43747 );
not ( n43749 , n43748 );
not ( n43750 , n204815 );
not ( n43751 , n205068 );
or ( n43752 , n43750 , n43751 );
not ( n221514 , n204815 );
nand ( n221515 , n221514 , n205074 );
nand ( n43755 , n43752 , n221515 );
not ( n43756 , n43755 );
buf ( n43757 , n33178 );
not ( n43758 , n43757 );
not ( n43759 , n43758 );
and ( n221521 , n43756 , n43759 );
and ( n221522 , n43755 , n43758 );
nor ( n43762 , n221521 , n221522 );
not ( n43763 , n43762 );
nand ( n43764 , n43749 , n43763 );
not ( n43765 , n43764 );
or ( n43766 , n43738 , n43765 );
or ( n43767 , n43764 , n43737 );
nand ( n43768 , n43766 , n43767 );
not ( n43769 , n43768 );
buf ( n43770 , n204965 );
not ( n43771 , n43770 );
not ( n43772 , n36025 );
or ( n43773 , n43771 , n43772 );
or ( n221535 , n36025 , n43770 );
nand ( n221536 , n43773 , n221535 );
and ( n221537 , n221536 , n40862 );
not ( n221538 , n221536 );
and ( n43778 , n221538 , n221434 );
nor ( n43779 , n221537 , n43778 );
not ( n43780 , n43779 );
not ( n43781 , n32148 );
not ( n221543 , n33614 );
or ( n221544 , n43781 , n221543 );
not ( n43784 , n32148 );
nand ( n221546 , n43784 , n33618 );
nand ( n221547 , n221544 , n221546 );
not ( n43787 , n41520 );
and ( n43788 , n221547 , n43787 );
not ( n43789 , n221547 );
and ( n43790 , n43789 , n41520 );
nor ( n43791 , n43788 , n43790 );
not ( n43792 , n43791 );
nand ( n221554 , n43780 , n43792 );
not ( n221555 , n221554 );
not ( n43795 , n35773 );
not ( n43796 , n39481 );
or ( n43797 , n43795 , n43796 );
not ( n43798 , n35773 );
nand ( n43799 , n43798 , n40607 );
nand ( n43800 , n43797 , n43799 );
and ( n43801 , n43800 , n43554 );
not ( n43802 , n43800 );
not ( n43803 , n43554 );
and ( n43804 , n43802 , n43803 );
nor ( n221566 , n43801 , n43804 );
not ( n221567 , n221566 );
not ( n43807 , n221567 );
and ( n43808 , n221555 , n43807 );
and ( n43809 , n221554 , n221567 );
nor ( n43810 , n43808 , n43809 );
not ( n43811 , n43810 );
and ( n43812 , n43769 , n43811 );
and ( n43813 , n43768 , n43810 );
nor ( n43814 , n43812 , n43813 );
not ( n43815 , n43814 );
not ( n43816 , n43815 );
not ( n221578 , n43636 );
not ( n221579 , n35273 );
not ( n43819 , n36934 );
or ( n43820 , n221579 , n43819 );
not ( n43821 , n35273 );
nand ( n43822 , n43821 , n221403 );
nand ( n43823 , n43820 , n43822 );
not ( n43824 , n43823 );
or ( n43825 , n221578 , n43824 );
or ( n43826 , n43823 , n43636 );
nand ( n43827 , n43825 , n43826 );
not ( n43828 , n43827 );
not ( n221590 , n32209 );
not ( n221591 , n42512 );
or ( n43831 , n221590 , n221591 );
not ( n43832 , n32209 );
nand ( n43833 , n43832 , n220278 );
nand ( n43834 , n43831 , n43833 );
xor ( n221596 , n37328 , n215106 );
buf ( n221597 , n37336 );
xnor ( n43837 , n221596 , n221597 );
not ( n43838 , n43837 );
not ( n43839 , n43838 );
and ( n43840 , n43834 , n43839 );
not ( n43841 , n43834 );
not ( n43842 , n37346 );
not ( n221604 , n43842 );
and ( n221605 , n43841 , n221604 );
nor ( n43845 , n43840 , n221605 );
nand ( n43846 , n43828 , n43845 );
not ( n43847 , n43846 );
xor ( n43848 , n39694 , n39701 );
xnor ( n43849 , n43848 , n39705 );
not ( n43850 , n43849 );
buf ( n43851 , n32727 );
not ( n43852 , n43851 );
and ( n221614 , n43850 , n43852 );
and ( n221615 , n43849 , n43851 );
nor ( n43855 , n221614 , n221615 );
and ( n43856 , n43855 , n36377 );
not ( n43857 , n43855 );
and ( n43858 , n43857 , n35787 );
nor ( n43859 , n43856 , n43858 );
not ( n43860 , n43859 );
not ( n43861 , n43860 );
not ( n43862 , n43861 );
or ( n221624 , n43847 , n43862 );
nand ( n221625 , n43828 , n43845 );
or ( n43865 , n43861 , n221625 );
nand ( n43866 , n221624 , n43865 );
not ( n221628 , n43866 );
xor ( n221629 , n30822 , n36423 );
xnor ( n43869 , n221629 , n36456 );
not ( n43870 , n43869 );
not ( n43871 , n25994 );
not ( n43872 , n43270 );
or ( n43873 , n43871 , n43872 );
or ( n43874 , n43270 , n25994 );
nand ( n43875 , n43873 , n43874 );
and ( n43876 , n43875 , n32903 );
not ( n43877 , n43875 );
and ( n43878 , n43877 , n32900 );
nor ( n43879 , n43876 , n43878 );
not ( n221641 , n43879 );
nand ( n221642 , n43870 , n221641 );
not ( n43882 , n221642 );
buf ( n221644 , n28592 );
xor ( n221645 , n215140 , n37387 );
xnor ( n43885 , n221645 , n37396 );
and ( n43886 , n221644 , n43885 );
not ( n43887 , n221644 );
not ( n43888 , n37397 );
and ( n43889 , n43887 , n43888 );
nor ( n43890 , n43886 , n43889 );
xor ( n221652 , n30810 , n43890 );
not ( n221653 , n221652 );
not ( n43893 , n221653 );
and ( n43894 , n43882 , n43893 );
nand ( n43895 , n43870 , n221641 );
and ( n43896 , n43895 , n221653 );
nor ( n221658 , n43894 , n43896 );
not ( n221659 , n221658 );
or ( n43899 , n221628 , n221659 );
or ( n43900 , n221658 , n43866 );
nand ( n43901 , n43899 , n43900 );
not ( n43902 , n43901 );
not ( n43903 , n33875 );
not ( n43904 , n205216 );
or ( n43905 , n43903 , n43904 );
not ( n43906 , n205221 );
or ( n221668 , n43906 , n33875 );
nand ( n221669 , n43905 , n221668 );
not ( n43909 , n221669 );
buf ( n43910 , n35200 );
not ( n43911 , n43910 );
and ( n43912 , n43909 , n43911 );
buf ( n43913 , n35199 );
not ( n43914 , n43913 );
and ( n43915 , n221669 , n43914 );
nor ( n43916 , n43912 , n43915 );
not ( n43917 , n43916 );
buf ( n43918 , n37059 );
not ( n221680 , n43918 );
not ( n221681 , n43695 );
or ( n43921 , n221680 , n221681 );
or ( n43922 , n40814 , n43918 );
nand ( n43923 , n43921 , n43922 );
not ( n43924 , n43923 );
not ( n43925 , n29372 );
and ( n43926 , n43924 , n43925 );
and ( n43927 , n43923 , n221463 );
nor ( n43928 , n43926 , n43927 );
nand ( n43929 , n43917 , n43928 );
not ( n43930 , n43929 );
not ( n221692 , n205518 );
not ( n221693 , n25508 );
or ( n43933 , n221692 , n221693 );
or ( n43934 , n25508 , n205518 );
nand ( n43935 , n43933 , n43934 );
buf ( n43936 , n37449 );
not ( n43937 , n43936 );
and ( n43938 , n43935 , n43937 );
not ( n43939 , n43935 );
and ( n43940 , n43939 , n43936 );
nor ( n221702 , n43938 , n43940 );
not ( n221703 , n221702 );
and ( n43943 , n43930 , n221703 );
and ( n43944 , n43929 , n221702 );
nor ( n43945 , n43943 , n43944 );
not ( n43946 , n43945 );
and ( n43947 , n43902 , n43946 );
and ( n43948 , n43901 , n43945 );
nor ( n43949 , n43947 , n43948 );
not ( n43950 , n43949 );
or ( n43951 , n43816 , n43950 );
not ( n43952 , n43949 );
nand ( n221714 , n43952 , n43814 );
nand ( n221715 , n43951 , n221714 );
not ( n43955 , n221715 );
not ( n43956 , n43955 );
and ( n43957 , n43728 , n43956 );
not ( n43958 , n43728 );
and ( n43959 , n43949 , n43815 );
not ( n43960 , n43949 );
and ( n43961 , n43960 , n43814 );
nor ( n43962 , n43959 , n43961 );
not ( n43963 , n43962 );
not ( n43964 , n43963 );
and ( n221726 , n43958 , n43964 );
nor ( n221727 , n43957 , n221726 );
not ( n43967 , n221727 );
buf ( n43968 , n31571 );
not ( n43969 , n43968 );
nand ( n43970 , n43967 , n43969 );
nand ( n43971 , n42970 , n42990 );
buf ( n43972 , RI19a952a0_2646);
nand ( n43973 , n25851 , n43972 );
not ( n43974 , RI1747b7c8_1134);
and ( n43975 , n43973 , n43974 );
not ( n43976 , n43973 );
buf ( n221738 , RI1747b7c8_1134);
and ( n221739 , n43976 , n221738 );
nor ( n43979 , n43975 , n221739 );
not ( n43980 , n43979 );
not ( n43981 , n33134 );
or ( n43982 , n43980 , n43981 );
not ( n43983 , n43979 );
nand ( n43984 , n43983 , n33140 );
nand ( n43985 , n43982 , n43984 );
and ( n43986 , n43985 , n214235 );
not ( n43987 , n43985 );
and ( n43988 , n43987 , n30689 );
nor ( n43989 , n43986 , n43988 );
not ( n43990 , n43989 );
and ( n43991 , n43971 , n43990 );
not ( n43992 , n43971 );
and ( n43993 , n43992 , n43989 );
nor ( n43994 , n43991 , n43993 );
not ( n43995 , n43994 );
not ( n43996 , n43849 );
not ( n43997 , n43996 );
not ( n43998 , n32708 );
and ( n43999 , n43997 , n43998 );
not ( n221761 , n39706 );
and ( n221762 , n221761 , n32708 );
nor ( n44002 , n43999 , n221762 );
not ( n44003 , n35787 );
and ( n44004 , n44002 , n44003 );
not ( n44005 , n44002 );
not ( n44006 , n36377 );
and ( n44007 , n44005 , n44006 );
nor ( n221769 , n44004 , n44007 );
buf ( n221770 , n221769 );
not ( n44010 , n221770 );
nand ( n44011 , n43989 , n42991 );
not ( n44012 , n44011 );
or ( n44013 , n44010 , n44012 );
or ( n221775 , n44011 , n221770 );
nand ( n221776 , n44013 , n221775 );
buf ( n44016 , n39312 );
not ( n221778 , n44016 );
buf ( n221779 , n205029 );
not ( n44019 , n221779 );
or ( n44020 , n221778 , n44019 );
not ( n44021 , n44016 );
nand ( n44022 , n30896 , n44021 );
nand ( n221784 , n44020 , n44022 );
and ( n221785 , n221784 , n205074 );
not ( n221786 , n221784 );
buf ( n221787 , n205068 );
and ( n44027 , n221786 , n221787 );
nor ( n44028 , n221785 , n44027 );
not ( n44029 , n44028 );
nand ( n44030 , n44029 , n42885 );
not ( n44031 , n44030 );
not ( n44032 , n204321 );
not ( n221794 , n30405 );
or ( n221795 , n44032 , n221794 );
not ( n44035 , n33891 );
or ( n44036 , n44035 , n204321 );
nand ( n44037 , n221795 , n44036 );
and ( n44038 , n44037 , n33886 );
not ( n44039 , n44037 );
not ( n44040 , n33886 );
and ( n44041 , n44039 , n44040 );
nor ( n44042 , n44038 , n44041 );
not ( n221804 , n44042 );
not ( n221805 , n221804 );
and ( n44045 , n44031 , n221805 );
and ( n221807 , n44030 , n221804 );
nor ( n221808 , n44045 , n221807 );
and ( n44048 , n221776 , n221808 );
not ( n44049 , n221776 );
not ( n44050 , n221808 );
and ( n44051 , n44049 , n44050 );
nor ( n44052 , n44048 , n44051 );
not ( n44053 , n44052 );
not ( n221815 , n41751 );
not ( n221816 , n35274 );
or ( n44056 , n221815 , n221816 );
or ( n44057 , n41751 , n35274 );
nand ( n44058 , n44056 , n44057 );
and ( n44059 , n44058 , n213041 );
not ( n44060 , n44058 );
not ( n44061 , n213041 );
and ( n221823 , n44060 , n44061 );
nor ( n221824 , n44059 , n221823 );
nand ( n44064 , n221824 , n42866 );
not ( n221826 , n44064 );
not ( n221827 , n25676 );
not ( n44067 , n221827 );
not ( n44068 , n37843 );
not ( n44069 , n38130 );
or ( n44070 , n44068 , n44069 );
or ( n44071 , n38130 , n37843 );
nand ( n44072 , n44070 , n44071 );
not ( n44073 , n44072 );
or ( n44074 , n44067 , n44073 );
or ( n221836 , n44072 , n38141 );
nand ( n221837 , n44074 , n221836 );
not ( n44077 , n221837 );
and ( n44078 , n221826 , n44077 );
and ( n44079 , n44064 , n221837 );
nor ( n44080 , n44078 , n44079 );
not ( n221842 , n29990 );
not ( n221843 , n36683 );
not ( n44083 , n42284 );
not ( n44084 , n44083 );
or ( n44085 , n221843 , n44084 );
or ( n44086 , n44083 , n36683 );
nand ( n44087 , n44085 , n44086 );
not ( n44088 , n44087 );
and ( n44089 , n221842 , n44088 );
and ( n44090 , n29990 , n44087 );
nor ( n221852 , n44089 , n44090 );
nand ( n221853 , n221852 , n220589 );
not ( n44093 , n221853 );
not ( n44094 , n32188 );
not ( n44095 , n42512 );
or ( n44096 , n44094 , n44095 );
or ( n44097 , n42512 , n32188 );
nand ( n44098 , n44096 , n44097 );
and ( n44099 , n44098 , n221604 );
not ( n44100 , n44098 );
and ( n44101 , n44100 , n43839 );
nor ( n44102 , n44099 , n44101 );
not ( n221864 , n44102 );
not ( n221865 , n221864 );
and ( n44105 , n44093 , n221865 );
and ( n44106 , n221853 , n221864 );
nor ( n44107 , n44105 , n44106 );
xor ( n44108 , n44080 , n44107 );
not ( n44109 , n41359 );
and ( n44110 , n30146 , n44109 );
not ( n221872 , n30146 );
and ( n221873 , n221872 , n219115 );
nor ( n44113 , n44110 , n221873 );
and ( n44114 , n44113 , n27716 );
not ( n44115 , n44113 );
and ( n44116 , n44115 , n27721 );
nor ( n44117 , n44114 , n44116 );
buf ( n44118 , n44117 );
not ( n221880 , n44118 );
not ( n221881 , n34561 );
buf ( n44121 , RI174a51e0_931);
buf ( n221883 , RI1740a938_1456);
not ( n221884 , n221883 );
not ( n44124 , RI173c1c48_1811);
not ( n44125 , n44124 );
or ( n44126 , n221884 , n44125 );
not ( n44127 , RI1740a938_1456);
buf ( n44128 , RI173c1c48_1811);
nand ( n44129 , n44127 , n44128 );
nand ( n221891 , n44126 , n44129 );
xor ( n221892 , n44121 , n221891 );
buf ( n44132 , RI173386c8_2166);
xor ( n44133 , n44132 , n33060 );
xnor ( n44134 , n44133 , n33056 );
xnor ( n44135 , n221892 , n44134 );
not ( n44136 , n44135 );
not ( n44137 , n44136 );
or ( n44138 , n221881 , n44137 );
not ( n44139 , n34561 );
nand ( n44140 , n44139 , n44135 );
nand ( n44141 , n44138 , n44140 );
not ( n44142 , n35947 );
not ( n44143 , RI173964a8_2023);
not ( n44144 , n44143 );
or ( n44145 , n44142 , n44144 );
not ( n44146 , RI173df198_1668);
nand ( n44147 , n44146 , n34605 );
nand ( n44148 , n44145 , n44147 );
not ( n44149 , RI17456c70_1313);
and ( n44150 , n44148 , n44149 );
not ( n44151 , n44148 );
and ( n44152 , n44151 , n41058 );
nor ( n44153 , n44150 , n44152 );
xor ( n44154 , n44153 , n36467 );
xor ( n221916 , n44154 , n43979 );
not ( n221917 , n221916 );
not ( n44157 , n221917 );
buf ( n44158 , n44157 );
and ( n44159 , n44141 , n44158 );
not ( n44160 , n44141 );
not ( n44161 , n44158 );
and ( n44162 , n44160 , n44161 );
nor ( n44163 , n44159 , n44162 );
not ( n44164 , n44163 );
nand ( n44165 , n220481 , n44164 );
not ( n44166 , n44165 );
or ( n221928 , n221880 , n44166 );
or ( n221929 , n44165 , n44118 );
nand ( n44169 , n221928 , n221929 );
xor ( n44170 , n44108 , n44169 );
not ( n44171 , n44170 );
or ( n44172 , n44053 , n44171 );
not ( n44173 , n44170 );
not ( n44174 , n44052 );
nand ( n44175 , n44173 , n44174 );
nand ( n44176 , n44172 , n44175 );
not ( n44177 , n44176 );
or ( n44178 , n43995 , n44177 );
or ( n221940 , n44176 , n43994 );
nand ( n221941 , n44178 , n221940 );
not ( n44181 , n37810 );
buf ( n44182 , RI17359008_2091);
not ( n44183 , n44182 );
not ( n44184 , n25626 );
or ( n44185 , n44183 , n44184 );
or ( n44186 , n25626 , n44182 );
nand ( n44187 , n44185 , n44186 );
and ( n44188 , n44187 , n37464 );
not ( n221950 , n44187 );
and ( n221951 , n221950 , n28877 );
nor ( n44191 , n44188 , n221951 );
not ( n44192 , n32402 );
not ( n44193 , n39336 );
and ( n44194 , n44192 , n44193 );
and ( n44195 , n32402 , n39336 );
nor ( n44196 , n44194 , n44195 );
and ( n221958 , n44196 , n34575 );
not ( n221959 , n44196 );
and ( n44199 , n221959 , n32442 );
nor ( n44200 , n221958 , n44199 );
nand ( n44201 , n44191 , n44200 );
not ( n44202 , n44201 );
or ( n44203 , n44181 , n44202 );
or ( n44204 , n44201 , n37810 );
nand ( n44205 , n44203 , n44204 );
not ( n44206 , n44205 );
not ( n44207 , n40314 );
not ( n44208 , n207296 );
not ( n221970 , n38435 );
or ( n221971 , n44208 , n221970 );
or ( n44211 , n38435 , n207296 );
nand ( n44212 , n221971 , n44211 );
not ( n44213 , n44212 );
and ( n44214 , n44207 , n44213 );
and ( n44215 , n40314 , n44212 );
nor ( n44216 , n44214 , n44215 );
not ( n221978 , n34004 );
not ( n221979 , n38267 );
not ( n44219 , n30888 );
or ( n221981 , n221979 , n44219 );
or ( n221982 , n30888 , n38267 );
nand ( n44222 , n221981 , n221982 );
not ( n44223 , n44222 );
and ( n44224 , n221978 , n44223 );
and ( n44225 , n34004 , n44222 );
nor ( n44226 , n44224 , n44225 );
not ( n44227 , n44226 );
nand ( n44228 , n44216 , n44227 );
not ( n44229 , n44228 );
not ( n44230 , n37906 );
and ( n44231 , n44229 , n44230 );
and ( n221993 , n44228 , n37906 );
nor ( n221994 , n44231 , n221993 );
not ( n44234 , n221994 );
or ( n44235 , n44206 , n44234 );
or ( n44236 , n44205 , n221994 );
nand ( n44237 , n44235 , n44236 );
not ( n44238 , n40413 );
not ( n44239 , n44238 );
xor ( n222001 , n29821 , n44239 );
xnor ( n222002 , n222001 , n41878 );
not ( n44242 , n222002 );
not ( n44243 , n37782 );
nand ( n44244 , n44242 , n44243 );
not ( n44245 , n44244 );
not ( n44246 , n37958 );
and ( n44247 , n44245 , n44246 );
and ( n44248 , n44244 , n37958 );
nor ( n44249 , n44247 , n44248 );
not ( n222011 , n44249 );
and ( n222012 , n44237 , n222011 );
not ( n44252 , n44237 );
and ( n222014 , n44252 , n44249 );
nor ( n222015 , n222012 , n222014 );
not ( n44255 , n222015 );
not ( n222017 , n44255 );
not ( n222018 , n27931 );
not ( n44258 , n33849 );
or ( n44259 , n222018 , n44258 );
or ( n44260 , n33849 , n27931 );
nand ( n44261 , n44259 , n44260 );
not ( n222023 , n44261 );
not ( n222024 , n33812 );
or ( n44264 , n222023 , n222024 );
or ( n222026 , n33859 , n44261 );
nand ( n222027 , n44264 , n222026 );
not ( n44267 , n222027 );
not ( n44268 , n27725 );
not ( n44269 , n25502 );
not ( n44270 , n44269 );
or ( n222032 , n44268 , n44270 );
not ( n222033 , n25502 );
or ( n44273 , n222033 , n27725 );
nand ( n44274 , n222032 , n44273 );
and ( n44275 , n44274 , n43936 );
not ( n44276 , n44274 );
and ( n44277 , n44276 , n43937 );
nor ( n44278 , n44275 , n44277 );
not ( n44279 , n44278 );
nand ( n44280 , n44267 , n44279 );
not ( n44281 , n44280 );
not ( n44282 , n38038 );
and ( n222044 , n44281 , n44282 );
and ( n222045 , n44280 , n38038 );
nor ( n44285 , n222044 , n222045 );
not ( n44286 , n44285 );
xor ( n44287 , n33387 , n37106 );
xnor ( n44288 , n44287 , n38570 );
and ( n44289 , n31359 , n40057 );
not ( n44290 , n31359 );
and ( n44291 , n44290 , n40053 );
or ( n44292 , n44289 , n44291 );
not ( n222054 , n44292 );
not ( n222055 , n39320 );
or ( n44295 , n222054 , n222055 );
or ( n222057 , n39320 , n44292 );
nand ( n222058 , n44295 , n222057 );
buf ( n44298 , n222058 );
not ( n222060 , n44298 );
nand ( n222061 , n44288 , n222060 );
and ( n44301 , n222061 , n38209 );
not ( n44302 , n222061 );
not ( n44303 , n38209 );
and ( n44304 , n44302 , n44303 );
nor ( n44305 , n44301 , n44304 );
not ( n44306 , n44305 );
or ( n44307 , n44286 , n44306 );
not ( n44308 , n44305 );
not ( n44309 , n44285 );
nand ( n44310 , n44308 , n44309 );
nand ( n222072 , n44307 , n44310 );
not ( n222073 , n222072 );
and ( n44313 , n222017 , n222073 );
and ( n44314 , n44255 , n222072 );
nor ( n44315 , n44313 , n44314 );
buf ( n44316 , n44315 );
and ( n44317 , n221941 , n44316 );
not ( n44318 , n221941 );
not ( n222080 , n222015 );
not ( n222081 , n222072 );
not ( n44321 , n222081 );
or ( n44322 , n222080 , n44321 );
nand ( n44323 , n44255 , n222072 );
nand ( n44324 , n44322 , n44323 );
buf ( n44325 , n44324 );
and ( n44326 , n44318 , n44325 );
nor ( n44327 , n44317 , n44326 );
not ( n44328 , n204381 );
not ( n222090 , n37123 );
or ( n222091 , n44328 , n222090 );
nand ( n44331 , n37128 , n204377 );
nand ( n44332 , n222091 , n44331 );
buf ( n44333 , n34299 );
buf ( n44334 , n44333 );
and ( n44335 , n44332 , n44334 );
not ( n44336 , n44332 );
not ( n44337 , n44333 );
buf ( n44338 , n44337 );
and ( n44339 , n44336 , n44338 );
nor ( n44340 , n44335 , n44339 );
not ( n222102 , n44340 );
not ( n222103 , n33199 );
not ( n44343 , n25771 );
or ( n44344 , n222103 , n44343 );
or ( n44345 , n25771 , n33199 );
nand ( n44346 , n44344 , n44345 );
buf ( n44347 , n33362 );
buf ( n44348 , n44347 );
and ( n44349 , n44346 , n44348 );
not ( n44350 , n44346 );
buf ( n44351 , n33366 );
buf ( n44352 , n44351 );
and ( n44353 , n44350 , n44352 );
nor ( n44354 , n44349 , n44353 );
nand ( n222116 , n222102 , n44354 );
not ( n222117 , n222116 );
xor ( n44357 , n35739 , n30200 );
xnor ( n44358 , n44357 , n32916 );
not ( n44359 , n44358 );
not ( n44360 , n44359 );
or ( n222122 , n222117 , n44360 );
or ( n222123 , n44359 , n222116 );
nand ( n44363 , n222122 , n222123 );
not ( n222125 , n44363 );
not ( n222126 , n220493 );
not ( n44366 , n35923 );
or ( n44367 , n222126 , n44366 );
not ( n44368 , n220493 );
nand ( n44369 , n44368 , n43340 );
nand ( n44370 , n44367 , n44369 );
not ( n44371 , n44370 );
not ( n222133 , n41395 );
and ( n222134 , n44371 , n222133 );
and ( n44374 , n44370 , n41395 );
nor ( n222136 , n222134 , n44374 );
not ( n222137 , n222136 );
not ( n44377 , n36445 );
not ( n44378 , n26260 );
not ( n44379 , n44378 );
or ( n44380 , n44377 , n44379 );
or ( n44381 , n44378 , n36445 );
nand ( n44382 , n44380 , n44381 );
and ( n44383 , n44382 , n26310 );
not ( n44384 , n44382 );
and ( n222146 , n44384 , n26318 );
nor ( n222147 , n44383 , n222146 );
nand ( n44387 , n222137 , n222147 );
not ( n44388 , n44387 );
buf ( n44389 , n29843 );
not ( n44390 , n44389 );
buf ( n44391 , RI17406ae0_1475);
xor ( n44392 , n44391 , n35540 );
xor ( n44393 , n44392 , n35547 );
not ( n44394 , n44393 );
or ( n44395 , n44390 , n44394 );
or ( n44396 , n44393 , n44389 );
nand ( n222158 , n44395 , n44396 );
not ( n222159 , n40414 );
and ( n44399 , n222158 , n222159 );
not ( n222161 , n222158 );
and ( n222162 , n222161 , n44239 );
nor ( n44402 , n44399 , n222162 );
not ( n44403 , n44402 );
and ( n44404 , n44388 , n44403 );
and ( n44405 , n44387 , n44402 );
nor ( n44406 , n44404 , n44405 );
not ( n44407 , n44406 );
not ( n44408 , n32291 );
not ( n44409 , n37260 );
or ( n44410 , n44408 , n44409 );
not ( n44411 , n32291 );
not ( n44412 , n37260 );
nand ( n44413 , n44411 , n44412 );
nand ( n222175 , n44410 , n44413 );
and ( n222176 , n222175 , n39361 );
not ( n44416 , n222175 );
not ( n44417 , n217118 );
not ( n44418 , n38367 );
or ( n44419 , n44417 , n44418 );
or ( n44420 , n217118 , n38367 );
nand ( n44421 , n44419 , n44420 );
xnor ( n222183 , n44421 , n39349 );
buf ( n222184 , n222183 );
and ( n44424 , n44416 , n222184 );
nor ( n44425 , n222176 , n44424 );
not ( n44426 , n32230 );
not ( n44427 , n37346 );
or ( n222189 , n44426 , n44427 );
not ( n222190 , n32230 );
nand ( n44430 , n222190 , n43837 );
nand ( n44431 , n222189 , n44430 );
xnor ( n44432 , n44431 , n37352 );
nand ( n44433 , n44425 , n44432 );
not ( n44434 , n41258 );
not ( n44435 , n34024 );
not ( n44436 , n41303 );
or ( n44437 , n44435 , n44436 );
not ( n44438 , n34024 );
nand ( n44439 , n44438 , n219052 );
nand ( n222201 , n44437 , n44439 );
not ( n222202 , n222201 );
or ( n44442 , n44434 , n222202 );
or ( n222204 , n41258 , n222201 );
nand ( n222205 , n44442 , n222204 );
buf ( n44445 , n222205 );
xnor ( n44446 , n44433 , n44445 );
not ( n44447 , n44446 );
or ( n44448 , n44407 , n44447 );
or ( n44449 , n44446 , n44406 );
nand ( n44450 , n44448 , n44449 );
not ( n44451 , n34630 );
not ( n44452 , n43936 );
or ( n44453 , n44451 , n44452 );
or ( n44454 , n43936 , n34630 );
nand ( n222216 , n44453 , n44454 );
and ( n222217 , n222216 , n37455 );
not ( n44457 , n222216 );
buf ( n44458 , n32729 );
and ( n44459 , n44457 , n44458 );
nor ( n44460 , n222217 , n44459 );
buf ( n44461 , n35526 );
not ( n44462 , n44461 );
not ( n44463 , n33957 );
or ( n44464 , n44462 , n44463 );
not ( n44465 , n44461 );
nand ( n44466 , n44465 , n33954 );
nand ( n222228 , n44464 , n44466 );
xor ( n222229 , n222228 , n31344 );
nand ( n44469 , n44460 , n222229 );
not ( n44470 , n44469 );
not ( n44471 , n29815 );
xor ( n44472 , n26461 , n44471 );
xnor ( n44473 , n44472 , n36710 );
not ( n44474 , n44473 );
or ( n44475 , n44470 , n44474 );
or ( n44476 , n44473 , n44469 );
nand ( n44477 , n44475 , n44476 );
and ( n44478 , n44450 , n44477 );
not ( n222240 , n44450 );
not ( n222241 , n44477 );
and ( n44481 , n222240 , n222241 );
nor ( n44482 , n44478 , n44481 );
not ( n44483 , n39902 );
not ( n44484 , n38140 );
or ( n44485 , n44483 , n44484 );
or ( n44486 , n221827 , n39902 );
nand ( n222248 , n44485 , n44486 );
and ( n222249 , n222248 , n25683 );
not ( n44489 , n222248 );
and ( n222251 , n44489 , n25684 );
nor ( n222252 , n222249 , n222251 );
not ( n44492 , n29608 );
and ( n44493 , n35356 , n44492 );
not ( n44494 , n35356 );
and ( n44495 , n44494 , n29608 );
nor ( n44496 , n44493 , n44495 );
and ( n44497 , n44496 , n207409 );
not ( n44498 , n44496 );
and ( n44499 , n44498 , n29647 );
nor ( n44500 , n44497 , n44499 );
nand ( n44501 , n222252 , n44500 );
not ( n44502 , n44501 );
not ( n44503 , n40412 );
not ( n222265 , n29519 );
or ( n222266 , n44503 , n222265 );
not ( n44506 , n40412 );
nand ( n44507 , n44506 , n29525 );
nand ( n222269 , n222266 , n44507 );
and ( n222270 , n222269 , n29567 );
not ( n44510 , n222269 );
and ( n44511 , n44510 , n207325 );
nor ( n44512 , n222270 , n44511 );
not ( n44513 , n44512 );
not ( n44514 , n44513 );
and ( n44515 , n44502 , n44514 );
and ( n44516 , n44501 , n44513 );
nor ( n44517 , n44515 , n44516 );
not ( n44518 , n44517 );
xor ( n44519 , n29686 , n34700 );
xor ( n222281 , n44519 , n36859 );
not ( n222282 , n222281 );
not ( n44522 , n44354 );
nand ( n44523 , n44358 , n44522 );
not ( n44524 , n44523 );
or ( n44525 , n222282 , n44524 );
not ( n44526 , n44354 );
nand ( n44527 , n44526 , n44358 );
or ( n44528 , n44527 , n222281 );
nand ( n44529 , n44525 , n44528 );
not ( n44530 , n44529 );
or ( n44531 , n44518 , n44530 );
or ( n222293 , n44529 , n44517 );
nand ( n222294 , n44531 , n222293 );
and ( n44534 , n44482 , n222294 );
not ( n44535 , n44482 );
not ( n44536 , n222294 );
and ( n44537 , n44535 , n44536 );
nor ( n44538 , n44534 , n44537 );
buf ( n44539 , n44538 );
not ( n222301 , n44539 );
not ( n222302 , n222301 );
or ( n44542 , n222125 , n222302 );
not ( n222304 , n44363 );
nand ( n222305 , n222304 , n44539 );
nand ( n44545 , n44542 , n222305 );
not ( n44546 , n208623 );
not ( n44547 , n36455 );
or ( n44548 , n44546 , n44547 );
not ( n44549 , n208623 );
nand ( n44550 , n44549 , n36456 );
nand ( n44551 , n44548 , n44550 );
and ( n44552 , n44551 , n39212 );
not ( n222314 , n44551 );
and ( n222315 , n222314 , n39211 );
nor ( n44555 , n44552 , n222315 );
not ( n44556 , n44555 );
not ( n44557 , n44556 );
not ( n44558 , n33063 );
not ( n44559 , n36812 );
or ( n44560 , n44558 , n44559 );
or ( n44561 , n36812 , n33063 );
nand ( n44562 , n44560 , n44561 );
and ( n222324 , n39023 , n44562 );
not ( n222325 , n39023 );
not ( n44565 , n44562 );
and ( n222327 , n222325 , n44565 );
nor ( n222328 , n222324 , n222327 );
not ( n44568 , n222328 );
not ( n44569 , n33868 );
not ( n44570 , n205219 );
or ( n44571 , n44569 , n44570 );
not ( n44572 , n33868 );
nand ( n44573 , n44572 , n205220 );
nand ( n44574 , n44571 , n44573 );
and ( n44575 , n44574 , n43913 );
not ( n44576 , n44574 );
and ( n44577 , n44576 , n43910 );
nor ( n222339 , n44575 , n44577 );
nand ( n222340 , n44568 , n222339 );
not ( n44580 , n222340 );
or ( n44581 , n44557 , n44580 );
or ( n44582 , n222340 , n44556 );
nand ( n44583 , n44581 , n44582 );
not ( n44584 , n44583 );
not ( n44585 , n30005 );
not ( n44586 , n35888 );
or ( n44587 , n44585 , n44586 );
not ( n222349 , n30005 );
nand ( n222350 , n222349 , n35882 );
nand ( n44590 , n44587 , n222350 );
and ( n44591 , n44590 , n42391 );
not ( n44592 , n44590 );
and ( n44593 , n44592 , n42394 );
nor ( n44594 , n44591 , n44593 );
not ( n44595 , n38340 );
not ( n222357 , n32322 );
or ( n222358 , n44595 , n222357 );
not ( n44598 , n38340 );
nand ( n44599 , n44598 , n37900 );
nand ( n44600 , n222358 , n44599 );
and ( n44601 , n44600 , n220574 );
not ( n44602 , n44600 );
and ( n44603 , n44602 , n37397 );
nor ( n44604 , n44601 , n44603 );
nand ( n44605 , n44594 , n44604 );
not ( n222367 , n44605 );
not ( n222368 , n39696 );
not ( n44608 , n30756 );
or ( n222370 , n222368 , n44608 );
not ( n222371 , n39696 );
nand ( n44611 , n222371 , n30769 );
nand ( n44612 , n222370 , n44611 );
and ( n44613 , n44612 , n39480 );
not ( n44614 , n44612 );
not ( n44615 , n39480 );
and ( n44616 , n44614 , n44615 );
nor ( n44617 , n44613 , n44616 );
not ( n44618 , n44617 );
not ( n44619 , n44618 );
and ( n44620 , n222367 , n44619 );
and ( n222382 , n44605 , n44618 );
nor ( n222383 , n44620 , n222382 );
not ( n44623 , n222383 );
or ( n44624 , n44584 , n44623 );
or ( n44625 , n222383 , n44583 );
nand ( n44626 , n44624 , n44625 );
not ( n44627 , n44626 );
not ( n44628 , n44627 );
xor ( n44629 , n26450 , n29815 );
xnor ( n44630 , n44629 , n36710 );
not ( n222392 , n44630 );
not ( n222393 , n42956 );
not ( n44633 , n222393 );
not ( n44634 , n44633 );
not ( n222396 , n35997 );
not ( n222397 , n39246 );
or ( n44637 , n222396 , n222397 );
or ( n44638 , n39246 , n35997 );
nand ( n44639 , n44637 , n44638 );
not ( n44640 , n44639 );
or ( n222402 , n44634 , n44640 );
buf ( n222403 , n44633 );
or ( n44643 , n44639 , n222403 );
nand ( n44644 , n222402 , n44643 );
not ( n44645 , n44644 );
nand ( n44646 , n222392 , n44645 );
not ( n44647 , n44646 );
and ( n44648 , n32375 , n36187 );
not ( n44649 , n32375 );
and ( n44650 , n44649 , n36188 );
or ( n222412 , n44648 , n44650 );
not ( n222413 , n33525 );
xnor ( n44653 , n222412 , n222413 );
not ( n44654 , n44653 );
not ( n44655 , n44654 );
and ( n44656 , n44647 , n44655 );
and ( n44657 , n44646 , n44654 );
nor ( n222419 , n44656 , n44657 );
not ( n222420 , n222419 );
not ( n44660 , n222420 );
or ( n44661 , n44628 , n44660 );
nand ( n44662 , n222419 , n44626 );
nand ( n44663 , n44661 , n44662 );
not ( n44664 , n30553 );
not ( n44665 , n27802 );
or ( n44666 , n44664 , n44665 );
not ( n44667 , n30553 );
nand ( n222429 , n44667 , n27801 );
nand ( n222430 , n44666 , n222429 );
and ( n44670 , n222430 , n38771 );
not ( n44671 , n222430 );
and ( n44672 , n44671 , n38775 );
nor ( n44673 , n44670 , n44672 );
not ( n222435 , n44673 );
not ( n222436 , n222435 );
not ( n44676 , n222436 );
not ( n44677 , n25556 );
not ( n222439 , n36663 );
or ( n222440 , n44677 , n222439 );
or ( n44680 , n25556 , n36663 );
nand ( n222442 , n222440 , n44680 );
not ( n222443 , n206537 );
not ( n44683 , n222443 );
and ( n44684 , n222442 , n44683 );
not ( n44685 , n222442 );
not ( n44686 , n44683 );
and ( n44687 , n44685 , n44686 );
nor ( n44688 , n44684 , n44687 );
not ( n44689 , n44688 );
buf ( n44690 , n29117 );
not ( n44691 , n44690 );
not ( n44692 , n32586 );
not ( n222454 , n28502 );
or ( n222455 , n44692 , n222454 );
or ( n44695 , n28502 , n32586 );
nand ( n44696 , n222455 , n44695 );
not ( n44697 , n44696 );
and ( n44698 , n44691 , n44697 );
and ( n44699 , n44690 , n44696 );
nor ( n44700 , n44698 , n44699 );
not ( n222462 , n44700 );
nand ( n222463 , n44689 , n222462 );
not ( n44703 , n222463 );
or ( n44704 , n44676 , n44703 );
or ( n44705 , n222463 , n222436 );
nand ( n44706 , n44704 , n44705 );
not ( n44707 , n44706 );
not ( n44708 , n44707 );
not ( n222470 , n41713 );
buf ( n222471 , RI17460d38_1264);
xor ( n44711 , n222471 , n28138 );
xnor ( n44712 , n44711 , n28145 );
not ( n44713 , n44712 );
or ( n44714 , n222470 , n44713 );
not ( n44715 , n41713 );
nand ( n44716 , n44715 , n28146 );
nand ( n222478 , n44714 , n44716 );
and ( n222479 , n222478 , n35275 );
not ( n44719 , n222478 );
not ( n44720 , n35275 );
and ( n44721 , n44719 , n44720 );
nor ( n44722 , n222479 , n44721 );
not ( n44723 , n44722 );
buf ( n44724 , RI17407b48_1470);
not ( n222486 , n44724 );
not ( n222487 , n25762 );
or ( n44727 , n222486 , n222487 );
not ( n44728 , n44724 );
nand ( n44729 , n44728 , n25765 );
nand ( n44730 , n44727 , n44729 );
and ( n44731 , n44730 , n34331 );
not ( n44732 , n44730 );
and ( n44733 , n44732 , n34328 );
nor ( n44734 , n44731 , n44733 );
nand ( n222496 , n44723 , n44734 );
not ( n222497 , n222496 );
not ( n44737 , n37602 );
not ( n44738 , n35481 );
or ( n44739 , n44737 , n44738 );
or ( n44740 , n35481 , n37602 );
nand ( n44741 , n44739 , n44740 );
and ( n44742 , n44741 , n31137 );
not ( n222504 , n44741 );
and ( n222505 , n222504 , n29694 );
nor ( n44745 , n44742 , n222505 );
not ( n44746 , n44745 );
not ( n44747 , n44746 );
and ( n44748 , n222497 , n44747 );
and ( n44749 , n222496 , n44746 );
nor ( n44750 , n44748 , n44749 );
not ( n222512 , n44750 );
not ( n222513 , n222512 );
or ( n44753 , n44708 , n222513 );
nand ( n44754 , n44750 , n44706 );
nand ( n44755 , n44753 , n44754 );
and ( n44756 , n44663 , n44755 );
not ( n44757 , n44663 );
not ( n44758 , n44755 );
and ( n44759 , n44757 , n44758 );
nor ( n44760 , n44756 , n44759 );
not ( n44761 , n44760 );
and ( n44762 , n44545 , n44761 );
not ( n222524 , n44545 );
not ( n222525 , n44761 );
and ( n44765 , n222524 , n222525 );
nor ( n44766 , n44762 , n44765 );
not ( n44767 , n44766 );
nand ( n44768 , n44327 , n44767 );
or ( n44769 , n43970 , n44768 );
not ( n222531 , n35427 );
buf ( n222532 , n222531 );
not ( n222533 , n222532 );
nor ( n222534 , n43967 , n222533 );
nand ( n44774 , n222534 , n44768 );
nand ( n222536 , n39767 , n42337 );
nand ( n222537 , n44769 , n44774 , n222536 );
buf ( n44777 , n222537 );
not ( n44778 , n35551 );
buf ( n44779 , n40523 );
not ( n44780 , n44779 );
or ( n44781 , n44778 , n44780 );
not ( n44782 , n35551 );
nand ( n44783 , n44782 , n41040 );
nand ( n44784 , n44781 , n44783 );
buf ( n44785 , n40569 );
and ( n44786 , n44784 , n44785 );
not ( n222548 , n44784 );
buf ( n222549 , n40564 );
and ( n44789 , n222548 , n222549 );
nor ( n44790 , n44786 , n44789 );
not ( n44791 , n44790 );
not ( n44792 , n208497 );
not ( n44793 , n31637 );
or ( n44794 , n44792 , n44793 );
or ( n222556 , n31637 , n208497 );
nand ( n222557 , n44794 , n222556 );
and ( n44797 , n222557 , n37506 );
not ( n44798 , n222557 );
and ( n44799 , n44798 , n37507 );
nor ( n44800 , n44797 , n44799 );
nand ( n44801 , n44791 , n44800 );
not ( n44802 , n44801 );
not ( n44803 , n33292 );
not ( n44804 , n36414 );
or ( n222566 , n44803 , n44804 );
not ( n222567 , n33292 );
nand ( n44807 , n222567 , n35021 );
nand ( n44808 , n222566 , n44807 );
xor ( n44809 , n44808 , n26047 );
not ( n44810 , n44809 );
not ( n44811 , n44810 );
and ( n44812 , n44802 , n44811 );
and ( n44813 , n44801 , n44810 );
nor ( n44814 , n44812 , n44813 );
not ( n222576 , n44814 );
not ( n222577 , n29721 );
not ( n44817 , n39850 );
or ( n222579 , n222577 , n44817 );
or ( n222580 , n39850 , n29721 );
nand ( n44820 , n222579 , n222580 );
and ( n222582 , n44820 , n39845 );
not ( n222583 , n44820 );
buf ( n44823 , n41797 );
and ( n222585 , n222583 , n44823 );
nor ( n222586 , n222582 , n222585 );
not ( n44826 , n222586 );
not ( n222588 , n44826 );
not ( n222589 , n26222 );
not ( n44829 , n34575 );
not ( n44830 , n38854 );
and ( n44831 , n44829 , n44830 );
and ( n44832 , n34575 , n38854 );
nor ( n44833 , n44831 , n44832 );
and ( n44834 , n222589 , n44833 );
not ( n222596 , n222589 );
not ( n222597 , n44833 );
and ( n44837 , n222596 , n222597 );
nor ( n222599 , n44834 , n44837 );
not ( n222600 , n222599 );
not ( n44840 , n38783 );
not ( n222602 , n204830 );
and ( n222603 , n44840 , n222602 );
and ( n44843 , n37464 , n204830 );
nor ( n44844 , n222603 , n44843 );
and ( n44845 , n44844 , n211807 );
not ( n44846 , n44844 );
and ( n44847 , n44846 , n37472 );
nor ( n44848 , n44845 , n44847 );
not ( n44849 , n44848 );
nand ( n44850 , n222600 , n44849 );
not ( n44851 , n44850 );
or ( n44852 , n222588 , n44851 );
or ( n222614 , n44850 , n44826 );
nand ( n222615 , n44852 , n222614 );
not ( n44855 , n222615 );
not ( n44856 , n36211 );
not ( n44857 , RI173e9260_1619);
not ( n44858 , n29981 );
xor ( n44859 , n44857 , n44858 );
xnor ( n44860 , n44859 , n207749 );
not ( n222622 , n44860 );
or ( n222623 , n44856 , n222622 );
or ( n44863 , n29989 , n36211 );
nand ( n222625 , n222623 , n44863 );
and ( n222626 , n222625 , n28340 );
not ( n44866 , n222625 );
not ( n222628 , n28340 );
and ( n222629 , n44866 , n222628 );
nor ( n44869 , n222626 , n222629 );
not ( n222631 , n38154 );
not ( n222632 , n34102 );
or ( n44872 , n222631 , n222632 );
or ( n44873 , n34102 , n38154 );
nand ( n44874 , n44872 , n44873 );
and ( n44875 , n44874 , n40170 );
not ( n44876 , n44874 );
and ( n44877 , n44876 , n40169 );
nor ( n44878 , n44875 , n44877 );
not ( n44879 , n44878 );
nand ( n44880 , n44869 , n44879 );
not ( n44881 , n44880 );
buf ( n222643 , n28555 );
not ( n222644 , n222643 );
not ( n44884 , RI17334528_2186);
not ( n44885 , n44884 );
not ( n44886 , n28593 );
not ( n44887 , n44886 );
not ( n44888 , n44887 );
or ( n44889 , n44885 , n44888 );
nand ( n44890 , n28594 , n36181 );
nand ( n44891 , n44889 , n44890 );
not ( n44892 , n44891 );
or ( n44893 , n222644 , n44892 );
or ( n222655 , n44891 , n28557 );
nand ( n222656 , n44893 , n222655 );
not ( n44896 , n222656 );
not ( n44897 , n44896 );
not ( n44898 , n44897 );
and ( n44899 , n44881 , n44898 );
and ( n44900 , n44880 , n44897 );
nor ( n44901 , n44899 , n44900 );
not ( n44902 , n44901 );
or ( n44903 , n44855 , n44902 );
or ( n44904 , n44901 , n222615 );
nand ( n44905 , n44903 , n44904 );
buf ( n222667 , n38130 );
not ( n222668 , n222667 );
not ( n44908 , n37869 );
buf ( n44909 , RI173fc6d0_1525);
not ( n44910 , n44909 );
not ( n44911 , RI173b3698_1881);
not ( n44912 , n44911 );
or ( n44913 , n44910 , n44912 );
not ( n44914 , RI173fc6d0_1525);
buf ( n44915 , RI173b3698_1881);
nand ( n44916 , n44914 , n44915 );
nand ( n44917 , n44913 , n44916 );
and ( n222679 , n44917 , n39414 );
not ( n222680 , n44917 );
and ( n44920 , n222680 , n39409 );
nor ( n44921 , n222679 , n44920 );
buf ( n44922 , RI19a91c40_2670);
nand ( n44923 , n25416 , n44922 );
buf ( n44924 , RI175298b8_637);
and ( n44925 , n44923 , n44924 );
not ( n222687 , n44923 );
not ( n222688 , RI175298b8_637);
and ( n44928 , n222687 , n222688 );
nor ( n44929 , n44925 , n44928 );
xor ( n44930 , n44921 , n44929 );
xnor ( n44931 , n44930 , n32617 );
buf ( n44932 , n44931 );
not ( n44933 , n44932 );
or ( n44934 , n44908 , n44933 );
or ( n44935 , n44932 , n37869 );
nand ( n44936 , n44934 , n44935 );
not ( n44937 , n44936 );
or ( n222699 , n222668 , n44937 );
buf ( n222700 , n38130 );
or ( n44940 , n44936 , n222700 );
nand ( n44941 , n222699 , n44940 );
buf ( n44942 , n44941 );
not ( n44943 , n44942 );
xor ( n44944 , n37976 , n34179 );
not ( n44945 , n34139 );
xnor ( n44946 , n44944 , n44945 );
not ( n44947 , n44946 );
nand ( n222709 , n44943 , n44947 );
buf ( n222710 , n37439 );
not ( n44950 , n222710 );
not ( n44951 , n31905 );
or ( n44952 , n44950 , n44951 );
or ( n44953 , n31905 , n222710 );
nand ( n44954 , n44952 , n44953 );
xor ( n44955 , n39707 , n44954 );
and ( n222717 , n222709 , n44955 );
not ( n222718 , n222709 );
not ( n44958 , n44955 );
and ( n222720 , n222718 , n44958 );
nor ( n222721 , n222717 , n222720 );
not ( n44961 , n222721 );
and ( n44962 , n44905 , n44961 );
not ( n44963 , n44905 );
and ( n44964 , n44963 , n222721 );
nor ( n44965 , n44962 , n44964 );
not ( n44966 , n37211 );
xor ( n222728 , n30271 , n44966 );
xor ( n222729 , n222728 , n204621 );
not ( n44969 , n222729 );
not ( n44970 , n44969 );
not ( n44971 , n40007 );
not ( n44972 , n25732 );
and ( n44973 , n44971 , n44972 );
buf ( n44974 , n40005 );
and ( n44975 , n44974 , n25732 );
nor ( n44976 , n44973 , n44975 );
not ( n44977 , n44976 );
not ( n44978 , n30608 );
or ( n222740 , n44977 , n44978 );
or ( n222741 , n30608 , n44976 );
nand ( n44981 , n222740 , n222741 );
not ( n44982 , n44981 );
not ( n44983 , n31327 );
buf ( n44984 , n35821 );
not ( n44985 , n44984 );
or ( n44986 , n44983 , n44985 );
not ( n44987 , n35821 );
not ( n44988 , n44987 );
or ( n44989 , n44988 , n31327 );
nand ( n44990 , n44986 , n44989 );
buf ( n222752 , n37526 );
not ( n222753 , n222752 );
not ( n44993 , n222753 );
and ( n44994 , n44990 , n44993 );
not ( n44995 , n44990 );
and ( n44996 , n44995 , n222753 );
nor ( n44997 , n44994 , n44996 );
not ( n44998 , n44997 );
nand ( n44999 , n44982 , n44998 );
not ( n222761 , n44999 );
or ( n222762 , n44970 , n222761 );
or ( n45002 , n44999 , n44969 );
nand ( n45003 , n222762 , n45002 );
not ( n45004 , n45003 );
and ( n45005 , n44790 , n44809 );
buf ( n45006 , n36932 );
xor ( n45007 , n45006 , n37746 );
xnor ( n45008 , n45007 , n32240 );
and ( n45009 , n45005 , n45008 );
not ( n45010 , n45005 );
not ( n45011 , n45008 );
and ( n222773 , n45010 , n45011 );
nor ( n222774 , n45009 , n222773 );
not ( n45014 , n222774 );
and ( n45015 , n45004 , n45014 );
and ( n45016 , n45003 , n222774 );
nor ( n45017 , n45015 , n45016 );
and ( n45018 , n44965 , n45017 );
not ( n45019 , n44965 );
not ( n45020 , n45017 );
and ( n222782 , n45019 , n45020 );
nor ( n222783 , n45018 , n222782 );
not ( n45023 , n222783 );
not ( n45024 , n45023 );
or ( n45025 , n222576 , n45024 );
buf ( n45026 , n222783 );
not ( n45027 , n45026 );
or ( n45028 , n45027 , n44814 );
nand ( n222790 , n45025 , n45028 );
not ( n222791 , n34194 );
not ( n45031 , n32136 );
or ( n222793 , n222791 , n45031 );
or ( n222794 , n32136 , n34194 );
nand ( n45034 , n222793 , n222794 );
and ( n222796 , n45034 , n32183 );
not ( n222797 , n45034 );
and ( n45037 , n222797 , n32177 );
nor ( n45038 , n222796 , n45037 );
not ( n45039 , n45038 );
not ( n45040 , n45039 );
not ( n45041 , n26124 );
buf ( n45042 , n32766 );
not ( n45043 , n45042 );
or ( n45044 , n45041 , n45043 );
not ( n45045 , n32767 );
or ( n45046 , n45045 , n26124 );
nand ( n222808 , n45044 , n45046 );
and ( n222809 , n222808 , n39569 );
not ( n45049 , n222808 );
and ( n45050 , n45049 , n40480 );
nor ( n45051 , n222809 , n45050 );
not ( n45052 , n45051 );
buf ( n222814 , n205417 );
not ( n222815 , n222814 );
not ( n45055 , n205414 );
and ( n222817 , n222815 , n45055 );
and ( n222818 , n222814 , n205414 );
nor ( n45058 , n222817 , n222818 );
xor ( n222820 , n45058 , n39558 );
and ( n45060 , n222820 , n37303 );
not ( n45061 , n222820 );
and ( n45062 , n45061 , n36751 );
nor ( n45063 , n45060 , n45062 );
nand ( n45064 , n45052 , n45063 );
not ( n45065 , n45064 );
or ( n222827 , n45040 , n45065 );
or ( n222828 , n45064 , n45039 );
nand ( n45068 , n222827 , n222828 );
xor ( n45069 , n32298 , n222184 );
xnor ( n45070 , n45069 , n215032 );
not ( n45071 , n204811 );
not ( n45072 , n205068 );
or ( n45073 , n45071 , n45072 );
not ( n45074 , n204811 );
nand ( n45075 , n45074 , n205074 );
nand ( n45076 , n45073 , n45075 );
and ( n45077 , n45076 , n43757 );
not ( n222839 , n45076 );
and ( n222840 , n222839 , n43758 );
nor ( n45080 , n45077 , n222840 );
nand ( n45081 , n45070 , n45080 );
not ( n45082 , n45081 );
not ( n45083 , n205079 );
not ( n45084 , n32608 );
or ( n45085 , n45083 , n45084 );
or ( n45086 , n34759 , n205079 );
nand ( n45087 , n45085 , n45086 );
and ( n45088 , n45087 , n36414 );
not ( n45089 , n45087 );
and ( n222851 , n45089 , n36415 );
nor ( n222852 , n45088 , n222851 );
not ( n45092 , n222852 );
not ( n45093 , n45092 );
and ( n45094 , n45082 , n45093 );
and ( n45095 , n45081 , n45092 );
nor ( n45096 , n45094 , n45095 );
and ( n45097 , n45068 , n45096 );
not ( n222859 , n45068 );
not ( n222860 , n45096 );
and ( n45100 , n222859 , n222860 );
nor ( n45101 , n45097 , n45100 );
not ( n45102 , n45101 );
not ( n45103 , n30319 );
not ( n222865 , n41148 );
not ( n222866 , n222865 );
or ( n45106 , n45103 , n222866 );
not ( n45107 , n30319 );
not ( n45108 , n222865 );
nand ( n45109 , n45107 , n45108 );
nand ( n45110 , n45106 , n45109 );
not ( n45111 , n218917 );
and ( n45112 , n45110 , n45111 );
not ( n45113 , n45110 );
not ( n45114 , n37120 );
and ( n45115 , n45113 , n45114 );
nor ( n222877 , n45112 , n45115 );
not ( n222878 , n222877 );
not ( n45118 , n204952 );
not ( n45119 , n213777 );
or ( n45120 , n45118 , n45119 );
not ( n45121 , n204952 );
nand ( n222883 , n45121 , n36024 );
nand ( n222884 , n45120 , n222883 );
and ( n45124 , n222884 , n40862 );
not ( n222886 , n222884 );
and ( n222887 , n222886 , n221434 );
nor ( n45127 , n45124 , n222887 );
not ( n45128 , n45127 );
nand ( n45129 , n222878 , n45128 );
not ( n45130 , n45129 );
not ( n45131 , n40813 );
not ( n45132 , n38532 );
not ( n45133 , n33474 );
or ( n45134 , n45132 , n45133 );
nand ( n45135 , n33473 , n38528 );
nand ( n45136 , n45134 , n45135 );
not ( n222898 , n45136 );
and ( n222899 , n45131 , n222898 );
not ( n45139 , n43695 );
and ( n45140 , n45139 , n45136 );
nor ( n45141 , n222899 , n45140 );
not ( n45142 , n45141 );
not ( n45143 , n45142 );
and ( n45144 , n45130 , n45143 );
nand ( n45145 , n222878 , n45128 );
and ( n45146 , n45145 , n45142 );
nor ( n222908 , n45144 , n45146 );
not ( n222909 , n222908 );
buf ( n45149 , n31414 );
not ( n222911 , n45149 );
not ( n222912 , n39501 );
or ( n45152 , n222911 , n222912 );
not ( n45153 , n45149 );
nand ( n45154 , n45153 , n39319 );
nand ( n45155 , n45152 , n45154 );
and ( n45156 , n45155 , n39327 );
not ( n45157 , n45155 );
and ( n45158 , n45157 , n204825 );
nor ( n45159 , n45156 , n45158 );
not ( n222921 , n26479 );
not ( n222922 , n29815 );
or ( n45162 , n222921 , n222922 );
not ( n45163 , n26479 );
nand ( n45164 , n45163 , n36534 );
nand ( n45165 , n45162 , n45164 );
and ( n45166 , n45165 , n29856 );
not ( n45167 , n45165 );
and ( n222929 , n45167 , n29859 );
nor ( n222930 , n45166 , n222929 );
nand ( n45170 , n45159 , n222930 );
and ( n45171 , n33531 , n35357 );
not ( n45172 , n33531 );
and ( n45173 , n45172 , n38255 );
nor ( n45174 , n45171 , n45173 );
xnor ( n45175 , n35390 , n45174 );
and ( n45176 , n45170 , n45175 );
not ( n45177 , n45170 );
not ( n222939 , n45175 );
and ( n222940 , n45177 , n222939 );
nor ( n45180 , n45176 , n222940 );
not ( n45181 , n45180 );
or ( n45182 , n222909 , n45181 );
or ( n45183 , n45180 , n222908 );
nand ( n45184 , n45182 , n45183 );
not ( n45185 , n28222 );
not ( n45186 , n36238 );
or ( n45187 , n45185 , n45186 );
nand ( n222949 , n36243 , n28225 );
nand ( n222950 , n45187 , n222949 );
buf ( n45190 , RI173e5de0_1635);
not ( n45191 , n45190 );
not ( n45192 , RI1739cda8_1991);
not ( n45193 , n45192 );
or ( n45194 , n45191 , n45193 );
not ( n45195 , RI173e5de0_1635);
buf ( n45196 , RI1739cda8_1991);
nand ( n45197 , n45195 , n45196 );
nand ( n45198 , n45194 , n45197 );
buf ( n45199 , RI1745d8b8_1280);
and ( n222961 , n45198 , n45199 );
not ( n222962 , n45198 );
not ( n45202 , RI1745d8b8_1280);
and ( n45203 , n222962 , n45202 );
nor ( n45204 , n222961 , n45203 );
buf ( n45205 , RI19a843b0_2764);
nand ( n45206 , n206902 , n45205 );
buf ( n45207 , RI17506188_747);
and ( n222969 , n45206 , n45207 );
not ( n222970 , n45206 );
not ( n45210 , RI17506188_747);
and ( n45211 , n222970 , n45210 );
nor ( n45212 , n222969 , n45211 );
xor ( n45213 , n45204 , n45212 );
xnor ( n45214 , n45213 , n28305 );
buf ( n45215 , n45214 );
and ( n45216 , n222950 , n45215 );
not ( n45217 , n222950 );
not ( n45218 , n45214 );
and ( n45219 , n45217 , n45218 );
nor ( n222981 , n45216 , n45219 );
not ( n222982 , n222981 );
not ( n45222 , n42931 );
not ( n45223 , n43261 );
or ( n45224 , n45222 , n45223 );
not ( n45225 , n43260 );
not ( n45226 , n42931 );
nand ( n45227 , n45225 , n45226 );
nand ( n45228 , n45224 , n45227 );
not ( n45229 , n45228 );
buf ( n45230 , n40267 );
not ( n45231 , n45230 );
and ( n222993 , n45229 , n45231 );
not ( n222994 , n42675 );
and ( n45234 , n45228 , n222994 );
nor ( n222996 , n222993 , n45234 );
not ( n222997 , n222996 );
nand ( n45237 , n222982 , n222997 );
not ( n45238 , n45237 );
buf ( n45239 , RI173d15c0_1735);
xor ( n45240 , n45239 , n28877 );
xnor ( n45241 , n45240 , n25683 );
not ( n45242 , n45241 );
not ( n223004 , n45242 );
or ( n223005 , n45238 , n223004 );
or ( n45245 , n45242 , n45237 );
nand ( n45246 , n223005 , n45245 );
xor ( n45247 , n45184 , n45246 );
not ( n45248 , n45247 );
or ( n45249 , n45102 , n45248 );
not ( n45250 , n45247 );
not ( n45251 , n45101 );
nand ( n45252 , n45250 , n45251 );
nand ( n45253 , n45249 , n45252 );
not ( n223015 , n45253 );
not ( n223016 , n223015 );
and ( n45256 , n222790 , n223016 );
not ( n223018 , n222790 );
and ( n223019 , n45250 , n45251 );
not ( n45259 , n45250 );
and ( n45260 , n45259 , n45101 );
nor ( n45261 , n223019 , n45260 );
buf ( n45262 , n45261 );
and ( n45263 , n223018 , n45262 );
nor ( n45264 , n45256 , n45263 );
not ( n223026 , n45264 );
nor ( n223027 , n37652 , n28852 );
not ( n45267 , n223027 );
not ( n45268 , n37649 );
nand ( n45269 , n45268 , n28852 );
nand ( n45270 , n45267 , n45269 );
and ( n45271 , n45270 , n43073 );
not ( n45272 , n45270 );
and ( n223034 , n45272 , n220845 );
nor ( n223035 , n45271 , n223034 );
not ( n45275 , n223035 );
not ( n45276 , n32650 );
not ( n45277 , n221917 );
or ( n45278 , n45276 , n45277 );
not ( n45279 , n32650 );
not ( n45280 , n221916 );
not ( n45281 , n45280 );
nand ( n45282 , n45279 , n45281 );
nand ( n45283 , n45278 , n45282 );
buf ( n45284 , RI173fca18_1524);
not ( n45285 , n45284 );
not ( n45286 , RI173b39e0_1880);
not ( n223048 , n45286 );
or ( n223049 , n45285 , n223048 );
not ( n45289 , RI173fca18_1524);
buf ( n45290 , RI173b39e0_1880);
nand ( n45291 , n45289 , n45290 );
nand ( n45292 , n223049 , n45291 );
buf ( n45293 , RI173ab9e8_1919);
and ( n45294 , n45292 , n45293 );
not ( n223056 , n45292 );
not ( n223057 , RI173ab9e8_1919);
and ( n45297 , n223056 , n223057 );
nor ( n45298 , n45294 , n45297 );
buf ( n45299 , RI19aa8da0_2504);
nand ( n45300 , n33787 , n45299 );
buf ( n45301 , RI17498d00_991);
and ( n45302 , n45300 , n45301 );
not ( n223064 , n45300 );
not ( n223065 , RI17498d00_991);
and ( n45305 , n223064 , n223065 );
nor ( n45306 , n45302 , n45305 );
xor ( n45307 , n45298 , n45306 );
xor ( n45308 , n45307 , n30649 );
buf ( n45309 , n45308 );
not ( n45310 , n45309 );
and ( n45311 , n45283 , n45310 );
not ( n45312 , n45283 );
not ( n45313 , n45308 );
not ( n45314 , n45313 );
and ( n223076 , n45312 , n45314 );
nor ( n223077 , n45311 , n223076 );
nand ( n45317 , n45275 , n223077 );
not ( n45318 , n45317 );
not ( n45319 , n38347 );
not ( n45320 , n45319 );
xor ( n45321 , n40989 , n45320 );
not ( n45322 , n41520 );
xnor ( n45323 , n45321 , n45322 );
not ( n45324 , n45323 );
not ( n45325 , n45324 );
and ( n45326 , n45318 , n45325 );
and ( n223088 , n45317 , n45324 );
nor ( n223089 , n45326 , n223088 );
not ( n45329 , n223089 );
not ( n45330 , n45329 );
not ( n45331 , n206513 );
not ( n45332 , n205322 );
or ( n45333 , n45331 , n45332 );
or ( n45334 , n205322 , n206513 );
nand ( n45335 , n45333 , n45334 );
buf ( n45336 , n34381 );
and ( n223098 , n45335 , n45336 );
not ( n223099 , n45335 );
and ( n45339 , n223099 , n34391 );
nor ( n45340 , n223098 , n45339 );
not ( n45341 , n31616 );
not ( n45342 , n42372 );
or ( n223104 , n45341 , n45342 );
or ( n223105 , n42372 , n31616 );
nand ( n45345 , n223104 , n223105 );
and ( n223107 , n45345 , n26146 );
not ( n223108 , n45345 );
and ( n45348 , n223108 , n26149 );
nor ( n223110 , n223107 , n45348 );
nand ( n223111 , n45340 , n223110 );
not ( n45351 , n223111 );
not ( n45352 , n204484 );
not ( n45353 , n25927 );
or ( n45354 , n45352 , n45353 );
not ( n223116 , n25927 );
nand ( n223117 , n223116 , n204480 );
nand ( n45357 , n45354 , n223117 );
and ( n45358 , n45357 , n25978 );
not ( n45359 , n45357 );
and ( n45360 , n45359 , n25965 );
nor ( n45361 , n45358 , n45360 );
not ( n45362 , n45361 );
and ( n223124 , n45351 , n45362 );
and ( n223125 , n223111 , n45361 );
nor ( n45365 , n223124 , n223125 );
not ( n45366 , n45365 );
buf ( n45367 , RI1740d098_1444);
xor ( n45368 , n45367 , n28043 );
xnor ( n45369 , n45368 , n25868 );
not ( n45370 , n36455 );
not ( n45371 , n45370 );
xor ( n45372 , n30825 , n45371 );
not ( n45373 , n35107 );
xnor ( n45374 , n45372 , n45373 );
not ( n223136 , n45374 );
nand ( n223137 , n45369 , n223136 );
not ( n45377 , n31150 );
not ( n223139 , n42285 );
or ( n223140 , n45377 , n223139 );
or ( n45380 , n42285 , n31150 );
nand ( n45381 , n223140 , n45380 );
not ( n45382 , n29990 );
and ( n45383 , n45381 , n45382 );
not ( n45384 , n45381 );
and ( n45385 , n45384 , n29991 );
nor ( n45386 , n45383 , n45385 );
not ( n45387 , n45386 );
and ( n45388 , n223137 , n45387 );
not ( n45389 , n223137 );
and ( n45390 , n45389 , n45386 );
nor ( n223152 , n45388 , n45390 );
not ( n223153 , n223152 );
or ( n45393 , n45366 , n223153 );
or ( n223155 , n223152 , n45365 );
nand ( n223156 , n45393 , n223155 );
not ( n45396 , n29573 );
not ( n45397 , n38908 );
or ( n45398 , n45396 , n45397 );
not ( n45399 , n38911 );
or ( n45400 , n45399 , n29573 );
nand ( n45401 , n45398 , n45400 );
and ( n223163 , n45401 , n43469 );
not ( n223164 , n45401 );
not ( n45404 , n221233 );
not ( n223166 , n45404 );
not ( n223167 , n223166 );
and ( n45407 , n223164 , n223167 );
nor ( n45408 , n223163 , n45407 );
not ( n45409 , n36791 );
xor ( n45410 , n42612 , n42621 );
xnor ( n223172 , n45410 , n220226 );
not ( n223173 , n223172 );
or ( n45413 , n45409 , n223173 );
not ( n45414 , n36791 );
not ( n45415 , n223172 );
nand ( n45416 , n45414 , n45415 );
nand ( n45417 , n45413 , n45416 );
not ( n45418 , n44932 );
and ( n45419 , n45417 , n45418 );
not ( n45420 , n45417 );
and ( n45421 , n45420 , n44932 );
nor ( n45422 , n45419 , n45421 );
nand ( n223184 , n45408 , n45422 );
not ( n223185 , n223184 );
xor ( n45425 , n34673 , n204890 );
and ( n45426 , n45425 , n40218 );
not ( n45427 , n45425 );
and ( n45428 , n45427 , n40215 );
nor ( n223190 , n45426 , n45428 );
not ( n223191 , n223190 );
not ( n45431 , n223191 );
and ( n223193 , n223185 , n45431 );
and ( n223194 , n223184 , n223191 );
nor ( n45434 , n223193 , n223194 );
not ( n45435 , n45434 );
not ( n45436 , n38978 );
not ( n45437 , n204975 );
not ( n45438 , n45437 );
or ( n45439 , n45436 , n45438 );
or ( n45440 , n45437 , n38978 );
nand ( n45441 , n45439 , n45440 );
and ( n45442 , n36887 , n45441 );
not ( n45443 , n36887 );
not ( n223205 , n45441 );
and ( n223206 , n45443 , n223205 );
nor ( n45446 , n45442 , n223206 );
not ( n45447 , n45446 );
not ( n223209 , n37449 );
not ( n223210 , n42363 );
and ( n45450 , n223209 , n223210 );
and ( n45451 , n37449 , n42363 );
nor ( n45452 , n45450 , n45451 );
and ( n45453 , n45452 , n37458 );
not ( n45454 , n45452 );
and ( n45455 , n45454 , n37455 );
nor ( n45456 , n45453 , n45455 );
nand ( n45457 , n45447 , n45456 );
not ( n45458 , n37371 );
not ( n223220 , n222183 );
or ( n223221 , n45458 , n223220 );
nand ( n45461 , n39359 , n37367 );
nand ( n45462 , n223221 , n45461 );
not ( n45463 , n45462 );
buf ( n45464 , n38877 );
not ( n45465 , n45464 );
not ( n45466 , n45465 );
and ( n45467 , n45463 , n45466 );
not ( n45468 , n45464 );
and ( n223230 , n45462 , n45468 );
nor ( n223231 , n45467 , n223230 );
and ( n45471 , n45457 , n223231 );
not ( n45472 , n45457 );
not ( n45473 , n223231 );
and ( n45474 , n45472 , n45473 );
nor ( n45475 , n45471 , n45474 );
not ( n45476 , n45475 );
or ( n45477 , n45435 , n45476 );
or ( n45478 , n45475 , n45434 );
nand ( n223240 , n45477 , n45478 );
nand ( n223241 , n45323 , n223035 );
not ( n45481 , n223241 );
not ( n45482 , n29519 );
not ( n45483 , n35538 );
not ( n45484 , n40569 );
or ( n45485 , n45483 , n45484 );
nand ( n45486 , n40562 , n35535 );
nand ( n45487 , n45485 , n45486 );
not ( n45488 , n45487 );
or ( n45489 , n45482 , n45488 );
or ( n45490 , n45487 , n29519 );
nand ( n223252 , n45489 , n45490 );
not ( n223253 , n223252 );
and ( n45493 , n45481 , n223253 );
and ( n223255 , n223241 , n223252 );
nor ( n223256 , n45493 , n223255 );
and ( n45496 , n223240 , n223256 );
not ( n45497 , n223240 );
not ( n45498 , n223256 );
and ( n45499 , n45497 , n45498 );
nor ( n45500 , n45496 , n45499 );
and ( n45501 , n223156 , n45500 );
not ( n45502 , n223156 );
not ( n45503 , n45500 );
and ( n223265 , n45502 , n45503 );
nor ( n223266 , n45501 , n223265 );
not ( n45506 , n223266 );
not ( n45507 , n45506 );
not ( n45508 , n45507 );
or ( n45509 , n45330 , n45508 );
not ( n223271 , n45329 );
nand ( n223272 , n223271 , n45506 );
nand ( n45512 , n45509 , n223272 );
not ( n45513 , n39006 );
not ( n45514 , n28398 );
and ( n45515 , n45513 , n45514 );
and ( n45516 , n39006 , n28398 );
nor ( n45517 , n45515 , n45516 );
buf ( n45518 , n41855 );
xor ( n45519 , n45517 , n45518 );
not ( n45520 , n45519 );
not ( n45521 , n41405 );
buf ( n223283 , n25372 );
not ( n223284 , n223283 );
not ( n45524 , n30281 );
not ( n223286 , n45524 );
or ( n223287 , n223284 , n223286 );
or ( n45527 , n45524 , n223283 );
nand ( n45528 , n223287 , n45527 );
not ( n45529 , n45528 );
and ( n45530 , n45521 , n45529 );
not ( n45531 , n30247 );
and ( n45532 , n45531 , n45528 );
nor ( n45533 , n45530 , n45532 );
nand ( n45534 , n45520 , n45533 );
not ( n45535 , n45534 );
not ( n45536 , n32628 );
not ( n223298 , n45280 );
or ( n223299 , n45536 , n223298 );
or ( n45539 , n221917 , n32628 );
nand ( n45540 , n223299 , n45539 );
and ( n45541 , n45540 , n45314 );
not ( n45542 , n45540 );
and ( n45543 , n45542 , n45313 );
nor ( n45544 , n45541 , n45543 );
not ( n45545 , n45544 );
not ( n45546 , n45545 );
and ( n45547 , n45535 , n45546 );
and ( n45548 , n45534 , n45545 );
nor ( n223310 , n45547 , n45548 );
not ( n223311 , n223310 );
buf ( n45551 , RI19a8b700_2715);
nand ( n223313 , n25851 , n45551 );
buf ( n223314 , RI1746d8a8_1202);
and ( n45554 , n223313 , n223314 );
not ( n45555 , n223313 );
not ( n45556 , RI1746d8a8_1202);
and ( n45557 , n45555 , n45556 );
nor ( n45558 , n45554 , n45557 );
not ( n45559 , n45558 );
not ( n223321 , n25683 );
or ( n223322 , n45559 , n223321 );
or ( n45562 , n25683 , n45558 );
nand ( n45563 , n223322 , n45562 );
and ( n45564 , n45563 , n28878 );
not ( n45565 , n45563 );
and ( n45566 , n45565 , n28877 );
nor ( n45567 , n45564 , n45566 );
buf ( n223329 , n29595 );
not ( n223330 , n223329 );
not ( n45570 , n38911 );
or ( n45571 , n223330 , n45570 );
not ( n45572 , n38908 );
or ( n45573 , n45572 , n223329 );
nand ( n45574 , n45571 , n45573 );
and ( n45575 , n45574 , n43473 );
not ( n223337 , n45574 );
and ( n223338 , n223337 , n223167 );
nor ( n45578 , n45575 , n223338 );
not ( n45579 , n45578 );
nand ( n45580 , n45567 , n45579 );
not ( n45581 , n39694 );
not ( n45582 , n30756 );
or ( n45583 , n45581 , n45582 );
not ( n45584 , n39694 );
nand ( n45585 , n45584 , n30769 );
nand ( n45586 , n45583 , n45585 );
and ( n45587 , n45586 , n39481 );
not ( n45588 , n45586 );
and ( n45589 , n45588 , n44615 );
nor ( n45590 , n45587 , n45589 );
and ( n45591 , n45580 , n45590 );
not ( n45592 , n45580 );
not ( n45593 , n45590 );
and ( n223355 , n45592 , n45593 );
nor ( n223356 , n45591 , n223355 );
not ( n45596 , n223356 );
or ( n45597 , n223311 , n45596 );
or ( n45598 , n223356 , n223310 );
nand ( n45599 , n45597 , n45598 );
not ( n45600 , n39922 );
buf ( n45601 , n30674 );
not ( n45602 , n45601 );
not ( n45603 , n45602 );
not ( n45604 , n40619 );
or ( n45605 , n45603 , n45604 );
nand ( n45606 , n37865 , n45601 );
nand ( n223368 , n45605 , n45606 );
not ( n223369 , n223368 );
or ( n45609 , n45600 , n223369 );
or ( n45610 , n223368 , n39922 );
nand ( n45611 , n45609 , n45610 );
not ( n45612 , n45611 );
not ( n45613 , n34381 );
buf ( n45614 , n28765 );
and ( n45615 , n45614 , n34384 );
not ( n45616 , n45614 );
xor ( n45617 , n205303 , n205311 );
not ( n45618 , n205320 );
xnor ( n45619 , n45617 , n45618 );
and ( n223381 , n45616 , n45619 );
nor ( n223382 , n45615 , n223381 );
not ( n45622 , n223382 );
and ( n45623 , n45613 , n45622 );
and ( n45624 , n34381 , n223382 );
nor ( n45625 , n45623 , n45624 );
not ( n45626 , n45625 );
nand ( n45627 , n45612 , n45626 );
not ( n45628 , n29711 );
not ( n45629 , n34700 );
or ( n45630 , n45628 , n45629 );
or ( n45631 , n34700 , n29711 );
nand ( n223393 , n45630 , n45631 );
and ( n223394 , n223393 , n39845 );
not ( n45634 , n223393 );
and ( n223396 , n45634 , n44823 );
nor ( n223397 , n223394 , n223396 );
not ( n45637 , n223397 );
and ( n223399 , n45627 , n45637 );
not ( n223400 , n45627 );
and ( n45640 , n223400 , n223397 );
nor ( n45641 , n223399 , n45640 );
not ( n45642 , n45641 );
and ( n45643 , n45599 , n45642 );
not ( n45644 , n45599 );
and ( n45645 , n45644 , n45641 );
nor ( n223407 , n45643 , n45645 );
not ( n223408 , n205230 );
and ( n45648 , n25813 , n37169 );
not ( n45649 , n25813 );
and ( n45650 , n45649 , n38688 );
or ( n45651 , n45648 , n45650 );
not ( n45652 , n45651 );
and ( n45653 , n223408 , n45652 );
and ( n223415 , n205230 , n45651 );
nor ( n223416 , n45653 , n223415 );
not ( n45656 , n223416 );
not ( n45657 , n28875 );
not ( n45658 , n37652 );
or ( n45659 , n45657 , n45658 );
not ( n223421 , n28875 );
nand ( n223422 , n223421 , n37649 );
nand ( n45662 , n45659 , n223422 );
and ( n223424 , n45662 , n43073 );
not ( n223425 , n45662 );
and ( n45665 , n223425 , n220845 );
nor ( n45666 , n223424 , n45665 );
not ( n45667 , n45666 );
nand ( n45668 , n45656 , n45667 );
not ( n45669 , n45668 );
not ( n45670 , n45669 );
xor ( n45671 , n26236 , n43122 );
buf ( n45672 , n220543 );
xor ( n45673 , n45671 , n45672 );
not ( n45674 , n45673 );
or ( n223436 , n45670 , n45674 );
not ( n223437 , n45673 );
nand ( n45677 , n223437 , n45668 );
nand ( n45678 , n223436 , n45677 );
buf ( n45679 , n204580 );
not ( n45680 , n45679 );
not ( n45681 , n28381 );
or ( n45682 , n45680 , n45681 );
or ( n223444 , n28381 , n45679 );
nand ( n223445 , n45682 , n223444 );
and ( n45685 , n223445 , n30140 );
not ( n45686 , n223445 );
and ( n45687 , n45686 , n30137 );
nor ( n45688 , n45685 , n45687 );
not ( n45689 , n45688 );
not ( n45690 , n26396 );
not ( n45691 , n45690 );
xor ( n45692 , n45691 , n41040 );
buf ( n223454 , RI174022b0_1497);
xor ( n223455 , n223454 , n41049 );
xnor ( n45695 , n223455 , n41053 );
buf ( n45696 , n45695 );
xnor ( n45697 , n45692 , n45696 );
nand ( n45698 , n45689 , n45697 );
not ( n45699 , n45698 );
not ( n45700 , n37004 );
not ( n45701 , n41592 );
not ( n45702 , n45701 );
not ( n223464 , n45702 );
or ( n223465 , n45700 , n223464 );
or ( n45705 , n41593 , n37004 );
nand ( n223467 , n223465 , n45705 );
and ( n223468 , n223467 , n36093 );
not ( n45708 , n223467 );
and ( n45709 , n45708 , n44712 );
nor ( n45710 , n223468 , n45709 );
not ( n45711 , n45710 );
not ( n223473 , n45711 );
and ( n223474 , n45699 , n223473 );
not ( n45714 , n45688 );
nand ( n45715 , n45714 , n45697 );
and ( n45716 , n45715 , n45711 );
nor ( n45717 , n223474 , n45716 );
and ( n45718 , n45678 , n45717 );
not ( n45719 , n45678 );
not ( n45720 , n45717 );
and ( n45721 , n45719 , n45720 );
nor ( n45722 , n45718 , n45721 );
and ( n45723 , n223407 , n45722 );
not ( n223485 , n223407 );
not ( n223486 , n45722 );
and ( n45726 , n223485 , n223486 );
nor ( n45727 , n45723 , n45726 );
buf ( n45728 , n45727 );
xor ( n45729 , n45512 , n45728 );
not ( n45730 , n45729 );
nand ( n45731 , n223026 , n45730 );
not ( n45732 , n28567 );
not ( n45733 , n37398 );
or ( n45734 , n45732 , n45733 );
or ( n45735 , n37398 , n28567 );
nand ( n223497 , n45734 , n45735 );
and ( n223498 , n223497 , n30809 );
not ( n45738 , n223497 );
and ( n45739 , n45738 , n30810 );
nor ( n45740 , n223498 , n45739 );
not ( n45741 , n45740 );
not ( n223503 , n29973 );
buf ( n223504 , n204791 );
not ( n45744 , n223504 );
not ( n223506 , n45744 );
or ( n223507 , n223503 , n223506 );
or ( n45747 , n204792 , n29973 );
nand ( n223509 , n223507 , n45747 );
buf ( n223510 , n36309 );
not ( n45750 , n223510 );
and ( n45751 , n223509 , n45750 );
not ( n45752 , n223509 );
and ( n45753 , n45752 , n223510 );
nor ( n45754 , n45751 , n45753 );
nand ( n45755 , n45741 , n45754 );
not ( n45756 , n45755 );
not ( n45757 , n36688 );
and ( n223519 , n45756 , n45757 );
and ( n223520 , n45755 , n36688 );
nor ( n45760 , n223519 , n223520 );
buf ( n45761 , n45760 );
not ( n45762 , n45761 );
not ( n45763 , n36378 );
not ( n45764 , n34358 );
not ( n45765 , n219430 );
or ( n45766 , n45764 , n45765 );
nand ( n45767 , n37023 , n34354 );
nand ( n223529 , n45766 , n45767 );
buf ( n223530 , n41723 );
buf ( n45770 , n223530 );
and ( n45771 , n223529 , n45770 );
not ( n45772 , n223529 );
buf ( n45773 , n42348 );
not ( n223535 , n45773 );
not ( n223536 , n223535 );
and ( n45776 , n45772 , n223536 );
nor ( n45777 , n45771 , n45776 );
not ( n45778 , n45777 );
nand ( n45779 , n36382 , n45778 );
not ( n45780 , n45779 );
or ( n45781 , n45763 , n45780 );
not ( n45782 , n45777 );
nand ( n45783 , n45782 , n36382 );
or ( n45784 , n45783 , n36378 );
nand ( n223546 , n45781 , n45784 );
not ( n223547 , n223546 );
not ( n45787 , n36540 );
not ( n45788 , n39221 );
not ( n45789 , RI173ddaa0_1675);
not ( n45790 , n28396 );
xor ( n45791 , n45789 , n45790 );
xnor ( n45792 , n45791 , n28403 );
not ( n45793 , n45792 );
or ( n45794 , n45788 , n45793 );
or ( n45795 , n45792 , n39221 );
nand ( n45796 , n45794 , n45795 );
and ( n223558 , n45796 , n43262 );
not ( n223559 , n45796 );
not ( n45799 , n45225 );
and ( n223561 , n223559 , n45799 );
nor ( n223562 , n223558 , n223561 );
nand ( n45802 , n45787 , n223562 );
not ( n45803 , n45802 );
not ( n45804 , n36528 );
and ( n45805 , n45803 , n45804 );
not ( n45806 , n36540 );
nand ( n45807 , n45806 , n223562 );
and ( n45808 , n45807 , n36528 );
nor ( n45809 , n45805 , n45808 );
not ( n45810 , n45809 );
not ( n45811 , n36779 );
not ( n223573 , n42623 );
or ( n223574 , n45811 , n223573 );
not ( n45814 , n36779 );
nand ( n45815 , n45814 , n45415 );
nand ( n45816 , n223574 , n45815 );
buf ( n45817 , n44932 );
not ( n45818 , n45817 );
and ( n45819 , n45816 , n45818 );
not ( n45820 , n45816 );
and ( n45821 , n45820 , n45817 );
nor ( n223583 , n45819 , n45821 );
nand ( n223584 , n223583 , n36478 );
and ( n45824 , n223584 , n36459 );
not ( n45825 , n223584 );
and ( n45826 , n45825 , n36458 );
nor ( n45827 , n45824 , n45826 );
not ( n45828 , n45827 );
and ( n45829 , n45810 , n45828 );
and ( n45830 , n45809 , n45827 );
nor ( n45831 , n45829 , n45830 );
not ( n45832 , n45831 );
or ( n45833 , n223547 , n45832 );
or ( n223595 , n223546 , n45831 );
nand ( n223596 , n45833 , n223595 );
not ( n45836 , n36698 );
not ( n45837 , n45836 );
nand ( n45838 , n36687 , n45740 );
not ( n45839 , n45838 );
or ( n45840 , n45837 , n45839 );
or ( n45841 , n45838 , n45836 );
nand ( n223603 , n45840 , n45841 );
not ( n223604 , n223603 );
not ( n45844 , n31050 );
not ( n45845 , n34914 );
or ( n45846 , n45844 , n45845 );
nand ( n45847 , n34917 , n31046 );
nand ( n45848 , n45846 , n45847 );
not ( n45849 , n45524 );
not ( n45850 , n45849 );
and ( n45851 , n45848 , n45850 );
not ( n223613 , n45848 );
buf ( n223614 , n45849 );
not ( n45854 , n223614 );
not ( n45855 , n45854 );
and ( n45856 , n223613 , n45855 );
nor ( n45857 , n45851 , n45856 );
nand ( n45858 , n36666 , n45857 );
not ( n45859 , n45858 );
not ( n223621 , n36628 );
and ( n223622 , n45859 , n223621 );
and ( n45862 , n45858 , n36628 );
nor ( n45863 , n223622 , n45862 );
not ( n45864 , n45863 );
or ( n45865 , n223604 , n45864 );
or ( n223627 , n45863 , n223603 );
nand ( n223628 , n45865 , n223627 );
and ( n45868 , n223596 , n223628 );
not ( n223630 , n223596 );
not ( n223631 , n223628 );
and ( n45871 , n223630 , n223631 );
nor ( n45872 , n45868 , n45871 );
buf ( n45873 , n45872 );
not ( n45874 , n45873 );
or ( n45875 , n45762 , n45874 );
not ( n45876 , n45872 );
not ( n45877 , n45876 );
or ( n45878 , n45877 , n45761 );
nand ( n45879 , n45875 , n45878 );
and ( n45880 , n32142 , n33613 );
not ( n223642 , n32142 );
and ( n223643 , n223642 , n33618 );
nor ( n45883 , n45880 , n223643 );
not ( n45884 , n45883 );
not ( n45885 , n41520 );
or ( n45886 , n45884 , n45885 );
or ( n45887 , n41520 , n45883 );
nand ( n45888 , n45886 , n45887 );
not ( n223650 , n45888 );
not ( n223651 , n29121 );
not ( n45891 , n36262 );
or ( n223653 , n223651 , n45891 );
not ( n223654 , n29121 );
nand ( n45894 , n223654 , n210587 );
nand ( n45895 , n223653 , n45894 );
xor ( n45896 , n39395 , n38035 );
xnor ( n45897 , n45896 , n32516 );
buf ( n45898 , n45897 );
and ( n45899 , n45895 , n45898 );
not ( n223661 , n45895 );
and ( n223662 , n223661 , n39401 );
nor ( n45902 , n45899 , n223662 );
nand ( n45903 , n223650 , n45902 );
not ( n45904 , n45903 );
not ( n45905 , n32619 );
not ( n45906 , n45280 );
or ( n45907 , n45905 , n45906 );
or ( n223669 , n221917 , n32619 );
nand ( n223670 , n45907 , n223669 );
and ( n45910 , n223670 , n45308 );
not ( n45911 , n223670 );
and ( n45912 , n45911 , n45313 );
nor ( n45913 , n45910 , n45912 );
not ( n45914 , n45913 );
not ( n45915 , n45914 );
and ( n45916 , n45904 , n45915 );
and ( n45917 , n45903 , n45914 );
nor ( n223679 , n45916 , n45917 );
not ( n223680 , n223679 );
not ( n45920 , n223680 );
not ( n45921 , n36816 );
not ( n45922 , n42593 );
or ( n45923 , n45921 , n45922 );
or ( n45924 , n42593 , n36816 );
nand ( n45925 , n45923 , n45924 );
buf ( n45926 , n42624 );
not ( n45927 , n45926 );
and ( n45928 , n45925 , n45927 );
not ( n45929 , n45925 );
and ( n223691 , n45929 , n45926 );
nor ( n223692 , n45928 , n223691 );
not ( n45932 , n36006 );
buf ( n45933 , n39244 );
not ( n45934 , n45933 );
or ( n45935 , n45932 , n45934 );
not ( n45936 , n36006 );
nand ( n45937 , n45936 , n39250 );
nand ( n223699 , n45935 , n45937 );
and ( n223700 , n223699 , n44633 );
not ( n45940 , n223699 );
xor ( n45941 , n42950 , n42922 );
xnor ( n45942 , n45941 , n45226 );
not ( n45943 , n45942 );
not ( n45944 , n45943 );
and ( n45945 , n45940 , n45944 );
nor ( n45946 , n223700 , n45945 );
not ( n45947 , n45946 );
nand ( n45948 , n223692 , n45947 );
not ( n45949 , n45948 );
buf ( n223711 , n221403 );
xor ( n223712 , n28133 , n223711 );
xnor ( n45952 , n223712 , n40976 );
not ( n45953 , n45952 );
or ( n45954 , n45949 , n45953 );
or ( n45955 , n45952 , n45948 );
nand ( n45956 , n45954 , n45955 );
not ( n45957 , n45956 );
not ( n223719 , n45957 );
or ( n223720 , n45920 , n223719 );
nand ( n45960 , n45956 , n223679 );
nand ( n45961 , n223720 , n45960 );
xor ( n45962 , n32746 , n35754 );
xnor ( n45963 , n45962 , n36377 );
not ( n45964 , n35481 );
not ( n45965 , n40103 );
not ( n223727 , n37991 );
or ( n223728 , n45965 , n223727 );
or ( n45968 , n37991 , n40103 );
nand ( n223730 , n223728 , n45968 );
not ( n223731 , n223730 );
or ( n45971 , n45964 , n223731 );
or ( n45972 , n223730 , n38000 );
nand ( n45973 , n45971 , n45972 );
not ( n45974 , n45973 );
nand ( n223736 , n45963 , n45974 );
not ( n223737 , n41837 );
not ( n45977 , n43063 );
or ( n45978 , n223737 , n45977 );
or ( n45979 , n28906 , n41837 );
nand ( n45980 , n45978 , n45979 );
and ( n45981 , n45980 , n30943 );
not ( n45982 , n45980 );
and ( n45983 , n45982 , n30936 );
nor ( n45984 , n45981 , n45983 );
buf ( n223746 , n45984 );
xnor ( n223747 , n223736 , n223746 );
not ( n45987 , n223747 );
and ( n45988 , n45961 , n45987 );
not ( n45989 , n45961 );
and ( n45990 , n45989 , n223747 );
nor ( n223752 , n45988 , n45990 );
not ( n223753 , n223752 );
not ( n45993 , n219094 );
not ( n45994 , n25965 );
or ( n45995 , n45993 , n45994 );
nand ( n45996 , n25978 , n41330 );
nand ( n45997 , n45995 , n45996 );
and ( n45998 , n45997 , n25456 );
not ( n45999 , n45997 );
and ( n46000 , n45999 , n25457 );
nor ( n46001 , n45998 , n46000 );
not ( n46002 , n26013 );
not ( n223764 , n29175 );
or ( n223765 , n46002 , n223764 );
or ( n46005 , n29175 , n26013 );
nand ( n46006 , n223765 , n46005 );
and ( n46007 , n46006 , n33937 );
not ( n46008 , n46006 );
and ( n46009 , n46008 , n33936 );
nor ( n46010 , n46007 , n46009 );
not ( n46011 , n46010 );
nand ( n46012 , n46001 , n46011 );
not ( n46013 , n46012 );
not ( n223775 , n204612 );
not ( n223776 , n30137 );
or ( n46016 , n223775 , n223776 );
nand ( n46017 , n43577 , n204615 );
nand ( n46018 , n46016 , n46017 );
and ( n46019 , n46018 , n33957 );
not ( n46020 , n46018 );
and ( n46021 , n46020 , n33954 );
nor ( n46022 , n46019 , n46021 );
not ( n223784 , n46022 );
not ( n223785 , n223784 );
and ( n46025 , n46013 , n223785 );
and ( n46026 , n46012 , n223784 );
nor ( n46027 , n46025 , n46026 );
not ( n46028 , n46027 );
not ( n223790 , n31026 );
not ( n223791 , n34115 );
or ( n46031 , n223790 , n223791 );
buf ( n223793 , n42023 );
nand ( n46033 , n223793 , n31022 );
nand ( n46034 , n46031 , n46033 );
buf ( n46035 , n34917 );
and ( n46036 , n46034 , n46035 );
not ( n46037 , n46034 );
not ( n46038 , n46035 );
and ( n46039 , n46037 , n46038 );
nor ( n46040 , n46036 , n46039 );
not ( n46041 , n46040 );
xor ( n46042 , n26386 , n41041 );
xnor ( n223804 , n46042 , n41055 );
not ( n223805 , n223804 );
nand ( n46045 , n46041 , n223805 );
not ( n46046 , n38860 );
not ( n46047 , n34575 );
or ( n46048 , n46046 , n46047 );
or ( n223810 , n34575 , n38860 );
nand ( n223811 , n46048 , n223810 );
xnor ( n46051 , n223811 , n35188 );
not ( n46052 , n46051 );
and ( n46053 , n46045 , n46052 );
not ( n46054 , n46045 );
and ( n223816 , n46054 , n46051 );
nor ( n223817 , n46053 , n223816 );
not ( n46057 , n223817 );
or ( n46058 , n46028 , n46057 );
not ( n46059 , n46027 );
not ( n46060 , n223817 );
nand ( n46061 , n46059 , n46060 );
nand ( n46062 , n46058 , n46061 );
not ( n46063 , n46062 );
and ( n46064 , n223753 , n46063 );
and ( n223826 , n223752 , n46062 );
nor ( n223827 , n46064 , n223826 );
buf ( n46067 , n223827 );
and ( n46068 , n45879 , n46067 );
not ( n46069 , n45879 );
not ( n46070 , n46062 );
and ( n46071 , n223752 , n46070 );
not ( n46072 , n223752 );
and ( n46073 , n46072 , n46062 );
nor ( n46074 , n46071 , n46073 );
buf ( n223836 , n46074 );
and ( n223837 , n46069 , n223836 );
nor ( n46077 , n46068 , n223837 );
not ( n223839 , n31572 );
nand ( n223840 , n46077 , n223839 );
or ( n46080 , n45731 , n223840 );
nor ( n46081 , n46077 , n43968 );
nand ( n46082 , n46081 , n45731 );
buf ( n46083 , n35431 );
buf ( n46084 , RI173f01f0_1585);
nand ( n46085 , n46083 , n46084 );
nand ( n223847 , n46080 , n46082 , n46085 );
buf ( n223848 , n223847 );
not ( n46088 , n35045 );
nand ( n223850 , n35109 , n35157 );
not ( n223851 , n206887 );
not ( n46091 , n39400 );
or ( n46092 , n223851 , n46091 );
not ( n46093 , n206887 );
nand ( n46094 , n46093 , n45897 );
nand ( n46095 , n46092 , n46094 );
and ( n46096 , n46095 , n43589 );
not ( n223858 , n46095 );
not ( n223859 , n43589 );
and ( n46099 , n223858 , n223859 );
nor ( n46100 , n46096 , n46099 );
and ( n46101 , n223850 , n46100 );
not ( n46102 , n223850 );
not ( n46103 , n46100 );
and ( n46104 , n46102 , n46103 );
nor ( n46105 , n46101 , n46104 );
not ( n46106 , n46105 );
nand ( n223868 , n35042 , n35018 );
not ( n223869 , n29053 );
not ( n46109 , n28004 );
or ( n46110 , n223869 , n46109 );
or ( n46111 , n28004 , n29053 );
nand ( n46112 , n46110 , n46111 );
and ( n46113 , n46112 , n32916 );
not ( n46114 , n46112 );
and ( n46115 , n46114 , n32915 );
nor ( n46116 , n46113 , n46115 );
and ( n46117 , n223868 , n46116 );
not ( n46118 , n223868 );
not ( n223880 , n46116 );
and ( n223881 , n46118 , n223880 );
nor ( n46121 , n46117 , n223881 );
not ( n46122 , n46121 );
or ( n46123 , n46106 , n46122 );
or ( n46124 , n46121 , n46105 );
nand ( n223886 , n46123 , n46124 );
not ( n223887 , n41405 );
not ( n46127 , n25390 );
and ( n223889 , n223887 , n46127 );
and ( n223890 , n41405 , n25390 );
nor ( n46130 , n223889 , n223890 );
and ( n223892 , n46130 , n41415 );
not ( n223893 , n46130 );
and ( n46133 , n223893 , n41411 );
nor ( n46134 , n223892 , n46133 );
not ( n46135 , n46134 );
nand ( n46136 , n35170 , n35206 );
not ( n46137 , n46136 );
and ( n46138 , n46135 , n46137 );
nand ( n46139 , n35206 , n35170 );
and ( n46140 , n46134 , n46139 );
nor ( n46141 , n46138 , n46140 );
and ( n46142 , n223886 , n46141 );
not ( n223904 , n223886 );
not ( n223905 , n46141 );
and ( n46145 , n223904 , n223905 );
nor ( n46146 , n46142 , n46145 );
not ( n46147 , n46146 );
nand ( n46148 , n35293 , n35231 );
not ( n223910 , n46148 );
nor ( n223911 , n33096 , n221883 );
not ( n46151 , n223911 );
nand ( n46152 , n33096 , n221883 );
nand ( n46153 , n46151 , n46152 );
and ( n46154 , n46153 , n33142 );
not ( n46155 , n46153 );
and ( n46156 , n46155 , n33135 );
nor ( n46157 , n46154 , n46156 );
not ( n46158 , n46157 );
and ( n223920 , n223910 , n46158 );
not ( n223921 , n35232 );
nand ( n46161 , n223921 , n35293 );
and ( n223923 , n46161 , n46157 );
nor ( n223924 , n223920 , n223923 );
not ( n46164 , n223924 );
nand ( n46165 , n35395 , n35320 );
not ( n46166 , n217588 );
not ( n46167 , n40218 );
or ( n46168 , n46166 , n46167 );
or ( n46169 , n40218 , n217588 );
nand ( n46170 , n46168 , n46169 );
buf ( n46171 , n29411 );
and ( n46172 , n46170 , n46171 );
not ( n46173 , n46170 );
not ( n46174 , n46171 );
and ( n46175 , n46173 , n46174 );
nor ( n46176 , n46172 , n46175 );
not ( n223938 , n46176 );
and ( n223939 , n46165 , n223938 );
not ( n46179 , n46165 );
and ( n46180 , n46179 , n46176 );
nor ( n46181 , n223939 , n46180 );
not ( n46182 , n46181 );
and ( n46183 , n46164 , n46182 );
and ( n46184 , n223924 , n46181 );
nor ( n46185 , n46183 , n46184 );
not ( n46186 , n46185 );
not ( n46187 , n46186 );
and ( n46188 , n46147 , n46187 );
and ( n223950 , n46146 , n46186 );
nor ( n223951 , n46188 , n223950 );
not ( n46191 , n223951 );
not ( n46192 , n46191 );
or ( n46193 , n46088 , n46192 );
nand ( n46194 , n223951 , n35044 );
nand ( n46195 , n46193 , n46194 );
not ( n46196 , n46195 );
buf ( n46197 , n204660 );
not ( n46198 , n46197 );
not ( n46199 , n42756 );
or ( n46200 , n46198 , n46199 );
or ( n46201 , n42756 , n46197 );
nand ( n46202 , n46200 , n46201 );
nor ( n46203 , n42779 , n46202 );
not ( n46204 , n46203 );
nand ( n223966 , n220543 , n46202 );
nand ( n223967 , n46204 , n223966 );
not ( n46207 , n223967 );
not ( n223969 , n31227 );
not ( n223970 , n209722 );
not ( n46210 , n29061 );
not ( n46211 , n46210 );
or ( n46212 , n223970 , n46211 );
or ( n46213 , n46210 , n209722 );
nand ( n46214 , n46212 , n46213 );
not ( n46215 , n46214 );
not ( n223977 , RI174a9d58_908);
and ( n223978 , n29086 , n223977 );
not ( n46218 , n29086 );
and ( n46219 , n46218 , n29052 );
nor ( n46220 , n223978 , n46219 );
not ( n46221 , n46220 );
or ( n46222 , n46215 , n46221 );
or ( n46223 , n46220 , n46214 );
nand ( n223985 , n46222 , n46223 );
not ( n223986 , n223985 );
and ( n46226 , n223969 , n223986 );
and ( n46227 , n31227 , n223985 );
nor ( n46228 , n46226 , n46227 );
not ( n46229 , n28785 );
not ( n223991 , n34360 );
or ( n46231 , n46229 , n223991 );
or ( n46232 , n34360 , n28785 );
nand ( n46233 , n46231 , n46232 );
not ( n46234 , n46233 );
not ( n46235 , n34375 );
or ( n46236 , n46234 , n46235 );
or ( n46237 , n34375 , n46233 );
nand ( n46238 , n46236 , n46237 );
not ( n224000 , n46238 );
buf ( n224001 , n42512 );
not ( n46241 , n224001 );
and ( n224003 , n224000 , n46241 );
and ( n224004 , n224001 , n46238 );
nor ( n46244 , n224003 , n224004 );
not ( n46245 , n46244 );
nand ( n46246 , n46228 , n46245 );
not ( n46247 , n46246 );
and ( n46248 , n46207 , n46247 );
and ( n46249 , n223967 , n46246 );
nor ( n224011 , n46248 , n46249 );
not ( n224012 , n224011 );
buf ( n46252 , n25537 );
not ( n46253 , n46252 );
not ( n46254 , n33885 );
or ( n46255 , n46253 , n46254 );
or ( n46256 , n33885 , n46252 );
nand ( n46257 , n46255 , n46256 );
buf ( n46258 , n36662 );
and ( n46259 , n46257 , n46258 );
not ( n224021 , n46257 );
not ( n224022 , n46258 );
and ( n46262 , n224021 , n224022 );
nor ( n224024 , n46259 , n46262 );
not ( n224025 , n224024 );
not ( n46265 , n33284 );
nand ( n46266 , n33294 , n30047 );
not ( n46267 , n46266 );
nor ( n46268 , n33294 , n30047 );
nor ( n46269 , n46267 , n46268 );
not ( n46270 , n46269 );
and ( n46271 , n46265 , n46270 );
and ( n46272 , n33284 , n46269 );
nor ( n224034 , n46271 , n46272 );
not ( n224035 , n224034 );
not ( n46275 , n40726 );
and ( n46276 , n224035 , n46275 );
and ( n46277 , n224034 , n40726 );
nor ( n46278 , n46276 , n46277 );
not ( n46279 , n46278 );
not ( n46280 , n29160 );
not ( n224042 , n39400 );
or ( n224043 , n46280 , n224042 );
not ( n46283 , n29160 );
nand ( n224045 , n46283 , n45897 );
nand ( n224046 , n224043 , n224045 );
and ( n46286 , n224046 , n223859 );
not ( n46287 , n224046 );
and ( n46288 , n46287 , n204728 );
nor ( n46289 , n46286 , n46288 );
nand ( n46290 , n46279 , n46289 );
not ( n46291 , n46290 );
or ( n224053 , n224025 , n46291 );
or ( n224054 , n46290 , n224024 );
nand ( n46294 , n224053 , n224054 );
not ( n46295 , n46294 );
or ( n46296 , n224012 , n46295 );
or ( n46297 , n46294 , n224011 );
nand ( n224059 , n46296 , n46297 );
nor ( n224060 , n38255 , n33553 );
not ( n46300 , n224060 );
nand ( n224062 , n33553 , n38255 );
nand ( n224063 , n46300 , n224062 );
not ( n46303 , n35390 );
and ( n46304 , n224063 , n46303 );
not ( n46305 , n224063 );
and ( n46306 , n46305 , n35393 );
nor ( n224068 , n46304 , n46306 );
not ( n224069 , n224068 );
not ( n46309 , n28061 );
not ( n46310 , n25385 );
or ( n46311 , n46309 , n46310 );
not ( n46312 , n28061 );
nand ( n46313 , n46312 , n39811 );
nand ( n46314 , n46311 , n46313 );
and ( n224076 , n46314 , n25426 );
not ( n224077 , n46314 );
and ( n46317 , n224077 , n25429 );
nor ( n46318 , n224076 , n46317 );
not ( n46319 , n46318 );
nand ( n46320 , n224069 , n46319 );
not ( n46321 , n46320 );
not ( n46322 , n204350 );
xor ( n224084 , n41138 , n46322 );
xnor ( n224085 , n224084 , n205436 );
not ( n46325 , n224085 );
and ( n46326 , n46321 , n46325 );
and ( n46327 , n46320 , n224085 );
nor ( n46328 , n46326 , n46327 );
and ( n224090 , n224059 , n46328 );
not ( n224091 , n224059 );
not ( n46331 , n46328 );
and ( n224093 , n224091 , n46331 );
nor ( n224094 , n224090 , n224093 );
not ( n46334 , n224094 );
not ( n46335 , n214422 );
not ( n46336 , n35199 );
or ( n46337 , n46335 , n46336 );
or ( n224099 , n43913 , n214422 );
nand ( n224100 , n46337 , n224099 );
xnor ( n46340 , n224100 , n205322 );
not ( n46341 , n46340 );
not ( n46342 , n43634 );
not ( n46343 , n46342 );
not ( n46344 , n36070 );
or ( n46345 , n46343 , n46344 );
or ( n224107 , n37749 , n46342 );
nand ( n224108 , n46345 , n224107 );
buf ( n46348 , n33096 );
not ( n46349 , n46348 );
and ( n46350 , n224108 , n46349 );
not ( n46351 , n224108 );
and ( n46352 , n46351 , n46348 );
nor ( n46353 , n46350 , n46352 );
not ( n224115 , n46353 );
not ( n224116 , n30730 );
not ( n46356 , n31637 );
or ( n224118 , n224116 , n46356 );
or ( n224119 , n31637 , n30730 );
nand ( n46359 , n224118 , n224119 );
not ( n224121 , n46359 );
not ( n224122 , n37510 );
and ( n46362 , n224121 , n224122 );
and ( n46363 , n46359 , n37507 );
nor ( n46364 , n46362 , n46363 );
not ( n46365 , n46364 );
nand ( n46366 , n224115 , n46365 );
not ( n46367 , n46366 );
or ( n224129 , n46341 , n46367 );
not ( n224130 , n46340 );
not ( n46370 , n46366 );
nand ( n46371 , n224130 , n46370 );
nand ( n46372 , n224129 , n46371 );
xor ( n46373 , n36236 , n29970 );
xnor ( n46374 , n46373 , n29990 );
not ( n46375 , n46374 );
not ( n224137 , n40109 );
not ( n224138 , n37991 );
or ( n46378 , n224137 , n224138 );
not ( n224140 , n40109 );
nand ( n224141 , n224140 , n37996 );
nand ( n46381 , n46378 , n224141 );
not ( n46382 , n46381 );
not ( n46383 , n38000 );
and ( n46384 , n46382 , n46383 );
and ( n46385 , n46381 , n35481 );
nor ( n46386 , n46384 , n46385 );
not ( n224148 , n46386 );
nand ( n224149 , n46375 , n224148 );
not ( n46389 , n224149 );
buf ( n46390 , n35880 );
not ( n46391 , n46390 );
not ( n46392 , n35877 );
and ( n46393 , n46391 , n46392 );
and ( n46394 , n46390 , n35877 );
nor ( n46395 , n46393 , n46394 );
not ( n46396 , n46395 );
not ( n46397 , n35754 );
or ( n46398 , n46396 , n46397 );
or ( n224160 , n35754 , n46395 );
nand ( n224161 , n46398 , n224160 );
and ( n46401 , n224161 , n30971 );
not ( n46402 , n224161 );
and ( n46403 , n46402 , n208776 );
nor ( n46404 , n46401 , n46403 );
not ( n46405 , n46404 );
and ( n46406 , n46389 , n46405 );
and ( n46407 , n224149 , n46404 );
nor ( n46408 , n46406 , n46407 );
and ( n224170 , n46372 , n46408 );
not ( n224171 , n46372 );
not ( n46411 , n46408 );
and ( n46412 , n224171 , n46411 );
nor ( n46413 , n224170 , n46412 );
not ( n46414 , n46413 );
not ( n46415 , n46414 );
or ( n46416 , n46334 , n46415 );
not ( n46417 , n224094 );
nand ( n224179 , n46417 , n46413 );
nand ( n224180 , n46416 , n224179 );
not ( n46420 , n224180 );
not ( n224182 , n46420 );
and ( n224183 , n46196 , n224182 );
and ( n46423 , n46195 , n46420 );
nor ( n46424 , n224183 , n46423 );
not ( n46425 , n222532 );
nor ( n46426 , n46424 , n46425 );
nand ( n46427 , n36378 , n36399 );
not ( n46428 , n46427 );
xor ( n46429 , n36901 , n37746 );
xnor ( n46430 , n46429 , n32236 );
not ( n46431 , n46430 );
not ( n46432 , n46431 );
and ( n46433 , n46428 , n46432 );
nand ( n46434 , n36378 , n36399 );
and ( n224196 , n46434 , n46431 );
nor ( n224197 , n46433 , n224196 );
not ( n46437 , n224197 );
not ( n46438 , n46437 );
not ( n46439 , n37831 );
not ( n46440 , n38130 );
or ( n46441 , n46439 , n46440 );
not ( n46442 , n37831 );
nand ( n46443 , n46442 , n38129 );
nand ( n46444 , n46441 , n46443 );
and ( n224206 , n46444 , n221827 );
not ( n224207 , n46444 );
and ( n46447 , n224207 , n38137 );
nor ( n46448 , n224206 , n46447 );
nand ( n46449 , n46448 , n36551 );
not ( n46450 , n46449 );
not ( n46451 , n223562 );
and ( n46452 , n46450 , n46451 );
and ( n224214 , n46449 , n223562 );
nor ( n224215 , n46452 , n224214 );
not ( n46455 , n40529 );
not ( n224217 , n34225 );
or ( n224218 , n46455 , n224217 );
not ( n46458 , n40529 );
nand ( n46459 , n46458 , n34218 );
nand ( n46460 , n224218 , n46459 );
xor ( n46461 , n216225 , n46460 );
not ( n46462 , n46461 );
nand ( n46463 , n46462 , n36418 );
not ( n224225 , n223583 );
and ( n224226 , n46463 , n224225 );
not ( n46466 , n46463 );
and ( n46467 , n46466 , n223583 );
nor ( n46468 , n224226 , n46467 );
xor ( n46469 , n224215 , n46468 );
nand ( n46470 , n46430 , n36396 );
and ( n46471 , n46470 , n45777 );
not ( n224233 , n46470 );
and ( n224234 , n224233 , n45778 );
nor ( n46474 , n46471 , n224234 );
xnor ( n224236 , n46469 , n46474 );
not ( n224237 , n224236 );
not ( n46477 , n45740 );
not ( n46478 , n45754 );
nand ( n46479 , n36716 , n46478 );
not ( n46480 , n46479 );
or ( n46481 , n46477 , n46480 );
not ( n46482 , n45754 );
nand ( n46483 , n46482 , n36716 );
or ( n224245 , n46483 , n45740 );
nand ( n224246 , n46481 , n224245 );
xor ( n46486 , n30045 , n42400 );
xor ( n224248 , n46486 , n33300 );
not ( n224249 , n224248 );
nand ( n46489 , n224249 , n36579 );
not ( n46490 , n46489 );
not ( n46491 , n45857 );
not ( n46492 , n46491 );
not ( n224254 , n46492 );
and ( n224255 , n46490 , n224254 );
and ( n46495 , n46489 , n46492 );
nor ( n46496 , n224255 , n46495 );
and ( n46497 , n224246 , n46496 );
not ( n46498 , n224246 );
not ( n46499 , n46496 );
and ( n46500 , n46498 , n46499 );
nor ( n46501 , n46497 , n46500 );
not ( n46502 , n46501 );
and ( n224264 , n224237 , n46502 );
not ( n224265 , n224237 );
and ( n46505 , n224265 , n46501 );
nor ( n46506 , n224264 , n46505 );
not ( n46507 , n46506 );
or ( n46508 , n46438 , n46507 );
not ( n46509 , n46437 );
not ( n46510 , n46501 );
not ( n224272 , n224236 );
or ( n224273 , n46510 , n224272 );
nand ( n46513 , n224237 , n46502 );
nand ( n46514 , n224273 , n46513 );
nand ( n46515 , n46509 , n46514 );
nand ( n46516 , n46508 , n46515 );
buf ( n46517 , n26250 );
not ( n46518 , n46517 );
not ( n224280 , RI173d9270_1697);
xor ( n224281 , n224280 , n42772 );
xor ( n46521 , n224281 , n42778 );
not ( n46522 , n46521 );
or ( n46523 , n46518 , n46522 );
or ( n46524 , n46521 , n46517 );
nand ( n46525 , n46523 , n46524 );
and ( n46526 , n46525 , n43122 );
not ( n46527 , n46525 );
and ( n46528 , n46527 , n38973 );
nor ( n46529 , n46526 , n46528 );
not ( n46530 , n46529 );
not ( n224292 , n37862 );
not ( n224293 , n38130 );
or ( n46533 , n224292 , n224293 );
not ( n46534 , n37862 );
nand ( n46535 , n46534 , n38129 );
nand ( n46536 , n46533 , n46535 );
and ( n224298 , n46536 , n221827 );
not ( n224299 , n46536 );
not ( n46539 , n38140 );
and ( n46540 , n224299 , n46539 );
nor ( n46541 , n224298 , n46540 );
not ( n46542 , n46541 );
nand ( n46543 , n46530 , n46542 );
not ( n46544 , n46543 );
not ( n224306 , n45902 );
and ( n224307 , n46544 , n224306 );
not ( n46547 , n46541 );
nand ( n46548 , n46547 , n46530 );
and ( n46549 , n46548 , n45902 );
nor ( n46550 , n224307 , n46549 );
not ( n46551 , n46550 );
not ( n46552 , n46551 );
not ( n224314 , n41448 );
buf ( n224315 , RI173ea610_1613);
not ( n46555 , n224315 );
not ( n46556 , RI173a1920_1968);
not ( n46557 , n46556 );
or ( n46558 , n46555 , n46557 );
not ( n46559 , RI173ea610_1613);
buf ( n46560 , RI173a1920_1968);
nand ( n224322 , n46559 , n46560 );
nand ( n224323 , n46558 , n224322 );
not ( n46563 , RI1746c4f8_1208);
and ( n46564 , n224323 , n46563 );
not ( n46565 , n224323 );
buf ( n46566 , RI1746c4f8_1208);
and ( n46567 , n46565 , n46566 );
nor ( n46568 , n46564 , n46567 );
buf ( n224330 , RI19a82790_2777);
nand ( n224331 , n29151 , n224330 );
buf ( n46571 , RI1750d2f8_725);
and ( n46572 , n224331 , n46571 );
not ( n46573 , n224331 );
not ( n46574 , RI1750d2f8_725);
and ( n46575 , n46573 , n46574 );
nor ( n46576 , n46572 , n46575 );
xor ( n46577 , n46568 , n46576 );
buf ( n46578 , RI19aa1618_2557);
nand ( n46579 , n26325 , n46578 );
not ( n46580 , RI174868f8_1080);
and ( n224342 , n46579 , n46580 );
not ( n224343 , n46579 );
buf ( n46583 , RI174868f8_1080);
and ( n46584 , n224343 , n46583 );
nor ( n46585 , n224342 , n46584 );
xnor ( n46586 , n46577 , n46585 );
not ( n46587 , n46586 );
not ( n46588 , n46587 );
not ( n224350 , n30531 );
and ( n224351 , n46588 , n224350 );
and ( n46591 , n46587 , n30531 );
nor ( n46592 , n224351 , n46591 );
not ( n46593 , n46592 );
and ( n46594 , n224314 , n46593 );
buf ( n46595 , n41447 );
not ( n46596 , n46595 );
and ( n46597 , n46596 , n46592 );
nor ( n46598 , n46594 , n46597 );
and ( n224360 , n35542 , n40562 );
not ( n224361 , n35542 );
and ( n46601 , n224361 , n40568 );
nor ( n224363 , n224360 , n46601 );
not ( n224364 , n224363 );
not ( n46604 , n29525 );
and ( n46605 , n224364 , n46604 );
and ( n46606 , n224363 , n29525 );
nor ( n46607 , n46605 , n46606 );
not ( n224369 , n46607 );
nand ( n224370 , n46598 , n224369 );
not ( n46610 , n224370 );
not ( n224372 , n45963 );
or ( n224373 , n46610 , n224372 );
or ( n46613 , n45963 , n224370 );
nand ( n46614 , n224373 , n46613 );
not ( n46615 , n46614 );
not ( n46616 , n46615 );
or ( n46617 , n46552 , n46616 );
nand ( n46618 , n46614 , n46550 );
nand ( n224380 , n46617 , n46618 );
not ( n224381 , n29080 );
not ( n46621 , n36568 );
or ( n224383 , n224381 , n46621 );
not ( n46623 , n29080 );
nand ( n46624 , n46623 , n205766 );
nand ( n46625 , n224383 , n46624 );
not ( n46626 , n46625 );
not ( n46627 , n32916 );
and ( n46628 , n46626 , n46627 );
and ( n46629 , n46625 , n32916 );
nor ( n46630 , n46628 , n46629 );
not ( n46631 , n46630 );
not ( n46632 , n35096 );
not ( n46633 , n39873 );
not ( n46634 , n46633 );
or ( n224396 , n46632 , n46634 );
not ( n224397 , n35096 );
nand ( n46637 , n224397 , n39874 );
nand ( n46638 , n224396 , n46637 );
not ( n46639 , n204672 );
and ( n46640 , n46638 , n46639 );
not ( n224402 , n46638 );
and ( n224403 , n224402 , n204672 );
nor ( n46643 , n46640 , n224403 );
not ( n46644 , n46643 );
nand ( n46645 , n46631 , n46644 );
and ( n46646 , n46645 , n45946 );
not ( n46647 , n46645 );
and ( n46648 , n46647 , n45947 );
nor ( n46649 , n46646 , n46648 );
not ( n46650 , n46649 );
and ( n224412 , n224380 , n46650 );
not ( n224413 , n224380 );
and ( n46653 , n224413 , n46649 );
nor ( n224415 , n224412 , n46653 );
not ( n224416 , n224415 );
not ( n46656 , n221323 );
xor ( n46657 , n205279 , n46656 );
xnor ( n46658 , n46657 , n31778 );
not ( n46659 , n46658 );
buf ( n46660 , n35382 );
not ( n46661 , n46660 );
not ( n46662 , n29647 );
or ( n46663 , n46661 , n46662 );
not ( n46664 , n29645 );
not ( n46665 , n46664 );
or ( n224427 , n46665 , n46660 );
nand ( n224428 , n46663 , n224427 );
buf ( n46668 , n39968 );
and ( n46669 , n224428 , n46668 );
not ( n46670 , n224428 );
buf ( n46671 , n39974 );
and ( n46672 , n46670 , n46671 );
nor ( n46673 , n46669 , n46672 );
nand ( n224435 , n46659 , n46673 );
not ( n224436 , n224435 );
not ( n46676 , n46001 );
and ( n46677 , n224436 , n46676 );
and ( n46678 , n224435 , n46001 );
nor ( n46679 , n46677 , n46678 );
not ( n46680 , n38970 );
not ( n46681 , n204935 );
not ( n224443 , n46681 );
not ( n224444 , n224443 );
or ( n46684 , n46680 , n224444 );
not ( n46685 , n224443 );
not ( n46686 , n38970 );
nand ( n46687 , n46685 , n46686 );
nand ( n224449 , n46684 , n46687 );
not ( n224450 , n204981 );
and ( n46690 , n224449 , n224450 );
not ( n224452 , n224449 );
and ( n224453 , n224452 , n204977 );
nor ( n46693 , n46690 , n224453 );
not ( n46694 , n46693 );
xor ( n46695 , n42283 , n45744 );
xnor ( n46696 , n46695 , n204825 );
not ( n46697 , n46696 );
nand ( n46698 , n46694 , n46697 );
and ( n46699 , n46698 , n223804 );
not ( n46700 , n46698 );
and ( n224462 , n46700 , n223805 );
nor ( n224463 , n46699 , n224462 );
xor ( n46703 , n46679 , n224463 );
not ( n46704 , n46703 );
not ( n46705 , n46704 );
and ( n46706 , n224416 , n46705 );
and ( n46707 , n46704 , n224415 );
nor ( n46708 , n46706 , n46707 );
and ( n46709 , n46516 , n46708 );
not ( n46710 , n46516 );
not ( n224472 , n46703 );
not ( n224473 , n224415 );
not ( n46713 , n224473 );
or ( n46714 , n224472 , n46713 );
nand ( n46715 , n224415 , n46704 );
nand ( n46716 , n46714 , n46715 );
buf ( n224478 , n46716 );
and ( n224479 , n46710 , n224478 );
nor ( n46719 , n46709 , n224479 );
not ( n46720 , n210564 );
not ( n46721 , n37533 );
or ( n46722 , n46720 , n46721 );
or ( n46723 , n37533 , n210564 );
nand ( n46724 , n46722 , n46723 );
and ( n46725 , n46724 , n30100 );
not ( n46726 , n46724 );
and ( n46727 , n46726 , n38037 );
nor ( n46728 , n46725 , n46727 );
not ( n224490 , n46728 );
not ( n224491 , n205295 );
buf ( n46731 , n34873 );
not ( n46732 , n46731 );
or ( n46733 , n224491 , n46732 );
not ( n46734 , n46731 );
nand ( n46735 , n46734 , n205291 );
nand ( n46736 , n46733 , n46735 );
buf ( n46737 , n219430 );
and ( n46738 , n46736 , n46737 );
not ( n46739 , n46736 );
not ( n46740 , n46737 );
and ( n224502 , n46739 , n46740 );
nor ( n224503 , n46738 , n224502 );
nand ( n46743 , n224490 , n224503 );
not ( n46744 , n46743 );
not ( n46745 , n30330 );
not ( n46746 , n29335 );
not ( n46747 , n46746 );
or ( n46748 , n46745 , n46747 );
or ( n224510 , n29336 , n30330 );
nand ( n224511 , n46748 , n224510 );
and ( n46751 , n224511 , n41149 );
not ( n46752 , n224511 );
not ( n46753 , n41149 );
and ( n46754 , n46752 , n46753 );
nor ( n46755 , n46751 , n46754 );
not ( n46756 , n46755 );
and ( n46757 , n46744 , n46756 );
and ( n46758 , n46743 , n46755 );
nor ( n224520 , n46757 , n46758 );
not ( n224521 , n224520 );
not ( n46761 , n224521 );
not ( n46762 , n44909 );
not ( n46763 , n32652 );
or ( n46764 , n46762 , n46763 );
or ( n46765 , n32652 , n44909 );
nand ( n46766 , n46764 , n46765 );
nor ( n46767 , n40963 , n46766 );
not ( n224529 , n46767 );
nand ( n224530 , n40963 , n46766 );
nand ( n46770 , n224529 , n224530 );
not ( n46771 , n26295 );
not ( n46772 , n38971 );
or ( n46773 , n46771 , n46772 );
not ( n224535 , n26295 );
nand ( n224536 , n224535 , n219976 );
nand ( n46776 , n46773 , n224536 );
and ( n46777 , n46776 , n39007 );
not ( n46778 , n46776 );
and ( n46779 , n46778 , n39002 );
nor ( n46780 , n46777 , n46779 );
nand ( n46781 , n46770 , n46780 );
not ( n46782 , n36023 );
not ( n46783 , n39244 );
or ( n46784 , n46782 , n46783 );
not ( n46785 , n36023 );
nand ( n224547 , n46785 , n39250 );
nand ( n224548 , n46784 , n224547 );
and ( n46788 , n224548 , n42956 );
not ( n46789 , n224548 );
and ( n46790 , n46789 , n45942 );
nor ( n46791 , n46788 , n46790 );
and ( n46792 , n46781 , n46791 );
not ( n46793 , n46781 );
not ( n224555 , n46791 );
and ( n224556 , n46793 , n224555 );
nor ( n46796 , n46792 , n224556 );
not ( n46797 , n46796 );
not ( n224559 , n28528 );
not ( n224560 , n37406 );
or ( n46800 , n224559 , n224560 );
or ( n46801 , n37406 , n28528 );
nand ( n46802 , n46800 , n46801 );
and ( n46803 , n46802 , n29608 );
not ( n46804 , n46802 );
and ( n46805 , n46804 , n44492 );
nor ( n46806 , n46803 , n46805 );
not ( n46807 , n43228 );
not ( n224569 , n41856 );
or ( n224570 , n46807 , n224569 );
not ( n46810 , n41855 );
or ( n46811 , n46810 , n43228 );
nand ( n46812 , n224570 , n46811 );
and ( n46813 , n46812 , n217819 );
not ( n46814 , n46812 );
not ( n46815 , n40057 );
not ( n46816 , n46815 );
and ( n46817 , n46814 , n46816 );
nor ( n46818 , n46813 , n46817 );
not ( n46819 , n46818 );
nand ( n224581 , n46806 , n46819 );
not ( n224582 , n224581 );
not ( n46822 , n41063 );
not ( n46823 , n44132 );
not ( n46824 , n33095 );
or ( n46825 , n46823 , n46824 );
or ( n46826 , n33095 , n44132 );
nand ( n46827 , n46825 , n46826 );
not ( n46828 , n46827 );
or ( n46829 , n46822 , n46828 );
or ( n46830 , n46827 , n33135 );
nand ( n46831 , n46829 , n46830 );
buf ( n46832 , n46831 );
not ( n46833 , n46832 );
and ( n224595 , n224582 , n46833 );
and ( n224596 , n224581 , n46832 );
nor ( n46836 , n224595 , n224596 );
not ( n46837 , n46836 );
or ( n46838 , n46797 , n46837 );
or ( n46839 , n46836 , n46796 );
nand ( n46840 , n46838 , n46839 );
not ( n46841 , n30034 );
not ( n46842 , n37496 );
not ( n46843 , n40072 );
or ( n224605 , n46842 , n46843 );
or ( n224606 , n26145 , n37496 );
nand ( n46846 , n224605 , n224606 );
not ( n224608 , n46846 );
or ( n224609 , n46841 , n224608 );
or ( n46849 , n46846 , n30034 );
nand ( n46850 , n224609 , n46849 );
not ( n46851 , n46850 );
xor ( n46852 , n208577 , n36457 );
xnor ( n46853 , n46852 , n40935 );
not ( n46854 , n46853 );
nand ( n46855 , n46851 , n46854 );
not ( n46856 , n44690 );
not ( n46857 , n32606 );
nor ( n46858 , n28508 , n46857 );
not ( n224620 , n46858 );
nand ( n224621 , n28508 , n46857 );
nand ( n46861 , n224620 , n224621 );
not ( n224623 , n46861 );
and ( n224624 , n46856 , n224623 );
and ( n46864 , n44690 , n46861 );
nor ( n224626 , n224624 , n46864 );
and ( n224627 , n46855 , n224626 );
not ( n46867 , n46855 );
not ( n46868 , n224626 );
and ( n46869 , n46867 , n46868 );
nor ( n46870 , n224627 , n46869 );
xnor ( n46871 , n46840 , n46870 );
not ( n46872 , n46755 );
not ( n224634 , n224503 );
nand ( n224635 , n46872 , n224634 );
not ( n46875 , n224635 );
not ( n46876 , n46875 );
buf ( n46877 , n31868 );
xor ( n46878 , n46877 , n205385 );
buf ( n46879 , RI173cb680_1764);
xor ( n46880 , n46879 , n205341 );
xnor ( n224642 , n46880 , n205349 );
buf ( n224643 , n224642 );
xnor ( n46883 , n46878 , n224643 );
not ( n46884 , n46883 );
not ( n46885 , n46884 );
or ( n46886 , n46876 , n46885 );
nand ( n46887 , n46883 , n224635 );
nand ( n46888 , n46886 , n46887 );
not ( n46889 , n204860 );
not ( n46890 , n34708 );
and ( n46891 , n46889 , n46890 );
and ( n46892 , n204860 , n34708 );
nor ( n46893 , n46891 , n46892 );
not ( n46894 , n204895 );
and ( n224656 , n46893 , n46894 );
not ( n224657 , n46893 );
and ( n46897 , n224657 , n204895 );
nor ( n224659 , n224656 , n46897 );
not ( n224660 , n224659 );
buf ( n46900 , RI17407e90_1469);
not ( n46901 , n46900 );
not ( n46902 , n27842 );
or ( n46903 , n46901 , n46902 );
nand ( n46904 , n32454 , n30584 );
nand ( n46905 , n46903 , n46904 );
and ( n224667 , n46905 , n43155 );
not ( n224668 , n46905 );
and ( n46908 , n224668 , n27802 );
nor ( n46909 , n224667 , n46908 );
nand ( n46910 , n224660 , n46909 );
not ( n46911 , n46910 );
buf ( n224673 , n46576 );
not ( n224674 , n224673 );
not ( n46914 , n224674 );
not ( n46915 , n35703 );
not ( n46916 , n46915 );
not ( n46917 , n46916 );
or ( n46918 , n46914 , n46917 );
nand ( n46919 , n38829 , n224673 );
nand ( n46920 , n46918 , n46919 );
not ( n46921 , n25766 );
and ( n46922 , n46920 , n46921 );
not ( n46923 , n46920 );
not ( n224685 , n25762 );
not ( n224686 , n224685 );
and ( n46926 , n46923 , n224686 );
nor ( n46927 , n46922 , n46926 );
not ( n46928 , n46927 );
and ( n46929 , n46911 , n46928 );
and ( n224691 , n46910 , n46927 );
nor ( n224692 , n46929 , n224691 );
and ( n46932 , n46888 , n224692 );
not ( n46933 , n46888 );
not ( n46934 , n224692 );
and ( n46935 , n46933 , n46934 );
nor ( n46936 , n46932 , n46935 );
not ( n46937 , n46936 );
and ( n224699 , n46871 , n46937 );
not ( n224700 , n46871 );
and ( n46940 , n224700 , n46936 );
nor ( n46941 , n224699 , n46940 );
not ( n46942 , n46941 );
or ( n46943 , n46761 , n46942 );
not ( n46944 , n224521 );
not ( n46945 , n46936 );
not ( n224707 , n46871 );
not ( n224708 , n224707 );
or ( n46948 , n46945 , n224708 );
nand ( n46949 , n46871 , n46937 );
nand ( n46950 , n46948 , n46949 );
nand ( n46951 , n46944 , n46950 );
nand ( n46952 , n46943 , n46951 );
not ( n46953 , n37899 );
not ( n224715 , n37261 );
or ( n224716 , n46953 , n224715 );
not ( n46956 , n37899 );
nand ( n46957 , n46956 , n37260 );
nand ( n46958 , n224716 , n46957 );
and ( n46959 , n46958 , n39361 );
not ( n46960 , n46958 );
and ( n46961 , n46960 , n222184 );
nor ( n224723 , n46959 , n46961 );
buf ( n224724 , RI1745c508_1286);
xor ( n46964 , n28757 , n206535 );
xor ( n46965 , n46964 , n28765 );
not ( n46966 , n46965 );
and ( n46967 , n224724 , n46966 );
not ( n46968 , n224724 );
and ( n46969 , n46968 , n46965 );
nor ( n46970 , n46967 , n46969 );
not ( n46971 , n46970 );
not ( n46972 , n28816 );
and ( n46973 , n46971 , n46972 );
and ( n224735 , n46970 , n28816 );
nor ( n224736 , n46973 , n224735 );
nand ( n46976 , n224723 , n224736 );
not ( n46977 , n46976 );
not ( n46978 , n45284 );
not ( n46979 , n30685 );
or ( n46980 , n46978 , n46979 );
or ( n46981 , n30685 , n45284 );
nand ( n46982 , n46980 , n46981 );
xor ( n46983 , n34139 , n46982 );
not ( n46984 , n46983 );
and ( n46985 , n46977 , n46984 );
and ( n224747 , n46976 , n46983 );
nor ( n224748 , n46985 , n224747 );
not ( n46988 , n224748 );
not ( n46989 , n37068 );
not ( n46990 , n43695 );
or ( n46991 , n46989 , n46990 );
xor ( n46992 , n31475 , n40788 );
xnor ( n46993 , n46992 , n40811 );
not ( n46994 , n46993 );
or ( n46995 , n46994 , n37068 );
nand ( n224757 , n46991 , n46995 );
and ( n224758 , n224757 , n221462 );
not ( n224759 , n224757 );
and ( n224760 , n224759 , n29371 );
nor ( n47000 , n224758 , n224760 );
not ( n224762 , n34203 );
not ( n224763 , n40944 );
or ( n47003 , n224762 , n224763 );
or ( n47004 , n40944 , n34203 );
nand ( n47005 , n47003 , n47004 );
and ( n47006 , n47005 , n32175 );
not ( n224768 , n47005 );
and ( n224769 , n224768 , n32176 );
nor ( n47009 , n47006 , n224769 );
nand ( n47010 , n47000 , n47009 );
not ( n47011 , n30902 );
xor ( n47012 , n40880 , n40884 );
xnor ( n47013 , n47012 , n40893 );
not ( n47014 , n47013 );
or ( n224776 , n47011 , n47014 );
or ( n224777 , n47013 , n30902 );
nand ( n47017 , n224776 , n224777 );
and ( n47018 , n47017 , n32053 );
not ( n47019 , n47017 );
and ( n47020 , n47019 , n32050 );
nor ( n47021 , n47018 , n47020 );
and ( n47022 , n47010 , n47021 );
not ( n47023 , n47010 );
not ( n47024 , n47021 );
and ( n47025 , n47023 , n47024 );
nor ( n47026 , n47022 , n47025 );
not ( n224788 , n47026 );
or ( n224789 , n46988 , n224788 );
or ( n47029 , n47026 , n224748 );
nand ( n47030 , n224789 , n47029 );
not ( n47031 , n32284 );
buf ( n47032 , n33602 );
and ( n47033 , n47032 , n40413 );
not ( n47034 , n47032 );
and ( n47035 , n47034 , n43459 );
nor ( n47036 , n47033 , n47035 );
not ( n47037 , n47036 );
or ( n47038 , n47031 , n47037 );
or ( n224800 , n47036 , n42300 );
nand ( n224801 , n47038 , n224800 );
buf ( n47041 , n224801 );
not ( n224803 , n47041 );
not ( n224804 , n33500 );
not ( n47044 , n28555 );
or ( n224806 , n224804 , n47044 );
not ( n224807 , n33500 );
nand ( n47047 , n224807 , n38250 );
nand ( n47048 , n224806 , n47047 );
and ( n47049 , n47048 , n38257 );
not ( n47050 , n47048 );
and ( n47051 , n47050 , n35358 );
nor ( n47052 , n47049 , n47051 );
nor ( n224814 , n224803 , n47052 );
not ( n224815 , n224814 );
xor ( n47055 , n26227 , n38973 );
xor ( n47056 , n47055 , n45672 );
not ( n47057 , n47056 );
not ( n47058 , n47057 );
or ( n224820 , n224815 , n47058 );
not ( n224821 , n224814 );
nand ( n47061 , n224821 , n47056 );
nand ( n47062 , n224820 , n47061 );
and ( n47063 , n47030 , n47062 );
not ( n47064 , n47030 );
not ( n47065 , n47062 );
and ( n47066 , n47064 , n47065 );
nor ( n47067 , n47063 , n47066 );
and ( n47068 , n40710 , n26050 );
not ( n47069 , n40710 );
and ( n47070 , n47069 , n26047 );
nor ( n224832 , n47068 , n47070 );
and ( n224833 , n224832 , n26009 );
not ( n47073 , n224832 );
and ( n47074 , n47073 , n38587 );
nor ( n47075 , n224833 , n47074 );
buf ( n47076 , n32360 );
not ( n47077 , n47076 );
not ( n47078 , n210118 );
and ( n224840 , n47077 , n47078 );
and ( n224841 , n47076 , n210118 );
nor ( n47081 , n224840 , n224841 );
not ( n224843 , n47081 );
not ( n224844 , n38204 );
or ( n47084 , n224843 , n224844 );
or ( n47085 , n29411 , n47081 );
nand ( n47086 , n47084 , n47085 );
and ( n47087 , n47086 , n29457 );
not ( n47088 , n47086 );
and ( n224850 , n47088 , n29460 );
nor ( n224851 , n47087 , n224850 );
not ( n47091 , n224851 );
nand ( n224853 , n47075 , n47091 );
not ( n224854 , n42325 );
not ( n47094 , n28159 );
and ( n224856 , n224854 , n47094 );
and ( n224857 , n42325 , n28159 );
nor ( n224858 , n224856 , n224857 );
buf ( n224859 , n40976 );
and ( n47099 , n224858 , n224859 );
not ( n47100 , n224858 );
not ( n47101 , n224859 );
and ( n47102 , n47100 , n47101 );
nor ( n47103 , n47099 , n47102 );
not ( n224865 , n47103 );
and ( n224866 , n224853 , n224865 );
not ( n47106 , n224853 );
and ( n47107 , n47106 , n47103 );
nor ( n47108 , n224866 , n47107 );
not ( n47109 , n47108 );
not ( n47110 , n47109 );
xor ( n47111 , n36825 , n42623 );
not ( n47112 , n42593 );
not ( n224874 , n47112 );
xnor ( n224875 , n47111 , n224874 );
not ( n47115 , n32442 );
buf ( n224877 , n217118 );
not ( n224878 , n224877 );
not ( n47118 , n32405 );
or ( n47119 , n224878 , n47118 );
or ( n47120 , n32405 , n224877 );
nand ( n47121 , n47119 , n47120 );
not ( n224883 , n47121 );
not ( n224884 , n224883 );
or ( n47124 , n47115 , n224884 );
nand ( n47125 , n47121 , n32443 );
nand ( n47126 , n47124 , n47125 );
nand ( n47127 , n224875 , n47126 );
not ( n47128 , n47127 );
not ( n47129 , n31244 );
not ( n47130 , n33195 );
or ( n47131 , n47129 , n47130 );
or ( n224893 , n33195 , n31244 );
nand ( n224894 , n47131 , n224893 );
buf ( n47134 , n46746 );
not ( n47135 , n47134 );
and ( n47136 , n224894 , n47135 );
not ( n47137 , n224894 );
and ( n47138 , n47137 , n29336 );
nor ( n47139 , n47136 , n47138 );
not ( n47140 , n47139 );
and ( n47141 , n47128 , n47140 );
not ( n224903 , n47126 );
not ( n224904 , n224903 );
nand ( n47144 , n224904 , n224875 );
and ( n47145 , n47144 , n47139 );
nor ( n47146 , n47141 , n47145 );
not ( n47147 , n47146 );
not ( n47148 , n47147 );
or ( n47149 , n47110 , n47148 );
nand ( n224911 , n47146 , n47108 );
nand ( n224912 , n47149 , n224911 );
and ( n47152 , n47067 , n224912 );
not ( n224914 , n47067 );
not ( n224915 , n224912 );
and ( n47155 , n224914 , n224915 );
nor ( n47156 , n47152 , n47155 );
buf ( n47157 , n47156 );
and ( n47158 , n46952 , n47157 );
not ( n47159 , n46952 );
and ( n47160 , n47067 , n224915 );
not ( n47161 , n47067 );
and ( n47162 , n47161 , n224912 );
nor ( n224924 , n47160 , n47162 );
buf ( n224925 , n224924 );
and ( n47165 , n47159 , n224925 );
nor ( n47166 , n47158 , n47165 );
not ( n47167 , n47166 );
nand ( n47168 , n46426 , n46719 , n47167 );
not ( n47169 , n46424 );
not ( n47170 , n47169 );
not ( n47171 , n46719 );
or ( n47172 , n47170 , n47171 );
buf ( n47173 , n31571 );
nor ( n47174 , n47167 , n47173 );
nand ( n47175 , n47172 , n47174 );
buf ( n224937 , n35431 );
nand ( n224938 , n224937 , n204758 );
nand ( n47178 , n47168 , n47175 , n224938 );
buf ( n47179 , n47178 );
not ( n47180 , n37020 );
not ( n47181 , n205298 );
not ( n47182 , n34873 );
or ( n47183 , n47181 , n47182 );
nand ( n47184 , n36990 , n205301 );
nand ( n224946 , n47183 , n47184 );
not ( n224947 , n224946 );
or ( n47187 , n47180 , n224947 );
or ( n224949 , n224946 , n37020 );
nand ( n224950 , n47187 , n224949 );
not ( n47190 , n224950 );
nand ( n47191 , n47190 , n40637 );
not ( n47192 , n47191 );
not ( n47193 , n40383 );
not ( n47194 , n29518 );
or ( n47195 , n47193 , n47194 );
or ( n47196 , n29518 , n40383 );
nand ( n47197 , n47195 , n47196 );
and ( n224959 , n47197 , n29563 );
not ( n224960 , n47197 );
and ( n47200 , n224960 , n29562 );
nor ( n47201 , n224959 , n47200 );
not ( n47202 , n47201 );
not ( n47203 , n47202 );
and ( n47204 , n47192 , n47203 );
and ( n47205 , n47191 , n47202 );
nor ( n224967 , n47204 , n47205 );
not ( n224968 , n224967 );
not ( n47208 , n224968 );
nand ( n224970 , n224950 , n47201 );
not ( n224971 , n224970 );
not ( n47211 , n40626 );
and ( n47212 , n224971 , n47211 );
and ( n47213 , n224970 , n40626 );
nor ( n47214 , n47212 , n47213 );
xor ( n47215 , n204456 , n27926 );
buf ( n47216 , n25926 );
xnor ( n47217 , n47215 , n47216 );
not ( n47218 , n47217 );
not ( n224980 , n40491 );
nand ( n224981 , n47218 , n224980 );
and ( n224982 , n224981 , n40572 );
not ( n224983 , n224981 );
and ( n47223 , n224983 , n40571 );
nor ( n47224 , n224982 , n47223 );
xor ( n47225 , n47214 , n47224 );
not ( n47226 , n210628 );
not ( n47227 , n36702 );
or ( n47228 , n47226 , n47227 );
or ( n224990 , n36705 , n210628 );
nand ( n224991 , n47228 , n224990 );
not ( n47231 , n36710 );
and ( n224993 , n224991 , n47231 );
not ( n224994 , n224991 );
and ( n47234 , n224994 , n214472 );
nor ( n47235 , n224993 , n47234 );
not ( n47236 , n47235 );
not ( n47237 , n42610 );
not ( n224999 , n34564 );
or ( n225000 , n47237 , n224999 );
nand ( n47240 , n43326 , n42607 );
nand ( n225002 , n225000 , n47240 );
and ( n225003 , n225002 , n42473 );
not ( n47243 , n225002 );
and ( n47244 , n47243 , n42472 );
nor ( n47245 , n225003 , n47244 );
nand ( n47246 , n47236 , n47245 );
buf ( n47247 , n40736 );
not ( n47248 , n47247 );
and ( n47249 , n47246 , n47248 );
not ( n47250 , n47246 );
and ( n225012 , n47250 , n47247 );
nor ( n225013 , n47249 , n225012 );
xnor ( n47253 , n47225 , n225013 );
not ( n47254 , n47253 );
not ( n47255 , n47254 );
not ( n47256 , n27979 );
not ( n47257 , n204505 );
or ( n47258 , n47256 , n47257 );
nand ( n225020 , n204508 , n27975 );
nand ( n225021 , n47258 , n225020 );
not ( n47261 , n219115 );
not ( n47262 , n47261 );
xor ( n47263 , n225021 , n47262 );
not ( n47264 , n47263 );
not ( n225026 , n35133 );
not ( n225027 , n38775 );
or ( n47267 , n225026 , n225027 );
nand ( n47268 , n38774 , n35136 );
nand ( n47269 , n47267 , n47268 );
not ( n47270 , n47269 );
not ( n225032 , n206777 );
and ( n225033 , n47270 , n225032 );
and ( n47273 , n206777 , n47269 );
nor ( n47274 , n225033 , n47273 );
not ( n47275 , n47274 );
nand ( n47276 , n47264 , n47275 );
not ( n225038 , n47276 );
not ( n225039 , n40818 );
and ( n47279 , n225038 , n225039 );
and ( n47280 , n47276 , n40818 );
nor ( n47281 , n47279 , n47280 );
buf ( n47282 , RI1740c030_1449);
not ( n225044 , n47282 );
not ( n225045 , n211807 );
or ( n47285 , n225044 , n225045 );
nand ( n47286 , n37472 , n204868 );
nand ( n47287 , n47285 , n47286 );
and ( n47288 , n47287 , n34090 );
not ( n47289 , n47287 );
and ( n47290 , n47289 , n34104 );
nor ( n225052 , n47288 , n47290 );
not ( n225053 , n225052 );
xor ( n47293 , n31846 , n205389 );
xnor ( n47294 , n47293 , n224643 );
nand ( n47295 , n225053 , n47294 );
not ( n47296 , n47295 );
not ( n47297 , n40669 );
and ( n47298 , n47296 , n47297 );
and ( n225060 , n47295 , n40669 );
nor ( n225061 , n47298 , n225060 );
not ( n47301 , n225061 );
and ( n47302 , n47281 , n47301 );
not ( n47303 , n47281 );
and ( n47304 , n47303 , n225061 );
nor ( n47305 , n47302 , n47304 );
not ( n47306 , n47305 );
not ( n47307 , n47306 );
and ( n47308 , n47255 , n47307 );
and ( n47309 , n47254 , n47306 );
nor ( n47310 , n47308 , n47309 );
not ( n47311 , n47310 );
or ( n47312 , n47208 , n47311 );
not ( n47313 , n224968 );
not ( n225075 , n47305 );
not ( n225076 , n47253 );
or ( n47316 , n225075 , n225076 );
not ( n47317 , n47253 );
nand ( n47318 , n47317 , n47306 );
nand ( n47319 , n47316 , n47318 );
nand ( n47320 , n47313 , n47319 );
nand ( n47321 , n47312 , n47320 );
buf ( n225083 , n220460 );
and ( n225084 , n47321 , n225083 );
not ( n47324 , n47321 );
buf ( n225086 , n220467 );
and ( n225087 , n47324 , n225086 );
nor ( n47327 , n225084 , n225087 );
xor ( n225089 , n34534 , n45280 );
buf ( n225090 , n44135 );
not ( n47330 , n225090 );
xnor ( n47331 , n225089 , n47330 );
not ( n47332 , n47331 );
not ( n47333 , n47332 );
buf ( n47334 , n33753 );
xor ( n47335 , n47334 , n33195 );
not ( n47336 , n34825 );
xnor ( n47337 , n47335 , n47336 );
not ( n47338 , n47337 );
not ( n47339 , n33523 );
not ( n225101 , n28555 );
or ( n225102 , n47339 , n225101 );
not ( n47342 , n33523 );
buf ( n225104 , n38250 );
nand ( n225105 , n47342 , n225104 );
nand ( n47345 , n225102 , n225105 );
buf ( n47346 , n35358 );
and ( n47347 , n47345 , n47346 );
not ( n225109 , n47345 );
and ( n225110 , n225109 , n38257 );
nor ( n225111 , n47347 , n225110 );
nand ( n225112 , n47338 , n225111 );
not ( n47352 , n225112 );
or ( n47353 , n47333 , n47352 );
not ( n47354 , n225111 );
not ( n47355 , n47354 );
nand ( n47356 , n47355 , n47338 );
or ( n47357 , n47356 , n47332 );
nand ( n225119 , n47353 , n47357 );
not ( n225120 , n225119 );
and ( n47360 , n31513 , n37171 );
not ( n47361 , n31513 );
and ( n47362 , n47361 , n38690 );
nor ( n47363 , n47360 , n47362 );
and ( n47364 , n47363 , n37196 );
not ( n47365 , n47363 );
and ( n225127 , n47365 , n37193 );
nor ( n225128 , n47364 , n225127 );
not ( n47368 , n33592 );
not ( n47369 , n43460 );
or ( n47370 , n47368 , n47369 );
not ( n47371 , n33592 );
nand ( n47372 , n47371 , n44238 );
nand ( n47373 , n47370 , n47372 );
and ( n47374 , n47373 , n32280 );
not ( n47375 , n47373 );
and ( n225137 , n47375 , n210046 );
nor ( n225138 , n47374 , n225137 );
nand ( n47378 , n225128 , n225138 );
not ( n47379 , n47378 );
not ( n47380 , n31180 );
not ( n47381 , n31424 );
not ( n225143 , n47381 );
or ( n225144 , n47380 , n225143 );
or ( n47384 , n47381 , n31180 );
nand ( n225146 , n225144 , n47384 );
and ( n225147 , n225146 , n42285 );
not ( n47387 , n225146 );
and ( n47388 , n47387 , n220896 );
nor ( n47389 , n225147 , n47388 );
not ( n47390 , n47389 );
not ( n47391 , n47390 );
and ( n47392 , n47379 , n47391 );
and ( n225154 , n47378 , n47390 );
nor ( n225155 , n47392 , n225154 );
not ( n47395 , n225155 );
buf ( n225157 , n32391 );
not ( n225158 , n225157 );
not ( n47398 , n36188 );
or ( n47399 , n225158 , n47398 );
or ( n47400 , n36188 , n225157 );
nand ( n47401 , n47399 , n47400 );
and ( n47402 , n47401 , n40178 );
not ( n47403 , n47401 );
not ( n225165 , n33524 );
buf ( n225166 , n225165 );
and ( n47406 , n47403 , n225166 );
nor ( n47407 , n47402 , n47406 );
buf ( n47408 , RI1745e920_1275);
not ( n47409 , n47408 );
not ( n47410 , n41668 );
or ( n47411 , n47409 , n47410 );
or ( n47412 , n41668 , n47408 );
nand ( n47413 , n47411 , n47412 );
and ( n225175 , n47413 , n223530 );
not ( n225176 , n47413 );
and ( n225177 , n225176 , n45773 );
nor ( n225178 , n225175 , n225177 );
nand ( n47418 , n47407 , n225178 );
not ( n47419 , n25675 );
not ( n47420 , n39896 );
and ( n47421 , n47419 , n47420 );
and ( n47422 , n25675 , n39896 );
nor ( n47423 , n47421 , n47422 );
xor ( n225185 , n25683 , n47423 );
and ( n225186 , n47418 , n225185 );
not ( n47426 , n47418 );
not ( n47427 , n225185 );
and ( n47428 , n47426 , n47427 );
nor ( n47429 , n225186 , n47428 );
not ( n47430 , n47429 );
or ( n47431 , n47395 , n47430 );
or ( n47432 , n47429 , n225155 );
nand ( n47433 , n47431 , n47432 );
buf ( n47434 , n29551 );
not ( n47435 , n47434 );
not ( n47436 , n47435 );
not ( n47437 , n38435 );
or ( n225199 , n47436 , n47437 );
not ( n225200 , n38435 );
nand ( n47440 , n225200 , n47434 );
nand ( n47441 , n225199 , n47440 );
not ( n47442 , n47441 );
not ( n47443 , n43735 );
or ( n47444 , n47442 , n47443 );
or ( n47445 , n33047 , n47441 );
nand ( n47446 , n47444 , n47445 );
not ( n47447 , n29582 );
not ( n225209 , n38908 );
or ( n225210 , n47447 , n225209 );
not ( n47450 , n38912 );
or ( n47451 , n47450 , n29582 );
nand ( n47452 , n225210 , n47451 );
not ( n47453 , n47452 );
not ( n47454 , n43473 );
and ( n47455 , n47453 , n47454 );
not ( n225217 , n43473 );
not ( n225218 , n225217 );
and ( n47458 , n47452 , n225218 );
nor ( n47459 , n47455 , n47458 );
nand ( n47460 , n47446 , n47459 );
xor ( n47461 , n204901 , n36018 );
xnor ( n225223 , n47461 , n34004 );
and ( n225224 , n47460 , n225223 );
not ( n47464 , n47460 );
not ( n47465 , n225223 );
and ( n47466 , n47464 , n47465 );
nor ( n47467 , n225224 , n47466 );
xor ( n225229 , n47433 , n47467 );
not ( n225230 , n225229 );
not ( n47470 , n225230 );
not ( n225232 , n225111 );
nand ( n225233 , n225232 , n47331 );
not ( n47473 , n225233 );
not ( n47474 , n205403 );
not ( n47475 , n39558 );
or ( n47476 , n47474 , n47475 );
or ( n47477 , n39558 , n205403 );
nand ( n225239 , n47476 , n47477 );
and ( n225240 , n225239 , n37303 );
not ( n47480 , n225239 );
and ( n47481 , n47480 , n36751 );
nor ( n225243 , n225240 , n47481 );
not ( n225244 , n225243 );
and ( n47484 , n47473 , n225244 );
nand ( n47485 , n47331 , n47354 );
and ( n47486 , n47485 , n225243 );
nor ( n47487 , n47484 , n47486 );
not ( n47488 , n47487 );
and ( n47489 , n33401 , n33398 );
not ( n225251 , n33401 );
buf ( n225252 , RI174a9038_912);
and ( n47492 , n225251 , n225252 );
nor ( n47493 , n47489 , n47492 );
not ( n47494 , n39267 );
xor ( n47495 , n47493 , n47494 );
xnor ( n225257 , n47495 , n38570 );
not ( n225258 , n33914 );
not ( n47498 , n204723 );
or ( n47499 , n225258 , n47498 );
or ( n47500 , n204727 , n33914 );
nand ( n47501 , n47499 , n47500 );
not ( n225263 , n47501 );
not ( n225264 , n36702 );
and ( n47504 , n225263 , n225264 );
and ( n47505 , n47501 , n204745 );
nor ( n47506 , n47504 , n47505 );
nand ( n47507 , n225257 , n47506 );
not ( n225269 , n32208 );
buf ( n225270 , n220278 );
not ( n47510 , n225270 );
or ( n47511 , n225269 , n47510 );
or ( n47512 , n225270 , n32208 );
nand ( n47513 , n47511 , n47512 );
and ( n47514 , n47513 , n221604 );
not ( n47515 , n47513 );
and ( n47516 , n47515 , n43839 );
nor ( n47517 , n47514 , n47516 );
and ( n225279 , n47507 , n47517 );
not ( n225280 , n47507 );
not ( n47520 , n47517 );
and ( n225282 , n225280 , n47520 );
nor ( n47522 , n225279 , n225282 );
not ( n225284 , n47522 );
or ( n225285 , n47488 , n225284 );
or ( n47525 , n47522 , n47487 );
nand ( n47526 , n225285 , n47525 );
buf ( n47527 , n47526 );
not ( n47528 , n47527 );
and ( n47529 , n47470 , n47528 );
and ( n47530 , n225230 , n47527 );
nor ( n47531 , n47529 , n47530 );
not ( n47532 , n47531 );
or ( n47533 , n225120 , n47532 );
not ( n47534 , n225119 );
not ( n47535 , n225229 );
not ( n225297 , n47526 );
not ( n225298 , n225297 );
or ( n47538 , n47535 , n225298 );
nand ( n47539 , n225230 , n47526 );
nand ( n225301 , n47538 , n47539 );
nand ( n225302 , n47534 , n225301 );
nand ( n47542 , n47533 , n225302 );
buf ( n47543 , n31197 );
not ( n47544 , n47543 );
not ( n47545 , n31425 );
or ( n47546 , n47544 , n47545 );
or ( n47547 , n31425 , n47543 );
nand ( n225309 , n47546 , n47547 );
and ( n225310 , n225309 , n220896 );
not ( n47550 , n225309 );
and ( n47551 , n47550 , n42285 );
nor ( n47552 , n225310 , n47551 );
not ( n47553 , n40024 );
not ( n47554 , n30936 );
or ( n47555 , n47553 , n47554 );
or ( n47556 , n30936 , n40024 );
nand ( n47557 , n47555 , n47556 );
and ( n225319 , n47557 , n30897 );
not ( n225320 , n47557 );
not ( n47560 , n205033 );
not ( n47561 , n47560 );
and ( n47562 , n225320 , n47561 );
nor ( n47563 , n225319 , n47562 );
nor ( n47564 , n47552 , n47563 );
xor ( n47565 , n28545 , n30781 );
xnor ( n47566 , n47565 , n37407 );
not ( n225328 , n47566 );
and ( n225329 , n47564 , n225328 );
not ( n225330 , n47564 );
and ( n225331 , n225330 , n47566 );
nor ( n47571 , n225329 , n225331 );
not ( n47572 , n47571 );
not ( n47573 , n47572 );
not ( n47574 , n39943 );
not ( n47575 , n206425 );
or ( n47576 , n47574 , n47575 );
or ( n47577 , n206425 , n39943 );
nand ( n47578 , n47576 , n47577 );
and ( n225340 , n47578 , n28646 );
not ( n225341 , n47578 );
buf ( n47581 , n38747 );
and ( n225343 , n225341 , n47581 );
nor ( n225344 , n225340 , n225343 );
not ( n47584 , n225344 );
not ( n47585 , n30632 );
not ( n47586 , n39922 );
or ( n47587 , n47585 , n47586 );
not ( n47588 , n30632 );
nand ( n47589 , n47588 , n39921 );
nand ( n225351 , n47587 , n47589 );
not ( n225352 , n45239 );
not ( n47592 , RI17359008_2091);
not ( n47593 , n47592 );
or ( n47594 , n225352 , n47593 );
not ( n47595 , RI173d15c0_1735);
nand ( n47596 , n47595 , n44182 );
nand ( n47597 , n47594 , n47596 );
not ( n225359 , RI17449098_1380);
and ( n225360 , n47597 , n225359 );
not ( n47600 , n47597 );
buf ( n47601 , RI17449098_1380);
and ( n47602 , n47600 , n47601 );
nor ( n47603 , n225360 , n47602 );
xor ( n47604 , n47603 , n28841 );
xnor ( n47605 , n47604 , n45558 );
buf ( n47606 , n47605 );
not ( n47607 , n47606 );
and ( n47608 , n225351 , n47607 );
not ( n47609 , n225351 );
not ( n225371 , n47606 );
not ( n225372 , n225371 );
buf ( n47612 , n225372 );
and ( n47613 , n47609 , n47612 );
nor ( n47614 , n47608 , n47613 );
nand ( n47615 , n47584 , n47614 );
not ( n47616 , n47615 );
not ( n47617 , n25848 );
buf ( n225379 , n37579 );
xor ( n225380 , n47617 , n225379 );
xnor ( n47620 , n225380 , n38839 );
not ( n225382 , n47620 );
or ( n225383 , n47616 , n225382 );
nand ( n47623 , n47584 , n47614 );
or ( n47624 , n47620 , n47623 );
nand ( n47625 , n225383 , n47624 );
not ( n47626 , n47625 );
not ( n225388 , n47626 );
or ( n225389 , n47573 , n225388 );
nand ( n47629 , n47625 , n47571 );
nand ( n47630 , n225389 , n47629 );
not ( n47631 , n47630 );
buf ( n47632 , n29605 );
not ( n47633 , n47632 );
not ( n47634 , n38911 );
or ( n47635 , n47633 , n47634 );
or ( n47636 , n38911 , n47632 );
nand ( n47637 , n47635 , n47636 );
and ( n47638 , n47637 , n225217 );
not ( n47639 , n47637 );
and ( n47640 , n47639 , n43469 );
nor ( n47641 , n47638 , n47640 );
not ( n225403 , n47641 );
buf ( n225404 , n33361 );
not ( n47644 , n225404 );
not ( n47645 , n30580 );
or ( n47646 , n47644 , n47645 );
or ( n47647 , n30580 , n225404 );
nand ( n47648 , n47646 , n47647 );
and ( n47649 , n47648 , n39558 );
not ( n47650 , n47648 );
and ( n47651 , n47650 , n39559 );
nor ( n225413 , n47649 , n47651 );
not ( n225414 , n33404 );
not ( n47654 , n29383 );
not ( n47655 , n40369 );
or ( n47656 , n47654 , n47655 );
or ( n47657 , n40369 , n29383 );
nand ( n47658 , n47656 , n47657 );
not ( n47659 , n47658 );
or ( n47660 , n225414 , n47659 );
or ( n47661 , n33404 , n47658 );
nand ( n225423 , n47660 , n47661 );
nand ( n225424 , n225413 , n225423 );
not ( n47664 , n225424 );
or ( n47665 , n225403 , n47664 );
or ( n47666 , n225424 , n47641 );
nand ( n47667 , n47665 , n47666 );
not ( n225429 , n47667 );
not ( n225430 , n31735 );
not ( n47670 , n33925 );
not ( n47671 , n204726 );
or ( n47672 , n47670 , n47671 );
not ( n47673 , n43269 );
or ( n225435 , n43589 , n47673 );
nand ( n225436 , n47672 , n225435 );
not ( n47676 , n225436 );
and ( n225438 , n225430 , n47676 );
and ( n225439 , n36705 , n225436 );
nor ( n47679 , n225438 , n225439 );
not ( n47680 , n224443 );
not ( n47681 , n42764 );
not ( n47682 , n216052 );
or ( n47683 , n47681 , n47682 );
or ( n47684 , n216052 , n42764 );
nand ( n225446 , n47683 , n47684 );
not ( n225447 , n225446 );
or ( n47687 , n47680 , n225447 );
or ( n47688 , n225446 , n204936 );
nand ( n47689 , n47687 , n47688 );
nand ( n225451 , n47679 , n47689 );
not ( n225452 , n225451 );
not ( n47692 , n36158 );
not ( n47693 , n38347 );
or ( n47694 , n47692 , n47693 );
not ( n47695 , n36158 );
not ( n47696 , n38322 );
xor ( n47697 , n38342 , n47696 );
xnor ( n225459 , n47697 , n37893 );
nand ( n225460 , n47695 , n225459 );
nand ( n47700 , n47694 , n225460 );
not ( n47701 , n47700 );
not ( n47702 , n38353 );
and ( n47703 , n47701 , n47702 );
not ( n47704 , n44887 );
and ( n47705 , n47700 , n47704 );
nor ( n225467 , n47703 , n47705 );
not ( n225468 , n225467 );
not ( n47708 , n225468 );
and ( n47709 , n225452 , n47708 );
and ( n47710 , n225451 , n225468 );
nor ( n47711 , n47709 , n47710 );
not ( n225473 , n47711 );
or ( n225474 , n225429 , n225473 );
or ( n47714 , n47711 , n47667 );
nand ( n47715 , n225474 , n47714 );
not ( n47716 , n39478 );
not ( n47717 , n37507 );
or ( n47718 , n47716 , n47717 );
not ( n47719 , n39478 );
nand ( n225481 , n47719 , n37506 );
nand ( n225482 , n47718 , n225481 );
buf ( n47722 , n39875 );
xor ( n47723 , n225482 , n47722 );
not ( n47724 , n35229 );
not ( n47725 , n34992 );
not ( n225487 , n25550 );
or ( n225488 , n47725 , n225487 );
or ( n47728 , n25550 , n34992 );
nand ( n47729 , n225488 , n47728 );
not ( n47730 , n47729 );
or ( n47731 , n47724 , n47730 );
or ( n47732 , n47729 , n35229 );
nand ( n47733 , n47731 , n47732 );
nand ( n225495 , n47723 , n47733 );
not ( n225496 , n225495 );
not ( n47736 , n29366 );
not ( n47737 , n29369 );
or ( n47738 , n47736 , n47737 );
or ( n47739 , n29369 , n29366 );
nand ( n225501 , n47738 , n47739 );
not ( n225502 , n225501 );
not ( n47742 , n31514 );
or ( n47743 , n225502 , n47742 );
not ( n47744 , n225501 );
nand ( n47745 , n47744 , n31527 );
nand ( n47746 , n47743 , n47745 );
and ( n47747 , n47746 , n33853 );
not ( n225509 , n47746 );
and ( n225510 , n225509 , n33849 );
nor ( n47750 , n47747 , n225510 );
buf ( n225512 , n47750 );
not ( n47752 , n225512 );
and ( n225514 , n225496 , n47752 );
and ( n225515 , n225495 , n225512 );
nor ( n47755 , n225514 , n225515 );
and ( n225517 , n47715 , n47755 );
not ( n225518 , n47715 );
not ( n47758 , n47755 );
and ( n47759 , n225518 , n47758 );
nor ( n47760 , n225517 , n47759 );
not ( n47761 , n47760 );
and ( n47762 , n47631 , n47761 );
and ( n47763 , n47630 , n47760 );
nor ( n225525 , n47762 , n47763 );
and ( n225526 , n47542 , n225525 );
not ( n47766 , n47542 );
not ( n47767 , n47760 );
not ( n47768 , n47630 );
or ( n47769 , n47767 , n47768 );
not ( n47770 , n47630 );
not ( n47771 , n47760 );
nand ( n47772 , n47770 , n47771 );
nand ( n47773 , n47769 , n47772 );
not ( n225535 , n47773 );
not ( n225536 , n225535 );
and ( n47776 , n47766 , n225536 );
nor ( n47777 , n225526 , n47776 );
nand ( n47778 , n47327 , n47777 );
buf ( n47779 , n207783 );
xor ( n47780 , n47779 , n35926 );
xnor ( n47781 , n47780 , n39569 );
not ( n47782 , n47781 );
not ( n47783 , n36635 );
not ( n47784 , n35200 );
or ( n47785 , n47783 , n47784 );
nand ( n225547 , n35199 , n36631 );
nand ( n225548 , n47785 , n225547 );
not ( n47788 , n225548 );
not ( n225550 , n205322 );
and ( n225551 , n47788 , n225550 );
and ( n47791 , n225548 , n205322 );
nor ( n47792 , n225551 , n47791 );
not ( n47793 , n47792 );
nand ( n47794 , n47782 , n47793 );
not ( n47795 , RI174a96c8_910);
and ( n47796 , n37190 , n47795 );
not ( n47797 , n37190 );
and ( n47798 , n47797 , n37187 );
nor ( n225560 , n47796 , n47798 );
xor ( n225561 , n225560 , n28043 );
xnor ( n47801 , n225561 , n205230 );
and ( n225563 , n47794 , n47801 );
not ( n225564 , n47794 );
not ( n47804 , n47801 );
and ( n47805 , n225564 , n47804 );
nor ( n47806 , n225563 , n47805 );
not ( n47807 , n47806 );
not ( n47808 , n47807 );
not ( n47809 , n37396 );
not ( n47810 , n222183 );
or ( n225572 , n47809 , n47810 );
not ( n225573 , n37396 );
nand ( n47813 , n225573 , n39359 );
nand ( n47814 , n225572 , n47813 );
not ( n47815 , n47814 );
not ( n47816 , n38877 );
not ( n47817 , n47816 );
and ( n47818 , n47815 , n47817 );
and ( n225580 , n47814 , n45465 );
nor ( n225581 , n47818 , n225580 );
not ( n47821 , n41055 );
buf ( n47822 , n26354 );
not ( n47823 , n29872 );
not ( n47824 , n32987 );
or ( n47825 , n47823 , n47824 );
or ( n47826 , n29872 , n32987 );
nand ( n47827 , n47825 , n47826 );
not ( n47828 , n32978 );
and ( n47829 , n47827 , n47828 );
not ( n47830 , n47827 );
and ( n47831 , n47830 , n32978 );
nor ( n225593 , n47829 , n47831 );
and ( n225594 , n47822 , n225593 );
not ( n47834 , n47822 );
and ( n225596 , n47834 , n32988 );
nor ( n225597 , n225594 , n225596 );
not ( n47837 , n225597 );
not ( n47838 , n47837 );
or ( n47839 , n47821 , n47838 );
nand ( n47840 , n225597 , n45696 );
nand ( n47841 , n47839 , n47840 );
nand ( n47842 , n225581 , n47841 );
not ( n225604 , n47842 );
not ( n225605 , n35684 );
not ( n47845 , n39968 );
or ( n225607 , n225605 , n47845 );
or ( n225608 , n39968 , n35684 );
nand ( n47848 , n225607 , n225608 );
and ( n47849 , n47848 , n40007 );
not ( n47850 , n47848 );
and ( n47851 , n47850 , n40006 );
nor ( n47852 , n47849 , n47851 );
not ( n47853 , n47852 );
not ( n47854 , n47853 );
and ( n47855 , n225604 , n47854 );
and ( n47856 , n47842 , n47853 );
nor ( n47857 , n47855 , n47856 );
not ( n225619 , n47857 );
buf ( n225620 , n204802 );
not ( n47860 , n225620 );
not ( n225622 , n205072 );
or ( n225623 , n47860 , n225622 );
or ( n47863 , n205072 , n225620 );
nand ( n47864 , n225623 , n47863 );
and ( n47865 , n47864 , n33183 );
not ( n47866 , n47864 );
and ( n47867 , n47866 , n43757 );
nor ( n47868 , n47865 , n47867 );
not ( n225630 , n47868 );
buf ( n225631 , n38905 );
not ( n47871 , n225631 );
buf ( n47872 , RI174146b8_1408);
xor ( n47873 , n47872 , n26214 );
xor ( n47874 , n47873 , n26221 );
not ( n47875 , n47874 );
or ( n47876 , n47871 , n47875 );
or ( n225638 , n47874 , n225631 );
nand ( n225639 , n47876 , n225638 );
buf ( n47879 , n40224 );
and ( n47880 , n225639 , n47879 );
not ( n47881 , n225639 );
and ( n47882 , n47881 , n26205 );
nor ( n225644 , n47880 , n47882 );
nand ( n225645 , n225630 , n225644 );
not ( n47885 , n32221 );
not ( n47886 , n37346 );
or ( n47887 , n47885 , n47886 );
not ( n47888 , n32221 );
nand ( n47889 , n47888 , n43837 );
nand ( n47890 , n47887 , n47889 );
and ( n225652 , n47890 , n37353 );
not ( n225653 , n47890 );
and ( n47893 , n225653 , n37356 );
nor ( n47894 , n225652 , n47893 );
and ( n225656 , n225645 , n47894 );
not ( n225657 , n225645 );
not ( n47897 , n47894 );
and ( n47898 , n225657 , n47897 );
nor ( n47899 , n225656 , n47898 );
not ( n47900 , n47899 );
or ( n47901 , n225619 , n47900 );
or ( n225663 , n47899 , n47857 );
nand ( n225664 , n47901 , n225663 );
buf ( n47904 , n29005 );
not ( n47905 , n47904 );
not ( n47906 , n31263 );
or ( n47907 , n47905 , n47906 );
or ( n47908 , n31263 , n47904 );
nand ( n47909 , n47907 , n47908 );
and ( n47910 , n47909 , n30321 );
not ( n47911 , n47909 );
and ( n225673 , n47911 , n35169 );
nor ( n225674 , n47910 , n225673 );
not ( n47914 , n225674 );
not ( n225676 , n26203 );
not ( n225677 , n225676 );
not ( n47917 , n36626 );
or ( n225679 , n225677 , n47917 );
nand ( n225680 , n36620 , n26203 );
nand ( n47920 , n225679 , n225680 );
not ( n225682 , n46586 );
buf ( n225683 , n225682 );
not ( n47923 , n225683 );
and ( n47924 , n47920 , n47923 );
not ( n47925 , n47920 );
and ( n47926 , n47925 , n225683 );
nor ( n225688 , n47924 , n47926 );
nand ( n225689 , n47914 , n225688 );
not ( n47929 , n225689 );
not ( n225691 , n40963 );
not ( n225692 , n38109 );
and ( n47932 , n225691 , n225692 );
and ( n47933 , n39417 , n38109 );
nor ( n225695 , n47932 , n47933 );
not ( n225696 , n40111 );
not ( n47936 , n40131 );
or ( n47937 , n225696 , n47936 );
nand ( n47938 , n47937 , n40135 );
not ( n47939 , n47938 );
and ( n47940 , n225695 , n47939 );
not ( n47941 , n225695 );
and ( n47942 , n47941 , n47938 );
nor ( n47943 , n47940 , n47942 );
not ( n225705 , n47943 );
and ( n225706 , n47929 , n225705 );
and ( n47946 , n225689 , n47943 );
nor ( n47947 , n225706 , n47946 );
and ( n47948 , n225664 , n47947 );
not ( n47949 , n225664 );
not ( n47950 , n47947 );
and ( n47951 , n47949 , n47950 );
nor ( n225713 , n47948 , n47951 );
buf ( n225714 , n225713 );
not ( n47954 , n225714 );
xor ( n225716 , n27911 , n36380 );
xnor ( n225717 , n225716 , n36258 );
not ( n47957 , n25619 );
not ( n47958 , n40101 );
not ( n47959 , n47958 );
or ( n47960 , n47957 , n47959 );
not ( n47961 , n25619 );
nand ( n47962 , n47961 , n40101 );
nand ( n47963 , n47960 , n47962 );
not ( n47964 , n37652 );
and ( n225726 , n47963 , n47964 );
not ( n225727 , n47963 );
and ( n47967 , n225727 , n45268 );
nor ( n47968 , n225726 , n47967 );
nand ( n47969 , n225717 , n47968 );
not ( n47970 , n47969 );
not ( n47971 , n47704 );
not ( n47972 , n213927 );
not ( n47973 , n225459 );
or ( n47974 , n47972 , n47973 );
not ( n225736 , n213927 );
nand ( n225737 , n225736 , n38347 );
nand ( n225738 , n47974 , n225737 );
not ( n225739 , n225738 );
or ( n47979 , n47971 , n225739 );
or ( n225741 , n225738 , n38356 );
nand ( n225742 , n47979 , n225741 );
buf ( n47982 , n225742 );
not ( n47983 , n47982 );
and ( n47984 , n47970 , n47983 );
not ( n47985 , n47968 );
not ( n47986 , n47985 );
nand ( n47987 , n47986 , n225717 );
and ( n47988 , n47987 , n47982 );
nor ( n47989 , n47984 , n47988 );
not ( n47990 , n47989 );
not ( n47991 , n47990 );
nand ( n225753 , n47801 , n47781 );
not ( n225754 , n29941 );
not ( n47994 , n32909 );
or ( n225756 , n225754 , n47994 );
nand ( n225757 , n32910 , n29938 );
nand ( n47997 , n225756 , n225757 );
and ( n47998 , n47997 , n204258 );
not ( n47999 , n47997 );
and ( n48000 , n47999 , n204259 );
nor ( n225762 , n47998 , n48000 );
not ( n225763 , n225762 );
and ( n48003 , n225753 , n225763 );
not ( n48004 , n225753 );
and ( n48005 , n48004 , n225762 );
nor ( n48006 , n48003 , n48005 );
not ( n48007 , n48006 );
not ( n48008 , n48007 );
or ( n225770 , n47991 , n48008 );
nand ( n225771 , n48006 , n47989 );
nand ( n48011 , n225770 , n225771 );
not ( n48012 , n48011 );
or ( n48013 , n47954 , n48012 );
or ( n48014 , n48011 , n225714 );
nand ( n48015 , n48013 , n48014 );
not ( n48016 , n48015 );
or ( n225778 , n47808 , n48016 );
not ( n225779 , n47807 );
xor ( n48019 , n48011 , n225713 );
nand ( n225781 , n225779 , n48019 );
nand ( n225782 , n225778 , n225781 );
not ( n48022 , n204820 );
not ( n48023 , n42258 );
and ( n48024 , n48022 , n48023 );
and ( n48025 , n204820 , n42258 );
nor ( n48026 , n48024 , n48025 );
not ( n48027 , n48026 );
not ( n48028 , n204812 );
or ( n48029 , n48027 , n48028 );
or ( n48030 , n204812 , n48026 );
nand ( n48031 , n48029 , n48030 );
and ( n225793 , n48031 , n204792 );
not ( n225794 , n48031 );
and ( n48034 , n225794 , n223504 );
nor ( n225796 , n225793 , n48034 );
not ( n225797 , RI173cda98_1753);
xor ( n48037 , n225797 , n41241 );
xnor ( n48038 , n48037 , n41256 );
not ( n48039 , n48038 );
not ( n48040 , n48039 );
not ( n48041 , n34029 );
not ( n48042 , n41303 );
or ( n225804 , n48041 , n48042 );
or ( n225805 , n41303 , n34029 );
nand ( n48045 , n225804 , n225805 );
not ( n48046 , n48045 );
or ( n48047 , n48040 , n48046 );
or ( n48048 , n48045 , n41258 );
nand ( n48049 , n48047 , n48048 );
nand ( n48050 , n225796 , n48049 );
not ( n225812 , n48050 );
not ( n225813 , n28246 );
not ( n48053 , n36237 );
or ( n48054 , n225813 , n48053 );
not ( n48055 , n28246 );
nand ( n48056 , n48055 , n36242 );
nand ( n48057 , n48054 , n48056 );
not ( n48058 , n45215 );
and ( n225820 , n48057 , n48058 );
not ( n225821 , n48057 );
not ( n48061 , n45218 );
and ( n48062 , n225821 , n48061 );
nor ( n48063 , n225820 , n48062 );
not ( n48064 , n48063 );
not ( n48065 , n48064 );
and ( n225827 , n225812 , n48065 );
and ( n225828 , n48050 , n48064 );
nor ( n225829 , n225827 , n225828 );
not ( n225830 , n225829 );
not ( n48070 , n36286 );
xor ( n48071 , n36303 , n48070 );
buf ( n48072 , n36277 );
xnor ( n48073 , n48071 , n48072 );
xor ( n225835 , n28307 , n48073 );
not ( n225836 , n36347 );
xnor ( n48076 , n225835 , n225836 );
not ( n48077 , n48076 );
not ( n48078 , n25693 );
not ( n48079 , n208349 );
or ( n48080 , n48078 , n48079 );
or ( n225842 , n208349 , n25693 );
nand ( n225843 , n48080 , n225842 );
not ( n48083 , n225843 );
not ( n48084 , n30602 );
or ( n48085 , n48083 , n48084 );
or ( n48086 , n30602 , n225843 );
nand ( n225848 , n48085 , n48086 );
not ( n225849 , n225848 );
not ( n48089 , n30580 );
and ( n48090 , n225849 , n48089 );
and ( n48091 , n225848 , n39554 );
nor ( n48092 , n48090 , n48091 );
nand ( n48093 , n48077 , n48092 );
not ( n48094 , n29690 );
not ( n48095 , n34733 );
or ( n225857 , n48094 , n48095 );
nand ( n225858 , n34710 , n29677 );
nand ( n48098 , n225857 , n225858 );
not ( n48099 , n48098 );
buf ( n48100 , n34729 );
not ( n48101 , n48100 );
or ( n225863 , n48099 , n48101 );
or ( n225864 , n48100 , n48098 );
nand ( n48104 , n225863 , n225864 );
and ( n225866 , n48104 , n34700 );
not ( n225867 , n48104 );
and ( n48107 , n225867 , n39850 );
nor ( n225869 , n225866 , n48107 );
and ( n225870 , n48093 , n225869 );
not ( n48110 , n48093 );
not ( n48111 , n225869 );
and ( n48112 , n48110 , n48111 );
nor ( n48113 , n225870 , n48112 );
not ( n48114 , n48113 );
or ( n48115 , n225830 , n48114 );
or ( n48116 , n48113 , n225829 );
nand ( n48117 , n48115 , n48116 );
not ( n48118 , n40872 );
not ( n48119 , n42966 );
or ( n225881 , n48118 , n48119 );
not ( n225882 , n40872 );
nand ( n48122 , n225882 , n38657 );
nand ( n48123 , n225881 , n48122 );
and ( n48124 , n48123 , n38677 );
not ( n48125 , n48123 );
and ( n225887 , n48125 , n38662 );
nor ( n225888 , n48124 , n225887 );
not ( n48128 , n28394 );
not ( n48129 , n39007 );
or ( n48130 , n48128 , n48129 );
nand ( n48131 , n39002 , n28390 );
nand ( n48132 , n48130 , n48131 );
not ( n48133 , n48132 );
not ( n225895 , n41857 );
and ( n225896 , n48133 , n225895 );
and ( n48136 , n48132 , n41857 );
nor ( n48137 , n225896 , n48136 );
nand ( n48138 , n225888 , n48137 );
not ( n48139 , n48138 );
not ( n225901 , n204259 );
not ( n225902 , n37775 );
not ( n48142 , n32906 );
or ( n48143 , n225902 , n48142 );
not ( n48144 , n37775 );
nand ( n48145 , n48144 , n32910 );
nand ( n225907 , n48143 , n48145 );
not ( n225908 , n225907 );
or ( n48148 , n225901 , n225908 );
or ( n48149 , n204259 , n225907 );
nand ( n48150 , n48148 , n48149 );
not ( n48151 , n48150 );
and ( n225913 , n48139 , n48151 );
and ( n225914 , n48138 , n48150 );
nor ( n48154 , n225913 , n225914 );
and ( n48155 , n48117 , n48154 );
not ( n48156 , n48117 );
not ( n48157 , n48154 );
and ( n225919 , n48156 , n48157 );
nor ( n225920 , n48155 , n225919 );
not ( n48160 , n225920 );
not ( n48161 , n48160 );
not ( n48162 , n31486 );
not ( n48163 , n38690 );
or ( n225925 , n48162 , n48163 );
not ( n225926 , n31486 );
nand ( n48166 , n225926 , n38691 );
nand ( n48167 , n225925 , n48166 );
not ( n48168 , n48167 );
not ( n48169 , n38795 );
and ( n48170 , n48168 , n48169 );
and ( n48171 , n48167 , n38795 );
nor ( n48172 , n48170 , n48171 );
not ( n48173 , n33869 );
buf ( n48174 , n205219 );
not ( n48175 , n48174 );
or ( n225937 , n48173 , n48175 );
not ( n225938 , n33869 );
nand ( n48178 , n225938 , n205215 );
nand ( n48179 , n225937 , n48178 );
not ( n48180 , n43910 );
and ( n48181 , n48179 , n48180 );
not ( n48182 , n48179 );
and ( n48183 , n48182 , n43914 );
nor ( n48184 , n48181 , n48183 );
nand ( n48185 , n48172 , n48184 );
not ( n225947 , n48185 );
not ( n225948 , n42174 );
not ( n48188 , n225948 );
xor ( n48189 , n41147 , n48188 );
xnor ( n48190 , n48189 , n205436 );
not ( n48191 , n48190 );
not ( n225953 , n48191 );
or ( n225954 , n225947 , n225953 );
or ( n48194 , n48191 , n48185 );
nand ( n225956 , n225954 , n48194 );
not ( n225957 , n225956 );
not ( n48197 , n225957 );
xor ( n48198 , n30847 , n45371 );
xnor ( n48199 , n48198 , n35107 );
not ( n48200 , n48199 );
not ( n48201 , n48200 );
not ( n48202 , n41594 );
xor ( n48203 , n34846 , n34264 );
not ( n225965 , n48203 );
or ( n225966 , n48202 , n225965 );
or ( n48206 , n48203 , n41594 );
nand ( n48207 , n225966 , n48206 );
not ( n48208 , n36785 );
not ( n48209 , n42623 );
or ( n48210 , n48208 , n48209 );
nand ( n48211 , n42624 , n36781 );
nand ( n48212 , n48210 , n48211 );
not ( n225974 , n48212 );
not ( n225975 , n45817 );
and ( n48215 , n225974 , n225975 );
and ( n48216 , n48212 , n45817 );
nor ( n48217 , n48215 , n48216 );
nor ( n48218 , n48207 , n48217 );
not ( n225980 , n48218 );
and ( n225981 , n48201 , n225980 );
and ( n48221 , n48200 , n48218 );
nor ( n48222 , n225981 , n48221 );
not ( n48223 , n48222 );
not ( n48224 , n48223 );
or ( n225986 , n48197 , n48224 );
nand ( n225987 , n48222 , n225956 );
nand ( n48227 , n225986 , n225987 );
not ( n225989 , n48227 );
not ( n225990 , n225989 );
or ( n48230 , n48161 , n225990 );
nand ( n48231 , n225920 , n48227 );
nand ( n48232 , n48230 , n48231 );
not ( n48233 , n48232 );
not ( n48234 , n48233 );
and ( n48235 , n225782 , n48234 );
not ( n225997 , n225782 );
buf ( n225998 , n48232 );
not ( n48238 , n225998 );
and ( n226000 , n225997 , n48238 );
nor ( n226001 , n48235 , n226000 );
not ( n48241 , n226001 );
buf ( n226003 , n27886 );
buf ( n226004 , n226003 );
nor ( n48244 , n48241 , n226004 );
not ( n48245 , n48244 );
or ( n48246 , n47778 , n48245 );
nand ( n48247 , n226001 , n47777 );
not ( n48248 , n47327 );
buf ( n226010 , n222531 );
nand ( n226011 , n48247 , n48248 , n226010 );
buf ( n48251 , n35431 );
nand ( n48252 , n48251 , n38166 );
nand ( n48253 , n48246 , n226011 , n48252 );
buf ( n48254 , n48253 );
not ( n48255 , n225138 );
nand ( n48256 , n48255 , n47389 );
not ( n48257 , n36599 );
not ( n226019 , n38817 );
or ( n226020 , n48257 , n226019 );
not ( n48260 , n36599 );
nand ( n48261 , n48260 , n38823 );
nand ( n48262 , n226020 , n48261 );
and ( n48263 , n48262 , n38830 );
not ( n48264 , n48262 );
and ( n48265 , n48264 , n38826 );
nor ( n48266 , n48263 , n48265 );
not ( n48267 , n48266 );
and ( n48268 , n48256 , n48267 );
not ( n48269 , n48256 );
and ( n226031 , n48269 , n48266 );
nor ( n226032 , n48268 , n226031 );
buf ( n48272 , n226032 );
not ( n226034 , n48272 );
not ( n226035 , n42942 );
not ( n48275 , n43261 );
or ( n226037 , n226035 , n48275 );
not ( n226038 , n42942 );
nand ( n48278 , n226038 , n45225 );
nand ( n226040 , n226037 , n48278 );
and ( n226041 , n226040 , n42675 );
not ( n48281 , n226040 );
and ( n48282 , n48281 , n45230 );
nor ( n48283 , n226041 , n48282 );
not ( n48284 , n48283 );
nand ( n48285 , n47427 , n48284 );
not ( n48286 , n30941 );
not ( n48287 , n48286 );
not ( n48288 , n47013 );
not ( n48289 , n48288 );
or ( n48290 , n48287 , n48289 );
not ( n48291 , n218655 );
or ( n226053 , n48291 , n48286 );
nand ( n226054 , n48290 , n226053 );
and ( n48294 , n226054 , n32053 );
not ( n48295 , n226054 );
and ( n48296 , n48295 , n32050 );
nor ( n48297 , n48294 , n48296 );
not ( n48298 , n48297 );
not ( n48299 , n48298 );
and ( n226061 , n48285 , n48299 );
not ( n226062 , n48285 );
and ( n48302 , n226062 , n48298 );
nor ( n48303 , n226061 , n48302 );
nand ( n48304 , n48266 , n47390 );
not ( n48305 , n48304 );
not ( n48306 , n32671 );
xor ( n48307 , n45298 , n45306 );
xor ( n48308 , n48307 , n30649 );
not ( n48309 , n48308 );
or ( n48310 , n48306 , n48309 );
not ( n48311 , n32671 );
not ( n48312 , n48308 );
nand ( n226074 , n48311 , n48312 );
nand ( n226075 , n48310 , n226074 );
and ( n48315 , n226075 , n37996 );
not ( n48316 , n226075 );
buf ( n48317 , n37991 );
and ( n48318 , n48316 , n48317 );
nor ( n48319 , n48315 , n48318 );
not ( n48320 , n48319 );
and ( n48321 , n48305 , n48320 );
and ( n48322 , n48304 , n48319 );
nor ( n226084 , n48321 , n48322 );
or ( n226085 , n48303 , n226084 );
nand ( n48325 , n226084 , n48303 );
nand ( n226087 , n226085 , n48325 );
buf ( n226088 , n218484 );
not ( n48328 , n226088 );
not ( n48329 , n26050 );
or ( n48330 , n48328 , n48329 );
not ( n48331 , n26047 );
or ( n226093 , n48331 , n226088 );
nand ( n226094 , n48330 , n226093 );
not ( n48334 , n226094 );
not ( n226096 , n26009 );
and ( n226097 , n48334 , n226096 );
and ( n48337 , n26009 , n226094 );
nor ( n226099 , n226097 , n48337 );
not ( n226100 , n226099 );
not ( n48340 , n226100 );
not ( n48341 , n35048 );
not ( n48342 , n204671 );
or ( n48343 , n48341 , n48342 );
or ( n48344 , n204671 , n35048 );
nand ( n48345 , n48343 , n48344 );
and ( n48346 , n48345 , n26261 );
not ( n48347 , n48345 );
and ( n226109 , n48347 , n204681 );
nor ( n226110 , n48346 , n226109 );
buf ( n48350 , n226110 );
nand ( n48351 , n47465 , n48350 );
not ( n48352 , n48351 );
or ( n48353 , n48340 , n48352 );
nand ( n48354 , n47465 , n226099 , n48350 );
nand ( n48355 , n48353 , n48354 );
and ( n226117 , n226087 , n48355 );
not ( n226118 , n226087 );
not ( n48358 , n48355 );
and ( n48359 , n226118 , n48358 );
nor ( n48360 , n226117 , n48359 );
not ( n48361 , n39707 );
buf ( n226123 , n32718 );
not ( n226124 , n226123 );
and ( n48364 , n48361 , n226124 );
and ( n226126 , n39707 , n226123 );
nor ( n226127 , n48364 , n226126 );
and ( n48367 , n226127 , n36377 );
not ( n48368 , n226127 );
and ( n48369 , n48368 , n44006 );
nor ( n48370 , n48367 , n48369 );
not ( n226132 , n48370 );
not ( n226133 , n226132 );
and ( n48373 , n205157 , n204439 );
not ( n48374 , n205157 );
and ( n48375 , n48374 , n204436 );
nor ( n48376 , n48373 , n48375 );
and ( n48377 , n48376 , n204391 );
not ( n48378 , n48376 );
and ( n48379 , n48378 , n34477 );
nor ( n48380 , n48377 , n48379 );
nor ( n48381 , n47517 , n48380 );
not ( n48382 , n48381 );
and ( n226144 , n226133 , n48382 );
and ( n226145 , n48381 , n226132 );
nor ( n48385 , n226144 , n226145 );
not ( n226147 , n48385 );
not ( n226148 , n226147 );
not ( n48388 , n33417 );
not ( n48389 , n39845 );
or ( n48390 , n48388 , n48389 );
or ( n48391 , n39845 , n33417 );
nand ( n48392 , n48390 , n48391 );
and ( n48393 , n48392 , n32363 );
not ( n226155 , n48392 );
not ( n226156 , n32363 );
and ( n48396 , n226155 , n226156 );
nor ( n48397 , n48393 , n48396 );
nand ( n48398 , n48397 , n225243 );
not ( n48399 , n48398 );
not ( n48400 , n47338 );
or ( n48401 , n48399 , n48400 );
or ( n226163 , n47338 , n48398 );
nand ( n226164 , n48401 , n226163 );
not ( n48404 , n226164 );
not ( n48405 , n48404 );
or ( n48406 , n226148 , n48405 );
nand ( n48407 , n226164 , n48385 );
nand ( n226169 , n48406 , n48407 );
not ( n226170 , n226169 );
and ( n48410 , n48360 , n226170 );
not ( n48411 , n48360 );
and ( n48412 , n48411 , n226169 );
nor ( n48413 , n48410 , n48412 );
not ( n48414 , n48413 );
not ( n48415 , n48414 );
or ( n226177 , n226034 , n48415 );
or ( n226178 , n48414 , n48272 );
nand ( n48418 , n226177 , n226178 );
not ( n48419 , n26183 );
not ( n48420 , n36626 );
or ( n48421 , n48419 , n48420 );
not ( n226183 , n26183 );
nand ( n226184 , n226183 , n36618 );
nand ( n48424 , n48421 , n226184 );
and ( n226186 , n48424 , n225683 );
not ( n226187 , n48424 );
buf ( n48427 , n46587 );
not ( n48428 , n48427 );
and ( n48429 , n226187 , n48428 );
nor ( n48430 , n226186 , n48429 );
not ( n48431 , n48430 );
nand ( n48432 , n48431 , n225468 );
not ( n226194 , n48432 );
not ( n226195 , n226194 );
xor ( n48435 , n39215 , n45799 );
xnor ( n48436 , n48435 , n28405 );
not ( n48437 , n48436 );
or ( n48438 , n226195 , n48437 );
not ( n226200 , n48436 );
nand ( n226201 , n226200 , n48432 );
nand ( n48441 , n48438 , n226201 );
not ( n226203 , n29538 );
not ( n226204 , n38435 );
or ( n48444 , n226203 , n226204 );
or ( n48445 , n38435 , n29538 );
nand ( n48446 , n48444 , n48445 );
not ( n48447 , n48446 );
not ( n48448 , n43735 );
or ( n48449 , n48447 , n48448 );
or ( n48450 , n33047 , n48446 );
nand ( n48451 , n48449 , n48450 );
not ( n48452 , n48451 );
nand ( n48453 , n48452 , n47620 );
not ( n226215 , n48453 );
not ( n226216 , n205068 );
buf ( n48456 , RI173d6b10_1709);
not ( n226218 , n48456 );
and ( n226219 , n226216 , n226218 );
and ( n48459 , n205068 , n48456 );
nor ( n48460 , n226219 , n48459 );
not ( n48461 , n43757 );
and ( n48462 , n48460 , n48461 );
not ( n226224 , n48460 );
and ( n226225 , n226224 , n43757 );
nor ( n48465 , n48462 , n226225 );
buf ( n48466 , n48465 );
not ( n48467 , n48466 );
and ( n48468 , n226215 , n48467 );
not ( n48469 , n48451 );
nand ( n48470 , n48469 , n47620 );
and ( n226232 , n48470 , n48466 );
nor ( n226233 , n48468 , n226232 );
xor ( n48473 , n48441 , n226233 );
not ( n226235 , n48473 );
not ( n226236 , n41730 );
not ( n48476 , n35275 );
or ( n226238 , n226236 , n48476 );
or ( n226239 , n35275 , n41730 );
nand ( n48479 , n226238 , n226239 );
and ( n48480 , n48479 , n215580 );
not ( n48481 , n48479 );
and ( n48482 , n48481 , n37820 );
nor ( n48483 , n48480 , n48482 );
not ( n48484 , n48483 );
not ( n226246 , n32988 );
not ( n226247 , n26344 );
and ( n48487 , n226246 , n226247 );
and ( n48488 , n32988 , n26344 );
nor ( n48489 , n48487 , n48488 );
not ( n48490 , n48489 );
not ( n48491 , n45696 );
and ( n48492 , n48490 , n48491 );
and ( n226254 , n48489 , n45696 );
nor ( n226255 , n48492 , n226254 );
nand ( n48495 , n226255 , n47750 );
not ( n48496 , n48495 );
or ( n48497 , n48484 , n48496 );
or ( n226259 , n48495 , n48483 );
nand ( n226260 , n48497 , n226259 );
not ( n226261 , n226260 );
not ( n226262 , n33111 );
not ( n48502 , n37882 );
or ( n48503 , n226262 , n48502 );
not ( n48504 , n33111 );
nand ( n48505 , n48504 , n39019 );
nand ( n48506 , n48503 , n48505 );
and ( n48507 , n48506 , n40619 );
not ( n226269 , n48506 );
and ( n226270 , n226269 , n40620 );
nor ( n48510 , n48507 , n226270 );
nand ( n48511 , n48510 , n47641 );
not ( n48512 , n48511 );
not ( n48513 , n28952 );
not ( n226275 , n30321 );
or ( n226276 , n48513 , n226275 );
or ( n48516 , n30321 , n28952 );
nand ( n226278 , n226276 , n48516 );
not ( n226279 , n204436 );
and ( n48519 , n226278 , n226279 );
not ( n48520 , n226278 );
not ( n48521 , n226279 );
and ( n48522 , n48520 , n48521 );
nor ( n226284 , n48519 , n48522 );
not ( n226285 , n226284 );
and ( n48525 , n48512 , n226285 );
and ( n48526 , n48511 , n226284 );
nor ( n48527 , n48525 , n48526 );
not ( n48528 , n48527 );
or ( n48529 , n226261 , n48528 );
or ( n48530 , n48527 , n226260 );
nand ( n226292 , n48529 , n48530 );
xor ( n226293 , n222471 , n223711 );
xnor ( n48533 , n226293 , n40976 );
not ( n48534 , n48533 );
nand ( n48535 , n47566 , n48534 );
and ( n48536 , n37596 , n31126 );
not ( n48537 , n37596 );
and ( n48538 , n48537 , n35481 );
nor ( n226300 , n48536 , n48538 );
and ( n226301 , n226300 , n29694 );
not ( n48541 , n226300 );
and ( n226303 , n48541 , n31137 );
nor ( n226304 , n226301 , n226303 );
not ( n48544 , n226304 );
and ( n48545 , n48535 , n48544 );
not ( n48546 , n48535 );
and ( n48547 , n48546 , n226304 );
nor ( n48548 , n48545 , n48547 );
and ( n48549 , n226292 , n48548 );
not ( n48550 , n226292 );
not ( n48551 , n48548 );
and ( n226313 , n48550 , n48551 );
nor ( n226314 , n48549 , n226313 );
not ( n48554 , n226314 );
and ( n48555 , n226235 , n48554 );
and ( n48556 , n48473 , n226314 );
nor ( n48557 , n48555 , n48556 );
buf ( n226319 , n48557 );
not ( n226320 , n226319 );
and ( n226321 , n48418 , n226320 );
not ( n226322 , n48418 );
and ( n48562 , n226322 , n226319 );
nor ( n48563 , n226321 , n48562 );
not ( n48564 , n48563 );
nand ( n48565 , n48564 , n223839 );
not ( n226327 , n48006 );
not ( n226328 , n225581 );
nand ( n48568 , n226328 , n47852 );
not ( n48569 , n41831 );
not ( n48570 , n28906 );
or ( n48571 , n48569 , n48570 );
not ( n226333 , n41831 );
nand ( n226334 , n226333 , n28907 );
nand ( n48574 , n48571 , n226334 );
and ( n48575 , n48574 , n30943 );
not ( n48576 , n48574 );
and ( n48577 , n48576 , n36890 );
nor ( n226339 , n48575 , n48577 );
and ( n226340 , n48568 , n226339 );
not ( n48580 , n48568 );
not ( n48581 , n226339 );
and ( n48582 , n48580 , n48581 );
nor ( n48583 , n226340 , n48582 );
not ( n48584 , n48583 );
not ( n48585 , n225644 );
nand ( n48586 , n48585 , n47894 );
not ( n48587 , n34702 );
not ( n226349 , n204858 );
not ( n226350 , n226349 );
or ( n48590 , n48587 , n226350 );
or ( n48591 , n226349 , n34702 );
nand ( n48592 , n48590 , n48591 );
not ( n48593 , n204891 );
and ( n48594 , n48592 , n48593 );
not ( n48595 , n48592 );
and ( n226357 , n48595 , n204891 );
nor ( n226358 , n48594 , n226357 );
not ( n48598 , n226358 );
and ( n226360 , n48586 , n48598 );
not ( n226361 , n48586 );
and ( n48601 , n226361 , n226358 );
nor ( n226363 , n226360 , n48601 );
not ( n226364 , n226363 );
or ( n48604 , n48584 , n226364 );
or ( n48605 , n226363 , n48583 );
nand ( n48606 , n48604 , n48605 );
not ( n48607 , n225717 );
not ( n226369 , n47982 );
nand ( n226370 , n48607 , n226369 );
not ( n48610 , n226370 );
not ( n48611 , n28213 );
not ( n48612 , n36237 );
or ( n48613 , n48611 , n48612 );
not ( n48614 , n28213 );
nand ( n48615 , n48614 , n36242 );
nand ( n226377 , n48613 , n48615 );
and ( n226378 , n226377 , n48058 );
not ( n48618 , n226377 );
and ( n48619 , n48618 , n48061 );
nor ( n48620 , n226378 , n48619 );
not ( n48621 , n48620 );
not ( n226383 , n48621 );
and ( n226384 , n48610 , n226383 );
and ( n48624 , n226370 , n48621 );
nor ( n226386 , n226384 , n48624 );
and ( n48626 , n48606 , n226386 );
not ( n48627 , n48606 );
not ( n48628 , n226386 );
and ( n48629 , n48627 , n48628 );
nor ( n48630 , n48626 , n48629 );
not ( n48631 , n48630 );
not ( n48632 , n47943 );
not ( n48633 , n225688 );
nand ( n48634 , n48632 , n48633 );
not ( n48635 , n34976 );
not ( n226397 , n31926 );
not ( n226398 , n226397 );
or ( n48638 , n48635 , n226398 );
or ( n48639 , n42174 , n34976 );
nand ( n48640 , n48638 , n48639 );
not ( n48641 , n48640 );
not ( n48642 , n25550 );
and ( n48643 , n48641 , n48642 );
and ( n48644 , n48640 , n31932 );
nor ( n48645 , n48643 , n48644 );
not ( n226407 , n48645 );
and ( n226408 , n48634 , n226407 );
not ( n48648 , n48634 );
and ( n48649 , n48648 , n48645 );
nor ( n226411 , n226408 , n48649 );
not ( n48651 , n226411 );
not ( n48652 , n48651 );
nand ( n48653 , n47804 , n225763 );
not ( n48654 , n43611 );
not ( n226416 , n36071 );
or ( n226417 , n48654 , n226416 );
or ( n48657 , n37746 , n43611 );
nand ( n48658 , n226417 , n48657 );
and ( n48659 , n48658 , n46349 );
not ( n48660 , n48658 );
and ( n48661 , n48660 , n46348 );
nor ( n48662 , n48659 , n48661 );
not ( n226424 , n48662 );
and ( n226425 , n48653 , n226424 );
not ( n48665 , n48653 );
and ( n48666 , n48665 , n48662 );
nor ( n48667 , n226425 , n48666 );
not ( n48668 , n48667 );
not ( n226430 , n48668 );
or ( n226431 , n48652 , n226430 );
nand ( n48671 , n48667 , n226411 );
nand ( n226433 , n226431 , n48671 );
not ( n226434 , n226433 );
and ( n48674 , n48631 , n226434 );
and ( n48675 , n48630 , n226433 );
nor ( n48676 , n48674 , n48675 );
not ( n48677 , n48676 );
or ( n226439 , n226327 , n48677 );
not ( n226440 , n48006 );
not ( n48680 , n226433 );
not ( n226442 , n48680 );
not ( n226443 , n48630 );
not ( n48683 , n226443 );
or ( n48684 , n226442 , n48683 );
nand ( n48685 , n48630 , n226433 );
nand ( n48686 , n48684 , n48685 );
nand ( n48687 , n226440 , n48686 );
nand ( n48688 , n226439 , n48687 );
not ( n48689 , n48172 );
nand ( n48690 , n48190 , n48689 );
buf ( n48691 , n35693 );
not ( n48692 , n48691 );
not ( n226454 , n48692 );
not ( n226455 , n46668 );
or ( n48695 , n226454 , n226455 );
nand ( n48696 , n46671 , n48691 );
nand ( n48697 , n48695 , n48696 );
not ( n48698 , n44974 );
and ( n226460 , n48697 , n48698 );
not ( n226461 , n48697 );
and ( n48701 , n226461 , n44974 );
nor ( n226463 , n226460 , n48701 );
not ( n226464 , n226463 );
and ( n48704 , n48690 , n226464 );
not ( n226466 , n48690 );
and ( n226467 , n226466 , n226463 );
nor ( n48707 , n48704 , n226467 );
not ( n48708 , n48707 );
not ( n48709 , n48708 );
nand ( n48710 , n48200 , n48207 );
not ( n226472 , n48710 );
not ( n226473 , n204471 );
not ( n48713 , n204468 );
and ( n226475 , n226473 , n48713 );
and ( n226476 , n204471 , n204468 );
nor ( n48716 , n226475 , n226476 );
xor ( n48717 , n48716 , n47216 );
xnor ( n48718 , n48717 , n27968 );
not ( n48719 , n48718 );
not ( n48720 , n48719 );
and ( n48721 , n226472 , n48720 );
and ( n226483 , n48710 , n48719 );
nor ( n226484 , n48721 , n226483 );
not ( n48724 , n226484 );
not ( n48725 , n48724 );
or ( n48726 , n48709 , n48725 );
nand ( n48727 , n226484 , n48707 );
nand ( n226489 , n48726 , n48727 );
not ( n226490 , n226489 );
not ( n48730 , n36624 );
not ( n48731 , n48730 );
not ( n48732 , n38823 );
not ( n48733 , n48732 );
or ( n48734 , n48731 , n48733 );
not ( n48735 , n48730 );
nand ( n48736 , n48735 , n38823 );
nand ( n48737 , n48734 , n48736 );
and ( n48738 , n48737 , n46915 );
not ( n48739 , n48737 );
and ( n226501 , n48739 , n35704 );
nor ( n226502 , n48738 , n226501 );
not ( n48742 , n226502 );
not ( n48743 , n225796 );
nand ( n48744 , n48743 , n48063 );
not ( n48745 , n48744 );
and ( n48746 , n48742 , n48745 );
and ( n48747 , n48744 , n226502 );
nor ( n48748 , n48746 , n48747 );
not ( n48749 , n48748 );
not ( n48750 , n48749 );
not ( n226512 , n48092 );
nand ( n226513 , n225869 , n226512 );
not ( n48753 , n226513 );
buf ( n48754 , n206832 );
xor ( n48755 , n48754 , n28004 );
and ( n48756 , n48755 , n32915 );
not ( n48757 , n48755 );
and ( n48758 , n48757 , n32916 );
nor ( n48759 , n48756 , n48758 );
not ( n226521 , n48759 );
or ( n226522 , n48753 , n226521 );
or ( n48762 , n48759 , n226513 );
nand ( n226524 , n226522 , n48762 );
not ( n226525 , n226524 );
not ( n48765 , n226525 );
or ( n226527 , n48750 , n48765 );
nand ( n226528 , n226524 , n48748 );
nand ( n48768 , n226527 , n226528 );
not ( n48769 , n48137 );
not ( n48770 , n48150 );
nand ( n48771 , n48769 , n48770 );
not ( n48772 , n48771 );
not ( n48773 , n32440 );
not ( n226535 , n225165 );
or ( n226536 , n48773 , n226535 );
not ( n48776 , n32440 );
nand ( n48777 , n48776 , n33524 );
nand ( n48778 , n226536 , n48777 );
not ( n48779 , n33563 );
not ( n48780 , n48779 );
not ( n48781 , n48780 );
xor ( n226543 , n48778 , n48781 );
not ( n226544 , n226543 );
not ( n48784 , n226544 );
and ( n48785 , n48772 , n48784 );
and ( n48786 , n48771 , n226544 );
nor ( n48787 , n48785 , n48786 );
and ( n48788 , n48768 , n48787 );
not ( n226550 , n48768 );
not ( n226551 , n48787 );
and ( n48791 , n226550 , n226551 );
nor ( n48792 , n48788 , n48791 );
not ( n48793 , n48792 );
and ( n48794 , n226490 , n48793 );
and ( n226556 , n226489 , n48792 );
nor ( n226557 , n48794 , n226556 );
buf ( n48797 , n226557 );
and ( n48798 , n48688 , n48797 );
not ( n48799 , n48688 );
not ( n48800 , n48792 );
and ( n48801 , n226489 , n48800 );
not ( n48802 , n226489 );
and ( n48803 , n48802 , n48792 );
nor ( n48804 , n48801 , n48803 );
not ( n48805 , n48804 );
not ( n48806 , n48805 );
and ( n226568 , n48799 , n48806 );
nor ( n226569 , n48798 , n226568 );
not ( n48809 , n226569 );
not ( n48810 , n44288 );
nand ( n48811 , n38093 , n38143 );
not ( n48812 , n48811 );
or ( n226574 , n48810 , n48812 );
nand ( n226575 , n38143 , n38093 );
or ( n48815 , n226575 , n44288 );
nand ( n48816 , n226574 , n48815 );
not ( n48817 , n48816 );
not ( n48818 , n44216 );
not ( n48819 , n48818 );
nand ( n48820 , n44226 , n37947 );
not ( n226582 , n48820 );
or ( n226583 , n48819 , n226582 );
or ( n48823 , n48820 , n48818 );
nand ( n226585 , n226583 , n48823 );
not ( n226586 , n226585 );
not ( n48826 , n44200 );
nand ( n48827 , n48826 , n37825 );
not ( n48828 , n48827 );
not ( n48829 , n44191 );
not ( n48830 , n48829 );
and ( n48831 , n48828 , n48830 );
not ( n48832 , n44200 );
nand ( n48833 , n48832 , n37825 );
and ( n226595 , n48833 , n48829 );
nor ( n226596 , n48831 , n226595 );
not ( n48836 , n226596 );
and ( n48837 , n226586 , n48836 );
and ( n48838 , n226585 , n226596 );
nor ( n48839 , n48837 , n48838 );
not ( n48840 , n48839 );
nand ( n48841 , n222002 , n38005 );
and ( n226603 , n48841 , n44243 );
not ( n226604 , n48841 );
and ( n48844 , n226604 , n37782 );
nor ( n226606 , n226603 , n48844 );
not ( n226607 , n226606 );
and ( n48847 , n48840 , n226607 );
and ( n226609 , n48839 , n226606 );
nor ( n226610 , n48847 , n226609 );
not ( n48850 , n226610 );
not ( n226612 , n48850 );
nand ( n226613 , n38025 , n44278 );
not ( n48853 , n226613 );
not ( n226615 , n44267 );
not ( n226616 , n226615 );
and ( n48856 , n48853 , n226616 );
and ( n226618 , n226613 , n226615 );
nor ( n226619 , n48856 , n226618 );
not ( n48859 , n226619 );
not ( n48860 , n44288 );
nand ( n48861 , n48860 , n38092 );
and ( n48862 , n48861 , n222060 );
not ( n226624 , n48861 );
and ( n226625 , n226624 , n44298 );
nor ( n48865 , n48862 , n226625 );
not ( n48866 , n48865 );
or ( n48867 , n48859 , n48866 );
or ( n48868 , n48865 , n226619 );
nand ( n48869 , n48867 , n48868 );
not ( n48870 , n48869 );
not ( n226632 , n48870 );
and ( n226633 , n226612 , n226632 );
not ( n48873 , n226610 );
and ( n48874 , n48873 , n48870 );
nor ( n48875 , n226633 , n48874 );
not ( n48876 , n48875 );
or ( n48877 , n48817 , n48876 );
not ( n48878 , n48816 );
not ( n226640 , n48869 );
not ( n226641 , n226610 );
or ( n48881 , n226640 , n226641 );
nand ( n48882 , n48850 , n48870 );
nand ( n48883 , n48881 , n48882 );
nand ( n48884 , n48878 , n48883 );
nand ( n48885 , n48877 , n48884 );
not ( n48886 , n38378 );
not ( n226648 , n38128 );
not ( n226649 , n39417 );
or ( n48889 , n226648 , n226649 );
not ( n48890 , n38128 );
nand ( n48891 , n48890 , n32688 );
nand ( n48892 , n48889 , n48891 );
and ( n48893 , n48892 , n47938 );
not ( n48894 , n48892 );
and ( n48895 , n48894 , n47939 );
nor ( n48896 , n48893 , n48895 );
not ( n48897 , n48896 );
nand ( n226659 , n48886 , n48897 );
not ( n226660 , n226659 );
not ( n48900 , n31673 );
not ( n48901 , n46879 );
not ( n48902 , n31828 );
not ( n48903 , n48902 );
or ( n48904 , n48901 , n48903 );
not ( n48905 , n31828 );
or ( n226667 , n48905 , n46879 );
nand ( n226668 , n48904 , n226667 );
not ( n48908 , n226668 );
or ( n48909 , n48900 , n48908 );
or ( n48910 , n226668 , n38709 );
nand ( n48911 , n48909 , n48910 );
not ( n48912 , n48911 );
and ( n48913 , n226660 , n48912 );
not ( n48914 , n48911 );
not ( n48915 , n48914 );
and ( n48916 , n226659 , n48915 );
nor ( n48917 , n48913 , n48916 );
not ( n48918 , n48917 );
buf ( n226680 , n43622 );
not ( n226681 , n226680 );
not ( n48921 , n36071 );
or ( n48922 , n226681 , n48921 );
or ( n48923 , n36074 , n226680 );
nand ( n48924 , n48922 , n48923 );
and ( n226686 , n48924 , n33096 );
not ( n226687 , n48924 );
and ( n48927 , n226687 , n33099 );
nor ( n226689 , n226686 , n48927 );
not ( n226690 , n226689 );
not ( n48930 , n226690 );
buf ( n48931 , n28287 );
not ( n48932 , n48931 );
not ( n48933 , n45214 );
or ( n48934 , n48932 , n48933 );
or ( n48935 , n45214 , n48931 );
nand ( n48936 , n48934 , n48935 );
and ( n48937 , n48936 , n34416 );
not ( n48938 , n48936 );
and ( n48939 , n48938 , n204586 );
nor ( n226701 , n48937 , n48939 );
not ( n226702 , n226701 );
nand ( n48942 , n226702 , n38299 );
not ( n48943 , n48942 );
or ( n48944 , n48930 , n48943 );
or ( n48945 , n48942 , n226690 );
nand ( n226707 , n48944 , n48945 );
not ( n226708 , n226707 );
not ( n48948 , n226708 );
buf ( n48949 , n36801 );
not ( n48950 , n48949 );
not ( n48951 , n45415 );
or ( n48952 , n48950 , n48951 );
or ( n48953 , n42624 , n48949 );
nand ( n48954 , n48952 , n48953 );
and ( n48955 , n48954 , n45817 );
not ( n48956 , n48954 );
and ( n48957 , n48956 , n45418 );
nor ( n226719 , n48955 , n48957 );
nand ( n226720 , n38479 , n226719 );
not ( n48960 , n47606 );
and ( n48961 , n34154 , n48960 );
not ( n48962 , n34154 );
and ( n48963 , n48962 , n47606 );
nor ( n48964 , n48961 , n48963 );
not ( n48965 , n48964 );
and ( n48966 , n204860 , n48965 );
not ( n48967 , n204860 );
and ( n226729 , n48967 , n48964 );
nor ( n226730 , n48966 , n226729 );
not ( n48970 , n226730 );
and ( n48971 , n226720 , n48970 );
not ( n48972 , n226720 );
and ( n48973 , n48972 , n226730 );
nor ( n48974 , n48971 , n48973 );
not ( n48975 , n48974 );
not ( n48976 , n48975 );
or ( n48977 , n48948 , n48976 );
nand ( n48978 , n48974 , n226707 );
nand ( n48979 , n48977 , n48978 );
not ( n226741 , n48979 );
or ( n226742 , n48918 , n226741 );
or ( n48982 , n48979 , n48917 );
nand ( n48983 , n226742 , n48982 );
not ( n48984 , n37996 );
buf ( n48985 , n40120 );
not ( n48986 , n48985 );
and ( n48987 , n48984 , n48986 );
and ( n48988 , n37996 , n48985 );
nor ( n226750 , n48987 , n48988 );
and ( n226751 , n226750 , n35481 );
not ( n48991 , n226750 );
and ( n48992 , n48991 , n38001 );
nor ( n48993 , n226751 , n48992 );
not ( n48994 , n48993 );
nand ( n226756 , n38573 , n48994 );
not ( n226757 , n226756 );
xor ( n48997 , n30012 , n35926 );
xnor ( n48998 , n48997 , n40480 );
not ( n48999 , n48998 );
or ( n49000 , n226757 , n48999 );
or ( n226762 , n48998 , n226756 );
nand ( n226763 , n49000 , n226762 );
not ( n49003 , n226763 );
not ( n226765 , n36309 );
buf ( n226766 , n29987 );
xor ( n49006 , n226766 , n29984 );
not ( n226768 , n49006 );
not ( n226769 , n204791 );
or ( n49009 , n226768 , n226769 );
or ( n226771 , n204791 , n49006 );
nand ( n226772 , n49009 , n226771 );
not ( n49012 , n226772 );
or ( n49013 , n226765 , n49012 );
or ( n49014 , n226772 , n36309 );
nand ( n49015 , n49013 , n49014 );
not ( n226777 , n49015 );
nand ( n226778 , n38588 , n226777 );
not ( n49018 , n226778 );
not ( n49019 , n34276 );
not ( n49020 , n25597 );
or ( n49021 , n49019 , n49020 );
or ( n49022 , n25597 , n34276 );
nand ( n49023 , n49021 , n49022 );
and ( n226785 , n49023 , n29773 );
not ( n226786 , n49023 );
not ( n49026 , n32483 );
and ( n49027 , n226786 , n49026 );
or ( n49028 , n226785 , n49027 );
not ( n49029 , n49028 );
not ( n49030 , n49029 );
and ( n49031 , n49018 , n49030 );
and ( n226793 , n226778 , n49029 );
nor ( n226794 , n49031 , n226793 );
not ( n49034 , n226794 );
or ( n49035 , n49003 , n49034 );
or ( n49036 , n226794 , n226763 );
nand ( n49037 , n49035 , n49036 );
not ( n49038 , n49037 );
and ( n49039 , n48983 , n49038 );
not ( n226801 , n48983 );
and ( n226802 , n226801 , n49037 );
nor ( n49042 , n49039 , n226802 );
buf ( n49043 , n49042 );
and ( n49044 , n48885 , n49043 );
not ( n49045 , n48885 );
not ( n226807 , n49043 );
and ( n226808 , n49045 , n226807 );
nor ( n49048 , n49044 , n226808 );
nand ( n226810 , n48809 , n49048 );
or ( n226811 , n48565 , n226810 );
buf ( n49051 , n37724 );
nor ( n49052 , n48564 , n49051 );
nand ( n49053 , n49052 , n226810 );
buf ( n49054 , n35431 );
nand ( n49055 , n49054 , n31692 );
nand ( n49056 , n226811 , n49053 , n49055 );
buf ( n226818 , n49056 );
buf ( n226819 , n25328 );
not ( n49059 , RI19aa29c8_2548);
or ( n226821 , n226819 , n49059 );
buf ( n226822 , n25335 );
not ( n49062 , RI19acf680_2215);
or ( n49063 , n226822 , n49062 );
nand ( n49064 , n226821 , n49063 );
buf ( n49065 , n49064 );
not ( n49066 , n216226 );
nand ( n49067 , n49066 , n48970 );
not ( n49068 , n49067 );
not ( n49069 , n38400 );
and ( n49070 , n49068 , n49069 );
not ( n49071 , n226730 );
nand ( n49072 , n49071 , n49066 );
and ( n226834 , n49072 , n38400 );
nor ( n226835 , n49070 , n226834 );
not ( n49075 , n226835 );
not ( n49076 , n49075 );
not ( n49077 , n38633 );
or ( n49078 , n49076 , n49077 );
not ( n49079 , n49075 );
nand ( n49080 , n49079 , n38625 );
nand ( n49081 , n49078 , n49080 );
not ( n49082 , n36348 );
buf ( n49083 , n28379 );
not ( n226845 , n49083 );
and ( n226846 , n49082 , n226845 );
and ( n49086 , n225836 , n49083 );
nor ( n226848 , n226846 , n49086 );
xor ( n226849 , n205846 , n226848 );
not ( n49089 , n226849 );
not ( n226851 , n45422 );
nand ( n226852 , n49089 , n226851 );
not ( n49092 , n226852 );
not ( n49093 , n45408 );
not ( n49094 , n49093 );
and ( n49095 , n49092 , n49094 );
and ( n49096 , n226852 , n49093 );
nor ( n49097 , n49095 , n49096 );
not ( n226859 , n49097 );
buf ( n226860 , n37995 );
not ( n49100 , n226860 );
not ( n49101 , n220558 );
or ( n49102 , n49100 , n49101 );
or ( n49103 , n220558 , n226860 );
nand ( n226865 , n49102 , n49103 );
and ( n226866 , n226865 , n34179 );
not ( n49106 , n226865 );
and ( n226868 , n49106 , n42802 );
nor ( n226869 , n226866 , n226868 );
not ( n49109 , n226869 );
not ( n226871 , n45456 );
nand ( n226872 , n49109 , n226871 );
and ( n49112 , n226872 , n45447 );
not ( n226874 , n226872 );
and ( n226875 , n226874 , n45446 );
nor ( n49115 , n49112 , n226875 );
not ( n226877 , n49115 );
or ( n226878 , n226859 , n226877 );
or ( n49118 , n49115 , n49097 );
nand ( n49119 , n226878 , n49118 );
and ( n49120 , n49119 , n223089 );
not ( n49121 , n49119 );
and ( n49122 , n49121 , n45329 );
nor ( n49123 , n49120 , n49122 );
not ( n226885 , n49123 );
not ( n226886 , n226885 );
not ( n49126 , n226886 );
buf ( n49127 , n34167 );
not ( n49128 , n49127 );
not ( n49129 , n49128 );
not ( n226891 , n47607 );
or ( n226892 , n49129 , n226891 );
buf ( n49132 , n47606 );
nand ( n49133 , n49132 , n49127 );
nand ( n49134 , n226892 , n49133 );
and ( n49135 , n49134 , n204860 );
not ( n49136 , n49134 );
not ( n49137 , n226349 );
and ( n226899 , n49136 , n49137 );
nor ( n226900 , n49135 , n226899 );
not ( n49140 , n226900 );
nand ( n226902 , n49140 , n45374 );
not ( n226903 , n226902 );
not ( n49143 , n45369 );
not ( n49144 , n49143 );
and ( n49145 , n226903 , n49144 );
and ( n49146 , n226902 , n49143 );
nor ( n49147 , n49145 , n49146 );
not ( n49148 , n49147 );
not ( n49149 , n223110 );
not ( n49150 , n49149 );
not ( n49151 , n45340 );
buf ( n49152 , n31034 );
buf ( n226914 , RI1749f2b8_960);
and ( n226915 , n49152 , n226914 );
not ( n49155 , n49152 );
and ( n49156 , n49155 , n208792 );
nor ( n226918 , n226915 , n49156 );
not ( n226919 , n226918 );
not ( n49159 , n226919 );
not ( n49160 , n34115 );
or ( n49161 , n49159 , n49160 );
nand ( n49162 , n223793 , n226918 );
nand ( n49163 , n49161 , n49162 );
and ( n226925 , n49163 , n46035 );
not ( n226926 , n49163 );
and ( n226927 , n226926 , n46038 );
nor ( n226928 , n226925 , n226927 );
nand ( n49168 , n49151 , n226928 );
not ( n49169 , n49168 );
or ( n49170 , n49150 , n49169 );
or ( n49171 , n49168 , n49149 );
nand ( n226933 , n49170 , n49171 );
not ( n226934 , n226933 );
and ( n49174 , n49148 , n226934 );
and ( n226936 , n49147 , n226933 );
nor ( n226937 , n49174 , n226936 );
not ( n49177 , n226937 );
not ( n49178 , n49177 );
and ( n49179 , n49126 , n49178 );
and ( n49180 , n226886 , n49177 );
nor ( n49181 , n49179 , n49180 );
buf ( n49182 , n49181 );
and ( n49183 , n49081 , n49182 );
not ( n49184 , n49081 );
not ( n49185 , n226937 );
not ( n226947 , n49185 );
not ( n226948 , n49123 );
or ( n49188 , n226947 , n226948 );
nand ( n49189 , n226885 , n226937 );
nand ( n49190 , n49188 , n49189 );
buf ( n49191 , n49190 );
and ( n49192 , n49184 , n49191 );
nor ( n49193 , n49183 , n49192 );
buf ( n226955 , n33252 );
nor ( n226956 , n49193 , n226955 );
not ( n49196 , n32219 );
not ( n226958 , n39615 );
not ( n226959 , n206591 );
or ( n49199 , n226958 , n226959 );
or ( n49200 , n206591 , n39615 );
nand ( n49201 , n49199 , n49200 );
not ( n49202 , n49201 );
and ( n49203 , n49196 , n49202 );
and ( n49204 , n32219 , n49201 );
nor ( n226966 , n49203 , n49204 );
not ( n226967 , n32625 );
not ( n49207 , n45280 );
or ( n49208 , n226967 , n49207 );
nand ( n49209 , n44157 , n32621 );
nand ( n49210 , n49208 , n49209 );
and ( n49211 , n49210 , n45314 );
not ( n49212 , n49210 );
and ( n226974 , n49212 , n45310 );
or ( n226975 , n49211 , n226974 );
nand ( n49215 , n226966 , n226975 );
not ( n49216 , n49215 );
xor ( n49217 , n26259 , n43122 );
xnor ( n49218 , n49217 , n45672 );
not ( n49219 , n49218 );
and ( n49220 , n49216 , n49219 );
and ( n226982 , n49215 , n49218 );
nor ( n226983 , n49220 , n226982 );
not ( n49223 , n226983 );
not ( n226985 , n49223 );
buf ( n226986 , n31965 );
not ( n49226 , n226986 );
not ( n49227 , n31962 );
and ( n49228 , n49226 , n49227 );
and ( n49229 , n226986 , n31962 );
nor ( n226991 , n49228 , n49229 );
xor ( n226992 , n226991 , n31227 );
xnor ( n49232 , n226992 , n29088 );
buf ( n49233 , n49232 );
not ( n49234 , n49233 );
not ( n49235 , n49218 );
not ( n49236 , n226966 );
nand ( n49237 , n49235 , n49236 );
not ( n49238 , n49237 );
or ( n49239 , n49234 , n49238 );
or ( n227001 , n49237 , n49233 );
nand ( n227002 , n49239 , n227001 );
not ( n49242 , n227002 );
xor ( n227004 , n30403 , n48174 );
xnor ( n227005 , n227004 , n33002 );
not ( n49245 , n227005 );
xor ( n227007 , n25836 , n37580 );
xnor ( n227008 , n227007 , n38839 );
not ( n49248 , n227008 );
nand ( n49249 , n49245 , n49248 );
not ( n227011 , n49249 );
buf ( n227012 , n28645 );
not ( n49252 , n227012 );
not ( n49253 , n208303 );
or ( n49254 , n49252 , n49253 );
or ( n49255 , n208303 , n227012 );
nand ( n49256 , n49254 , n49255 );
buf ( n227018 , n33759 );
and ( n227019 , n49256 , n227018 );
not ( n49259 , n49256 );
and ( n49260 , n49259 , n33760 );
nor ( n49261 , n227019 , n49260 );
not ( n49262 , n49261 );
and ( n227024 , n227011 , n49262 );
and ( n227025 , n49249 , n49261 );
nor ( n49265 , n227024 , n227025 );
not ( n49266 , n49265 );
or ( n49267 , n49242 , n49266 );
not ( n49268 , n227002 );
not ( n227030 , n49265 );
nand ( n227031 , n49268 , n227030 );
nand ( n49271 , n49267 , n227031 );
not ( n49272 , n29813 );
not ( n49273 , n35584 );
or ( n49274 , n49272 , n49273 );
not ( n49275 , n29813 );
nand ( n49276 , n49275 , n35590 );
nand ( n227038 , n49274 , n49276 );
not ( n227039 , n227038 );
not ( n49279 , n35940 );
and ( n49280 , n227039 , n49279 );
and ( n49281 , n41878 , n227038 );
nor ( n49282 , n49280 , n49281 );
not ( n227044 , n218656 );
nor ( n227045 , n43672 , n206656 );
not ( n49285 , n227045 );
nand ( n49286 , n43672 , n206656 );
nand ( n49287 , n49285 , n49286 );
not ( n227049 , n49287 );
or ( n227050 , n227044 , n227049 );
or ( n49290 , n49287 , n218656 );
nand ( n49291 , n227050 , n49290 );
nand ( n49292 , n49282 , n49291 );
not ( n49293 , n38254 );
not ( n49294 , n29607 );
or ( n49295 , n49293 , n49294 );
not ( n49296 , n38254 );
nand ( n49297 , n49296 , n30781 );
nand ( n49298 , n49295 , n49297 );
and ( n49299 , n49298 , n207409 );
not ( n227061 , n49298 );
and ( n227062 , n227061 , n29647 );
nor ( n49302 , n49299 , n227062 );
and ( n49303 , n49292 , n49302 );
not ( n49304 , n49292 );
not ( n49305 , n49302 );
and ( n49306 , n49304 , n49305 );
nor ( n49307 , n49303 , n49306 );
not ( n49308 , n49307 );
not ( n227070 , n49308 );
buf ( n227071 , n28329 );
not ( n227072 , n227071 );
not ( n227073 , n48073 );
or ( n49313 , n227072 , n227073 );
or ( n227075 , n36308 , n227071 );
nand ( n227076 , n49313 , n227075 );
and ( n49316 , n227076 , n36349 );
not ( n49317 , n227076 );
not ( n49318 , n36349 );
and ( n49319 , n49317 , n49318 );
nor ( n227081 , n49316 , n49319 );
not ( n227082 , n227081 );
not ( n49322 , n33147 );
not ( n49323 , n28247 );
or ( n49324 , n49322 , n49323 );
or ( n49325 , n28247 , n33147 );
nand ( n227087 , n49324 , n49325 );
not ( n227088 , n227087 );
not ( n49328 , n28288 );
and ( n227090 , n227088 , n49328 );
and ( n227091 , n227087 , n28288 );
nor ( n49331 , n227090 , n227091 );
not ( n49332 , n49331 );
nand ( n49333 , n227082 , n49332 );
not ( n49334 , n49333 );
not ( n227096 , n39972 );
buf ( n227097 , RI17447ce8_1386);
not ( n49337 , n28656 );
xor ( n49338 , n227097 , n49337 );
xnor ( n49339 , n49338 , n28663 );
not ( n49340 , n49339 );
or ( n49341 , n227096 , n49340 );
or ( n49342 , n49339 , n39972 );
nand ( n49343 , n49341 , n49342 );
and ( n49344 , n49343 , n28646 );
not ( n49345 , n49343 );
and ( n49346 , n49345 , n47581 );
nor ( n49347 , n49344 , n49346 );
not ( n49348 , n49347 );
not ( n49349 , n49348 );
and ( n227111 , n49334 , n49349 );
not ( n227112 , n227081 );
nand ( n49352 , n227112 , n49332 );
and ( n49353 , n49352 , n49348 );
nor ( n49354 , n227111 , n49353 );
not ( n49355 , n49354 );
not ( n49356 , n49355 );
or ( n227118 , n227070 , n49356 );
nand ( n227119 , n49354 , n49307 );
nand ( n49359 , n227118 , n227119 );
not ( n49360 , n204876 );
not ( n49361 , n211806 );
or ( n49362 , n49360 , n49361 );
not ( n49363 , n204876 );
nand ( n49364 , n49363 , n34051 );
nand ( n49365 , n49362 , n49364 );
and ( n49366 , n49365 , n34089 );
not ( n49367 , n49365 );
and ( n227129 , n49367 , n34103 );
nor ( n227130 , n49366 , n227129 );
buf ( n49370 , n227130 );
not ( n49371 , n49370 );
not ( n49372 , n27775 );
not ( n227134 , RI1744e930_1353);
xor ( n227135 , n227134 , n31246 );
xor ( n49375 , n227135 , n31252 );
not ( n49376 , n49375 );
not ( n49377 , n49376 );
or ( n49378 , n49372 , n49377 );
or ( n49379 , n49376 , n27775 );
nand ( n49380 , n49378 , n49379 );
and ( n227142 , n49380 , n31264 );
not ( n227143 , n49380 );
and ( n49383 , n227143 , n31273 );
nor ( n227145 , n227142 , n49383 );
not ( n227146 , n227145 );
nand ( n49386 , n49371 , n227146 );
not ( n49387 , n49386 );
not ( n49388 , n219113 );
not ( n49389 , n25963 );
or ( n227151 , n49388 , n49389 );
not ( n227152 , n219113 );
nand ( n49392 , n227152 , n25977 );
nand ( n49393 , n227151 , n49392 );
not ( n49394 , n49393 );
not ( n49395 , n25457 );
and ( n49396 , n49394 , n49395 );
and ( n49397 , n36983 , n49393 );
nor ( n227159 , n49396 , n49397 );
not ( n227160 , n227159 );
not ( n49400 , n227160 );
and ( n227162 , n49387 , n49400 );
and ( n227163 , n49386 , n227160 );
nor ( n49403 , n227162 , n227163 );
and ( n227165 , n49359 , n49403 );
not ( n227166 , n49359 );
not ( n49406 , n49403 );
and ( n49407 , n227166 , n49406 );
nor ( n49408 , n227165 , n49407 );
and ( n49409 , n49271 , n49408 );
not ( n49410 , n49271 );
not ( n49411 , n49408 );
and ( n227173 , n49410 , n49411 );
nor ( n227174 , n49409 , n227173 );
not ( n49414 , n227174 );
or ( n49415 , n226985 , n49414 );
not ( n49416 , n49223 );
and ( n49417 , n49271 , n49411 );
not ( n227179 , n49271 );
and ( n227180 , n227179 , n49408 );
nor ( n49420 , n49417 , n227180 );
nand ( n49421 , n49416 , n49420 );
nand ( n49422 , n49415 , n49421 );
buf ( n49423 , RI173d7b78_1704);
not ( n49424 , n49423 );
not ( n49425 , n33947 );
or ( n49426 , n49424 , n49425 );
or ( n49427 , n33947 , n49423 );
nand ( n49428 , n49426 , n49427 );
and ( n49429 , n49428 , n33957 );
not ( n227191 , n49428 );
and ( n227192 , n227191 , n33954 );
nor ( n49432 , n49429 , n227192 );
not ( n49433 , n35336 );
not ( n49434 , n29607 );
or ( n49435 , n49433 , n49434 );
or ( n227197 , n29607 , n35336 );
nand ( n227198 , n49435 , n227197 );
and ( n49438 , n227198 , n207407 );
not ( n49439 , n227198 );
and ( n49440 , n49439 , n46665 );
nor ( n49441 , n49438 , n49440 );
not ( n227203 , n49441 );
nand ( n227204 , n49432 , n227203 );
not ( n49444 , n227204 );
xor ( n49445 , n29308 , n205420 );
and ( n49446 , n49445 , n205436 );
not ( n49447 , n49445 );
and ( n49448 , n49447 , n205435 );
nor ( n49449 , n49446 , n49448 );
not ( n227211 , n49449 );
not ( n227212 , n227211 );
and ( n49452 , n49444 , n227212 );
and ( n49453 , n227204 , n227211 );
nor ( n49454 , n49452 , n49453 );
not ( n49455 , n49454 );
not ( n49456 , n219841 );
not ( n49457 , n29377 );
not ( n49458 , n40369 );
or ( n49459 , n49457 , n49458 );
or ( n227221 , n40369 , n29377 );
nand ( n227222 , n49459 , n227221 );
not ( n49462 , n227222 );
or ( n49463 , n49456 , n49462 );
not ( n49464 , n227222 );
nand ( n49465 , n49464 , n42159 );
nand ( n49466 , n49463 , n49465 );
not ( n49467 , n49466 );
not ( n227229 , n37867 );
not ( n227230 , n44932 );
or ( n49470 , n227229 , n227230 );
not ( n49471 , n37867 );
nand ( n49472 , n49471 , n45418 );
nand ( n49473 , n49470 , n49472 );
and ( n49474 , n49473 , n222700 );
not ( n49475 , n49473 );
not ( n227237 , n222667 );
and ( n227238 , n49475 , n227237 );
nor ( n49478 , n49474 , n227238 );
not ( n227240 , n49478 );
nand ( n227241 , n49467 , n227240 );
not ( n49481 , n45196 );
xor ( n49482 , n28321 , n28338 );
xor ( n49483 , n49482 , n28329 );
not ( n49484 , n49483 );
or ( n227246 , n49481 , n49484 );
not ( n227247 , n45192 );
or ( n49487 , n49483 , n227247 );
nand ( n227249 , n227246 , n49487 );
and ( n227250 , n227249 , n28382 );
not ( n49490 , n227249 );
not ( n49491 , n39671 );
and ( n49492 , n49490 , n49491 );
nor ( n49493 , n227250 , n49492 );
buf ( n49494 , n49493 );
and ( n49495 , n227241 , n49494 );
not ( n49496 , n227241 );
not ( n49497 , n49494 );
and ( n49498 , n49496 , n49497 );
nor ( n49499 , n49495 , n49498 );
not ( n227261 , n49499 );
or ( n227262 , n49455 , n227261 );
or ( n49502 , n49499 , n49454 );
nand ( n49503 , n227262 , n49502 );
buf ( n49504 , n28251 );
xor ( n49505 , n205036 , n49504 );
xnor ( n49506 , n49505 , n32082 );
not ( n49507 , n208320 );
not ( n227269 , n38764 );
or ( n227270 , n49507 , n227269 );
or ( n49510 , n27802 , n208320 );
nand ( n49511 , n227270 , n49510 );
and ( n49512 , n49511 , n38774 );
not ( n49513 , n49511 );
and ( n49514 , n49513 , n38770 );
nor ( n49515 , n49512 , n49514 );
nand ( n49516 , n49506 , n49515 );
not ( n49517 , n49516 );
not ( n49518 , n38643 );
not ( n49519 , n220435 );
or ( n227281 , n49518 , n49519 );
not ( n227282 , n38643 );
nand ( n49522 , n227282 , n220432 );
nand ( n49523 , n227281 , n49522 );
and ( n49524 , n49523 , n31428 );
not ( n49525 , n49523 );
and ( n49526 , n49525 , n42680 );
nor ( n49527 , n49524 , n49526 );
not ( n49528 , n49527 );
not ( n49529 , n49528 );
and ( n227291 , n49517 , n49529 );
and ( n227292 , n49516 , n49528 );
nor ( n49532 , n227291 , n227292 );
and ( n49533 , n49503 , n49532 );
not ( n49534 , n49503 );
not ( n49535 , n49532 );
and ( n227297 , n49534 , n49535 );
nor ( n227298 , n49533 , n227297 );
not ( n49538 , n227298 );
not ( n227300 , n208419 );
buf ( n227301 , n37864 );
not ( n49541 , n227301 );
or ( n227303 , n227300 , n49541 );
nand ( n227304 , n40620 , n30654 );
nand ( n49544 , n227303 , n227304 );
not ( n227306 , n39922 );
and ( n227307 , n49544 , n227306 );
not ( n49547 , n49544 );
and ( n49548 , n49547 , n39922 );
nor ( n49549 , n227307 , n49548 );
not ( n49550 , n49549 );
not ( n49551 , n32151 );
not ( n49552 , n33614 );
or ( n49553 , n49551 , n49552 );
or ( n49554 , n33614 , n32151 );
nand ( n49555 , n49553 , n49554 );
and ( n49556 , n49555 , n43787 );
not ( n227318 , n49555 );
and ( n227319 , n227318 , n41520 );
nor ( n49559 , n49556 , n227319 );
not ( n49560 , n49559 );
nand ( n49561 , n49550 , n49560 );
not ( n49562 , n49561 );
not ( n49563 , n42494 );
not ( n49564 , n223530 );
or ( n49565 , n49563 , n49564 );
or ( n49566 , n223530 , n42494 );
nand ( n49567 , n49565 , n49566 );
not ( n49568 , n41754 );
buf ( n227330 , n49568 );
and ( n227331 , n49567 , n227330 );
not ( n49571 , n49567 );
and ( n49572 , n49571 , n42356 );
nor ( n49573 , n227331 , n49572 );
not ( n49574 , n49573 );
not ( n49575 , n49574 );
and ( n49576 , n49562 , n49575 );
and ( n49577 , n49561 , n49574 );
nor ( n49578 , n49576 , n49577 );
not ( n49579 , n49578 );
not ( n49580 , n49579 );
not ( n227342 , n37636 );
not ( n227343 , n31136 );
or ( n49583 , n227342 , n227343 );
or ( n49584 , n31136 , n37636 );
nand ( n49585 , n49583 , n49584 );
and ( n49586 , n49585 , n34589 );
not ( n49587 , n49585 );
and ( n49588 , n49587 , n207493 );
nor ( n49589 , n49586 , n49588 );
not ( n49590 , n49589 );
not ( n227352 , n29753 );
not ( n227353 , n46966 );
or ( n49593 , n227352 , n227353 );
or ( n49594 , n222443 , n29753 );
nand ( n49595 , n49593 , n49594 );
and ( n49596 , n49595 , n206591 );
not ( n49597 , n49595 );
and ( n49598 , n49597 , n28817 );
nor ( n227360 , n49596 , n49598 );
nand ( n227361 , n49590 , n227360 );
not ( n49601 , n227361 );
xor ( n49602 , n27897 , n36255 );
xnor ( n49603 , n49602 , n36258 );
not ( n49604 , n49603 );
or ( n49605 , n49601 , n49604 );
or ( n49606 , n49603 , n227361 );
nand ( n227368 , n49605 , n49606 );
not ( n227369 , n227368 );
not ( n49609 , n227369 );
or ( n227371 , n49580 , n49609 );
nand ( n227372 , n227368 , n49578 );
nand ( n49612 , n227371 , n227372 );
not ( n49613 , n49612 );
and ( n227375 , n49538 , n49613 );
not ( n227376 , n49538 );
and ( n49616 , n227376 , n49612 );
nor ( n49617 , n227375 , n49616 );
buf ( n49618 , n49617 );
and ( n49619 , n49422 , n49618 );
not ( n227381 , n49422 );
not ( n227382 , n49613 );
not ( n49622 , n227298 );
not ( n227384 , n49622 );
or ( n227385 , n227382 , n227384 );
nand ( n49625 , n227298 , n49612 );
nand ( n49626 , n227385 , n49625 );
buf ( n49627 , n49626 );
and ( n49628 , n227381 , n49627 );
nor ( n49629 , n49619 , n49628 );
not ( n49630 , n38696 );
buf ( n49631 , n25957 );
not ( n49632 , n49631 );
not ( n227394 , n35622 );
or ( n227395 , n49632 , n227394 );
or ( n49635 , n35622 , n49631 );
nand ( n49636 , n227395 , n49635 );
and ( n49637 , n49636 , n42058 );
not ( n49638 , n49636 );
and ( n49639 , n49638 , n42057 );
nor ( n49640 , n49637 , n49639 );
nand ( n49641 , n38935 , n49640 );
not ( n49642 , n49641 );
or ( n227404 , n49630 , n49642 );
or ( n227405 , n49641 , n38696 );
nand ( n49645 , n227404 , n227405 );
not ( n49646 , n49645 );
buf ( n49647 , n36261 );
not ( n49648 , n49647 );
not ( n227410 , n37537 );
or ( n227411 , n49648 , n227410 );
or ( n49651 , n37537 , n49647 );
nand ( n49652 , n227411 , n49651 );
and ( n49653 , n38037 , n49652 );
not ( n49654 , n38037 );
not ( n227416 , n49652 );
and ( n227417 , n49654 , n227416 );
nor ( n49657 , n49653 , n227417 );
not ( n49658 , n49657 );
not ( n49659 , n32066 );
not ( n49660 , n31176 );
or ( n227422 , n49659 , n49660 );
not ( n227423 , n32066 );
nand ( n49663 , n227423 , n36684 );
nand ( n49664 , n227422 , n49663 );
and ( n49665 , n49664 , n36243 );
not ( n49666 , n49664 );
and ( n49667 , n49666 , n36238 );
nor ( n49668 , n49665 , n49667 );
nand ( n227430 , n49658 , n49668 );
not ( n227431 , n227430 );
not ( n49671 , n38792 );
and ( n49672 , n227431 , n49671 );
and ( n49673 , n227430 , n38792 );
nor ( n49674 , n49672 , n49673 );
not ( n227436 , n49674 );
buf ( n227437 , n33471 );
not ( n49677 , n227437 );
not ( n227439 , n32362 );
not ( n227440 , n227439 );
or ( n49680 , n49677 , n227440 );
or ( n49681 , n227439 , n227437 );
nand ( n49682 , n49680 , n49681 );
not ( n227444 , n37296 );
and ( n227445 , n49682 , n227444 );
not ( n227446 , n49682 );
and ( n227447 , n227446 , n37296 );
nor ( n49687 , n227445 , n227447 );
buf ( n49688 , n33214 );
not ( n49689 , n49688 );
not ( n49690 , n25721 );
or ( n227452 , n49689 , n49690 );
or ( n227453 , n25772 , n49688 );
nand ( n49693 , n227452 , n227453 );
and ( n49694 , n49693 , n44351 );
not ( n49695 , n49693 );
and ( n49696 , n49695 , n44347 );
nor ( n49697 , n49694 , n49696 );
nand ( n49698 , n49687 , n49697 );
not ( n227460 , n38738 );
and ( n227461 , n49698 , n227460 );
not ( n49701 , n49698 );
and ( n49702 , n49701 , n38738 );
nor ( n49703 , n227461 , n49702 );
not ( n49704 , n49703 );
or ( n49705 , n227436 , n49704 );
or ( n49706 , n49674 , n49703 );
nand ( n49707 , n49705 , n49706 );
buf ( n49708 , n41290 );
not ( n49709 , n49708 );
not ( n49710 , n207493 );
or ( n227472 , n49709 , n49710 );
or ( n227473 , n207493 , n49708 );
nand ( n49713 , n227472 , n227473 );
xor ( n49714 , n49713 , n33444 );
buf ( n49715 , n34515 );
and ( n49716 , n49715 , n43635 );
not ( n49717 , n49715 );
xor ( n49718 , n43624 , n43633 );
xnor ( n227480 , n49718 , n37742 );
and ( n227481 , n49717 , n227480 );
nor ( n49721 , n49716 , n227481 );
not ( n227483 , n49721 );
not ( n227484 , n44135 );
or ( n49724 , n227483 , n227484 );
not ( n49725 , n44136 );
or ( n49726 , n49725 , n49721 );
nand ( n49727 , n49724 , n49726 );
buf ( n227489 , n49727 );
nand ( n227490 , n49714 , n227489 );
not ( n49730 , n227490 );
not ( n49731 , n38851 );
and ( n49732 , n49730 , n49731 );
and ( n49733 , n227490 , n38851 );
nor ( n227495 , n49732 , n49733 );
not ( n227496 , n227495 );
and ( n227497 , n49707 , n227496 );
not ( n227498 , n49707 );
and ( n49738 , n227498 , n227495 );
nor ( n49739 , n227497 , n49738 );
not ( n49740 , n34807 );
buf ( n49741 , RI174a0320_955);
not ( n227503 , n49741 );
not ( n227504 , n205093 );
or ( n49744 , n227503 , n227504 );
not ( n227506 , n205093 );
nand ( n227507 , n227506 , n205090 );
nand ( n49747 , n49744 , n227507 );
not ( n49748 , n49747 );
nor ( n49749 , n49748 , n34763 );
not ( n49750 , n49749 );
not ( n49751 , n49747 );
nand ( n49752 , n49751 , n34763 );
nand ( n227514 , n49750 , n49752 );
not ( n227515 , n227514 );
or ( n49755 , n49740 , n227515 );
or ( n49756 , n227514 , n36411 );
nand ( n49757 , n49755 , n49756 );
not ( n49758 , n49757 );
xor ( n227520 , n41016 , n41520 );
buf ( n227521 , n225459 );
xnor ( n49761 , n227520 , n227521 );
not ( n227523 , n49761 );
nand ( n227524 , n49758 , n227523 );
and ( n49764 , n227524 , n39025 );
not ( n49765 , n227524 );
and ( n49766 , n49765 , n39026 );
nor ( n227528 , n49764 , n49766 );
not ( n49768 , n227528 );
not ( n49769 , n49768 );
not ( n49770 , n38696 );
not ( n49771 , n49640 );
nand ( n49772 , n49770 , n49771 );
and ( n49773 , n49772 , n38923 );
not ( n49774 , n49772 );
and ( n49775 , n49774 , n38679 );
nor ( n227537 , n49773 , n49775 );
not ( n227538 , n227537 );
not ( n49778 , n227538 );
or ( n227540 , n49769 , n49778 );
nand ( n227541 , n227537 , n227528 );
nand ( n49781 , n227540 , n227541 );
and ( n49782 , n49739 , n49781 );
not ( n49783 , n49739 );
not ( n49784 , n49781 );
and ( n49785 , n49783 , n49784 );
nor ( n49786 , n49782 , n49785 );
not ( n227548 , n49786 );
not ( n227549 , n227548 );
or ( n49789 , n49646 , n227549 );
not ( n49790 , n49645 );
not ( n49791 , n49739 );
and ( n49792 , n49791 , n49784 );
not ( n49793 , n49791 );
and ( n49794 , n49793 , n49781 );
nor ( n227556 , n49792 , n49794 );
nand ( n227557 , n49790 , n227556 );
nand ( n49797 , n49789 , n227557 );
not ( n227559 , n28008 );
not ( n227560 , n37579 );
or ( n49800 , n227559 , n227560 );
not ( n49801 , n28008 );
nand ( n49802 , n49801 , n37580 );
nand ( n49803 , n49800 , n49802 );
and ( n49804 , n49803 , n204505 );
not ( n49805 , n49803 );
and ( n227567 , n49805 , n204508 );
nor ( n227568 , n49804 , n227567 );
not ( n49808 , n208085 );
not ( n49809 , n29334 );
or ( n49810 , n49808 , n49809 );
or ( n49811 , n29334 , n208085 );
nand ( n227573 , n49810 , n49811 );
and ( n227574 , n227573 , n41149 );
not ( n49814 , n227573 );
and ( n227576 , n49814 , n46753 );
nor ( n227577 , n227574 , n227576 );
nand ( n49817 , n227568 , n227577 );
not ( n49818 , n49817 );
not ( n49819 , n39147 );
not ( n49820 , n49819 );
and ( n49821 , n49818 , n49820 );
and ( n49822 , n49817 , n49819 );
nor ( n49823 , n49821 , n49822 );
not ( n49824 , n28256 );
not ( n227586 , n45218 );
or ( n227587 , n49824 , n227586 );
not ( n49827 , n28256 );
nand ( n227589 , n49827 , n45214 );
nand ( n227590 , n227587 , n227589 );
not ( n49830 , n227590 );
not ( n49831 , n204586 );
and ( n49832 , n49830 , n49831 );
and ( n49833 , n204586 , n227590 );
nor ( n227595 , n49832 , n49833 );
not ( n227596 , n227595 );
not ( n49836 , n33728 );
not ( n227598 , n33203 );
or ( n227599 , n49836 , n227598 );
or ( n49839 , n33203 , n33728 );
nand ( n49840 , n227599 , n49839 );
not ( n49841 , n49840 );
not ( n49842 , n33225 );
or ( n227604 , n49841 , n49842 );
or ( n227605 , n33225 , n49840 );
nand ( n49845 , n227604 , n227605 );
not ( n227607 , n49845 );
not ( n227608 , n33195 );
and ( n49848 , n227607 , n227608 );
and ( n227610 , n49845 , n33195 );
nor ( n227611 , n49848 , n227610 );
nand ( n49851 , n227596 , n227611 );
not ( n49852 , n39180 );
and ( n49853 , n49851 , n49852 );
not ( n49854 , n49851 );
and ( n49855 , n49854 , n39180 );
nor ( n49856 , n49853 , n49855 );
xor ( n227618 , n49823 , n49856 );
not ( n227619 , n227618 );
xor ( n49859 , n39937 , n47581 );
xnor ( n49860 , n49859 , n28665 );
not ( n49861 , n26209 );
not ( n49862 , n48779 );
or ( n227624 , n49861 , n49862 );
or ( n227625 , n26209 , n48779 );
nand ( n49865 , n227624 , n227625 );
and ( n49866 , n49865 , n36620 );
not ( n49867 , n49865 );
and ( n49868 , n49867 , n36626 );
nor ( n49869 , n49866 , n49868 );
not ( n227631 , n49869 );
nand ( n227632 , n49860 , n227631 );
not ( n49872 , n39075 );
and ( n49873 , n227632 , n49872 );
not ( n49874 , n227632 );
and ( n49875 , n49874 , n39075 );
nor ( n49876 , n49873 , n49875 );
not ( n49877 , n49876 );
and ( n227639 , n227619 , n49877 );
and ( n227640 , n227618 , n49876 );
nor ( n49880 , n227639 , n227640 );
not ( n49881 , n39289 );
not ( n49882 , n40285 );
not ( n49883 , n209347 );
not ( n49884 , n206437 );
or ( n49885 , n49883 , n49884 );
not ( n227647 , n209347 );
nand ( n227648 , n227647 , n37229 );
nand ( n49888 , n49885 , n227648 );
not ( n49889 , n49888 );
or ( n49890 , n49882 , n49889 );
or ( n49891 , n205096 , n49888 );
nand ( n49892 , n49890 , n49891 );
not ( n49893 , n49892 );
buf ( n227655 , RI174001e0_1507);
not ( n227656 , n227655 );
not ( n49896 , n43936 );
or ( n49897 , n227656 , n49896 );
or ( n49898 , n43936 , n227655 );
nand ( n49899 , n49897 , n49898 );
and ( n49900 , n49899 , n37455 );
not ( n49901 , n49899 );
and ( n49902 , n49901 , n44458 );
nor ( n49903 , n49900 , n49902 );
nand ( n227665 , n49893 , n49903 );
not ( n227666 , n227665 );
or ( n49906 , n49881 , n227666 );
or ( n49907 , n227665 , n39289 );
nand ( n49908 , n49906 , n49907 );
not ( n49909 , n49908 );
not ( n49910 , n39363 );
not ( n49911 , n35777 );
not ( n227673 , n39480 );
or ( n227674 , n49911 , n227673 );
or ( n49914 , n39481 , n35777 );
nand ( n49915 , n227674 , n49914 );
not ( n49916 , n49915 );
not ( n49917 , n43554 );
and ( n49918 , n49916 , n49917 );
and ( n49919 , n49915 , n43554 );
nor ( n227681 , n49918 , n49919 );
not ( n227682 , n204943 );
buf ( n49922 , n213777 );
not ( n227684 , n49922 );
or ( n227685 , n227682 , n227684 );
not ( n49925 , n204943 );
nand ( n227687 , n49925 , n36025 );
nand ( n227688 , n227685 , n227687 );
and ( n49928 , n227688 , n40862 );
not ( n49929 , n227688 );
and ( n49930 , n49929 , n221434 );
nor ( n49931 , n49928 , n49930 );
nand ( n227693 , n227681 , n49931 );
not ( n227694 , n227693 );
and ( n49934 , n49910 , n227694 );
and ( n49935 , n39363 , n227693 );
nor ( n49936 , n49934 , n49935 );
not ( n227698 , n49936 );
or ( n227699 , n49909 , n227698 );
or ( n49939 , n49936 , n49908 );
nand ( n49940 , n227699 , n49939 );
not ( n49941 , n49940 );
and ( n49942 , n49880 , n49941 );
not ( n49943 , n49880 );
and ( n49944 , n49943 , n49940 );
nor ( n227706 , n49942 , n49944 );
buf ( n227707 , n227706 );
buf ( n49947 , n227707 );
and ( n49948 , n49797 , n49947 );
not ( n49949 , n49797 );
not ( n49950 , n227707 );
and ( n227712 , n49949 , n49950 );
nor ( n227713 , n49948 , n227712 );
not ( n49953 , n227713 );
nand ( n49954 , n226956 , n49629 , n49953 );
not ( n49955 , n49193 );
not ( n49956 , n49955 );
not ( n227718 , n49629 );
or ( n227719 , n49956 , n227718 );
buf ( n49959 , n33253 );
nor ( n49960 , n49953 , n49959 );
nand ( n49961 , n227719 , n49960 );
nand ( n49962 , n35431 , n204839 );
nand ( n49963 , n49954 , n49961 , n49962 );
buf ( n49964 , n49963 );
nand ( n49965 , n221864 , n42815 );
not ( n49966 , n49965 );
not ( n49967 , n42804 );
not ( n49968 , n49967 );
or ( n227730 , n49966 , n49968 );
or ( n227731 , n49967 , n49965 );
nand ( n49971 , n227730 , n227731 );
buf ( n49972 , n49971 );
not ( n49973 , n49972 );
not ( n49974 , n43010 );
or ( n49975 , n49973 , n49974 );
or ( n49976 , n43010 , n49972 );
nand ( n227738 , n49975 , n49976 );
not ( n227739 , n48816 );
not ( n49979 , n38048 );
nand ( n49980 , n38024 , n49979 );
not ( n49981 , n49980 );
not ( n49982 , n44279 );
and ( n227744 , n49981 , n49982 );
and ( n227745 , n49980 , n44279 );
nor ( n49985 , n227744 , n227745 );
not ( n49986 , n49985 );
and ( n49987 , n227739 , n49986 );
and ( n49988 , n48816 , n49985 );
nor ( n227750 , n49987 , n49988 );
not ( n227751 , n227750 );
not ( n49991 , n37799 );
nand ( n49992 , n49991 , n37824 );
not ( n49993 , n49992 );
not ( n49994 , n44200 );
and ( n227756 , n49993 , n49994 );
not ( n227757 , n48832 );
and ( n49997 , n49992 , n227757 );
nor ( n49998 , n227756 , n49997 );
not ( n49999 , n49998 );
not ( n50000 , n37883 );
nand ( n227762 , n50000 , n37948 );
and ( n227763 , n227762 , n44226 );
not ( n50003 , n227762 );
and ( n50004 , n50003 , n44227 );
nor ( n50005 , n227763 , n50004 );
not ( n50006 , n50005 );
or ( n50007 , n49999 , n50006 );
or ( n50008 , n50005 , n49998 );
nand ( n50009 , n50007 , n50008 );
not ( n50010 , n38005 );
nand ( n227772 , n50010 , n37755 );
not ( n227773 , n227772 );
not ( n50013 , n44242 );
or ( n227775 , n227773 , n50013 );
or ( n227776 , n44242 , n227772 );
nand ( n50016 , n227775 , n227776 );
and ( n50017 , n50009 , n50016 );
not ( n50018 , n50009 );
not ( n50019 , n50016 );
and ( n50020 , n50018 , n50019 );
nor ( n50021 , n50017 , n50020 );
not ( n50022 , n50021 );
or ( n50023 , n227751 , n50022 );
not ( n227785 , n50021 );
not ( n227786 , n227750 );
nand ( n50026 , n227785 , n227786 );
nand ( n50027 , n50023 , n50026 );
buf ( n50028 , n50027 );
and ( n50029 , n227738 , n50028 );
not ( n50030 , n227738 );
and ( n50031 , n50021 , n227750 );
not ( n50032 , n50021 );
and ( n50033 , n50032 , n227786 );
nor ( n227795 , n50031 , n50033 );
buf ( n227796 , n227795 );
and ( n50036 , n50030 , n227796 );
nor ( n50037 , n50029 , n50036 );
nand ( n50038 , n50037 , n205649 );
buf ( n50039 , n29898 );
not ( n227801 , n50039 );
not ( n227802 , n32899 );
or ( n50042 , n227801 , n227802 );
or ( n50043 , n32899 , n50039 );
nand ( n50044 , n50042 , n50043 );
and ( n50045 , n50044 , n32906 );
not ( n50046 , n50044 );
and ( n50047 , n50046 , n32910 );
nor ( n227809 , n50045 , n50047 );
not ( n227810 , n227809 );
not ( n50050 , n227810 );
not ( n50051 , n31796 );
not ( n50052 , n27759 );
or ( n50053 , n50051 , n50052 );
or ( n50054 , n27762 , n31796 );
nand ( n50055 , n50053 , n50054 );
not ( n50056 , n50055 );
not ( n50057 , n34654 );
or ( n50058 , n50056 , n50057 );
or ( n50059 , n220878 , n50055 );
nand ( n227821 , n50058 , n50059 );
not ( n227822 , n204697 );
not ( n50062 , n28721 );
or ( n50063 , n227822 , n50062 );
not ( n50064 , n204697 );
nand ( n50065 , n50064 , n206479 );
nand ( n50066 , n50063 , n50065 );
and ( n50067 , n50066 , n28725 );
not ( n227829 , n50066 );
buf ( n227830 , n42844 );
not ( n50070 , n227830 );
and ( n50071 , n227829 , n50070 );
nor ( n50072 , n50067 , n50071 );
nand ( n50073 , n227821 , n50072 );
not ( n50074 , n50073 );
or ( n50075 , n50050 , n50074 );
or ( n227837 , n50073 , n227810 );
nand ( n227838 , n50075 , n227837 );
not ( n50078 , n227838 );
not ( n50079 , n50072 );
nand ( n50080 , n50079 , n227809 );
not ( n50081 , n50080 );
buf ( n50082 , n34253 );
xor ( n50083 , n50082 , n40743 );
xnor ( n227845 , n50083 , n49026 );
not ( n227846 , n227845 );
or ( n50086 , n50081 , n227846 );
or ( n227848 , n227845 , n50080 );
nand ( n227849 , n50086 , n227848 );
not ( n50089 , n227849 );
not ( n227851 , n50089 );
not ( n50091 , n46587 );
buf ( n50092 , n30522 );
not ( n50093 , n50092 );
and ( n50094 , n50091 , n50093 );
and ( n227856 , n225682 , n50092 );
nor ( n227857 , n50094 , n227856 );
not ( n50097 , n227857 );
not ( n50098 , n46596 );
or ( n50099 , n50097 , n50098 );
or ( n50100 , n46596 , n227857 );
nand ( n227862 , n50099 , n50100 );
not ( n227863 , n227862 );
not ( n50103 , n44993 );
not ( n50104 , n31333 );
not ( n50105 , n35821 );
or ( n50106 , n50104 , n50105 );
or ( n227868 , n44984 , n31333 );
nand ( n227869 , n50106 , n227868 );
not ( n50109 , n227869 );
or ( n50110 , n50103 , n50109 );
buf ( n50111 , n35861 );
or ( n50112 , n227869 , n50111 );
nand ( n227874 , n50110 , n50112 );
nand ( n227875 , n227863 , n227874 );
not ( n50115 , n204361 );
not ( n50116 , n37127 );
or ( n50117 , n50115 , n50116 );
or ( n50118 , n37127 , n204361 );
nand ( n227880 , n50117 , n50118 );
buf ( n227881 , n34303 );
not ( n50121 , n227881 );
and ( n50122 , n227880 , n50121 );
not ( n50123 , n227880 );
and ( n50124 , n50123 , n44337 );
nor ( n50125 , n50122 , n50124 );
not ( n50126 , n50125 );
and ( n50127 , n227875 , n50126 );
not ( n50128 , n227875 );
and ( n50129 , n50128 , n50125 );
nor ( n50130 , n50127 , n50129 );
not ( n227892 , n50130 );
not ( n227893 , n227892 );
or ( n50133 , n227851 , n227893 );
nand ( n50134 , n227849 , n50130 );
nand ( n50135 , n50133 , n50134 );
not ( n50136 , n25447 );
not ( n50137 , n41113 );
or ( n50138 , n50136 , n50137 );
not ( n50139 , n25447 );
nand ( n50140 , n50139 , n42057 );
nand ( n227902 , n50138 , n50140 );
not ( n227903 , n40418 );
and ( n50143 , n227902 , n227903 );
not ( n50144 , n227902 );
and ( n50145 , n50144 , n37946 );
nor ( n50146 , n50143 , n50145 );
not ( n50147 , n50146 );
not ( n50148 , n36903 );
not ( n50149 , n32240 );
or ( n227911 , n50148 , n50149 );
not ( n227912 , n36903 );
nand ( n50152 , n227912 , n32236 );
nand ( n50153 , n227911 , n50152 );
xor ( n50154 , n50153 , n36071 );
not ( n50155 , n50154 );
nand ( n227917 , n50147 , n50155 );
not ( n227918 , n227917 );
buf ( n50158 , n39204 );
not ( n227920 , n50158 );
not ( n227921 , n227920 );
not ( n50161 , n26310 );
or ( n50162 , n227921 , n50161 );
nand ( n50163 , n26318 , n50158 );
nand ( n50164 , n50162 , n50163 );
and ( n50165 , n50164 , n38305 );
not ( n50166 , n50164 );
not ( n227928 , n38305 );
and ( n227929 , n50166 , n227928 );
nor ( n50169 , n50165 , n227929 );
not ( n50170 , n50169 );
not ( n50171 , n50170 );
not ( n50172 , n50171 );
and ( n50173 , n227918 , n50172 );
and ( n50174 , n227917 , n50171 );
nor ( n227936 , n50173 , n50174 );
and ( n227937 , n50135 , n227936 );
not ( n50177 , n50135 );
not ( n50178 , n227936 );
and ( n50179 , n50177 , n50178 );
nor ( n50180 , n227937 , n50179 );
not ( n50181 , n35107 );
not ( n50182 , n30982 );
not ( n227944 , n43553 );
or ( n227945 , n50182 , n227944 );
buf ( n50185 , n35098 );
nand ( n50186 , n50185 , n30978 );
nand ( n50187 , n227945 , n50186 );
not ( n50188 , n50187 );
not ( n50189 , n50188 );
or ( n50190 , n50181 , n50189 );
nand ( n50191 , n45373 , n50187 );
nand ( n50192 , n50190 , n50191 );
not ( n227954 , n45314 );
not ( n227955 , n32641 );
not ( n50195 , n44157 );
or ( n50196 , n227955 , n50195 );
or ( n50197 , n44157 , n32641 );
nand ( n50198 , n50196 , n50197 );
not ( n227960 , n50198 );
or ( n227961 , n227954 , n227960 );
or ( n50201 , n50198 , n45309 );
nand ( n50202 , n227961 , n50201 );
not ( n50203 , n50202 );
nand ( n50204 , n50192 , n50203 );
not ( n227966 , n39640 );
not ( n227967 , n227966 );
not ( n50207 , n28829 );
or ( n50208 , n227967 , n50207 );
nand ( n50209 , n28816 , n39640 );
nand ( n50210 , n50208 , n50209 );
not ( n227972 , n50210 );
not ( n227973 , n32219 );
or ( n50213 , n227972 , n227973 );
or ( n50214 , n32219 , n50210 );
nand ( n50215 , n50213 , n50214 );
and ( n50216 , n50204 , n50215 );
not ( n50217 , n50204 );
not ( n50218 , n50215 );
and ( n227980 , n50217 , n50218 );
nor ( n227981 , n50216 , n227980 );
not ( n50221 , n227981 );
buf ( n50222 , n34911 );
not ( n50223 , n50222 );
not ( n50224 , n34416 );
or ( n227986 , n50223 , n50224 );
or ( n227987 , n34416 , n50222 );
nand ( n50227 , n227986 , n227987 );
and ( n50228 , n50227 , n204622 );
not ( n50229 , n50227 );
and ( n50230 , n50229 , n204632 );
nor ( n50231 , n50228 , n50230 );
not ( n50232 , n28849 );
not ( n50233 , n37652 );
or ( n50234 , n50232 , n50233 );
not ( n227996 , n28849 );
nand ( n227997 , n227996 , n37649 );
nand ( n50237 , n50234 , n227997 );
and ( n50238 , n50237 , n220845 );
not ( n50239 , n50237 );
and ( n50240 , n50239 , n43073 );
nor ( n50241 , n50238 , n50240 );
not ( n50242 , n50241 );
nand ( n228004 , n50231 , n50242 );
not ( n228005 , n228004 );
not ( n50245 , n204936 );
not ( n228007 , n220535 );
not ( n228008 , n42777 );
or ( n50248 , n228007 , n228008 );
or ( n50249 , n42777 , n220535 );
nand ( n50250 , n50248 , n50249 );
not ( n50251 , n50250 );
not ( n50252 , n216493 );
or ( n50253 , n50251 , n50252 );
or ( n228015 , n50250 , n216493 );
nand ( n228016 , n50253 , n228015 );
not ( n50256 , n228016 );
or ( n50257 , n50245 , n50256 );
or ( n50258 , n228016 , n204936 );
nand ( n50259 , n50257 , n50258 );
not ( n50260 , n50259 );
and ( n50261 , n228005 , n50260 );
and ( n228023 , n228004 , n50259 );
nor ( n228024 , n50261 , n228023 );
not ( n50264 , n228024 );
not ( n50265 , n50264 );
or ( n228027 , n50221 , n50265 );
not ( n228028 , n227981 );
nand ( n50268 , n228028 , n228024 );
nand ( n50269 , n228027 , n50268 );
and ( n50270 , n50180 , n50269 );
not ( n50271 , n50180 );
not ( n228033 , n50269 );
and ( n228034 , n50271 , n228033 );
nor ( n50274 , n50270 , n228034 );
not ( n50275 , n50274 );
or ( n50276 , n50078 , n50275 );
not ( n50277 , n227838 );
and ( n50278 , n50180 , n228033 );
not ( n50279 , n50180 );
and ( n228041 , n50279 , n50269 );
nor ( n228042 , n50278 , n228041 );
nand ( n50282 , n50277 , n228042 );
nand ( n50283 , n50276 , n50282 );
not ( n50284 , n29354 );
not ( n50285 , n31514 );
or ( n228047 , n50284 , n50285 );
not ( n228048 , n29354 );
nand ( n50288 , n228048 , n31527 );
nand ( n50289 , n228047 , n50288 );
and ( n50290 , n50289 , n33849 );
not ( n50291 , n50289 );
not ( n228053 , n33849 );
and ( n228054 , n50291 , n228053 );
nor ( n50294 , n50290 , n228054 );
not ( n50295 , n50294 );
not ( n50296 , n43165 );
not ( n50297 , n37417 );
not ( n50298 , n31899 );
or ( n50299 , n50297 , n50298 );
or ( n228061 , n31899 , n37417 );
nand ( n228062 , n50299 , n228061 );
not ( n50302 , n228062 );
and ( n50303 , n50296 , n50302 );
and ( n50304 , n43165 , n228062 );
nor ( n50305 , n50303 , n50304 );
nand ( n50306 , n50295 , n50305 );
not ( n50307 , n50306 );
not ( n228069 , n32970 );
not ( n228070 , n29908 );
not ( n50310 , n228070 );
or ( n228072 , n228069 , n50310 );
not ( n228073 , n29909 );
or ( n50313 , n228073 , n32970 );
nand ( n50314 , n228072 , n50313 );
and ( n50315 , n50314 , n29948 );
not ( n50316 , n50314 );
and ( n228078 , n50316 , n207706 );
nor ( n228079 , n50315 , n228078 );
not ( n50319 , n228079 );
not ( n50320 , n50319 );
not ( n50321 , n50320 );
and ( n50322 , n50307 , n50321 );
and ( n228084 , n50306 , n50320 );
nor ( n228085 , n50322 , n228084 );
not ( n50325 , n228085 );
xor ( n50326 , n39381 , n206479 );
xor ( n50327 , n50326 , n30099 );
not ( n50328 , n35251 );
not ( n228090 , n36934 );
or ( n228091 , n50328 , n228090 );
or ( n50331 , n36934 , n35251 );
nand ( n228093 , n228091 , n50331 );
and ( n228094 , n228093 , n43636 );
not ( n50334 , n228093 );
buf ( n50335 , n227480 );
and ( n50336 , n50334 , n50335 );
nor ( n50337 , n228094 , n50336 );
not ( n228099 , n50337 );
nand ( n228100 , n50327 , n228099 );
not ( n50340 , n205085 );
not ( n50341 , n32607 );
or ( n50342 , n50340 , n50341 );
not ( n50343 , n205085 );
nand ( n228105 , n50343 , n34763 );
nand ( n228106 , n50342 , n228105 );
and ( n50346 , n228106 , n36415 );
not ( n50347 , n228106 );
and ( n50348 , n50347 , n36411 );
nor ( n50349 , n50346 , n50348 );
not ( n228111 , n50349 );
and ( n228112 , n228100 , n228111 );
not ( n50352 , n228100 );
and ( n50353 , n50352 , n50349 );
nor ( n50354 , n228112 , n50353 );
not ( n50355 , n50354 );
or ( n50356 , n50325 , n50355 );
or ( n50357 , n50354 , n228085 );
nand ( n50358 , n50356 , n50357 );
not ( n228120 , n33657 );
not ( n228121 , n40492 );
and ( n50361 , n228120 , n228121 );
and ( n50362 , n211419 , n40492 );
nor ( n50363 , n50361 , n50362 );
and ( n50364 , n50363 , n34227 );
not ( n50365 , n50363 );
and ( n50366 , n50365 , n34220 );
nor ( n50367 , n50364 , n50366 );
not ( n228129 , n50367 );
not ( n228130 , n204387 );
not ( n50370 , n35017 );
or ( n228132 , n228130 , n50370 );
not ( n228133 , n204387 );
nand ( n50373 , n228133 , n37127 );
nand ( n50374 , n228132 , n50373 );
and ( n50375 , n50374 , n50121 );
not ( n50376 , n50374 );
and ( n228138 , n50376 , n44337 );
nor ( n228139 , n50375 , n228138 );
not ( n50379 , n228139 );
nand ( n50380 , n228129 , n50379 );
not ( n50381 , n50380 );
not ( n50382 , n50381 );
xor ( n228144 , n36822 , n42627 );
buf ( n228145 , n42593 );
xor ( n50385 , n228144 , n228145 );
not ( n50386 , n50385 );
not ( n50387 , n50386 );
or ( n50388 , n50382 , n50387 );
nand ( n228150 , n50385 , n50380 );
nand ( n228151 , n50388 , n228150 );
not ( n50391 , n228151 );
and ( n50392 , n50358 , n50391 );
not ( n50393 , n50358 );
and ( n50394 , n50393 , n228151 );
nor ( n228156 , n50392 , n50394 );
not ( n228157 , n228156 );
not ( n50397 , n207466 );
not ( n50398 , n34700 );
or ( n50399 , n50397 , n50398 );
or ( n50400 , n34700 , n207466 );
nand ( n50401 , n50399 , n50400 );
and ( n50402 , n50401 , n39845 );
not ( n50403 , n50401 );
and ( n50404 , n50403 , n44823 );
nor ( n50405 , n50402 , n50404 );
not ( n50406 , n50405 );
not ( n50407 , n50406 );
not ( n228169 , n27968 );
nor ( n228170 , n27961 , n46084 );
not ( n50410 , n228170 );
not ( n50411 , n37562 );
nand ( n50412 , n50411 , n27961 );
nand ( n50413 , n50410 , n50412 );
not ( n228175 , n50413 );
and ( n228176 , n228169 , n228175 );
and ( n50416 , n27968 , n50413 );
nor ( n50417 , n228176 , n50416 );
not ( n50418 , n27839 );
not ( n50419 , n33760 );
or ( n50420 , n50418 , n50419 );
nand ( n228182 , n33759 , n205597 );
nand ( n228183 , n50420 , n228182 );
not ( n50423 , n228183 );
not ( n50424 , n33764 );
and ( n50425 , n50423 , n50424 );
and ( n50426 , n33764 , n228183 );
nor ( n50427 , n50425 , n50426 );
not ( n50428 , n50427 );
nand ( n50429 , n50417 , n50428 );
not ( n50430 , n50429 );
or ( n50431 , n50407 , n50430 );
or ( n50432 , n50429 , n50406 );
nand ( n228194 , n50431 , n50432 );
not ( n228195 , n228194 );
xor ( n50435 , n29228 , n30200 );
xnor ( n50436 , n50435 , n32916 );
not ( n50437 , n50436 );
not ( n50438 , n25609 );
not ( n228200 , n47958 );
or ( n228201 , n50438 , n228200 );
or ( n50441 , n47958 , n25609 );
nand ( n50442 , n228201 , n50441 );
not ( n50443 , n50442 );
not ( n50444 , n45268 );
and ( n50445 , n50443 , n50444 );
and ( n50446 , n50442 , n45268 );
nor ( n228208 , n50445 , n50446 );
nand ( n228209 , n50437 , n228208 );
not ( n50449 , n228209 );
not ( n228211 , n45672 );
not ( n228212 , n204644 );
buf ( n50452 , n42756 );
not ( n50453 , n50452 );
not ( n50454 , n50453 );
or ( n50455 , n228212 , n50454 );
or ( n50456 , n42760 , n204644 );
nand ( n50457 , n50455 , n50456 );
not ( n50458 , n50457 );
or ( n50459 , n228211 , n50458 );
or ( n228221 , n50457 , n45672 );
nand ( n228222 , n50459 , n228221 );
not ( n50462 , n228222 );
and ( n50463 , n50449 , n50462 );
and ( n50464 , n228209 , n228222 );
nor ( n50465 , n50463 , n50464 );
not ( n50466 , n50465 );
or ( n50467 , n228195 , n50466 );
or ( n50468 , n50465 , n228194 );
nand ( n50469 , n50467 , n50468 );
not ( n228231 , n50469 );
and ( n228232 , n228157 , n228231 );
not ( n50472 , n228157 );
and ( n50473 , n50472 , n50469 );
nor ( n50474 , n228232 , n50473 );
buf ( n50475 , n50474 );
and ( n228237 , n50283 , n50475 );
not ( n228238 , n50283 );
not ( n50478 , n50469 );
not ( n50479 , n228156 );
or ( n50480 , n50478 , n50479 );
nand ( n50481 , n228157 , n228231 );
nand ( n50482 , n50480 , n50481 );
buf ( n50483 , n50482 );
and ( n50484 , n228238 , n50483 );
nor ( n50485 , n228237 , n50484 );
not ( n50486 , n205223 );
nand ( n50487 , n50486 , n205145 );
not ( n228249 , n50487 );
not ( n228250 , n35647 );
and ( n50490 , n228249 , n228250 );
and ( n50491 , n50487 , n35647 );
nor ( n50492 , n50490 , n50491 );
not ( n50493 , n50492 );
nand ( n228255 , n205391 , n205327 );
and ( n228256 , n228255 , n35530 );
not ( n50496 , n228255 );
and ( n228258 , n50496 , n35529 );
nor ( n228259 , n228256 , n228258 );
not ( n50499 , n228259 );
or ( n228261 , n50493 , n50499 );
or ( n228262 , n228259 , n50492 );
nand ( n50502 , n228261 , n228262 );
not ( n228264 , n27855 );
nand ( n228265 , n228264 , n27679 );
not ( n50505 , n35489 );
xor ( n50506 , n228265 , n50505 );
and ( n50507 , n50502 , n50506 );
not ( n50508 , n50502 );
not ( n228270 , n50506 );
and ( n228271 , n50508 , n228270 );
nor ( n50511 , n50507 , n228271 );
not ( n50512 , n50511 );
not ( n50513 , n50512 );
not ( n50514 , n204750 );
nand ( n228276 , n50514 , n204685 );
and ( n228277 , n228276 , n35789 );
not ( n50517 , n228276 );
and ( n50518 , n50517 , n35788 );
nor ( n228280 , n228277 , n50518 );
not ( n228281 , n228280 );
not ( n50521 , n228281 );
not ( n50522 , n204983 );
nand ( n50523 , n204826 , n50522 );
not ( n50524 , n50523 );
not ( n50525 , n35707 );
not ( n228287 , n50525 );
and ( n228288 , n50524 , n228287 );
and ( n50528 , n50523 , n50525 );
nor ( n50529 , n228288 , n50528 );
not ( n50530 , n50529 );
not ( n50531 , n50530 );
or ( n50532 , n50521 , n50531 );
nand ( n50533 , n50529 , n228280 );
nand ( n50534 , n50532 , n50533 );
not ( n50535 , n50534 );
not ( n228297 , n50535 );
or ( n228298 , n50513 , n228297 );
nand ( n50538 , n50511 , n50534 );
nand ( n50539 , n228298 , n50538 );
buf ( n50540 , n50539 );
not ( n50541 , n50540 );
buf ( n50542 , n25876 );
not ( n50543 , n50542 );
not ( n228305 , n31430 );
nand ( n228306 , n204510 , n204445 );
not ( n50546 , n228306 );
or ( n50547 , n228305 , n50546 );
not ( n50548 , n31431 );
or ( n50549 , n228306 , n50548 );
nand ( n228311 , n50547 , n50549 );
not ( n228312 , n228311 );
not ( n50552 , n35441 );
or ( n50553 , n228312 , n50552 );
or ( n50554 , n35441 , n228311 );
nand ( n50555 , n50553 , n50554 );
not ( n228317 , n25872 );
not ( n228318 , n25686 );
nand ( n50558 , n228317 , n228318 );
not ( n50559 , n31235 );
and ( n50560 , n50558 , n50559 );
not ( n50561 , n50558 );
and ( n50562 , n50561 , n31235 );
nor ( n50563 , n50560 , n50562 );
not ( n228325 , n50563 );
and ( n228326 , n50555 , n228325 );
not ( n50566 , n50555 );
and ( n50567 , n50566 , n50563 );
nor ( n50568 , n228326 , n50567 );
not ( n50569 , n50568 );
not ( n228331 , n31083 );
not ( n228332 , n26151 );
nand ( n50572 , n25980 , n228332 );
not ( n228334 , n50572 );
or ( n228335 , n228331 , n228334 );
or ( n50575 , n50572 , n31083 );
nand ( n50576 , n228335 , n50575 );
not ( n50577 , n50576 );
not ( n50578 , n50577 );
nand ( n50579 , n26223 , n26413 );
not ( n50580 , n50579 );
not ( n50581 , n31139 );
and ( n50582 , n50580 , n50581 );
and ( n50583 , n50579 , n31139 );
nor ( n228345 , n50582 , n50583 );
not ( n228346 , n228345 );
not ( n50586 , n228346 );
or ( n50587 , n50578 , n50586 );
nand ( n50588 , n228345 , n50576 );
nand ( n50589 , n50587 , n50588 );
not ( n228351 , n50589 );
not ( n228352 , n228351 );
and ( n50592 , n50569 , n228352 );
and ( n50593 , n50568 , n228351 );
nor ( n50594 , n50592 , n50593 );
not ( n50595 , n50594 );
not ( n228357 , n50595 );
or ( n228358 , n50543 , n228357 );
or ( n50598 , n50595 , n50542 );
nand ( n50599 , n228358 , n50598 );
not ( n50600 , n50599 );
not ( n50601 , n50600 );
or ( n228363 , n50541 , n50601 );
xor ( n228364 , n50534 , n50511 );
buf ( n50604 , n228364 );
nand ( n228366 , n50604 , n50599 );
nand ( n228367 , n228363 , n228366 );
not ( n50607 , n228367 );
nand ( n50608 , n50485 , n50607 );
or ( n50609 , n50038 , n50608 );
not ( n50610 , n50485 );
not ( n228372 , n50037 );
or ( n228373 , n50610 , n228372 );
nor ( n50613 , n50607 , n33254 );
nand ( n50614 , n228373 , n50613 );
buf ( n50615 , n41944 );
nand ( n228377 , n50615 , n31765 );
nand ( n228378 , n50609 , n50614 , n228377 );
buf ( n228379 , n228378 );
not ( n228380 , n46832 );
not ( n50620 , n46806 );
nand ( n228382 , n228380 , n50620 );
not ( n228383 , n33404 );
not ( n50623 , n29408 );
not ( n228385 , n40168 );
or ( n228386 , n50623 , n228385 );
or ( n50626 , n40168 , n29408 );
nand ( n50627 , n228386 , n50626 );
not ( n50628 , n50627 );
or ( n50629 , n228383 , n50628 );
not ( n228391 , n50627 );
nand ( n228392 , n228391 , n42159 );
nand ( n50632 , n50629 , n228392 );
not ( n50633 , n50632 );
and ( n50634 , n228382 , n50633 );
not ( n50635 , n228382 );
and ( n228397 , n50635 , n50632 );
nor ( n228398 , n50634 , n228397 );
not ( n50638 , n228398 );
buf ( n50639 , RI1745a0f0_1297);
nor ( n50640 , n34299 , n50639 );
not ( n50641 , n50640 );
nand ( n228403 , n34299 , n50639 );
nand ( n228404 , n50641 , n228403 );
not ( n50644 , n228404 );
not ( n50645 , n34265 );
and ( n50646 , n50644 , n50645 );
not ( n50647 , n34264 );
and ( n50648 , n228404 , n50647 );
nor ( n50649 , n50646 , n50648 );
not ( n50650 , n50649 );
not ( n228412 , n50650 );
xor ( n228413 , n41007 , n41519 );
xnor ( n50653 , n228413 , n225459 );
not ( n50654 , n50653 );
nand ( n50655 , n50654 , n224555 );
not ( n50656 , n50655 );
or ( n50657 , n228412 , n50656 );
not ( n50658 , n46791 );
nand ( n228420 , n50658 , n50654 );
or ( n228421 , n228420 , n50650 );
nand ( n50661 , n50657 , n228421 );
not ( n50662 , n50661 );
nand ( n50663 , n50633 , n46831 );
not ( n50664 , n50663 );
not ( n50665 , n40562 );
not ( n228427 , n35563 );
not ( n228428 , n40523 );
or ( n50668 , n228427 , n228428 );
or ( n50669 , n40523 , n35563 );
nand ( n50670 , n50668 , n50669 );
not ( n50671 , n50670 );
or ( n228433 , n50665 , n50671 );
or ( n228434 , n50670 , n40564 );
nand ( n50674 , n228433 , n228434 );
not ( n50675 , n50674 );
and ( n50676 , n50664 , n50675 );
and ( n50677 , n50663 , n50674 );
nor ( n228439 , n50676 , n50677 );
not ( n228440 , n228439 );
or ( n50680 , n50662 , n228440 );
or ( n50681 , n228439 , n50661 );
nand ( n50682 , n50680 , n50681 );
not ( n50683 , n34224 );
not ( n228445 , n32135 );
or ( n228446 , n50683 , n228445 );
not ( n50686 , n34224 );
nand ( n50687 , n50686 , n32139 );
nand ( n50688 , n228446 , n50687 );
and ( n50689 , n50688 , n32182 );
not ( n50690 , n50688 );
not ( n50691 , n32176 );
and ( n50692 , n50690 , n50691 );
nor ( n50693 , n50689 , n50692 );
not ( n50694 , n50693 );
nand ( n228456 , n50694 , n46868 );
not ( n228457 , n39344 );
not ( n50697 , n32406 );
or ( n228459 , n228457 , n50697 );
nand ( n228460 , n33013 , n39347 );
nand ( n50700 , n228459 , n228460 );
not ( n50701 , n50700 );
not ( n50702 , n32443 );
and ( n50703 , n50701 , n50702 );
and ( n228465 , n50700 , n32443 );
nor ( n228466 , n50703 , n228465 );
and ( n50706 , n228456 , n228466 );
not ( n50707 , n228456 );
not ( n228469 , n228466 );
and ( n228470 , n50707 , n228469 );
nor ( n228471 , n50706 , n228470 );
not ( n228472 , n228471 );
and ( n50712 , n50682 , n228472 );
not ( n50713 , n50682 );
and ( n50714 , n50713 , n228471 );
nor ( n50715 , n50712 , n50714 );
not ( n50716 , n50715 );
not ( n50717 , n47696 );
not ( n228479 , n32323 );
or ( n228480 , n50717 , n228479 );
not ( n50720 , n47696 );
nand ( n50721 , n50720 , n32326 );
nand ( n50722 , n228480 , n50721 );
not ( n50723 , n50722 );
not ( n228485 , n37398 );
and ( n228486 , n50723 , n228485 );
and ( n50726 , n50722 , n37398 );
nor ( n50727 , n228486 , n50726 );
nand ( n50728 , n46927 , n50727 );
not ( n50729 , n50728 );
xor ( n50730 , n36913 , n37746 );
xnor ( n50731 , n50730 , n32236 );
not ( n228493 , n50731 );
not ( n228494 , n228493 );
or ( n50734 , n50729 , n228494 );
or ( n50735 , n228493 , n50728 );
nand ( n50736 , n50734 , n50735 );
not ( n50737 , n50736 );
not ( n228499 , n50737 );
buf ( n228500 , n41250 );
not ( n50740 , n228500 );
not ( n50741 , n50740 );
not ( n50742 , n33444 );
or ( n50743 , n50741 , n50742 );
nand ( n50744 , n34594 , n228500 );
nand ( n50745 , n50743 , n50744 );
and ( n228507 , n50745 , n40772 );
not ( n228508 , n50745 );
and ( n50748 , n228508 , n40773 );
nor ( n50749 , n228507 , n50748 );
not ( n50750 , n50749 );
nand ( n50751 , n46883 , n50750 );
not ( n228513 , n50751 );
not ( n228514 , n224490 );
and ( n50754 , n228513 , n228514 );
nand ( n50755 , n46883 , n50750 );
and ( n50756 , n50755 , n224490 );
nor ( n50757 , n50754 , n50756 );
not ( n50758 , n50757 );
not ( n50759 , n50758 );
or ( n228521 , n228499 , n50759 );
nand ( n228522 , n50757 , n50736 );
nand ( n50762 , n228521 , n228522 );
not ( n50763 , n50762 );
and ( n50764 , n50716 , n50763 );
and ( n228526 , n50762 , n50715 );
nor ( n228527 , n50764 , n228526 );
not ( n50767 , n228527 );
or ( n50768 , n50638 , n50767 );
not ( n50769 , n228398 );
not ( n50770 , n50762 );
not ( n228532 , n50715 );
or ( n228533 , n50770 , n228532 );
not ( n50773 , n50715 );
not ( n50774 , n50762 );
nand ( n50775 , n50773 , n50774 );
nand ( n50776 , n228533 , n50775 );
nand ( n228538 , n50769 , n50776 );
nand ( n228539 , n50768 , n228538 );
buf ( n50779 , n39995 );
not ( n50780 , n50779 );
not ( n50781 , n38747 );
or ( n50782 , n50780 , n50781 );
or ( n50783 , n38747 , n50779 );
nand ( n50784 , n50782 , n50783 );
and ( n228546 , n50784 , n32457 );
not ( n228547 , n50784 );
and ( n50787 , n228547 , n32454 );
nor ( n50788 , n228546 , n50787 );
not ( n50789 , n50788 );
not ( n50790 , n50789 );
not ( n50791 , n41258 );
not ( n50792 , n34035 );
not ( n228554 , n41303 );
or ( n228555 , n50792 , n228554 );
nand ( n50795 , n219052 , n34031 );
nand ( n50796 , n228555 , n50795 );
not ( n50797 , n50796 );
or ( n50798 , n50791 , n50797 );
or ( n228560 , n41258 , n50796 );
nand ( n228561 , n50798 , n228560 );
not ( n50801 , n228561 );
nand ( n50802 , n50801 , n47139 );
not ( n50803 , n50802 );
or ( n50804 , n50790 , n50803 );
or ( n228566 , n50802 , n50789 );
nand ( n228567 , n50804 , n228566 );
not ( n50807 , n204277 );
not ( n228569 , n36751 );
or ( n228570 , n50807 , n228569 );
not ( n50810 , n204277 );
nand ( n50811 , n50810 , n37303 );
nand ( n50812 , n228570 , n50811 );
and ( n50813 , n50812 , n36758 );
not ( n50814 , n50812 );
and ( n50815 , n50814 , n208210 );
nor ( n228577 , n50813 , n50815 );
not ( n228578 , n228577 );
nand ( n50818 , n47103 , n228578 );
not ( n50819 , n31671 );
not ( n50820 , n34654 );
or ( n50821 , n50819 , n50820 );
not ( n50822 , n31671 );
nand ( n50823 , n50822 , n34644 );
nand ( n50824 , n50821 , n50823 );
not ( n50825 , n42372 );
and ( n228587 , n50824 , n50825 );
not ( n228588 , n50824 );
and ( n50828 , n228588 , n42372 );
nor ( n50829 , n228587 , n50828 );
not ( n50830 , n50829 );
and ( n228592 , n50818 , n50830 );
not ( n228593 , n50818 );
and ( n50833 , n228593 , n50829 );
nor ( n50834 , n228592 , n50833 );
not ( n50835 , n50834 );
and ( n50836 , n228567 , n50835 );
not ( n50837 , n228567 );
and ( n50838 , n50837 , n50834 );
nor ( n50839 , n50836 , n50838 );
not ( n50840 , n50839 );
not ( n228602 , n213777 );
not ( n228603 , n204949 );
and ( n50843 , n228602 , n228603 );
and ( n50844 , n213777 , n204949 );
nor ( n228606 , n50843 , n50844 );
and ( n228607 , n228606 , n221434 );
not ( n50847 , n228606 );
and ( n50848 , n50847 , n40862 );
nor ( n50849 , n228607 , n50848 );
not ( n228611 , n50849 );
nand ( n228612 , n46983 , n228611 );
not ( n50852 , n228612 );
not ( n50853 , n43259 );
not ( n50854 , n41856 );
or ( n50855 , n50853 , n50854 );
or ( n50856 , n46810 , n43259 );
nand ( n50857 , n50855 , n50856 );
not ( n228619 , n50857 );
not ( n228620 , n46815 );
and ( n50860 , n228619 , n228620 );
and ( n50861 , n50857 , n217819 );
nor ( n50862 , n50860 , n50861 );
not ( n50863 , n50862 );
not ( n228625 , n50863 );
and ( n228626 , n50852 , n228625 );
and ( n50866 , n228612 , n50863 );
nor ( n50867 , n228626 , n50866 );
not ( n50868 , n50867 );
not ( n50869 , n38889 );
not ( n228631 , n26222 );
or ( n228632 , n50869 , n228631 );
or ( n50872 , n26222 , n38889 );
nand ( n50873 , n228632 , n50872 );
and ( n50874 , n50873 , n47879 );
not ( n50875 , n50873 );
and ( n228637 , n50875 , n26205 );
nor ( n228638 , n50874 , n228637 );
nand ( n50878 , n228638 , n47024 );
not ( n50879 , n37876 );
not ( n50880 , n44932 );
or ( n50881 , n50879 , n50880 );
or ( n228643 , n44932 , n37876 );
nand ( n228644 , n50881 , n228643 );
not ( n50884 , n38130 );
and ( n50885 , n228644 , n50884 );
not ( n228647 , n228644 );
and ( n228648 , n228647 , n222700 );
nor ( n50888 , n50885 , n228648 );
not ( n50889 , n50888 );
xor ( n50890 , n50878 , n50889 );
not ( n50891 , n50890 );
or ( n228653 , n50868 , n50891 );
or ( n228654 , n50890 , n50867 );
nand ( n50894 , n228653 , n228654 );
not ( n50895 , n30971 );
and ( n50896 , n35872 , n31008 );
not ( n50897 , n35872 );
and ( n228659 , n50897 , n35753 );
nor ( n228660 , n50896 , n228659 );
not ( n50900 , n228660 );
or ( n50901 , n50895 , n50900 );
not ( n50902 , n30853 );
or ( n50903 , n228660 , n50902 );
nand ( n228665 , n50901 , n50903 );
not ( n228666 , n228665 );
nand ( n50906 , n47056 , n228666 );
buf ( n228668 , n32825 );
not ( n228669 , n228668 );
not ( n50909 , n37537 );
or ( n50910 , n228669 , n50909 );
or ( n50911 , n37537 , n228668 );
nand ( n50912 , n50910 , n50911 );
and ( n228674 , n38037 , n50912 );
not ( n228675 , n38037 );
not ( n50915 , n50912 );
and ( n50916 , n228675 , n50915 );
nor ( n50917 , n228674 , n50916 );
buf ( n50918 , n50917 );
xor ( n228680 , n50906 , n50918 );
not ( n228681 , n228680 );
and ( n50921 , n50894 , n228681 );
not ( n228683 , n50894 );
and ( n228684 , n228683 , n228680 );
nor ( n50924 , n50921 , n228684 );
not ( n50925 , n50924 );
or ( n50926 , n50840 , n50925 );
not ( n50927 , n50839 );
not ( n228689 , n50924 );
nand ( n228690 , n50927 , n228689 );
nand ( n50930 , n50926 , n228690 );
buf ( n50931 , n50930 );
and ( n50932 , n228539 , n50931 );
not ( n50933 , n228539 );
not ( n228695 , n50924 );
not ( n228696 , n228695 );
not ( n50936 , n50839 );
not ( n50937 , n50936 );
and ( n50938 , n228696 , n50937 );
and ( n50939 , n228695 , n50936 );
nor ( n50940 , n50938 , n50939 );
buf ( n50941 , n50940 );
and ( n50942 , n50933 , n50941 );
nor ( n50943 , n50932 , n50942 );
buf ( n50944 , n35427 );
not ( n50945 , n50944 );
nand ( n228707 , n50943 , n50945 );
not ( n228708 , n205095 );
not ( n50948 , n35856 );
and ( n50949 , n228708 , n50948 );
not ( n50950 , n205096 );
and ( n50951 , n50950 , n35856 );
nor ( n50952 , n50949 , n50951 );
and ( n50953 , n50952 , n33300 );
not ( n228715 , n50952 );
not ( n228716 , n33300 );
and ( n50956 , n228715 , n228716 );
nor ( n50957 , n50953 , n50956 );
not ( n50958 , n50957 );
not ( n50959 , n30204 );
not ( n228721 , n50959 );
not ( n228722 , n27721 );
or ( n50962 , n228721 , n228722 );
or ( n228724 , n27721 , n50959 );
nand ( n228725 , n50962 , n228724 );
and ( n50965 , n228725 , n27759 );
not ( n50966 , n228725 );
and ( n50967 , n50966 , n27763 );
nor ( n50968 , n50965 , n50967 );
not ( n50969 , n50968 );
nand ( n50970 , n50958 , n50969 );
not ( n228732 , n46664 );
not ( n228733 , n38821 );
and ( n50973 , n228732 , n228733 );
and ( n50974 , n46664 , n38821 );
nor ( n50975 , n50973 , n50974 );
and ( n50976 , n50975 , n46668 );
not ( n228738 , n50975 );
and ( n228739 , n228738 , n46671 );
nor ( n50979 , n50976 , n228739 );
not ( n50980 , n50979 );
and ( n50981 , n50970 , n50980 );
not ( n50982 , n50970 );
and ( n50983 , n50982 , n50979 );
nor ( n50984 , n50981 , n50983 );
not ( n228746 , n50984 );
xor ( n228747 , n30258 , n37212 );
xnor ( n50987 , n228747 , n204631 );
buf ( n228749 , n34506 );
not ( n228750 , n228749 );
not ( n50990 , n228750 );
not ( n50991 , n43635 );
or ( n50992 , n50990 , n50991 );
nand ( n50993 , n227480 , n228749 );
nand ( n50994 , n50992 , n50993 );
xor ( n50995 , n44135 , n50994 );
nand ( n50996 , n50987 , n50995 );
not ( n228758 , n50996 );
not ( n228759 , n31869 );
not ( n228760 , n25463 );
and ( n228761 , n228759 , n228760 );
and ( n51001 , n40418 , n25463 );
nor ( n51002 , n228761 , n51001 );
and ( n51003 , n51002 , n31900 );
not ( n51004 , n51002 );
and ( n228766 , n51004 , n31907 );
nor ( n228767 , n51003 , n228766 );
not ( n51007 , n228767 );
and ( n51008 , n228758 , n51007 );
and ( n51009 , n50996 , n228767 );
nor ( n51010 , n51008 , n51009 );
not ( n228772 , n51010 );
nand ( n228773 , n50957 , n50980 );
not ( n51013 , n204312 );
not ( n228775 , n208165 );
or ( n228776 , n51013 , n228775 );
not ( n51016 , n204312 );
nand ( n51017 , n51016 , n37762 );
nand ( n51018 , n228776 , n51017 );
not ( n51019 , n51018 );
not ( n51020 , n33886 );
and ( n51021 , n51019 , n51020 );
and ( n228783 , n33886 , n51018 );
nor ( n228784 , n51021 , n228783 );
and ( n51024 , n228773 , n228784 );
not ( n51025 , n228773 );
not ( n51026 , n228784 );
and ( n51027 , n51025 , n51026 );
nor ( n228789 , n51024 , n51027 );
not ( n228790 , n228789 );
or ( n51030 , n228772 , n228790 );
or ( n51031 , n228789 , n51010 );
nand ( n51032 , n51030 , n51031 );
buf ( n51033 , n31613 );
xor ( n228795 , n31316 , n51033 );
xnor ( n228796 , n228795 , n28122 );
not ( n51036 , n223859 );
not ( n51037 , n29135 );
not ( n51038 , n39400 );
or ( n51039 , n51037 , n51038 );
or ( n228801 , n39400 , n29135 );
nand ( n228802 , n51039 , n228801 );
not ( n51042 , n228802 );
or ( n51043 , n51036 , n51042 );
or ( n51044 , n228802 , n223859 );
nand ( n51045 , n51043 , n51044 );
not ( n228807 , n51045 );
nand ( n228808 , n228796 , n228807 );
not ( n51048 , n228808 );
not ( n51049 , n28011 );
not ( n51050 , n204473 );
or ( n51051 , n51049 , n51050 );
or ( n51052 , n28011 , n204473 );
nand ( n51053 , n51051 , n51052 );
xor ( n51054 , n51053 , n204505 );
not ( n51055 , n51054 );
not ( n228817 , n51055 );
and ( n228818 , n51048 , n228817 );
nand ( n51058 , n228796 , n228807 );
and ( n228820 , n51058 , n51055 );
nor ( n51060 , n228818 , n228820 );
not ( n51061 , n51060 );
and ( n51062 , n51032 , n51061 );
not ( n51063 , n51032 );
and ( n51064 , n51063 , n51060 );
nor ( n51065 , n51062 , n51064 );
buf ( n228827 , n51065 );
not ( n228828 , n38438 );
not ( n51068 , n209942 );
or ( n51069 , n228828 , n51068 );
or ( n51070 , n32175 , n38438 );
nand ( n51071 , n51069 , n51070 );
and ( n228833 , n51071 , n42097 );
not ( n228834 , n51071 );
and ( n51074 , n228834 , n42092 );
nor ( n51075 , n228833 , n51074 );
not ( n51076 , n51075 );
not ( n51077 , n51076 );
not ( n51078 , n31254 );
not ( n51079 , n27781 );
and ( n51080 , n51078 , n51079 );
and ( n51081 , n31254 , n27781 );
nor ( n228843 , n51080 , n51081 );
and ( n228844 , n228843 , n31264 );
not ( n51084 , n228843 );
and ( n51085 , n51084 , n31273 );
nor ( n51086 , n228844 , n51085 );
not ( n51087 , n51086 );
buf ( n51088 , n33283 );
not ( n51089 , n51088 );
not ( n228851 , n51089 );
not ( n228852 , n36411 );
or ( n51092 , n228851 , n228852 );
nand ( n51093 , n36415 , n51088 );
nand ( n51094 , n51092 , n51093 );
and ( n51095 , n51094 , n26047 );
not ( n228857 , n51094 );
and ( n228858 , n228857 , n35028 );
nor ( n51098 , n51095 , n228858 );
not ( n51099 , n51098 );
nand ( n51100 , n51087 , n51099 );
not ( n51101 , n51100 );
or ( n228863 , n51077 , n51101 );
not ( n228864 , n51098 );
nand ( n51104 , n228864 , n51087 );
or ( n51105 , n51104 , n51076 );
nand ( n51106 , n228863 , n51105 );
not ( n51107 , n51106 );
not ( n228869 , n32082 );
and ( n228870 , n205007 , n32053 );
not ( n51110 , n205007 );
and ( n51111 , n51110 , n32050 );
nor ( n51112 , n228870 , n51111 );
not ( n51113 , n51112 );
and ( n51114 , n228869 , n51113 );
and ( n51115 , n32082 , n51112 );
nor ( n228877 , n51114 , n51115 );
not ( n228878 , RI174a68d8_924);
and ( n51118 , n32234 , n228878 );
not ( n51119 , n32234 );
and ( n51120 , n51119 , n32231 );
nor ( n51121 , n51118 , n51120 );
not ( n51122 , n51121 );
not ( n51123 , n37346 );
or ( n51124 , n51122 , n51123 );
not ( n51125 , n51121 );
nand ( n51126 , n51125 , n43839 );
nand ( n228888 , n51124 , n51126 );
and ( n228889 , n228888 , n37356 );
not ( n51129 , n228888 );
and ( n51130 , n51129 , n37353 );
nor ( n51131 , n228889 , n51130 );
nand ( n51132 , n228877 , n51131 );
not ( n228894 , n51132 );
not ( n228895 , n224315 );
not ( n51135 , n35704 );
or ( n51136 , n228895 , n51135 );
or ( n51137 , n35704 , n224315 );
nand ( n51138 , n51136 , n51137 );
and ( n228900 , n51138 , n224686 );
not ( n228901 , n51138 );
and ( n51141 , n228901 , n46921 );
nor ( n51142 , n228900 , n51141 );
not ( n51143 , n51142 );
not ( n51144 , n51143 );
and ( n51145 , n228894 , n51144 );
and ( n51146 , n51132 , n51143 );
nor ( n228908 , n51145 , n51146 );
not ( n228909 , n228908 );
and ( n51149 , n51107 , n228909 );
and ( n51150 , n51106 , n228908 );
nor ( n51151 , n51149 , n51150 );
buf ( n51152 , n51151 );
and ( n51153 , n228827 , n51152 );
not ( n51154 , n228827 );
not ( n51155 , n51152 );
and ( n228917 , n51154 , n51155 );
nor ( n228918 , n51153 , n228917 );
not ( n51158 , n228918 );
or ( n51159 , n228746 , n51158 );
not ( n51160 , n50984 );
not ( n51161 , n51151 );
not ( n228923 , n51065 );
or ( n228924 , n51161 , n228923 );
not ( n51164 , n51065 );
not ( n51165 , n51151 );
nand ( n51166 , n51164 , n51165 );
nand ( n51167 , n228924 , n51166 );
nand ( n228929 , n51160 , n51167 );
nand ( n228930 , n51159 , n228929 );
not ( n51170 , n31834 );
nand ( n51171 , n51170 , n31909 );
not ( n51172 , n51171 );
not ( n51173 , n34806 );
not ( n228935 , n29117 );
or ( n228936 , n51173 , n228935 );
not ( n51176 , n34806 );
nand ( n51177 , n51176 , n29123 );
nand ( n51178 , n228936 , n51177 );
and ( n51179 , n51178 , n29175 );
not ( n51180 , n51178 );
and ( n51181 , n51180 , n29162 );
nor ( n51182 , n51179 , n51181 );
not ( n228944 , n51182 );
not ( n228945 , n228944 );
and ( n51185 , n51172 , n228945 );
and ( n51186 , n51171 , n228944 );
nor ( n51187 , n51185 , n51186 );
nand ( n51188 , n31744 , n31937 );
not ( n228950 , n51188 );
not ( n228951 , n33094 );
not ( n51191 , n39065 );
or ( n51192 , n228951 , n51191 );
or ( n51193 , n39065 , n33094 );
nand ( n51194 , n51192 , n51193 );
not ( n228956 , n51194 );
not ( n228957 , n39020 );
and ( n51197 , n228956 , n228957 );
and ( n51198 , n51194 , n39020 );
nor ( n51199 , n51197 , n51198 );
not ( n51200 , n51199 );
not ( n51201 , n51200 );
and ( n51202 , n228950 , n51201 );
and ( n228964 , n51188 , n51200 );
nor ( n228965 , n51202 , n228964 );
xor ( n51205 , n51187 , n228965 );
buf ( n51206 , n34763 );
xor ( n51207 , n205133 , n51206 );
xnor ( n51208 , n51207 , n41415 );
not ( n228970 , n51208 );
not ( n228971 , n228970 );
not ( n51211 , n32087 );
nand ( n228973 , n51211 , n31947 );
not ( n228974 , n228973 );
or ( n51214 , n228971 , n228974 );
or ( n51215 , n228973 , n228970 );
nand ( n51216 , n51214 , n51215 );
xnor ( n51217 , n51205 , n51216 );
not ( n51218 , n32447 );
nand ( n51219 , n51218 , n32364 );
not ( n228981 , n51219 );
buf ( n228982 , RI174a6c20_923);
and ( n51222 , n42590 , n228982 );
not ( n51223 , n42590 );
and ( n51224 , n51223 , n42587 );
nor ( n51225 , n51222 , n51224 );
not ( n228987 , n51225 );
not ( n228988 , n215580 );
or ( n51228 , n228987 , n228988 );
or ( n51229 , n44061 , n51225 );
nand ( n51230 , n51228 , n51229 );
buf ( n51231 , n34564 );
and ( n51232 , n51230 , n51231 );
not ( n51233 , n51230 );
and ( n228995 , n51233 , n43326 );
nor ( n228996 , n51232 , n228995 );
not ( n51236 , n228996 );
not ( n51237 , n51236 );
and ( n51238 , n228981 , n51237 );
and ( n51239 , n51219 , n51236 );
nor ( n51240 , n51238 , n51239 );
not ( n51241 , n51240 );
not ( n229003 , n32185 );
not ( n229004 , n32243 );
nand ( n51244 , n229003 , n229004 );
not ( n51245 , n29149 );
not ( n51246 , n45898 );
or ( n51247 , n51245 , n51246 );
or ( n51248 , n45898 , n29149 );
nand ( n51249 , n51247 , n51248 );
and ( n229011 , n51249 , n223859 );
not ( n229012 , n51249 );
not ( n51252 , n223859 );
and ( n229014 , n229012 , n51252 );
nor ( n229015 , n229011 , n229014 );
and ( n51255 , n51244 , n229015 );
not ( n51256 , n51244 );
not ( n51257 , n229015 );
and ( n51258 , n51256 , n51257 );
nor ( n229020 , n51255 , n51258 );
not ( n229021 , n229020 );
or ( n51261 , n51241 , n229021 );
or ( n51262 , n229020 , n51240 );
nand ( n51263 , n51261 , n51262 );
and ( n51264 , n51217 , n51263 );
not ( n51265 , n51217 );
not ( n51266 , n51263 );
and ( n229028 , n51265 , n51266 );
nor ( n229029 , n51264 , n229028 );
buf ( n51269 , n229029 );
and ( n51270 , n228930 , n51269 );
not ( n51271 , n228930 );
not ( n51272 , n51269 );
and ( n51273 , n51271 , n51272 );
nor ( n51274 , n51270 , n51273 );
not ( n229036 , n221837 );
not ( n229037 , n221824 );
nand ( n51277 , n229036 , n229037 );
not ( n229039 , n51277 );
not ( n229040 , n220602 );
or ( n51280 , n229039 , n229040 );
or ( n51281 , n220602 , n51277 );
nand ( n51282 , n51280 , n51281 );
not ( n51283 , n51282 );
not ( n51284 , n51283 );
not ( n51285 , n220545 );
nand ( n51286 , n51285 , n44117 );
not ( n51287 , n51286 );
not ( n229049 , n42730 );
not ( n229050 , n229049 );
and ( n51290 , n51287 , n229050 );
and ( n51291 , n51286 , n229049 );
nor ( n51292 , n51290 , n51291 );
not ( n51293 , n51292 );
not ( n51294 , n51293 );
not ( n51295 , n49971 );
not ( n229057 , n51295 );
or ( n229058 , n51294 , n229057 );
nand ( n51298 , n49971 , n51292 );
nand ( n229060 , n229058 , n51298 );
or ( n229061 , n220602 , n229036 );
and ( n51301 , n229061 , n42854 );
not ( n229063 , n229061 );
and ( n229064 , n229063 , n220614 );
nor ( n51304 , n51301 , n229064 );
and ( n51305 , n229060 , n51304 );
not ( n51306 , n229060 );
not ( n51307 , n51304 );
and ( n229069 , n51306 , n51307 );
nor ( n229070 , n51305 , n229069 );
not ( n51310 , n42896 );
not ( n51311 , n51310 );
nand ( n51312 , n221804 , n220667 );
not ( n51313 , n51312 );
or ( n51314 , n51311 , n51313 );
or ( n51315 , n51312 , n51310 );
nand ( n229077 , n51314 , n51315 );
not ( n229078 , n229077 );
not ( n51318 , n229078 );
not ( n229080 , n42982 );
nand ( n229081 , n221769 , n229080 );
not ( n51321 , n229081 );
not ( n51322 , n42970 );
and ( n51323 , n51321 , n51322 );
and ( n229085 , n229081 , n42970 );
nor ( n229086 , n51323 , n229085 );
not ( n229087 , n229086 );
not ( n229088 , n229087 );
or ( n51328 , n51318 , n229088 );
nand ( n51329 , n229086 , n229077 );
nand ( n51330 , n51328 , n51329 );
not ( n51331 , n51330 );
and ( n229093 , n229070 , n51331 );
not ( n229094 , n229070 );
and ( n51334 , n229094 , n51330 );
nor ( n51335 , n229093 , n51334 );
not ( n51336 , n51335 );
not ( n229098 , n51336 );
or ( n229099 , n51284 , n229098 );
and ( n51339 , n229070 , n51331 );
not ( n51340 , n229070 );
and ( n51341 , n51340 , n51330 );
nor ( n51342 , n51339 , n51341 );
not ( n51343 , n51342 );
or ( n229105 , n51343 , n51283 );
nand ( n229106 , n229099 , n229105 );
not ( n51346 , n229106 );
not ( n51347 , n38222 );
and ( n51348 , n51346 , n51347 );
buf ( n51349 , n38222 );
and ( n229111 , n229106 , n51349 );
nor ( n229112 , n51348 , n229111 );
nand ( n51352 , n51274 , n229112 );
or ( n51353 , n228707 , n51352 );
not ( n51354 , n50943 );
not ( n51355 , n51274 );
or ( n51356 , n51354 , n51355 );
nor ( n51357 , n229112 , n31571 );
nand ( n51358 , n51356 , n51357 );
nand ( n51359 , n31577 , n42972 );
nand ( n229121 , n51353 , n51358 , n51359 );
buf ( n229122 , n229121 );
and ( n51362 , n25326 , RI1754a798_67);
and ( n51363 , n25325 , n25319 , n51362 );
not ( n51364 , RI1754a6a8_69);
nand ( n51365 , n51364 , RI1754a720_68);
nand ( n229127 , n51363 , n51365 );
and ( n229128 , n51363 , RI1754a630_70);
not ( n51368 , n229128 );
and ( n51369 , n229127 , n51368 );
not ( n51370 , RI1754bad0_26);
or ( n51371 , n51369 , n51370 );
not ( n229133 , n226822 );
not ( n229134 , n49059 );
and ( n51374 , n229133 , n229134 );
nor ( n51375 , n51365 , RI1754a5b8_71);
and ( n51376 , n229128 , n51375 );
nor ( n51377 , n51374 , n51376 );
nand ( n229139 , n51371 , n51377 );
buf ( n229140 , n229139 );
not ( n51380 , n26212 );
buf ( n51381 , n31577 );
not ( n51382 , n51381 );
or ( n51383 , n51380 , n51382 );
not ( n229145 , n38817 );
buf ( n229146 , n33562 );
not ( n51386 , n229146 );
not ( n229148 , n51386 );
not ( n229149 , n35357 );
or ( n51389 , n229148 , n229149 );
nand ( n51390 , n38255 , n229146 );
nand ( n51391 , n51389 , n51390 );
not ( n51392 , n51391 );
and ( n229154 , n229145 , n51392 );
and ( n229155 , n35390 , n51391 );
nor ( n51395 , n229154 , n229155 );
not ( n51396 , n51395 );
not ( n51397 , n51396 );
not ( n51398 , n41051 );
not ( n51399 , n37776 );
or ( n51400 , n51398 , n51399 );
or ( n51401 , n37776 , n41051 );
nand ( n51402 , n51400 , n51401 );
and ( n51403 , n51402 , n34191 );
not ( n229165 , n51402 );
and ( n229166 , n229165 , n211419 );
nor ( n51406 , n51403 , n229166 );
not ( n51407 , n51406 );
nand ( n51408 , n51407 , n36028 );
not ( n51409 , n51408 );
or ( n51410 , n51397 , n51409 );
not ( n51411 , n51406 );
nand ( n51412 , n51411 , n36028 );
or ( n229174 , n51412 , n51396 );
nand ( n229175 , n51410 , n229174 );
not ( n51415 , n229175 );
not ( n229177 , n35969 );
nand ( n229178 , n51395 , n51406 );
not ( n51418 , n229178 );
or ( n51419 , n229177 , n51418 );
or ( n51420 , n229178 , n35969 );
nand ( n51421 , n51419 , n51420 );
not ( n51422 , n51421 );
not ( n51423 , n42622 );
not ( n51424 , n51423 );
not ( n51425 , n34557 );
or ( n229187 , n51424 , n51425 );
or ( n229188 , n34557 , n51423 );
nand ( n51428 , n229187 , n229188 );
and ( n229190 , n51428 , n39411 );
not ( n229191 , n51428 );
not ( n51431 , n32652 );
and ( n229193 , n229191 , n51431 );
nor ( n229194 , n229190 , n229193 );
not ( n51434 , n229194 );
nand ( n51435 , n35928 , n51434 );
not ( n51436 , n51435 );
not ( n51437 , n35863 );
and ( n229199 , n51436 , n51437 );
and ( n229200 , n51435 , n35863 );
nor ( n51440 , n229199 , n229200 );
not ( n51441 , n51440 );
or ( n51442 , n51422 , n51441 );
or ( n51443 , n51440 , n51421 );
nand ( n51444 , n51442 , n51443 );
not ( n51445 , n51444 );
not ( n51446 , n26149 );
not ( n51447 , n41169 );
buf ( n229209 , n31634 );
not ( n229210 , n229209 );
and ( n51450 , n51447 , n229210 );
not ( n51451 , n42372 );
and ( n51452 , n51451 , n229209 );
nor ( n51453 , n51450 , n51452 );
not ( n51454 , n51453 );
or ( n51455 , n51446 , n51454 );
or ( n229217 , n51453 , n26149 );
nand ( n229218 , n51455 , n229217 );
not ( n51458 , n229218 );
xor ( n51459 , n25859 , n225379 );
xnor ( n51460 , n51459 , n38839 );
nand ( n51461 , n51458 , n51460 );
not ( n51462 , n51461 );
not ( n51463 , n36104 );
not ( n229225 , n51463 );
not ( n229226 , n229225 );
and ( n51466 , n51462 , n229226 );
not ( n51467 , n229218 );
nand ( n51468 , n51467 , n51460 );
and ( n51469 , n51468 , n229225 );
nor ( n229231 , n51466 , n51469 );
not ( n229232 , n229231 );
or ( n51472 , n51445 , n229232 );
or ( n229234 , n229231 , n51444 );
nand ( n229235 , n51472 , n229234 );
not ( n51475 , n229235 );
not ( n51476 , n51475 );
not ( n51477 , n40041 );
not ( n51478 , n30943 );
or ( n229240 , n51477 , n51478 );
or ( n229241 , n30943 , n40041 );
nand ( n51481 , n229240 , n229241 );
xnor ( n51482 , n51481 , n30898 );
buf ( n51483 , n35912 );
not ( n51484 , n51483 );
not ( n229246 , n30971 );
or ( n229247 , n51484 , n229246 );
or ( n51487 , n30971 , n51483 );
nand ( n229249 , n229247 , n51487 );
buf ( n229250 , n30888 );
and ( n51490 , n229249 , n229250 );
not ( n51491 , n229249 );
not ( n51492 , n229250 );
and ( n51493 , n51491 , n51492 );
nor ( n229255 , n51490 , n51493 );
nand ( n229256 , n51482 , n229255 );
and ( n51496 , n229256 , n36198 );
not ( n229258 , n229256 );
and ( n229259 , n229258 , n36197 );
nor ( n51499 , n51496 , n229259 );
not ( n51500 , n51499 );
not ( n51501 , n36259 );
buf ( n51502 , n204424 );
and ( n51503 , n51502 , n37120 );
not ( n229265 , n51502 );
and ( n229266 , n229265 , n218917 );
nor ( n229267 , n51503 , n229266 );
and ( n229268 , n229267 , n37123 );
not ( n51508 , n229267 );
and ( n51509 , n51508 , n37128 );
nor ( n51510 , n229268 , n51509 );
not ( n51511 , n51510 );
buf ( n51512 , n30803 );
not ( n51513 , n51512 );
not ( n229275 , n45468 );
or ( n229276 , n51513 , n229275 );
not ( n51516 , n51512 );
not ( n51517 , n45465 );
nand ( n51518 , n51516 , n51517 );
nand ( n51519 , n229276 , n51518 );
not ( n229281 , n38912 );
buf ( n229282 , n229281 );
and ( n51522 , n51519 , n229282 );
not ( n51523 , n51519 );
and ( n51524 , n51523 , n38912 );
nor ( n51525 , n51522 , n51524 );
nand ( n229287 , n51511 , n51525 );
not ( n229288 , n229287 );
or ( n51528 , n51501 , n229288 );
or ( n51529 , n229287 , n36259 );
nand ( n51530 , n51528 , n51529 );
not ( n51531 , n51530 );
or ( n229293 , n51500 , n51531 );
or ( n229294 , n51530 , n51499 );
nand ( n51534 , n229293 , n229294 );
buf ( n51535 , n51534 );
not ( n51536 , n51535 );
and ( n51537 , n51476 , n51536 );
and ( n229299 , n51475 , n51535 );
nor ( n229300 , n51537 , n229299 );
not ( n51540 , n229300 );
or ( n51541 , n51415 , n51540 );
not ( n51542 , n229175 );
not ( n51543 , n51534 );
not ( n229305 , n51543 );
not ( n229306 , n229235 );
or ( n51546 , n229305 , n229306 );
not ( n51547 , n229235 );
nand ( n51548 , n51547 , n51534 );
nand ( n51549 , n51546 , n51548 );
nand ( n229311 , n51542 , n51549 );
nand ( n229312 , n51541 , n229311 );
nand ( n51552 , n224248 , n46491 );
not ( n51553 , n51552 );
not ( n51554 , n36667 );
and ( n229316 , n51553 , n51554 );
not ( n229317 , n45857 );
nand ( n229318 , n229317 , n224248 );
and ( n229319 , n229318 , n36667 );
nor ( n51559 , n229316 , n229319 );
xnor ( n51560 , n45760 , n51559 );
not ( n51561 , n51560 );
not ( n51562 , n223562 );
not ( n51563 , n46448 );
nand ( n51564 , n51562 , n51563 );
not ( n229326 , n51564 );
not ( n229327 , n36540 );
and ( n51567 , n229326 , n229327 );
not ( n51568 , n46448 );
nand ( n51569 , n51568 , n51562 );
and ( n51570 , n51569 , n36540 );
nor ( n51571 , n51567 , n51570 );
not ( n51572 , n51571 );
nand ( n51573 , n46461 , n224225 );
and ( n51574 , n51573 , n36478 );
not ( n51575 , n51573 );
and ( n229337 , n51575 , n36479 );
nor ( n229338 , n51574 , n229337 );
not ( n229339 , n229338 );
or ( n229340 , n51572 , n229339 );
or ( n51580 , n229338 , n51571 );
nand ( n51581 , n229340 , n51580 );
nand ( n51582 , n46431 , n45777 );
and ( n51583 , n51582 , n36382 );
not ( n51584 , n51582 );
and ( n51585 , n51584 , n36383 );
nor ( n229347 , n51583 , n51585 );
and ( n229348 , n51581 , n229347 );
not ( n51588 , n51581 );
not ( n51589 , n229347 );
and ( n51590 , n51588 , n51589 );
nor ( n51591 , n229348 , n51590 );
not ( n51592 , n51591 );
or ( n51593 , n51561 , n51592 );
not ( n229355 , n51591 );
not ( n229356 , n51560 );
nand ( n51596 , n229355 , n229356 );
nand ( n51597 , n51593 , n51596 );
buf ( n51598 , n51597 );
and ( n51599 , n229312 , n51598 );
not ( n229361 , n229312 );
not ( n229362 , n51591 );
not ( n51602 , n229362 );
not ( n229364 , n229356 );
and ( n229365 , n51602 , n229364 );
and ( n51605 , n229362 , n229356 );
nor ( n51606 , n229365 , n51605 );
buf ( n51607 , n51606 );
and ( n51608 , n229361 , n51607 );
nor ( n229370 , n51599 , n51608 );
xor ( n229371 , n37178 , n37184 );
xnor ( n51611 , n229371 , n37191 );
xor ( n51612 , n33847 , n51611 );
xnor ( n51613 , n51612 , n38805 );
nand ( n51614 , n51613 , n208212 );
not ( n229376 , n51614 );
not ( n229377 , n28888 );
not ( n51617 , n43672 );
or ( n51618 , n229377 , n51617 );
not ( n51619 , n28888 );
nand ( n51620 , n51619 , n40861 );
nand ( n51621 , n51618 , n51620 );
and ( n51622 , n51621 , n218656 );
not ( n229384 , n51621 );
and ( n229385 , n229384 , n220953 );
nor ( n51625 , n51622 , n229385 );
not ( n229387 , n51625 );
not ( n229388 , n229387 );
and ( n51628 , n229376 , n229388 );
and ( n229390 , n51614 , n229387 );
nor ( n229391 , n51628 , n229390 );
not ( n51631 , n229391 );
not ( n229393 , n51631 );
not ( n229394 , n51613 );
nand ( n51634 , n51625 , n229394 );
not ( n51635 , n51634 );
not ( n51636 , n30287 );
and ( n51637 , n51635 , n51636 );
and ( n51638 , n51634 , n30287 );
nor ( n51639 , n51637 , n51638 );
not ( n229401 , n38514 );
not ( n229402 , n40156 );
xor ( n51642 , n38540 , n38557 );
not ( n229404 , n38548 );
xnor ( n229405 , n51642 , n229404 );
not ( n51645 , n229405 );
or ( n51646 , n229402 , n51645 );
or ( n51647 , n229405 , n40156 );
nand ( n51648 , n51646 , n51647 );
not ( n51649 , n51648 );
and ( n229411 , n229401 , n51649 );
and ( n229412 , n38514 , n51648 );
nor ( n51652 , n229411 , n229412 );
not ( n51653 , n225593 );
not ( n51654 , n26363 );
and ( n51655 , n51653 , n51654 );
and ( n51656 , n225593 , n26363 );
nor ( n229418 , n51655 , n51656 );
and ( n229419 , n229418 , n41055 );
not ( n51659 , n229418 );
and ( n229421 , n51659 , n45696 );
nor ( n229422 , n229419 , n229421 );
nand ( n51662 , n51652 , n229422 );
buf ( n51663 , n30222 );
xnor ( n51664 , n51662 , n51663 );
xor ( n51665 , n51639 , n51664 );
not ( n51666 , n208370 );
not ( n229428 , n51666 );
not ( n229429 , n204490 );
not ( n51669 , n25927 );
or ( n51670 , n229429 , n51669 );
nand ( n51671 , n47216 , n204487 );
nand ( n51672 , n51670 , n51671 );
and ( n229434 , n51672 , n25978 );
not ( n229435 , n51672 );
and ( n51675 , n229435 , n25965 );
nor ( n229437 , n229434 , n51675 );
buf ( n229438 , n40807 );
not ( n51678 , n229438 );
not ( n51679 , n37297 );
or ( n229441 , n51678 , n51679 );
not ( n229442 , n229438 );
nand ( n51682 , n229442 , n37296 );
nand ( n51683 , n229441 , n51682 );
and ( n51684 , n51683 , n31515 );
not ( n51685 , n51683 );
and ( n51686 , n51685 , n31528 );
nor ( n51687 , n51684 , n51686 );
nor ( n51688 , n229437 , n51687 );
not ( n51689 , n51688 );
and ( n229451 , n229428 , n51689 );
and ( n229452 , n51666 , n51688 );
nor ( n51692 , n229451 , n229452 );
xnor ( n51693 , n51665 , n51692 );
not ( n51694 , n39908 );
not ( n51695 , n38140 );
or ( n229457 , n51694 , n51695 );
or ( n229458 , n221827 , n39908 );
nand ( n51698 , n229457 , n229458 );
and ( n51699 , n51698 , n25684 );
not ( n51700 , n51698 );
and ( n51701 , n51700 , n25683 );
nor ( n229463 , n51699 , n51701 );
buf ( n229464 , n26003 );
nor ( n51704 , n43274 , n229464 );
not ( n229466 , n51704 );
nand ( n229467 , n229464 , n33937 );
nand ( n51707 , n229466 , n229467 );
and ( n51708 , n51707 , n43279 );
not ( n51709 , n51707 );
and ( n51710 , n51709 , n41082 );
nor ( n229472 , n51708 , n51710 );
nand ( n229473 , n229463 , n229472 );
and ( n51713 , n229473 , n208710 );
not ( n51714 , n229473 );
not ( n51715 , n208710 );
and ( n51716 , n51714 , n51715 );
or ( n229478 , n51713 , n51716 );
not ( n229479 , n229478 );
not ( n51719 , n29045 );
xor ( n229481 , n205781 , n204453 );
xnor ( n229482 , n229481 , n28029 );
nor ( n51722 , n51719 , n229482 );
not ( n51723 , n51722 );
not ( n51724 , n29045 );
nand ( n51725 , n51724 , n229482 );
nand ( n229487 , n51723 , n51725 );
and ( n229488 , n229487 , n205766 );
not ( n51728 , n229487 );
and ( n51729 , n51728 , n36568 );
nor ( n51730 , n229488 , n51729 );
nand ( n51731 , n29992 , n51730 );
not ( n229493 , n51731 );
not ( n229494 , n30040 );
and ( n51734 , n229493 , n229494 );
and ( n51735 , n51731 , n30040 );
nor ( n51736 , n51734 , n51735 );
not ( n51737 , n51736 );
or ( n229499 , n229479 , n51737 );
not ( n229500 , n229478 );
not ( n51740 , n51736 );
nand ( n51741 , n229500 , n51740 );
nand ( n51742 , n229499 , n51741 );
and ( n51743 , n51693 , n51742 );
not ( n229505 , n51693 );
not ( n229506 , n51742 );
and ( n51746 , n229505 , n229506 );
nor ( n51747 , n51743 , n51746 );
not ( n51748 , n51747 );
or ( n51749 , n229393 , n51748 );
or ( n51750 , n51747 , n51631 );
nand ( n229512 , n51749 , n51750 );
not ( n229513 , n204544 );
not ( n51753 , n229513 );
and ( n51754 , n229512 , n51753 );
not ( n51755 , n229512 );
not ( n51756 , n204553 );
not ( n229518 , n51756 );
and ( n229519 , n51755 , n229518 );
nor ( n51759 , n51754 , n229519 );
nand ( n229521 , n229370 , n51759 );
buf ( n229522 , n204722 );
not ( n51762 , n229522 );
not ( n229524 , n51762 );
not ( n229525 , n28721 );
or ( n51765 , n229524 , n229525 );
nand ( n51766 , n28722 , n229522 );
nand ( n51767 , n51765 , n51766 );
and ( n51768 , n51767 , n50070 );
not ( n51769 , n51767 );
and ( n229531 , n51769 , n227830 );
nor ( n229532 , n51768 , n229531 );
not ( n51772 , n33614 );
not ( n51773 , n32119 );
not ( n51774 , n29854 );
or ( n51775 , n51773 , n51774 );
or ( n229537 , n29854 , n32119 );
nand ( n229538 , n51775 , n229537 );
not ( n51778 , n229538 );
or ( n229540 , n51772 , n51778 );
or ( n229541 , n229538 , n33614 );
nand ( n51781 , n229540 , n229541 );
not ( n51782 , n51781 );
nand ( n51783 , n229532 , n51782 );
not ( n51784 , n31640 );
not ( n51785 , n34643 );
or ( n229547 , n51784 , n51785 );
or ( n229548 , n34643 , n31640 );
nand ( n51788 , n229547 , n229548 );
and ( n51789 , n51788 , n42372 );
not ( n229551 , n51788 );
and ( n229552 , n229551 , n50825 );
nor ( n51792 , n51789 , n229552 );
and ( n51793 , n51783 , n51792 );
not ( n51794 , n51783 );
not ( n51795 , n51792 );
and ( n51796 , n51794 , n51795 );
nor ( n51797 , n51793 , n51796 );
buf ( n229559 , n51797 );
not ( n229560 , n229559 );
not ( n51800 , n32740 );
not ( n51801 , n35782 );
or ( n51802 , n51800 , n51801 );
or ( n51803 , n35782 , n32740 );
nand ( n51804 , n51802 , n51803 );
not ( n51805 , n51804 );
not ( n51806 , n35774 );
not ( n51807 , n51806 );
or ( n229569 , n51805 , n51807 );
not ( n229570 , n35774 );
or ( n51810 , n229570 , n51804 );
nand ( n51811 , n229569 , n51810 );
and ( n51812 , n51811 , n35753 );
not ( n51813 , n51811 );
and ( n51814 , n51813 , n31008 );
nor ( n51815 , n51812 , n51814 );
not ( n229577 , n51815 );
not ( n229578 , n32240 );
not ( n51818 , n36936 );
not ( n51819 , n32214 );
or ( n51820 , n51818 , n51819 );
not ( n51821 , n32214 );
nand ( n229583 , n51821 , n36940 );
nand ( n229584 , n51820 , n229583 );
buf ( n51824 , n32206 );
xnor ( n51825 , n229584 , n51824 );
not ( n51826 , n51825 );
and ( n51827 , n229578 , n51826 );
and ( n229589 , n32240 , n51825 );
nor ( n229590 , n51827 , n229589 );
not ( n51830 , n30442 );
and ( n51831 , n205402 , n41227 );
not ( n51832 , n205402 );
not ( n51833 , n41227 );
and ( n229595 , n51832 , n51833 );
nor ( n229596 , n51831 , n229595 );
not ( n51836 , n229596 );
or ( n229598 , n51830 , n51836 );
or ( n229599 , n229596 , n37303 );
nand ( n51839 , n229598 , n229599 );
nand ( n51840 , n229590 , n51839 );
not ( n51841 , n51840 );
or ( n229603 , n229577 , n51841 );
or ( n229604 , n51840 , n51815 );
nand ( n51844 , n229603 , n229604 );
not ( n51845 , n51844 );
not ( n51846 , n51845 );
not ( n51847 , n29174 );
not ( n229609 , n26022 );
and ( n229610 , n51847 , n229609 );
and ( n51850 , n29174 , n26022 );
nor ( n51851 , n229610 , n51850 );
and ( n51852 , n51851 , n33936 );
not ( n51853 , n51851 );
and ( n51854 , n51853 , n33937 );
nor ( n51855 , n51852 , n51854 );
not ( n229617 , n30848 );
xor ( n229618 , n35891 , n229617 );
xnor ( n51858 , n229618 , n30889 );
nand ( n51859 , n51855 , n51858 );
not ( n51860 , n51859 );
and ( n51861 , n38446 , n29488 );
not ( n229623 , n38446 );
and ( n229624 , n229623 , n29492 );
nor ( n51864 , n51861 , n229624 );
not ( n51865 , n51864 );
not ( n51866 , n51865 );
not ( n51867 , n38460 );
not ( n229629 , n51867 );
or ( n229630 , n51866 , n229629 );
nand ( n51870 , n38460 , n51864 );
nand ( n229632 , n229630 , n51870 );
and ( n229633 , n229632 , n225200 );
not ( n51873 , n229632 );
and ( n51874 , n51873 , n38435 );
nor ( n51875 , n229633 , n51874 );
not ( n51876 , n51875 );
and ( n229638 , n51860 , n51876 );
and ( n229639 , n51859 , n51875 );
nor ( n51879 , n229638 , n229639 );
not ( n51880 , n51879 );
not ( n51881 , n51880 );
or ( n51882 , n51846 , n51881 );
nand ( n51883 , n51879 , n51844 );
nand ( n51884 , n51882 , n51883 );
nand ( n51885 , n51792 , n51781 );
not ( n51886 , n25443 );
not ( n229648 , n41113 );
or ( n229649 , n51886 , n229648 );
not ( n51889 , n25443 );
nand ( n51890 , n51889 , n42057 );
nand ( n51891 , n229649 , n51890 );
and ( n51892 , n51891 , n37946 );
not ( n229654 , n51891 );
and ( n229655 , n229654 , n227903 );
nor ( n51895 , n51892 , n229655 );
and ( n51896 , n51885 , n51895 );
not ( n51897 , n51885 );
not ( n51898 , n51895 );
and ( n229660 , n51897 , n51898 );
nor ( n229661 , n51896 , n229660 );
not ( n51901 , n229661 );
and ( n51902 , n51884 , n51901 );
not ( n51903 , n51884 );
and ( n51904 , n51903 , n229661 );
nor ( n51905 , n51902 , n51904 );
not ( n51906 , n44915 );
not ( n51907 , n32652 );
or ( n51908 , n51906 , n51907 );
not ( n229670 , n44915 );
nand ( n229671 , n229670 , n32651 );
nand ( n51911 , n51908 , n229671 );
not ( n229673 , n51911 );
not ( n51913 , n39417 );
and ( n51914 , n229673 , n51913 );
and ( n51915 , n32689 , n51911 );
nor ( n51916 , n51914 , n51915 );
not ( n229678 , n51916 );
not ( n229679 , n229678 );
not ( n51919 , n205256 );
not ( n51920 , n31777 );
or ( n51921 , n51919 , n51920 );
not ( n51922 , n205256 );
nand ( n229684 , n51922 , n33684 );
nand ( n229685 , n51921 , n229684 );
and ( n51925 , n229685 , n46734 );
not ( n51926 , n229685 );
and ( n51927 , n51926 , n46731 );
nor ( n51928 , n51925 , n51927 );
not ( n51929 , n26212 );
not ( n51930 , n48779 );
or ( n229692 , n51929 , n51930 );
or ( n229693 , n33565 , n26212 );
nand ( n51933 , n229692 , n229693 );
not ( n51934 , n51933 );
not ( n51935 , n36625 );
not ( n51936 , n51935 );
not ( n229698 , n51936 );
and ( n229699 , n51934 , n229698 );
and ( n51939 , n51933 , n51936 );
nor ( n51940 , n229699 , n51939 );
nand ( n51941 , n51928 , n51940 );
not ( n51942 , n51941 );
or ( n229704 , n229679 , n51942 );
or ( n229705 , n51941 , n229678 );
nand ( n51945 , n229704 , n229705 );
not ( n51946 , n51945 );
not ( n51947 , n51946 );
not ( n51948 , n41121 );
not ( n229710 , n205434 );
or ( n229711 , n51948 , n229710 );
not ( n51951 , n204279 );
not ( n229713 , n204306 );
or ( n229714 , n51951 , n229713 );
nand ( n51954 , n229714 , n205433 );
not ( n51955 , n51954 );
nand ( n51956 , n51955 , n41117 );
nand ( n51957 , n229711 , n51956 );
and ( n51958 , n51957 , n42174 );
not ( n229720 , n51957 );
not ( n229721 , n42174 );
and ( n51961 , n229720 , n229721 );
nor ( n51962 , n51958 , n51961 );
not ( n51963 , n41405 );
not ( n51964 , n25355 );
not ( n229726 , n45849 );
or ( n229727 , n51964 , n229726 );
or ( n51967 , n45849 , n25355 );
nand ( n51968 , n229727 , n51967 );
not ( n51969 , n51968 );
or ( n51970 , n51963 , n51969 );
or ( n51971 , n45531 , n51968 );
nand ( n51972 , n51970 , n51971 );
nand ( n229734 , n51962 , n51972 );
not ( n229735 , n229734 );
not ( n51975 , n35681 );
not ( n51976 , n39968 );
or ( n51977 , n51975 , n51976 );
not ( n51978 , n35681 );
nand ( n229740 , n51978 , n39974 );
nand ( n229741 , n51977 , n229740 );
and ( n51981 , n229741 , n48698 );
not ( n229743 , n229741 );
and ( n229744 , n229743 , n40007 );
nor ( n51984 , n51981 , n229744 );
not ( n229746 , n51984 );
and ( n229747 , n229735 , n229746 );
and ( n51987 , n229734 , n51984 );
nor ( n229749 , n229747 , n51987 );
not ( n51989 , n229749 );
not ( n51990 , n51989 );
or ( n51991 , n51947 , n51990 );
nand ( n51992 , n229749 , n51945 );
nand ( n229754 , n51991 , n51992 );
and ( n229755 , n51905 , n229754 );
not ( n51995 , n51905 );
not ( n51996 , n229754 );
and ( n51997 , n51995 , n51996 );
nor ( n51998 , n229755 , n51997 );
not ( n51999 , n51998 );
or ( n52000 , n229560 , n51999 );
xor ( n229762 , n229661 , n51884 );
xnor ( n229763 , n229762 , n229754 );
or ( n52003 , n229763 , n229559 );
nand ( n229765 , n52000 , n52003 );
not ( n229766 , n40393 );
not ( n52006 , n29518 );
or ( n52007 , n229766 , n52006 );
not ( n52008 , n40393 );
nand ( n52009 , n52008 , n207285 );
nand ( n229771 , n52007 , n52009 );
not ( n229772 , n229771 );
not ( n52012 , n29563 );
and ( n52013 , n229772 , n52012 );
and ( n52014 , n229771 , n29563 );
nor ( n52015 , n52013 , n52014 );
not ( n229777 , n52015 );
not ( n229778 , n229777 );
not ( n52018 , n45531 );
not ( n52019 , n25384 );
not ( n52020 , n45849 );
or ( n52021 , n52019 , n52020 );
not ( n229783 , n25384 );
nand ( n229784 , n229783 , n45524 );
nand ( n52024 , n52021 , n229784 );
not ( n52025 , n52024 );
or ( n52026 , n52018 , n52025 );
or ( n52027 , n45531 , n52024 );
nand ( n52028 , n52026 , n52027 );
not ( n52029 , n32987 );
not ( n229791 , n29909 );
not ( n229792 , n229791 );
or ( n52032 , n52029 , n229792 );
not ( n52033 , n32987 );
nand ( n52034 , n52033 , n29909 );
nand ( n52035 , n52032 , n52034 );
and ( n229797 , n52035 , n207706 );
not ( n229798 , n52035 );
and ( n52038 , n229798 , n29948 );
nor ( n52039 , n229797 , n52038 );
nand ( n52040 , n52028 , n52039 );
not ( n52041 , n52040 );
or ( n52042 , n229778 , n52041 );
or ( n52043 , n52040 , n229777 );
nand ( n229805 , n52042 , n52043 );
not ( n229806 , n229805 );
buf ( n52046 , n34728 );
not ( n52047 , n52046 );
not ( n52048 , n204858 );
or ( n52049 , n52047 , n52048 );
or ( n52050 , n204858 , n52046 );
nand ( n52051 , n52049 , n52050 );
and ( n52052 , n52051 , n204891 );
not ( n52053 , n52051 );
and ( n52054 , n52053 , n48593 );
nor ( n229816 , n52052 , n52054 );
not ( n229817 , n28140 );
not ( n52057 , n36967 );
or ( n52058 , n229817 , n52057 );
not ( n52059 , RI17337cf0_2169);
nand ( n52060 , n36943 , n52059 );
nand ( n229822 , n52058 , n52060 );
not ( n229823 , n229822 );
buf ( n52063 , n36963 );
not ( n52064 , n52063 );
or ( n52065 , n229823 , n52064 );
or ( n52066 , n52063 , n229822 );
nand ( n229828 , n52065 , n52066 );
and ( n229829 , n229828 , n223711 );
not ( n52069 , n229828 );
buf ( n52070 , n36934 );
and ( n52071 , n52069 , n52070 );
nor ( n52072 , n229829 , n52071 );
nand ( n52073 , n229816 , n52072 );
not ( n52074 , n52073 );
not ( n229836 , n204703 );
not ( n229837 , n28717 );
or ( n52077 , n229836 , n229837 );
or ( n229839 , n28717 , n204703 );
nand ( n229840 , n52077 , n229839 );
and ( n52080 , n229840 , n227830 );
not ( n52081 , n229840 );
and ( n52082 , n52081 , n26366 );
nor ( n52083 , n52080 , n52082 );
not ( n52084 , n52083 );
not ( n229846 , n52084 );
and ( n229847 , n52074 , n229846 );
and ( n52087 , n52073 , n52084 );
nor ( n52088 , n229847 , n52087 );
not ( n52089 , n52088 );
or ( n52090 , n229806 , n52089 );
or ( n229852 , n52088 , n229805 );
nand ( n229853 , n52090 , n229852 );
not ( n52093 , n33647 );
not ( n52094 , n204257 );
not ( n52095 , n52094 );
or ( n52096 , n52093 , n52095 );
not ( n52097 , n33647 );
nand ( n52098 , n52097 , n204257 );
nand ( n229860 , n52096 , n52098 );
xnor ( n229861 , n229860 , n32136 );
not ( n52101 , n229861 );
not ( n52102 , n35921 );
not ( n52103 , n208610 );
not ( n52104 , n52103 );
or ( n229866 , n52102 , n52104 );
not ( n229867 , n35921 );
nand ( n52107 , n229867 , n208610 );
nand ( n229869 , n229866 , n52107 );
and ( n229870 , n229869 , n229250 );
not ( n52110 , n229869 );
and ( n52111 , n52110 , n51492 );
nor ( n52112 , n229870 , n52111 );
not ( n52113 , n52112 );
nand ( n52114 , n52101 , n52113 );
not ( n52115 , n52114 );
not ( n229877 , n28951 );
not ( n229878 , n30320 );
or ( n52118 , n229877 , n229878 );
or ( n52119 , n30320 , n28951 );
nand ( n52120 , n52118 , n52119 );
and ( n52121 , n52120 , n204436 );
not ( n229883 , n52120 );
and ( n229884 , n229883 , n226279 );
nor ( n52124 , n52121 , n229884 );
not ( n52125 , n52124 );
not ( n52126 , n52125 );
and ( n52127 , n52115 , n52126 );
and ( n52128 , n52114 , n52125 );
nor ( n52129 , n52127 , n52128 );
and ( n229891 , n229853 , n52129 );
not ( n229892 , n229853 );
not ( n52132 , n52129 );
and ( n52133 , n229892 , n52132 );
nor ( n52134 , n229891 , n52133 );
buf ( n52135 , n209886 );
not ( n52136 , n52135 );
not ( n52137 , n52136 );
not ( n229899 , n38396 );
or ( n229900 , n52137 , n229899 );
nand ( n52140 , n38386 , n52135 );
nand ( n52141 , n229900 , n52140 );
and ( n52142 , n52141 , n33614 );
not ( n52143 , n52141 );
and ( n229905 , n52143 , n33619 );
nor ( n229906 , n52142 , n229905 );
buf ( n52146 , n32431 );
not ( n52147 , n52146 );
not ( n52148 , n52147 );
not ( n52149 , n40177 );
or ( n229911 , n52148 , n52149 );
nand ( n229912 , n222413 , n52146 );
nand ( n52152 , n229911 , n229912 );
and ( n229914 , n52152 , n33566 );
not ( n229915 , n52152 );
and ( n52155 , n229915 , n33567 );
nor ( n52156 , n229914 , n52155 );
not ( n52157 , n52156 );
nand ( n52158 , n229906 , n52157 );
not ( n229920 , n52158 );
xor ( n229921 , n34240 , n40743 );
xnor ( n52161 , n229921 , n207535 );
not ( n229923 , n52161 );
not ( n229924 , n229923 );
or ( n52164 , n229920 , n229924 );
or ( n52165 , n229923 , n52158 );
nand ( n52166 , n52164 , n52165 );
not ( n52167 , n52166 );
buf ( n229929 , n25912 );
not ( n229930 , n229929 );
not ( n52170 , n36255 );
or ( n52171 , n229930 , n52170 );
or ( n52172 , n36255 , n229929 );
nand ( n52173 , n52171 , n52172 );
and ( n229935 , n52173 , n32011 );
not ( n229936 , n52173 );
and ( n52176 , n229936 , n35624 );
nor ( n229938 , n229935 , n52176 );
not ( n229939 , n229938 );
not ( n52179 , RI174a7fd0_917);
and ( n52180 , n25624 , n52179 );
not ( n52181 , n25624 );
and ( n52182 , n52181 , n25620 );
or ( n52183 , n52180 , n52182 );
not ( n52184 , n52183 );
not ( n52185 , n37619 );
not ( n52186 , n52185 );
or ( n52187 , n52184 , n52186 );
or ( n52188 , n52185 , n52183 );
nand ( n229950 , n52187 , n52188 );
not ( n229951 , n229950 );
not ( n52191 , n37652 );
and ( n52192 , n229951 , n52191 );
and ( n52193 , n229950 , n37652 );
nor ( n52194 , n52192 , n52193 );
nand ( n229956 , n229939 , n52194 );
not ( n229957 , n229956 );
not ( n52197 , n35504 );
not ( n52198 , n33957 );
or ( n52199 , n52197 , n52198 );
not ( n52200 , n35504 );
nand ( n52201 , n52200 , n33954 );
nand ( n52202 , n52199 , n52201 );
not ( n229964 , n52202 );
not ( n229965 , n31344 );
and ( n229966 , n229964 , n229965 );
and ( n229967 , n52202 , n31344 );
nor ( n52207 , n229966 , n229967 );
not ( n52208 , n52207 );
not ( n52209 , n52208 );
and ( n52210 , n229957 , n52209 );
and ( n52211 , n229956 , n52208 );
nor ( n52212 , n52210 , n52211 );
not ( n229974 , n52212 );
and ( n229975 , n52167 , n229974 );
and ( n52215 , n52166 , n52212 );
nor ( n52216 , n229975 , n52215 );
not ( n52217 , n52216 );
and ( n52218 , n52134 , n52217 );
not ( n229980 , n52134 );
and ( n229981 , n229980 , n52216 );
nor ( n52221 , n52218 , n229981 );
not ( n52222 , n52221 );
not ( n52223 , n52222 );
and ( n52224 , n229765 , n52223 );
not ( n52225 , n229765 );
and ( n52226 , n52134 , n52216 );
not ( n52227 , n52134 );
and ( n52228 , n52227 , n52217 );
nor ( n52229 , n52226 , n52228 );
buf ( n229991 , n52229 );
and ( n229992 , n52225 , n229991 );
nor ( n52232 , n52224 , n229992 );
not ( n52233 , n52232 );
and ( n52234 , n229521 , n52233 );
not ( n52235 , n229521 );
and ( n229997 , n52235 , n52232 );
nor ( n229998 , n52234 , n229997 );
or ( n52238 , n229998 , n49959 );
nand ( n52239 , n51383 , n52238 );
buf ( n52240 , n52239 );
nand ( n52241 , n45952 , n46630 );
and ( n230003 , n52241 , n46644 );
not ( n230004 , n52241 );
and ( n52244 , n230004 , n46643 );
nor ( n230006 , n230003 , n52244 );
not ( n230007 , n230006 );
not ( n52247 , n230007 );
not ( n52248 , n46716 );
or ( n52249 , n52247 , n52248 );
or ( n52250 , n46716 , n230007 );
nand ( n52251 , n52249 , n52250 );
not ( n52252 , n52251 );
not ( n52253 , n204559 );
not ( n52254 , n39671 );
or ( n52255 , n52253 , n52254 );
not ( n52256 , n28381 );
or ( n230018 , n52256 , n204559 );
nand ( n230019 , n52255 , n230018 );
and ( n52259 , n230019 , n30140 );
not ( n52260 , n230019 );
and ( n52261 , n52260 , n39679 );
nor ( n52262 , n52259 , n52261 );
not ( n230024 , n33537 );
not ( n230025 , n35357 );
or ( n52265 , n230024 , n230025 );
or ( n52266 , n35357 , n33537 );
nand ( n52267 , n52265 , n52266 );
not ( n52268 , n52267 );
not ( n52269 , n35390 );
or ( n230031 , n52268 , n52269 );
or ( n230032 , n35390 , n52267 );
nand ( n52272 , n230031 , n230032 );
not ( n52273 , n52272 );
nand ( n52274 , n52262 , n52273 );
buf ( n52275 , n33167 );
not ( n230037 , n52275 );
not ( n230038 , n28251 );
or ( n52278 , n230037 , n230038 );
or ( n52279 , n28251 , n52275 );
nand ( n52280 , n52278 , n52279 );
xnor ( n52281 , n52280 , n223793 );
xor ( n230043 , n52274 , n52281 );
not ( n230044 , n230043 );
not ( n52284 , n230044 );
not ( n52285 , n205875 );
not ( n52286 , n25426 );
or ( n52287 , n52285 , n52286 );
or ( n52288 , n25426 , n205875 );
nand ( n52289 , n52287 , n52288 );
and ( n230051 , n52289 , n28680 );
not ( n230052 , n52289 );
not ( n52292 , n28680 );
and ( n52293 , n230052 , n52292 );
nor ( n52294 , n230051 , n52293 );
not ( n52295 , n28725 );
and ( n230057 , n204691 , n206479 );
not ( n230058 , n204691 );
and ( n52298 , n230058 , n28721 );
nor ( n52299 , n230057 , n52298 );
not ( n52300 , n52299 );
or ( n52301 , n52295 , n52300 );
or ( n230063 , n52299 , n227830 );
nand ( n230064 , n52301 , n230063 );
nand ( n52304 , n52294 , n230064 );
not ( n52305 , n52304 );
xor ( n52306 , n34262 , n40743 );
xnor ( n52307 , n52306 , n49026 );
not ( n230069 , n52307 );
or ( n230070 , n52305 , n230069 );
nand ( n52310 , n52294 , n230064 );
or ( n52311 , n52307 , n52310 );
nand ( n230073 , n230070 , n52311 );
not ( n230074 , n230073 );
or ( n52314 , n52284 , n230074 );
or ( n52315 , n230073 , n230044 );
nand ( n52316 , n52314 , n52315 );
not ( n52317 , n52316 );
not ( n52318 , n39922 );
not ( n52319 , n30652 );
not ( n230081 , n40619 );
or ( n230082 , n52319 , n230081 );
or ( n52322 , n40619 , n30652 );
nand ( n52323 , n230082 , n52322 );
not ( n52324 , n52323 );
or ( n52325 , n52318 , n52324 );
or ( n52326 , n52323 , n39922 );
nand ( n230088 , n52325 , n52326 );
not ( n230089 , n230088 );
not ( n52329 , n32252 );
xor ( n52330 , n29543 , n29560 );
xnor ( n52331 , n52330 , n47434 );
not ( n52332 , n52331 );
not ( n230094 , n52332 );
or ( n230095 , n52329 , n230094 );
nand ( n52335 , n52331 , n32248 );
nand ( n52336 , n230095 , n52335 );
not ( n52337 , n52336 );
not ( n52338 , n37261 );
and ( n52339 , n52337 , n52338 );
not ( n52340 , n37260 );
and ( n230102 , n52340 , n52336 );
nor ( n230103 , n52339 , n230102 );
not ( n52343 , n230103 );
nand ( n52344 , n230089 , n52343 );
not ( n52345 , n52344 );
buf ( n52346 , n40129 );
not ( n52347 , n52346 );
not ( n52348 , n37991 );
or ( n52349 , n52347 , n52348 );
not ( n52350 , n52346 );
nand ( n230112 , n52350 , n37996 );
nand ( n230113 , n52349 , n230112 );
and ( n52353 , n230113 , n35482 );
not ( n52354 , n230113 );
and ( n52355 , n52354 , n38000 );
nor ( n52356 , n52353 , n52355 );
not ( n230118 , n52356 );
and ( n230119 , n52345 , n230118 );
and ( n52359 , n52344 , n52356 );
nor ( n52360 , n230119 , n52359 );
not ( n52361 , n52360 );
not ( n52362 , n40869 );
not ( n230124 , n220726 );
or ( n230125 , n52362 , n230124 );
not ( n52365 , n40869 );
nand ( n52366 , n52365 , n216417 );
nand ( n52367 , n230125 , n52366 );
and ( n52368 , n52367 , n31213 );
not ( n230130 , n52367 );
and ( n230131 , n230130 , n38677 );
nor ( n52371 , n52368 , n230131 );
not ( n52372 , n226349 );
xnor ( n52373 , n34145 , n47605 );
not ( n52374 , n52373 );
not ( n52375 , n52374 );
or ( n52376 , n52372 , n52375 );
nand ( n52377 , n52373 , n204858 );
nand ( n52378 , n52376 , n52377 );
nand ( n52379 , n52371 , n52378 );
not ( n230141 , n38449 );
not ( n230142 , n32174 );
or ( n230143 , n230141 , n230142 );
or ( n230144 , n32174 , n38449 );
nand ( n52384 , n230143 , n230144 );
not ( n52385 , n219851 );
and ( n52386 , n52384 , n52385 );
not ( n52387 , n52384 );
and ( n230149 , n52387 , n219851 );
nor ( n230150 , n52386 , n230149 );
buf ( n52390 , n230150 );
xor ( n230152 , n52379 , n52390 );
not ( n230153 , n230152 );
or ( n52393 , n52361 , n230153 );
or ( n230155 , n230152 , n52360 );
nand ( n230156 , n52393 , n230155 );
xor ( n52396 , n34525 , n45281 );
xnor ( n52397 , n52396 , n44136 );
not ( n52398 , n37346 );
not ( n52399 , n32223 );
and ( n230161 , n52398 , n52399 );
and ( n230162 , n37346 , n32223 );
nor ( n52402 , n230161 , n230162 );
and ( n52403 , n52402 , n37353 );
not ( n52404 , n52402 );
and ( n52405 , n52404 , n37356 );
nor ( n230167 , n52403 , n52405 );
not ( n230168 , n230167 );
nand ( n52408 , n52397 , n230168 );
not ( n52409 , n52408 );
not ( n52410 , n25457 );
not ( n52411 , n25977 );
buf ( n52412 , n41343 );
not ( n52413 , n52412 );
and ( n230175 , n52411 , n52413 );
and ( n230176 , n25977 , n52412 );
nor ( n52416 , n230175 , n230176 );
not ( n230178 , n52416 );
not ( n230179 , n230178 );
or ( n52419 , n52410 , n230179 );
nand ( n52420 , n52416 , n36982 );
nand ( n52421 , n52419 , n52420 );
not ( n52422 , n52421 );
and ( n230184 , n52409 , n52422 );
not ( n230185 , n230167 );
nand ( n52425 , n230185 , n52397 );
and ( n52426 , n52425 , n52421 );
nor ( n52427 , n230184 , n52426 );
and ( n52428 , n230156 , n52427 );
not ( n52429 , n230156 );
not ( n52430 , n52427 );
and ( n52431 , n52429 , n52430 );
nor ( n52432 , n52428 , n52431 );
not ( n52433 , n52432 );
or ( n230195 , n52317 , n52433 );
not ( n230196 , n52316 );
not ( n52436 , n52432 );
nand ( n230198 , n230196 , n52436 );
nand ( n230199 , n230195 , n230198 );
buf ( n52439 , n230199 );
not ( n230201 , n52439 );
not ( n230202 , n230201 );
and ( n52442 , n52252 , n230202 );
and ( n230204 , n52251 , n230201 );
nor ( n230205 , n52442 , n230204 );
buf ( n52445 , n43517 );
not ( n230207 , n52445 );
nand ( n230208 , n230205 , n230207 );
not ( n230209 , n35330 );
not ( n230210 , n29607 );
or ( n52450 , n230209 , n230210 );
or ( n52451 , n29607 , n35330 );
nand ( n52452 , n52450 , n52451 );
and ( n52453 , n52452 , n207407 );
not ( n230215 , n52452 );
and ( n230216 , n230215 , n29647 );
nor ( n52456 , n52453 , n230216 );
nand ( n52457 , n40068 , n52456 );
buf ( n52458 , n26193 );
not ( n52459 , n52458 );
not ( n230221 , n36618 );
or ( n230222 , n52459 , n230221 );
or ( n52462 , n36618 , n52458 );
nand ( n52463 , n230222 , n52462 );
and ( n52464 , n52463 , n48427 );
not ( n52465 , n52463 );
not ( n230227 , n225682 );
and ( n230228 , n52465 , n230227 );
nor ( n52468 , n52464 , n230228 );
buf ( n52469 , n52468 );
not ( n52470 , n52469 );
and ( n52471 , n52457 , n52470 );
not ( n230233 , n52457 );
and ( n230234 , n230233 , n52469 );
nor ( n52474 , n52471 , n230234 );
buf ( n230236 , n52474 );
not ( n230237 , n230236 );
not ( n52477 , n33455 );
buf ( n230239 , RI173e46e8_1642);
xor ( n230240 , n230239 , n32354 );
xor ( n52480 , n230240 , n32361 );
not ( n230242 , n52480 );
or ( n230243 , n52477 , n230242 );
or ( n52483 , n52480 , n33455 );
nand ( n52484 , n230243 , n52483 );
and ( n52485 , n52484 , n227444 );
not ( n52486 , n52484 );
not ( n230248 , n37297 );
and ( n230249 , n52486 , n230248 );
nor ( n52489 , n52485 , n230249 );
not ( n52490 , n52489 );
xor ( n52491 , n28899 , n40861 );
xnor ( n52492 , n52491 , n218655 );
not ( n230254 , n52492 );
nand ( n230255 , n52490 , n230254 );
not ( n52495 , n230255 );
buf ( n52496 , n39933 );
not ( n52497 , n52496 );
and ( n52498 , n52495 , n52497 );
not ( n230260 , n52492 );
nand ( n230261 , n230260 , n52490 );
and ( n52501 , n230261 , n52496 );
nor ( n52502 , n52498 , n52501 );
not ( n52503 , n52502 );
not ( n52504 , n37018 );
not ( n52505 , n41593 );
or ( n52506 , n52504 , n52505 );
not ( n230268 , n37018 );
nand ( n230269 , n230268 , n28188 );
nand ( n52509 , n52506 , n230269 );
not ( n230271 , n52509 );
not ( n230272 , n36093 );
and ( n52512 , n230271 , n230272 );
and ( n52513 , n52509 , n36093 );
nor ( n52514 , n52512 , n52513 );
not ( n52515 , n32323 );
not ( n52516 , n41498 );
not ( n52517 , n32284 );
or ( n230279 , n52516 , n52517 );
not ( n230280 , n32279 );
nand ( n52520 , n230280 , n41495 );
nand ( n52521 , n230279 , n52520 );
not ( n52522 , n52521 );
or ( n52523 , n52515 , n52522 );
not ( n230285 , n32326 );
or ( n230286 , n52521 , n230285 );
nand ( n52526 , n52523 , n230286 );
nand ( n230288 , n52514 , n52526 );
not ( n230289 , n230288 );
not ( n52529 , n40138 );
or ( n52530 , n230289 , n52529 );
or ( n52531 , n40138 , n230288 );
nand ( n52532 , n52530 , n52531 );
not ( n230294 , n52532 );
or ( n230295 , n52503 , n230294 );
or ( n52535 , n52532 , n52502 );
nand ( n52536 , n230295 , n52535 );
not ( n52537 , RI17538c00_591);
and ( n52538 , n52537 , n35629 );
nand ( n230300 , n204524 , n52538 , n204517 , n204525 );
not ( n230301 , n40090 );
xor ( n52541 , n230300 , n230301 );
not ( n52542 , n52456 );
nand ( n52543 , n52542 , n52470 );
xnor ( n230305 , n52541 , n52543 );
and ( n230306 , n52536 , n230305 );
not ( n230307 , n52536 );
not ( n230308 , n230305 );
and ( n52548 , n230307 , n230308 );
nor ( n52549 , n230306 , n52548 );
not ( n52550 , n39817 );
not ( n52551 , n30175 );
not ( n230313 , n27716 );
or ( n230314 , n52551 , n230313 );
or ( n52554 , n27716 , n30175 );
nand ( n52555 , n230314 , n52554 );
not ( n52556 , n52555 );
not ( n52557 , n27759 );
and ( n230319 , n52556 , n52557 );
and ( n230320 , n52555 , n27759 );
nor ( n52560 , n230319 , n230320 );
not ( n52561 , n52560 );
nand ( n52562 , n39788 , n52561 );
not ( n52563 , n52562 );
or ( n230325 , n52550 , n52563 );
or ( n230326 , n52562 , n39817 );
nand ( n52566 , n230325 , n230326 );
not ( n52567 , n52566 );
not ( n52568 , n52567 );
not ( n52569 , n28262 );
not ( n52570 , n48058 );
or ( n52571 , n52569 , n52570 );
or ( n230333 , n48058 , n28262 );
nand ( n230334 , n52571 , n230333 );
and ( n52574 , n230334 , n204586 );
not ( n52575 , n230334 );
and ( n52576 , n52575 , n34416 );
nor ( n52577 , n52574 , n52576 );
not ( n230339 , n52577 );
buf ( n230340 , n37557 );
not ( n52580 , n230340 );
not ( n52581 , n35291 );
or ( n52582 , n52580 , n52581 );
or ( n52583 , n35291 , n230340 );
nand ( n52584 , n52582 , n52583 );
not ( n52585 , n52584 );
not ( n230347 , n27968 );
or ( n230348 , n52585 , n230347 );
or ( n52588 , n27968 , n52584 );
nand ( n52589 , n230348 , n52588 );
not ( n52590 , n52589 );
nand ( n52591 , n230339 , n52590 );
not ( n230353 , n52591 );
not ( n230354 , n39859 );
and ( n52594 , n230353 , n230354 );
and ( n52595 , n52591 , n39859 );
nor ( n52596 , n52594 , n52595 );
not ( n52597 , n52596 );
not ( n52598 , n52597 );
or ( n52599 , n52568 , n52598 );
nand ( n230361 , n52596 , n52566 );
nand ( n230362 , n52599 , n230361 );
and ( n52602 , n52549 , n230362 );
not ( n52603 , n52549 );
not ( n52604 , n230362 );
and ( n52605 , n52603 , n52604 );
nor ( n230367 , n52602 , n52605 );
not ( n230368 , n230367 );
or ( n52608 , n230237 , n230368 );
not ( n52609 , n230236 );
and ( n52610 , n52549 , n52604 );
not ( n52611 , n52549 );
and ( n230373 , n52611 , n230362 );
nor ( n230374 , n52610 , n230373 );
nand ( n52614 , n52609 , n230374 );
nand ( n52615 , n52608 , n52614 );
not ( n52616 , n52615 );
not ( n52617 , n29608 );
not ( n52618 , n28522 );
not ( n230380 , n37406 );
or ( n230381 , n52618 , n230380 );
or ( n52621 , n37406 , n28522 );
nand ( n52622 , n230381 , n52621 );
not ( n52623 , n52622 );
or ( n52624 , n52617 , n52623 );
or ( n230386 , n52622 , n29608 );
nand ( n230387 , n52624 , n230386 );
not ( n52627 , n40813 );
not ( n52628 , n38538 );
not ( n52629 , n33474 );
or ( n52630 , n52628 , n52629 );
or ( n52631 , n33474 , n38538 );
nand ( n52632 , n52630 , n52631 );
not ( n230394 , n52632 );
and ( n230395 , n52627 , n230394 );
not ( n52635 , n43695 );
and ( n52636 , n52635 , n52632 );
nor ( n52637 , n230395 , n52636 );
nor ( n52638 , n230387 , n52637 );
and ( n52639 , n52638 , n40315 );
not ( n230401 , n52638 );
and ( n230402 , n230401 , n40316 );
nor ( n52642 , n52639 , n230402 );
not ( n52643 , n52642 );
xor ( n52644 , n204995 , n216262 );
not ( n52645 , n52644 );
not ( n230407 , n32082 );
or ( n230408 , n52645 , n230407 );
or ( n52648 , n32082 , n52644 );
nand ( n52649 , n230408 , n52648 );
not ( n52650 , n52649 );
not ( n52651 , n35866 );
not ( n230413 , n31008 );
or ( n230414 , n52651 , n230413 );
not ( n52654 , n35866 );
nand ( n230416 , n52654 , n35753 );
nand ( n230417 , n230414 , n230416 );
and ( n52657 , n230417 , n30972 );
not ( n52658 , n230417 );
and ( n52659 , n52658 , n50902 );
nor ( n52660 , n52657 , n52659 );
not ( n230422 , n52660 );
nand ( n230423 , n52650 , n230422 );
not ( n52663 , n40236 );
and ( n52664 , n230423 , n52663 );
not ( n52665 , n230423 );
and ( n52666 , n52665 , n40236 );
nor ( n230428 , n52664 , n52666 );
not ( n230429 , n230428 );
or ( n52669 , n52643 , n230429 );
or ( n52670 , n230428 , n52642 );
nand ( n52671 , n52669 , n52670 );
xor ( n52672 , n25649 , n52185 );
xnor ( n230434 , n52672 , n40969 );
not ( n230435 , n28613 );
xor ( n52675 , n30476 , n30484 );
xnor ( n230437 , n52675 , n30493 );
not ( n230438 , n230437 );
not ( n52678 , n230438 );
or ( n52679 , n230435 , n52678 );
or ( n52680 , n30495 , n28613 );
nand ( n52681 , n52679 , n52680 );
xnor ( n230443 , n52681 , n227018 );
buf ( n230444 , n230443 );
nand ( n52684 , n230434 , n230444 );
not ( n52685 , n52684 );
not ( n52686 , n40262 );
and ( n52687 , n52685 , n52686 );
and ( n230449 , n52684 , n40262 );
nor ( n230450 , n52687 , n230449 );
and ( n52690 , n52671 , n230450 );
not ( n230452 , n52671 );
not ( n230453 , n230450 );
and ( n52693 , n230452 , n230453 );
nor ( n230455 , n52690 , n52693 );
not ( n230456 , n40350 );
xor ( n52696 , n39227 , n45799 );
xnor ( n230458 , n52696 , n28405 );
not ( n230459 , n230458 );
not ( n52699 , n30153 );
not ( n230461 , n47261 );
or ( n230462 , n52699 , n230461 );
nand ( n52702 , n41359 , n30149 );
nand ( n52703 , n230462 , n52702 );
not ( n52704 , n27721 );
not ( n52705 , n52704 );
and ( n52706 , n52703 , n52705 );
not ( n230468 , n52703 );
and ( n230469 , n230468 , n27716 );
nor ( n52709 , n52706 , n230469 );
not ( n52710 , n52709 );
nand ( n52711 , n230459 , n52710 );
not ( n52712 , n52711 );
or ( n52713 , n230456 , n52712 );
not ( n52714 , n52709 );
nand ( n52715 , n52714 , n230459 );
or ( n230477 , n52715 , n40350 );
nand ( n230478 , n52713 , n230477 );
not ( n52718 , n230478 );
not ( n230480 , n42738 );
not ( n230481 , n35923 );
or ( n52721 , n230480 , n230481 );
nand ( n52722 , n42394 , n42734 );
nand ( n52723 , n52721 , n52722 );
and ( n52724 , n52723 , n41398 );
not ( n52725 , n52723 );
and ( n230487 , n52725 , n41395 );
nor ( n230488 , n52724 , n230487 );
not ( n52728 , n230488 );
not ( n52729 , n37326 );
not ( n52730 , n41756 );
or ( n52731 , n52729 , n52730 );
or ( n230493 , n227330 , n37326 );
nand ( n230494 , n52731 , n230493 );
and ( n52734 , n230494 , n228145 );
not ( n52735 , n230494 );
not ( n230497 , n228145 );
and ( n230498 , n52735 , n230497 );
nor ( n52738 , n52734 , n230498 );
not ( n52739 , n52738 );
nand ( n52740 , n52728 , n52739 );
not ( n52741 , n52740 );
not ( n52742 , n40428 );
not ( n230504 , n52742 );
not ( n230505 , n230504 );
and ( n52745 , n52741 , n230505 );
and ( n52746 , n52740 , n230504 );
nor ( n52747 , n52745 , n52746 );
not ( n52748 , n52747 );
and ( n52749 , n52718 , n52748 );
and ( n230511 , n230478 , n52747 );
nor ( n230512 , n52749 , n230511 );
not ( n52752 , n230512 );
and ( n52753 , n230455 , n52752 );
not ( n52754 , n230455 );
and ( n52755 , n52754 , n230512 );
nor ( n52756 , n52753 , n52755 );
buf ( n52757 , n52756 );
not ( n230519 , n52757 );
and ( n230520 , n52616 , n230519 );
and ( n52760 , n52615 , n52757 );
nor ( n52761 , n230520 , n52760 );
not ( n52762 , n25890 );
not ( n52763 , n31967 );
or ( n52764 , n52762 , n52763 );
or ( n52765 , n31967 , n25890 );
nand ( n52766 , n52764 , n52765 );
not ( n52767 , n52766 );
not ( n52768 , n32011 );
and ( n52769 , n52767 , n52768 );
and ( n52770 , n52766 , n32011 );
nor ( n52771 , n52769 , n52770 );
not ( n230533 , n52771 );
not ( n230534 , n230533 );
not ( n52774 , n39836 );
not ( n230536 , n38188 );
or ( n230537 , n52774 , n230536 );
not ( n52777 , n39836 );
nand ( n52778 , n52777 , n38201 );
nand ( n52779 , n230537 , n52778 );
and ( n52780 , n52779 , n29411 );
not ( n230542 , n52779 );
and ( n230543 , n230542 , n38205 );
nor ( n52783 , n52780 , n230543 );
not ( n230545 , n204271 );
not ( n230546 , n36750 );
or ( n52786 , n230545 , n230546 );
or ( n52787 , n36750 , n204271 );
nand ( n52788 , n52786 , n52787 );
and ( n52789 , n52788 , n44035 );
not ( n230551 , n52788 );
not ( n230552 , n30405 );
and ( n52792 , n230551 , n230552 );
nor ( n52793 , n52789 , n52792 );
nand ( n52794 , n52783 , n52793 );
not ( n52795 , n52794 );
or ( n230557 , n230534 , n52795 );
or ( n230558 , n52794 , n230533 );
nand ( n52798 , n230557 , n230558 );
not ( n52799 , n52798 );
not ( n52800 , n30467 );
not ( n52801 , n41448 );
or ( n230563 , n52800 , n52801 );
or ( n230564 , n46596 , n30467 );
nand ( n52804 , n230563 , n230564 );
buf ( n52805 , n33229 );
not ( n52806 , n52805 );
and ( n52807 , n52804 , n52806 );
not ( n52808 , n52804 );
and ( n52809 , n52808 , n52805 );
nor ( n230571 , n52807 , n52809 );
not ( n230572 , n230571 );
not ( n52812 , n207407 );
not ( n230574 , n35371 );
and ( n230575 , n52812 , n230574 );
and ( n52815 , n46664 , n35371 );
nor ( n52816 , n230575 , n52815 );
and ( n52817 , n52816 , n46668 );
not ( n52818 , n52816 );
and ( n52819 , n52818 , n46671 );
nor ( n52820 , n52817 , n52819 );
not ( n230582 , n52820 );
nand ( n230583 , n230572 , n230582 );
not ( n52823 , n44929 );
not ( n52824 , n32655 );
or ( n52825 , n52823 , n52824 );
or ( n52826 , n32655 , n44929 );
nand ( n230588 , n52825 , n52826 );
not ( n230589 , n230588 );
not ( n52829 , n230589 );
not ( n230591 , n32688 );
or ( n230592 , n52829 , n230591 );
nand ( n52832 , n39417 , n230588 );
nand ( n230594 , n230592 , n52832 );
not ( n230595 , n230594 );
and ( n52835 , n230583 , n230595 );
not ( n230597 , n230583 );
and ( n52837 , n230597 , n230594 );
nor ( n52838 , n52835 , n52837 );
not ( n52839 , n52838 );
not ( n52840 , n41150 );
not ( n230602 , n30359 );
not ( n230603 , n46746 );
or ( n52843 , n230602 , n230603 );
not ( n52844 , n30359 );
nand ( n52845 , n29335 , n52844 );
nand ( n52846 , n52843 , n52845 );
not ( n230608 , n52846 );
or ( n230609 , n52840 , n230608 );
or ( n52849 , n52846 , n46753 );
nand ( n52850 , n230609 , n52849 );
not ( n52851 , n52850 );
not ( n52852 , n28071 );
not ( n230614 , n36347 );
not ( n230615 , n28348 );
and ( n52855 , n230614 , n230615 );
and ( n230617 , n36347 , n28348 );
nor ( n230618 , n52855 , n230617 );
and ( n52858 , n52852 , n230618 );
not ( n52859 , n52852 );
not ( n52860 , n230618 );
and ( n52861 , n52859 , n52860 );
nor ( n230623 , n52858 , n52861 );
not ( n230624 , n230623 );
not ( n52864 , n33328 );
not ( n52865 , n39554 );
or ( n52866 , n52864 , n52865 );
not ( n52867 , n33328 );
nand ( n230629 , n52867 , n39553 );
nand ( n230630 , n52866 , n230629 );
and ( n52870 , n230630 , n39558 );
not ( n52871 , n230630 );
and ( n52872 , n52871 , n39559 );
nor ( n52873 , n52870 , n52872 );
nand ( n230635 , n230624 , n52873 );
not ( n230636 , n230635 );
or ( n52876 , n52851 , n230636 );
or ( n52877 , n230635 , n52850 );
nand ( n52878 , n52876 , n52877 );
not ( n52879 , n52878 );
not ( n52880 , n52793 );
nand ( n52881 , n52771 , n52880 );
not ( n230643 , n52881 );
xor ( n230644 , n31030 , n42023 );
not ( n52884 , n34913 );
xnor ( n52885 , n230644 , n52884 );
not ( n52886 , n52885 );
not ( n52887 , n52886 );
and ( n230649 , n230643 , n52887 );
and ( n230650 , n52881 , n52886 );
nor ( n52890 , n230649 , n230650 );
not ( n52891 , n52890 );
or ( n52892 , n52879 , n52891 );
or ( n52893 , n52890 , n52878 );
nand ( n52894 , n52892 , n52893 );
not ( n52895 , n52894 );
not ( n230657 , n52895 );
or ( n230658 , n52839 , n230657 );
not ( n52898 , n52838 );
nand ( n52899 , n52898 , n52894 );
nand ( n52900 , n230658 , n52899 );
not ( n52901 , n52900 );
buf ( n230663 , RI17400528_1506);
not ( n230664 , n230663 );
not ( n52904 , n30757 );
or ( n230666 , n230664 , n52904 );
nand ( n230667 , n30771 , n39695 );
nand ( n52907 , n230666 , n230667 );
and ( n230669 , n52907 , n40607 );
not ( n230670 , n52907 );
and ( n52910 , n230670 , n39481 );
nor ( n52911 , n230669 , n52910 );
not ( n52912 , n32580 );
not ( n230674 , n28502 );
or ( n230675 , n52912 , n230674 );
nand ( n52915 , n28508 , n32576 );
nand ( n52916 , n230675 , n52915 );
not ( n52917 , n52916 );
not ( n52918 , n44690 );
or ( n230680 , n52917 , n52918 );
or ( n230681 , n44690 , n52916 );
nand ( n52921 , n230680 , n230681 );
not ( n52922 , n52921 );
nand ( n52923 , n52911 , n52922 );
not ( n52924 , n52923 );
not ( n230686 , n27747 );
not ( n230687 , n25508 );
or ( n52927 , n230686 , n230687 );
or ( n230689 , n25508 , n27747 );
nand ( n230690 , n52927 , n230689 );
not ( n52930 , n230690 );
not ( n230692 , n37450 );
not ( n230693 , n230692 );
and ( n52933 , n52930 , n230693 );
and ( n52934 , n230690 , n230692 );
nor ( n52935 , n52933 , n52934 );
not ( n52936 , n52935 );
not ( n52937 , n52936 );
and ( n52938 , n52924 , n52937 );
and ( n230700 , n52923 , n52936 );
nor ( n230701 , n52938 , n230700 );
not ( n52941 , n230701 );
not ( n52942 , n52941 );
not ( n52943 , n42936 );
not ( n52944 , n43261 );
or ( n230706 , n52943 , n52944 );
or ( n230707 , n45799 , n42936 );
nand ( n52947 , n230706 , n230707 );
xor ( n52948 , n52947 , n45230 );
not ( n52949 , n52948 );
not ( n52950 , n38062 );
not ( n230712 , n30034 );
or ( n230713 , n52950 , n230712 );
not ( n52953 , n30038 );
nand ( n52954 , n52953 , n38058 );
nand ( n52955 , n230713 , n52954 );
not ( n52956 , n52955 );
not ( n230718 , n50452 );
not ( n230719 , n230718 );
and ( n52959 , n52956 , n230719 );
and ( n52960 , n52955 , n230718 );
nor ( n52961 , n52959 , n52960 );
nand ( n52962 , n52949 , n52961 );
not ( n52963 , n52962 );
buf ( n230725 , n32400 );
xor ( n230726 , n230725 , n40178 );
xnor ( n52966 , n230726 , n36189 );
not ( n52967 , n52966 );
or ( n52968 , n52963 , n52967 );
not ( n52969 , n52966 );
not ( n230731 , n52969 );
or ( n230732 , n230731 , n52962 );
nand ( n52972 , n52968 , n230732 );
not ( n52973 , n52972 );
not ( n52974 , n52973 );
or ( n52975 , n52942 , n52974 );
nand ( n230737 , n52972 , n230701 );
nand ( n230738 , n52975 , n230737 );
not ( n52978 , n230738 );
not ( n230740 , n52978 );
and ( n52980 , n52901 , n230740 );
and ( n52981 , n52900 , n52978 );
nor ( n52982 , n52980 , n52981 );
not ( n52983 , n52982 );
or ( n230745 , n52799 , n52983 );
not ( n230746 , n52798 );
and ( n52986 , n52900 , n230738 );
not ( n52987 , n52900 );
and ( n52988 , n52987 , n52978 );
nor ( n52989 , n52986 , n52988 );
nand ( n52990 , n230746 , n52989 );
nand ( n52991 , n230745 , n52990 );
and ( n230753 , n51693 , n51742 );
not ( n230754 , n51693 );
and ( n52994 , n230754 , n229506 );
nor ( n52995 , n230753 , n52994 );
buf ( n52996 , n52995 );
not ( n52997 , n52996 );
and ( n52998 , n52991 , n52997 );
not ( n52999 , n52991 );
and ( n53000 , n52999 , n52996 );
nor ( n53001 , n52998 , n53000 );
nand ( n53002 , n52761 , n53001 );
or ( n230764 , n230208 , n53002 );
nor ( n230765 , n230205 , n221279 );
nand ( n230766 , n230765 , n53002 );
nand ( n230767 , n31576 , n25615 );
nand ( n53007 , n230764 , n230766 , n230767 );
buf ( n53008 , n53007 );
not ( n53009 , RI19aad468_2473);
or ( n53010 , n25328 , n53009 );
not ( n53011 , RI19aa3238_2544);
or ( n53012 , n226822 , n53011 );
nand ( n53013 , n53010 , n53012 );
buf ( n53014 , n53013 );
not ( n53015 , n42016 );
not ( n230777 , n41649 );
buf ( n230778 , n41673 );
not ( n230779 , n230778 );
nand ( n230780 , n230777 , n230779 );
not ( n53020 , n230780 );
or ( n230782 , n53015 , n53020 );
or ( n230783 , n230780 , n42016 );
nand ( n53023 , n230782 , n230783 );
not ( n230785 , n53023 );
not ( n230786 , n230785 );
nand ( n53026 , n219882 , n41829 );
not ( n53027 , n53026 );
not ( n53028 , n42132 );
not ( n53029 , n53028 );
or ( n230791 , n53027 , n53029 );
or ( n230792 , n53028 , n53026 );
nand ( n53032 , n230791 , n230792 );
not ( n53033 , n53032 );
not ( n53034 , n42099 );
nand ( n53035 , n41892 , n53034 );
not ( n230797 , n53035 );
not ( n230798 , n42081 );
not ( n53038 , n230798 );
and ( n53039 , n230797 , n53038 );
nand ( n53040 , n41892 , n53034 );
and ( n53041 , n53040 , n230798 );
nor ( n53042 , n53039 , n53041 );
not ( n53043 , n53042 );
or ( n53044 , n53033 , n53043 );
not ( n53045 , n53032 );
not ( n230807 , n53042 );
nand ( n230808 , n53045 , n230807 );
nand ( n230809 , n53044 , n230808 );
not ( n230810 , n230809 );
not ( n53050 , n230810 );
not ( n230812 , n41993 );
nand ( n230813 , n42015 , n41649 );
and ( n53053 , n230813 , n42029 );
not ( n53054 , n230813 );
not ( n53055 , n42029 );
and ( n53056 , n53054 , n53055 );
nor ( n230818 , n53053 , n53056 );
not ( n230819 , n230818 );
or ( n53059 , n230812 , n230819 );
or ( n230821 , n230818 , n41993 );
nand ( n230822 , n53059 , n230821 );
nand ( n53062 , n219823 , n41806 );
and ( n53063 , n53062 , n42049 );
not ( n53064 , n53062 );
not ( n53065 , n42049 );
and ( n230827 , n53064 , n53065 );
nor ( n230828 , n53063 , n230827 );
and ( n53068 , n230822 , n230828 );
not ( n53069 , n230822 );
not ( n53070 , n230828 );
and ( n53071 , n53069 , n53070 );
nor ( n230833 , n53068 , n53071 );
not ( n230834 , n230833 );
and ( n53074 , n53050 , n230834 );
and ( n53075 , n230810 , n230833 );
nor ( n53076 , n53074 , n53075 );
not ( n53077 , n53076 );
not ( n230839 , n53077 );
or ( n230840 , n230786 , n230839 );
xnor ( n53080 , n230809 , n230833 );
not ( n53081 , n53080 );
or ( n53082 , n53081 , n230785 );
nand ( n53083 , n230840 , n53082 );
not ( n230845 , n53083 );
not ( n230846 , n42409 );
nand ( n53086 , n220157 , n43648 );
not ( n53087 , n53086 );
or ( n53088 , n230846 , n53087 );
or ( n53089 , n53086 , n42409 );
nand ( n230851 , n53088 , n53089 );
not ( n230852 , n230851 );
nand ( n53092 , n42333 , n43596 );
not ( n230854 , n53092 );
not ( n230855 , n42359 );
not ( n53095 , n230855 );
and ( n230857 , n230854 , n53095 );
and ( n230858 , n53092 , n230855 );
nor ( n53098 , n230857 , n230858 );
not ( n53099 , n53098 );
or ( n53100 , n230852 , n53099 );
or ( n53101 , n230851 , n53098 );
nand ( n230863 , n53100 , n53101 );
not ( n230864 , n43564 );
not ( n53104 , n230864 );
buf ( n53105 , n42180 );
nand ( n53106 , n53104 , n53105 );
xnor ( n53107 , n53106 , n42170 );
not ( n230869 , n53107 );
and ( n230870 , n230863 , n230869 );
not ( n53110 , n230863 );
and ( n53111 , n53110 , n53107 );
nor ( n53112 , n230870 , n53111 );
buf ( n53113 , n42211 );
not ( n230875 , n53113 );
nand ( n230876 , n230875 , n43682 );
not ( n53116 , n230876 );
not ( n53117 , n219982 );
not ( n53118 , n53117 );
and ( n53119 , n53116 , n53118 );
and ( n230881 , n230876 , n53117 );
nor ( n230882 , n53119 , n230881 );
not ( n53122 , n230882 );
not ( n53123 , n53122 );
not ( n53124 , n42295 );
nand ( n53125 , n43691 , n53124 );
not ( n230887 , n53125 );
not ( n230888 , n42251 );
and ( n53128 , n230887 , n230888 );
and ( n53129 , n53125 , n42251 );
nor ( n53130 , n53128 , n53129 );
not ( n53131 , n53130 );
or ( n230893 , n53123 , n53131 );
not ( n230894 , n53130 );
nand ( n53134 , n230894 , n230882 );
nand ( n53135 , n230893 , n53134 );
and ( n53136 , n53112 , n53135 );
not ( n53137 , n53112 );
not ( n230899 , n53135 );
and ( n230900 , n53137 , n230899 );
nor ( n53140 , n53136 , n230900 );
not ( n230902 , n53140 );
not ( n230903 , n230902 );
not ( n53143 , n230903 );
and ( n230905 , n230845 , n53143 );
not ( n230906 , n230902 );
and ( n53146 , n53083 , n230906 );
nor ( n53147 , n230905 , n53146 );
nor ( n53148 , n53147 , n35427 );
not ( n53149 , n33236 );
not ( n230911 , n205492 );
not ( n230912 , n25501 );
or ( n53152 , n230911 , n230912 );
not ( n230914 , n205492 );
nand ( n230915 , n230914 , n25508 );
nand ( n53155 , n53152 , n230915 );
and ( n53156 , n53155 , n37450 );
not ( n53157 , n53155 );
and ( n53158 , n53157 , n43936 );
nor ( n230920 , n53156 , n53158 );
not ( n230921 , n230920 );
nand ( n53161 , n32495 , n32507 );
not ( n53162 , n53161 );
or ( n53163 , n230921 , n53162 );
or ( n53164 , n53161 , n230920 );
nand ( n230926 , n53163 , n53164 );
not ( n230927 , n230926 );
not ( n53167 , n32609 );
nand ( n53168 , n53167 , n32785 );
not ( n53169 , n53168 );
not ( n53170 , n26376 );
not ( n53171 , n45695 );
or ( n230933 , n53170 , n53171 );
not ( n230934 , n26376 );
nand ( n53174 , n230934 , n41054 );
nand ( n53175 , n230933 , n53174 );
and ( n53176 , n53175 , n41041 );
not ( n53177 , n53175 );
and ( n53178 , n53177 , n41040 );
nor ( n230940 , n53176 , n53178 );
not ( n230941 , n230940 );
not ( n53181 , n230941 );
and ( n53182 , n53169 , n53181 );
and ( n53183 , n53168 , n230941 );
nor ( n53184 , n53182 , n53183 );
not ( n53185 , n53184 );
or ( n53186 , n230927 , n53185 );
or ( n53187 , n230926 , n53184 );
nand ( n53188 , n53186 , n53187 );
not ( n53189 , n32912 );
nand ( n53190 , n32918 , n53189 );
xor ( n230952 , n204463 , n47216 );
xnor ( n230953 , n230952 , n27968 );
not ( n53193 , n230953 );
and ( n53194 , n53190 , n53193 );
not ( n230956 , n53190 );
and ( n230957 , n230956 , n230953 );
nor ( n53197 , n53194 , n230957 );
and ( n53198 , n53188 , n53197 );
not ( n53199 , n53188 );
not ( n53200 , n53197 );
and ( n53201 , n53199 , n53200 );
nor ( n53202 , n53198 , n53201 );
not ( n53203 , n53202 );
not ( n230965 , n53203 );
nand ( n230966 , n33048 , n33008 );
not ( n53206 , n230966 );
not ( n230968 , n224874 );
not ( n230969 , n37320 );
not ( n53209 , n42355 );
or ( n53210 , n230969 , n53209 );
or ( n53211 , n41756 , n37320 );
nand ( n53212 , n53210 , n53211 );
not ( n53213 , n53212 );
or ( n53214 , n230968 , n53213 );
or ( n53215 , n53212 , n228145 );
nand ( n53216 , n53214 , n53215 );
buf ( n53217 , n53216 );
not ( n53218 , n53217 );
and ( n230980 , n53206 , n53218 );
and ( n230981 , n230966 , n53217 );
nor ( n53221 , n230980 , n230981 );
not ( n53222 , n53221 );
not ( n53223 , n33191 );
nand ( n53224 , n33231 , n53223 );
not ( n230986 , n33497 );
not ( n230987 , n28555 );
or ( n53227 , n230986 , n230987 );
nand ( n53228 , n225104 , n33493 );
nand ( n53229 , n53227 , n53228 );
and ( n53230 , n53229 , n38257 );
not ( n230992 , n53229 );
and ( n230993 , n230992 , n47346 );
nor ( n53233 , n53230 , n230993 );
not ( n230995 , n53233 );
and ( n230996 , n53224 , n230995 );
not ( n53236 , n53224 );
and ( n230998 , n53236 , n53233 );
nor ( n230999 , n230996 , n230998 );
not ( n53239 , n230999 );
or ( n231001 , n53222 , n53239 );
not ( n231002 , n230999 );
not ( n53242 , n53221 );
nand ( n53243 , n231002 , n53242 );
nand ( n53244 , n231001 , n53243 );
not ( n53245 , n53244 );
and ( n231007 , n230965 , n53245 );
and ( n231008 , n53203 , n53244 );
nor ( n53248 , n231007 , n231008 );
not ( n53249 , n53248 );
or ( n53250 , n53149 , n53249 );
not ( n53251 , n33236 );
not ( n231013 , n53202 );
not ( n231014 , n53244 );
not ( n53254 , n231014 );
or ( n53255 , n231013 , n53254 );
nand ( n53256 , n53203 , n53244 );
nand ( n53257 , n53255 , n53256 );
nand ( n231019 , n53251 , n53257 );
nand ( n231020 , n53250 , n231019 );
not ( n53260 , n218918 );
not ( n53261 , n204411 );
and ( n53262 , n53260 , n53261 );
and ( n53263 , n45111 , n204411 );
nor ( n231025 , n53262 , n53263 );
and ( n231026 , n231025 , n37123 );
not ( n53266 , n231025 );
and ( n53267 , n53266 , n37128 );
nor ( n53268 , n231026 , n53267 );
buf ( n53269 , n53268 );
not ( n231031 , n53269 );
not ( n231032 , n43735 );
buf ( n53272 , n29560 );
not ( n53273 , n53272 );
nor ( n53274 , n53273 , n225200 );
not ( n53275 , n53274 );
not ( n231037 , n53272 );
nand ( n231038 , n231037 , n43201 );
nand ( n53278 , n53275 , n231038 );
not ( n231040 , n53278 );
and ( n231041 , n231032 , n231040 );
and ( n53281 , n33047 , n53278 );
nor ( n53282 , n231041 , n53281 );
not ( n53283 , n53282 );
not ( n53284 , n29907 );
not ( n231046 , n41082 );
or ( n231047 , n53284 , n231046 );
or ( n53287 , n32900 , n29907 );
nand ( n53288 , n231047 , n53287 );
and ( n53289 , n53288 , n32906 );
not ( n53290 , n53288 );
and ( n231052 , n53290 , n32910 );
nor ( n231053 , n53289 , n231052 );
nand ( n53293 , n53283 , n231053 );
not ( n53294 , n53293 );
or ( n53295 , n231031 , n53294 );
or ( n53296 , n53293 , n53269 );
nand ( n53297 , n53295 , n53296 );
buf ( n53298 , n37095 );
xor ( n231060 , n53298 , n35291 );
xnor ( n231061 , n231060 , n221462 );
buf ( n53301 , n37880 );
not ( n53302 , RI174a72b0_921);
and ( n53303 , n53301 , n53302 );
not ( n53304 , n53301 );
and ( n231066 , n53304 , n37877 );
nor ( n231067 , n53303 , n231066 );
not ( n53307 , n231067 );
not ( n53308 , n45817 );
or ( n53309 , n53307 , n53308 );
not ( n53310 , n231067 );
nand ( n231072 , n53310 , n45418 );
nand ( n231073 , n53309 , n231072 );
xor ( n53313 , n231073 , n222667 );
nand ( n53314 , n231061 , n53313 );
not ( n53315 , n53314 );
not ( n53316 , n28265 );
not ( n231078 , n48058 );
or ( n231079 , n53316 , n231078 );
nand ( n53319 , n48061 , n206029 );
nand ( n53320 , n231079 , n53319 );
and ( n53321 , n53320 , n34416 );
not ( n53322 , n53320 );
and ( n53323 , n53322 , n204586 );
nor ( n53324 , n53321 , n53323 );
not ( n231086 , n53324 );
and ( n231087 , n53315 , n231086 );
and ( n53327 , n53314 , n53324 );
nor ( n53328 , n231087 , n53327 );
and ( n53329 , n53297 , n53328 );
not ( n53330 , n53297 );
not ( n53331 , n53328 );
and ( n53332 , n53330 , n53331 );
nor ( n231094 , n53329 , n53332 );
not ( n231095 , n231094 );
xor ( n231096 , n28482 , n32862 );
xor ( n231097 , n231096 , n36262 );
not ( n53337 , n231097 );
not ( n53338 , n30638 );
buf ( n53339 , n45306 );
not ( n53340 , n53339 );
not ( n231102 , n53340 );
not ( n231103 , n30685 );
or ( n53343 , n231102 , n231103 );
nand ( n53344 , n208445 , n53339 );
nand ( n53345 , n53343 , n53344 );
not ( n53346 , n53345 );
and ( n231108 , n53338 , n53346 );
and ( n231109 , n30638 , n53345 );
nor ( n53349 , n231108 , n231109 );
not ( n53350 , n31750 );
not ( n53351 , n34299 );
or ( n53352 , n53350 , n53351 );
not ( n231114 , n31750 );
nand ( n231115 , n231114 , n34303 );
nand ( n53355 , n53352 , n231115 );
and ( n53356 , n53355 , n34264 );
not ( n53357 , n53355 );
and ( n53358 , n53357 , n34308 );
nor ( n231120 , n53356 , n53358 );
nand ( n231121 , n53349 , n231120 );
not ( n53361 , n231121 );
or ( n53362 , n53337 , n53361 );
or ( n53363 , n231121 , n231097 );
nand ( n53364 , n53362 , n53363 );
not ( n231126 , n53364 );
and ( n231127 , n210489 , n26100 );
not ( n53367 , n210489 );
and ( n53368 , n53367 , n26101 );
or ( n53369 , n231127 , n53368 );
and ( n53370 , n53369 , n45045 );
not ( n231132 , n53369 );
and ( n231133 , n231132 , n32783 );
nor ( n53373 , n53370 , n231133 );
not ( n231135 , n53373 );
buf ( n231136 , n32960 );
not ( n231137 , n231136 );
not ( n231138 , n38585 );
or ( n53378 , n231137 , n231138 );
or ( n53379 , n38585 , n231136 );
nand ( n53380 , n53378 , n53379 );
not ( n231142 , n38581 );
and ( n231143 , n53380 , n231142 );
not ( n231144 , n53380 );
and ( n231145 , n231144 , n29909 );
nor ( n53385 , n231143 , n231145 );
nand ( n53386 , n231135 , n53385 );
not ( n53387 , n53386 );
not ( n53388 , n27802 );
not ( n53389 , n30591 );
not ( n53390 , n27848 );
or ( n231152 , n53389 , n53390 );
buf ( n231153 , RI1744c518_1364);
nand ( n53393 , n27842 , n231153 );
nand ( n231155 , n231152 , n53393 );
not ( n231156 , n231155 );
or ( n53396 , n53388 , n231156 );
or ( n231158 , n231155 , n27802 );
nand ( n231159 , n53396 , n231158 );
not ( n53399 , n231159 );
and ( n53400 , n53387 , n53399 );
and ( n53401 , n53386 , n231159 );
nor ( n53402 , n53400 , n53401 );
not ( n231164 , n53402 );
or ( n231165 , n231126 , n231164 );
or ( n53405 , n53402 , n53364 );
nand ( n53406 , n231165 , n53405 );
not ( n53407 , n53406 );
and ( n53408 , n204780 , n43757 );
not ( n231170 , n204780 );
and ( n231171 , n231170 , n33183 );
or ( n53411 , n53408 , n231171 );
and ( n53412 , n53411 , n33187 );
not ( n53413 , n53411 );
and ( n53414 , n53413 , n33186 );
nor ( n231176 , n53412 , n53414 );
not ( n231177 , n231176 );
buf ( n53417 , n40725 );
buf ( n231179 , n53417 );
xor ( n231180 , n30068 , n231179 );
xnor ( n53420 , n231180 , n33303 );
nand ( n231182 , n231177 , n53420 );
not ( n231183 , n231182 );
not ( n53423 , n31719 );
not ( n53424 , n26409 );
or ( n53425 , n53423 , n53424 );
not ( n53426 , n26409 );
nand ( n53427 , n53426 , n31722 );
nand ( n53428 , n53425 , n53427 );
buf ( n231190 , n35590 );
and ( n231191 , n53428 , n231190 );
not ( n53431 , n53428 );
buf ( n53432 , n35584 );
and ( n53433 , n53431 , n53432 );
nor ( n53434 , n231191 , n53433 );
not ( n53435 , n53434 );
and ( n53436 , n231183 , n53435 );
not ( n231198 , n231176 );
nand ( n231199 , n53420 , n231198 );
and ( n53439 , n231199 , n53434 );
nor ( n53440 , n53436 , n53439 );
not ( n53441 , n53440 );
and ( n53442 , n53407 , n53441 );
and ( n231204 , n53406 , n53440 );
nor ( n231205 , n53442 , n231204 );
not ( n53445 , n231205 );
not ( n231207 , n53445 );
or ( n231208 , n231095 , n231207 );
not ( n53448 , n231094 );
nand ( n231210 , n231205 , n53448 );
nand ( n231211 , n231208 , n231210 );
buf ( n53451 , n231211 );
and ( n53452 , n231020 , n53451 );
not ( n53453 , n231020 );
not ( n53454 , n53451 );
and ( n231216 , n53453 , n53454 );
nor ( n231217 , n53452 , n231216 );
xor ( n53457 , n220035 , n223504 );
xnor ( n53458 , n53457 , n204825 );
not ( n53459 , n53458 );
not ( n53460 , n204669 );
not ( n231222 , n230718 );
or ( n231223 , n53460 , n231222 );
or ( n53463 , n230718 , n204669 );
nand ( n53464 , n231223 , n53463 );
not ( n53465 , n45672 );
and ( n53466 , n53464 , n53465 );
not ( n53467 , n53464 );
and ( n53468 , n53467 , n45672 );
nor ( n231230 , n53466 , n53468 );
nand ( n231231 , n53459 , n231230 );
not ( n53471 , n204591 );
not ( n53472 , n43577 );
not ( n53473 , n53472 );
or ( n53474 , n53471 , n53473 );
or ( n231236 , n53472 , n204591 );
nand ( n231237 , n53474 , n231236 );
not ( n53477 , n231237 );
not ( n231239 , n33957 );
and ( n53479 , n53477 , n231239 );
and ( n53480 , n231237 , n33957 );
nor ( n53481 , n53479 , n53480 );
and ( n53482 , n231231 , n53481 );
not ( n231244 , n231231 );
not ( n231245 , n53481 );
and ( n53485 , n231244 , n231245 );
nor ( n53486 , n53482 , n53485 );
not ( n53487 , n53486 );
nand ( n53488 , n53458 , n53481 );
xor ( n53489 , n34054 , n229405 );
xnor ( n53490 , n53489 , n41258 );
and ( n53491 , n53488 , n53490 );
not ( n53492 , n53488 );
not ( n231254 , n53490 );
and ( n231255 , n53492 , n231254 );
nor ( n53495 , n53491 , n231255 );
not ( n231257 , n48072 );
not ( n231258 , RI173eb678_1608);
not ( n53498 , n31028 );
xor ( n53499 , n231258 , n53498 );
xnor ( n53500 , n53499 , n31035 );
not ( n53501 , n53500 );
or ( n231263 , n231257 , n53501 );
or ( n231264 , n53500 , n48072 );
nand ( n53504 , n231263 , n231264 );
not ( n53505 , n53504 );
not ( n53506 , n53505 );
not ( n53507 , n31072 );
not ( n231269 , n31053 );
and ( n231270 , n53507 , n231269 );
and ( n53510 , n31072 , n31053 );
nor ( n53511 , n231270 , n53510 );
not ( n53512 , n53511 );
not ( n53513 , n53512 );
or ( n231275 , n53506 , n53513 );
nand ( n231276 , n53511 , n53504 );
nand ( n53516 , n231275 , n231276 );
buf ( n53517 , RI1740b310_1453);
not ( n53518 , n53517 );
not ( n53519 , n32278 );
not ( n231281 , n53519 );
or ( n231282 , n53518 , n231281 );
or ( n53522 , n53519 , n53517 );
nand ( n53523 , n231282 , n53522 );
not ( n231285 , n53523 );
not ( n231286 , n230285 );
and ( n53526 , n231285 , n231286 );
and ( n53527 , n53523 , n230285 );
nor ( n53528 , n53526 , n53527 );
nand ( n53529 , n53516 , n53528 );
not ( n231291 , n53529 );
not ( n231292 , n25726 );
not ( n53532 , n40007 );
or ( n53533 , n231292 , n53532 );
or ( n53534 , n40007 , n25726 );
nand ( n53535 , n53533 , n53534 );
not ( n231297 , n53535 );
not ( n231298 , n30607 );
or ( n53538 , n231297 , n231298 );
not ( n53539 , n53535 );
nand ( n53540 , n53539 , n41891 );
nand ( n53541 , n53538 , n53540 );
not ( n231303 , n53541 );
or ( n231304 , n231291 , n231303 );
or ( n53544 , n53541 , n53529 );
nand ( n53545 , n231304 , n53544 );
not ( n53546 , n53545 );
not ( n53547 , n53546 );
nand ( n231309 , n25592 , n34298 );
not ( n231310 , n231309 );
nor ( n53550 , n25592 , n34298 );
nor ( n53551 , n231310 , n53550 );
not ( n53552 , n53551 );
not ( n53553 , n32483 );
or ( n231315 , n53552 , n53553 );
or ( n231316 , n29773 , n53551 );
nand ( n53556 , n231315 , n231316 );
xor ( n53557 , n32029 , n38676 );
xnor ( n53558 , n53557 , n36685 );
nand ( n53559 , n53556 , n53558 );
not ( n231321 , n27933 );
nand ( n231322 , n231321 , n33848 );
not ( n53562 , n231322 );
nor ( n231324 , n33848 , n27937 );
nor ( n231325 , n53562 , n231324 );
not ( n231326 , n231325 );
not ( n231327 , n36258 );
not ( n53567 , n231327 );
or ( n231329 , n231326 , n53567 );
not ( n231330 , n231325 );
nand ( n53570 , n231330 , n36258 );
nand ( n231332 , n231329 , n53570 );
and ( n53572 , n53559 , n231332 );
not ( n231334 , n53559 );
not ( n231335 , n231332 );
and ( n53575 , n231334 , n231335 );
nor ( n53576 , n53572 , n53575 );
not ( n53577 , n53576 );
not ( n53578 , n53577 );
or ( n231340 , n53547 , n53578 );
nand ( n231341 , n53576 , n53545 );
nand ( n53581 , n231340 , n231341 );
xor ( n53582 , n53495 , n53581 );
xor ( n53583 , n38892 , n47879 );
xnor ( n53584 , n53583 , n26222 );
not ( n231346 , n31071 );
not ( n231347 , n34914 );
or ( n53587 , n231346 , n231347 );
not ( n53588 , n31071 );
nand ( n53589 , n53588 , n52884 );
nand ( n53590 , n53587 , n53589 );
and ( n231352 , n53590 , n45854 );
not ( n231353 , n53590 );
and ( n53593 , n231353 , n45849 );
nor ( n53594 , n231352 , n53593 );
nand ( n53595 , n53584 , n53594 );
not ( n53596 , n53595 );
not ( n231358 , n25990 );
not ( n231359 , n33935 );
or ( n53599 , n231358 , n231359 );
nand ( n231361 , n41076 , n25986 );
nand ( n231362 , n53599 , n231361 );
and ( n53602 , n231362 , n43279 );
not ( n53603 , n231362 );
and ( n53604 , n53603 , n41071 );
nor ( n53605 , n53602 , n53604 );
not ( n231367 , n53605 );
and ( n231368 , n53596 , n231367 );
and ( n53608 , n53595 , n53605 );
nor ( n53609 , n231368 , n53608 );
not ( n53610 , n53609 );
not ( n53611 , n36135 );
not ( n231373 , n38347 );
or ( n231374 , n53611 , n231373 );
nand ( n53614 , n227521 , n36131 );
nand ( n53615 , n231374 , n53614 );
not ( n53616 , n38356 );
and ( n53617 , n53615 , n53616 );
not ( n231379 , n53615 );
and ( n231380 , n231379 , n38356 );
nor ( n53620 , n53617 , n231380 );
not ( n53621 , n53620 );
and ( n53622 , n38279 , n30889 );
not ( n53623 , n38279 );
and ( n231385 , n53623 , n30890 );
nor ( n231386 , n53622 , n231385 );
not ( n53626 , n231386 );
not ( n53627 , n33986 );
and ( n53628 , n53626 , n53627 );
and ( n53629 , n231386 , n34004 );
nor ( n231391 , n53628 , n53629 );
not ( n231392 , n33880 );
not ( n53632 , n33883 );
or ( n53633 , n231392 , n53632 );
not ( n53634 , n33883 );
not ( n53635 , RI174a5870_929);
nand ( n231397 , n53634 , n53635 );
nand ( n231398 , n53633 , n231397 );
not ( n53638 , n231398 );
nor ( n53639 , n53638 , n205214 );
not ( n53640 , n53639 );
not ( n53641 , n231398 );
nand ( n231403 , n53641 , n205214 );
nand ( n231404 , n53640 , n231403 );
and ( n53644 , n231404 , n43913 );
not ( n53645 , n231404 );
and ( n53646 , n53645 , n35200 );
nor ( n53647 , n53644 , n53646 );
nand ( n53648 , n231391 , n53647 );
not ( n231410 , n53648 );
or ( n231411 , n53621 , n231410 );
or ( n231412 , n53648 , n53620 );
nand ( n231413 , n231411 , n231412 );
not ( n53653 , n231413 );
and ( n53654 , n53610 , n53653 );
and ( n53655 , n53609 , n231413 );
nor ( n53656 , n53654 , n53655 );
xor ( n53657 , n53582 , n53656 );
not ( n53658 , n53657 );
or ( n53659 , n53487 , n53658 );
not ( n231421 , n53657 );
not ( n231422 , n53486 );
nand ( n231423 , n231421 , n231422 );
nand ( n231424 , n53659 , n231423 );
not ( n53664 , n34448 );
not ( n53665 , n53664 );
and ( n53666 , n231424 , n53665 );
not ( n53667 , n231424 );
not ( n53668 , n34439 );
not ( n53669 , n53668 );
and ( n53670 , n53667 , n53669 );
nor ( n231432 , n53666 , n53670 );
nor ( n231433 , n231217 , n231432 );
nand ( n53673 , n53148 , n231433 );
not ( n53674 , n231432 );
not ( n53675 , n53674 );
not ( n53676 , n53147 );
not ( n231438 , n53676 );
or ( n231439 , n53675 , n231438 );
not ( n53679 , n231217 );
buf ( n53680 , n47173 );
nor ( n53681 , n53679 , n53680 );
nand ( n53682 , n231439 , n53681 );
buf ( n231444 , n35431 );
nand ( n231445 , n231444 , n31822 );
nand ( n53685 , n53673 , n53682 , n231445 );
buf ( n53686 , n53685 );
not ( n53687 , n32925 );
not ( n53688 , n53687 );
not ( n231450 , n53248 );
or ( n231451 , n53688 , n231450 );
not ( n53691 , n53687 );
nand ( n53692 , n53691 , n53257 );
nand ( n53693 , n231451 , n53692 );
not ( n53694 , n53451 );
and ( n53695 , n53693 , n53694 );
not ( n53696 , n53693 );
and ( n53697 , n53696 , n53451 );
nor ( n231459 , n53695 , n53697 );
not ( n231460 , n231459 );
not ( n53700 , n228194 );
not ( n53701 , n50305 );
nand ( n53702 , n53701 , n50319 );
not ( n53703 , n53702 );
not ( n231465 , n31703 );
xor ( n231466 , n26388 , n26406 );
xor ( n53706 , n231466 , n45690 );
not ( n231468 , n53706 );
or ( n231469 , n231465 , n231468 );
or ( n53709 , n53706 , n31703 );
nand ( n53710 , n231469 , n53709 );
and ( n53711 , n53710 , n35590 );
not ( n53712 , n53710 );
and ( n231474 , n53712 , n53432 );
nor ( n231475 , n53711 , n231474 );
buf ( n53715 , n231475 );
not ( n53716 , n53715 );
and ( n53717 , n53703 , n53716 );
and ( n53718 , n53702 , n53715 );
nor ( n231480 , n53717 , n53718 );
not ( n231481 , n231480 );
not ( n53721 , n50327 );
nand ( n231483 , n53721 , n228111 );
nand ( n231484 , n40006 , n25749 );
not ( n53724 , n231484 );
nor ( n53725 , n40006 , n25749 );
nor ( n53726 , n53724 , n53725 );
and ( n53727 , n53726 , n30607 );
not ( n231489 , n53726 );
and ( n231490 , n231489 , n41891 );
or ( n53730 , n53727 , n231490 );
and ( n53731 , n231483 , n53730 );
not ( n53732 , n231483 );
not ( n53733 , n53730 );
and ( n53734 , n53732 , n53733 );
nor ( n53735 , n53731 , n53734 );
not ( n53736 , n53735 );
or ( n53737 , n231481 , n53736 );
or ( n231499 , n53735 , n231480 );
nand ( n231500 , n53737 , n231499 );
nand ( n53740 , n50386 , n50367 );
not ( n231502 , n31673 );
not ( n231503 , n205344 );
not ( n53743 , n31829 );
or ( n231505 , n231503 , n53743 );
or ( n231506 , n48905 , n205344 );
nand ( n53746 , n231505 , n231506 );
not ( n231508 , n53746 );
or ( n231509 , n231502 , n231508 );
or ( n53749 , n53746 , n38709 );
nand ( n53750 , n231509 , n53749 );
not ( n53751 , n53750 );
and ( n53752 , n53740 , n53751 );
not ( n231514 , n53740 );
and ( n231515 , n231514 , n53750 );
nor ( n53755 , n53752 , n231515 );
not ( n53756 , n53755 );
and ( n53757 , n231500 , n53756 );
not ( n53758 , n231500 );
and ( n231520 , n53758 , n53755 );
nor ( n231521 , n53757 , n231520 );
not ( n53761 , n228222 );
not ( n53762 , n228208 );
nand ( n53763 , n53761 , n53762 );
buf ( n53764 , n30683 );
not ( n53765 , n53764 );
not ( n53766 , n227301 );
or ( n231528 , n53765 , n53766 );
not ( n231529 , n53764 );
nand ( n231530 , n231529 , n40620 );
nand ( n231531 , n231528 , n231530 );
and ( n53771 , n231531 , n39922 );
not ( n53772 , n231531 );
and ( n53773 , n53772 , n227306 );
nor ( n53774 , n53771 , n53773 );
buf ( n231536 , n53774 );
and ( n231537 , n53763 , n231536 );
not ( n53777 , n53763 );
not ( n53778 , n231536 );
and ( n53779 , n53777 , n53778 );
nor ( n53780 , n231537 , n53779 );
not ( n231542 , n53780 );
not ( n231543 , n231542 );
not ( n53783 , n50417 );
nand ( n53784 , n53783 , n50405 );
not ( n53785 , n53784 );
not ( n53786 , n52852 );
buf ( n53787 , n30134 );
not ( n53788 , n53787 );
and ( n53789 , n53786 , n53788 );
and ( n231551 , n205833 , n53787 );
nor ( n231552 , n53789 , n231551 );
and ( n231553 , n231552 , n28122 );
not ( n231554 , n231552 );
and ( n53794 , n231554 , n28125 );
nor ( n53795 , n231553 , n53794 );
not ( n53796 , n53795 );
not ( n53797 , n53796 );
not ( n231559 , n53797 );
and ( n231560 , n53785 , n231559 );
and ( n53800 , n53784 , n53797 );
nor ( n53801 , n231560 , n53800 );
not ( n53802 , n53801 );
not ( n53803 , n53802 );
or ( n231565 , n231543 , n53803 );
nand ( n231566 , n53801 , n53780 );
nand ( n53806 , n231565 , n231566 );
and ( n53807 , n231521 , n53806 );
not ( n53808 , n231521 );
not ( n53809 , n53806 );
and ( n53810 , n53808 , n53809 );
nor ( n53811 , n53807 , n53810 );
not ( n231573 , n53811 );
or ( n231574 , n53700 , n231573 );
not ( n53814 , n228194 );
not ( n53815 , n53809 );
not ( n53816 , n231521 );
not ( n53817 , n53816 );
or ( n231579 , n53815 , n53817 );
nand ( n231580 , n231521 , n53806 );
nand ( n53820 , n231579 , n231580 );
nand ( n53821 , n53814 , n53820 );
nand ( n53822 , n231574 , n53821 );
xor ( n53823 , n36642 , n36660 );
not ( n231585 , n36651 );
xnor ( n231586 , n53823 , n231585 );
xor ( n53826 , n25568 , n231586 );
and ( n53827 , n53826 , n28780 );
not ( n231589 , n53826 );
and ( n231590 , n231589 , n222443 );
nor ( n231591 , n53827 , n231590 );
not ( n231592 , n231591 );
not ( n53832 , n45942 );
not ( n53833 , n221432 );
and ( n53834 , n53832 , n53833 );
and ( n53835 , n45942 , n221432 );
nor ( n231597 , n53834 , n53835 );
and ( n231598 , n42966 , n231597 );
not ( n53838 , n42966 );
not ( n53839 , n231597 );
and ( n53840 , n53838 , n53839 );
nor ( n53841 , n231598 , n53840 );
not ( n231603 , n53841 );
nand ( n231604 , n231592 , n231603 );
not ( n53844 , n231604 );
not ( n53845 , n32107 );
not ( n53846 , n29853 );
or ( n53847 , n53845 , n53846 );
not ( n231609 , n29859 );
or ( n231610 , n231609 , n32107 );
nand ( n53850 , n53847 , n231610 );
and ( n53851 , n53850 , n33614 );
not ( n53852 , n53850 );
and ( n53853 , n53852 , n33618 );
nor ( n231615 , n53851 , n53853 );
not ( n231616 , n231615 );
not ( n53856 , n231616 );
and ( n53857 , n53844 , n53856 );
not ( n53858 , n231591 );
nand ( n53859 , n53858 , n231603 );
and ( n231621 , n53859 , n231616 );
nor ( n231622 , n53857 , n231621 );
xor ( n53862 , n37178 , n229482 );
xnor ( n53863 , n53862 , n205230 );
not ( n53864 , n53863 );
not ( n53865 , n42346 );
not ( n231627 , n28146 );
or ( n231628 , n53865 , n231627 );
not ( n53868 , n42346 );
nand ( n53869 , n53868 , n44712 );
nand ( n53870 , n231628 , n53869 );
and ( n53871 , n53870 , n35275 );
not ( n231633 , n53870 );
and ( n231634 , n231633 , n44720 );
nor ( n53874 , n53871 , n231634 );
not ( n53875 , n53874 );
nand ( n53876 , n53864 , n53875 );
not ( n53877 , n30724 );
not ( n231639 , n31636 );
or ( n231640 , n53877 , n231639 );
or ( n53880 , n31636 , n30724 );
nand ( n53881 , n231640 , n53880 );
xor ( n53882 , n37506 , n53881 );
not ( n53883 , n53882 );
and ( n231645 , n53876 , n53883 );
not ( n231646 , n53876 );
and ( n53886 , n231646 , n53882 );
nor ( n231648 , n231645 , n53886 );
xor ( n231649 , n231622 , n231648 );
not ( n53889 , n36050 );
not ( n53890 , n37353 );
or ( n53891 , n53889 , n53890 );
nand ( n53892 , n37356 , n36047 );
nand ( n231654 , n53891 , n53892 );
and ( n231655 , n231654 , n36813 );
not ( n53895 , n231654 );
and ( n231657 , n53895 , n40678 );
nor ( n231658 , n231655 , n231657 );
not ( n53898 , n219430 );
buf ( n53899 , n205320 );
not ( n53900 , n53899 );
nor ( n53901 , n53900 , n36990 );
not ( n231663 , n53901 );
not ( n231664 , n53899 );
nand ( n53904 , n231664 , n34872 );
nand ( n53905 , n231663 , n53904 );
not ( n53906 , n53905 );
or ( n53907 , n53898 , n53906 );
or ( n231669 , n53905 , n219430 );
nand ( n231670 , n53907 , n231669 );
nand ( n53910 , n231658 , n231670 );
not ( n53911 , n53910 );
not ( n53912 , n53911 );
xor ( n53913 , n32929 , n29909 );
xnor ( n231675 , n53913 , n26009 );
not ( n231676 , n231675 );
not ( n53916 , n231676 );
or ( n53917 , n53912 , n53916 );
nand ( n53918 , n231675 , n53910 );
nand ( n53919 , n53917 , n53918 );
xor ( n231681 , n231649 , n53919 );
xor ( n231682 , n29667 , n34700 );
xnor ( n53922 , n231682 , n36859 );
not ( n53923 , n53922 );
xor ( n53924 , n27694 , n25509 );
not ( n53925 , n25457 );
not ( n231687 , n53925 );
xnor ( n231688 , n53924 , n231687 );
not ( n53928 , n231688 );
buf ( n231690 , n35264 );
not ( n231691 , n231690 );
not ( n53931 , n231691 );
not ( n231693 , n52070 );
or ( n231694 , n53931 , n231693 );
nand ( n53934 , n223711 , n231690 );
nand ( n53935 , n231694 , n53934 );
not ( n53936 , n53935 );
not ( n53937 , n43635 );
not ( n231699 , n53937 );
not ( n231700 , n231699 );
and ( n53940 , n53936 , n231700 );
and ( n231702 , n53935 , n231699 );
nor ( n231703 , n53940 , n231702 );
not ( n53943 , n231703 );
nand ( n53944 , n53928 , n53943 );
not ( n53945 , n53944 );
or ( n53946 , n53923 , n53945 );
not ( n231708 , n231703 );
nand ( n231709 , n231708 , n53928 );
or ( n53949 , n231709 , n53922 );
nand ( n53950 , n53946 , n53949 );
not ( n53951 , n53950 );
not ( n53952 , n29277 );
not ( n231714 , n44347 );
or ( n231715 , n53952 , n231714 );
nand ( n53955 , n44351 , n29274 );
nand ( n53956 , n231715 , n53955 );
and ( n53957 , n53956 , n40697 );
not ( n53958 , n53956 );
and ( n53959 , n53958 , n205420 );
nor ( n53960 , n53957 , n53959 );
not ( n231722 , n41857 );
not ( n231723 , n206160 );
buf ( n53963 , n28402 );
not ( n53964 , n53963 );
or ( n53965 , n231723 , n53964 );
or ( n53966 , n53963 , n206160 );
nand ( n231728 , n53965 , n53966 );
not ( n231729 , n231728 );
not ( n53969 , n39007 );
or ( n53970 , n231729 , n53969 );
not ( n53971 , n231728 );
nand ( n53972 , n53971 , n39002 );
nand ( n231734 , n53970 , n53972 );
not ( n231735 , n231734 );
or ( n53975 , n231722 , n231735 );
or ( n53976 , n231734 , n41857 );
nand ( n53977 , n53975 , n53976 );
buf ( n53978 , n53977 );
nand ( n231740 , n53960 , n53978 );
not ( n231741 , n231740 );
buf ( n53981 , RI173f0538_1584);
not ( n53982 , n53981 );
not ( n53983 , n38806 );
not ( n53984 , n53983 );
or ( n231746 , n53982 , n53984 );
or ( n231747 , n38801 , n53981 );
nand ( n231748 , n231746 , n231747 );
and ( n231749 , n231748 , n40359 );
not ( n53989 , n231748 );
buf ( n53990 , n29088 );
and ( n53991 , n53989 , n53990 );
nor ( n53992 , n231749 , n53991 );
not ( n231754 , n53992 );
not ( n231755 , n231754 );
not ( n53995 , n231755 );
and ( n53996 , n231741 , n53995 );
and ( n53997 , n231740 , n231755 );
nor ( n53998 , n53996 , n53997 );
not ( n231760 , n53998 );
and ( n231761 , n53951 , n231760 );
and ( n54001 , n53950 , n53998 );
nor ( n54002 , n231761 , n54001 );
and ( n54003 , n231681 , n54002 );
not ( n54004 , n231681 );
not ( n54005 , n54002 );
and ( n54006 , n54004 , n54005 );
nor ( n231768 , n54003 , n54006 );
buf ( n231769 , n231768 );
and ( n54009 , n53822 , n231769 );
not ( n54010 , n53822 );
and ( n54011 , n231681 , n54005 );
not ( n54012 , n231681 );
and ( n54013 , n54012 , n54002 );
nor ( n231775 , n54011 , n54013 );
buf ( n231776 , n231775 );
and ( n54016 , n54010 , n231776 );
nor ( n54017 , n54009 , n54016 );
not ( n54018 , n54017 );
nand ( n54019 , n231460 , n54018 );
nand ( n231781 , n34656 , n34566 );
not ( n231782 , n231781 );
not ( n231783 , n37347 );
not ( n231784 , n32205 );
not ( n54024 , n42512 );
or ( n231786 , n231784 , n54024 );
not ( n231787 , n32205 );
nand ( n54027 , n231787 , n220278 );
nand ( n231789 , n231786 , n54027 );
not ( n231790 , n231789 );
or ( n54030 , n231783 , n231790 );
or ( n54031 , n231789 , n221604 );
nand ( n54032 , n54030 , n54031 );
not ( n54033 , n54032 );
and ( n231795 , n231782 , n54033 );
and ( n231796 , n231781 , n54032 );
nor ( n54036 , n231795 , n231796 );
buf ( n54037 , n54036 );
not ( n54038 , n54037 );
not ( n54039 , n37186 );
not ( n54040 , n25864 );
or ( n231802 , n54039 , n54040 );
not ( n231803 , RI1733ae28_2154);
nand ( n54043 , n25838 , n231803 );
nand ( n54044 , n231802 , n54043 );
not ( n54045 , n54044 );
not ( n54046 , n25861 );
or ( n54047 , n54045 , n54046 );
or ( n231809 , n25861 , n54044 );
nand ( n231810 , n54047 , n231809 );
and ( n54050 , n231810 , n28030 );
not ( n54051 , n231810 );
and ( n54052 , n54051 , n28043 );
nor ( n54053 , n54050 , n54052 );
not ( n231815 , n54053 );
nand ( n231816 , n231815 , n34879 );
not ( n54056 , n231816 );
not ( n54057 , n39579 );
and ( n54058 , n54056 , n54057 );
and ( n54059 , n231816 , n39579 );
nor ( n231821 , n54058 , n54059 );
not ( n231822 , n231821 );
not ( n54062 , n39537 );
not ( n231824 , n32837 );
not ( n231825 , n35857 );
or ( n54065 , n231824 , n231825 );
or ( n231827 , n35857 , n32837 );
nand ( n231828 , n54065 , n231827 );
and ( n54068 , n231828 , n30078 );
not ( n54069 , n231828 );
and ( n54070 , n54069 , n37537 );
nor ( n54071 , n54068 , n54070 );
nand ( n231833 , n54071 , n34768 );
not ( n231834 , n231833 );
and ( n54074 , n54062 , n231834 );
and ( n54075 , n39537 , n231833 );
nor ( n54076 , n54074 , n54075 );
not ( n54077 , n54076 );
not ( n231839 , n54077 );
or ( n231840 , n231822 , n231839 );
not ( n54080 , n231821 );
nand ( n54081 , n54076 , n54080 );
nand ( n54082 , n231840 , n54081 );
buf ( n54083 , n28583 );
not ( n231845 , n54083 );
not ( n231846 , n231845 );
not ( n54086 , n37397 );
or ( n54087 , n231846 , n54086 );
nand ( n54088 , n43888 , n54083 );
nand ( n54089 , n54087 , n54088 );
not ( n231851 , n54089 );
not ( n231852 , n30810 );
and ( n54092 , n231851 , n231852 );
and ( n231854 , n37407 , n54089 );
nor ( n231855 , n54092 , n231854 );
nand ( n54095 , n231855 , n34920 );
not ( n54096 , n39563 );
and ( n54097 , n54095 , n54096 );
not ( n54098 , n54095 );
and ( n231860 , n54098 , n39563 );
nor ( n231861 , n54097 , n231860 );
not ( n54101 , n231861 );
and ( n54102 , n54082 , n54101 );
not ( n54103 , n54082 );
and ( n54104 , n54103 , n231861 );
nor ( n54105 , n54102 , n54104 );
not ( n54106 , n54105 );
not ( n231868 , n54106 );
buf ( n231869 , n39498 );
not ( n54109 , n231869 );
not ( n54110 , n39510 );
nand ( n54111 , n54110 , n34616 );
not ( n54112 , n54111 );
or ( n231874 , n54109 , n54112 );
or ( n231875 , n54111 , n231869 );
nand ( n54115 , n231874 , n231875 );
not ( n54116 , n54115 );
not ( n54117 , n54032 );
nand ( n54118 , n54117 , n34657 );
not ( n231880 , n54118 );
not ( n231881 , n212240 );
not ( n54121 , n231881 );
not ( n54122 , n54121 );
and ( n54123 , n231880 , n54122 );
and ( n54124 , n54118 , n54121 );
nor ( n54125 , n54123 , n54124 );
not ( n54126 , n54125 );
and ( n54127 , n54116 , n54126 );
and ( n54128 , n54115 , n54125 );
nor ( n54129 , n54127 , n54128 );
not ( n231891 , n54129 );
or ( n231892 , n231868 , n231891 );
not ( n231893 , n54129 );
nand ( n231894 , n231893 , n54105 );
nand ( n54134 , n231892 , n231894 );
not ( n231896 , n54134 );
or ( n231897 , n54038 , n231896 );
or ( n54137 , n54134 , n54037 );
nand ( n54138 , n231897 , n54137 );
nand ( n54139 , n46103 , n35158 );
not ( n54140 , n54139 );
not ( n231902 , n39643 );
and ( n231903 , n54140 , n231902 );
nand ( n54143 , n46103 , n35158 );
and ( n54144 , n54143 , n39643 );
nor ( n54145 , n231903 , n54144 );
not ( n54146 , n54145 );
nand ( n54147 , n46116 , n35043 );
not ( n54148 , n39657 );
and ( n231910 , n54147 , n54148 );
not ( n231911 , n54147 );
and ( n54151 , n231911 , n39657 );
nor ( n54152 , n231910 , n54151 );
not ( n54153 , n54152 );
or ( n54154 , n54146 , n54153 );
or ( n54155 , n54152 , n54145 );
nand ( n231917 , n54154 , n54155 );
not ( n231918 , n46134 );
nand ( n54158 , n231918 , n35209 );
not ( n231920 , n54158 );
not ( n231921 , n39681 );
and ( n54161 , n231920 , n231921 );
and ( n231923 , n54158 , n39681 );
nor ( n231924 , n54161 , n231923 );
not ( n54164 , n231924 );
and ( n54165 , n231917 , n54164 );
not ( n54166 , n231917 );
and ( n54167 , n54166 , n231924 );
nor ( n231929 , n54165 , n54167 );
nand ( n231930 , n35396 , n223938 );
not ( n54170 , n231930 );
not ( n54171 , n39735 );
not ( n54172 , n54171 );
not ( n54173 , n54172 );
and ( n54174 , n54170 , n54173 );
and ( n54175 , n231930 , n54172 );
nor ( n54176 , n54174 , n54175 );
not ( n54177 , n46157 );
nand ( n231939 , n54177 , n35294 );
buf ( n231940 , n217478 );
not ( n54180 , n231940 );
and ( n54181 , n231939 , n54180 );
not ( n54182 , n231939 );
and ( n54183 , n54182 , n231940 );
nor ( n231945 , n54181 , n54183 );
xor ( n231946 , n54176 , n231945 );
and ( n54186 , n231929 , n231946 );
not ( n54187 , n231929 );
not ( n54188 , n231946 );
and ( n54189 , n54187 , n54188 );
nor ( n231951 , n54186 , n54189 );
not ( n231952 , n231951 );
not ( n54192 , n231952 );
and ( n54193 , n54138 , n54192 );
not ( n54194 , n54138 );
buf ( n54195 , n231951 );
buf ( n231957 , n54195 );
not ( n231958 , n231957 );
and ( n54198 , n54194 , n231958 );
nor ( n54199 , n54193 , n54198 );
not ( n54200 , n40465 );
nand ( n54201 , n54199 , n54200 );
or ( n231963 , n54019 , n54201 );
nor ( n231964 , n54199 , n219702 );
nand ( n54204 , n54019 , n231964 );
nand ( n231966 , n31577 , n36135 );
nand ( n54206 , n231963 , n54204 , n231966 );
buf ( n54207 , n54206 );
buf ( n54208 , n35427 );
nor ( n54209 , n51759 , n54208 );
not ( n54210 , n41167 );
not ( n54211 , n40952 );
nand ( n231973 , n54211 , n40937 );
not ( n231974 , n231973 );
not ( n54214 , n42642 );
and ( n231976 , n231974 , n54214 );
and ( n231977 , n231973 , n42642 );
nor ( n54217 , n231976 , n231977 );
not ( n54218 , n54217 );
nand ( n54219 , n41028 , n40973 );
not ( n54220 , n42564 );
and ( n54221 , n54219 , n54220 );
not ( n54222 , n54219 );
and ( n231984 , n54222 , n42564 );
nor ( n231985 , n54221 , n231984 );
not ( n54225 , n231985 );
or ( n54226 , n54218 , n54225 );
or ( n54227 , n231985 , n54217 );
nand ( n54228 , n54226 , n54227 );
not ( n231990 , n41056 );
nand ( n231991 , n231990 , n41085 );
not ( n54231 , n42536 );
and ( n54232 , n231991 , n54231 );
not ( n54233 , n231991 );
and ( n54234 , n54233 , n42536 );
nor ( n231996 , n54232 , n54234 );
not ( n231997 , n231996 );
and ( n54237 , n54228 , n231997 );
not ( n54238 , n54228 );
and ( n54239 , n54238 , n231996 );
nor ( n54240 , n54237 , n54239 );
not ( n232002 , n54240 );
nand ( n232003 , n41197 , n41201 );
and ( n54243 , n232003 , n42454 );
not ( n54244 , n232003 );
and ( n54245 , n54244 , n220214 );
or ( n54246 , n54243 , n54245 );
not ( n232008 , n54246 );
not ( n232009 , n42664 );
not ( n54249 , n41115 );
nand ( n232011 , n41105 , n54249 );
not ( n232012 , n232011 );
or ( n54252 , n232009 , n232012 );
or ( n232014 , n42664 , n232011 );
nand ( n54254 , n54252 , n232014 );
not ( n54255 , n54254 );
or ( n54256 , n232008 , n54255 );
or ( n54257 , n54254 , n54246 );
nand ( n54258 , n54256 , n54257 );
not ( n232020 , n54258 );
and ( n232021 , n232002 , n232020 );
not ( n54261 , n232002 );
and ( n54262 , n54261 , n54258 );
nor ( n54263 , n232021 , n54262 );
not ( n54264 , n54263 );
or ( n54265 , n54210 , n54264 );
not ( n54266 , n41167 );
not ( n232028 , n54258 );
not ( n232029 , n54240 );
or ( n54269 , n232028 , n232029 );
not ( n54270 , n54258 );
not ( n54271 , n54240 );
nand ( n54272 , n54270 , n54271 );
nand ( n54273 , n54269 , n54272 );
nand ( n232035 , n54266 , n54273 );
nand ( n232036 , n54265 , n232035 );
not ( n54276 , n232036 );
not ( n54277 , n221852 );
nand ( n54278 , n54277 , n44102 );
and ( n54279 , n54278 , n42815 );
not ( n232041 , n54278 );
and ( n232042 , n232041 , n220577 );
nor ( n54282 , n54279 , n232042 );
not ( n54283 , n54282 );
not ( n54284 , n54283 );
not ( n54285 , n44117 );
nand ( n232047 , n44163 , n54285 );
not ( n232048 , n232047 );
not ( n54288 , n42788 );
and ( n54289 , n232048 , n54288 );
and ( n54290 , n232047 , n42788 );
nor ( n54291 , n54289 , n54290 );
not ( n232053 , n54291 );
not ( n232054 , n232053 );
or ( n54294 , n54284 , n232054 );
nand ( n54295 , n54291 , n54282 );
nand ( n54296 , n54294 , n54295 );
and ( n54297 , n54296 , n51282 );
not ( n232059 , n54296 );
and ( n232060 , n232059 , n51283 );
nor ( n54300 , n54297 , n232060 );
not ( n54301 , n54300 );
nand ( n54302 , n44028 , n44042 );
not ( n54303 , n54302 );
not ( n232065 , n220668 );
and ( n232066 , n54303 , n232065 );
and ( n54306 , n54302 , n220668 );
nor ( n54307 , n232066 , n54306 );
not ( n54308 , n54307 );
not ( n54309 , n54308 );
not ( n232071 , n221769 );
nand ( n232072 , n232071 , n43990 );
and ( n54312 , n232072 , n229080 );
not ( n54313 , n232072 );
and ( n54314 , n54313 , n42982 );
nor ( n54315 , n54312 , n54314 );
not ( n232077 , n54315 );
not ( n232078 , n232077 );
or ( n54318 , n54309 , n232078 );
nand ( n54319 , n54315 , n54307 );
nand ( n54320 , n54318 , n54319 );
and ( n54321 , n54301 , n54320 );
not ( n232083 , n54301 );
not ( n232084 , n54320 );
and ( n54324 , n232083 , n232084 );
nor ( n54325 , n54321 , n54324 );
not ( n54326 , n54325 );
and ( n54327 , n54276 , n54326 );
and ( n232089 , n232036 , n54325 );
nor ( n232090 , n54327 , n232089 );
nand ( n54330 , n54209 , n232090 , n52232 );
not ( n54331 , n232090 );
not ( n54332 , n51759 );
nand ( n54333 , n54332 , n52232 );
nand ( n232095 , n54331 , n54333 , n223839 );
nand ( n232096 , n41944 , n33531 );
nand ( n54336 , n54330 , n232095 , n232096 );
buf ( n54337 , n54336 );
buf ( n54338 , n31057 );
buf ( n54339 , n204329 );
buf ( n232101 , n26248 );
not ( n232102 , n25778 );
not ( n54342 , n39267 );
or ( n54343 , n232102 , n54342 );
or ( n54344 , n39267 , n25778 );
nand ( n54345 , n54343 , n54344 );
not ( n54346 , n54345 );
not ( n232108 , n38839 );
or ( n232109 , n54346 , n232108 );
or ( n232110 , n38839 , n54345 );
nand ( n232111 , n232109 , n232110 );
not ( n54351 , n232111 );
not ( n232113 , n40027 );
not ( n232114 , n30936 );
or ( n54354 , n232113 , n232114 );
nand ( n54355 , n30942 , n40030 );
nand ( n54356 , n54354 , n54355 );
not ( n54357 , n54356 );
not ( n232119 , n221779 );
and ( n232120 , n54357 , n232119 );
and ( n54360 , n54356 , n221779 );
nor ( n232122 , n232120 , n54360 );
not ( n232123 , n232122 );
nand ( n54363 , n54351 , n232123 );
and ( n54364 , n30116 , n28071 );
not ( n54365 , n30116 );
and ( n54366 , n54365 , n28070 );
nor ( n232128 , n54364 , n54366 );
and ( n232129 , n232128 , n28121 );
not ( n54369 , n232128 );
not ( n54370 , n28121 );
and ( n54371 , n54369 , n54370 );
nor ( n54372 , n232129 , n54371 );
not ( n232134 , n54372 );
and ( n232135 , n54363 , n232134 );
not ( n54375 , n54363 );
and ( n54376 , n54375 , n54372 );
nor ( n54377 , n232135 , n54376 );
not ( n54378 , n54377 );
not ( n232140 , n54378 );
buf ( n232141 , RI17408ef8_1464);
not ( n54381 , n232141 );
not ( n54382 , n32174 );
or ( n54383 , n54381 , n54382 );
not ( n54384 , n232141 );
nand ( n232146 , n54384 , n32180 );
nand ( n232147 , n54383 , n232146 );
not ( n54387 , n232147 );
not ( n232149 , n42091 );
and ( n232150 , n54387 , n232149 );
and ( n54390 , n232147 , n42091 );
nor ( n232152 , n232150 , n54390 );
not ( n232153 , n232152 );
not ( n54393 , n46586 );
not ( n232155 , n30500 );
and ( n232156 , n54393 , n232155 );
and ( n54396 , n46586 , n30500 );
nor ( n54397 , n232156 , n54396 );
not ( n54398 , n54397 );
not ( n54399 , n46595 );
not ( n232161 , n54399 );
or ( n232162 , n54398 , n232161 );
not ( n54402 , n46595 );
or ( n54403 , n54402 , n54397 );
nand ( n54404 , n232162 , n54403 );
not ( n54405 , n54404 );
nand ( n232167 , n232153 , n54405 );
not ( n232168 , n232167 );
not ( n54408 , n38514 );
not ( n54409 , n40150 );
not ( n54410 , n229405 );
or ( n54411 , n54409 , n54410 );
nand ( n232173 , n38558 , n40146 );
nand ( n232174 , n54411 , n232173 );
not ( n54414 , n232174 );
and ( n54415 , n54408 , n54414 );
and ( n54416 , n38514 , n232174 );
nor ( n54417 , n54415 , n54416 );
not ( n232179 , n54417 );
not ( n232180 , n232179 );
and ( n54420 , n232168 , n232180 );
and ( n54421 , n232167 , n232179 );
nor ( n54422 , n54420 , n54421 );
not ( n54423 , n54422 );
not ( n232185 , n54423 );
or ( n232186 , n232140 , n232185 );
nand ( n54426 , n54377 , n54422 );
nand ( n54427 , n232186 , n54426 );
buf ( n54428 , n54427 );
xor ( n54429 , n34667 , n40218 );
xnor ( n232191 , n54429 , n204892 );
not ( n232192 , n31054 );
not ( n54432 , n34914 );
or ( n54433 , n232192 , n54432 );
not ( n54434 , RI1744f308_1350);
nand ( n54435 , n34917 , n54434 );
nand ( n232197 , n54433 , n54435 );
and ( n232198 , n232197 , n45850 );
not ( n54438 , n232197 );
and ( n54439 , n54438 , n45855 );
nor ( n54440 , n232198 , n54439 );
nand ( n54441 , n232191 , n54440 );
not ( n232203 , n54441 );
not ( n232204 , n25615 );
not ( n54444 , n47958 );
or ( n54445 , n232204 , n54444 );
or ( n54446 , n47958 , n25615 );
nand ( n54447 , n54445 , n54446 );
not ( n232209 , n54447 );
not ( n232210 , n45268 );
and ( n54450 , n232209 , n232210 );
and ( n54451 , n54447 , n45268 );
nor ( n54452 , n54450 , n54451 );
not ( n54453 , n54452 );
not ( n232215 , n54453 );
and ( n232216 , n232203 , n232215 );
and ( n54456 , n54441 , n54453 );
nor ( n54457 , n232216 , n54456 );
buf ( n54458 , n54457 );
not ( n54459 , n54458 );
and ( n232221 , n54428 , n54459 );
not ( n232222 , n54428 );
and ( n54462 , n232222 , n54458 );
nor ( n232224 , n232221 , n54462 );
not ( n232225 , n33047 );
not ( n54465 , n29529 );
not ( n232227 , n38435 );
or ( n232228 , n54465 , n232227 );
or ( n54468 , n38436 , n29529 );
nand ( n54469 , n232228 , n54468 );
not ( n54470 , n54469 );
and ( n54471 , n232225 , n54470 );
and ( n232233 , n43735 , n54469 );
nor ( n232234 , n54471 , n232233 );
not ( n54474 , n204650 );
not ( n54475 , n42760 );
or ( n54476 , n54474 , n54475 );
nand ( n54477 , n50452 , n204647 );
nand ( n232239 , n54476 , n54477 );
and ( n232240 , n232239 , n53465 );
not ( n54480 , n232239 );
and ( n232242 , n54480 , n45672 );
nor ( n232243 , n232240 , n232242 );
nand ( n54483 , n232234 , n232243 );
not ( n54484 , n29881 );
not ( n54485 , n32900 );
or ( n54486 , n54484 , n54485 );
nand ( n232248 , n32903 , n29877 );
nand ( n232249 , n54486 , n232248 );
and ( n54489 , n232249 , n26475 );
not ( n54490 , n232249 );
and ( n54491 , n54490 , n32909 );
nor ( n54492 , n54489 , n54491 );
not ( n232254 , n54492 );
and ( n232255 , n54483 , n232254 );
not ( n54495 , n54483 );
and ( n54496 , n54495 , n54492 );
nor ( n54497 , n232255 , n54496 );
not ( n54498 , n54497 );
xor ( n232260 , n28531 , n30781 );
xnor ( n232261 , n232260 , n37407 );
buf ( n54501 , RI17404a10_1485);
not ( n54502 , n54501 );
not ( n54503 , n53417 );
or ( n54504 , n54502 , n54503 );
or ( n232266 , n53417 , n54501 );
nand ( n232267 , n54504 , n232266 );
and ( n54507 , n232267 , n42397 );
not ( n54508 , n232267 );
not ( n54509 , n42397 );
and ( n54510 , n54508 , n54509 );
nor ( n232272 , n54507 , n54510 );
nand ( n232273 , n232261 , n232272 );
not ( n54513 , n232273 );
not ( n54514 , n35126 );
not ( n54515 , n38770 );
or ( n54516 , n54514 , n54515 );
or ( n232278 , n38775 , n35126 );
nand ( n232279 , n54516 , n232278 );
and ( n54519 , n232279 , n29015 );
not ( n232281 , n232279 );
and ( n232282 , n232281 , n206777 );
nor ( n54522 , n54519 , n232282 );
not ( n232284 , n54522 );
and ( n232285 , n54513 , n232284 );
nand ( n54525 , n232272 , n232261 );
and ( n54526 , n54525 , n54522 );
nor ( n54527 , n232285 , n54526 );
not ( n54528 , n54527 );
or ( n232290 , n54498 , n54528 );
or ( n232291 , n54527 , n54497 );
nand ( n54531 , n232290 , n232291 );
buf ( n232293 , n54531 );
not ( n232294 , n232293 );
and ( n54534 , n232224 , n232294 );
not ( n54535 , n232224 );
and ( n54536 , n54535 , n232293 );
nor ( n54537 , n54534 , n54536 );
buf ( n232299 , n54537 );
not ( n232300 , n232299 );
not ( n54540 , n204621 );
and ( n54541 , n34896 , n204585 );
not ( n54542 , n34896 );
and ( n54543 , n54542 , n34415 );
nor ( n232305 , n54541 , n54543 );
not ( n232306 , n232305 );
not ( n54546 , n232306 );
or ( n54547 , n54540 , n54546 );
nand ( n54548 , n232305 , n204631 );
nand ( n54549 , n54547 , n54548 );
not ( n232311 , n54549 );
not ( n232312 , n31440 );
not ( n54552 , n29454 );
or ( n54553 , n232312 , n54552 );
not ( n54554 , n31440 );
nand ( n54555 , n54554 , n38682 );
nand ( n232317 , n54553 , n54555 );
and ( n232318 , n232317 , n38694 );
not ( n232319 , n232317 );
and ( n232320 , n232319 , n38691 );
nor ( n54560 , n232318 , n232320 );
not ( n54561 , n54560 );
nand ( n54562 , n232311 , n54561 );
not ( n54563 , n36626 );
not ( n232325 , n26216 );
not ( n232326 , n48779 );
or ( n54566 , n232325 , n232326 );
or ( n54567 , n48779 , n26216 );
nand ( n54568 , n54566 , n54567 );
not ( n54569 , n54568 );
or ( n232331 , n54563 , n54569 );
or ( n232332 , n54568 , n51936 );
nand ( n54572 , n232331 , n232332 );
not ( n54573 , n54572 );
and ( n54574 , n54562 , n54573 );
not ( n54575 , n54562 );
and ( n232337 , n54575 , n54572 );
nor ( n232338 , n54574 , n232337 );
not ( n54578 , n232338 );
not ( n54579 , n54578 );
buf ( n54580 , n28236 );
not ( n54581 , n54580 );
not ( n232343 , n36243 );
or ( n232344 , n54581 , n232343 );
or ( n54584 , n36243 , n54580 );
nand ( n54585 , n232344 , n54584 );
not ( n54586 , n54585 );
not ( n54587 , n45218 );
and ( n232349 , n54586 , n54587 );
buf ( n232350 , n48058 );
and ( n54590 , n54585 , n232350 );
nor ( n232352 , n232349 , n54590 );
not ( n232353 , n232352 );
not ( n54593 , n232353 );
buf ( n54594 , n205122 );
xor ( n54595 , n54594 , n41411 );
xor ( n54596 , n54595 , n34759 );
not ( n54597 , n54596 );
not ( n54598 , n29265 );
not ( n54599 , n44347 );
or ( n54600 , n54598 , n54599 );
or ( n54601 , n44347 , n29265 );
nand ( n54602 , n54600 , n54601 );
and ( n54603 , n54602 , n40697 );
not ( n232365 , n54602 );
and ( n232366 , n232365 , n205420 );
nor ( n232367 , n54603 , n232366 );
not ( n232368 , n232367 );
nand ( n54608 , n54597 , n232368 );
not ( n54609 , n54608 );
or ( n54610 , n54593 , n54609 );
or ( n54611 , n54608 , n232353 );
nand ( n232373 , n54610 , n54611 );
not ( n232374 , n232373 );
not ( n54614 , n232374 );
xor ( n54615 , n34556 , n44158 );
xnor ( n54616 , n54615 , n47330 );
not ( n54617 , n54616 );
not ( n232379 , n28691 );
not ( n232380 , n32962 );
or ( n54620 , n232379 , n232380 );
or ( n54621 , n32962 , n28691 );
nand ( n54622 , n54620 , n54621 );
buf ( n54623 , n225593 );
and ( n232385 , n54622 , n54623 );
not ( n232386 , n54622 );
and ( n54626 , n232386 , n32989 );
nor ( n54627 , n232385 , n54626 );
nand ( n54628 , n54617 , n54627 );
not ( n54629 , n54628 );
buf ( n232391 , RI174a4b50_933);
and ( n232392 , n28966 , n232391 );
not ( n54632 , n28966 );
and ( n54633 , n54632 , n28963 );
nor ( n54634 , n232392 , n54633 );
xor ( n54635 , n54634 , n30321 );
not ( n232397 , n54635 );
not ( n232398 , n204436 );
and ( n54638 , n232397 , n232398 );
and ( n54639 , n54635 , n48521 );
nor ( n54640 , n54638 , n54639 );
not ( n54641 , n54640 );
not ( n232403 , n54641 );
and ( n232404 , n54629 , n232403 );
and ( n54644 , n54628 , n54641 );
nor ( n54645 , n232404 , n54644 );
not ( n54646 , n54645 );
not ( n54647 , n54646 );
or ( n232409 , n54614 , n54647 );
nand ( n232410 , n54645 , n232373 );
nand ( n54650 , n232409 , n232410 );
not ( n232412 , n54650 );
not ( n232413 , n232412 );
not ( n54653 , n39569 );
not ( n54654 , n32781 );
not ( n54655 , n26143 );
and ( n54656 , n54654 , n54655 );
not ( n232418 , n26144 );
and ( n232419 , n32781 , n232418 );
nor ( n54659 , n54656 , n232419 );
not ( n54660 , n54659 );
or ( n54661 , n54653 , n54660 );
or ( n54662 , n54659 , n39569 );
nand ( n54663 , n54661 , n54662 );
not ( n54664 , n54663 );
xor ( n232426 , n39910 , n39919 );
xor ( n232427 , n232426 , n25637 );
not ( n54667 , n232427 );
not ( n54668 , n54667 );
not ( n54669 , n208380 );
and ( n54670 , n54668 , n54669 );
and ( n232432 , n39922 , n208380 );
nor ( n232433 , n54670 , n232432 );
and ( n54673 , n232433 , n47607 );
not ( n232435 , n232433 );
and ( n232436 , n232435 , n47612 );
nor ( n54676 , n54673 , n232436 );
nand ( n54677 , n54664 , n54676 );
not ( n54678 , n54677 );
not ( n54679 , n40051 );
not ( n232441 , n30942 );
or ( n232442 , n54679 , n232441 );
or ( n54682 , n30942 , n40051 );
nand ( n232444 , n232442 , n54682 );
xor ( n232445 , n232444 , n221779 );
not ( n54685 , n232445 );
not ( n232447 , n54685 );
and ( n232448 , n54678 , n232447 );
and ( n54688 , n54677 , n54685 );
nor ( n54689 , n232448 , n54688 );
not ( n54690 , n54689 );
not ( n54691 , n45139 );
not ( n54692 , n229404 );
not ( n232454 , n54692 );
not ( n232455 , n40772 );
or ( n54695 , n232454 , n232455 );
or ( n54696 , n40772 , n54692 );
nand ( n54697 , n54695 , n54696 );
not ( n54698 , n54697 );
and ( n54699 , n54691 , n54698 );
and ( n232461 , n40813 , n54697 );
nor ( n232462 , n54699 , n232461 );
not ( n54702 , n39833 );
not ( n54703 , n38188 );
or ( n54704 , n54702 , n54703 );
nand ( n54705 , n38201 , n39829 );
nand ( n54706 , n54704 , n54705 );
not ( n54707 , n54706 );
not ( n54708 , n38205 );
and ( n232470 , n54707 , n54708 );
and ( n232471 , n54706 , n38205 );
nor ( n54711 , n232470 , n232471 );
not ( n54712 , n54711 );
nand ( n54713 , n232462 , n54712 );
buf ( n54714 , n205067 );
and ( n232476 , n54714 , n28251 );
not ( n232477 , n54714 );
and ( n54717 , n232477 , n28247 );
nor ( n54718 , n232476 , n54717 );
not ( n54719 , n54718 );
not ( n54720 , n54719 );
not ( n232482 , n209844 );
or ( n232483 , n54720 , n232482 );
nand ( n54723 , n32082 , n54718 );
nand ( n54724 , n232483 , n54723 );
not ( n54725 , n54724 );
and ( n54726 , n54713 , n54725 );
not ( n232488 , n54713 );
and ( n232489 , n232488 , n54724 );
nor ( n54729 , n54726 , n232489 );
not ( n54730 , n54729 );
or ( n54731 , n54690 , n54730 );
or ( n54732 , n54729 , n54689 );
nand ( n54733 , n54731 , n54732 );
nand ( n54734 , n54549 , n54573 );
buf ( n232496 , n204334 );
not ( n232497 , n232496 );
not ( n54737 , n37762 );
or ( n54738 , n232497 , n54737 );
or ( n54739 , n37762 , n232496 );
nand ( n54740 , n54738 , n54739 );
xnor ( n232502 , n54740 , n33886 );
not ( n232503 , n232502 );
xor ( n54743 , n54734 , n232503 );
not ( n54744 , n54743 );
and ( n54745 , n54733 , n54744 );
not ( n54746 , n54733 );
and ( n54747 , n54746 , n54743 );
nor ( n54748 , n54745 , n54747 );
not ( n54749 , n54748 );
not ( n54750 , n54749 );
or ( n232512 , n232413 , n54750 );
nand ( n232513 , n54748 , n54650 );
nand ( n232514 , n232512 , n232513 );
not ( n232515 , n232514 );
or ( n54755 , n54579 , n232515 );
and ( n232517 , n54748 , n54650 );
not ( n232518 , n54748 );
and ( n54758 , n232518 , n232412 );
nor ( n232520 , n232517 , n54758 );
nand ( n232521 , n232520 , n232338 );
nand ( n54761 , n54755 , n232521 );
not ( n232523 , n54761 );
and ( n232524 , n232300 , n232523 );
and ( n54764 , n232299 , n54761 );
nor ( n54765 , n232524 , n54764 );
not ( n232527 , n54765 );
not ( n232528 , n45070 );
nand ( n54768 , n232528 , n222852 );
not ( n54769 , n27833 );
not ( n54770 , n33756 );
or ( n54771 , n54769 , n54770 );
nand ( n54772 , n227018 , n27829 );
nand ( n54773 , n54771 , n54772 );
and ( n54774 , n54773 , n33764 );
not ( n54775 , n54773 );
and ( n232537 , n54775 , n31253 );
nor ( n232538 , n54774 , n232537 );
and ( n54778 , n54768 , n232538 );
not ( n54779 , n54768 );
not ( n54780 , n232538 );
and ( n54781 , n54779 , n54780 );
nor ( n232543 , n54778 , n54781 );
not ( n232544 , n232543 );
not ( n54784 , n47450 );
buf ( n54785 , RI17334bb8_2184);
not ( n54786 , n54785 );
not ( n54787 , n47816 );
or ( n232549 , n54786 , n54787 );
nand ( n232550 , n45464 , n30794 );
nand ( n54790 , n232549 , n232550 );
not ( n54791 , n54790 );
or ( n54792 , n54784 , n54791 );
or ( n54793 , n54790 , n229281 );
nand ( n232555 , n54792 , n54793 );
buf ( n232556 , n232555 );
not ( n54796 , n232556 );
not ( n232558 , n53511 );
and ( n232559 , n35432 , n53500 );
not ( n54799 , n35432 );
and ( n232561 , n54799 , n31037 );
nor ( n232562 , n232559 , n232561 );
not ( n54802 , n232562 );
and ( n54803 , n232558 , n54802 );
and ( n54804 , n31078 , n232562 );
nor ( n54805 , n54803 , n54804 );
nand ( n232567 , n54805 , n45142 );
not ( n232568 , n232567 );
or ( n54808 , n54796 , n232568 );
or ( n54809 , n232567 , n232556 );
nand ( n54810 , n54808 , n54809 );
not ( n54811 , n54810 );
not ( n232573 , n41265 );
not ( n232574 , n34589 );
or ( n54814 , n232573 , n232574 );
or ( n54815 , n29733 , n41265 );
nand ( n54816 , n54814 , n54815 );
and ( n54817 , n54816 , n34594 );
not ( n232579 , n54816 );
and ( n232580 , n232579 , n34598 );
nor ( n54820 , n54817 , n232580 );
not ( n232582 , n54820 );
nand ( n232583 , n222939 , n232582 );
not ( n54823 , n232583 );
not ( n54824 , n38177 );
not ( n54825 , n34088 );
or ( n54826 , n54824 , n54825 );
or ( n232588 , n34088 , n38177 );
nand ( n232589 , n54826 , n232588 );
and ( n54829 , n232589 , n40369 );
not ( n54830 , n232589 );
and ( n54831 , n54830 , n40370 );
nor ( n54832 , n54829 , n54831 );
not ( n232594 , n54832 );
not ( n232595 , n232594 );
and ( n54835 , n54823 , n232595 );
and ( n54836 , n232583 , n232594 );
nor ( n54837 , n54835 , n54836 );
not ( n54838 , n54837 );
or ( n232600 , n54811 , n54838 );
or ( n232601 , n54837 , n54810 );
nand ( n54841 , n232600 , n232601 );
not ( n54842 , n32667 );
not ( n54843 , n48308 );
or ( n54844 , n54842 , n54843 );
not ( n232606 , n32667 );
nand ( n232607 , n232606 , n48312 );
nand ( n54847 , n54844 , n232607 );
not ( n54848 , n37996 );
not ( n54849 , n54848 );
and ( n54850 , n54847 , n54849 );
not ( n54851 , n54847 );
and ( n54852 , n54851 , n48317 );
nor ( n54853 , n54850 , n54852 );
not ( n54854 , n54853 );
nand ( n54855 , n45242 , n54854 );
not ( n232617 , n54855 );
not ( n232618 , n37507 );
not ( n54858 , n30755 );
not ( n54859 , n31636 );
or ( n54860 , n54858 , n54859 );
not ( n54861 , n30755 );
nand ( n232623 , n54861 , n37488 );
nand ( n232624 , n54860 , n232623 );
not ( n54864 , n232624 );
and ( n232626 , n232618 , n54864 );
and ( n232627 , n37507 , n232624 );
nor ( n54867 , n232626 , n232627 );
not ( n54868 , n54867 );
not ( n54869 , n54868 );
and ( n54870 , n232617 , n54869 );
and ( n54871 , n54855 , n54868 );
nor ( n232633 , n54870 , n54871 );
and ( n232634 , n54841 , n232633 );
not ( n54874 , n54841 );
not ( n54875 , n232633 );
and ( n54876 , n54874 , n54875 );
nor ( n54877 , n232634 , n54876 );
xor ( n232639 , n36847 , n42624 );
xnor ( n232640 , n232639 , n224874 );
not ( n54880 , n232640 );
not ( n54881 , n54880 );
not ( n232643 , n29132 );
not ( n232644 , n39401 );
or ( n54884 , n232643 , n232644 );
nand ( n54885 , n45898 , n29128 );
nand ( n54886 , n54884 , n54885 );
and ( n54887 , n54886 , n51252 );
not ( n232649 , n54886 );
and ( n232650 , n232649 , n223859 );
nor ( n54890 , n54887 , n232650 );
nor ( n54891 , n45038 , n54890 );
not ( n54892 , n54891 );
and ( n54893 , n54881 , n54892 );
and ( n232655 , n54891 , n54880 );
nor ( n232656 , n54893 , n232655 );
not ( n54896 , n232656 );
not ( n232658 , n54896 );
nand ( n232659 , n232538 , n45092 );
not ( n54899 , n232659 );
not ( n54900 , n31322 );
xor ( n54901 , n54900 , n51033 );
xnor ( n54902 , n54901 , n28122 );
not ( n232664 , n54902 );
not ( n232665 , n232664 );
or ( n54905 , n54899 , n232665 );
or ( n54906 , n232664 , n232659 );
nand ( n54907 , n54905 , n54906 );
not ( n54908 , n54907 );
not ( n232670 , n54908 );
or ( n232671 , n232658 , n232670 );
nand ( n54911 , n54907 , n232656 );
nand ( n54912 , n232671 , n54911 );
and ( n54913 , n54877 , n54912 );
not ( n54914 , n54877 );
not ( n232676 , n54912 );
and ( n232677 , n54914 , n232676 );
nor ( n54917 , n54913 , n232677 );
not ( n54918 , n54917 );
or ( n54919 , n232544 , n54918 );
not ( n54920 , n232543 );
not ( n232682 , n232676 );
not ( n232683 , n54877 );
not ( n54923 , n232683 );
or ( n54924 , n232682 , n54923 );
nand ( n54925 , n54877 , n54912 );
nand ( n54926 , n54924 , n54925 );
nand ( n54927 , n54920 , n54926 );
nand ( n232689 , n54919 , n54927 );
not ( n232690 , n43260 );
not ( n232691 , n42948 );
and ( n232692 , n232690 , n232691 );
and ( n54932 , n43260 , n42948 );
nor ( n232694 , n232692 , n54932 );
and ( n232695 , n232694 , n220435 );
not ( n54935 , n232694 );
and ( n232697 , n54935 , n220432 );
nor ( n232698 , n232695 , n232697 );
not ( n54938 , n232698 );
nand ( n54939 , n54938 , n232502 );
not ( n54940 , n54939 );
not ( n54941 , n54561 );
and ( n232703 , n54940 , n54941 );
and ( n232704 , n54939 , n54561 );
nor ( n54944 , n232703 , n232704 );
not ( n54945 , n54944 );
not ( n232707 , n28665 );
not ( n232708 , n29613 );
not ( n54948 , n221233 );
or ( n54949 , n232708 , n54948 );
or ( n54950 , n221233 , n29613 );
nand ( n54951 , n54949 , n54950 );
not ( n232713 , n54951 );
and ( n232714 , n232707 , n232713 );
and ( n54954 , n28665 , n54951 );
nor ( n54955 , n232714 , n54954 );
not ( n54956 , n54955 );
not ( n54957 , n54956 );
xor ( n232719 , n44391 , n40568 );
xnor ( n232720 , n232719 , n29518 );
not ( n54960 , n232720 );
nand ( n54961 , n54960 , n54724 );
not ( n54962 , n54961 );
or ( n54963 , n54957 , n54962 );
or ( n232725 , n54961 , n54956 );
nand ( n232726 , n54963 , n232725 );
not ( n54966 , n232726 );
or ( n232728 , n54945 , n54966 );
or ( n232729 , n54944 , n232726 );
nand ( n54969 , n232728 , n232729 );
not ( n54970 , n28319 );
not ( n54971 , n36309 );
or ( n54972 , n54970 , n54971 );
not ( n232734 , n28319 );
nand ( n232735 , n232734 , n36308 );
nand ( n54975 , n54972 , n232735 );
and ( n54976 , n54975 , n36350 );
not ( n54977 , n54975 );
and ( n54978 , n54977 , n36349 );
nor ( n232740 , n54976 , n54978 );
nand ( n232741 , n232740 , n54685 );
not ( n54981 , n232741 );
not ( n54982 , n37624 );
not ( n54983 , n31136 );
or ( n54984 , n54982 , n54983 );
or ( n232746 , n31136 , n37624 );
nand ( n232747 , n54984 , n232746 );
and ( n54987 , n232747 , n29733 );
not ( n232749 , n232747 );
and ( n54989 , n232749 , n207493 );
nor ( n54990 , n54987 , n54989 );
not ( n54991 , n54990 );
not ( n54992 , n54991 );
and ( n54993 , n54981 , n54992 );
and ( n54994 , n232741 , n54991 );
nor ( n232756 , n54993 , n54994 );
and ( n232757 , n54969 , n232756 );
not ( n54997 , n54969 );
not ( n54998 , n232756 );
and ( n54999 , n54997 , n54998 );
nor ( n55000 , n232757 , n54999 );
not ( n232762 , n40935 );
not ( n232763 , n30985 );
not ( n55003 , n43553 );
or ( n55004 , n232763 , n55003 );
not ( n55005 , n30985 );
nand ( n55006 , n55005 , n50185 );
nand ( n55007 , n55004 , n55006 );
not ( n55008 , n55007 );
or ( n55009 , n232762 , n55008 );
or ( n55010 , n40935 , n55007 );
nand ( n55011 , n55009 , n55010 );
not ( n232773 , n55011 );
nand ( n232774 , n232773 , n54641 );
not ( n232775 , n33580 );
not ( n232776 , n40414 );
or ( n55016 , n232775 , n232776 );
or ( n232778 , n44239 , n33580 );
nand ( n232779 , n55016 , n232778 );
not ( n55019 , n232779 );
not ( n55020 , n32284 );
and ( n55021 , n55019 , n55020 );
and ( n55022 , n232779 , n32280 );
nor ( n232784 , n55021 , n55022 );
not ( n232785 , n232784 );
and ( n55025 , n232774 , n232785 );
not ( n55026 , n232774 );
and ( n55027 , n55026 , n232784 );
nor ( n55028 , n55025 , n55027 );
not ( n232790 , n55028 );
not ( n232791 , n232790 );
not ( n55031 , n32378 );
not ( n55032 , n36187 );
or ( n55033 , n55031 , n55032 );
or ( n55034 , n36187 , n32378 );
nand ( n232796 , n55033 , n55034 );
not ( n232797 , n225166 );
and ( n55037 , n232796 , n232797 );
not ( n55038 , n232796 );
and ( n55039 , n55038 , n225166 );
nor ( n55040 , n55037 , n55039 );
not ( n232802 , n55040 );
nand ( n232803 , n232802 , n232353 );
not ( n55043 , n29107 );
not ( n55044 , n36262 );
or ( n55045 , n55043 , n55044 );
nand ( n55046 , n32827 , n29103 );
nand ( n55047 , n55045 , n55046 );
and ( n55048 , n55047 , n39402 );
not ( n232810 , n55047 );
and ( n232811 , n232810 , n45898 );
nor ( n232812 , n55048 , n232811 );
and ( n232813 , n232803 , n232812 );
not ( n55053 , n232803 );
not ( n232815 , n232812 );
and ( n232816 , n55053 , n232815 );
nor ( n55056 , n232813 , n232816 );
not ( n232818 , n55056 );
not ( n232819 , n232818 );
or ( n55059 , n232791 , n232819 );
nand ( n55060 , n55056 , n55028 );
nand ( n55061 , n55059 , n55060 );
not ( n55062 , n55061 );
and ( n55063 , n55000 , n55062 );
not ( n232825 , n55000 );
and ( n232826 , n232825 , n55061 );
nor ( n55066 , n55063 , n232826 );
not ( n55067 , n55066 );
buf ( n55068 , n55067 );
xnor ( n55069 , n232689 , n55068 );
not ( n55070 , n55069 );
or ( n55071 , n232527 , n55070 );
not ( n232833 , n32023 );
not ( n232834 , n38674 );
or ( n55074 , n232833 , n232834 );
or ( n55075 , n38674 , n32023 );
nand ( n55076 , n55074 , n55075 );
not ( n55077 , n55076 );
not ( n232839 , n38670 );
not ( n232840 , n232839 );
or ( n55080 , n55077 , n232840 );
or ( n55081 , n232839 , n55076 );
nand ( n55082 , n55080 , n55081 );
and ( n55083 , n55082 , n36684 );
not ( n232845 , n55082 );
and ( n232846 , n232845 , n31176 );
nor ( n55086 , n55083 , n232846 );
nand ( n55087 , n55086 , n47868 );
not ( n55088 , n55087 );
not ( n55089 , n48585 );
and ( n232851 , n55088 , n55089 );
and ( n232852 , n55087 , n48585 );
nor ( n55092 , n232851 , n232852 );
not ( n55093 , n55092 );
not ( n55094 , n48015 );
or ( n55095 , n55093 , n55094 );
not ( n232857 , n55092 );
nand ( n232858 , n232857 , n48019 );
nand ( n55098 , n55095 , n232858 );
not ( n55099 , n55098 );
not ( n55100 , n48238 );
and ( n55101 , n55099 , n55100 );
and ( n232863 , n55098 , n48233 );
nor ( n232864 , n55101 , n232863 );
buf ( n55104 , n37724 );
nor ( n55105 , n232864 , n55104 );
nand ( n55106 , n55071 , n55105 );
not ( n55107 , n54765 );
not ( n55108 , n226010 );
nor ( n232870 , n55107 , n55108 );
nand ( n232871 , n232870 , n232864 , n55069 );
nand ( n55111 , n31577 , n38903 );
nand ( n55112 , n55106 , n232871 , n55111 );
buf ( n55113 , n55112 );
not ( n55114 , n46566 );
xor ( n232876 , n35689 , n35693 );
xor ( n232877 , n232876 , n35702 );
not ( n55117 , n232877 );
or ( n55118 , n55114 , n55117 );
or ( n55119 , n232877 , n46566 );
nand ( n55120 , n55118 , n55119 );
and ( n55121 , n55120 , n25762 );
not ( n232883 , n55120 );
and ( n232884 , n232883 , n25765 );
nor ( n55124 , n55121 , n232884 );
not ( n55125 , n55124 );
nand ( n232887 , n55125 , n37139 );
not ( n232888 , n232887 );
not ( n55128 , n37130 );
not ( n55129 , n55128 );
and ( n55130 , n232888 , n55129 );
and ( n55131 , n232887 , n55128 );
nor ( n232893 , n55130 , n55131 );
not ( n232894 , n232893 );
not ( n55134 , n232894 );
not ( n55135 , n37288 );
not ( n55136 , n55135 );
or ( n55137 , n55134 , n55136 );
buf ( n232899 , n37288 );
not ( n232900 , n232899 );
or ( n55140 , n232900 , n232894 );
nand ( n55141 , n55137 , n55140 );
and ( n55142 , n55141 , n37715 );
not ( n55143 , n55141 );
and ( n232905 , n55143 , n37709 );
nor ( n232906 , n55142 , n232905 );
buf ( n55146 , n35427 );
not ( n55147 , n55146 );
nand ( n55148 , n232906 , n55147 );
not ( n55149 , n39757 );
nand ( n232911 , n39447 , n55149 );
or ( n232912 , n55148 , n232911 );
buf ( n55152 , n226003 );
nor ( n232914 , n232906 , n55152 );
nand ( n232915 , n232914 , n232911 );
nand ( n55155 , n49054 , n33497 );
nand ( n55156 , n232912 , n232915 , n55155 );
buf ( n55157 , n55156 );
not ( n55158 , n41491 );
not ( n55159 , n219315 );
not ( n55160 , n41530 );
nand ( n232922 , n55159 , n55160 );
not ( n232923 , n232922 );
not ( n55163 , n32219 );
nor ( n55164 , n28829 , n39609 );
not ( n55165 , n55164 );
nand ( n55166 , n28829 , n39609 );
nand ( n55167 , n55165 , n55166 );
not ( n232929 , n55167 );
and ( n232930 , n55163 , n232929 );
and ( n55170 , n32219 , n55167 );
nor ( n55171 , n232930 , n55170 );
not ( n55172 , n55171 );
not ( n55173 , n55172 );
and ( n232935 , n232923 , n55173 );
and ( n232936 , n232922 , n55172 );
nor ( n55176 , n232935 , n232936 );
not ( n55177 , n55176 );
not ( n55178 , n41617 );
nand ( n55179 , n55178 , n41589 );
not ( n232941 , n30100 );
not ( n232942 , n32795 );
not ( n55182 , n30078 );
or ( n55183 , n232942 , n55182 );
or ( n55184 , n30078 , n32795 );
nand ( n55185 , n55183 , n55184 );
not ( n232947 , n55185 );
and ( n232948 , n232941 , n232947 );
and ( n55188 , n30100 , n55185 );
nor ( n55189 , n232948 , n55188 );
and ( n55190 , n55179 , n55189 );
not ( n55191 , n55179 );
not ( n232953 , n55189 );
and ( n232954 , n55191 , n232953 );
nor ( n55194 , n55190 , n232954 );
not ( n232956 , n55194 );
or ( n232957 , n55177 , n232956 );
or ( n55197 , n55194 , n55176 );
nand ( n55198 , n232957 , n55197 );
not ( n55199 , n41573 );
nand ( n55200 , n55199 , n41364 );
not ( n232962 , n204407 );
not ( n232963 , n218917 );
or ( n55203 , n232962 , n232963 );
not ( n55204 , n204407 );
nand ( n55205 , n55204 , n37120 );
nand ( n55206 , n55203 , n55205 );
and ( n232968 , n55206 , n37128 );
not ( n232969 , n55206 );
and ( n55209 , n232969 , n37123 );
nor ( n232971 , n232968 , n55209 );
not ( n232972 , n232971 );
xor ( n55212 , n55200 , n232972 );
not ( n55213 , n55212 );
and ( n55214 , n55198 , n55213 );
not ( n55215 , n55198 );
and ( n232977 , n55215 , n55212 );
nor ( n232978 , n55214 , n232977 );
not ( n55218 , n41475 );
nand ( n55219 , n41487 , n55218 );
not ( n55220 , n52256 );
not ( n55221 , n45190 );
not ( n232983 , n49483 );
or ( n232984 , n55221 , n232983 );
not ( n55224 , n28344 );
or ( n55225 , n55224 , n45190 );
nand ( n55226 , n232984 , n55225 );
not ( n55227 , n55226 );
or ( n232989 , n55220 , n55227 );
or ( n232990 , n55226 , n28382 );
nand ( n55230 , n232989 , n232990 );
and ( n55231 , n55219 , n55230 );
not ( n55232 , n55219 );
not ( n55233 , n55230 );
and ( n232995 , n55232 , n55233 );
or ( n232996 , n55231 , n232995 );
not ( n55236 , n232996 );
not ( n232998 , n41381 );
nand ( n232999 , n41419 , n232998 );
not ( n55239 , n33975 );
not ( n55240 , n39207 );
or ( n55241 , n55239 , n55240 );
not ( n55242 , n39207 );
nand ( n55243 , n55242 , n33971 );
nand ( n55244 , n55241 , n55243 );
and ( n55245 , n55244 , n39251 );
not ( n55246 , n55244 );
buf ( n233008 , n45933 );
and ( n233009 , n55246 , n233008 );
nor ( n55249 , n55245 , n233009 );
not ( n55250 , n55249 );
and ( n55251 , n232999 , n55250 );
not ( n55252 , n232999 );
and ( n233014 , n55252 , n55249 );
nor ( n233015 , n55251 , n233014 );
not ( n55255 , n233015 );
not ( n55256 , n55255 );
or ( n55257 , n55236 , n55256 );
not ( n55258 , n232996 );
nand ( n233020 , n55258 , n233015 );
nand ( n233021 , n55257 , n233020 );
and ( n55261 , n232978 , n233021 );
not ( n55262 , n232978 );
not ( n55263 , n233021 );
and ( n55264 , n55262 , n55263 );
nor ( n233026 , n55261 , n55264 );
not ( n233027 , n233026 );
or ( n55267 , n55158 , n233027 );
not ( n55268 , n41491 );
not ( n55269 , n233021 );
not ( n55270 , n232978 );
or ( n55271 , n55269 , n55270 );
not ( n55272 , n232978 );
nand ( n233034 , n55272 , n55263 );
nand ( n233035 , n55271 , n233034 );
nand ( n55275 , n55268 , n233035 );
nand ( n55276 , n55267 , n55275 );
not ( n55277 , n219824 );
nand ( n55278 , n41805 , n41789 );
not ( n233040 , n55278 );
or ( n233041 , n55277 , n233040 );
or ( n55281 , n55278 , n219824 );
nand ( n233043 , n233041 , n55281 );
not ( n233044 , n233043 );
nand ( n55284 , n41880 , n41828 );
not ( n233046 , n55284 );
not ( n233047 , n219881 );
and ( n55287 , n233046 , n233047 );
and ( n55288 , n55284 , n219881 );
nor ( n55289 , n55287 , n55288 );
not ( n55290 , n55289 );
or ( n233052 , n233044 , n55290 );
or ( n233053 , n55289 , n233043 );
nand ( n55293 , n233052 , n233053 );
not ( n55294 , n55293 );
not ( n55295 , n41892 );
nand ( n55296 , n55295 , n41912 );
and ( n233058 , n55296 , n53034 );
not ( n233059 , n55296 );
and ( n55299 , n233059 , n42099 );
nor ( n55300 , n233058 , n55299 );
not ( n55301 , n55300 );
not ( n55302 , n55301 );
or ( n55303 , n55294 , n55302 );
not ( n55304 , n55293 );
nand ( n233066 , n55304 , n55300 );
nand ( n233067 , n55303 , n233066 );
not ( n55307 , n230785 );
not ( n55308 , n41768 );
not ( n55309 , n41683 );
nand ( n55310 , n55308 , n55309 );
not ( n233072 , n55310 );
not ( n233073 , n41996 );
and ( n55313 , n233072 , n233073 );
and ( n55314 , n55310 , n41996 );
nor ( n55315 , n55313 , n55314 );
not ( n55316 , n55315 );
not ( n233078 , n55316 );
or ( n233079 , n55307 , n233078 );
nand ( n55319 , n53023 , n55315 );
nand ( n55320 , n233079 , n55319 );
not ( n55321 , n55320 );
xnor ( n55322 , n233067 , n55321 );
buf ( n233084 , n55322 );
and ( n233085 , n55276 , n233084 );
not ( n55325 , n55276 );
and ( n55326 , n233067 , n55321 );
not ( n55327 , n233067 );
and ( n55328 , n55327 , n55320 );
nor ( n233090 , n55326 , n55328 );
buf ( n233091 , n233090 );
and ( n55331 , n55325 , n233091 );
nor ( n55332 , n233085 , n55331 );
not ( n55333 , n55332 );
nand ( n55334 , n206427 , n28682 );
not ( n233096 , n55334 );
buf ( n233097 , n33669 );
not ( n55337 , n233097 );
and ( n55338 , n233096 , n55337 );
and ( n55339 , n55334 , n233097 );
nor ( n55340 , n55338 , n55339 );
not ( n233102 , n55340 );
and ( n233103 , n33489 , n33706 );
not ( n55343 , n33489 );
and ( n55344 , n55343 , n33703 );
nor ( n55345 , n233103 , n55344 );
not ( n55346 , n55345 );
or ( n233108 , n233102 , n55346 );
not ( n233109 , n55340 );
nand ( n55349 , n233109 , n33708 );
nand ( n55350 , n233108 , n55349 );
not ( n55351 , n30471 );
not ( n55352 , n54399 );
or ( n233114 , n55351 , n55352 );
or ( n233115 , n54402 , n30471 );
nand ( n55355 , n233114 , n233115 );
and ( n55356 , n55355 , n33229 );
not ( n55357 , n55355 );
and ( n55358 , n55357 , n33230 );
nor ( n233120 , n55356 , n55358 );
not ( n233121 , n233120 );
not ( n55361 , n233121 );
buf ( n55362 , n32565 );
not ( n55363 , n55362 );
not ( n55364 , n55363 );
not ( n233126 , n28463 );
or ( n233127 , n55364 , n233126 );
nand ( n55367 , n28466 , n55362 );
nand ( n55368 , n233127 , n55367 );
and ( n55369 , n55368 , n28511 );
not ( n55370 , n55368 );
and ( n233132 , n55370 , n28503 );
nor ( n233133 , n55369 , n233132 );
nor ( n55373 , n29950 , n233133 );
not ( n55374 , n55373 );
and ( n55375 , n55361 , n55374 );
and ( n55376 , n233121 , n55373 );
nor ( n233138 , n55375 , n55376 );
not ( n233139 , n233138 );
buf ( n55379 , n34373 );
not ( n55380 , n55379 );
not ( n55381 , n37020 );
or ( n55382 , n55380 , n55381 );
not ( n233144 , n55379 );
nand ( n233145 , n233144 , n37023 );
nand ( n55385 , n55382 , n233145 );
and ( n55386 , n55385 , n45770 );
not ( n55387 , n55385 );
and ( n55388 , n55387 , n223536 );
nor ( n233150 , n55386 , n55388 );
nand ( n233151 , n29738 , n233150 );
not ( n55391 , n40837 );
not ( n55392 , n44633 );
or ( n55393 , n55391 , n55392 );
nand ( n55394 , n45944 , n40840 );
nand ( n233156 , n55393 , n55394 );
and ( n233157 , n233156 , n42966 );
not ( n55397 , n233156 );
and ( n233159 , n55397 , n38657 );
nor ( n233160 , n233157 , n233159 );
not ( n55400 , n233160 );
and ( n55401 , n233151 , n55400 );
not ( n55402 , n233151 );
and ( n55403 , n55402 , n233160 );
nor ( n233165 , n55401 , n55403 );
not ( n233166 , n233165 );
and ( n55406 , n233139 , n233166 );
and ( n55407 , n233138 , n233165 );
nor ( n55408 , n55406 , n55407 );
not ( n55409 , n55408 );
not ( n55410 , n32218 );
xor ( n55411 , n36962 , n55410 );
xor ( n55412 , n55411 , n32240 );
not ( n55413 , n55412 );
not ( n55414 , n29341 );
nand ( n55415 , n55413 , n55414 );
not ( n233177 , n55415 );
not ( n233178 , n45199 );
not ( n55418 , n49483 );
or ( n55419 , n233178 , n55418 );
or ( n55420 , n49483 , n45199 );
nand ( n55421 , n55419 , n55420 );
and ( n55422 , n55421 , n52256 );
not ( n55423 , n55421 );
and ( n233185 , n55423 , n49491 );
nor ( n233186 , n55422 , n233185 );
not ( n55426 , n233186 );
not ( n233188 , n55426 );
and ( n233189 , n233177 , n233188 );
nand ( n55429 , n55413 , n29342 );
and ( n233191 , n55429 , n55426 );
nor ( n233192 , n233189 , n233191 );
not ( n55432 , n233192 );
not ( n55433 , n37221 );
not ( n55434 , RI173f22c0_1575);
not ( n55435 , n207999 );
xor ( n233197 , n55434 , n55435 );
xnor ( n233198 , n233197 , n30245 );
not ( n55438 , n233198 );
or ( n55439 , n55433 , n55438 );
not ( n55440 , n37221 );
not ( n55441 , n233198 );
nand ( n233203 , n55440 , n55441 );
nand ( n233204 , n55439 , n233203 );
and ( n55444 , n233204 , n41411 );
not ( n233206 , n233204 );
not ( n233207 , n41411 );
and ( n55447 , n233206 , n233207 );
nor ( n55448 , n55444 , n55447 );
not ( n55449 , n55448 );
nand ( n55450 , n55449 , n28949 );
not ( n233212 , n47450 );
not ( n233213 , n30783 );
not ( n55453 , n45464 );
or ( n55454 , n233213 , n55453 );
buf ( n55455 , RI174122a0_1419);
nand ( n55456 , n47816 , n55455 );
nand ( n233218 , n55454 , n55456 );
not ( n233219 , n233218 );
or ( n55459 , n233212 , n233219 );
or ( n55460 , n233218 , n47450 );
nand ( n55461 , n55459 , n55460 );
buf ( n55462 , n55461 );
not ( n233224 , n55462 );
and ( n233225 , n55450 , n233224 );
not ( n55465 , n55450 );
and ( n55466 , n55465 , n55462 );
nor ( n55467 , n233225 , n55466 );
not ( n55468 , n55467 );
or ( n233230 , n55432 , n55468 );
or ( n233231 , n55467 , n233192 );
nand ( n55471 , n233230 , n233231 );
xor ( n233233 , n36337 , n41894 );
xnor ( n233234 , n233233 , n31078 );
not ( n55474 , n233234 );
nand ( n55475 , n55474 , n29473 );
buf ( n55476 , RI17450028_1346);
not ( n55477 , n55476 );
not ( n233239 , n35861 );
or ( n233240 , n55477 , n233239 );
not ( n55480 , n222752 );
not ( n55481 , n55480 );
or ( n55482 , n55481 , n55476 );
nand ( n55483 , n233240 , n55482 );
and ( n233245 , n55483 , n37539 );
not ( n233246 , n55483 );
and ( n55486 , n233246 , n37533 );
nor ( n55487 , n233245 , n55486 );
not ( n55488 , n55487 );
and ( n55489 , n55475 , n55488 );
not ( n233251 , n55475 );
and ( n233252 , n233251 , n55487 );
nor ( n55492 , n55489 , n233252 );
and ( n55493 , n55471 , n55492 );
not ( n55494 , n55471 );
not ( n55495 , n55492 );
and ( n55496 , n55494 , n55495 );
nor ( n233258 , n55493 , n55496 );
not ( n233259 , n233258 );
or ( n55499 , n55409 , n233259 );
not ( n55500 , n233258 );
not ( n55501 , n55408 );
nand ( n55502 , n55500 , n55501 );
nand ( n233264 , n55499 , n55502 );
buf ( n233265 , n233264 );
and ( n55505 , n55350 , n233265 );
not ( n55506 , n55350 );
and ( n55507 , n55500 , n55501 );
not ( n55508 , n55500 );
and ( n233270 , n55508 , n55408 );
nor ( n233271 , n55507 , n233270 );
buf ( n55511 , n233271 );
and ( n55512 , n55506 , n55511 );
nor ( n55513 , n55505 , n55512 );
not ( n55514 , n55513 );
not ( n233276 , n55514 );
or ( n233277 , n55333 , n233276 );
not ( n55517 , n205397 );
not ( n55518 , n228364 );
or ( n55519 , n55517 , n55518 );
not ( n55520 , n205397 );
nand ( n233282 , n55520 , n50539 );
nand ( n233283 , n55519 , n233282 );
and ( n55523 , n32574 , n28502 );
not ( n55524 , n32574 );
and ( n55525 , n55524 , n28508 );
nor ( n55526 , n55523 , n55525 );
and ( n233288 , n29117 , n55526 );
not ( n233289 , n29117 );
not ( n55529 , n55526 );
and ( n55530 , n233289 , n55529 );
nor ( n55531 , n233288 , n55530 );
not ( n55532 , n55531 );
not ( n55533 , n55532 );
not ( n55534 , n55533 );
not ( n233296 , n29250 );
not ( n233297 , n30163 );
or ( n55537 , n233296 , n233297 );
or ( n55538 , n30163 , n29250 );
nand ( n233300 , n55537 , n55538 );
and ( n233301 , n233300 , n30207 );
not ( n55541 , n233300 );
and ( n55542 , n55541 , n30200 );
nor ( n55543 , n233301 , n55542 );
buf ( n55544 , RI173e6e48_1630);
not ( n233306 , n55544 );
not ( n233307 , n31176 );
or ( n55547 , n233306 , n233307 );
not ( n55548 , n55544 );
nand ( n55549 , n55548 , n36684 );
nand ( n55550 , n55547 , n55549 );
and ( n233312 , n55550 , n36238 );
not ( n233313 , n55550 );
and ( n55553 , n233313 , n36243 );
nor ( n233315 , n233312 , n55553 );
nand ( n233316 , n55543 , n233315 );
not ( n55556 , n233316 );
or ( n233318 , n55534 , n55556 );
not ( n233319 , n233315 );
not ( n55559 , n233319 );
nand ( n55560 , n55559 , n55543 );
or ( n55561 , n55560 , n55533 );
nand ( n55562 , n233318 , n55561 );
not ( n233324 , n55562 );
not ( n233325 , n37549 );
not ( n55565 , n27960 );
or ( n55566 , n233325 , n55565 );
or ( n55567 , n27960 , n37549 );
nand ( n55568 , n55566 , n55567 );
not ( n233330 , n55568 );
not ( n233331 , n233330 );
not ( n55571 , n27926 );
or ( n55572 , n233331 , n55571 );
nand ( n55573 , n205688 , n55568 );
nand ( n55574 , n55572 , n55573 );
not ( n233336 , n55574 );
not ( n233337 , n220964 );
not ( n55577 , n40552 );
not ( n55578 , n55577 );
not ( n55579 , n34225 );
or ( n55580 , n55578 , n55579 );
nand ( n233342 , n34218 , n40552 );
nand ( n233343 , n55580 , n233342 );
not ( n55583 , n233343 );
and ( n233345 , n233337 , n55583 );
and ( n233346 , n220964 , n233343 );
nor ( n55586 , n233345 , n233346 );
not ( n233348 , n55586 );
nand ( n233349 , n233336 , n233348 );
not ( n55589 , n41593 );
not ( n55590 , n34840 );
not ( n55591 , n34263 );
not ( n55592 , n55591 );
or ( n233354 , n55590 , n55592 );
or ( n233355 , n55591 , n34840 );
nand ( n55595 , n233354 , n233355 );
not ( n55596 , n55595 );
or ( n55597 , n55589 , n55596 );
or ( n55598 , n55595 , n45702 );
nand ( n233360 , n55597 , n55598 );
buf ( n233361 , n233360 );
xor ( n55601 , n233349 , n233361 );
not ( n55602 , n55601 );
or ( n55603 , n233324 , n55602 );
or ( n55604 , n55562 , n55601 );
nand ( n233366 , n55603 , n55604 );
not ( n233367 , n33795 );
not ( n55607 , n38801 );
or ( n233369 , n233367 , n55607 );
not ( n233370 , n33795 );
nand ( n55610 , n233370 , n38806 );
nand ( n55611 , n233369 , n55610 );
and ( n55612 , n55611 , n219311 );
not ( n55613 , n55611 );
and ( n233375 , n55613 , n53990 );
nor ( n233376 , n55612 , n233375 );
not ( n55616 , n25472 );
not ( n233378 , n37946 );
or ( n233379 , n55616 , n233378 );
or ( n55619 , n40418 , n25472 );
nand ( n55620 , n233379 , n55619 );
not ( n55621 , n55620 );
not ( n55622 , n40426 );
and ( n55623 , n55621 , n55622 );
and ( n233385 , n55620 , n40426 );
nor ( n233386 , n55623 , n233385 );
nand ( n55626 , n233376 , n233386 );
not ( n55627 , n55626 );
not ( n55628 , n28969 );
not ( n55629 , n30409 );
and ( n55630 , n55628 , n55629 );
and ( n233392 , n206777 , n30409 );
nor ( n233393 , n55630 , n233392 );
buf ( n55633 , n33002 );
xnor ( n55634 , n233393 , n55633 );
not ( n55635 , n55634 );
or ( n55636 , n55627 , n55635 );
or ( n233398 , n55634 , n55626 );
nand ( n233399 , n55636 , n233398 );
and ( n55639 , n233366 , n233399 );
not ( n55640 , n233366 );
not ( n55641 , n233399 );
and ( n55642 , n55640 , n55641 );
nor ( n233404 , n55639 , n55642 );
not ( n233405 , n34038 );
not ( n55645 , n220845 );
or ( n55646 , n233405 , n55645 );
or ( n55647 , n220845 , n34038 );
nand ( n55648 , n55646 , n55647 );
and ( n233410 , n55648 , n41258 );
not ( n233411 , n55648 );
and ( n55651 , n233411 , n41257 );
nor ( n55652 , n233410 , n55651 );
buf ( n55653 , RI174a1a18_948);
not ( n55654 , n55653 );
not ( n233416 , n204255 );
or ( n233417 , n55654 , n233416 );
or ( n55657 , n204255 , n55653 );
nand ( n55658 , n233417 , n55657 );
and ( n55659 , n29815 , n55658 );
not ( n55660 , n55659 );
or ( n233422 , n55658 , n29815 );
nand ( n233423 , n55660 , n233422 );
and ( n55663 , n233423 , n29855 );
not ( n55664 , n233423 );
and ( n55665 , n55664 , n29860 );
nor ( n55666 , n55663 , n55665 );
nand ( n233428 , n55652 , n55666 );
not ( n233429 , n233428 );
not ( n55669 , n33153 );
not ( n233431 , n28247 );
or ( n233432 , n55669 , n233431 );
nand ( n55672 , n49504 , n33149 );
nand ( n233434 , n233432 , n55672 );
and ( n233435 , n233434 , n223793 );
not ( n55675 , n233434 );
and ( n233437 , n55675 , n34115 );
nor ( n55677 , n233435 , n233437 );
not ( n233439 , n55677 );
and ( n233440 , n233429 , n233439 );
and ( n55680 , n233428 , n55677 );
nor ( n55681 , n233440 , n55680 );
not ( n55682 , n55681 );
not ( n55683 , n30125 );
not ( n233445 , n40345 );
or ( n233446 , n55683 , n233445 );
not ( n55686 , n205846 );
or ( n55687 , n55686 , n30125 );
nand ( n55688 , n233446 , n55687 );
and ( n55689 , n55688 , n28122 );
not ( n233451 , n55688 );
and ( n233452 , n233451 , n28125 );
nor ( n55692 , n55689 , n233452 );
and ( n55693 , n30198 , n52704 );
not ( n55694 , n30198 );
and ( n55695 , n55694 , n27721 );
nor ( n233457 , n55693 , n55695 );
not ( n233458 , n233457 );
not ( n55698 , n27762 );
and ( n55699 , n233458 , n55698 );
and ( n55700 , n233457 , n27759 );
nor ( n55701 , n55699 , n55700 );
not ( n233463 , n55701 );
nand ( n233464 , n55692 , n233463 );
not ( n55704 , n220531 );
not ( n233466 , n41395 );
or ( n233467 , n55704 , n233466 );
nand ( n55707 , n41398 , n42766 );
nand ( n233469 , n233467 , n55707 );
buf ( n233470 , n204936 );
xnor ( n55710 , n233469 , n233470 );
not ( n55711 , n55710 );
and ( n55712 , n233464 , n55711 );
not ( n55713 , n233464 );
and ( n55714 , n55713 , n55710 );
nor ( n233476 , n55712 , n55714 );
not ( n233477 , n233476 );
or ( n55717 , n55682 , n233477 );
or ( n55718 , n233476 , n55681 );
nand ( n55719 , n55717 , n55718 );
and ( n55720 , n233404 , n55719 );
not ( n55721 , n233404 );
not ( n233483 , n55719 );
and ( n233484 , n55721 , n233483 );
nor ( n55724 , n55720 , n233484 );
not ( n55725 , n55724 );
not ( n55726 , n55725 );
not ( n55727 , n55726 );
and ( n233489 , n233283 , n55727 );
not ( n233490 , n233283 );
not ( n55730 , n55725 );
and ( n55731 , n233490 , n55730 );
nor ( n55732 , n233489 , n55731 );
nor ( n55733 , n55732 , n31572 );
nand ( n233495 , n233277 , n55733 );
nor ( n233496 , n55513 , n54208 );
not ( n55736 , n55732 );
not ( n55737 , n55332 );
nor ( n55738 , n55736 , n55737 );
nand ( n55739 , n233496 , n55738 );
buf ( n233501 , n35431 );
nand ( n233502 , n233501 , n38160 );
nand ( n55742 , n233495 , n55739 , n233502 );
buf ( n55743 , n55742 );
buf ( n55744 , n40793 );
buf ( n55745 , n35759 );
buf ( n233507 , n25328 );
not ( n233508 , RI19aaa858_2492);
or ( n55748 , n233507 , n233508 );
not ( n55749 , RI19a82538_2778);
or ( n55750 , n25336 , n55749 );
nand ( n55751 , n55748 , n55750 );
buf ( n233513 , n55751 );
not ( n233514 , RI19a88e38_2732);
or ( n233515 , n233507 , n233514 );
not ( n233516 , RI19accea8_2232);
or ( n55756 , n25335 , n233516 );
nand ( n233518 , n233515 , n55756 );
buf ( n233519 , n233518 );
not ( n55759 , n39914 );
buf ( n55760 , n31577 );
not ( n55761 , n55760 );
or ( n55762 , n55759 , n55761 );
nand ( n55763 , n42193 , n42170 );
and ( n55764 , n55763 , n221320 );
not ( n55765 , n55763 );
not ( n55766 , n221320 );
and ( n55767 , n55765 , n55766 );
nor ( n55768 , n55764 , n55767 );
not ( n55769 , n55768 );
not ( n55770 , n55769 );
not ( n233532 , n43722 );
or ( n233533 , n55770 , n233532 );
not ( n55773 , n55769 );
not ( n55774 , n43722 );
nand ( n55775 , n55773 , n55774 );
nand ( n55776 , n233533 , n55775 );
and ( n233538 , n55776 , n43956 );
not ( n233539 , n55776 );
and ( n55779 , n233539 , n43964 );
nor ( n55780 , n233538 , n55779 );
not ( n55781 , n55780 );
not ( n55782 , n33513 );
not ( n55783 , n55782 );
not ( n55784 , n55783 );
not ( n55785 , n38250 );
or ( n55786 , n55784 , n55785 );
or ( n55787 , n38250 , n55783 );
nand ( n233549 , n55786 , n55787 );
and ( n233550 , n233549 , n35358 );
not ( n233551 , n233549 );
and ( n233552 , n233551 , n38257 );
nor ( n55792 , n233550 , n233552 );
nand ( n55793 , n45473 , n55792 );
and ( n55794 , n55793 , n226869 );
not ( n55795 , n55793 );
and ( n233557 , n55795 , n49109 );
nor ( n233558 , n55794 , n233557 );
not ( n55798 , n233558 );
not ( n55799 , n33979 );
not ( n55800 , n39207 );
or ( n55801 , n55799 , n55800 );
or ( n233563 , n39207 , n33979 );
nand ( n233564 , n55801 , n233563 );
xnor ( n55804 , n233564 , n39251 );
not ( n55805 , n55804 );
nand ( n55806 , n55805 , n226849 );
not ( n55807 , n55806 );
not ( n233569 , n45422 );
and ( n233570 , n55807 , n233569 );
and ( n55810 , n55806 , n45422 );
nor ( n233572 , n233570 , n55810 );
not ( n233573 , n233572 );
not ( n55813 , n55792 );
nand ( n55814 , n226869 , n55813 );
and ( n55815 , n55814 , n226871 );
not ( n55816 , n55814 );
and ( n233578 , n55816 , n45456 );
nor ( n233579 , n55815 , n233578 );
not ( n55819 , n233579 );
or ( n55820 , n233573 , n55819 );
or ( n55821 , n233579 , n233572 );
nand ( n55822 , n55820 , n55821 );
not ( n233584 , n29773 );
not ( n233585 , n25592 );
buf ( n55825 , n34289 );
not ( n55826 , n55825 );
and ( n55827 , n233585 , n55826 );
and ( n55828 , n35635 , n55825 );
nor ( n233590 , n55827 , n55828 );
not ( n233591 , n233590 );
and ( n55831 , n233584 , n233591 );
and ( n55832 , n207535 , n233590 );
nor ( n55833 , n55831 , n55832 );
not ( n55834 , n55833 );
not ( n55835 , n223077 );
nand ( n55836 , n55834 , n55835 );
and ( n55837 , n55836 , n45275 );
not ( n233599 , n55836 );
and ( n233600 , n233599 , n223035 );
nor ( n233601 , n55837 , n233600 );
and ( n233602 , n55822 , n233601 );
not ( n55842 , n55822 );
not ( n55843 , n233601 );
and ( n55844 , n55842 , n55843 );
nor ( n55845 , n233602 , n55844 );
not ( n233607 , n55845 );
buf ( n233608 , n210649 );
not ( n55848 , n233608 );
not ( n55849 , n204744 );
or ( n55850 , n55848 , n55849 );
or ( n55851 , n204744 , n233608 );
nand ( n233613 , n55850 , n55851 );
and ( n233614 , n233613 , n214472 );
not ( n55854 , n233613 );
and ( n55855 , n55854 , n47231 );
nor ( n55856 , n233614 , n55855 );
not ( n55857 , n55856 );
not ( n233619 , n226928 );
nand ( n233620 , n55857 , n233619 );
and ( n55860 , n233620 , n49151 );
not ( n55861 , n233620 );
and ( n55862 , n55861 , n45340 );
nor ( n55863 , n55860 , n55862 );
not ( n233625 , n55863 );
buf ( n233626 , n40798 );
not ( n55866 , n233626 );
not ( n55867 , n32347 );
or ( n55868 , n55866 , n55867 );
or ( n55869 , n230248 , n233626 );
nand ( n233631 , n55868 , n55869 );
buf ( n233632 , n31528 );
and ( n55872 , n233631 , n233632 );
not ( n233634 , n233631 );
and ( n233635 , n233634 , n31515 );
nor ( n233636 , n55872 , n233635 );
nand ( n233637 , n226900 , n233636 );
not ( n55877 , n233637 );
not ( n55878 , n223136 );
and ( n233640 , n55877 , n55878 );
and ( n233641 , n233637 , n223136 );
nor ( n55881 , n233640 , n233641 );
not ( n55882 , n55881 );
and ( n55883 , n233625 , n55882 );
and ( n55884 , n55863 , n55881 );
nor ( n233646 , n55883 , n55884 );
not ( n233647 , n233646 );
and ( n55887 , n233607 , n233647 );
and ( n55888 , n55845 , n233646 );
nor ( n55889 , n55887 , n55888 );
not ( n55890 , n55889 );
or ( n233652 , n55798 , n55890 );
not ( n233653 , n233558 );
not ( n55893 , n233646 );
not ( n55894 , n55845 );
or ( n55895 , n55893 , n55894 );
not ( n55896 , n55845 );
not ( n55897 , n233646 );
nand ( n55898 , n55896 , n55897 );
nand ( n233660 , n55895 , n55898 );
nand ( n233661 , n233653 , n233660 );
nand ( n233662 , n233652 , n233661 );
not ( n233663 , n32409 );
xor ( n55903 , n33505 , n33522 );
xnor ( n233665 , n55903 , n55782 );
not ( n233666 , n233665 );
not ( n55906 , n233666 );
or ( n233668 , n233663 , n55906 );
or ( n233669 , n225165 , n32409 );
nand ( n55909 , n233668 , n233669 );
and ( n55910 , n55909 , n48780 );
not ( n55911 , n55909 );
and ( n55912 , n55911 , n48781 );
nor ( n233674 , n55910 , n55912 );
not ( n233675 , n233674 );
not ( n55915 , n38657 );
not ( n55916 , n40828 );
not ( n55917 , n42956 );
or ( n55918 , n55916 , n55917 );
or ( n233680 , n42956 , n40828 );
nand ( n233681 , n55918 , n233680 );
not ( n55921 , n233681 );
or ( n233683 , n55915 , n55921 );
not ( n55923 , n233681 );
nand ( n233685 , n55923 , n220726 );
nand ( n233686 , n233683 , n233685 );
nand ( n55926 , n233675 , n233686 );
not ( n55927 , n55926 );
not ( n55928 , n45579 );
and ( n55929 , n55927 , n55928 );
and ( n233691 , n55926 , n45579 );
nor ( n233692 , n55929 , n233691 );
not ( n55932 , n233692 );
not ( n55933 , n34060 );
not ( n55934 , n48039 );
or ( n55935 , n55933 , n55934 );
or ( n233697 , n48039 , n34060 );
nand ( n233698 , n55935 , n233697 );
buf ( n55938 , n229405 );
and ( n55939 , n233698 , n55938 );
not ( n55940 , n233698 );
buf ( n55941 , n38558 );
and ( n233703 , n55940 , n55941 );
nor ( n233704 , n55939 , n233703 );
not ( n55944 , n26171 );
not ( n55945 , n36625 );
or ( n55946 , n55944 , n55945 );
or ( n55947 , n36625 , n26171 );
nand ( n233709 , n55946 , n55947 );
and ( n233710 , n233709 , n230227 );
not ( n55950 , n233709 );
and ( n55951 , n55950 , n225682 );
nor ( n55952 , n233710 , n55951 );
not ( n55953 , n55952 );
nand ( n233715 , n233704 , n55953 );
buf ( n233716 , n45519 );
and ( n55956 , n233715 , n233716 );
not ( n55957 , n233715 );
not ( n55958 , n233716 );
and ( n55959 , n55957 , n55958 );
nor ( n233721 , n55956 , n55959 );
not ( n233722 , n233721 );
or ( n55962 , n55932 , n233722 );
or ( n55963 , n233721 , n233692 );
nand ( n55964 , n55962 , n55963 );
not ( n55965 , n32180 );
not ( n233727 , n55965 );
not ( n233728 , n38444 );
and ( n55968 , n233727 , n233728 );
and ( n233730 , n32175 , n38444 );
nor ( n233731 , n55968 , n233730 );
and ( n55971 , n233731 , n42091 );
not ( n55972 , n233731 );
and ( n55973 , n55972 , n42096 );
nor ( n55974 , n55971 , n55973 );
buf ( n233736 , n55974 );
not ( n233737 , n233736 );
xor ( n55977 , n32289 , n39361 );
xnor ( n55978 , n55977 , n41971 );
nand ( n55979 , n233737 , n55978 );
and ( n55980 , n55979 , n45625 );
not ( n233742 , n55979 );
and ( n233743 , n233742 , n45626 );
nor ( n55983 , n55980 , n233743 );
and ( n233745 , n55964 , n55983 );
not ( n55985 , n55964 );
not ( n55986 , n55983 );
and ( n55987 , n55985 , n55986 );
nor ( n55988 , n233745 , n55987 );
not ( n233750 , n55988 );
not ( n233751 , n45656 );
xor ( n55991 , n204457 , n47216 );
xnor ( n55992 , n55991 , n27968 );
not ( n55993 , n204764 );
not ( n55994 , n33182 );
or ( n233756 , n55993 , n55994 );
or ( n233757 , n210940 , n204764 );
nand ( n55997 , n233756 , n233757 );
and ( n55998 , n55997 , n31037 );
not ( n55999 , n55997 );
and ( n56000 , n55999 , n33186 );
or ( n233762 , n55998 , n56000 );
not ( n233763 , n233762 );
nand ( n56003 , n55992 , n233763 );
not ( n56004 , n56003 );
or ( n56005 , n233751 , n56004 );
or ( n56006 , n56003 , n45656 );
nand ( n233768 , n56005 , n56006 );
not ( n233769 , n233768 );
not ( n56009 , n31981 );
not ( n56010 , n31227 );
or ( n56011 , n56009 , n56010 );
or ( n56012 , n31227 , n31981 );
nand ( n56013 , n56011 , n56012 );
not ( n56014 , n56013 );
not ( n233776 , n29258 );
and ( n233777 , n56014 , n233776 );
and ( n56017 , n56013 , n29258 );
nor ( n56018 , n233777 , n56017 );
xor ( n56019 , n32734 , n35754 );
xnor ( n56020 , n56019 , n44003 );
nand ( n56021 , n56018 , n56020 );
not ( n233783 , n56021 );
not ( n233784 , n45697 );
and ( n56024 , n233783 , n233784 );
not ( n233786 , n56018 );
not ( n233787 , n233786 );
nand ( n56027 , n233787 , n56020 );
and ( n56028 , n56027 , n45697 );
nor ( n56029 , n56024 , n56028 );
not ( n56030 , n56029 );
or ( n233792 , n233769 , n56030 );
or ( n233793 , n56029 , n233768 );
nand ( n56033 , n233792 , n233793 );
not ( n56034 , n56033 );
not ( n56035 , n56034 );
or ( n56036 , n233750 , n56035 );
not ( n233798 , n55988 );
nand ( n233799 , n56033 , n233798 );
nand ( n56039 , n56036 , n233799 );
not ( n56040 , n56039 );
not ( n56041 , n56040 );
and ( n56042 , n233662 , n56041 );
not ( n233804 , n233662 );
buf ( n233805 , n56040 );
and ( n56045 , n233804 , n233805 );
nor ( n56046 , n56042 , n56045 );
nand ( n56047 , n55781 , n56046 );
not ( n56048 , n221191 );
not ( n233810 , n56048 );
buf ( n233811 , n41441 );
not ( n56051 , n233811 );
not ( n233813 , n224685 );
or ( n233814 , n56051 , n233813 );
or ( n56054 , n25765 , n233811 );
nand ( n233816 , n233814 , n56054 );
and ( n233817 , n233816 , n25772 );
not ( n56057 , n233816 );
and ( n56058 , n56057 , n25773 );
nor ( n56059 , n233817 , n56058 );
nand ( n56060 , n56059 , n43419 );
not ( n233822 , n56060 );
or ( n233823 , n233810 , n233822 );
or ( n56063 , n56060 , n56048 );
nand ( n56064 , n233823 , n56063 );
not ( n56065 , n56064 );
not ( n56066 , n43497 );
or ( n233828 , n56065 , n56066 );
not ( n233829 , n56064 );
nand ( n56069 , n233829 , n43504 );
nand ( n56070 , n233828 , n56069 );
not ( n56071 , n56070 );
not ( n56072 , n43220 );
and ( n233834 , n56071 , n56072 );
and ( n233835 , n56070 , n43220 );
nor ( n56075 , n233834 , n233835 );
not ( n233837 , n56075 );
and ( n233838 , n56047 , n233837 );
not ( n56078 , n56047 );
and ( n233840 , n56078 , n56075 );
nor ( n233841 , n233838 , n233840 );
or ( n233842 , n233841 , n39763 );
nand ( n233843 , n55762 , n233842 );
buf ( n233844 , n233843 );
buf ( n233845 , n28458 );
not ( n233846 , n33485 );
not ( n233847 , n233846 );
not ( n233848 , n33372 );
nand ( n233849 , n27970 , n233848 );
and ( n233850 , n233849 , n28052 );
not ( n233851 , n233849 );
and ( n233852 , n233851 , n28051 );
nor ( n233853 , n233850 , n233852 );
not ( n233854 , n233853 );
not ( n233855 , n233854 );
not ( n233856 , n33317 );
nand ( n233857 , n33305 , n233856 );
not ( n233858 , n233857 );
buf ( n233859 , n28208 );
not ( n233860 , n233859 );
and ( n233861 , n233858 , n233860 );
and ( n233862 , n233857 , n233859 );
nor ( n233863 , n233861 , n233862 );
not ( n233864 , n233863 );
not ( n233865 , n233864 );
or ( n233866 , n233855 , n233865 );
nand ( n233867 , n233863 , n233853 );
nand ( n233868 , n233866 , n233867 );
nand ( n233869 , n33405 , n33480 );
not ( n233870 , n233869 );
not ( n233871 , n28425 );
and ( n233872 , n233870 , n233871 );
and ( n233873 , n233869 , n28425 );
nor ( n233874 , n233872 , n233873 );
not ( n233875 , n233874 );
and ( n233876 , n233868 , n233875 );
not ( n233877 , n233868 );
and ( n233878 , n233877 , n233874 );
nor ( n233879 , n233876 , n233878 );
nand ( n233880 , n33669 , n33690 );
not ( n233881 , n233880 );
not ( n233882 , n28726 );
not ( n233883 , n233882 );
and ( n233884 , n233881 , n233883 );
and ( n233885 , n233880 , n233882 );
nor ( n233886 , n233884 , n233885 );
not ( n233887 , n233886 );
not ( n233888 , n28881 );
nand ( n233889 , n33621 , n33571 );
not ( n233890 , n233889 );
or ( n233891 , n233888 , n233890 );
nand ( n233892 , n33621 , n33571 );
or ( n233893 , n233892 , n28881 );
nand ( n233894 , n233891 , n233893 );
not ( n233895 , n233894 );
or ( n233896 , n233887 , n233895 );
or ( n233897 , n233894 , n233886 );
nand ( n233898 , n233896 , n233897 );
buf ( n233899 , n233898 );
xnor ( n233900 , n233879 , n233899 );
not ( n233901 , n233900 );
or ( n233902 , n233847 , n233901 );
not ( n233903 , n233846 );
not ( n233904 , n233900 );
nand ( n233905 , n233903 , n233904 );
nand ( n233906 , n233902 , n233905 );
not ( n233907 , n233150 );
nand ( n233908 , n55400 , n233907 );
buf ( n233909 , n29652 );
xor ( n233910 , n233908 , n233909 );
not ( n233911 , n233910 );
nand ( n233912 , n233121 , n233133 );
not ( n233913 , n233912 );
not ( n233914 , n29863 );
and ( n233915 , n233913 , n233914 );
and ( n233916 , n233912 , n29863 );
nor ( n233917 , n233915 , n233916 );
not ( n233918 , n233917 );
or ( n233919 , n233911 , n233918 );
not ( n233920 , n233910 );
not ( n233921 , n233917 );
nand ( n233922 , n233920 , n233921 );
nand ( n233923 , n233919 , n233922 );
not ( n233924 , n233923 );
nand ( n233925 , n55412 , n233186 );
not ( n233926 , n233925 );
not ( n233927 , n29260 );
and ( n233928 , n233926 , n233927 );
not ( n233929 , n55426 );
nand ( n233930 , n233929 , n55412 );
and ( n233931 , n233930 , n29260 );
nor ( n233932 , n233928 , n233931 );
not ( n233933 , n233932 );
not ( n233934 , n55461 );
nand ( n233935 , n233934 , n55448 );
buf ( n233936 , n206779 );
and ( n233937 , n233935 , n233936 );
not ( n233938 , n233935 );
not ( n233939 , n233936 );
and ( n233940 , n233938 , n233939 );
nor ( n233941 , n233937 , n233940 );
not ( n233942 , n233941 );
or ( n233943 , n233933 , n233942 );
or ( n233944 , n233941 , n233932 );
nand ( n233945 , n233943 , n233944 );
nand ( n233946 , n233234 , n55488 );
and ( n233947 , n233946 , n29373 );
not ( n233948 , n233946 );
and ( n233949 , n233948 , n29374 );
nor ( n233950 , n233947 , n233949 );
not ( n233951 , n233950 );
and ( n233952 , n233945 , n233951 );
not ( n233953 , n233945 );
and ( n233954 , n233953 , n233950 );
nor ( n233955 , n233952 , n233954 );
not ( n233956 , n233955 );
or ( n233957 , n233924 , n233956 );
or ( n233958 , n233955 , n233923 );
nand ( n233959 , n233957 , n233958 );
buf ( n233960 , n233959 );
and ( n233961 , n233906 , n233960 );
not ( n233962 , n233906 );
and ( n233963 , n233955 , n233923 );
not ( n233964 , n233955 );
not ( n233965 , n233923 );
and ( n233966 , n233964 , n233965 );
nor ( n233967 , n233963 , n233966 );
buf ( n233968 , n233967 );
and ( n233969 , n233962 , n233968 );
nor ( n233970 , n233961 , n233969 );
buf ( n233971 , n27886 );
buf ( n233972 , n233971 );
not ( n233973 , n233972 );
nand ( n233974 , n233970 , n233973 );
nand ( n233975 , n40923 , n42629 );
not ( n233976 , n233975 );
not ( n233977 , n40937 );
and ( n233978 , n233976 , n233977 );
and ( n233979 , n233975 , n40937 );
nor ( n233980 , n233978 , n233979 );
not ( n233981 , n233980 );
not ( n233982 , n233981 );
not ( n233983 , n41216 );
or ( n233984 , n233982 , n233983 );
not ( n233985 , n233981 );
xor ( n233986 , n41089 , n41039 );
xnor ( n233987 , n233986 , n41211 );
nand ( n233988 , n233985 , n233987 );
nand ( n233989 , n233984 , n233988 );
buf ( n233990 , n44176 );
and ( n233991 , n233989 , n233990 );
not ( n233992 , n233989 );
and ( n233993 , n44173 , n44174 );
not ( n233994 , n44173 );
not ( n233995 , n44174 );
and ( n233996 , n233994 , n233995 );
nor ( n233997 , n233993 , n233996 );
and ( n233998 , n233992 , n233997 );
nor ( n233999 , n233991 , n233998 );
not ( n234000 , n34826 );
nor ( n234001 , n39579 , n231815 );
not ( n234002 , n234001 );
and ( n234003 , n234000 , n234002 );
and ( n234004 , n34826 , n234001 );
nor ( n234005 , n234003 , n234004 );
not ( n234006 , n234005 );
not ( n234007 , n234006 );
not ( n234008 , n39595 );
or ( n234009 , n234007 , n234008 );
not ( n234010 , n234006 );
nand ( n234011 , n234010 , n39598 );
nand ( n234012 , n234009 , n234011 );
not ( n234013 , n39749 );
and ( n234014 , n234012 , n234013 );
not ( n234015 , n234012 );
and ( n234016 , n234015 , n39755 );
nor ( n234017 , n234014 , n234016 );
nor ( n234018 , n233999 , n234017 );
or ( n234019 , n233974 , n234018 );
nor ( n234020 , n233970 , n233999 );
buf ( n234021 , n35427 );
nor ( n234022 , n234017 , n234021 );
nand ( n234023 , n234020 , n234022 );
buf ( n234024 , n31575 );
nand ( n234025 , n234024 , n205089 );
nand ( n234026 , n234019 , n234023 , n234025 );
buf ( n234027 , n234026 );
not ( n234028 , RI19a936f8_2658);
or ( n234029 , n25328 , n234028 );
not ( n234030 , RI19a894c8_2729);
or ( n234031 , n25335 , n234030 );
nand ( n234032 , n234029 , n234031 );
buf ( n234033 , n234032 );
buf ( n234034 , n31248 );
buf ( n234035 , n35094 );
buf ( n234036 , RI1747e5b8_1120);
buf ( n234037 , n234036 );
buf ( n234038 , n28231 );
buf ( n234039 , n34542 );
not ( n234040 , RI19a95b88_2642);
or ( n234041 , n25328 , n234040 );
not ( n234042 , RI19a8bbb0_2713);
or ( n234043 , n226822 , n234042 );
nand ( n234044 , n234041 , n234043 );
buf ( n234045 , n234044 );
not ( n234046 , n221776 );
not ( n234047 , n54325 );
or ( n234048 , n234046 , n234047 );
or ( n234049 , n54325 , n221776 );
nand ( n234050 , n234048 , n234049 );
not ( n234051 , n37787 );
nand ( n234052 , n222058 , n38209 );
not ( n234053 , n234052 );
not ( n234054 , n38143 );
and ( n234055 , n234053 , n234054 );
and ( n234056 , n234052 , n38143 );
nor ( n234057 , n234055 , n234056 );
not ( n234058 , n234057 );
or ( n234059 , n234051 , n234058 );
or ( n234060 , n234057 , n37787 );
nand ( n234061 , n234059 , n234060 );
not ( n234062 , n234061 );
not ( n234063 , n38038 );
nand ( n234064 , n234063 , n222027 );
not ( n234065 , n234064 );
not ( n234066 , n49979 );
and ( n234067 , n234065 , n234066 );
and ( n234068 , n234064 , n49979 );
nor ( n234069 , n234067 , n234068 );
not ( n234070 , n234069 );
or ( n234071 , n234062 , n234070 );
or ( n234072 , n234069 , n234061 );
nand ( n234073 , n234071 , n234072 );
buf ( n234074 , n234073 );
not ( n234075 , n37810 );
nand ( n234076 , n234075 , n48829 );
not ( n234077 , n234076 );
not ( n234078 , n49991 );
and ( n234079 , n234077 , n234078 );
and ( n234080 , n234076 , n49991 );
nor ( n234081 , n234079 , n234080 );
not ( n234082 , n234081 );
not ( n234083 , n234082 );
not ( n234084 , n37906 );
nand ( n234085 , n48818 , n234084 );
buf ( n234086 , n50000 );
xnor ( n234087 , n234085 , n234086 );
not ( n234088 , n234087 );
not ( n234089 , n234088 );
or ( n234090 , n234083 , n234089 );
nand ( n234091 , n234087 , n234081 );
nand ( n234092 , n234090 , n234091 );
not ( n234093 , n234092 );
and ( n234094 , n234074 , n234093 );
not ( n234095 , n234074 );
and ( n234096 , n234095 , n234092 );
nor ( n234097 , n234094 , n234096 );
buf ( n234098 , n234097 );
and ( n234099 , n234050 , n234098 );
not ( n234100 , n234050 );
not ( n234101 , n234093 );
not ( n234102 , n234073 );
or ( n234103 , n234101 , n234102 );
not ( n234104 , n234073 );
nand ( n234105 , n234104 , n234092 );
nand ( n234106 , n234103 , n234105 );
buf ( n234107 , n234106 );
and ( n234108 , n234100 , n234107 );
nor ( n234109 , n234099 , n234108 );
buf ( n234110 , n226003 );
not ( n234111 , n234110 );
nand ( n234112 , n234109 , n234111 );
not ( n234113 , n38588 );
not ( n234114 , n216359 );
nand ( n234115 , n234113 , n234114 );
and ( n234116 , n234115 , n226777 );
not ( n234117 , n234115 );
and ( n234118 , n234117 , n49015 );
nor ( n234119 , n234116 , n234118 );
not ( n234120 , n234119 );
not ( n234121 , n49042 );
and ( n234122 , n234120 , n234121 );
not ( n234123 , n234120 );
not ( n234124 , n49042 );
not ( n234125 , n234124 );
and ( n234126 , n234123 , n234125 );
or ( n234127 , n234122 , n234126 );
not ( n234128 , n234127 );
not ( n234129 , n45361 );
nand ( n234130 , n234129 , n49149 );
not ( n234131 , n234130 );
not ( n234132 , n55856 );
not ( n234133 , n234132 );
or ( n234134 , n234131 , n234133 );
or ( n234135 , n234132 , n234130 );
nand ( n234136 , n234134 , n234135 );
not ( n234137 , n234136 );
nand ( n234138 , n49143 , n45387 );
not ( n234139 , n234138 );
not ( n234140 , n233636 );
and ( n234141 , n234139 , n234140 );
and ( n234142 , n234138 , n233636 );
nor ( n234143 , n234141 , n234142 );
not ( n234144 , n234143 );
or ( n234145 , n234137 , n234144 );
not ( n234146 , n234136 );
not ( n234147 , n234143 );
nand ( n234148 , n234146 , n234147 );
nand ( n234149 , n234145 , n234148 );
not ( n234150 , n55813 );
nand ( n234151 , n45446 , n223231 );
not ( n234152 , n234151 );
or ( n234153 , n234150 , n234152 );
or ( n234154 , n234151 , n55813 );
nand ( n234155 , n234153 , n234154 );
not ( n234156 , n234155 );
nand ( n234157 , n223190 , n49093 );
not ( n234158 , n234157 );
not ( n234159 , n55804 );
not ( n234160 , n234159 );
and ( n234161 , n234158 , n234160 );
and ( n234162 , n234157 , n234159 );
nor ( n234163 , n234161 , n234162 );
not ( n234164 , n234163 );
or ( n234165 , n234156 , n234164 );
or ( n234166 , n234163 , n234155 );
nand ( n234167 , n234165 , n234166 );
not ( n234168 , n223252 );
nand ( n234169 , n234168 , n45324 );
not ( n234170 , n55834 );
and ( n234171 , n234169 , n234170 );
not ( n234172 , n234169 );
and ( n234173 , n234172 , n55834 );
nor ( n234174 , n234171 , n234173 );
and ( n234175 , n234167 , n234174 );
not ( n234176 , n234167 );
not ( n234177 , n234174 );
and ( n234178 , n234176 , n234177 );
nor ( n234179 , n234175 , n234178 );
and ( n234180 , n234149 , n234179 );
not ( n234181 , n234149 );
not ( n234182 , n234179 );
and ( n234183 , n234181 , n234182 );
nor ( n234184 , n234180 , n234183 );
buf ( n234185 , n234184 );
not ( n234186 , n234185 );
not ( n234187 , n234186 );
and ( n234188 , n234128 , n234187 );
and ( n234189 , n234127 , n234186 );
nor ( n234190 , n234188 , n234189 );
not ( n234191 , n234190 );
not ( n234192 , n42004 );
not ( n234193 , n234192 );
nand ( n234194 , n41989 , n219760 );
not ( n234195 , n234194 );
not ( n234196 , n55309 );
and ( n234197 , n234195 , n234196 );
nand ( n234198 , n41989 , n219760 );
and ( n234199 , n234198 , n55309 );
nor ( n234200 , n234197 , n234199 );
not ( n234201 , n234200 );
nand ( n234202 , n42031 , n53055 );
and ( n234203 , n234202 , n230778 );
not ( n234204 , n234202 );
and ( n234205 , n234204 , n230779 );
nor ( n234206 , n234203 , n234205 );
not ( n234207 , n234206 );
or ( n234208 , n234201 , n234207 );
or ( n234209 , n234206 , n234200 );
nand ( n234210 , n234208 , n234209 );
not ( n234211 , n41779 );
nand ( n234212 , n234211 , n53065 );
and ( n234213 , n234212 , n41790 );
not ( n234214 , n234212 );
and ( n234215 , n234214 , n41789 );
nor ( n234216 , n234213 , n234215 );
not ( n234217 , n234216 );
and ( n234218 , n234210 , n234217 );
not ( n234219 , n234210 );
and ( n234220 , n234219 , n234216 );
nor ( n234221 , n234218 , n234220 );
not ( n234222 , n234221 );
nand ( n234223 , n53028 , n42134 );
and ( n234224 , n234223 , n41881 );
not ( n234225 , n234223 );
and ( n234226 , n234225 , n41880 );
nor ( n234227 , n234224 , n234226 );
nand ( n234228 , n41896 , n230798 );
not ( n234229 , n234228 );
not ( n234230 , n41912 );
and ( n234231 , n234229 , n234230 );
and ( n234232 , n234228 , n41912 );
nor ( n234233 , n234231 , n234232 );
and ( n234234 , n234227 , n234233 );
not ( n234235 , n234227 );
not ( n234236 , n234233 );
and ( n234237 , n234235 , n234236 );
nor ( n234238 , n234234 , n234237 );
not ( n234239 , n234238 );
not ( n234240 , n234239 );
and ( n234241 , n234222 , n234240 );
and ( n234242 , n234221 , n234239 );
nor ( n234243 , n234241 , n234242 );
not ( n234244 , n234243 );
or ( n234245 , n234193 , n234244 );
not ( n234246 , n234192 );
not ( n234247 , n234239 );
not ( n234248 , n234221 );
or ( n234249 , n234247 , n234248 );
not ( n234250 , n234221 );
nand ( n234251 , n234250 , n234238 );
nand ( n234252 , n234249 , n234251 );
nand ( n234253 , n234246 , n234252 );
nand ( n234254 , n234245 , n234253 );
not ( n234255 , n43581 );
not ( n234256 , n42358 );
nand ( n234257 , n234256 , n42377 );
not ( n234258 , n234257 );
or ( n234259 , n234255 , n234258 );
not ( n234260 , n42358 );
nand ( n234261 , n234260 , n42377 );
or ( n234262 , n234261 , n43581 );
nand ( n234263 , n234259 , n234262 );
and ( n234264 , n234263 , n55768 );
not ( n234265 , n234263 );
and ( n234266 , n234265 , n55769 );
nor ( n234267 , n234264 , n234266 );
not ( n234268 , n234267 );
not ( n234269 , n43546 );
or ( n234270 , n234268 , n234269 );
or ( n234271 , n234267 , n43546 );
nand ( n234272 , n234270 , n234271 );
not ( n234273 , n43707 );
not ( n234274 , n234273 );
nand ( n234275 , n42251 , n42310 );
not ( n234276 , n234275 );
and ( n234277 , n234274 , n234276 );
and ( n234278 , n234273 , n234275 );
nor ( n234279 , n234277 , n234278 );
not ( n234280 , n234279 );
not ( n234281 , n234280 );
nand ( n234282 , n219993 , n53117 );
not ( n234283 , n234282 );
not ( n234284 , n43666 );
not ( n234285 , n234284 );
or ( n234286 , n234283 , n234285 );
or ( n234287 , n234284 , n234282 );
nand ( n234288 , n234286 , n234287 );
not ( n234289 , n234288 );
not ( n234290 , n234289 );
or ( n234291 , n234281 , n234290 );
nand ( n234292 , n234279 , n234288 );
nand ( n234293 , n234291 , n234292 );
and ( n234294 , n234272 , n234293 );
not ( n234295 , n234272 );
not ( n234296 , n234293 );
and ( n234297 , n234295 , n234296 );
nor ( n234298 , n234294 , n234297 );
buf ( n234299 , n234298 );
and ( n234300 , n234254 , n234299 );
not ( n234301 , n234254 );
and ( n234302 , n234272 , n234296 );
not ( n234303 , n234272 );
and ( n234304 , n234303 , n234293 );
nor ( n234305 , n234302 , n234304 );
buf ( n234306 , n234305 );
and ( n234307 , n234301 , n234306 );
nor ( n234308 , n234300 , n234307 );
not ( n234309 , n234308 );
nand ( n234310 , n234191 , n234309 );
or ( n234311 , n234112 , n234310 );
not ( n234312 , n234191 );
not ( n234313 , n234109 );
or ( n234314 , n234312 , n234313 );
nor ( n234315 , n234309 , n52445 );
nand ( n234316 , n234314 , n234315 );
nand ( n234317 , n31577 , n43240 );
nand ( n234318 , n234311 , n234316 , n234317 );
buf ( n234319 , n234318 );
not ( n234320 , n48397 );
not ( n234321 , n234320 );
not ( n234322 , n225243 );
nand ( n234323 , n234322 , n47332 );
not ( n234324 , n234323 );
or ( n234325 , n234321 , n234324 );
not ( n234326 , n225243 );
nand ( n234327 , n234326 , n47332 );
or ( n234328 , n234327 , n234320 );
nand ( n234329 , n234325 , n234328 );
not ( n234330 , n234329 );
not ( n234331 , n48413 );
or ( n234332 , n234330 , n234331 );
not ( n234333 , n234329 );
nand ( n234334 , n234333 , n48414 );
nand ( n234335 , n234332 , n234334 );
and ( n234336 , n234335 , n226320 );
not ( n234337 , n234335 );
and ( n234338 , n234337 , n226319 );
nor ( n234339 , n234336 , n234338 );
not ( n234340 , n234339 );
nand ( n234341 , n234340 , n233837 );
nand ( n234342 , n225742 , n48620 );
not ( n234343 , n234342 );
not ( n234344 , n47336 );
not ( n234345 , n208229 );
not ( n234346 , n41431 );
or ( n234347 , n234345 , n234346 );
not ( n234348 , n41431 );
nand ( n234349 , n234348 , n30464 );
nand ( n234350 , n234347 , n234349 );
xor ( n234351 , n32499 , n234350 );
xnor ( n234352 , n234351 , n41446 );
not ( n234353 , n234352 );
and ( n234354 , n234344 , n234353 );
and ( n234355 , n47336 , n234352 );
nor ( n234356 , n234354 , n234355 );
not ( n234357 , n234356 );
not ( n234358 , n234357 );
and ( n234359 , n234343 , n234358 );
and ( n234360 , n234342 , n234357 );
nor ( n234361 , n234359 , n234360 );
nand ( n234362 , n48598 , n47897 );
not ( n234363 , n55086 );
and ( n234364 , n234362 , n234363 );
not ( n234365 , n234362 );
not ( n234366 , n234363 );
and ( n234367 , n234365 , n234366 );
nor ( n234368 , n234364 , n234367 );
xor ( n234369 , n234361 , n234368 );
nand ( n234370 , n48581 , n47853 );
not ( n234371 , n234370 );
not ( n234372 , n39246 );
not ( n234373 , n33969 );
not ( n234374 , n39207 );
or ( n234375 , n234373 , n234374 );
or ( n234376 , n39207 , n33969 );
nand ( n234377 , n234375 , n234376 );
not ( n234378 , n234377 );
or ( n234379 , n234372 , n234378 );
or ( n234380 , n234377 , n39246 );
nand ( n234381 , n234379 , n234380 );
not ( n234382 , n234381 );
and ( n234383 , n234371 , n234382 );
and ( n234384 , n234370 , n234381 );
nor ( n234385 , n234383 , n234384 );
xor ( n234386 , n234369 , n234385 );
not ( n234387 , n37042 );
not ( n234388 , n45139 );
or ( n234389 , n234387 , n234388 );
nand ( n234390 , n43695 , n37038 );
nand ( n234391 , n234389 , n234390 );
not ( n234392 , n234391 );
not ( n234393 , n29372 );
and ( n234394 , n234392 , n234393 );
and ( n234395 , n234391 , n29372 );
nor ( n234396 , n234394 , n234395 );
not ( n234397 , n234396 );
not ( n234398 , n234397 );
nand ( n234399 , n47943 , n48645 );
not ( n234400 , n234399 );
or ( n234401 , n234398 , n234400 );
not ( n234402 , n226407 );
nand ( n234403 , n234402 , n47943 );
or ( n234404 , n234403 , n234397 );
nand ( n234405 , n234401 , n234404 );
not ( n234406 , n234405 );
nand ( n234407 , n225762 , n226424 );
and ( n234408 , n234407 , n47793 );
not ( n234409 , n234407 );
and ( n234410 , n234409 , n47792 );
nor ( n234411 , n234408 , n234410 );
not ( n234412 , n234411 );
and ( n234413 , n234406 , n234412 );
and ( n234414 , n234405 , n234411 );
nor ( n234415 , n234413 , n234414 );
and ( n234416 , n234386 , n234415 );
not ( n234417 , n234386 );
not ( n234418 , n234415 );
and ( n234419 , n234417 , n234418 );
nor ( n234420 , n234416 , n234419 );
not ( n234421 , n234420 );
nand ( n234422 , n225344 , n48465 );
and ( n234423 , n234422 , n47614 );
not ( n234424 , n234422 );
not ( n234425 , n47614 );
and ( n234426 , n234424 , n234425 );
nor ( n234427 , n234423 , n234426 );
buf ( n234428 , n234427 );
not ( n234429 , n234428 );
not ( n234430 , n225525 );
or ( n234431 , n234429 , n234430 );
not ( n234432 , n234428 );
nand ( n234433 , n234432 , n47773 );
nand ( n234434 , n234431 , n234433 );
not ( n234435 , n234434 );
or ( n234436 , n234421 , n234435 );
buf ( n234437 , n234420 );
or ( n234438 , n234434 , n234437 );
nand ( n234439 , n234436 , n234438 );
buf ( n234440 , n233971 );
nor ( n234441 , n234439 , n234440 );
not ( n234442 , n234441 );
or ( n234443 , n234341 , n234442 );
not ( n234444 , n234439 );
not ( n234445 , n205649 );
nor ( n234446 , n234444 , n234445 );
nand ( n234447 , n234341 , n234446 );
buf ( n234448 , n35431 );
nand ( n234449 , n234448 , n40115 );
nand ( n234450 , n234443 , n234447 , n234449 );
buf ( n234451 , n234450 );
not ( n234452 , n40002 );
buf ( n234453 , n234024 );
not ( n234454 , n234453 );
or ( n234455 , n234452 , n234454 );
not ( n234456 , n50027 );
not ( n234457 , n38009 );
and ( n234458 , n234456 , n234457 );
and ( n234459 , n50027 , n38009 );
nor ( n234460 , n234458 , n234459 );
not ( n234461 , n226719 );
not ( n234462 , n234461 );
nand ( n234463 , n38478 , n38399 );
not ( n234464 , n234463 );
or ( n234465 , n234462 , n234464 );
or ( n234466 , n234463 , n234461 );
nand ( n234467 , n234465 , n234466 );
not ( n234468 , n234467 );
nand ( n234469 , n38572 , n38510 );
not ( n234470 , n234469 );
not ( n234471 , n48993 );
and ( n234472 , n234470 , n234471 );
and ( n234473 , n234469 , n48993 );
nor ( n234474 , n234472 , n234473 );
not ( n234475 , n234474 );
or ( n234476 , n234468 , n234475 );
or ( n234477 , n234474 , n234467 );
nand ( n234478 , n234476 , n234477 );
and ( n234479 , n234478 , n234120 );
not ( n234480 , n234478 );
and ( n234481 , n234480 , n234119 );
nor ( n234482 , n234479 , n234481 );
not ( n234483 , n234482 );
buf ( n234484 , n226701 );
not ( n234485 , n234484 );
not ( n234486 , n38299 );
not ( n234487 , n38244 );
nand ( n234488 , n234486 , n234487 );
not ( n234489 , n234488 );
or ( n234490 , n234485 , n234489 );
or ( n234491 , n234488 , n234484 );
nand ( n234492 , n234490 , n234491 );
not ( n234493 , n234492 );
not ( n234494 , n38358 );
nand ( n234495 , n234494 , n38378 );
not ( n234496 , n234495 );
buf ( n234497 , n48896 );
not ( n234498 , n234497 );
or ( n234499 , n234496 , n234498 );
or ( n234500 , n234497 , n234495 );
nand ( n234501 , n234499 , n234500 );
not ( n234502 , n234501 );
not ( n234503 , n234502 );
or ( n234504 , n234493 , n234503 );
not ( n234505 , n234492 );
nand ( n234506 , n234505 , n234501 );
nand ( n234507 , n234504 , n234506 );
not ( n234508 , n234507 );
and ( n234509 , n234483 , n234508 );
not ( n234510 , n234483 );
not ( n234511 , n234508 );
and ( n234512 , n234510 , n234511 );
nor ( n234513 , n234509 , n234512 );
buf ( n234514 , n234513 );
and ( n234515 , n234460 , n234514 );
not ( n234516 , n234460 );
not ( n234517 , n234507 );
not ( n234518 , n234482 );
or ( n234519 , n234517 , n234518 );
nand ( n234520 , n234483 , n234508 );
nand ( n234521 , n234519 , n234520 );
buf ( n234522 , n234521 );
and ( n234523 , n234516 , n234522 );
nor ( n234524 , n234515 , n234523 );
not ( n234525 , n39011 );
nand ( n234526 , n39025 , n49757 );
not ( n234527 , n234526 );
or ( n234528 , n234525 , n234527 );
or ( n234529 , n234526 , n39011 );
nand ( n234530 , n234528 , n234529 );
not ( n234531 , n234530 );
not ( n234532 , n39052 );
or ( n234533 , n234531 , n234532 );
not ( n234534 , n234530 );
nand ( n234535 , n234534 , n39059 );
nand ( n234536 , n234533 , n234535 );
and ( n234537 , n234536 , n39435 );
not ( n234538 , n234536 );
and ( n234539 , n234538 , n39445 );
nor ( n234540 , n234537 , n234539 );
nand ( n234541 , n234524 , n234540 );
not ( n234542 , n234541 );
not ( n234543 , n53605 );
not ( n234544 , n53584 );
nand ( n234545 , n234543 , n234544 );
not ( n234546 , n234545 );
not ( n234547 , n30294 );
not ( n234548 , n222865 );
or ( n234549 , n234547 , n234548 );
or ( n234550 , n46753 , n30294 );
nand ( n234551 , n234549 , n234550 );
xor ( n234552 , n234551 , n45114 );
not ( n234553 , n234552 );
and ( n234554 , n234546 , n234553 );
and ( n234555 , n234545 , n234552 );
nor ( n234556 , n234554 , n234555 );
not ( n234557 , n234556 );
not ( n234558 , n234557 );
not ( n234559 , n38839 );
not ( n234560 , n25812 );
not ( n234561 , n234560 );
not ( n234562 , n47494 );
or ( n234563 , n234561 , n234562 );
or ( n234564 , n37106 , n234560 );
nand ( n234565 , n234563 , n234564 );
not ( n234566 , n234565 );
and ( n234567 , n234559 , n234566 );
and ( n234568 , n38839 , n234565 );
nor ( n234569 , n234567 , n234568 );
not ( n234570 , n234569 );
not ( n234571 , n234570 );
not ( n234572 , n31473 );
not ( n234573 , n40786 );
and ( n234574 , n234572 , n234573 );
and ( n234575 , n31473 , n40786 );
nor ( n234576 , n234574 , n234575 );
and ( n234577 , n234576 , n31515 );
not ( n234578 , n234576 );
and ( n234579 , n234578 , n31528 );
nor ( n234580 , n234577 , n234579 );
not ( n234581 , n234580 );
nand ( n234582 , n234581 , n53541 );
not ( n234583 , n234582 );
or ( n234584 , n234571 , n234583 );
or ( n234585 , n234582 , n234570 );
nand ( n234586 , n234584 , n234585 );
not ( n234587 , n234586 );
not ( n234588 , n233198 );
not ( n234589 , n25396 );
and ( n234590 , n234588 , n234589 );
and ( n234591 , n233198 , n25396 );
nor ( n234592 , n234590 , n234591 );
and ( n234593 , n234592 , n233207 );
not ( n234594 , n234592 );
and ( n234595 , n234594 , n41411 );
nor ( n234596 , n234593 , n234595 );
not ( n234597 , n234596 );
nand ( n234598 , n234597 , n231332 );
not ( n234599 , n234598 );
not ( n234600 , n28658 );
not ( n234601 , n30534 );
or ( n234602 , n234600 , n234601 );
or ( n234603 , n40230 , n28658 );
nand ( n234604 , n234602 , n234603 );
and ( n234605 , n234604 , n30497 );
not ( n234606 , n234604 );
and ( n234607 , n234606 , n208303 );
nor ( n234608 , n234605 , n234607 );
not ( n234609 , n234608 );
not ( n234610 , n234609 );
and ( n234611 , n234599 , n234610 );
and ( n234612 , n234598 , n234609 );
nor ( n234613 , n234611 , n234612 );
not ( n234614 , n234613 );
or ( n234615 , n234587 , n234614 );
or ( n234616 , n234613 , n234586 );
nand ( n234617 , n234615 , n234616 );
xor ( n234618 , n29673 , n34700 );
xnor ( n234619 , n234618 , n36859 );
not ( n234620 , n234619 );
nand ( n234621 , n234620 , n231254 );
not ( n234622 , n231230 );
and ( n234623 , n234621 , n234622 );
not ( n234624 , n234621 );
and ( n234625 , n234624 , n231230 );
nor ( n234626 , n234623 , n234625 );
and ( n234627 , n234617 , n234626 );
not ( n234628 , n234617 );
not ( n234629 , n234626 );
and ( n234630 , n234628 , n234629 );
nor ( n234631 , n234627 , n234630 );
not ( n234632 , n234631 );
not ( n234633 , n234632 );
not ( n234634 , n234552 );
nand ( n234635 , n234634 , n53605 );
not ( n234636 , n234635 );
xor ( n234637 , n30077 , n53417 );
xnor ( n234638 , n234637 , n33303 );
not ( n234639 , n234638 );
not ( n234640 , n234639 );
or ( n234641 , n234636 , n234640 );
or ( n234642 , n234639 , n234635 );
nand ( n234643 , n234641 , n234642 );
not ( n234644 , n234643 );
not ( n234645 , n31692 );
not ( n234646 , n26409 );
or ( n234647 , n234645 , n234646 );
not ( n234648 , n26409 );
nand ( n234649 , n234648 , n31688 );
nand ( n234650 , n234647 , n234649 );
and ( n234651 , n234650 , n53432 );
not ( n234652 , n234650 );
and ( n234653 , n234652 , n231190 );
nor ( n234654 , n234651 , n234653 );
and ( n234655 , n234654 , n53620 );
buf ( n234656 , n38119 );
not ( n234657 , n234656 );
not ( n234658 , n39417 );
not ( n234659 , n234658 );
or ( n234660 , n234657 , n234659 );
or ( n234661 , n234658 , n234656 );
nand ( n234662 , n234660 , n234661 );
and ( n234663 , n234662 , n47939 );
not ( n234664 , n234662 );
not ( n234665 , n47939 );
and ( n234666 , n234664 , n234665 );
nor ( n234667 , n234663 , n234666 );
not ( n234668 , n234667 );
not ( n234669 , n234668 );
and ( n234670 , n234655 , n234669 );
not ( n234671 , n234655 );
and ( n234672 , n234671 , n234668 );
nor ( n234673 , n234670 , n234672 );
not ( n234674 , n234673 );
and ( n234675 , n234644 , n234674 );
and ( n234676 , n234643 , n234673 );
nor ( n234677 , n234675 , n234676 );
not ( n234678 , n234677 );
not ( n234679 , n234678 );
and ( n234680 , n234633 , n234679 );
and ( n234681 , n234632 , n234678 );
nor ( n234682 , n234680 , n234681 );
not ( n234683 , n234682 );
or ( n234684 , n234558 , n234683 );
not ( n234685 , n234557 );
not ( n234686 , n234677 );
not ( n234687 , n234631 );
or ( n234688 , n234686 , n234687 );
not ( n234689 , n234631 );
nand ( n234690 , n234689 , n234678 );
nand ( n234691 , n234688 , n234690 );
nand ( n234692 , n234685 , n234691 );
nand ( n234693 , n234684 , n234692 );
not ( n234694 , n28088 );
not ( n234695 , n25426 );
or ( n234696 , n234694 , n234695 );
or ( n234697 , n25426 , n28088 );
nand ( n234698 , n234696 , n234697 );
and ( n234699 , n234698 , n28677 );
not ( n234700 , n234698 );
and ( n234701 , n234700 , n28680 );
nor ( n234702 , n234699 , n234701 );
not ( n234703 , n234702 );
nand ( n234704 , n234703 , n34120 );
not ( n234705 , n234704 );
xor ( n234706 , n33449 , n227444 );
xnor ( n234707 , n234706 , n32363 );
not ( n234708 , n234707 );
not ( n234709 , n234708 );
or ( n234710 , n234705 , n234709 );
or ( n234711 , n234708 , n234704 );
nand ( n234712 , n234710 , n234711 );
xor ( n234713 , n42261 , n45744 );
xnor ( n234714 , n234713 , n204825 );
nand ( n234715 , n234714 , n34393 );
not ( n234716 , n234715 );
not ( n234717 , n206789 );
not ( n234718 , n229482 );
not ( n234719 , n234718 );
or ( n234720 , n234717 , n234719 );
nand ( n234721 , n229482 , n29024 );
nand ( n234722 , n234720 , n234721 );
not ( n234723 , n234722 );
not ( n234724 , n36568 );
or ( n234725 , n234723 , n234724 );
or ( n234726 , n36568 , n234722 );
nand ( n234727 , n234725 , n234726 );
not ( n234728 , n234727 );
and ( n234729 , n234716 , n234728 );
and ( n234730 , n234715 , n234727 );
nor ( n234731 , n234729 , n234730 );
xor ( n234732 , n234712 , n234731 );
not ( n234733 , n234732 );
not ( n234734 , n37365 );
not ( n234735 , n222183 );
or ( n234736 , n234734 , n234735 );
not ( n234737 , n37365 );
nand ( n234738 , n234737 , n39359 );
nand ( n234739 , n234736 , n234738 );
not ( n234740 , n234739 );
not ( n234741 , n45468 );
and ( n234742 , n234740 , n234741 );
and ( n234743 , n234739 , n45465 );
nor ( n234744 , n234742 , n234743 );
not ( n234745 , n234744 );
not ( n234746 , n234745 );
not ( n234747 , n28405 );
nor ( n234748 , n26308 , n216952 );
not ( n234749 , n234748 );
nand ( n234750 , n26308 , n216952 );
nand ( n234751 , n234749 , n234750 );
not ( n234752 , n234751 );
and ( n234753 , n234747 , n234752 );
and ( n234754 , n227928 , n234751 );
nor ( n234755 , n234753 , n234754 );
nand ( n234756 , n234755 , n34310 );
not ( n234757 , n234756 );
or ( n234758 , n234746 , n234757 );
or ( n234759 , n234756 , n234745 );
nand ( n234760 , n234758 , n234759 );
not ( n234761 , n234760 );
xor ( n234762 , n36602 , n232877 );
xnor ( n234763 , n234762 , n38817 );
nand ( n234764 , n234763 , n33959 );
not ( n234765 , n204737 );
not ( n234766 , n26369 );
or ( n234767 , n234765 , n234766 );
nand ( n234768 , n26370 , n204733 );
nand ( n234769 , n234767 , n234768 );
not ( n234770 , n234769 );
not ( n234771 , n26409 );
and ( n234772 , n234770 , n234771 );
not ( n234773 , n43096 );
and ( n234774 , n234769 , n234773 );
nor ( n234775 , n234772 , n234774 );
not ( n234776 , n234775 );
and ( n234777 , n234764 , n234776 );
not ( n234778 , n234764 );
and ( n234779 , n234778 , n234775 );
nor ( n234780 , n234777 , n234779 );
not ( n234781 , n234780 );
or ( n234782 , n234761 , n234781 );
or ( n234783 , n234780 , n234760 );
nand ( n234784 , n234782 , n234783 );
xor ( n234785 , n37244 , n32406 );
xnor ( n234786 , n234785 , n33047 );
nand ( n234787 , n234786 , n34424 );
not ( n234788 , n33770 );
and ( n234789 , n234787 , n234788 );
not ( n234790 , n234787 );
and ( n234791 , n234790 , n33770 );
nor ( n234792 , n234789 , n234791 );
and ( n234793 , n234784 , n234792 );
not ( n234794 , n234784 );
not ( n234795 , n234792 );
and ( n234796 , n234794 , n234795 );
nor ( n234797 , n234793 , n234796 );
not ( n234798 , n234797 );
or ( n234799 , n234733 , n234798 );
not ( n234800 , n234797 );
not ( n234801 , n234732 );
nand ( n234802 , n234800 , n234801 );
nand ( n234803 , n234799 , n234802 );
buf ( n234804 , n234803 );
and ( n234805 , n234693 , n234804 );
not ( n234806 , n234693 );
and ( n234807 , n234797 , n234732 );
not ( n234808 , n234797 );
and ( n234809 , n234808 , n234801 );
nor ( n234810 , n234807 , n234809 );
buf ( n234811 , n234810 );
and ( n234812 , n234806 , n234811 );
nor ( n234813 , n234805 , n234812 );
not ( n234814 , n234813 );
and ( n234815 , n234542 , n234814 );
and ( n234816 , n234541 , n234813 );
nor ( n234817 , n234815 , n234816 );
buf ( n234818 , n226003 );
or ( n234819 , n234817 , n234818 );
nand ( n234820 , n234455 , n234819 );
buf ( n234821 , n234820 );
not ( n234822 , n30517 );
buf ( n234823 , n35431 );
not ( n234824 , n234823 );
or ( n234825 , n234822 , n234824 );
nand ( n234826 , n48436 , n48430 );
not ( n234827 , n234826 );
not ( n234828 , n47689 );
and ( n234829 , n234827 , n234828 );
and ( n234830 , n234826 , n47689 );
nor ( n234831 , n234829 , n234830 );
not ( n234832 , n234831 );
not ( n234833 , n234832 );
not ( n234834 , n234833 );
nand ( n234835 , n226304 , n47563 );
not ( n234836 , n234835 );
not ( n234837 , n47552 );
and ( n234838 , n234836 , n234837 );
and ( n234839 , n234835 , n47552 );
nor ( n234840 , n234838 , n234839 );
not ( n234841 , n234840 );
not ( n234842 , n234427 );
or ( n234843 , n234841 , n234842 );
or ( n234844 , n234427 , n234840 );
nand ( n234845 , n234843 , n234844 );
not ( n234846 , n47689 );
nand ( n234847 , n234846 , n226200 );
not ( n234848 , n234847 );
not ( n234849 , n47679 );
not ( n234850 , n234849 );
and ( n234851 , n234848 , n234850 );
and ( n234852 , n234847 , n234849 );
nor ( n234853 , n234851 , n234852 );
and ( n234854 , n234845 , n234853 );
not ( n234855 , n234845 );
not ( n234856 , n234853 );
and ( n234857 , n234855 , n234856 );
nor ( n234858 , n234854 , n234857 );
not ( n234859 , n225423 );
nand ( n234860 , n234859 , n226284 );
not ( n234861 , n225413 );
xnor ( n234862 , n234860 , n234861 );
not ( n234863 , n234862 );
not ( n234864 , n47733 );
nand ( n234865 , n234864 , n48483 );
not ( n234866 , n234865 );
not ( n234867 , n47723 );
not ( n234868 , n234867 );
and ( n234869 , n234866 , n234868 );
and ( n234870 , n234865 , n234867 );
nor ( n234871 , n234869 , n234870 );
not ( n234872 , n234871 );
or ( n234873 , n234863 , n234872 );
or ( n234874 , n234871 , n234862 );
nand ( n234875 , n234873 , n234874 );
not ( n234876 , n234875 );
and ( n234877 , n234858 , n234876 );
not ( n234878 , n234858 );
and ( n234879 , n234878 , n234875 );
nor ( n234880 , n234877 , n234879 );
not ( n234881 , n234880 );
not ( n234882 , n234881 );
not ( n234883 , n234882 );
or ( n234884 , n234834 , n234883 );
not ( n234885 , n234833 );
nand ( n234886 , n234885 , n234881 );
nand ( n234887 , n234884 , n234886 );
not ( n234888 , n48686 );
not ( n234889 , n234888 );
and ( n234890 , n234887 , n234889 );
not ( n234891 , n234887 );
and ( n234892 , n234891 , n48676 );
nor ( n234893 , n234890 , n234892 );
not ( n234894 , n234893 );
not ( n234895 , n55562 );
not ( n234896 , n204375 );
not ( n234897 , n35017 );
or ( n234898 , n234896 , n234897 );
or ( n234899 , n35017 , n204375 );
nand ( n234900 , n234898 , n234899 );
and ( n234901 , n234900 , n44337 );
not ( n234902 , n234900 );
and ( n234903 , n234902 , n44333 );
nor ( n234904 , n234901 , n234903 );
not ( n234905 , n234904 );
not ( n234906 , n234905 );
not ( n234907 , n234906 );
not ( n234908 , n233315 );
nand ( n234909 , n234908 , n55532 );
not ( n234910 , n234909 );
or ( n234911 , n234907 , n234910 );
or ( n234912 , n234909 , n234906 );
nand ( n234913 , n234911 , n234912 );
not ( n234914 , n234913 );
not ( n234915 , n233360 );
nand ( n234916 , n234915 , n55574 );
not ( n234917 , n31646 );
not ( n234918 , n220127 );
or ( n234919 , n234917 , n234918 );
or ( n234920 , n34643 , n31646 );
nand ( n234921 , n234919 , n234920 );
and ( n234922 , n234921 , n51451 );
not ( n234923 , n234921 );
and ( n234924 , n234923 , n42372 );
nor ( n234925 , n234922 , n234924 );
and ( n234926 , n234916 , n234925 );
not ( n234927 , n234916 );
not ( n234928 , n234925 );
and ( n234929 , n234927 , n234928 );
nor ( n234930 , n234926 , n234929 );
not ( n234931 , n234930 );
or ( n234932 , n234914 , n234931 );
or ( n234933 , n234930 , n234913 );
nand ( n234934 , n234932 , n234933 );
not ( n234935 , n234934 );
not ( n234936 , n233386 );
not ( n234937 , n233393 );
not ( n234938 , n234937 );
not ( n234939 , n33003 );
and ( n234940 , n234938 , n234939 );
and ( n234941 , n234937 , n33003 );
nor ( n234942 , n234940 , n234941 );
nand ( n234943 , n234936 , n234942 );
not ( n234944 , n234943 );
not ( n234945 , n29336 );
not ( n234946 , n31241 );
not ( n234947 , n33195 );
or ( n234948 , n234946 , n234947 );
or ( n234949 , n33195 , n31241 );
nand ( n234950 , n234948 , n234949 );
not ( n234951 , n234950 );
or ( n234952 , n234945 , n234951 );
or ( n234953 , n234950 , n29336 );
nand ( n234954 , n234952 , n234953 );
buf ( n234955 , n234954 );
not ( n234956 , n234955 );
and ( n234957 , n234944 , n234956 );
and ( n234958 , n234943 , n234955 );
nor ( n234959 , n234957 , n234958 );
not ( n234960 , n234959 );
and ( n234961 , n234935 , n234960 );
and ( n234962 , n234934 , n234959 );
nor ( n234963 , n234961 , n234962 );
not ( n234964 , n234963 );
not ( n234965 , n55652 );
not ( n234966 , n55677 );
nand ( n234967 , n234965 , n234966 );
not ( n234968 , n36003 );
not ( n234969 , n45933 );
or ( n234970 , n234968 , n234969 );
nand ( n234971 , n39251 , n35999 );
nand ( n234972 , n234970 , n234971 );
and ( n234973 , n234972 , n45944 );
not ( n234974 , n234972 );
and ( n234975 , n234974 , n222403 );
nor ( n234976 , n234973 , n234975 );
and ( n234977 , n234967 , n234976 );
not ( n234978 , n234967 );
not ( n234979 , n234976 );
and ( n234980 , n234978 , n234979 );
nor ( n234981 , n234977 , n234980 );
not ( n234982 , n234981 );
not ( n234983 , n234982 );
not ( n234984 , n55692 );
nand ( n234985 , n234984 , n55711 );
not ( n234986 , n234985 );
not ( n234987 , n26338 );
not ( n234988 , n32988 );
or ( n234989 , n234987 , n234988 );
nand ( n234990 , n54623 , n26334 );
nand ( n234991 , n234989 , n234990 );
and ( n234992 , n234991 , n45696 );
not ( n234993 , n234991 );
and ( n234994 , n234993 , n41055 );
nor ( n234995 , n234992 , n234994 );
not ( n234996 , n234995 );
and ( n234997 , n234986 , n234996 );
and ( n234998 , n234985 , n234995 );
nor ( n234999 , n234997 , n234998 );
not ( n235000 , n234999 );
or ( n235001 , n234983 , n235000 );
not ( n235002 , n234999 );
nand ( n235003 , n235002 , n234981 );
nand ( n235004 , n235001 , n235003 );
not ( n235005 , n235004 );
and ( n235006 , n234964 , n235005 );
and ( n235007 , n234963 , n235004 );
nor ( n235008 , n235006 , n235007 );
not ( n235009 , n235008 );
or ( n235010 , n234895 , n235009 );
not ( n235011 , n55562 );
not ( n235012 , n235004 );
and ( n235013 , n234963 , n235012 );
not ( n235014 , n234963 );
and ( n235015 , n235014 , n235004 );
nor ( n235016 , n235013 , n235015 );
nand ( n235017 , n235011 , n235016 );
nand ( n235018 , n235010 , n235017 );
buf ( n235019 , n41632 );
and ( n235020 , n235018 , n235019 );
not ( n235021 , n235018 );
not ( n235022 , n235019 );
and ( n235023 , n235021 , n235022 );
nor ( n235024 , n235020 , n235023 );
nand ( n235025 , n234894 , n235024 );
not ( n235026 , n34229 );
nand ( n235027 , n235026 , n234745 );
not ( n235028 , n235027 );
not ( n235029 , n34184 );
not ( n235030 , n235029 );
or ( n235031 , n235028 , n235030 );
or ( n235032 , n235029 , n235027 );
nand ( n235033 , n235031 , n235032 );
not ( n235034 , n235033 );
not ( n235035 , n34439 );
or ( n235036 , n235034 , n235035 );
not ( n235037 , n235033 );
nand ( n235038 , n235037 , n34448 );
nand ( n235039 , n235036 , n235038 );
and ( n235040 , n235039 , n33709 );
not ( n235041 , n235039 );
buf ( n235042 , n55345 );
and ( n235043 , n235041 , n235042 );
nor ( n235044 , n235040 , n235043 );
not ( n235045 , n235044 );
and ( n235046 , n235025 , n235045 );
not ( n235047 , n235025 );
and ( n235048 , n235047 , n235044 );
nor ( n235049 , n235046 , n235048 );
buf ( n235050 , n31571 );
not ( n235051 , n235050 );
not ( n235052 , n235051 );
or ( n235053 , n235049 , n235052 );
nand ( n235054 , n234825 , n235053 );
buf ( n235055 , n235054 );
not ( n235056 , RI19a87dd0_2739);
or ( n235057 , n25328 , n235056 );
not ( n235058 , RI19acc200_2238);
or ( n235059 , n25335 , n235058 );
nand ( n235060 , n235057 , n235059 );
buf ( n235061 , n235060 );
not ( n235062 , RI19ab29b8_2435);
or ( n235063 , n233507 , n235062 );
not ( n235064 , RI19aa8878_2506);
or ( n235065 , n25335 , n235064 );
nand ( n235066 , n235063 , n235065 );
buf ( n235067 , n235066 );
not ( n235068 , n230882 );
not ( n235069 , n42432 );
not ( n235070 , n42321 );
or ( n235071 , n235069 , n235070 );
nand ( n235072 , n235071 , n42435 );
not ( n235073 , n235072 );
or ( n235074 , n235068 , n235073 );
or ( n235075 , n235072 , n230882 );
nand ( n235076 , n235074 , n235075 );
not ( n235077 , n38068 );
not ( n235078 , n30038 );
or ( n235079 , n235077 , n235078 );
or ( n235080 , n30038 , n38068 );
nand ( n235081 , n235079 , n235080 );
xor ( n235082 , n235081 , n42760 );
not ( n235083 , n235082 );
xor ( n235084 , n34231 , n42325 );
xor ( n235085 , n235084 , n29773 );
nand ( n235086 , n235083 , n235085 );
not ( n235087 , n235086 );
not ( n235088 , n43916 );
not ( n235089 , n235088 );
and ( n235090 , n235087 , n235089 );
not ( n235091 , n235082 );
nand ( n235092 , n235085 , n235091 );
and ( n235093 , n235092 , n235088 );
nor ( n235094 , n235090 , n235093 );
not ( n235095 , n235094 );
not ( n235096 , n43870 );
not ( n235097 , n29188 );
not ( n235098 , n207960 );
or ( n235099 , n235097 , n235098 );
not ( n235100 , n29188 );
nand ( n235101 , n235100 , n30205 );
nand ( n235102 , n235099 , n235101 );
and ( n235103 , n235102 , n31832 );
not ( n235104 , n235102 );
not ( n235105 , n31832 );
and ( n235106 , n235104 , n235105 );
nor ( n235107 , n235103 , n235106 );
not ( n235108 , n36038 );
not ( n235109 , n36848 );
or ( n235110 , n235108 , n235109 );
or ( n235111 , n36848 , n36038 );
nand ( n235112 , n235110 , n235111 );
and ( n235113 , n235112 , n36813 );
not ( n235114 , n235112 );
and ( n235115 , n235114 , n39065 );
nor ( n235116 , n235113 , n235115 );
nand ( n235117 , n235107 , n235116 );
not ( n235118 , n235117 );
or ( n235119 , n235096 , n235118 );
or ( n235120 , n235117 , n43870 );
nand ( n235121 , n235119 , n235120 );
not ( n235122 , n235121 );
not ( n235123 , n41055 );
not ( n235124 , n26332 );
not ( n235125 , n32988 );
or ( n235126 , n235124 , n235125 );
not ( n235127 , n26332 );
nand ( n235128 , n235127 , n225593 );
nand ( n235129 , n235126 , n235128 );
not ( n235130 , n235129 );
and ( n235131 , n235123 , n235130 );
and ( n235132 , n41055 , n235129 );
nor ( n235133 , n235131 , n235132 );
not ( n235134 , n28054 );
not ( n235135 , n25385 );
or ( n235136 , n235134 , n235135 );
not ( n235137 , n28054 );
nand ( n235138 , n235137 , n39811 );
nand ( n235139 , n235136 , n235138 );
and ( n235140 , n235139 , n25429 );
not ( n235141 , n235139 );
and ( n235142 , n235141 , n25426 );
nor ( n235143 , n235140 , n235142 );
nand ( n235144 , n235133 , n235143 );
not ( n235145 , n235144 );
not ( n235146 , n43845 );
and ( n235147 , n235145 , n235146 );
and ( n235148 , n235144 , n43845 );
nor ( n235149 , n235147 , n235148 );
not ( n235150 , n235149 );
or ( n235151 , n235122 , n235150 );
or ( n235152 , n235149 , n235121 );
nand ( n235153 , n235151 , n235152 );
not ( n235154 , n235153 );
and ( n235155 , n235095 , n235154 );
and ( n235156 , n235094 , n235153 );
nor ( n235157 , n235155 , n235156 );
not ( n235158 , n43763 );
xor ( n235159 , n209045 , n51033 );
xor ( n235160 , n235159 , n28122 );
nor ( n235161 , n38690 , n31489 );
not ( n235162 , n235161 );
nand ( n235163 , n38690 , n31489 );
nand ( n235164 , n235162 , n235163 );
and ( n235165 , n235164 , n37192 );
not ( n235166 , n235164 );
and ( n235167 , n235166 , n38795 );
nor ( n235168 , n235165 , n235167 );
nand ( n235169 , n235160 , n235168 );
not ( n235170 , n235169 );
or ( n235171 , n235158 , n235170 );
or ( n235172 , n235169 , n43763 );
nand ( n235173 , n235171 , n235172 );
not ( n235174 , n235173 );
xor ( n235175 , n34787 , n29162 );
xnor ( n235176 , n235175 , n44690 );
and ( n235177 , n38646 , n40267 );
not ( n235178 , n38646 );
and ( n235179 , n235178 , n220432 );
or ( n235180 , n235177 , n235179 );
and ( n235181 , n235180 , n42681 );
not ( n235182 , n235180 );
and ( n235183 , n235182 , n40273 );
nor ( n235184 , n235181 , n235183 );
nand ( n235185 , n235176 , n235184 );
not ( n235186 , n235185 );
not ( n235187 , n43792 );
and ( n235188 , n235186 , n235187 );
not ( n235189 , n235184 );
not ( n235190 , n235189 );
nand ( n235191 , n235190 , n235176 );
and ( n235192 , n235191 , n43792 );
nor ( n235193 , n235188 , n235192 );
not ( n235194 , n235193 );
or ( n235195 , n235174 , n235194 );
or ( n235196 , n235193 , n235173 );
nand ( n235197 , n235195 , n235196 );
and ( n235198 , n235157 , n235197 );
not ( n235199 , n235157 );
not ( n235200 , n235197 );
and ( n235201 , n235199 , n235200 );
nor ( n235202 , n235198 , n235201 );
buf ( n235203 , n235202 );
and ( n235204 , n235076 , n235203 );
not ( n235205 , n235076 );
not ( n235206 , n235200 );
not ( n235207 , n235157 );
not ( n235208 , n235207 );
or ( n235209 , n235206 , n235208 );
nand ( n235210 , n235157 , n235197 );
nand ( n235211 , n235209 , n235210 );
and ( n235212 , n235205 , n235211 );
nor ( n235213 , n235204 , n235212 );
not ( n235214 , n235213 );
not ( n235215 , n235214 );
not ( n235216 , n220347 );
not ( n235217 , n213041 );
or ( n235218 , n235216 , n235217 );
not ( n235219 , n220347 );
nand ( n235220 , n235219 , n215580 );
nand ( n235221 , n235218 , n235220 );
and ( n235222 , n235221 , n43326 );
not ( n235223 , n235221 );
and ( n235224 , n235223 , n51231 );
nor ( n235225 , n235222 , n235224 );
not ( n235226 , n235225 );
nand ( n235227 , n44654 , n235226 );
not ( n235228 , n235227 );
not ( n235229 , n33442 );
not ( n235230 , n44823 );
or ( n235231 , n235229 , n235230 );
or ( n235232 , n44823 , n33442 );
nand ( n235233 , n235231 , n235232 );
and ( n235234 , n235233 , n226156 );
not ( n235235 , n235233 );
and ( n235236 , n235235 , n32363 );
nor ( n235237 , n235234 , n235236 );
not ( n235238 , n235237 );
and ( n235239 , n235228 , n235238 );
and ( n235240 , n235227 , n235237 );
nor ( n235241 , n235239 , n235240 );
not ( n235242 , n235241 );
not ( n235243 , n235242 );
not ( n235244 , n205143 );
buf ( n235245 , n35820 );
and ( n235246 , n235245 , n37229 );
not ( n235247 , n235245 );
and ( n235248 , n235247 , n205134 );
nor ( n235249 , n235246 , n235248 );
not ( n235250 , n235249 );
not ( n235251 , n235250 );
or ( n235252 , n235244 , n235251 );
nand ( n235253 , n205096 , n235249 );
nand ( n235254 , n235252 , n235253 );
not ( n235255 , n35589 );
not ( n235256 , n40523 );
or ( n235257 , n235255 , n235256 );
not ( n235258 , n35589 );
nand ( n235259 , n235258 , n41040 );
nand ( n235260 , n235257 , n235259 );
and ( n235261 , n235260 , n40564 );
not ( n235262 , n235260 );
and ( n235263 , n235262 , n44785 );
nor ( n235264 , n235261 , n235263 );
nand ( n235265 , n235254 , n235264 );
not ( n235266 , n235265 );
not ( n235267 , n44604 );
and ( n235268 , n235266 , n235267 );
and ( n235269 , n235265 , n44604 );
nor ( n235270 , n235268 , n235269 );
buf ( n235271 , n38433 );
not ( n235272 , n235271 );
not ( n235273 , n41017 );
not ( n235274 , n235273 );
or ( n235275 , n235272 , n235274 );
or ( n235276 , n235273 , n235271 );
nand ( n235277 , n235275 , n235276 );
not ( n235278 , n235277 );
not ( n235279 , n213924 );
or ( n235280 , n235278 , n235279 );
or ( n235281 , n36168 , n235277 );
nand ( n235282 , n235280 , n235281 );
not ( n235283 , n235282 );
not ( n235284 , n30537 );
not ( n235285 , n36519 );
not ( n235286 , n26204 );
or ( n235287 , n235285 , n235286 );
or ( n235288 , n26204 , n36519 );
nand ( n235289 , n235287 , n235288 );
not ( n235290 , n235289 );
or ( n235291 , n235284 , n235290 );
or ( n235292 , n235289 , n30534 );
nand ( n235293 , n235291 , n235292 );
nand ( n235294 , n235283 , n235293 );
and ( n235295 , n235294 , n44722 );
not ( n235296 , n235294 );
and ( n235297 , n235296 , n44723 );
nor ( n235298 , n235295 , n235297 );
xor ( n235299 , n235270 , n235298 );
buf ( n235300 , n27714 );
xor ( n235301 , n235300 , n222033 );
xnor ( n235302 , n235301 , n25457 );
not ( n235303 , n235302 );
not ( n235304 , n34103 );
buf ( n235305 , n204885 );
nor ( n235306 , n34051 , n235305 );
not ( n235307 , n235306 );
nand ( n235308 , n34051 , n235305 );
nand ( n235309 , n235307 , n235308 );
not ( n235310 , n235309 );
or ( n235311 , n235304 , n235310 );
or ( n235312 , n235309 , n34104 );
nand ( n235313 , n235311 , n235312 );
not ( n235314 , n235313 );
nand ( n235315 , n235303 , n235314 );
and ( n235316 , n235315 , n44700 );
not ( n235317 , n235315 );
and ( n235318 , n235317 , n222462 );
nor ( n235319 , n235316 , n235318 );
xnor ( n235320 , n235299 , n235319 );
not ( n235321 , n44630 );
nor ( n235322 , n235237 , n235226 );
not ( n235323 , n235322 );
and ( n235324 , n235321 , n235323 );
nor ( n235325 , n235237 , n235226 );
and ( n235326 , n44630 , n235325 );
nor ( n235327 , n235324 , n235326 );
not ( n235328 , n38436 );
xor ( n235329 , n29522 , n235328 );
xnor ( n235330 , n235329 , n220965 );
not ( n235331 , n204977 );
buf ( n235332 , n38961 );
not ( n235333 , n235332 );
not ( n235334 , n46681 );
or ( n235335 , n235333 , n235334 );
or ( n235336 , n46681 , n235332 );
nand ( n235337 , n235335 , n235336 );
not ( n235338 , n235337 );
or ( n235339 , n235331 , n235338 );
or ( n235340 , n235337 , n204981 );
nand ( n235341 , n235339 , n235340 );
nand ( n235342 , n235330 , n235341 );
not ( n235343 , n222339 );
and ( n235344 , n235342 , n235343 );
not ( n235345 , n235342 );
and ( n235346 , n235345 , n222339 );
nor ( n235347 , n235344 , n235346 );
and ( n235348 , n235327 , n235347 );
not ( n235349 , n235327 );
not ( n235350 , n235347 );
and ( n235351 , n235349 , n235350 );
nor ( n235352 , n235348 , n235351 );
and ( n235353 , n235320 , n235352 );
not ( n235354 , n235320 );
not ( n235355 , n235352 );
and ( n235356 , n235354 , n235355 );
nor ( n235357 , n235353 , n235356 );
not ( n235358 , n235357 );
or ( n235359 , n235243 , n235358 );
not ( n235360 , n235242 );
not ( n235361 , n235352 );
not ( n235362 , n235320 );
or ( n235363 , n235361 , n235362 );
not ( n235364 , n235320 );
nand ( n235365 , n235364 , n235355 );
nand ( n235366 , n235363 , n235365 );
nand ( n235367 , n235360 , n235366 );
nand ( n235368 , n235359 , n235367 );
buf ( n235369 , n46941 );
and ( n235370 , n235368 , n235369 );
not ( n235371 , n235368 );
buf ( n235372 , n46950 );
and ( n235373 , n235371 , n235372 );
nor ( n235374 , n235370 , n235373 );
not ( n235375 , n235374 );
or ( n235376 , n235215 , n235375 );
nand ( n235377 , n235376 , n226010 );
buf ( n235378 , n28451 );
not ( n235379 , n235378 );
not ( n235380 , n34338 );
or ( n235381 , n235379 , n235380 );
or ( n235382 , n34338 , n235378 );
nand ( n235383 , n235381 , n235382 );
not ( n235384 , n235383 );
not ( n235385 , n32863 );
or ( n235386 , n235384 , n235385 );
or ( n235387 , n32863 , n235383 );
nand ( n235388 , n235386 , n235387 );
not ( n235389 , n235388 );
not ( n235390 , n35621 );
not ( n235391 , n235390 );
not ( n235392 , n35740 );
or ( n235393 , n235391 , n235392 );
or ( n235394 , n35740 , n235390 );
nand ( n235395 , n235393 , n235394 );
and ( n235396 , n235395 , n206976 );
not ( n235397 , n235395 );
and ( n235398 , n235397 , n29214 );
nor ( n235399 , n235396 , n235398 );
not ( n235400 , n235399 );
nand ( n235401 , n235389 , n235400 );
not ( n235402 , n26207 );
not ( n235403 , n33564 );
or ( n235404 , n235402 , n235403 );
not ( n235405 , n26207 );
nand ( n235406 , n235405 , n48779 );
nand ( n235407 , n235404 , n235406 );
and ( n235408 , n235407 , n36620 );
not ( n235409 , n235407 );
and ( n235410 , n235409 , n51936 );
nor ( n235411 , n235408 , n235410 );
buf ( n235412 , n235411 );
not ( n235413 , n235412 );
and ( n235414 , n235401 , n235413 );
not ( n235415 , n235401 );
and ( n235416 , n235415 , n235412 );
nor ( n235417 , n235414 , n235416 );
not ( n235418 , n235417 );
not ( n235419 , n235411 );
nand ( n235420 , n235388 , n235419 );
not ( n235421 , n235420 );
not ( n235422 , n208049 );
not ( n235423 , n222865 );
or ( n235424 , n235422 , n235423 );
not ( n235425 , n208049 );
nand ( n235426 , n235425 , n41148 );
nand ( n235427 , n235424 , n235426 );
and ( n235428 , n235427 , n218917 );
not ( n235429 , n235427 );
not ( n235430 , n218917 );
and ( n235431 , n235429 , n235430 );
nor ( n235432 , n235428 , n235431 );
not ( n235433 , n235432 );
not ( n235434 , n235433 );
not ( n235435 , n235434 );
and ( n235436 , n235421 , n235435 );
and ( n235437 , n235420 , n235434 );
nor ( n235438 , n235436 , n235437 );
not ( n235439 , n235438 );
not ( n235440 , n235439 );
xor ( n235441 , n36324 , n41894 );
xnor ( n235442 , n235441 , n53512 );
not ( n235443 , n221597 );
not ( n235444 , n235443 );
not ( n235445 , n49568 );
or ( n235446 , n235444 , n235445 );
nand ( n235447 , n41754 , n221597 );
nand ( n235448 , n235446 , n235447 );
not ( n235449 , n235448 );
not ( n235450 , n228145 );
and ( n235451 , n235449 , n235450 );
and ( n235452 , n228145 , n235448 );
nor ( n235453 , n235451 , n235452 );
not ( n235454 , n235453 );
nand ( n235455 , n235442 , n235454 );
not ( n235456 , n207930 );
not ( n235457 , n205476 );
or ( n235458 , n235456 , n235457 );
or ( n235459 , n205476 , n207930 );
nand ( n235460 , n235458 , n235459 );
and ( n235461 , n235460 , n27759 );
not ( n235462 , n235460 );
and ( n235463 , n235462 , n27763 );
nor ( n235464 , n235461 , n235463 );
and ( n235465 , n235455 , n235464 );
not ( n235466 , n235455 );
not ( n235467 , n235464 );
and ( n235468 , n235466 , n235467 );
nor ( n235469 , n235465 , n235468 );
not ( n235470 , n235469 );
not ( n235471 , n235470 );
or ( n235472 , n235440 , n235471 );
nand ( n235473 , n235469 , n235438 );
nand ( n235474 , n235472 , n235473 );
xor ( n235475 , n30280 , n37212 );
xnor ( n235476 , n235475 , n204632 );
buf ( n235477 , RI17450370_1345);
not ( n235478 , n235477 );
not ( n235479 , n36411 );
or ( n235480 , n235478 , n235479 );
nand ( n235481 , n36415 , n33266 );
nand ( n235482 , n235480 , n235481 );
and ( n235483 , n235482 , n26047 );
not ( n235484 , n235482 );
and ( n235485 , n235484 , n35028 );
nor ( n235486 , n235483 , n235485 );
nand ( n235487 , n235476 , n235486 );
not ( n235488 , n235487 );
not ( n235489 , n33816 );
not ( n235490 , n38795 );
or ( n235491 , n235489 , n235490 );
or ( n235492 , n38795 , n33816 );
nand ( n235493 , n235491 , n235492 );
xor ( n235494 , n235493 , n38802 );
not ( n235495 , n235494 );
and ( n235496 , n235488 , n235495 );
and ( n235497 , n235487 , n235494 );
nor ( n235498 , n235496 , n235497 );
and ( n235499 , n235474 , n235498 );
not ( n235500 , n235474 );
not ( n235501 , n235498 );
and ( n235502 , n235500 , n235501 );
nor ( n235503 , n235499 , n235502 );
not ( n235504 , n235503 );
buf ( n235505 , RI17405a78_1480);
not ( n235506 , n235505 );
not ( n235507 , n40564 );
or ( n235508 , n235506 , n235507 );
nand ( n235509 , n40569 , n35534 );
nand ( n235510 , n235508 , n235509 );
and ( n235511 , n235510 , n29525 );
not ( n235512 , n235510 );
and ( n235513 , n235512 , n29519 );
nor ( n235514 , n235511 , n235513 );
not ( n235515 , n235514 );
xor ( n235516 , n25699 , n30582 );
xnor ( n235517 , n235516 , n30608 );
not ( n235518 , n235517 );
buf ( n235519 , n32846 );
not ( n235520 , n235519 );
not ( n235521 , n222753 );
or ( n235522 , n235520 , n235521 );
or ( n235523 , n222753 , n235519 );
nand ( n235524 , n235522 , n235523 );
and ( n235525 , n235524 , n37533 );
not ( n235526 , n235524 );
and ( n235527 , n235526 , n37539 );
nor ( n235528 , n235525 , n235527 );
not ( n235529 , n235528 );
nand ( n235530 , n235518 , n235529 );
not ( n235531 , n235530 );
or ( n235532 , n235515 , n235531 );
not ( n235533 , n235528 );
nand ( n235534 , n235533 , n235518 );
or ( n235535 , n235534 , n235514 );
nand ( n235536 , n235532 , n235535 );
not ( n235537 , n235536 );
not ( n235538 , RI174a6590_925);
and ( n235539 , n28144 , n235538 );
not ( n235540 , n28144 );
and ( n235541 , n235540 , n205902 );
nor ( n235542 , n235539 , n235541 );
xor ( n235543 , n235542 , n52070 );
xnor ( n235544 , n235543 , n224859 );
not ( n235545 , n235544 );
not ( n235546 , n46815 );
not ( n235547 , n31365 );
and ( n235548 , n235546 , n235547 );
and ( n235549 , n46815 , n31365 );
nor ( n235550 , n235548 , n235549 );
not ( n235551 , n235550 );
not ( n235552 , n40066 );
or ( n235553 , n235551 , n235552 );
or ( n235554 , n40066 , n235550 );
nand ( n235555 , n235553 , n235554 );
not ( n235556 , n235555 );
nand ( n235557 , n235545 , n235556 );
not ( n235558 , n235557 );
not ( n235559 , n36488 );
not ( n235560 , n47879 );
or ( n235561 , n235559 , n235560 );
or ( n235562 , n47879 , n36488 );
nand ( n235563 , n235561 , n235562 );
and ( n235564 , n235563 , n40231 );
not ( n235565 , n235563 );
and ( n235566 , n235565 , n40234 );
nor ( n235567 , n235564 , n235566 );
not ( n235568 , n235567 );
not ( n235569 , n235568 );
and ( n235570 , n235558 , n235569 );
and ( n235571 , n235557 , n235568 );
nor ( n235572 , n235570 , n235571 );
not ( n235573 , n235572 );
or ( n235574 , n235537 , n235573 );
or ( n235575 , n235536 , n235572 );
nand ( n235576 , n235574 , n235575 );
not ( n235577 , n235576 );
and ( n235578 , n235504 , n235577 );
and ( n235579 , n235503 , n235576 );
nor ( n235580 , n235578 , n235579 );
not ( n235581 , n235580 );
or ( n235582 , n235418 , n235581 );
not ( n235583 , n235417 );
not ( n235584 , n235503 );
not ( n235585 , n235584 );
not ( n235586 , n235576 );
not ( n235587 , n235586 );
or ( n235588 , n235585 , n235587 );
nand ( n235589 , n235503 , n235576 );
nand ( n235590 , n235588 , n235589 );
nand ( n235591 , n235583 , n235590 );
nand ( n235592 , n235582 , n235591 );
not ( n235593 , n50957 );
not ( n235594 , n25935 );
not ( n235595 , n32006 );
or ( n235596 , n235594 , n235595 );
or ( n235597 , n32006 , n25935 );
nand ( n235598 , n235596 , n235597 );
and ( n235599 , n235598 , n42057 );
not ( n235600 , n235598 );
and ( n235601 , n235600 , n42058 );
nor ( n235602 , n235599 , n235601 );
nand ( n235603 , n50968 , n235602 );
not ( n235604 , n235603 );
and ( n235605 , n235593 , n235604 );
and ( n235606 , n50957 , n235603 );
nor ( n235607 , n235605 , n235606 );
not ( n235608 , n235607 );
not ( n235609 , n32935 );
not ( n235610 , n26008 );
or ( n235611 , n235609 , n235610 );
or ( n235612 , n26008 , n32935 );
nand ( n235613 , n235611 , n235612 );
and ( n235614 , n235613 , n231142 );
not ( n235615 , n235613 );
and ( n235616 , n235615 , n29913 );
nor ( n235617 , n235614 , n235616 );
not ( n235618 , n235617 );
not ( n235619 , n206723 );
not ( n235620 , n30321 );
or ( n235621 , n235619 , n235620 );
or ( n235622 , n30321 , n206723 );
nand ( n235623 , n235621 , n235622 );
and ( n235624 , n235623 , n204436 );
not ( n235625 , n235623 );
and ( n235626 , n235625 , n41785 );
nor ( n235627 , n235624 , n235626 );
nand ( n235628 , n235618 , n235627 );
not ( n235629 , n50995 );
and ( n235630 , n235628 , n235629 );
not ( n235631 , n235628 );
and ( n235632 , n235631 , n50995 );
nor ( n235633 , n235630 , n235632 );
not ( n235634 , n235633 );
or ( n235635 , n235608 , n235634 );
or ( n235636 , n235633 , n235607 );
nand ( n235637 , n235635 , n235636 );
buf ( n235638 , n31375 );
and ( n235639 , n235638 , n46816 );
not ( n235640 , n235638 );
and ( n235641 , n235640 , n217819 );
nor ( n235642 , n235639 , n235641 );
not ( n235643 , n235642 );
not ( n235644 , n40066 );
or ( n235645 , n235643 , n235644 );
or ( n235646 , n40066 , n235642 );
nand ( n235647 , n235645 , n235646 );
not ( n235648 , n235647 );
not ( n235649 , n207116 );
not ( n235650 , n31514 );
or ( n235651 , n235649 , n235650 );
not ( n235652 , n207116 );
nand ( n235653 , n235652 , n31527 );
nand ( n235654 , n235651 , n235653 );
and ( n235655 , n235654 , n33853 );
not ( n235656 , n235654 );
and ( n235657 , n235656 , n33849 );
nor ( n235658 , n235655 , n235657 );
nand ( n235659 , n235648 , n235658 );
not ( n235660 , n228796 );
xor ( n235661 , n235659 , n235660 );
and ( n235662 , n235637 , n235661 );
not ( n235663 , n235637 );
not ( n235664 , n235661 );
and ( n235665 , n235663 , n235664 );
nor ( n235666 , n235662 , n235665 );
not ( n235667 , n51131 );
buf ( n235668 , n34087 );
xor ( n235669 , n235668 , n55938 );
xnor ( n235670 , n235669 , n41258 );
not ( n235671 , n38334 );
not ( n235672 , n32323 );
or ( n235673 , n235671 , n235672 );
or ( n235674 , n32323 , n38334 );
nand ( n235675 , n235673 , n235674 );
xor ( n235676 , n235675 , n37398 );
not ( n235677 , n235676 );
nand ( n235678 , n235670 , n235677 );
not ( n235679 , n235678 );
or ( n235680 , n235667 , n235679 );
or ( n235681 , n235678 , n51131 );
nand ( n235682 , n235680 , n235681 );
not ( n235683 , n235682 );
not ( n235684 , n37001 );
not ( n235685 , n41593 );
or ( n235686 , n235684 , n235685 );
or ( n235687 , n45702 , n37001 );
nand ( n235688 , n235686 , n235687 );
and ( n235689 , n235688 , n36093 );
not ( n235690 , n235688 );
and ( n235691 , n235690 , n44712 );
nor ( n235692 , n235689 , n235691 );
not ( n235693 , n235692 );
not ( n235694 , n35582 );
not ( n235695 , n41040 );
or ( n235696 , n235694 , n235695 );
not ( n235697 , n44779 );
or ( n235698 , n235697 , n35582 );
nand ( n235699 , n235696 , n235698 );
and ( n235700 , n235699 , n222549 );
not ( n235701 , n235699 );
and ( n235702 , n235701 , n44785 );
nor ( n235703 , n235700 , n235702 );
nand ( n235704 , n235693 , n235703 );
not ( n235705 , n235704 );
not ( n235706 , n51099 );
and ( n235707 , n235705 , n235706 );
and ( n235708 , n235704 , n51099 );
nor ( n235709 , n235707 , n235708 );
not ( n235710 , n235709 );
and ( n235711 , n235683 , n235710 );
and ( n235712 , n235682 , n235709 );
nor ( n235713 , n235711 , n235712 );
and ( n235714 , n235666 , n235713 );
not ( n235715 , n235666 );
not ( n235716 , n235713 );
and ( n235717 , n235715 , n235716 );
nor ( n235718 , n235714 , n235717 );
not ( n235719 , n235718 );
not ( n235720 , n235719 );
and ( n235721 , n235592 , n235720 );
not ( n235722 , n235592 );
not ( n235723 , n235716 );
not ( n235724 , n235666 );
not ( n235725 , n235724 );
or ( n235726 , n235723 , n235725 );
nand ( n235727 , n235666 , n235713 );
nand ( n235728 , n235726 , n235727 );
and ( n235729 , n235722 , n235728 );
nor ( n235730 , n235721 , n235729 );
or ( n235731 , n235377 , n235730 );
buf ( n235732 , n33252 );
nor ( n235733 , n235213 , n235732 );
nand ( n235734 , n235374 , n235733 , n235730 );
nand ( n235735 , n39766 , n34054 );
nand ( n235736 , n235731 , n235734 , n235735 );
buf ( n235737 , n235736 );
buf ( n235738 , RI19a25298_2780);
and ( n235739 , n25326 , n235738 );
buf ( n235740 , n235739 );
not ( n235741 , n55069 );
not ( n235742 , n39886 );
not ( n235743 , n39923 );
nand ( n235744 , n235743 , n40011 );
and ( n235745 , n235744 , n52489 );
not ( n235746 , n235744 );
and ( n235747 , n235746 , n52490 );
nor ( n235748 , n235745 , n235747 );
not ( n235749 , n235748 );
not ( n235750 , n235749 );
not ( n235751 , n40068 );
not ( n235752 , n40080 );
nand ( n235753 , n235751 , n235752 );
not ( n235754 , n235753 );
not ( n235755 , n52542 );
and ( n235756 , n235754 , n235755 );
and ( n235757 , n235753 , n52542 );
nor ( n235758 , n235756 , n235757 );
not ( n235759 , n235758 );
not ( n235760 , n235759 );
or ( n235761 , n235750 , n235760 );
nand ( n235762 , n235758 , n235748 );
nand ( n235763 , n235761 , n235762 );
not ( n235764 , n40180 );
not ( n235765 , n217935 );
nand ( n235766 , n235764 , n235765 );
not ( n235767 , n52526 );
and ( n235768 , n235766 , n235767 );
not ( n235769 , n235766 );
not ( n235770 , n235767 );
and ( n235771 , n235769 , n235770 );
nor ( n235772 , n235768 , n235771 );
and ( n235773 , n235763 , n235772 );
not ( n235774 , n235763 );
not ( n235775 , n235772 );
and ( n235776 , n235774 , n235775 );
nor ( n235777 , n235773 , n235776 );
not ( n235778 , n235777 );
not ( n235779 , n235778 );
not ( n235780 , n39880 );
not ( n235781 , n39780 );
nand ( n235782 , n235780 , n235781 );
not ( n235783 , n235782 );
not ( n235784 , n52561 );
and ( n235785 , n235783 , n235784 );
not ( n235786 , n39880 );
nand ( n235787 , n235786 , n235781 );
and ( n235788 , n235787 , n52561 );
nor ( n235789 , n235785 , n235788 );
not ( n235790 , n235789 );
not ( n235791 , n230339 );
not ( n235792 , n39826 );
nand ( n235793 , n235792 , n39863 );
not ( n235794 , n235793 );
or ( n235795 , n235791 , n235794 );
nand ( n235796 , n235792 , n39863 );
or ( n235797 , n235796 , n230339 );
nand ( n235798 , n235795 , n235797 );
not ( n235799 , n235798 );
and ( n235800 , n235790 , n235799 );
and ( n235801 , n235789 , n235798 );
nor ( n235802 , n235800 , n235801 );
not ( n235803 , n235802 );
not ( n235804 , n235803 );
and ( n235805 , n235779 , n235804 );
and ( n235806 , n235778 , n235803 );
nor ( n235807 , n235805 , n235806 );
not ( n235808 , n235807 );
or ( n235809 , n235742 , n235808 );
not ( n235810 , n39886 );
not ( n235811 , n235777 );
not ( n235812 , n235802 );
or ( n235813 , n235811 , n235812 );
nand ( n235814 , n235778 , n235803 );
nand ( n235815 , n235813 , n235814 );
nand ( n235816 , n235810 , n235815 );
nand ( n235817 , n235809 , n235816 );
not ( n235818 , n217981 );
not ( n235819 , n40246 );
nand ( n235820 , n235818 , n235819 );
not ( n235821 , n235820 );
not ( n235822 , n230422 );
and ( n235823 , n235821 , n235822 );
and ( n235824 , n235820 , n230422 );
nor ( n235825 , n235823 , n235824 );
not ( n235826 , n235825 );
not ( n235827 , n235826 );
not ( n235828 , n40275 );
nand ( n235829 , n40289 , n235828 );
not ( n235830 , n235829 );
not ( n235831 , n230434 );
or ( n235832 , n235830 , n235831 );
or ( n235833 , n230434 , n235829 );
nand ( n235834 , n235832 , n235833 );
not ( n235835 , n235834 );
not ( n235836 , n235835 );
or ( n235837 , n235827 , n235836 );
nand ( n235838 , n235834 , n235825 );
nand ( n235839 , n235837 , n235838 );
not ( n235840 , n40331 );
not ( n235841 , n40311 );
nand ( n235842 , n235840 , n235841 );
buf ( n235843 , n52637 );
and ( n235844 , n235842 , n235843 );
not ( n235845 , n235842 );
not ( n235846 , n235843 );
and ( n235847 , n235845 , n235846 );
nor ( n235848 , n235844 , n235847 );
and ( n235849 , n235839 , n235848 );
not ( n235850 , n235839 );
not ( n235851 , n235848 );
and ( n235852 , n235850 , n235851 );
nor ( n235853 , n235849 , n235852 );
not ( n235854 , n40446 );
not ( n235855 , n40416 );
nand ( n235856 , n235854 , n235855 );
not ( n235857 , n235856 );
not ( n235858 , n52739 );
and ( n235859 , n235857 , n235858 );
and ( n235860 , n235856 , n52739 );
nor ( n235861 , n235859 , n235860 );
not ( n235862 , n235861 );
not ( n235863 , n40361 );
nand ( n235864 , n235863 , n40375 );
not ( n235865 , n235864 );
not ( n235866 , n230459 );
or ( n235867 , n235865 , n235866 );
or ( n235868 , n230459 , n235864 );
nand ( n235869 , n235867 , n235868 );
not ( n235870 , n235869 );
and ( n235871 , n235862 , n235870 );
and ( n235872 , n235861 , n235869 );
nor ( n235873 , n235871 , n235872 );
and ( n235874 , n235853 , n235873 );
not ( n235875 , n235853 );
not ( n235876 , n235873 );
and ( n235877 , n235875 , n235876 );
nor ( n235878 , n235874 , n235877 );
buf ( n235879 , n235878 );
and ( n235880 , n235817 , n235879 );
not ( n235881 , n235817 );
not ( n235882 , n235873 );
not ( n235883 , n235853 );
or ( n235884 , n235882 , n235883 );
not ( n235885 , n235853 );
nand ( n235886 , n235885 , n235876 );
nand ( n235887 , n235884 , n235886 );
buf ( n235888 , n235887 );
and ( n235889 , n235881 , n235888 );
nor ( n235890 , n235880 , n235889 );
not ( n235891 , n235890 );
nand ( n235892 , n235741 , n235891 );
not ( n235893 , n232870 );
or ( n235894 , n235892 , n235893 );
not ( n235895 , n205649 );
nor ( n235896 , n54765 , n235895 );
nand ( n235897 , n235892 , n235896 );
nand ( n235898 , n49054 , n29600 );
nand ( n235899 , n235894 , n235897 , n235898 );
buf ( n235900 , n235899 );
buf ( n235901 , n206564 );
buf ( n235902 , n38457 );
not ( n235903 , RI19ac1490_2320);
or ( n235904 , n226819 , n235903 );
not ( n235905 , RI19ab8b38_2390);
or ( n235906 , n25335 , n235905 );
nand ( n235907 , n235904 , n235906 );
buf ( n235908 , n235907 );
buf ( n235909 , n32306 );
not ( n235910 , n28435 );
not ( n235911 , n55760 );
or ( n235912 , n235910 , n235911 );
not ( n235913 , n25899 );
not ( n235914 , n209733 );
or ( n235915 , n235913 , n235914 );
not ( n235916 , n25899 );
nand ( n235917 , n235916 , n31967 );
nand ( n235918 , n235915 , n235917 );
and ( n235919 , n235918 , n32007 );
not ( n235920 , n235918 );
and ( n235921 , n235920 , n35624 );
nor ( n235922 , n235919 , n235921 );
nand ( n235923 , n50215 , n235922 );
not ( n235924 , n235923 );
not ( n235925 , n30613 );
not ( n235926 , n54667 );
or ( n235927 , n235925 , n235926 );
or ( n235928 , n54667 , n30613 );
nand ( n235929 , n235927 , n235928 );
not ( n235930 , n49132 );
and ( n235931 , n235929 , n235930 );
not ( n235932 , n235929 );
not ( n235933 , n47607 );
and ( n235934 , n235932 , n235933 );
nor ( n235935 , n235931 , n235934 );
not ( n235936 , n235935 );
not ( n235937 , n235936 );
and ( n235938 , n235924 , n235937 );
and ( n235939 , n235923 , n235936 );
nor ( n235940 , n235938 , n235939 );
not ( n235941 , n235940 );
not ( n235942 , n235941 );
not ( n235943 , n50192 );
not ( n235944 , n235922 );
nand ( n235945 , n235944 , n235935 );
not ( n235946 , n235945 );
or ( n235947 , n235943 , n235946 );
or ( n235948 , n235945 , n50192 );
nand ( n235949 , n235947 , n235948 );
not ( n235950 , n235949 );
not ( n235951 , n205230 );
not ( n235952 , n37148 );
not ( n235953 , n205236 );
or ( n235954 , n235952 , n235953 );
or ( n235955 , n205236 , n37148 );
nand ( n235956 , n235954 , n235955 );
not ( n235957 , n235956 );
and ( n235958 , n235951 , n235957 );
and ( n235959 , n205230 , n235956 );
nor ( n235960 , n235958 , n235959 );
not ( n235961 , n41891 );
not ( n235962 , n44974 );
not ( n235963 , n25735 );
and ( n235964 , n235962 , n235963 );
and ( n235965 , n44974 , n25735 );
nor ( n235966 , n235964 , n235965 );
not ( n235967 , n235966 );
and ( n235968 , n235961 , n235967 );
and ( n235969 , n41891 , n235966 );
nor ( n235970 , n235968 , n235969 );
not ( n235971 , n235970 );
nand ( n235972 , n235960 , n235971 );
and ( n235973 , n235972 , n50242 );
not ( n235974 , n235972 );
and ( n235975 , n235974 , n50241 );
nor ( n235976 , n235973 , n235975 );
not ( n235977 , n235976 );
or ( n235978 , n235950 , n235977 );
or ( n235979 , n235949 , n235976 );
nand ( n235980 , n235978 , n235979 );
not ( n235981 , n235980 );
xor ( n235982 , n33386 , n38844 );
xnor ( n235983 , n235982 , n38570 );
not ( n235984 , n235983 );
not ( n235985 , n227821 );
nand ( n235986 , n235984 , n235985 );
not ( n235987 , n235986 );
not ( n235988 , n50079 );
and ( n235989 , n235987 , n235988 );
and ( n235990 , n235986 , n50079 );
nor ( n235991 , n235989 , n235990 );
not ( n235992 , n235991 );
and ( n235993 , n235981 , n235992 );
and ( n235994 , n235980 , n235991 );
nor ( n235995 , n235993 , n235994 );
not ( n235996 , n50155 );
not ( n235997 , n35584 );
not ( n235998 , n31686 );
not ( n235999 , n26408 );
or ( n236000 , n235998 , n235999 );
or ( n236001 , n26408 , n31686 );
nand ( n236002 , n236000 , n236001 );
not ( n236003 , n236002 );
or ( n236004 , n235997 , n236003 );
or ( n236005 , n236002 , n53432 );
nand ( n236006 , n236004 , n236005 );
not ( n236007 , n236006 );
xor ( n236008 , n208141 , n48174 );
xnor ( n236009 , n236008 , n39532 );
not ( n236010 , n236009 );
nand ( n236011 , n236007 , n236010 );
not ( n236012 , n236011 );
or ( n236013 , n235996 , n236012 );
not ( n236014 , n236006 );
nand ( n236015 , n236014 , n236010 );
or ( n236016 , n236015 , n50155 );
nand ( n236017 , n236013 , n236016 );
not ( n236018 , n236017 );
not ( n236019 , n34776 );
not ( n236020 , n29117 );
or ( n236021 , n236019 , n236020 );
not ( n236022 , n34776 );
nand ( n236023 , n236022 , n29123 );
nand ( n236024 , n236021 , n236023 );
and ( n236025 , n236024 , n29162 );
not ( n236026 , n236024 );
and ( n236027 , n236026 , n29175 );
nor ( n236028 , n236025 , n236027 );
not ( n236029 , n236028 );
not ( n236030 , n42500 );
not ( n236031 , n41723 );
or ( n236032 , n236030 , n236031 );
or ( n236033 , n41723 , n42500 );
nand ( n236034 , n236032 , n236033 );
and ( n236035 , n236034 , n42355 );
not ( n236036 , n236034 );
not ( n236037 , n227330 );
and ( n236038 , n236036 , n236037 );
nor ( n236039 , n236035 , n236038 );
not ( n236040 , n236039 );
nand ( n236041 , n236029 , n236040 );
and ( n236042 , n236041 , n227874 );
not ( n236043 , n236041 );
not ( n236044 , n227874 );
and ( n236045 , n236043 , n236044 );
nor ( n236046 , n236042 , n236045 );
not ( n236047 , n236046 );
and ( n236048 , n236018 , n236047 );
and ( n236049 , n236017 , n236046 );
nor ( n236050 , n236048 , n236049 );
and ( n236051 , n235995 , n236050 );
not ( n236052 , n235995 );
not ( n236053 , n236050 );
and ( n236054 , n236052 , n236053 );
nor ( n236055 , n236051 , n236054 );
not ( n236056 , n236055 );
not ( n236057 , n236056 );
or ( n236058 , n235942 , n236057 );
not ( n236059 , n235941 );
and ( n236060 , n235995 , n236050 );
not ( n236061 , n235995 );
and ( n236062 , n236061 , n236053 );
nor ( n236063 , n236060 , n236062 );
nand ( n236064 , n236059 , n236063 );
nand ( n236065 , n236058 , n236064 );
not ( n236066 , n34378 );
not ( n236067 , n34374 );
or ( n236068 , n236066 , n236067 );
or ( n236069 , n34374 , n34378 );
nand ( n236070 , n236068 , n236069 );
xor ( n236071 , n28815 , n236070 );
xnor ( n236072 , n236071 , n224001 );
nand ( n236073 , n236072 , n231475 );
not ( n236074 , n236073 );
not ( n236075 , n50294 );
not ( n236076 , n236075 );
and ( n236077 , n236074 , n236076 );
and ( n236078 , n236073 , n236075 );
nor ( n236079 , n236077 , n236078 );
not ( n236080 , n236079 );
not ( n236081 , n39000 );
not ( n236082 , n204975 );
or ( n236083 , n236081 , n236082 );
or ( n236084 , n204975 , n39000 );
nand ( n236085 , n236083 , n236084 );
and ( n236086 , n28907 , n236085 );
not ( n236087 , n28907 );
not ( n236088 , n236085 );
and ( n236089 , n236087 , n236088 );
nor ( n236090 , n236086 , n236089 );
not ( n236091 , n236090 );
nand ( n236092 , n236091 , n53750 );
and ( n236093 , n236092 , n228139 );
not ( n236094 , n236092 );
and ( n236095 , n236094 , n50379 );
nor ( n236096 , n236093 , n236095 );
not ( n236097 , n236096 );
or ( n236098 , n236080 , n236097 );
or ( n236099 , n236096 , n236079 );
nand ( n236100 , n236098 , n236099 );
not ( n236101 , n46966 );
not ( n236102 , n25591 );
not ( n236103 , n231586 );
or ( n236104 , n236102 , n236103 );
or ( n236105 , n231586 , n25591 );
nand ( n236106 , n236104 , n236105 );
not ( n236107 , n236106 );
or ( n236108 , n236101 , n236107 );
or ( n236109 , n236106 , n222443 );
nand ( n236110 , n236108 , n236109 );
not ( n236111 , n236110 );
nand ( n236112 , n53733 , n236111 );
xnor ( n236113 , n236112 , n228099 );
not ( n236114 , n236113 );
and ( n236115 , n236100 , n236114 );
not ( n236116 , n236100 );
and ( n236117 , n236116 , n236113 );
nor ( n236118 , n236115 , n236117 );
not ( n236119 , n236118 );
not ( n236120 , n236119 );
not ( n236121 , n53774 );
buf ( n236122 , n220277 );
not ( n236123 , n236122 );
not ( n236124 , n45773 );
or ( n236125 , n236123 , n236124 );
or ( n236126 , n45773 , n236122 );
nand ( n236127 , n236125 , n236126 );
and ( n236128 , n236127 , n227330 );
not ( n236129 , n236127 );
and ( n236130 , n236129 , n42356 );
nor ( n236131 , n236128 , n236130 );
nand ( n236132 , n236121 , n236131 );
and ( n236133 , n236132 , n50437 );
not ( n236134 , n236132 );
and ( n236135 , n236134 , n50436 );
nor ( n236136 , n236133 , n236135 );
not ( n236137 , n236136 );
and ( n236138 , n33983 , n33980 );
not ( n236139 , n33983 );
buf ( n236140 , RI1749d878_968);
and ( n236141 , n236139 , n236140 );
nor ( n236142 , n236138 , n236141 );
not ( n236143 , n236142 );
not ( n236144 , n39212 );
or ( n236145 , n236143 , n236144 );
not ( n236146 , n236142 );
nand ( n236147 , n236146 , n39211 );
nand ( n236148 , n236145 , n236147 );
and ( n236149 , n236148 , n233008 );
not ( n236150 , n236148 );
and ( n236151 , n236150 , n39251 );
nor ( n236152 , n236149 , n236151 );
nand ( n236153 , n53795 , n236152 );
and ( n236154 , n236153 , n50427 );
not ( n236155 , n236153 );
and ( n236156 , n236155 , n50428 );
nor ( n236157 , n236154 , n236156 );
not ( n236158 , n236157 );
or ( n236159 , n236137 , n236158 );
or ( n236160 , n236157 , n236136 );
nand ( n236161 , n236159 , n236160 );
not ( n236162 , n236161 );
not ( n236163 , n236162 );
or ( n236164 , n236120 , n236163 );
nand ( n236165 , n236161 , n236118 );
nand ( n236166 , n236164 , n236165 );
not ( n236167 , n236166 );
not ( n236168 , n236167 );
and ( n236169 , n236065 , n236168 );
not ( n236170 , n236065 );
buf ( n236171 , n236166 );
not ( n236172 , n236171 );
and ( n236173 , n236170 , n236172 );
nor ( n236174 , n236169 , n236173 );
xor ( n236175 , n30372 , n205221 );
xnor ( n236176 , n236175 , n39532 );
not ( n236177 , n52194 );
nand ( n236178 , n236177 , n52207 );
nand ( n236179 , n236176 , n236178 );
not ( n236180 , n236179 );
nor ( n236181 , n236176 , n236178 );
nor ( n236182 , n236180 , n236181 );
not ( n236183 , n236182 );
not ( n236184 , n229906 );
nand ( n236185 , n52161 , n236184 );
and ( n236186 , n35365 , n207407 );
not ( n236187 , n35365 );
and ( n236188 , n236187 , n29647 );
or ( n236189 , n236186 , n236188 );
and ( n236190 , n236189 , n46671 );
not ( n236191 , n236189 );
and ( n236192 , n236191 , n46668 );
nor ( n236193 , n236190 , n236192 );
not ( n236194 , n236193 );
and ( n236195 , n236185 , n236194 );
not ( n236196 , n236185 );
and ( n236197 , n236196 , n236193 );
nor ( n236198 , n236195 , n236197 );
not ( n236199 , n236198 );
or ( n236200 , n236183 , n236199 );
not ( n236201 , n236182 );
not ( n236202 , n236198 );
nand ( n236203 , n236201 , n236202 );
nand ( n236204 , n236200 , n236203 );
not ( n236205 , n228145 );
and ( n236206 , n37314 , n41753 );
not ( n236207 , n37314 );
and ( n236208 , n236207 , n41754 );
or ( n236209 , n236206 , n236208 );
not ( n236210 , n236209 );
and ( n236211 , n236205 , n236210 );
and ( n236212 , n228145 , n236209 );
nor ( n236213 , n236211 , n236212 );
not ( n236214 , n236213 );
not ( n236215 , n236214 );
nand ( n236216 , n229861 , n52124 );
not ( n236217 , n236216 );
or ( n236218 , n236215 , n236217 );
or ( n236219 , n236216 , n236214 );
nand ( n236220 , n236218 , n236219 );
not ( n236221 , n236220 );
not ( n236222 , n229816 );
nand ( n236223 , n236222 , n52083 );
not ( n236224 , n236223 );
not ( n236225 , n26260 );
not ( n236226 , n36425 );
and ( n236227 , n236225 , n236226 );
and ( n236228 , n26260 , n36425 );
nor ( n236229 , n236227 , n236228 );
and ( n236230 , n236229 , n26310 );
not ( n236231 , n236229 );
and ( n236232 , n236231 , n26318 );
nor ( n236233 , n236230 , n236232 );
not ( n236234 , n236233 );
and ( n236235 , n236224 , n236234 );
not ( n236236 , n52084 );
nand ( n236237 , n236236 , n236222 );
and ( n236238 , n236237 , n236233 );
nor ( n236239 , n236235 , n236238 );
not ( n236240 , n236239 );
or ( n236241 , n236221 , n236240 );
or ( n236242 , n236239 , n236220 );
nand ( n236243 , n236241 , n236242 );
not ( n236244 , n43996 );
not ( n236245 , n32696 );
and ( n236246 , n236244 , n236245 );
and ( n236247 , n221761 , n32696 );
nor ( n236248 , n236246 , n236247 );
and ( n236249 , n236248 , n36377 );
not ( n236250 , n236248 );
and ( n236251 , n236250 , n44006 );
nor ( n236252 , n236249 , n236251 );
not ( n236253 , n236252 );
not ( n236254 , n236253 );
buf ( n236255 , n52039 );
nor ( n236256 , n229777 , n236255 );
not ( n236257 , n236256 );
and ( n236258 , n236254 , n236257 );
nor ( n236259 , n229777 , n236255 );
and ( n236260 , n236253 , n236259 );
nor ( n236261 , n236258 , n236260 );
and ( n236262 , n236243 , n236261 );
not ( n236263 , n236243 );
not ( n236264 , n236261 );
and ( n236265 , n236263 , n236264 );
nor ( n236266 , n236262 , n236265 );
xor ( n236267 , n236204 , n236266 );
not ( n236268 , n236267 );
buf ( n236269 , n51879 );
not ( n236270 , n236269 );
buf ( n236271 , n45464 );
not ( n236272 , n236271 );
not ( n236273 , n236272 );
nor ( n236274 , n39359 , n37387 );
not ( n236275 , n236274 );
nand ( n236276 , n37387 , n39359 );
nand ( n236277 , n236275 , n236276 );
not ( n236278 , n236277 );
or ( n236279 , n236273 , n236278 );
or ( n236280 , n236277 , n236272 );
nand ( n236281 , n236279 , n236280 );
not ( n236282 , n236281 );
not ( n236283 , n51940 );
nand ( n236284 , n51916 , n236283 );
not ( n236285 , n236284 );
or ( n236286 , n236282 , n236285 );
or ( n236287 , n236284 , n236281 );
nand ( n236288 , n236286 , n236287 );
not ( n236289 , n236288 );
not ( n236290 , n51984 );
not ( n236291 , n51962 );
nand ( n236292 , n236290 , n236291 );
not ( n236293 , n204505 );
not ( n236294 , n28029 );
not ( n236295 , n37580 );
or ( n236296 , n236294 , n236295 );
not ( n236297 , n28029 );
nand ( n236298 , n236297 , n37579 );
nand ( n236299 , n236296 , n236298 );
not ( n236300 , n236299 );
or ( n236301 , n236293 , n236300 );
not ( n236302 , n204508 );
or ( n236303 , n236299 , n236302 );
nand ( n236304 , n236301 , n236303 );
and ( n236305 , n236292 , n236304 );
not ( n236306 , n236292 );
not ( n236307 , n236304 );
and ( n236308 , n236306 , n236307 );
nor ( n236309 , n236305 , n236308 );
not ( n236310 , n236309 );
or ( n236311 , n236289 , n236310 );
or ( n236312 , n236288 , n236309 );
nand ( n236313 , n236311 , n236312 );
not ( n236314 , n236313 );
not ( n236315 , n51815 );
not ( n236316 , n229590 );
nand ( n236317 , n236315 , n236316 );
buf ( n236318 , n38078 );
not ( n236319 , n236318 );
not ( n236320 , n30033 );
not ( n236321 , n236320 );
or ( n236322 , n236319 , n236321 );
or ( n236323 , n236320 , n236318 );
nand ( n236324 , n236322 , n236323 );
not ( n236325 , n236324 );
not ( n236326 , n50453 );
and ( n236327 , n236325 , n236326 );
and ( n236328 , n236324 , n230718 );
nor ( n236329 , n236327 , n236328 );
and ( n236330 , n236317 , n236329 );
not ( n236331 , n236317 );
not ( n236332 , n236329 );
and ( n236333 , n236331 , n236332 );
nor ( n236334 , n236330 , n236333 );
not ( n236335 , n236334 );
not ( n236336 , n236335 );
not ( n236337 , n51875 );
not ( n236338 , n51858 );
nand ( n236339 , n236337 , n236338 );
not ( n236340 , n34362 );
not ( n236341 , n41668 );
or ( n236342 , n236340 , n236341 );
or ( n236343 , n37020 , n34362 );
nand ( n236344 , n236342 , n236343 );
and ( n236345 , n236344 , n223530 );
not ( n236346 , n236344 );
and ( n236347 , n236346 , n45773 );
nor ( n236348 , n236345 , n236347 );
not ( n236349 , n236348 );
and ( n236350 , n236339 , n236349 );
not ( n236351 , n236339 );
and ( n236352 , n236351 , n236348 );
nor ( n236353 , n236350 , n236352 );
not ( n236354 , n236353 );
not ( n236355 , n236354 );
or ( n236356 , n236336 , n236355 );
nand ( n236357 , n236353 , n236334 );
nand ( n236358 , n236356 , n236357 );
nand ( n236359 , n51795 , n51895 );
not ( n236360 , n236359 );
buf ( n236361 , n28370 );
not ( n236362 , n236361 );
not ( n236363 , n36349 );
or ( n236364 , n236362 , n236363 );
or ( n236365 , n225836 , n236361 );
nand ( n236366 , n236364 , n236365 );
not ( n236367 , n236366 );
not ( n236368 , n40345 );
and ( n236369 , n236367 , n236368 );
and ( n236370 , n236366 , n55686 );
nor ( n236371 , n236369 , n236370 );
not ( n236372 , n236371 );
not ( n236373 , n236372 );
and ( n236374 , n236360 , n236373 );
and ( n236375 , n236359 , n236372 );
nor ( n236376 , n236374 , n236375 );
and ( n236377 , n236358 , n236376 );
not ( n236378 , n236358 );
not ( n236379 , n236376 );
and ( n236380 , n236378 , n236379 );
nor ( n236381 , n236377 , n236380 );
not ( n236382 , n236381 );
or ( n236383 , n236314 , n236382 );
or ( n236384 , n236381 , n236313 );
nand ( n236385 , n236383 , n236384 );
not ( n236386 , n236385 );
or ( n236387 , n236270 , n236386 );
or ( n236388 , n236385 , n236269 );
nand ( n236389 , n236387 , n236388 );
not ( n236390 , n236389 );
and ( n236391 , n236268 , n236390 );
buf ( n236392 , n236267 );
and ( n236393 , n236392 , n236389 );
nor ( n236394 , n236391 , n236393 );
nand ( n236395 , n236174 , n236394 );
not ( n236396 , n50969 );
not ( n236397 , n235602 );
nand ( n236398 , n236397 , n51026 );
not ( n236399 , n236398 );
or ( n236400 , n236396 , n236399 );
or ( n236401 , n236398 , n50969 );
nand ( n236402 , n236400 , n236401 );
not ( n236403 , n236402 );
not ( n236404 , n236403 );
not ( n236405 , n235728 );
or ( n236406 , n236404 , n236405 );
not ( n236407 , n236403 );
nand ( n236408 , n236407 , n235718 );
nand ( n236409 , n236406 , n236408 );
not ( n236410 , n236409 );
not ( n236411 , n32447 );
not ( n236412 , n236411 );
not ( n236413 , n32459 );
not ( n236414 , n31156 );
not ( n236415 , n42285 );
or ( n236416 , n236414 , n236415 );
or ( n236417 , n42285 , n31156 );
nand ( n236418 , n236416 , n236417 );
and ( n236419 , n236418 , n45382 );
not ( n236420 , n236418 );
and ( n236421 , n236420 , n29991 );
nor ( n236422 , n236419 , n236421 );
nand ( n236423 , n236413 , n236422 );
not ( n236424 , n236423 );
or ( n236425 , n236412 , n236424 );
or ( n236426 , n236423 , n236411 );
nand ( n236427 , n236425 , n236426 );
not ( n236428 , n236427 );
not ( n236429 , n29314 );
not ( n236430 , n205426 );
or ( n236431 , n236429 , n236430 );
or ( n236432 , n205421 , n29314 );
nand ( n236433 , n236431 , n236432 );
and ( n236434 , n236433 , n205436 );
not ( n236435 , n236433 );
and ( n236436 , n236435 , n205435 );
nor ( n236437 , n236434 , n236436 );
not ( n236438 , n236437 );
nand ( n236439 , n236438 , n32328 );
not ( n236440 , n236439 );
not ( n236441 , n229004 );
and ( n236442 , n236440 , n236441 );
and ( n236443 , n236439 , n229004 );
nor ( n236444 , n236442 , n236443 );
not ( n236445 , n236444 );
or ( n236446 , n236428 , n236445 );
or ( n236447 , n236444 , n236427 );
nand ( n236448 , n236446 , n236447 );
not ( n236449 , n236448 );
not ( n236450 , n236449 );
not ( n236451 , n227097 );
not ( n236452 , n40230 );
or ( n236453 , n236451 , n236452 );
not ( n236454 , n227097 );
nand ( n236455 , n236454 , n30533 );
nand ( n236456 , n236453 , n236455 );
and ( n236457 , n236456 , n30496 );
not ( n236458 , n236456 );
not ( n236459 , n208303 );
and ( n236460 , n236458 , n236459 );
nor ( n236461 , n236457 , n236460 );
nand ( n236462 , n31788 , n236461 );
not ( n236463 , n236462 );
not ( n236464 , n51170 );
and ( n236465 , n236463 , n236464 );
and ( n236466 , n236462 , n51170 );
nor ( n236467 , n236465 , n236466 );
not ( n236468 , n236467 );
not ( n236469 , n236468 );
not ( n236470 , n32989 );
not ( n236471 , n28697 );
not ( n236472 , n40733 );
not ( n236473 , n236472 );
or ( n236474 , n236471 , n236473 );
not ( n236475 , n28697 );
nand ( n236476 , n236475 , n40733 );
nand ( n236477 , n236474 , n236476 );
not ( n236478 , n236477 );
or ( n236479 , n236470 , n236478 );
or ( n236480 , n236477 , n32989 );
nand ( n236481 , n236479 , n236480 );
nand ( n236482 , n32013 , n236481 );
not ( n236483 , n236482 );
not ( n236484 , n31947 );
or ( n236485 , n236483 , n236484 );
or ( n236486 , n31947 , n236482 );
nand ( n236487 , n236485 , n236486 );
not ( n236488 , n236487 );
not ( n236489 , n236488 );
or ( n236490 , n236469 , n236489 );
nand ( n236491 , n236487 , n236467 );
nand ( n236492 , n236490 , n236491 );
and ( n236493 , n236492 , n31748 );
not ( n236494 , n236492 );
not ( n236495 , n31748 );
and ( n236496 , n236494 , n236495 );
nor ( n236497 , n236493 , n236496 );
not ( n236498 , n236497 );
not ( n236499 , n236498 );
or ( n236500 , n236450 , n236499 );
nand ( n236501 , n236497 , n236448 );
nand ( n236502 , n236500 , n236501 );
not ( n236503 , n236502 );
buf ( n236504 , n236503 );
not ( n236505 , n236504 );
and ( n236506 , n236410 , n236505 );
and ( n236507 , n236409 , n236504 );
nor ( n236508 , n236506 , n236507 );
not ( n236509 , n236508 );
and ( n236510 , n236395 , n236509 );
not ( n236511 , n236395 );
and ( n236512 , n236511 , n236508 );
nor ( n236513 , n236510 , n236512 );
or ( n236514 , n236513 , n226003 );
nand ( n236515 , n235912 , n236514 );
buf ( n236516 , n236515 );
not ( n236517 , n236338 );
not ( n236518 , n37618 );
not ( n236519 , n31126 );
or ( n236520 , n236518 , n236519 );
or ( n236521 , n31126 , n37618 );
nand ( n236522 , n236520 , n236521 );
and ( n236523 , n236522 , n31136 );
not ( n236524 , n236522 );
and ( n236525 , n236524 , n29694 );
nor ( n236526 , n236523 , n236525 );
not ( n236527 , n236526 );
not ( n236528 , n51855 );
nand ( n236529 , n236527 , n236528 );
not ( n236530 , n236529 );
or ( n236531 , n236517 , n236530 );
or ( n236532 , n236529 , n236338 );
nand ( n236533 , n236531 , n236532 );
buf ( n236534 , n236533 );
not ( n236535 , n236534 );
not ( n236536 , n51998 );
or ( n236537 , n236535 , n236536 );
or ( n236538 , n51998 , n236534 );
nand ( n236539 , n236537 , n236538 );
xor ( n236540 , n229991 , n236539 );
not ( n236541 , n236540 );
not ( n236542 , n236541 );
not ( n236543 , n43250 );
not ( n236544 , n236543 );
not ( n236545 , n46810 );
or ( n236546 , n236544 , n236545 );
nand ( n236547 , n45518 , n43250 );
nand ( n236548 , n236546 , n236547 );
not ( n236549 , n236548 );
not ( n236550 , n46815 );
and ( n236551 , n236549 , n236550 );
and ( n236552 , n236548 , n46815 );
nor ( n236553 , n236551 , n236552 );
buf ( n236554 , n45212 );
not ( n236555 , n236554 );
not ( n236556 , n28344 );
or ( n236557 , n236555 , n236556 );
or ( n236558 , n222628 , n236554 );
nand ( n236559 , n236557 , n236558 );
xor ( n236560 , n236559 , n39671 );
not ( n236561 , n236560 );
nand ( n236562 , n236553 , n236561 );
not ( n236563 , n236562 );
not ( n236564 , n43464 );
or ( n236565 , n236563 , n236564 );
or ( n236566 , n43464 , n236562 );
nand ( n236567 , n236565 , n236566 );
not ( n236568 , n236567 );
not ( n236569 , n221107 );
buf ( n236570 , n27847 );
not ( n236571 , n236570 );
not ( n236572 , n33755 );
or ( n236573 , n236571 , n236572 );
or ( n236574 , n33759 , n236570 );
nand ( n236575 , n236573 , n236574 );
xor ( n236576 , n31253 , n236575 );
nand ( n236577 , n236569 , n236576 );
not ( n236578 , n236577 );
not ( n236579 , n221116 );
not ( n236580 , n236579 );
and ( n236581 , n236578 , n236580 );
and ( n236582 , n236577 , n236579 );
nor ( n236583 , n236581 , n236582 );
not ( n236584 , n236583 );
not ( n236585 , n221062 );
or ( n236586 , n236584 , n236585 );
or ( n236587 , n221062 , n236583 );
nand ( n236588 , n236586 , n236587 );
not ( n236589 , n43304 );
not ( n236590 , n236589 );
buf ( n236591 , n30887 );
not ( n236592 , n236591 );
not ( n236593 , n236592 );
not ( n236594 , n36457 );
or ( n236595 , n236593 , n236594 );
nand ( n236596 , n45370 , n236591 );
nand ( n236597 , n236595 , n236596 );
and ( n236598 , n236597 , n39211 );
not ( n236599 , n236597 );
and ( n236600 , n236599 , n39212 );
or ( n236601 , n236598 , n236600 );
not ( n236602 , n236601 );
nand ( n236603 , n236602 , n43314 );
not ( n236604 , n236603 );
and ( n236605 , n236590 , n236604 );
and ( n236606 , n236589 , n236603 );
nor ( n236607 , n236605 , n236606 );
and ( n236608 , n236588 , n236607 );
not ( n236609 , n236588 );
not ( n236610 , n236607 );
and ( n236611 , n236609 , n236610 );
nor ( n236612 , n236608 , n236611 );
not ( n236613 , n236553 );
nand ( n236614 , n236613 , n43463 );
not ( n236615 , n236614 );
not ( n236616 , n43457 );
and ( n236617 , n236615 , n236616 );
not ( n236618 , n236553 );
nand ( n236619 , n43463 , n236618 );
and ( n236620 , n236619 , n43457 );
nor ( n236621 , n236617 , n236620 );
not ( n236622 , n236621 );
not ( n236623 , n56064 );
and ( n236624 , n236622 , n236623 );
and ( n236625 , n236621 , n56064 );
nor ( n236626 , n236624 , n236625 );
not ( n236627 , n236626 );
and ( n236628 , n236612 , n236627 );
not ( n236629 , n236612 );
and ( n236630 , n236629 , n236626 );
nor ( n236631 , n236628 , n236630 );
not ( n236632 , n236631 );
or ( n236633 , n236568 , n236632 );
and ( n236634 , n236612 , n236626 );
not ( n236635 , n236612 );
and ( n236636 , n236635 , n236627 );
nor ( n236637 , n236634 , n236636 );
not ( n236638 , n236567 );
nand ( n236639 , n236637 , n236638 );
nand ( n236640 , n236633 , n236639 );
not ( n236641 , n236640 );
not ( n236642 , n43051 );
not ( n236643 , n28247 );
not ( n236644 , n205042 );
not ( n236645 , n32064 );
or ( n236646 , n236644 , n236645 );
or ( n236647 , n32064 , n205042 );
nand ( n236648 , n236646 , n236647 );
not ( n236649 , n236648 );
not ( n236650 , n32077 );
not ( n236651 , n236650 );
or ( n236652 , n236649 , n236651 );
or ( n236653 , n236650 , n236648 );
nand ( n236654 , n236652 , n236653 );
not ( n236655 , n236654 );
and ( n236656 , n236643 , n236655 );
and ( n236657 , n236654 , n28247 );
nor ( n236658 , n236656 , n236657 );
not ( n236659 , n236658 );
nand ( n236660 , n236642 , n236659 );
not ( n236661 , n236660 );
not ( n236662 , n43037 );
not ( n236663 , n236662 );
and ( n236664 , n236661 , n236663 );
and ( n236665 , n236660 , n236662 );
nor ( n236666 , n236664 , n236665 );
not ( n236667 , n236666 );
not ( n236668 , n236667 );
not ( n236669 , n43072 );
not ( n236670 , n236669 );
not ( n236671 , n34736 );
and ( n236672 , n31099 , n34177 );
not ( n236673 , n31099 );
and ( n236674 , n236673 , n218085 );
nor ( n236675 , n236672 , n236674 );
not ( n236676 , n236675 );
not ( n236677 , n236676 );
or ( n236678 , n236671 , n236677 );
nand ( n236679 , n236675 , n34735 );
nand ( n236680 , n236678 , n236679 );
not ( n236681 , n43086 );
nand ( n236682 , n236680 , n236681 );
not ( n236683 , n236682 );
or ( n236684 , n236670 , n236683 );
or ( n236685 , n236682 , n236669 );
nand ( n236686 , n236684 , n236685 );
not ( n236687 , n236686 );
not ( n236688 , n236687 );
or ( n236689 , n236668 , n236688 );
nand ( n236690 , n236686 , n236666 );
nand ( n236691 , n236689 , n236690 );
not ( n236692 , n43119 );
not ( n236693 , n44128 );
not ( n236694 , n33096 );
or ( n236695 , n236693 , n236694 );
or ( n236696 , n33096 , n44128 );
nand ( n236697 , n236695 , n236696 );
and ( n236698 , n236697 , n33142 );
not ( n236699 , n236697 );
and ( n236700 , n236699 , n33135 );
nor ( n236701 , n236698 , n236700 );
nand ( n236702 , n236692 , n236701 );
and ( n236703 , n236702 , n220890 );
not ( n236704 , n236702 );
not ( n236705 , n220890 );
and ( n236706 , n236704 , n236705 );
nor ( n236707 , n236703 , n236706 );
not ( n236708 , n236707 );
and ( n236709 , n236691 , n236708 );
not ( n236710 , n236691 );
and ( n236711 , n236710 , n236707 );
nor ( n236712 , n236709 , n236711 );
not ( n236713 , n236712 );
not ( n236714 , n236713 );
not ( n236715 , n43162 );
not ( n236716 , n32855 );
not ( n236717 , n35861 );
or ( n236718 , n236716 , n236717 );
nand ( n236719 , n55480 , n32851 );
nand ( n236720 , n236718 , n236719 );
not ( n236721 , n236720 );
not ( n236722 , n37533 );
and ( n236723 , n236721 , n236722 );
and ( n236724 , n236720 , n37533 );
nor ( n236725 , n236723 , n236724 );
not ( n236726 , n236725 );
nand ( n236727 , n236715 , n236726 );
not ( n236728 , n236727 );
not ( n236729 , n43159 );
and ( n236730 , n236728 , n236729 );
and ( n236731 , n236727 , n43159 );
nor ( n236732 , n236730 , n236731 );
not ( n236733 , n43187 );
not ( n236734 , n41448 );
not ( n236735 , n236734 );
not ( n236736 , n236735 );
not ( n236737 , n230227 );
not ( n236738 , n30506 );
and ( n236739 , n236737 , n236738 );
and ( n236740 , n230227 , n30506 );
nor ( n236741 , n236739 , n236740 );
not ( n236742 , n236741 );
and ( n236743 , n236736 , n236742 );
and ( n236744 , n236735 , n236741 );
nor ( n236745 , n236743 , n236744 );
not ( n236746 , n236745 );
nand ( n236747 , n236733 , n236746 );
and ( n236748 , n236747 , n43199 );
not ( n236749 , n236747 );
not ( n236750 , n43199 );
and ( n236751 , n236749 , n236750 );
nor ( n236752 , n236748 , n236751 );
and ( n236753 , n236732 , n236752 );
not ( n236754 , n236732 );
not ( n236755 , n236752 );
and ( n236756 , n236754 , n236755 );
nor ( n236757 , n236753 , n236756 );
not ( n236758 , n236757 );
or ( n236759 , n236714 , n236758 );
not ( n236760 , n236757 );
nand ( n236761 , n236760 , n236712 );
nand ( n236762 , n236759 , n236761 );
not ( n236763 , n236762 );
not ( n236764 , n236763 );
and ( n236765 , n236641 , n236764 );
not ( n236766 , n236762 );
and ( n236767 , n236640 , n236766 );
nor ( n236768 , n236765 , n236767 );
not ( n236769 , n236768 );
not ( n236770 , n236769 );
or ( n236771 , n236542 , n236770 );
not ( n236772 , n226304 );
nand ( n236773 , n236772 , n48533 );
and ( n236774 , n236773 , n47563 );
not ( n236775 , n236773 );
not ( n236776 , n47563 );
and ( n236777 , n236775 , n236776 );
nor ( n236778 , n236774 , n236777 );
not ( n236779 , n236778 );
not ( n236780 , n236779 );
buf ( n236781 , n234880 );
not ( n236782 , n236781 );
or ( n236783 , n236780 , n236782 );
not ( n236784 , n236779 );
nand ( n236785 , n236784 , n234881 );
nand ( n236786 , n236783 , n236785 );
and ( n236787 , n236786 , n234889 );
not ( n236788 , n236786 );
buf ( n236789 , n48676 );
and ( n236790 , n236788 , n236789 );
nor ( n236791 , n236787 , n236790 );
not ( n236792 , n236791 );
nor ( n236793 , n236792 , n235050 );
nand ( n236794 , n236771 , n236793 );
buf ( n236795 , n31571 );
nor ( n236796 , n236540 , n236795 );
nand ( n236797 , n236796 , n236792 , n236769 );
buf ( n236798 , n35431 );
nand ( n236799 , n236798 , n36602 );
nand ( n236800 , n236794 , n236797 , n236799 );
buf ( n236801 , n236800 );
not ( n236802 , RI19a93fe0_2654);
or ( n236803 , n25328 , n236802 );
not ( n236804 , RI19a8a080_2724);
or ( n236805 , n25335 , n236804 );
nand ( n236806 , n236803 , n236805 );
buf ( n236807 , n236806 );
nor ( n236808 , n53556 , n234608 );
not ( n236809 , n236808 );
not ( n236810 , n53558 );
not ( n236811 , n236810 );
not ( n236812 , n236811 );
and ( n236813 , n236809 , n236812 );
and ( n236814 , n236808 , n236811 );
nor ( n236815 , n236813 , n236814 );
not ( n236816 , n236815 );
not ( n236817 , n231421 );
or ( n236818 , n236816 , n236817 );
or ( n236819 , n231421 , n236815 );
nand ( n236820 , n236818 , n236819 );
buf ( n236821 , n34439 );
and ( n236822 , n236820 , n236821 );
not ( n236823 , n236820 );
and ( n236824 , n236823 , n53665 );
nor ( n236825 , n236822 , n236824 );
nand ( n236826 , n236825 , n33255 );
not ( n236827 , n35795 );
nand ( n236828 , n35706 , n35729 );
not ( n236829 , n236828 );
not ( n236830 , n204897 );
or ( n236831 , n236829 , n236830 );
or ( n236832 , n204897 , n236828 );
nand ( n236833 , n236831 , n236832 );
not ( n236834 , n236833 );
nand ( n236835 , n35788 , n35748 );
not ( n236836 , n236835 );
not ( n236837 , n204635 );
and ( n236838 , n236836 , n236837 );
and ( n236839 , n236835 , n204635 );
nor ( n236840 , n236838 , n236839 );
not ( n236841 , n236840 );
or ( n236842 , n236834 , n236841 );
or ( n236843 , n236840 , n236833 );
nand ( n236844 , n236842 , n236843 );
not ( n236845 , n236844 );
nand ( n236846 , n35626 , n35646 );
not ( n236847 , n236846 );
not ( n236848 , n205076 );
not ( n236849 , n236848 );
and ( n236850 , n236847 , n236849 );
and ( n236851 , n236846 , n236848 );
nor ( n236852 , n236850 , n236851 );
not ( n236853 , n236852 );
not ( n236854 , n236853 );
nand ( n236855 , n35599 , n35529 );
not ( n236856 , n236855 );
not ( n236857 , n205246 );
or ( n236858 , n236856 , n236857 );
or ( n236859 , n205246 , n236855 );
nand ( n236860 , n236858 , n236859 );
not ( n236861 , n236860 );
not ( n236862 , n236861 );
or ( n236863 , n236854 , n236862 );
nand ( n236864 , n236860 , n236852 );
nand ( n236865 , n236863 , n236864 );
nand ( n236866 , n35466 , n50505 );
and ( n236867 , n236866 , n27766 );
not ( n236868 , n236866 );
and ( n236869 , n236868 , n27765 );
nor ( n236870 , n236867 , n236869 );
and ( n236871 , n236865 , n236870 );
not ( n236872 , n236865 );
not ( n236873 , n236870 );
and ( n236874 , n236872 , n236873 );
nor ( n236875 , n236871 , n236874 );
not ( n236876 , n236875 );
or ( n236877 , n236845 , n236876 );
not ( n236878 , n236844 );
not ( n236879 , n236875 );
nand ( n236880 , n236878 , n236879 );
nand ( n236881 , n236877 , n236880 );
not ( n236882 , n236881 );
not ( n236883 , n236882 );
not ( n236884 , n236883 );
or ( n236885 , n236827 , n236884 );
buf ( n236886 , n236881 );
or ( n236887 , n236886 , n35795 );
nand ( n236888 , n236885 , n236887 );
not ( n236889 , n236888 );
not ( n236890 , n231585 );
not ( n236891 , n236890 );
not ( n236892 , n205281 );
or ( n236893 , n236891 , n236892 );
or ( n236894 , n35199 , n236890 );
nand ( n236895 , n236893 , n236894 );
and ( n236896 , n236895 , n205322 );
not ( n236897 , n236895 );
and ( n236898 , n236897 , n205325 );
nor ( n236899 , n236896 , n236898 );
not ( n236900 , n236899 );
not ( n236901 , n236900 );
nand ( n236902 , n55531 , n234905 );
not ( n236903 , n236902 );
or ( n236904 , n236901 , n236903 );
or ( n236905 , n236902 , n236900 );
nand ( n236906 , n236904 , n236905 );
not ( n236907 , n236906 );
nand ( n236908 , n234928 , n233360 );
not ( n236909 , n236908 );
not ( n236910 , n31337 );
not ( n236911 , n35821 );
or ( n236912 , n236910 , n236911 );
not ( n236913 , n31337 );
nand ( n236914 , n236913 , n31613 );
nand ( n236915 , n236912 , n236914 );
and ( n236916 , n236915 , n35861 );
not ( n236917 , n236915 );
and ( n236918 , n236917 , n222753 );
nor ( n236919 , n236916 , n236918 );
not ( n236920 , n236919 );
not ( n236921 , n236920 );
and ( n236922 , n236909 , n236921 );
nand ( n236923 , n233360 , n234928 );
and ( n236924 , n236923 , n236920 );
nor ( n236925 , n236922 , n236924 );
not ( n236926 , n236925 );
or ( n236927 , n236907 , n236926 );
or ( n236928 , n236925 , n236906 );
nand ( n236929 , n236927 , n236928 );
not ( n236930 , n234954 );
nand ( n236931 , n236930 , n55634 );
not ( n236932 , n236931 );
buf ( n236933 , n34719 );
not ( n236934 , n236933 );
not ( n236935 , n204859 );
or ( n236936 , n236934 , n236935 );
or ( n236937 , n204859 , n236933 );
nand ( n236938 , n236936 , n236937 );
and ( n236939 , n236938 , n46894 );
not ( n236940 , n236938 );
and ( n236941 , n236940 , n204895 );
nor ( n236942 , n236939 , n236941 );
not ( n236943 , n236942 );
not ( n236944 , n236943 );
and ( n236945 , n236932 , n236944 );
not ( n236946 , n234954 );
nand ( n236947 , n236946 , n55634 );
and ( n236948 , n236947 , n236943 );
nor ( n236949 , n236945 , n236948 );
not ( n236950 , n236949 );
and ( n236951 , n236929 , n236950 );
not ( n236952 , n236929 );
and ( n236953 , n236952 , n236949 );
nor ( n236954 , n236951 , n236953 );
not ( n236955 , n236954 );
not ( n236956 , n234995 );
nand ( n236957 , n236956 , n55710 );
buf ( n236958 , n35087 );
and ( n236959 , n236958 , n39874 );
not ( n236960 , n236958 );
and ( n236961 , n236960 , n46633 );
or ( n236962 , n236959 , n236961 );
and ( n236963 , n236962 , n204672 );
not ( n236964 , n236962 );
and ( n236965 , n236964 , n46639 );
nor ( n236966 , n236963 , n236965 );
not ( n236967 , n236966 );
and ( n236968 , n236957 , n236967 );
not ( n236969 , n236957 );
and ( n236970 , n236969 , n236966 );
nor ( n236971 , n236968 , n236970 );
not ( n236972 , n236971 );
not ( n236973 , n236972 );
nand ( n236974 , n234979 , n55677 );
not ( n236975 , n236974 );
xor ( n236976 , n39967 , n28647 );
xnor ( n236977 , n236976 , n28665 );
not ( n236978 , n236977 );
not ( n236979 , n236978 );
or ( n236980 , n236975 , n236979 );
or ( n236981 , n236978 , n236974 );
nand ( n236982 , n236980 , n236981 );
not ( n236983 , n236982 );
not ( n236984 , n236983 );
or ( n236985 , n236973 , n236984 );
nand ( n236986 , n236982 , n236971 );
nand ( n236987 , n236985 , n236986 );
not ( n236988 , n236987 );
and ( n236989 , n236955 , n236988 );
not ( n236990 , n236955 );
and ( n236991 , n236990 , n236987 );
nor ( n236992 , n236989 , n236991 );
buf ( n236993 , n236992 );
not ( n236994 , n236993 );
not ( n236995 , n236994 );
and ( n236996 , n236889 , n236995 );
not ( n236997 , n236993 );
and ( n236998 , n236888 , n236997 );
nor ( n236999 , n236996 , n236998 );
not ( n237000 , n236999 );
not ( n237001 , n45619 );
not ( n237002 , n28743 );
and ( n237003 , n237001 , n237002 );
and ( n237004 , n45619 , n28743 );
nor ( n237005 , n237003 , n237004 );
not ( n237006 , n237005 );
not ( n237007 , n34381 );
or ( n237008 , n237006 , n237007 );
or ( n237009 , n34381 , n237005 );
nand ( n237010 , n237008 , n237009 );
buf ( n237011 , n237010 );
not ( n237012 , n237011 );
not ( n237013 , n231159 );
not ( n237014 , n53385 );
nand ( n237015 , n237013 , n237014 );
not ( n237016 , n237015 );
or ( n237017 , n237012 , n237016 );
not ( n237018 , n231159 );
nand ( n237019 , n237018 , n237014 );
or ( n237020 , n237019 , n237011 );
nand ( n237021 , n237017 , n237020 );
not ( n237022 , n237021 );
xor ( n237023 , n27683 , n222033 );
xnor ( n237024 , n237023 , n231687 );
nand ( n237025 , n237024 , n53434 );
not ( n237026 , n237025 );
xor ( n237027 , n31957 , n31227 );
xnor ( n237028 , n237027 , n29088 );
not ( n237029 , n237028 );
not ( n237030 , n237029 );
and ( n237031 , n237026 , n237030 );
and ( n237032 , n237025 , n237029 );
nor ( n237033 , n237031 , n237032 );
not ( n237034 , n237010 );
nand ( n237035 , n237034 , n231159 );
not ( n237036 , n31881 );
not ( n237037 , n35960 );
or ( n237038 , n237036 , n237037 );
or ( n237039 , n35960 , n31881 );
nand ( n237040 , n237038 , n237039 );
and ( n237041 , n237040 , n30756 );
not ( n237042 , n237040 );
and ( n237043 , n237042 , n30771 );
nor ( n237044 , n237041 , n237043 );
not ( n237045 , n237044 );
not ( n237046 , n237045 );
xnor ( n237047 , n237035 , n237046 );
not ( n237048 , n237047 );
not ( n237049 , n39480 );
buf ( n237050 , RI173d4d88_1718);
not ( n237051 , n237050 );
and ( n237052 , n237049 , n237051 );
and ( n237053 , n39480 , n237050 );
nor ( n237054 , n237052 , n237053 );
and ( n237055 , n237054 , n43554 );
not ( n237056 , n237054 );
and ( n237057 , n237056 , n43803 );
nor ( n237058 , n237055 , n237057 );
not ( n237059 , n237058 );
nand ( n237060 , n237059 , n231097 );
not ( n237061 , n33630 );
not ( n237062 , n52094 );
or ( n237063 , n237061 , n237062 );
not ( n237064 , n33630 );
nand ( n237065 , n237064 , n204257 );
nand ( n237066 , n237063 , n237065 );
xor ( n237067 , n237066 , n32136 );
and ( n237068 , n237060 , n237067 );
not ( n237069 , n237060 );
not ( n237070 , n237067 );
and ( n237071 , n237069 , n237070 );
nor ( n237072 , n237068 , n237071 );
not ( n237073 , n237072 );
or ( n237074 , n237048 , n237073 );
not ( n237075 , n237047 );
not ( n237076 , n237072 );
nand ( n237077 , n237075 , n237076 );
nand ( n237078 , n237074 , n237077 );
xor ( n237079 , n237033 , n237078 );
not ( n237080 , n36177 );
not ( n237081 , n38356 );
or ( n237082 , n237080 , n237081 );
not ( n237083 , n38353 );
nand ( n237084 , n237083 , n36173 );
nand ( n237085 , n237082 , n237084 );
and ( n237086 , n237085 , n28557 );
not ( n237087 , n237085 );
and ( n237088 , n237087 , n225104 );
nor ( n237089 , n237086 , n237088 );
nand ( n237090 , n53268 , n237089 );
not ( n237091 , n34490 );
not ( n237092 , n43636 );
or ( n237093 , n237091 , n237092 );
or ( n237094 , n43635 , n34490 );
nand ( n237095 , n237093 , n237094 );
and ( n237096 , n237095 , n47330 );
not ( n237097 , n237095 );
and ( n237098 , n237097 , n225090 );
nor ( n237099 , n237096 , n237098 );
and ( n237100 , n237090 , n237099 );
not ( n237101 , n237090 );
not ( n237102 , n237099 );
and ( n237103 , n237101 , n237102 );
nor ( n237104 , n237100 , n237103 );
not ( n237105 , n237104 );
not ( n237106 , n33334 );
not ( n237107 , n30580 );
or ( n237108 , n237106 , n237107 );
nand ( n237109 , n39555 , n33330 );
nand ( n237110 , n237108 , n237109 );
and ( n237111 , n237110 , n39558 );
not ( n237112 , n237110 );
and ( n237113 , n237112 , n39559 );
nor ( n237114 , n237111 , n237113 );
nand ( n237115 , n53324 , n237114 );
not ( n237116 , n237115 );
not ( n237117 , n207340 );
not ( n237118 , n229281 );
or ( n237119 , n237117 , n237118 );
nand ( n237120 , n38912 , n29575 );
nand ( n237121 , n237119 , n237120 );
and ( n237122 , n237121 , n225218 );
not ( n237123 , n237121 );
and ( n237124 , n237123 , n225217 );
nor ( n237125 , n237122 , n237124 );
not ( n237126 , n237125 );
not ( n237127 , n237126 );
and ( n237128 , n237116 , n237127 );
and ( n237129 , n237115 , n237126 );
nor ( n237130 , n237128 , n237129 );
not ( n237131 , n237130 );
and ( n237132 , n237105 , n237131 );
and ( n237133 , n237104 , n237130 );
nor ( n237134 , n237132 , n237133 );
xnor ( n237135 , n237079 , n237134 );
not ( n237136 , n237135 );
or ( n237137 , n237022 , n237136 );
not ( n237138 , n237021 );
not ( n237139 , n237033 );
and ( n237140 , n237078 , n237139 );
not ( n237141 , n237078 );
and ( n237142 , n237141 , n237033 );
nor ( n237143 , n237140 , n237142 );
not ( n237144 , n237134 );
and ( n237145 , n237143 , n237144 );
not ( n237146 , n237143 );
and ( n237147 , n237146 , n237134 );
nor ( n237148 , n237145 , n237147 );
nand ( n237149 , n237138 , n237148 );
nand ( n237150 , n237137 , n237149 );
buf ( n237151 , n26036 );
not ( n237152 , n237151 );
not ( n237153 , n29174 );
or ( n237154 , n237152 , n237153 );
not ( n237155 , n237151 );
nand ( n237156 , n237155 , n29161 );
nand ( n237157 , n237154 , n237156 );
not ( n237158 , n237157 );
not ( n237159 , n33936 );
and ( n237160 , n237158 , n237159 );
and ( n237161 , n237157 , n33936 );
nor ( n237162 , n237160 , n237161 );
not ( n237163 , n42022 );
not ( n237164 , n237163 );
not ( n237165 , n45214 );
or ( n237166 , n237164 , n237165 );
or ( n237167 , n45214 , n237163 );
nand ( n237168 , n237166 , n237167 );
and ( n237169 , n237168 , n34416 );
not ( n237170 , n237168 );
and ( n237171 , n237170 , n204586 );
nor ( n237172 , n237169 , n237171 );
nand ( n237173 , n237162 , n237172 );
not ( n237174 , n237173 );
not ( n237175 , n33657 );
not ( n237176 , n40503 );
and ( n237177 , n237175 , n237176 );
and ( n237178 , n33657 , n40503 );
nor ( n237179 , n237177 , n237178 );
and ( n237180 , n237179 , n34227 );
not ( n237181 , n237179 );
and ( n237182 , n237181 , n34218 );
nor ( n237183 , n237180 , n237182 );
not ( n237184 , n237183 );
and ( n237185 , n237174 , n237184 );
and ( n237186 , n237173 , n237183 );
nor ( n237187 , n237185 , n237186 );
not ( n237188 , n237187 );
not ( n237189 , n237188 );
not ( n237190 , n31712 );
not ( n237191 , n53706 );
or ( n237192 , n237190 , n237191 );
or ( n237193 , n43096 , n31712 );
nand ( n237194 , n237192 , n237193 );
and ( n237195 , n237194 , n35584 );
not ( n237196 , n237194 );
and ( n237197 , n237196 , n35590 );
nor ( n237198 , n237195 , n237197 );
not ( n237199 , n36147 );
not ( n237200 , n237199 );
not ( n237201 , n225459 );
or ( n237202 , n237200 , n237201 );
or ( n237203 , n225459 , n237199 );
nand ( n237204 , n237202 , n237203 );
and ( n237205 , n237204 , n237083 );
not ( n237206 , n237204 );
and ( n237207 , n237206 , n38356 );
nor ( n237208 , n237205 , n237207 );
nand ( n237209 , n237198 , n237208 );
not ( n237210 , n237209 );
xor ( n237211 , n25526 , n46258 );
xnor ( n237212 , n237211 , n33886 );
not ( n237213 , n237212 );
or ( n237214 , n237210 , n237213 );
or ( n237215 , n237212 , n237209 );
nand ( n237216 , n237214 , n237215 );
not ( n237217 , n237216 );
not ( n237218 , n237217 );
or ( n237219 , n237189 , n237218 );
nand ( n237220 , n237216 , n237187 );
nand ( n237221 , n237219 , n237220 );
and ( n237222 , n33838 , n37193 );
not ( n237223 , n33838 );
and ( n237224 , n237223 , n38795 );
or ( n237225 , n237222 , n237224 );
not ( n237226 , n38807 );
and ( n237227 , n237225 , n237226 );
not ( n237228 , n237225 );
and ( n237229 , n237228 , n38801 );
nor ( n237230 , n237227 , n237229 );
not ( n237231 , n32680 );
not ( n237232 , n45313 );
or ( n237233 , n237231 , n237232 );
or ( n237234 , n45313 , n32680 );
nand ( n237235 , n237233 , n237234 );
and ( n237236 , n237235 , n48317 );
not ( n237237 , n237235 );
and ( n237238 , n237237 , n54849 );
nor ( n237239 , n237236 , n237238 );
nand ( n237240 , n237230 , n237239 );
not ( n237241 , n237240 );
not ( n237242 , n28357 );
not ( n237243 , n225836 );
not ( n237244 , n237243 );
or ( n237245 , n237242 , n237244 );
or ( n237246 , n36350 , n28357 );
nand ( n237247 , n237245 , n237246 );
and ( n237248 , n237247 , n40345 );
not ( n237249 , n237247 );
and ( n237250 , n237249 , n205846 );
nor ( n237251 , n237248 , n237250 );
not ( n237252 , n237251 );
not ( n237253 , n237252 );
and ( n237254 , n237241 , n237253 );
and ( n237255 , n237240 , n237252 );
nor ( n237256 , n237254 , n237255 );
and ( n237257 , n237221 , n237256 );
not ( n237258 , n237221 );
not ( n237259 , n237256 );
and ( n237260 , n237258 , n237259 );
nor ( n237261 , n237257 , n237260 );
xor ( n237262 , n30054 , n33299 );
xor ( n237263 , n237262 , n53417 );
not ( n237264 , n237263 );
not ( n237265 , n237264 );
not ( n237266 , n237265 );
not ( n237267 , n39920 );
not ( n237268 , n38140 );
or ( n237269 , n237267 , n237268 );
nand ( n237270 , n25676 , n39919 );
nand ( n237271 , n237269 , n237270 );
not ( n237272 , n237271 );
not ( n237273 , n25684 );
and ( n237274 , n237272 , n237273 );
and ( n237275 , n25684 , n237271 );
nor ( n237276 , n237274 , n237275 );
not ( n237277 , n29764 );
not ( n237278 , n46966 );
or ( n237279 , n237277 , n237278 );
or ( n237280 , n46966 , n29764 );
nand ( n237281 , n237279 , n237280 );
and ( n237282 , n237281 , n206591 );
not ( n237283 , n237281 );
and ( n237284 , n237283 , n28817 );
nor ( n237285 , n237282 , n237284 );
not ( n237286 , n237285 );
nand ( n237287 , n237276 , n237286 );
not ( n237288 , n237287 );
or ( n237289 , n237266 , n237288 );
or ( n237290 , n237287 , n237265 );
nand ( n237291 , n237289 , n237290 );
not ( n237292 , n237291 );
not ( n237293 , n237292 );
not ( n237294 , n31734 );
not ( n237295 , n32897 );
and ( n237296 , n237294 , n237295 );
and ( n237297 , n31734 , n32897 );
nor ( n237298 , n237296 , n237297 );
and ( n237299 , n237298 , n36710 );
not ( n237300 , n237298 );
and ( n237301 , n237300 , n31730 );
nor ( n237302 , n237299 , n237301 );
not ( n237303 , n237302 );
buf ( n237304 , n35764 );
not ( n237305 , n237304 );
not ( n237306 , n44615 );
or ( n237307 , n237305 , n237306 );
or ( n237308 , n44615 , n237304 );
nand ( n237309 , n237307 , n237308 );
and ( n237310 , n237309 , n43554 );
not ( n237311 , n237309 );
and ( n237312 , n237311 , n43803 );
nor ( n237313 , n237310 , n237312 );
not ( n237314 , n237313 );
nand ( n237315 , n237303 , n237314 );
not ( n237316 , n237315 );
not ( n237317 , n227134 );
not ( n237318 , n34820 );
or ( n237319 , n237317 , n237318 );
or ( n237320 , n34820 , n227134 );
nand ( n237321 , n237319 , n237320 );
and ( n237322 , n237321 , n207100 );
not ( n237323 , n237321 );
and ( n237324 , n237323 , n47134 );
nor ( n237325 , n237322 , n237324 );
buf ( n237326 , n237325 );
not ( n237327 , n237326 );
and ( n237328 , n237316 , n237327 );
and ( n237329 , n237315 , n237326 );
nor ( n237330 , n237328 , n237329 );
not ( n237331 , n237330 );
not ( n237332 , n237331 );
or ( n237333 , n237293 , n237332 );
nand ( n237334 , n237330 , n237291 );
nand ( n237335 , n237333 , n237334 );
and ( n237336 , n237261 , n237335 );
not ( n237337 , n237261 );
not ( n237338 , n237335 );
and ( n237339 , n237337 , n237338 );
nor ( n237340 , n237336 , n237339 );
not ( n237341 , n237340 );
not ( n237342 , n237341 );
and ( n237343 , n237150 , n237342 );
not ( n237344 , n237150 );
not ( n237345 , n237338 );
not ( n237346 , n237261 );
not ( n237347 , n237346 );
or ( n237348 , n237345 , n237347 );
nand ( n237349 , n237261 , n237335 );
nand ( n237350 , n237348 , n237349 );
and ( n237351 , n237344 , n237350 );
nor ( n237352 , n237343 , n237351 );
nand ( n237353 , n237000 , n237352 );
or ( n237354 , n236826 , n237353 );
not ( n237355 , n237000 );
not ( n237356 , n236825 );
or ( n237357 , n237355 , n237356 );
buf ( n237358 , n43968 );
nor ( n237359 , n237352 , n237358 );
nand ( n237360 , n237357 , n237359 );
buf ( n237361 , n35431 );
nand ( n237362 , n237361 , n37090 );
nand ( n237363 , n237354 , n237360 , n237362 );
buf ( n237364 , n237363 );
not ( n237365 , n49668 );
nand ( n237366 , n38809 , n237365 );
not ( n237367 , n237366 );
buf ( n237368 , n49657 );
not ( n237369 , n237368 );
and ( n237370 , n237367 , n237369 );
and ( n237371 , n237366 , n237368 );
nor ( n237372 , n237370 , n237371 );
not ( n237373 , n237372 );
not ( n237374 , n237373 );
not ( n237375 , n227548 );
or ( n237376 , n237374 , n237375 );
not ( n237377 , n237373 );
nand ( n237378 , n237377 , n227556 );
nand ( n237379 , n237376 , n237378 );
and ( n237380 , n237379 , n49947 );
not ( n237381 , n237379 );
and ( n237382 , n237381 , n49950 );
nor ( n237383 , n237380 , n237382 );
buf ( n237384 , n33252 );
not ( n237385 , n237384 );
nand ( n237386 , n237383 , n237385 );
not ( n237387 , n232756 );
nand ( n237388 , n54560 , n232698 );
not ( n237389 , n237388 );
not ( n237390 , n54549 );
or ( n237391 , n237389 , n237390 );
or ( n237392 , n54549 , n237388 );
nand ( n237393 , n237391 , n237392 );
not ( n237394 , n237393 );
not ( n237395 , n237394 );
nand ( n237396 , n54955 , n232720 );
not ( n237397 , n237396 );
not ( n237398 , n54712 );
and ( n237399 , n237397 , n237398 );
and ( n237400 , n237396 , n54712 );
nor ( n237401 , n237399 , n237400 );
not ( n237402 , n237401 );
not ( n237403 , n237402 );
or ( n237404 , n237395 , n237403 );
nand ( n237405 , n237401 , n237393 );
nand ( n237406 , n237404 , n237405 );
not ( n237407 , n232740 );
nand ( n237408 , n54990 , n237407 );
not ( n237409 , n237408 );
buf ( n237410 , n54676 );
not ( n237411 , n237410 );
and ( n237412 , n237409 , n237411 );
and ( n237413 , n237408 , n237410 );
nor ( n237414 , n237412 , n237413 );
not ( n237415 , n237414 );
and ( n237416 , n237406 , n237415 );
not ( n237417 , n237406 );
and ( n237418 , n237417 , n237414 );
nor ( n237419 , n237416 , n237418 );
nand ( n237420 , n55011 , n232784 );
not ( n237421 , n237420 );
not ( n237422 , n54627 );
and ( n237423 , n237421 , n237422 );
and ( n237424 , n237420 , n54627 );
nor ( n237425 , n237423 , n237424 );
not ( n237426 , n237425 );
not ( n237427 , n237426 );
not ( n237428 , n232368 );
nand ( n237429 , n55040 , n232812 );
not ( n237430 , n237429 );
or ( n237431 , n237428 , n237430 );
or ( n237432 , n237429 , n232368 );
nand ( n237433 , n237431 , n237432 );
not ( n237434 , n237433 );
not ( n237435 , n237434 );
or ( n237436 , n237427 , n237435 );
nand ( n237437 , n237433 , n237425 );
nand ( n237438 , n237436 , n237437 );
not ( n237439 , n237438 );
and ( n237440 , n237419 , n237439 );
not ( n237441 , n237419 );
and ( n237442 , n237441 , n237438 );
nor ( n237443 , n237440 , n237442 );
not ( n237444 , n237443 );
not ( n237445 , n237444 );
or ( n237446 , n237387 , n237445 );
not ( n237447 , n237443 );
not ( n237448 , n54998 );
or ( n237449 , n237447 , n237448 );
nand ( n237450 , n237446 , n237449 );
not ( n237451 , n237450 );
buf ( n237452 , n205212 );
not ( n237453 , n237452 );
not ( n237454 , n30220 );
or ( n237455 , n237453 , n237454 );
not ( n237456 , n237452 );
nand ( n237457 , n237456 , n204390 );
nand ( n237458 , n237455 , n237457 );
and ( n237459 , n237458 , n33685 );
not ( n237460 , n237458 );
and ( n237461 , n237460 , n31778 );
nor ( n237462 , n237459 , n237461 );
not ( n237463 , n237462 );
not ( n237464 , n35384 );
not ( n237465 , n46664 );
or ( n237466 , n237464 , n237465 );
not ( n237467 , n35384 );
nand ( n237468 , n237467 , n29645 );
nand ( n237469 , n237466 , n237468 );
and ( n237470 , n237469 , n46671 );
not ( n237471 , n237469 );
and ( n237472 , n237471 , n46668 );
nor ( n237473 , n237470 , n237472 );
nand ( n237474 , n237463 , n237473 );
and ( n237475 , n237474 , n232123 );
not ( n237476 , n237474 );
and ( n237477 , n237476 , n232122 );
nor ( n237478 , n237475 , n237477 );
not ( n237479 , n237478 );
not ( n237480 , n237479 );
not ( n237481 , n36227 );
not ( n237482 , n44860 );
or ( n237483 , n237481 , n237482 );
or ( n237484 , n44860 , n36227 );
nand ( n237485 , n237483 , n237484 );
and ( n237486 , n237485 , n28340 );
not ( n237487 , n237485 );
and ( n237488 , n237487 , n222628 );
nor ( n237489 , n237486 , n237488 );
buf ( n237490 , n31462 );
not ( n237491 , n237490 );
not ( n237492 , n38682 );
or ( n237493 , n237491 , n237492 );
or ( n237494 , n38682 , n237490 );
nand ( n237495 , n237493 , n237494 );
and ( n237496 , n237495 , n38690 );
not ( n237497 , n237495 );
and ( n237498 , n237497 , n38691 );
nor ( n237499 , n237496 , n237498 );
not ( n237500 , n237499 );
nand ( n237501 , n237489 , n237500 );
buf ( n237502 , n232152 );
xor ( n237503 , n237501 , n237502 );
not ( n237504 , n237503 );
not ( n237505 , n237504 );
or ( n237506 , n237480 , n237505 );
nand ( n237507 , n237503 , n237478 );
nand ( n237508 , n237506 , n237507 );
xor ( n237509 , n32048 , n31177 );
xnor ( n237510 , n237509 , n38677 );
not ( n237511 , n31007 );
not ( n237512 , n43554 );
or ( n237513 , n237511 , n237512 );
not ( n237514 , n31007 );
nand ( n237515 , n237514 , n43557 );
nand ( n237516 , n237513 , n237515 );
and ( n237517 , n237516 , n35063 );
not ( n237518 , n237516 );
and ( n237519 , n237518 , n45373 );
nor ( n237520 , n237517 , n237519 );
nand ( n237521 , n237510 , n237520 );
not ( n237522 , n237521 );
not ( n237523 , n54440 );
and ( n237524 , n237522 , n237523 );
and ( n237525 , n237521 , n54440 );
nor ( n237526 , n237524 , n237525 );
and ( n237527 , n237508 , n237526 );
not ( n237528 , n237508 );
not ( n237529 , n237526 );
and ( n237530 , n237528 , n237529 );
nor ( n237531 , n237527 , n237530 );
not ( n237532 , n237531 );
not ( n237533 , n232243 );
not ( n237534 , n237533 );
not ( n237535 , n237534 );
buf ( n237536 , n34983 );
not ( n237537 , n237536 );
not ( n237538 , n34980 );
and ( n237539 , n237537 , n237538 );
and ( n237540 , n237536 , n34980 );
nor ( n237541 , n237539 , n237540 );
and ( n237542 , n237541 , n204347 );
not ( n237543 , n237541 );
and ( n237544 , n237543 , n229721 );
nor ( n237545 , n237542 , n237544 );
not ( n237546 , n31932 );
and ( n237547 , n237545 , n237546 );
not ( n237548 , n237545 );
and ( n237549 , n237548 , n31932 );
nor ( n237550 , n237547 , n237549 );
not ( n237551 , n237550 );
xor ( n237552 , n33133 , n227301 );
xnor ( n237553 , n237552 , n39020 );
not ( n237554 , n237553 );
nand ( n237555 , n237551 , n237554 );
not ( n237556 , n237555 );
or ( n237557 , n237535 , n237556 );
or ( n237558 , n237555 , n237534 );
nand ( n237559 , n237557 , n237558 );
not ( n237560 , n237559 );
buf ( n237561 , n28501 );
buf ( n237562 , n36262 );
xor ( n237563 , n237561 , n237562 );
xnor ( n237564 , n237563 , n32863 );
not ( n237565 , n237564 );
buf ( n237566 , n28338 );
not ( n237567 , n237566 );
not ( n237568 , n237567 );
not ( n237569 , n36309 );
or ( n237570 , n237568 , n237569 );
nand ( n237571 , n36312 , n237566 );
nand ( n237572 , n237570 , n237571 );
buf ( n237573 , n49318 );
xnor ( n237574 , n237572 , n237573 );
not ( n237575 , n237574 );
nand ( n237576 , n237565 , n237575 );
not ( n237577 , n237576 );
not ( n237578 , n232261 );
and ( n237579 , n237577 , n237578 );
and ( n237580 , n237576 , n232261 );
nor ( n237581 , n237579 , n237580 );
not ( n237582 , n237581 );
or ( n237583 , n237560 , n237582 );
or ( n237584 , n237581 , n237559 );
nand ( n237585 , n237583 , n237584 );
not ( n237586 , n237585 );
or ( n237587 , n237532 , n237586 );
or ( n237588 , n237585 , n237531 );
nand ( n237589 , n237587 , n237588 );
buf ( n237590 , n237589 );
not ( n237591 , n237590 );
not ( n237592 , n237591 );
and ( n237593 , n237451 , n237592 );
not ( n237594 , n237590 );
and ( n237595 , n237450 , n237594 );
nor ( n237596 , n237593 , n237595 );
not ( n237597 , n42644 );
not ( n237598 , n233980 );
not ( n237599 , n42554 );
nand ( n237600 , n237599 , n40986 );
and ( n237601 , n237600 , n41029 );
not ( n237602 , n237600 );
and ( n237603 , n237602 , n41028 );
nor ( n237604 , n237601 , n237603 );
not ( n237605 , n237604 );
or ( n237606 , n237598 , n237605 );
or ( n237607 , n237604 , n233980 );
nand ( n237608 , n237606 , n237607 );
not ( n237609 , n41069 );
nand ( n237610 , n237609 , n42523 );
not ( n237611 , n237610 );
not ( n237612 , n231990 );
or ( n237613 , n237611 , n237612 );
or ( n237614 , n231990 , n237610 );
nand ( n237615 , n237613 , n237614 );
and ( n237616 , n237608 , n237615 );
not ( n237617 , n237608 );
not ( n237618 , n237615 );
and ( n237619 , n237617 , n237618 );
nor ( n237620 , n237616 , n237619 );
not ( n237621 , n237620 );
nand ( n237622 , n41171 , n220238 );
xnor ( n237623 , n237622 , n41201 );
not ( n237624 , n237623 );
nand ( n237625 , n42683 , n41161 );
not ( n237626 , n237625 );
not ( n237627 , n54249 );
and ( n237628 , n237626 , n237627 );
and ( n237629 , n237625 , n54249 );
nor ( n237630 , n237628 , n237629 );
not ( n237631 , n237630 );
and ( n237632 , n237624 , n237631 );
and ( n237633 , n237623 , n237630 );
nor ( n237634 , n237632 , n237633 );
not ( n237635 , n237634 );
and ( n237636 , n237621 , n237635 );
not ( n237637 , n237621 );
and ( n237638 , n237637 , n237634 );
nor ( n237639 , n237636 , n237638 );
not ( n237640 , n237639 );
or ( n237641 , n237597 , n237640 );
not ( n237642 , n42644 );
not ( n237643 , n237634 );
not ( n237644 , n237620 );
or ( n237645 , n237643 , n237644 );
nand ( n237646 , n237621 , n237635 );
nand ( n237647 , n237645 , n237646 );
nand ( n237648 , n237642 , n237647 );
nand ( n237649 , n237641 , n237648 );
not ( n237650 , n54277 );
nand ( n237651 , n49967 , n42831 );
not ( n237652 , n237651 );
or ( n237653 , n237650 , n237652 );
not ( n237654 , n220589 );
nand ( n237655 , n237654 , n49967 );
or ( n237656 , n237655 , n54277 );
nand ( n237657 , n237653 , n237656 );
not ( n237658 , n237657 );
not ( n237659 , n220481 );
nand ( n237660 , n237659 , n229049 );
not ( n237661 , n237660 );
not ( n237662 , n44164 );
not ( n237663 , n237662 );
and ( n237664 , n237661 , n237663 );
and ( n237665 , n237660 , n237662 );
nor ( n237666 , n237664 , n237665 );
not ( n237667 , n237666 );
or ( n237668 , n237658 , n237667 );
or ( n237669 , n237666 , n237657 );
nand ( n237670 , n237668 , n237669 );
not ( n237671 , n237670 );
not ( n237672 , n237671 );
not ( n237673 , n43994 );
not ( n237674 , n229037 );
not ( n237675 , n42866 );
nand ( n237676 , n237675 , n220613 );
not ( n237677 , n237676 );
or ( n237678 , n237674 , n237677 );
or ( n237679 , n237676 , n229037 );
nand ( n237680 , n237678 , n237679 );
not ( n237681 , n237680 );
and ( n237682 , n237673 , n237681 );
and ( n237683 , n43994 , n237680 );
nor ( n237684 , n237682 , n237683 );
nand ( n237685 , n51310 , n42884 );
not ( n237686 , n237685 );
not ( n237687 , n44028 );
and ( n237688 , n237686 , n237687 );
and ( n237689 , n237685 , n44028 );
nor ( n237690 , n237688 , n237689 );
and ( n237691 , n237684 , n237690 );
not ( n237692 , n237684 );
not ( n237693 , n237690 );
and ( n237694 , n237692 , n237693 );
nor ( n237695 , n237691 , n237694 );
not ( n237696 , n237695 );
or ( n237697 , n237672 , n237696 );
or ( n237698 , n237695 , n237671 );
nand ( n237699 , n237697 , n237698 );
buf ( n237700 , n237699 );
not ( n237701 , n237700 );
and ( n237702 , n237649 , n237701 );
not ( n237703 , n237649 );
buf ( n237704 , n237700 );
and ( n237705 , n237703 , n237704 );
nor ( n237706 , n237702 , n237705 );
nand ( n237707 , n237596 , n237706 );
or ( n237708 , n237386 , n237707 );
not ( n237709 , n237706 );
not ( n237710 , n237383 );
or ( n237711 , n237709 , n237710 );
nor ( n237712 , n237596 , n235050 );
nand ( n237713 , n237711 , n237712 );
buf ( n237714 , n35431 );
nand ( n237715 , n237714 , n29107 );
nand ( n237716 , n237708 , n237713 , n237715 );
buf ( n237717 , n237716 );
buf ( n237718 , n41006 );
not ( n237719 , n54071 );
nand ( n237720 , n39536 , n237719 );
and ( n237721 , n237720 , n34737 );
not ( n237722 , n237720 );
not ( n237723 , n34737 );
and ( n237724 , n237722 , n237723 );
nor ( n237725 , n237721 , n237724 );
not ( n237726 , n237725 );
not ( n237727 , n39595 );
or ( n237728 , n237726 , n237727 );
not ( n237729 , n237725 );
nand ( n237730 , n237729 , n39598 );
nand ( n237731 , n237728 , n237730 );
and ( n237732 , n237731 , n217511 );
not ( n237733 , n237731 );
and ( n237734 , n237733 , n217515 );
nor ( n237735 , n237732 , n237734 );
nor ( n237736 , n237735 , n235050 );
nand ( n237737 , n229218 , n51463 );
not ( n237738 , n237737 );
not ( n237739 , n36094 );
not ( n237740 , n237739 );
and ( n237741 , n237738 , n237740 );
and ( n237742 , n237737 , n237739 );
nor ( n237743 , n237741 , n237742 );
not ( n237744 , n237743 );
not ( n237745 , n237744 );
not ( n237746 , n36372 );
not ( n237747 , n237746 );
or ( n237748 , n237745 , n237747 );
not ( n237749 , n237744 );
nand ( n237750 , n237749 , n36372 );
nand ( n237751 , n237748 , n237750 );
not ( n237752 , n237751 );
not ( n237753 , n36730 );
and ( n237754 , n237752 , n237753 );
and ( n237755 , n237751 , n36730 );
nor ( n237756 , n237754 , n237755 );
not ( n237757 , n44707 );
nand ( n237758 , n44688 , n222435 );
not ( n237759 , n237758 );
not ( n237760 , n235303 );
or ( n237761 , n237759 , n237760 );
or ( n237762 , n235303 , n237758 );
nand ( n237763 , n237761 , n237762 );
not ( n237764 , n237763 );
or ( n237765 , n44746 , n44734 );
not ( n237766 , n237765 );
not ( n237767 , n235293 );
and ( n237768 , n237766 , n237767 );
and ( n237769 , n237765 , n235293 );
nor ( n237770 , n237768 , n237769 );
not ( n237771 , n237770 );
and ( n237772 , n237764 , n237771 );
and ( n237773 , n237763 , n237770 );
nor ( n237774 , n237772 , n237773 );
not ( n237775 , n237774 );
not ( n237776 , n235341 );
nand ( n237777 , n222328 , n44555 );
not ( n237778 , n237777 );
or ( n237779 , n237776 , n237778 );
or ( n237780 , n237777 , n235341 );
nand ( n237781 , n237779 , n237780 );
not ( n237782 , n237781 );
nand ( n237783 , n44653 , n44644 );
not ( n237784 , n237783 );
not ( n237785 , n235225 );
and ( n237786 , n237784 , n237785 );
and ( n237787 , n237783 , n235225 );
nor ( n237788 , n237786 , n237787 );
not ( n237789 , n237788 );
or ( n237790 , n237782 , n237789 );
or ( n237791 , n237788 , n237781 );
nand ( n237792 , n237790 , n237791 );
not ( n237793 , n44594 );
nand ( n237794 , n237793 , n44617 );
not ( n237795 , n237794 );
not ( n237796 , n235254 );
and ( n237797 , n237795 , n237796 );
and ( n237798 , n237794 , n235254 );
nor ( n237799 , n237797 , n237798 );
and ( n237800 , n237792 , n237799 );
not ( n237801 , n237792 );
not ( n237802 , n237799 );
and ( n237803 , n237801 , n237802 );
nor ( n237804 , n237800 , n237803 );
not ( n237805 , n237804 );
not ( n237806 , n237805 );
or ( n237807 , n237775 , n237806 );
not ( n237808 , n237774 );
nand ( n237809 , n237804 , n237808 );
nand ( n237810 , n237807 , n237809 );
not ( n237811 , n237810 );
or ( n237812 , n237757 , n237811 );
not ( n237813 , n44707 );
and ( n237814 , n237804 , n237808 );
not ( n237815 , n237804 );
and ( n237816 , n237815 , n237774 );
nor ( n237817 , n237814 , n237816 );
nand ( n237818 , n237813 , n237817 );
nand ( n237819 , n237812 , n237818 );
not ( n237820 , n50674 );
nand ( n237821 , n237820 , n50632 );
not ( n237822 , n237821 );
not ( n237823 , n46819 );
and ( n237824 , n237822 , n237823 );
and ( n237825 , n237821 , n46819 );
nor ( n237826 , n237824 , n237825 );
not ( n237827 , n237826 );
nand ( n237828 , n50653 , n50649 );
not ( n237829 , n46770 );
and ( n237830 , n237828 , n237829 );
not ( n237831 , n237828 );
and ( n237832 , n237831 , n46770 );
nor ( n237833 , n237830 , n237832 );
not ( n237834 , n237833 );
or ( n237835 , n237827 , n237834 );
or ( n237836 , n237826 , n237833 );
nand ( n237837 , n237835 , n237836 );
not ( n237838 , n46854 );
nand ( n237839 , n228466 , n50693 );
not ( n237840 , n237839 );
and ( n237841 , n237838 , n237840 );
and ( n237842 , n46854 , n237839 );
nor ( n237843 , n237841 , n237842 );
and ( n237844 , n237837 , n237843 );
not ( n237845 , n237837 );
not ( n237846 , n237843 );
and ( n237847 , n237845 , n237846 );
nor ( n237848 , n237844 , n237847 );
not ( n237849 , n46909 );
not ( n237850 , n50727 );
nand ( n237851 , n50731 , n237850 );
not ( n237852 , n237851 );
or ( n237853 , n237849 , n237852 );
or ( n237854 , n237851 , n46909 );
nand ( n237855 , n237853 , n237854 );
not ( n237856 , n237855 );
nand ( n237857 , n46728 , n50749 );
not ( n237858 , n237857 );
not ( n237859 , n224634 );
and ( n237860 , n237858 , n237859 );
and ( n237861 , n237857 , n224634 );
nor ( n237862 , n237860 , n237861 );
not ( n237863 , n237862 );
and ( n237864 , n237856 , n237863 );
and ( n237865 , n237855 , n237862 );
nor ( n237866 , n237864 , n237865 );
xnor ( n237867 , n237848 , n237866 );
buf ( n237868 , n237867 );
not ( n237869 , n237868 );
and ( n237870 , n237819 , n237869 );
not ( n237871 , n237819 );
and ( n237872 , n237871 , n237868 );
nor ( n237873 , n237870 , n237872 );
not ( n237874 , n237873 );
nand ( n237875 , n237736 , n237756 , n237874 );
not ( n237876 , n237735 );
not ( n237877 , n237876 );
not ( n237878 , n237756 );
or ( n237879 , n237877 , n237878 );
nor ( n237880 , n237874 , n226955 );
nand ( n237881 , n237879 , n237880 );
nand ( n237882 , n237714 , n31144 );
nand ( n237883 , n237875 , n237881 , n237882 );
buf ( n237884 , n237883 );
not ( n237885 , n54810 );
nand ( n237886 , n54880 , n54890 );
not ( n237887 , n237886 );
not ( n237888 , n45063 );
and ( n237889 , n237887 , n237888 );
and ( n237890 , n237886 , n45063 );
nor ( n237891 , n237889 , n237890 );
nand ( n237892 , n54902 , n54780 );
buf ( n237893 , n45080 );
xnor ( n237894 , n237892 , n237893 );
and ( n237895 , n237891 , n237894 );
not ( n237896 , n237891 );
not ( n237897 , n237894 );
and ( n237898 , n237896 , n237897 );
nor ( n237899 , n237895 , n237898 );
not ( n237900 , n237899 );
not ( n237901 , n237900 );
nand ( n237902 , n54867 , n54853 );
not ( n237903 , n237902 );
not ( n237904 , n222997 );
and ( n237905 , n237903 , n237904 );
and ( n237906 , n237902 , n222997 );
nor ( n237907 , n237905 , n237906 );
not ( n237908 , n237907 );
nand ( n237909 , n54820 , n54832 );
not ( n237910 , n237909 );
not ( n237911 , n45159 );
or ( n237912 , n237910 , n237911 );
or ( n237913 , n45159 , n237909 );
nand ( n237914 , n237912 , n237913 );
not ( n237915 , n237914 );
or ( n237916 , n237908 , n237915 );
or ( n237917 , n237914 , n237907 );
nand ( n237918 , n237916 , n237917 );
not ( n237919 , n232556 );
not ( n237920 , n54805 );
nand ( n237921 , n237919 , n237920 );
not ( n237922 , n237921 );
not ( n237923 , n222878 );
and ( n237924 , n237922 , n237923 );
and ( n237925 , n237921 , n222878 );
nor ( n237926 , n237924 , n237925 );
not ( n237927 , n237926 );
and ( n237928 , n237918 , n237927 );
not ( n237929 , n237918 );
and ( n237930 , n237929 , n237926 );
nor ( n237931 , n237928 , n237930 );
not ( n237932 , n237931 );
not ( n237933 , n237932 );
and ( n237934 , n237901 , n237933 );
and ( n237935 , n237900 , n237932 );
nor ( n237936 , n237934 , n237935 );
not ( n237937 , n237936 );
or ( n237938 , n237885 , n237937 );
not ( n237939 , n54810 );
not ( n237940 , n237931 );
not ( n237941 , n237899 );
or ( n237942 , n237940 , n237941 );
nand ( n237943 , n237900 , n237932 );
nand ( n237944 , n237942 , n237943 );
nand ( n237945 , n237939 , n237944 );
nand ( n237946 , n237938 , n237945 );
not ( n237947 , n237447 );
not ( n237948 , n237947 );
and ( n237949 , n237946 , n237948 );
not ( n237950 , n237946 );
and ( n237951 , n237950 , n237947 );
nor ( n237952 , n237949 , n237951 );
not ( n237953 , n237952 );
not ( n237954 , n237953 );
buf ( n237955 , n38347 );
xor ( n237956 , n41001 , n237955 );
xnor ( n237957 , n237956 , n43787 );
not ( n237958 , n237957 );
nand ( n237959 , n237958 , n44997 );
and ( n237960 , n237959 , n44982 );
not ( n237961 , n237959 );
and ( n237962 , n237961 , n44981 );
nor ( n237963 , n237960 , n237962 );
not ( n237964 , n237963 );
not ( n237965 , n45026 );
or ( n237966 , n237964 , n237965 );
not ( n237967 , n237963 );
nand ( n237968 , n237967 , n45023 );
nand ( n237969 , n237966 , n237968 );
and ( n237970 , n237969 , n223016 );
not ( n237971 , n237969 );
and ( n237972 , n237971 , n45262 );
nor ( n237973 , n237970 , n237972 );
not ( n237974 , n237973 );
or ( n237975 , n237954 , n237974 );
not ( n237976 , n47572 );
not ( n237977 , n48510 );
not ( n237978 , n237977 );
not ( n237979 , n47641 );
nand ( n237980 , n237979 , n234861 );
not ( n237981 , n237980 );
or ( n237982 , n237978 , n237981 );
nand ( n237983 , n237979 , n234861 );
or ( n237984 , n237983 , n237977 );
nand ( n237985 , n237982 , n237984 );
not ( n237986 , n237985 );
nand ( n237987 , n234849 , n225467 );
not ( n237988 , n237987 );
not ( n237989 , n48430 );
and ( n237990 , n237988 , n237989 );
and ( n237991 , n237987 , n48430 );
nor ( n237992 , n237990 , n237991 );
not ( n237993 , n237992 );
or ( n237994 , n237986 , n237993 );
or ( n237995 , n237992 , n237985 );
nand ( n237996 , n237994 , n237995 );
not ( n237997 , n237996 );
not ( n237998 , n237997 );
not ( n237999 , n47620 );
nand ( n238000 , n237999 , n234425 );
not ( n238001 , n238000 );
buf ( n238002 , n48451 );
not ( n238003 , n238002 );
and ( n238004 , n238001 , n238003 );
and ( n238005 , n238000 , n238002 );
nor ( n238006 , n238004 , n238005 );
not ( n238007 , n238006 );
not ( n238008 , n238007 );
or ( n238009 , n237998 , n238008 );
nand ( n238010 , n238006 , n237996 );
nand ( n238011 , n238009 , n238010 );
not ( n238012 , n225512 );
nand ( n238013 , n234867 , n238012 );
not ( n238014 , n238013 );
not ( n238015 , n226255 );
not ( n238016 , n238015 );
and ( n238017 , n238014 , n238016 );
and ( n238018 , n238013 , n238015 );
nor ( n238019 , n238017 , n238018 );
not ( n238020 , n238019 );
not ( n238021 , n238020 );
nand ( n238022 , n225328 , n47552 );
xor ( n238023 , n238022 , n48534 );
not ( n238024 , n238023 );
not ( n238025 , n238024 );
or ( n238026 , n238021 , n238025 );
nand ( n238027 , n238023 , n238019 );
nand ( n238028 , n238026 , n238027 );
not ( n238029 , n238028 );
and ( n238030 , n238011 , n238029 );
not ( n238031 , n238011 );
and ( n238032 , n238031 , n238028 );
nor ( n238033 , n238030 , n238032 );
not ( n238034 , n238033 );
or ( n238035 , n237976 , n238034 );
not ( n238036 , n47572 );
and ( n238037 , n238011 , n238028 );
not ( n238038 , n238011 );
and ( n238039 , n238038 , n238029 );
nor ( n238040 , n238037 , n238039 );
nand ( n238041 , n238036 , n238040 );
nand ( n238042 , n238035 , n238041 );
nand ( n238043 , n234356 , n48621 );
and ( n238044 , n238043 , n47985 );
not ( n238045 , n238043 );
and ( n238046 , n238045 , n47968 );
nor ( n238047 , n238044 , n238046 );
not ( n238048 , n238047 );
not ( n238049 , n238048 );
nand ( n238050 , n226358 , n234363 );
not ( n238051 , n238050 );
not ( n238052 , n47868 );
not ( n238053 , n238052 );
and ( n238054 , n238051 , n238053 );
and ( n238055 , n238050 , n238052 );
nor ( n238056 , n238054 , n238055 );
not ( n238057 , n238056 );
not ( n238058 , n238057 );
or ( n238059 , n238049 , n238058 );
nand ( n238060 , n238056 , n238047 );
nand ( n238061 , n238059 , n238060 );
not ( n238062 , n234381 );
nand ( n238063 , n238062 , n226339 );
not ( n238064 , n238063 );
not ( n238065 , n47841 );
and ( n238066 , n238064 , n238065 );
not ( n238067 , n234381 );
nand ( n238068 , n238067 , n226339 );
and ( n238069 , n238068 , n47841 );
nor ( n238070 , n238066 , n238069 );
and ( n238071 , n238061 , n238070 );
not ( n238072 , n238061 );
not ( n238073 , n238070 );
and ( n238074 , n238072 , n238073 );
nor ( n238075 , n238071 , n238074 );
nand ( n238076 , n48662 , n47792 );
not ( n238077 , n238076 );
not ( n238078 , n47781 );
or ( n238079 , n238077 , n238078 );
nand ( n238080 , n48662 , n47792 );
or ( n238081 , n47781 , n238080 );
nand ( n238082 , n238079 , n238081 );
not ( n238083 , n238082 );
not ( n238084 , n238083 );
not ( n238085 , n48645 );
nand ( n238086 , n238085 , n234396 );
not ( n238087 , n238086 );
not ( n238088 , n47914 );
and ( n238089 , n238087 , n238088 );
and ( n238090 , n238086 , n47914 );
nor ( n238091 , n238089 , n238090 );
not ( n238092 , n238091 );
not ( n238093 , n238092 );
or ( n238094 , n238084 , n238093 );
nand ( n238095 , n238091 , n238082 );
nand ( n238096 , n238094 , n238095 );
and ( n238097 , n238075 , n238096 );
not ( n238098 , n238075 );
not ( n238099 , n238096 );
and ( n238100 , n238098 , n238099 );
nor ( n238101 , n238097 , n238100 );
buf ( n238102 , n238101 );
and ( n238103 , n238042 , n238102 );
not ( n238104 , n238042 );
xor ( n238105 , n238070 , n238061 );
xnor ( n238106 , n238105 , n238096 );
buf ( n238107 , n238106 );
and ( n238108 , n238104 , n238107 );
nor ( n238109 , n238103 , n238108 );
nor ( n238110 , n238109 , n49051 );
nand ( n238111 , n237975 , n238110 );
nor ( n238112 , n237952 , n49959 );
nand ( n238113 , n238112 , n237973 , n238109 );
buf ( n238114 , n35431 );
nand ( n238115 , n238114 , n28539 );
nand ( n238116 , n238111 , n238113 , n238115 );
buf ( n238117 , n238116 );
not ( n238118 , n33660 );
not ( n238119 , n51381 );
or ( n238120 , n238118 , n238119 );
not ( n238121 , n233579 );
not ( n238122 , n49181 );
or ( n238123 , n238121 , n238122 );
not ( n238124 , n233579 );
nand ( n238125 , n238124 , n49190 );
nand ( n238126 , n238123 , n238125 );
not ( n238127 , n45697 );
nand ( n238128 , n238127 , n233786 );
not ( n238129 , n238128 );
not ( n238130 , n45688 );
and ( n238131 , n238129 , n238130 );
and ( n238132 , n238128 , n45688 );
nor ( n238133 , n238131 , n238132 );
not ( n238134 , n238133 );
not ( n238135 , n238134 );
nand ( n238136 , n45625 , n55974 );
not ( n238137 , n238136 );
not ( n238138 , n45611 );
and ( n238139 , n238137 , n238138 );
and ( n238140 , n238136 , n45611 );
nor ( n238141 , n238139 , n238140 );
not ( n238142 , n238141 );
nand ( n238143 , n223416 , n233762 );
and ( n238144 , n238143 , n45667 );
not ( n238145 , n238143 );
and ( n238146 , n238145 , n45666 );
nor ( n238147 , n238144 , n238146 );
not ( n238148 , n238147 );
or ( n238149 , n238142 , n238148 );
or ( n238150 , n238147 , n238141 );
nand ( n238151 , n238149 , n238150 );
not ( n238152 , n238151 );
not ( n238153 , n238152 );
or ( n238154 , n238135 , n238153 );
nand ( n238155 , n238151 , n238133 );
nand ( n238156 , n238154 , n238155 );
not ( n238157 , n45533 );
not ( n238158 , n238157 );
not ( n238159 , n233704 );
nand ( n238160 , n238159 , n233716 );
not ( n238161 , n238160 );
or ( n238162 , n238158 , n238161 );
or ( n238163 , n238160 , n238157 );
nand ( n238164 , n238162 , n238163 );
not ( n238165 , n238164 );
buf ( n238166 , n233674 );
nand ( n238167 , n45578 , n238166 );
not ( n238168 , n238167 );
not ( n238169 , n45567 );
not ( n238170 , n238169 );
and ( n238171 , n238168 , n238170 );
and ( n238172 , n238167 , n238169 );
nor ( n238173 , n238171 , n238172 );
not ( n238174 , n238173 );
and ( n238175 , n238165 , n238174 );
and ( n238176 , n238164 , n238173 );
nor ( n238177 , n238175 , n238176 );
and ( n238178 , n238156 , n238177 );
not ( n238179 , n238156 );
not ( n238180 , n238177 );
and ( n238181 , n238179 , n238180 );
nor ( n238182 , n238178 , n238181 );
buf ( n238183 , n238182 );
and ( n238184 , n238126 , n238183 );
not ( n238185 , n238126 );
not ( n238186 , n238183 );
and ( n238187 , n238185 , n238186 );
nor ( n238188 , n238184 , n238187 );
not ( n238189 , n50540 );
not ( n238190 , n204267 );
not ( n238191 , n50595 );
or ( n238192 , n238190 , n238191 );
or ( n238193 , n50595 , n204267 );
nand ( n238194 , n238192 , n238193 );
not ( n238195 , n238194 );
not ( n238196 , n238195 );
or ( n238197 , n238189 , n238196 );
nand ( n238198 , n50604 , n238194 );
nand ( n238199 , n238197 , n238198 );
nand ( n238200 , n238188 , n238199 );
not ( n238201 , n33405 );
not ( n238202 , n28386 );
nand ( n238203 , n28513 , n238202 );
not ( n238204 , n238203 );
and ( n238205 , n238201 , n238204 );
and ( n238206 , n33405 , n238203 );
nor ( n238207 , n238205 , n238206 );
not ( n238208 , n238207 );
not ( n238209 , n55345 );
or ( n238210 , n238208 , n238209 );
not ( n238211 , n238207 );
nand ( n238212 , n238211 , n33708 );
nand ( n238213 , n238210 , n238212 );
and ( n238214 , n238213 , n55511 );
not ( n238215 , n238213 );
and ( n238216 , n238215 , n233265 );
nor ( n238217 , n238214 , n238216 );
not ( n238218 , n238217 );
and ( n238219 , n238200 , n238218 );
not ( n238220 , n238200 );
and ( n238221 , n238220 , n238217 );
nor ( n238222 , n238219 , n238221 );
buf ( n238223 , n40465 );
or ( n238224 , n238222 , n238223 );
nand ( n238225 , n238120 , n238224 );
buf ( n238226 , n238225 );
not ( n238227 , RI19a88a00_2734);
or ( n238228 , n25328 , n238227 );
not ( n238229 , RI19acc9f8_2234);
or ( n238230 , n25335 , n238229 );
nand ( n238231 , n238228 , n238230 );
buf ( n238232 , n238231 );
not ( n238233 , n53735 );
not ( n238234 , n231475 );
nand ( n238235 , n238234 , n228079 );
not ( n238236 , n238235 );
not ( n238237 , n236072 );
not ( n238238 , n238237 );
and ( n238239 , n238236 , n238238 );
and ( n238240 , n238235 , n238237 );
nor ( n238241 , n238239 , n238240 );
not ( n238242 , n238241 );
nand ( n238243 , n53730 , n50349 );
and ( n238244 , n238243 , n236111 );
not ( n238245 , n238243 );
and ( n238246 , n238245 , n236110 );
nor ( n238247 , n238244 , n238246 );
not ( n238248 , n238247 );
or ( n238249 , n238242 , n238248 );
or ( n238250 , n238247 , n238241 );
nand ( n238251 , n238249 , n238250 );
nand ( n238252 , n50385 , n53751 );
and ( n238253 , n238252 , n236091 );
not ( n238254 , n238252 );
and ( n238255 , n238254 , n236090 );
nor ( n238256 , n238253 , n238255 );
and ( n238257 , n238251 , n238256 );
not ( n238258 , n238251 );
not ( n238259 , n238256 );
and ( n238260 , n238258 , n238259 );
nor ( n238261 , n238257 , n238260 );
not ( n238262 , n238261 );
nand ( n238263 , n228222 , n53774 );
not ( n238264 , n238263 );
not ( n238265 , n236131 );
not ( n238266 , n238265 );
and ( n238267 , n238264 , n238266 );
and ( n238268 , n238263 , n238265 );
nor ( n238269 , n238267 , n238268 );
not ( n238270 , n238269 );
not ( n238271 , n236152 );
not ( n238272 , n238271 );
nand ( n238273 , n53796 , n50406 );
not ( n238274 , n238273 );
or ( n238275 , n238272 , n238274 );
not ( n238276 , n50405 );
nand ( n238277 , n238276 , n53796 );
or ( n238278 , n238277 , n238271 );
nand ( n238279 , n238275 , n238278 );
not ( n238280 , n238279 );
or ( n238281 , n238270 , n238280 );
or ( n238282 , n238279 , n238269 );
nand ( n238283 , n238281 , n238282 );
not ( n238284 , n238283 );
not ( n238285 , n238284 );
and ( n238286 , n238262 , n238285 );
and ( n238287 , n238261 , n238284 );
nor ( n238288 , n238286 , n238287 );
not ( n238289 , n238288 );
or ( n238290 , n238233 , n238289 );
not ( n238291 , n53735 );
not ( n238292 , n238284 );
not ( n238293 , n238261 );
or ( n238294 , n238292 , n238293 );
not ( n238295 , n238261 );
nand ( n238296 , n238295 , n238283 );
nand ( n238297 , n238294 , n238296 );
nand ( n238298 , n238291 , n238297 );
nand ( n238299 , n238290 , n238298 );
nand ( n238300 , n231615 , n231591 );
not ( n238301 , n238300 );
not ( n238302 , n34531 );
not ( n238303 , n44136 );
or ( n238304 , n238302 , n238303 );
not ( n238305 , n34531 );
nand ( n238306 , n238305 , n44135 );
nand ( n238307 , n238304 , n238306 );
and ( n238308 , n238307 , n44161 );
not ( n238309 , n238307 );
and ( n238310 , n238309 , n45281 );
nor ( n238311 , n238308 , n238310 );
not ( n238312 , n238311 );
not ( n238313 , n238312 );
and ( n238314 , n238301 , n238313 );
and ( n238315 , n238300 , n238312 );
nor ( n238316 , n238314 , n238315 );
nand ( n238317 , n53863 , n53883 );
not ( n238318 , n238317 );
not ( n238319 , n26444 );
not ( n238320 , n31695 );
or ( n238321 , n238319 , n238320 );
nand ( n238322 , n31694 , n26440 );
nand ( n238323 , n238321 , n238322 );
and ( n238324 , n238323 , n31727 );
not ( n238325 , n238323 );
and ( n238326 , n238325 , n31724 );
or ( n238327 , n238324 , n238326 );
and ( n238328 , n238327 , n29815 );
not ( n238329 , n238327 );
and ( n238330 , n238329 , n44471 );
nor ( n238331 , n238328 , n238330 );
not ( n238332 , n238331 );
not ( n238333 , n238332 );
and ( n238334 , n238318 , n238333 );
and ( n238335 , n238317 , n238332 );
nor ( n238336 , n238334 , n238335 );
xor ( n238337 , n238316 , n238336 );
not ( n238338 , n231658 );
nand ( n238339 , n231676 , n238338 );
not ( n238340 , n238339 );
not ( n238341 , n39401 );
not ( n238342 , n29104 );
not ( n238343 , n36262 );
or ( n238344 , n238342 , n238343 );
not ( n238345 , n29104 );
nand ( n238346 , n238345 , n210587 );
nand ( n238347 , n238344 , n238346 );
not ( n238348 , n238347 );
or ( n238349 , n238341 , n238348 );
or ( n238350 , n238347 , n39401 );
nand ( n238351 , n238349 , n238350 );
buf ( n238352 , n238351 );
not ( n238353 , n238352 );
and ( n238354 , n238340 , n238353 );
and ( n238355 , n238339 , n238352 );
nor ( n238356 , n238354 , n238355 );
xnor ( n238357 , n238337 , n238356 );
not ( n238358 , n238357 );
not ( n238359 , n53922 );
nand ( n238360 , n238359 , n231688 );
not ( n238361 , n238360 );
not ( n238362 , n38273 );
not ( n238363 , n229250 );
or ( n238364 , n238362 , n238363 );
nand ( n238365 , n30893 , n38269 );
nand ( n238366 , n238364 , n238365 );
xnor ( n238367 , n238366 , n34004 );
buf ( n238368 , n238367 );
not ( n238369 , n238368 );
and ( n238370 , n238361 , n238369 );
and ( n238371 , n238360 , n238368 );
nor ( n238372 , n238370 , n238371 );
not ( n238373 , n238372 );
not ( n238374 , n238373 );
not ( n238375 , n53960 );
nand ( n238376 , n238375 , n231754 );
not ( n238377 , n238376 );
not ( n238378 , n38160 );
not ( n238379 , n34103 );
or ( n238380 , n238378 , n238379 );
nand ( n238381 , n34089 , n38156 );
nand ( n238382 , n238380 , n238381 );
and ( n238383 , n238382 , n40369 );
not ( n238384 , n238382 );
and ( n238385 , n238384 , n40169 );
nor ( n238386 , n238383 , n238385 );
not ( n238387 , n238386 );
not ( n238388 , n238387 );
and ( n238389 , n238377 , n238388 );
and ( n238390 , n238376 , n238387 );
nor ( n238391 , n238389 , n238390 );
not ( n238392 , n238391 );
and ( n238393 , n238374 , n238392 );
and ( n238394 , n238373 , n238391 );
nor ( n238395 , n238393 , n238394 );
not ( n238396 , n238395 );
and ( n238397 , n238358 , n238396 );
not ( n238398 , n238358 );
and ( n238399 , n238398 , n238395 );
nor ( n238400 , n238397 , n238399 );
buf ( n238401 , n238400 );
and ( n238402 , n238299 , n238401 );
not ( n238403 , n238299 );
not ( n238404 , n238395 );
not ( n238405 , n238357 );
or ( n238406 , n238404 , n238405 );
nand ( n238407 , n238358 , n238396 );
nand ( n238408 , n238406 , n238407 );
buf ( n238409 , n238408 );
and ( n238410 , n238403 , n238409 );
nor ( n238411 , n238402 , n238410 );
not ( n238412 , n238411 );
not ( n238413 , n235682 );
not ( n238414 , n235627 );
nand ( n238415 , n235629 , n238414 );
not ( n238416 , n238415 );
not ( n238417 , n50987 );
not ( n238418 , n238417 );
and ( n238419 , n238416 , n238418 );
and ( n238420 , n238415 , n238417 );
nor ( n238421 , n238419 , n238420 );
not ( n238422 , n238421 );
not ( n238423 , n50984 );
or ( n238424 , n238422 , n238423 );
or ( n238425 , n50984 , n238421 );
nand ( n238426 , n238424 , n238425 );
nand ( n238427 , n235660 , n235647 );
and ( n238428 , n238427 , n228807 );
not ( n238429 , n238427 );
and ( n238430 , n238429 , n51045 );
nor ( n238431 , n238428 , n238430 );
and ( n238432 , n238426 , n238431 );
not ( n238433 , n238426 );
not ( n238434 , n238431 );
and ( n238435 , n238433 , n238434 );
nor ( n238436 , n238432 , n238435 );
not ( n238437 , n228877 );
not ( n238438 , n238437 );
not ( n238439 , n51131 );
not ( n238440 , n235670 );
nand ( n238441 , n238439 , n238440 );
not ( n238442 , n238441 );
or ( n238443 , n238438 , n238442 );
or ( n238444 , n238441 , n238437 );
nand ( n238445 , n238443 , n238444 );
not ( n238446 , n238445 );
not ( n238447 , n235703 );
and ( n238448 , n238447 , n51098 );
and ( n238449 , n238448 , n51087 );
not ( n238450 , n238448 );
and ( n238451 , n238450 , n51086 );
nor ( n238452 , n238449 , n238451 );
not ( n238453 , n238452 );
and ( n238454 , n238446 , n238453 );
and ( n238455 , n238445 , n238452 );
nor ( n238456 , n238454 , n238455 );
and ( n238457 , n238436 , n238456 );
not ( n238458 , n238436 );
not ( n238459 , n238456 );
and ( n238460 , n238458 , n238459 );
nor ( n238461 , n238457 , n238460 );
not ( n238462 , n238461 );
or ( n238463 , n238413 , n238462 );
not ( n238464 , n235682 );
not ( n238465 , n238456 );
not ( n238466 , n238436 );
or ( n238467 , n238465 , n238466 );
not ( n238468 , n238436 );
nand ( n238469 , n238468 , n238459 );
nand ( n238470 , n238467 , n238469 );
nand ( n238471 , n238464 , n238470 );
nand ( n238472 , n238463 , n238471 );
not ( n238473 , n32473 );
and ( n238474 , n238472 , n238473 );
not ( n238475 , n238472 );
buf ( n238476 , n32473 );
and ( n238477 , n238475 , n238476 );
nor ( n238478 , n238474 , n238477 );
nand ( n238479 , n238412 , n238478 );
not ( n238480 , n233138 );
nor ( n238481 , n238480 , n233967 );
not ( n238482 , n238481 );
not ( n238483 , n233138 );
nand ( n238484 , n238483 , n233967 );
nand ( n238485 , n238482 , n238484 );
not ( n238486 , n38657 );
not ( n238487 , n40860 );
not ( n238488 , n238487 );
not ( n238489 , n45944 );
or ( n238490 , n238488 , n238489 );
or ( n238491 , n45944 , n238487 );
nand ( n238492 , n238490 , n238491 );
not ( n238493 , n238492 );
or ( n238494 , n238486 , n238493 );
or ( n238495 , n38657 , n238492 );
nand ( n238496 , n238494 , n238495 );
not ( n238497 , n238496 );
not ( n238498 , n47494 );
xor ( n238499 , n33393 , n238498 );
xnor ( n238500 , n238499 , n38569 );
nand ( n238501 , n238497 , n238500 );
not ( n238502 , n238501 );
not ( n238503 , n235476 );
and ( n238504 , n238502 , n238503 );
and ( n238505 , n238501 , n235476 );
nor ( n238506 , n238504 , n238505 );
not ( n238507 , n238506 );
not ( n238508 , n235388 );
not ( n238509 , n27973 );
not ( n238510 , n204504 );
or ( n238511 , n238509 , n238510 );
not ( n238512 , n27973 );
nand ( n238513 , n238512 , n41319 );
nand ( n238514 , n238511 , n238513 );
and ( n238515 , n238514 , n41360 );
not ( n238516 , n238514 );
and ( n238517 , n238516 , n41361 );
nor ( n238518 , n238515 , n238517 );
not ( n238519 , n238518 );
nand ( n238520 , n238519 , n235399 );
not ( n238521 , n238520 );
or ( n238522 , n238508 , n238521 );
nand ( n238523 , n238519 , n235399 );
or ( n238524 , n235388 , n238523 );
nand ( n238525 , n238522 , n238524 );
not ( n238526 , n238525 );
not ( n238527 , n39383 );
not ( n238528 , n32524 );
or ( n238529 , n238527 , n238528 );
not ( n238530 , n39383 );
nand ( n238531 , n238530 , n30099 );
nand ( n238532 , n238529 , n238531 );
and ( n238533 , n238532 , n28721 );
not ( n238534 , n238532 );
and ( n238535 , n238534 , n28722 );
nor ( n238536 , n238533 , n238535 );
not ( n238537 , n238536 );
buf ( n238538 , RI173362b0_2177);
not ( n238539 , n238538 );
not ( n238540 , n35156 );
or ( n238541 , n238539 , n238540 );
nand ( n238542 , n51833 , n205413 );
nand ( n238543 , n238541 , n238542 );
not ( n238544 , n238543 );
not ( n238545 , n36751 );
and ( n238546 , n238544 , n238545 );
and ( n238547 , n238543 , n36751 );
nor ( n238548 , n238546 , n238547 );
nand ( n238549 , n238537 , n238548 );
not ( n238550 , n238549 );
not ( n238551 , n235454 );
and ( n238552 , n238550 , n238551 );
not ( n238553 , n238548 );
not ( n238554 , n238553 );
nand ( n238555 , n238554 , n238537 );
and ( n238556 , n238555 , n235454 );
nor ( n238557 , n238552 , n238556 );
not ( n238558 , n238557 );
or ( n238559 , n238526 , n238558 );
or ( n238560 , n238557 , n238525 );
nand ( n238561 , n238559 , n238560 );
not ( n238562 , n238561 );
and ( n238563 , n238507 , n238562 );
and ( n238564 , n238506 , n238561 );
nor ( n238565 , n238563 , n238564 );
not ( n238566 , n238565 );
not ( n238567 , n238566 );
buf ( n238568 , n34698 );
xor ( n238569 , n238568 , n40218 );
xnor ( n238570 , n238569 , n204892 );
not ( n238571 , n36168 );
not ( n238572 , n38408 );
not ( n238573 , n42091 );
or ( n238574 , n238572 , n238573 );
or ( n238575 , n42095 , n38408 );
nand ( n238576 , n238574 , n238575 );
not ( n238577 , n238576 );
and ( n238578 , n238571 , n238577 );
not ( n238579 , n41024 );
and ( n238580 , n238579 , n238576 );
nor ( n238581 , n238578 , n238580 );
not ( n238582 , n238581 );
nand ( n238583 , n238570 , n238582 );
not ( n238584 , n238583 );
not ( n238585 , n235545 );
and ( n238586 , n238584 , n238585 );
and ( n238587 , n238583 , n235545 );
nor ( n238588 , n238586 , n238587 );
not ( n238589 , n238588 );
not ( n238590 , n238589 );
xor ( n238591 , n26471 , n29815 );
xnor ( n238592 , n238591 , n36710 );
not ( n238593 , n28749 );
not ( n238594 , n205322 );
or ( n238595 , n238593 , n238594 );
or ( n238596 , n205322 , n28749 );
nand ( n238597 , n238595 , n238596 );
not ( n238598 , n45336 );
and ( n238599 , n238597 , n238598 );
not ( n238600 , n238597 );
and ( n238601 , n238600 , n45336 );
nor ( n238602 , n238599 , n238601 );
not ( n238603 , n238602 );
nand ( n238604 , n238592 , n238603 );
and ( n238605 , n238604 , n235528 );
not ( n238606 , n238604 );
and ( n238607 , n238606 , n235529 );
nor ( n238608 , n238605 , n238607 );
not ( n238609 , n238608 );
not ( n238610 , n238609 );
or ( n238611 , n238590 , n238610 );
nand ( n238612 , n238608 , n238588 );
nand ( n238613 , n238611 , n238612 );
not ( n238614 , n238613 );
not ( n238615 , n238614 );
or ( n238616 , n238567 , n238615 );
not ( n238617 , n238566 );
not ( n238618 , n238614 );
nand ( n238619 , n238617 , n238618 );
nand ( n238620 , n238616 , n238619 );
buf ( n238621 , n238620 );
and ( n238622 , n238485 , n238621 );
not ( n238623 , n238485 );
not ( n238624 , n238565 );
and ( n238625 , n238613 , n238624 );
not ( n238626 , n238613 );
and ( n238627 , n238626 , n238565 );
or ( n238628 , n238625 , n238627 );
buf ( n238629 , n238628 );
and ( n238630 , n238623 , n238629 );
nor ( n238631 , n238622 , n238630 );
not ( n238632 , n238631 );
nand ( n238633 , n238632 , n230207 );
or ( n238634 , n238479 , n238633 );
buf ( n238635 , n233971 );
nor ( n238636 , n238632 , n238635 );
nand ( n238637 , n238636 , n238479 );
buf ( n238638 , n35431 );
nand ( n238639 , n238638 , n25568 );
nand ( n238640 , n238634 , n238637 , n238639 );
buf ( n238641 , n238640 );
buf ( n238642 , n25760 );
not ( n238643 , n238642 );
not ( n238644 , n40006 );
or ( n238645 , n238643 , n238644 );
or ( n238646 , n40006 , n238642 );
nand ( n238647 , n238645 , n238646 );
not ( n238648 , n238647 );
not ( n238649 , n30607 );
or ( n238650 , n238648 , n238649 );
or ( n238651 , n30607 , n238647 );
nand ( n238652 , n238650 , n238651 );
nor ( n238653 , n238652 , n230150 );
not ( n238654 , n238653 );
not ( n238655 , n35077 );
not ( n238656 , n38088 );
or ( n238657 , n238655 , n238656 );
not ( n238658 , n35077 );
nand ( n238659 , n238658 , n39873 );
nand ( n238660 , n238657 , n238659 );
and ( n238661 , n238660 , n204676 );
not ( n238662 , n238660 );
not ( n238663 , n204671 );
and ( n238664 , n238662 , n238663 );
nor ( n238665 , n238661 , n238664 );
not ( n238666 , n238665 );
and ( n238667 , n238654 , n238666 );
and ( n238668 , n238653 , n238665 );
nor ( n238669 , n238667 , n238668 );
not ( n238670 , n238669 );
buf ( n238671 , n42755 );
not ( n238672 , n238671 );
not ( n238673 , n43340 );
or ( n238674 , n238672 , n238673 );
or ( n238675 , n43340 , n238671 );
nand ( n238676 , n238674 , n238675 );
xor ( n238677 , n238676 , n216493 );
nand ( n238678 , n52421 , n238677 );
not ( n238679 , n43240 );
not ( n238680 , n41856 );
or ( n238681 , n238679 , n238680 );
or ( n238682 , n46810 , n43240 );
nand ( n238683 , n238681 , n238682 );
and ( n238684 , n238683 , n217819 );
not ( n238685 , n238683 );
and ( n238686 , n238685 , n46816 );
nor ( n238687 , n238684 , n238686 );
and ( n238688 , n238678 , n238687 );
not ( n238689 , n238678 );
not ( n238690 , n238687 );
and ( n238691 , n238689 , n238690 );
nor ( n238692 , n238688 , n238691 );
not ( n238693 , n238692 );
or ( n238694 , n238670 , n238693 );
or ( n238695 , n238692 , n238669 );
nand ( n238696 , n238694 , n238695 );
not ( n238697 , n49922 );
buf ( n238698 , n204924 );
not ( n238699 , n238698 );
not ( n238700 , n33986 );
or ( n238701 , n238699 , n238700 );
or ( n238702 , n33986 , n238698 );
nand ( n238703 , n238701 , n238702 );
not ( n238704 , n238703 );
or ( n238705 , n238697 , n238704 );
or ( n238706 , n238703 , n49922 );
nand ( n238707 , n238705 , n238706 );
not ( n238708 , n238707 );
nand ( n238709 , n238708 , n52356 );
not ( n238710 , n238709 );
not ( n238711 , n40725 );
not ( n238712 , n32522 );
and ( n238713 , n238711 , n238712 );
and ( n238714 , n40725 , n32522 );
nor ( n238715 , n238713 , n238714 );
and ( n238716 , n238715 , n40734 );
not ( n238717 , n238715 );
not ( n238718 , n32962 );
and ( n238719 , n238717 , n238718 );
nor ( n238720 , n238716 , n238719 );
buf ( n238721 , n238720 );
not ( n238722 , n238721 );
and ( n238723 , n238710 , n238722 );
and ( n238724 , n238709 , n238721 );
nor ( n238725 , n238723 , n238724 );
and ( n238726 , n238696 , n238725 );
not ( n238727 , n238696 );
not ( n238728 , n238725 );
and ( n238729 , n238727 , n238728 );
nor ( n238730 , n238726 , n238729 );
not ( n238731 , n238730 );
not ( n238732 , n238731 );
not ( n238733 , n52281 );
buf ( n238734 , n36021 );
nor ( n238735 , n39250 , n238734 );
not ( n238736 , n238735 );
nand ( n238737 , n39250 , n238734 );
nand ( n238738 , n238736 , n238737 );
not ( n238739 , n238738 );
not ( n238740 , n44633 );
and ( n238741 , n238739 , n238740 );
and ( n238742 , n238738 , n44633 );
nor ( n238743 , n238741 , n238742 );
nand ( n238744 , n238733 , n238743 );
not ( n238745 , n238744 );
xor ( n238746 , n33633 , n32139 );
xnor ( n238747 , n238746 , n204259 );
not ( n238748 , n238747 );
or ( n238749 , n238745 , n238748 );
or ( n238750 , n238747 , n238744 );
nand ( n238751 , n238749 , n238750 );
not ( n238752 , n238751 );
not ( n238753 , n236459 );
and ( n238754 , n28662 , n28659 );
not ( n238755 , n28662 );
not ( n238756 , RI174a3ae8_938);
and ( n238757 , n238755 , n238756 );
nor ( n238758 , n238754 , n238757 );
nor ( n238759 , n30533 , n238758 );
not ( n238760 , n238759 );
nand ( n238761 , n30533 , n238758 );
nand ( n238762 , n238760 , n238761 );
not ( n238763 , n238762 );
or ( n238764 , n238753 , n238763 );
or ( n238765 , n238762 , n30543 );
nand ( n238766 , n238764 , n238765 );
not ( n238767 , n238766 );
nand ( n238768 , n238767 , n52307 );
not ( n238769 , n238768 );
not ( n238770 , n215681 );
not ( n238771 , n29213 );
or ( n238772 , n238770 , n238771 );
or ( n238773 , n206976 , n215681 );
nand ( n238774 , n238772 , n238773 );
not ( n238775 , n224643 );
and ( n238776 , n238774 , n238775 );
not ( n238777 , n238774 );
and ( n238778 , n238777 , n224643 );
nor ( n238779 , n238776 , n238778 );
not ( n238780 , n238779 );
and ( n238781 , n238769 , n238780 );
and ( n238782 , n238768 , n238779 );
nor ( n238783 , n238781 , n238782 );
not ( n238784 , n238783 );
or ( n238785 , n238752 , n238784 );
or ( n238786 , n238783 , n238751 );
nand ( n238787 , n238785 , n238786 );
not ( n238788 , n238787 );
not ( n238789 , n238788 );
or ( n238790 , n238732 , n238789 );
nand ( n238791 , n238787 , n238730 );
nand ( n238792 , n238790 , n238791 );
nand ( n238793 , n52272 , n52281 );
not ( n238794 , n238743 );
xor ( n238795 , n238793 , n238794 );
nor ( n238796 , n238792 , n238795 );
not ( n238797 , n238796 );
nand ( n238798 , n238795 , n238792 );
nand ( n238799 , n238797 , n238798 );
not ( n238800 , n238799 );
nand ( n238801 , n43372 , n236579 );
not ( n238802 , n41503 );
not ( n238803 , n53519 );
or ( n238804 , n238802 , n238803 );
or ( n238805 , n32279 , n41503 );
nand ( n238806 , n238804 , n238805 );
and ( n238807 , n238806 , n32323 );
not ( n238808 , n238806 );
and ( n238809 , n238808 , n32326 );
nor ( n238810 , n238807 , n238809 );
buf ( n238811 , n238810 );
xnor ( n238812 , n238801 , n238811 );
not ( n238813 , n238812 );
not ( n238814 , n238813 );
nand ( n238815 , n43296 , n43392 );
buf ( n238816 , n34176 );
not ( n238817 , n238816 );
not ( n238818 , n225371 );
or ( n238819 , n238817 , n238818 );
not ( n238820 , n238816 );
nand ( n238821 , n238820 , n47606 );
nand ( n238822 , n238819 , n238821 );
not ( n238823 , n238822 );
not ( n238824 , n204860 );
or ( n238825 , n238823 , n238824 );
or ( n238826 , n226349 , n238822 );
nand ( n238827 , n238825 , n238826 );
not ( n238828 , n238827 );
and ( n238829 , n238815 , n238828 );
not ( n238830 , n238815 );
and ( n238831 , n238830 , n238827 );
nor ( n238832 , n238829 , n238831 );
not ( n238833 , n238832 );
not ( n238834 , n238833 );
or ( n238835 , n238814 , n238834 );
nand ( n238836 , n238832 , n238812 );
nand ( n238837 , n238835 , n238836 );
nand ( n238838 , n236589 , n43329 );
not ( n238839 , n238838 );
buf ( n238840 , n37930 );
not ( n238841 , n238840 );
not ( n238842 , n29212 );
or ( n238843 , n238841 , n238842 );
or ( n238844 , n29214 , n238840 );
nand ( n238845 , n238843 , n238844 );
not ( n238846 , n238845 );
not ( n238847 , n224642 );
or ( n238848 , n238846 , n238847 );
or ( n238849 , n224643 , n238845 );
nand ( n238850 , n238848 , n238849 );
not ( n238851 , n238850 );
and ( n238852 , n238839 , n238851 );
and ( n238853 , n238838 , n238850 );
nor ( n238854 , n238852 , n238853 );
not ( n238855 , n238854 );
and ( n238856 , n238837 , n238855 );
not ( n238857 , n238837 );
and ( n238858 , n238857 , n238854 );
nor ( n238859 , n238856 , n238858 );
not ( n238860 , n236561 );
not ( n238861 , n43479 );
nand ( n238862 , n238861 , n43457 );
not ( n238863 , n238862 );
or ( n238864 , n238860 , n238863 );
or ( n238865 , n238862 , n236561 );
nand ( n238866 , n238864 , n238865 );
not ( n238867 , n238866 );
not ( n238868 , n221191 );
nand ( n238869 , n238868 , n43441 );
not ( n238870 , n28806 );
not ( n238871 , n34381 );
or ( n238872 , n238870 , n238871 );
or ( n238873 , n34381 , n28806 );
nand ( n238874 , n238872 , n238873 );
and ( n238875 , n238874 , n224001 );
not ( n238876 , n238874 );
and ( n238877 , n238876 , n225270 );
nor ( n238878 , n238875 , n238877 );
and ( n238879 , n238869 , n238878 );
not ( n238880 , n238869 );
not ( n238881 , n238878 );
and ( n238882 , n238880 , n238881 );
nor ( n238883 , n238879 , n238882 );
not ( n238884 , n238883 );
not ( n238885 , n238884 );
or ( n238886 , n238867 , n238885 );
not ( n238887 , n238866 );
nand ( n238888 , n238887 , n238883 );
nand ( n238889 , n238886 , n238888 );
not ( n238890 , n238889 );
and ( n238891 , n238859 , n238890 );
not ( n238892 , n238859 );
and ( n238893 , n238892 , n238889 );
nor ( n238894 , n238891 , n238893 );
buf ( n238895 , n238894 );
not ( n238896 , n238895 );
and ( n238897 , n238800 , n238896 );
and ( n238898 , n238799 , n238895 );
nor ( n238899 , n238897 , n238898 );
not ( n238900 , n205649 );
nor ( n238901 , n238899 , n238900 );
nand ( n238902 , n236526 , n236349 );
and ( n238903 , n238902 , n236528 );
not ( n238904 , n238902 );
not ( n238905 , n236528 );
and ( n238906 , n238904 , n238905 );
nor ( n238907 , n238903 , n238906 );
not ( n238908 , n238907 );
buf ( n238909 , n30630 );
not ( n238910 , n238909 );
not ( n238911 , n238910 );
not ( n238912 , n39922 );
or ( n238913 , n238911 , n238912 );
nand ( n238914 , n39921 , n238909 );
nand ( n238915 , n238913 , n238914 );
and ( n238916 , n238915 , n235930 );
not ( n238917 , n238915 );
and ( n238918 , n238917 , n47612 );
nor ( n238919 , n238916 , n238918 );
not ( n238920 , n238919 );
not ( n238921 , n51972 );
nand ( n238922 , n238920 , n238921 );
and ( n238923 , n238922 , n51962 );
not ( n238924 , n238922 );
and ( n238925 , n238924 , n236291 );
nor ( n238926 , n238923 , n238925 );
not ( n238927 , n238926 );
not ( n238928 , n238927 );
buf ( n238929 , n40522 );
not ( n238930 , n238929 );
not ( n238931 , n33657 );
or ( n238932 , n238930 , n238931 );
not ( n238933 , n238929 );
nand ( n238934 , n238933 , n34191 );
nand ( n238935 , n238932 , n238934 );
and ( n238936 , n238935 , n34220 );
not ( n238937 , n238935 );
and ( n238938 , n238937 , n34227 );
nor ( n238939 , n238936 , n238938 );
not ( n238940 , n51928 );
nand ( n238941 , n238939 , n238940 );
not ( n238942 , n238941 );
not ( n238943 , n236283 );
and ( n238944 , n238942 , n238943 );
and ( n238945 , n238941 , n236283 );
nor ( n238946 , n238944 , n238945 );
not ( n238947 , n238946 );
not ( n238948 , n238947 );
or ( n238949 , n238928 , n238948 );
nand ( n238950 , n238926 , n238946 );
nand ( n238951 , n238949 , n238950 );
xor ( n238952 , n51797 , n238951 );
not ( n238953 , n236534 );
not ( n238954 , n26407 );
not ( n238955 , n41054 );
or ( n238956 , n238954 , n238955 );
not ( n238957 , n26407 );
nand ( n238958 , n238957 , n45695 );
nand ( n238959 , n238956 , n238958 );
and ( n238960 , n238959 , n235697 );
not ( n238961 , n238959 );
and ( n238962 , n238961 , n44779 );
nor ( n238963 , n238960 , n238962 );
not ( n238964 , n51839 );
nand ( n238965 , n238963 , n238964 );
not ( n238966 , n238965 );
not ( n238967 , n236316 );
and ( n238968 , n238966 , n238967 );
and ( n238969 , n238965 , n236316 );
nor ( n238970 , n238968 , n238969 );
not ( n238971 , n238970 );
or ( n238972 , n238953 , n238971 );
or ( n238973 , n238970 , n236534 );
nand ( n238974 , n238972 , n238973 );
xnor ( n238975 , n238952 , n238974 );
not ( n238976 , n238975 );
or ( n238977 , n238908 , n238976 );
not ( n238978 , n238907 );
xor ( n238979 , n236533 , n238970 );
xor ( n238980 , n238979 , n51797 );
not ( n238981 , n238951 );
and ( n238982 , n238980 , n238981 );
not ( n238983 , n238980 );
and ( n238984 , n238983 , n238951 );
nor ( n238985 , n238982 , n238984 );
nand ( n238986 , n238978 , n238985 );
nand ( n238987 , n238977 , n238986 );
not ( n238988 , n45290 );
not ( n238989 , n214235 );
or ( n238990 , n238988 , n238989 );
or ( n238991 , n34603 , n45290 );
nand ( n238992 , n238990 , n238991 );
not ( n238993 , n238992 );
not ( n238994 , n30638 );
and ( n238995 , n238993 , n238994 );
and ( n238996 , n238992 , n44945 );
nor ( n238997 , n238995 , n238996 );
not ( n238998 , n238997 );
nand ( n238999 , n238998 , n52156 );
and ( n239000 , n238999 , n229906 );
not ( n239001 , n238999 );
and ( n239002 , n239001 , n236184 );
nor ( n239003 , n239000 , n239002 );
not ( n239004 , n239003 );
not ( n239005 , n239004 );
and ( n239006 , n28619 , n208303 );
not ( n239007 , n28619 );
and ( n239008 , n239007 , n30543 );
nor ( n239009 , n239006 , n239008 );
and ( n239010 , n239009 , n227018 );
not ( n239011 , n239009 );
and ( n239012 , n239011 , n33760 );
nor ( n239013 , n239010 , n239012 );
nand ( n239014 , n229938 , n239013 );
not ( n239015 , n239014 );
not ( n239016 , n236177 );
and ( n239017 , n239015 , n239016 );
and ( n239018 , n239014 , n236177 );
nor ( n239019 , n239017 , n239018 );
not ( n239020 , n239019 );
not ( n239021 , n239020 );
or ( n239022 , n239005 , n239021 );
nand ( n239023 , n239019 , n239003 );
nand ( n239024 , n239022 , n239023 );
not ( n239025 , n239024 );
not ( n239026 , n239025 );
not ( n239027 , n35065 );
not ( n239028 , n46633 );
or ( n239029 , n239027 , n239028 );
not ( n239030 , n35065 );
nand ( n239031 , n239030 , n39873 );
nand ( n239032 , n239029 , n239031 );
and ( n239033 , n239032 , n204672 );
not ( n239034 , n239032 );
and ( n239035 , n239034 , n204677 );
nor ( n239036 , n239033 , n239035 );
not ( n239037 , n239036 );
nand ( n239038 , n239037 , n52112 );
not ( n239039 , n239038 );
not ( n239040 , n229861 );
and ( n239041 , n239039 , n239040 );
and ( n239042 , n239038 , n229861 );
nor ( n239043 , n239041 , n239042 );
not ( n239044 , n52072 );
not ( n239045 , n40991 );
not ( n239046 , n41500 );
or ( n239047 , n239045 , n239046 );
or ( n239048 , n41500 , n40991 );
nand ( n239049 , n239047 , n239048 );
not ( n239050 , n239049 );
not ( n239051 , n41515 );
not ( n239052 , n239051 );
or ( n239053 , n239050 , n239052 );
or ( n239054 , n239051 , n239049 );
nand ( n239055 , n239053 , n239054 );
not ( n239056 , n239055 );
not ( n239057 , n38347 );
or ( n239058 , n239056 , n239057 );
or ( n239059 , n45320 , n239055 );
nand ( n239060 , n239058 , n239059 );
nand ( n239061 , n239044 , n239060 );
not ( n239062 , n239061 );
not ( n239063 , n236222 );
or ( n239064 , n239062 , n239063 );
or ( n239065 , n236222 , n239061 );
nand ( n239066 , n239064 , n239065 );
or ( n239067 , n239043 , n239066 );
nand ( n239068 , n239066 , n239043 );
nand ( n239069 , n239067 , n239068 );
not ( n239070 , n236255 );
not ( n239071 , n239070 );
not ( n239072 , n52028 );
not ( n239073 , n38709 );
not ( n239074 , n205333 );
not ( n239075 , n31832 );
not ( n239076 , n239075 );
or ( n239077 , n239074 , n239076 );
not ( n239078 , n205333 );
nand ( n239079 , n239078 , n31832 );
nand ( n239080 , n239077 , n239079 );
not ( n239081 , n239080 );
or ( n239082 , n239073 , n239081 );
or ( n239083 , n239080 , n38709 );
nand ( n239084 , n239082 , n239083 );
nand ( n239085 , n239072 , n239084 );
not ( n239086 , n239085 );
or ( n239087 , n239071 , n239086 );
or ( n239088 , n239085 , n239070 );
nand ( n239089 , n239087 , n239088 );
and ( n239090 , n239069 , n239089 );
not ( n239091 , n239069 );
not ( n239092 , n239089 );
and ( n239093 , n239091 , n239092 );
nor ( n239094 , n239090 , n239093 );
not ( n239095 , n239094 );
or ( n239096 , n239026 , n239095 );
not ( n239097 , n239094 );
nand ( n239098 , n239097 , n239024 );
nand ( n239099 , n239096 , n239098 );
buf ( n239100 , n239099 );
and ( n239101 , n238987 , n239100 );
not ( n239102 , n238987 );
not ( n239103 , n239097 );
not ( n239104 , n239024 );
and ( n239105 , n239103 , n239104 );
and ( n239106 , n239097 , n239024 );
nor ( n239107 , n239105 , n239106 );
buf ( n239108 , n239107 );
and ( n239109 , n239102 , n239108 );
nor ( n239110 , n239101 , n239109 );
not ( n239111 , n239110 );
not ( n239112 , n226363 );
not ( n239113 , n234420 );
or ( n239114 , n239112 , n239113 );
not ( n239115 , n226363 );
and ( n239116 , n234386 , n234418 );
not ( n239117 , n234386 );
and ( n239118 , n239117 , n234415 );
nor ( n239119 , n239116 , n239118 );
nand ( n239120 , n239115 , n239119 );
nand ( n239121 , n239114 , n239120 );
nand ( n239122 , n48150 , n226543 );
not ( n239123 , n239122 );
not ( n239124 , n30495 );
not ( n239125 , n28622 );
and ( n239126 , n239124 , n239125 );
not ( n239127 , n208303 );
and ( n239128 , n239127 , n28622 );
nor ( n239129 , n239126 , n239128 );
not ( n239130 , n227018 );
and ( n239131 , n239129 , n239130 );
not ( n239132 , n239129 );
and ( n239133 , n239132 , n33759 );
nor ( n239134 , n239131 , n239133 );
not ( n239135 , n239134 );
and ( n239136 , n239123 , n239135 );
and ( n239137 , n239122 , n239134 );
nor ( n239138 , n239136 , n239137 );
not ( n239139 , n239138 );
not ( n239140 , n239139 );
not ( n239141 , n48759 );
nand ( n239142 , n239141 , n48111 );
not ( n239143 , n222183 );
not ( n239144 , n37377 );
and ( n239145 , n239143 , n239144 );
and ( n239146 , n222183 , n37377 );
nor ( n239147 , n239145 , n239146 );
and ( n239148 , n239147 , n45468 );
not ( n239149 , n239147 );
and ( n239150 , n239149 , n236271 );
nor ( n239151 , n239148 , n239150 );
not ( n239152 , n239151 );
and ( n239153 , n239142 , n239152 );
not ( n239154 , n239142 );
and ( n239155 , n239154 , n239151 );
nor ( n239156 , n239153 , n239155 );
not ( n239157 , n239156 );
not ( n239158 , n239157 );
or ( n239159 , n239140 , n239158 );
nand ( n239160 , n239156 , n239138 );
nand ( n239161 , n239159 , n239160 );
nand ( n239162 , n48191 , n226464 );
not ( n239163 , n239162 );
not ( n239164 , n37988 );
not ( n239165 , n208398 );
or ( n239166 , n239164 , n239165 );
not ( n239167 , n37988 );
nand ( n239168 , n239167 , n30694 );
nand ( n239169 , n239166 , n239168 );
and ( n239170 , n239169 , n42802 );
not ( n239171 , n239169 );
and ( n239172 , n239171 , n34180 );
nor ( n239173 , n239170 , n239172 );
not ( n239174 , n239173 );
not ( n239175 , n239174 );
not ( n239176 , n239175 );
and ( n239177 , n239163 , n239176 );
and ( n239178 , n239162 , n239175 );
nor ( n239179 , n239177 , n239178 );
and ( n239180 , n239161 , n239179 );
not ( n239181 , n239161 );
not ( n239182 , n239179 );
and ( n239183 , n239181 , n239182 );
nor ( n239184 , n239180 , n239183 );
not ( n239185 , n239184 );
not ( n239186 , n226502 );
nand ( n239187 , n239186 , n48064 );
not ( n239188 , n239187 );
not ( n239189 , n42576 );
not ( n239190 , n34521 );
or ( n239191 , n239189 , n239190 );
or ( n239192 , n34521 , n42576 );
nand ( n239193 , n239191 , n239192 );
xnor ( n239194 , n239193 , n34558 );
not ( n239195 , n239194 );
not ( n239196 , n239195 );
and ( n239197 , n239188 , n239196 );
and ( n239198 , n239187 , n239195 );
nor ( n239199 , n239197 , n239198 );
nand ( n239200 , n48718 , n48199 );
not ( n239201 , n239200 );
not ( n239202 , n29791 );
not ( n239203 , n35584 );
or ( n239204 , n239202 , n239203 );
or ( n239205 , n53432 , n29791 );
nand ( n239206 , n239204 , n239205 );
nor ( n239207 , n239206 , n35940 );
not ( n239208 , n239207 );
nand ( n239209 , n239206 , n35940 );
nand ( n239210 , n239208 , n239209 );
not ( n239211 , n239210 );
and ( n239212 , n239201 , n239211 );
and ( n239213 , n239200 , n239210 );
nor ( n239214 , n239212 , n239213 );
xnor ( n239215 , n239199 , n239214 );
and ( n239216 , n239185 , n239215 );
not ( n239217 , n239185 );
not ( n239218 , n239215 );
and ( n239219 , n239217 , n239218 );
nor ( n239220 , n239216 , n239219 );
buf ( n239221 , n239220 );
and ( n239222 , n239121 , n239221 );
not ( n239223 , n239121 );
not ( n239224 , n239215 );
not ( n239225 , n239185 );
or ( n239226 , n239224 , n239225 );
nand ( n239227 , n239184 , n239218 );
nand ( n239228 , n239226 , n239227 );
buf ( n239229 , n239228 );
and ( n239230 , n239223 , n239229 );
nor ( n239231 , n239222 , n239230 );
nand ( n239232 , n238901 , n239111 , n239231 );
not ( n239233 , n238899 );
not ( n239234 , n239233 );
not ( n239235 , n239111 );
or ( n239236 , n239234 , n239235 );
buf ( n239237 , n226003 );
nor ( n239238 , n239231 , n239237 );
nand ( n239239 , n239236 , n239238 );
buf ( n239240 , n35431 );
nand ( n239241 , n239240 , n30017 );
nand ( n239242 , n239232 , n239239 , n239241 );
buf ( n239243 , n239242 );
not ( n239244 , n236972 );
nand ( n239245 , n234995 , n236966 );
and ( n239246 , n239245 , n55701 );
not ( n239247 , n239245 );
and ( n239248 , n239247 , n233463 );
nor ( n239249 , n239246 , n239248 );
not ( n239250 , n239249 );
not ( n239251 , n239250 );
not ( n239252 , n55666 );
nand ( n239253 , n236977 , n234976 );
not ( n239254 , n239253 );
or ( n239255 , n239252 , n239254 );
not ( n239256 , n234979 );
nand ( n239257 , n239256 , n236977 );
or ( n239258 , n239257 , n55666 );
nand ( n239259 , n239255 , n239258 );
not ( n239260 , n239259 );
or ( n239261 , n239251 , n239260 );
or ( n239262 , n239259 , n239250 );
nand ( n239263 , n239261 , n239262 );
not ( n239264 , n239263 );
nand ( n239265 , n234904 , n236899 );
not ( n239266 , n239265 );
not ( n239267 , n55543 );
and ( n239268 , n239266 , n239267 );
and ( n239269 , n239265 , n55543 );
nor ( n239270 , n239268 , n239269 );
not ( n239271 , n239270 );
nand ( n239272 , n234925 , n236919 );
and ( n239273 , n239272 , n55586 );
not ( n239274 , n239272 );
and ( n239275 , n239274 , n233348 );
nor ( n239276 , n239273 , n239275 );
not ( n239277 , n239276 );
or ( n239278 , n239271 , n239277 );
or ( n239279 , n239276 , n239270 );
nand ( n239280 , n239278 , n239279 );
nand ( n239281 , n236942 , n234954 );
not ( n239282 , n233376 );
and ( n239283 , n239281 , n239282 );
not ( n239284 , n239281 );
and ( n239285 , n239284 , n233376 );
nor ( n239286 , n239283 , n239285 );
not ( n239287 , n239286 );
and ( n239288 , n239280 , n239287 );
not ( n239289 , n239280 );
and ( n239290 , n239289 , n239286 );
nor ( n239291 , n239288 , n239290 );
not ( n239292 , n239291 );
or ( n239293 , n239264 , n239292 );
not ( n239294 , n239291 );
not ( n239295 , n239263 );
nand ( n239296 , n239294 , n239295 );
nand ( n239297 , n239293 , n239296 );
not ( n239298 , n239297 );
not ( n239299 , n239298 );
or ( n239300 , n239244 , n239299 );
not ( n239301 , n236972 );
nand ( n239302 , n239301 , n239297 );
nand ( n239303 , n239300 , n239302 );
nand ( n239304 , n41486 , n55233 );
not ( n239305 , n239304 );
not ( n239306 , n43234 );
not ( n239307 , n41856 );
or ( n239308 , n239306 , n239307 );
or ( n239309 , n41856 , n43234 );
nand ( n239310 , n239308 , n239309 );
and ( n239311 , n239310 , n46815 );
not ( n239312 , n239310 );
and ( n239313 , n239312 , n46816 );
nor ( n239314 , n239311 , n239313 );
not ( n239315 , n239314 );
not ( n239316 , n239315 );
and ( n239317 , n239305 , n239316 );
and ( n239318 , n239304 , n239315 );
nor ( n239319 , n239317 , n239318 );
nand ( n239320 , n41418 , n55250 );
not ( n239321 , n204259 );
not ( n239322 , n29935 );
not ( n239323 , n32909 );
or ( n239324 , n239322 , n239323 );
or ( n239325 , n32909 , n29935 );
nand ( n239326 , n239324 , n239325 );
not ( n239327 , n239326 );
and ( n239328 , n239321 , n239327 );
and ( n239329 , n204259 , n239326 );
nor ( n239330 , n239328 , n239329 );
and ( n239331 , n239320 , n239330 );
not ( n239332 , n239320 );
not ( n239333 , n239330 );
and ( n239334 , n239332 , n239333 );
nor ( n239335 , n239331 , n239334 );
and ( n239336 , n239319 , n239335 );
not ( n239337 , n239319 );
not ( n239338 , n239335 );
and ( n239339 , n239337 , n239338 );
nor ( n239340 , n239336 , n239339 );
not ( n239341 , n239340 );
nand ( n239342 , n41617 , n55189 );
not ( n239343 , n239342 );
not ( n239344 , n25562 );
not ( n239345 , n36663 );
or ( n239346 , n239344 , n239345 );
not ( n239347 , n25562 );
nand ( n239348 , n239347 , n36662 );
nand ( n239349 , n239346 , n239348 );
and ( n239350 , n239349 , n28780 );
not ( n239351 , n239349 );
and ( n239352 , n239351 , n28779 );
nor ( n239353 , n239350 , n239352 );
not ( n239354 , n239353 );
and ( n239355 , n239343 , n239354 );
and ( n239356 , n239342 , n239353 );
nor ( n239357 , n239355 , n239356 );
not ( n239358 , n239357 );
nand ( n239359 , n55171 , n219315 );
not ( n239360 , n32702 );
not ( n239361 , n43996 );
or ( n239362 , n239360 , n239361 );
or ( n239363 , n43996 , n32702 );
nand ( n239364 , n239362 , n239363 );
and ( n239365 , n239364 , n36377 );
not ( n239366 , n239364 );
and ( n239367 , n239366 , n35787 );
nor ( n239368 , n239365 , n239367 );
and ( n239369 , n239359 , n239368 );
not ( n239370 , n239359 );
not ( n239371 , n239368 );
and ( n239372 , n239370 , n239371 );
nor ( n239373 , n239369 , n239372 );
not ( n239374 , n239373 );
or ( n239375 , n239358 , n239374 );
or ( n239376 , n239373 , n239357 );
nand ( n239377 , n239375 , n239376 );
nand ( n239378 , n232972 , n41573 );
xor ( n239379 , n239378 , n41235 );
and ( n239380 , n239377 , n239379 );
not ( n239381 , n239377 );
not ( n239382 , n239379 );
and ( n239383 , n239381 , n239382 );
nor ( n239384 , n239380 , n239383 );
not ( n239385 , n239384 );
or ( n239386 , n239341 , n239385 );
not ( n239387 , n239384 );
not ( n239388 , n239340 );
nand ( n239389 , n239387 , n239388 );
nand ( n239390 , n239386 , n239389 );
buf ( n239391 , n239390 );
and ( n239392 , n239303 , n239391 );
not ( n239393 , n239303 );
buf ( n239394 , n239384 );
and ( n239395 , n239394 , n239340 );
not ( n239396 , n239394 );
and ( n239397 , n239396 , n239388 );
nor ( n239398 , n239395 , n239397 );
buf ( n239399 , n239398 );
and ( n239400 , n239393 , n239399 );
nor ( n239401 , n239392 , n239400 );
nor ( n239402 , n239401 , n47173 );
xor ( n239403 , n205100 , n51206 );
xnor ( n239404 , n239403 , n41415 );
not ( n239405 , n239404 );
xor ( n239406 , n25840 , n37580 );
xnor ( n239407 , n239406 , n38839 );
not ( n239408 , n239407 );
nand ( n239409 , n239405 , n239408 );
not ( n239410 , n239409 );
not ( n239411 , n48058 );
not ( n239412 , n28219 );
not ( n239413 , n36238 );
or ( n239414 , n239412 , n239413 );
or ( n239415 , n36238 , n28219 );
nand ( n239416 , n239414 , n239415 );
not ( n239417 , n239416 );
or ( n239418 , n239411 , n239417 );
or ( n239419 , n239416 , n232350 );
nand ( n239420 , n239418 , n239419 );
not ( n239421 , n239420 );
and ( n239422 , n239410 , n239421 );
and ( n239423 , n239409 , n239420 );
nor ( n239424 , n239422 , n239423 );
not ( n239425 , n239424 );
not ( n239426 , n28968 );
not ( n239427 , n30441 );
not ( n239428 , n239427 );
and ( n239429 , n239426 , n239428 );
and ( n239430 , n29015 , n239427 );
nor ( n239431 , n239429 , n239430 );
and ( n239432 , n239431 , n33003 );
not ( n239433 , n239431 );
and ( n239434 , n239433 , n33002 );
nor ( n239435 , n239432 , n239434 );
not ( n239436 , n239435 );
not ( n239437 , n239420 );
nand ( n239438 , n239437 , n239404 );
not ( n239439 , n239438 );
or ( n239440 , n239436 , n239439 );
not ( n239441 , n239420 );
nand ( n239442 , n239441 , n239404 );
or ( n239443 , n239442 , n239435 );
nand ( n239444 , n239440 , n239443 );
not ( n239445 , n239444 );
not ( n239446 , n215032 );
not ( n239447 , n32246 );
not ( n239448 , n41964 );
or ( n239449 , n239447 , n239448 );
or ( n239450 , n41964 , n32246 );
nand ( n239451 , n239449 , n239450 );
not ( n239452 , n239451 );
or ( n239453 , n239446 , n239452 );
or ( n239454 , n215032 , n239451 );
nand ( n239455 , n239453 , n239454 );
not ( n239456 , n239455 );
not ( n239457 , n39293 );
not ( n239458 , n47560 );
or ( n239459 , n239457 , n239458 );
not ( n239460 , n221779 );
nand ( n239461 , n239460 , n39298 );
nand ( n239462 , n239459 , n239461 );
and ( n239463 , n239462 , n205074 );
not ( n239464 , n239462 );
and ( n239465 , n239464 , n221787 );
nor ( n239466 , n239463 , n239465 );
nand ( n239467 , n239456 , n239466 );
not ( n239468 , n239467 );
buf ( n239469 , n42922 );
not ( n239470 , n239469 );
not ( n239471 , n45225 );
or ( n239472 , n239470 , n239471 );
or ( n239473 , n43262 , n239469 );
nand ( n239474 , n239472 , n239473 );
and ( n239475 , n239474 , n222994 );
not ( n239476 , n239474 );
not ( n239477 , n45230 );
and ( n239478 , n239476 , n239477 );
nor ( n239479 , n239475 , n239478 );
not ( n239480 , n239479 );
not ( n239481 , n239480 );
and ( n239482 , n239468 , n239481 );
and ( n239483 , n239467 , n239480 );
nor ( n239484 , n239482 , n239483 );
not ( n239485 , n239484 );
and ( n239486 , n239445 , n239485 );
and ( n239487 , n239444 , n239484 );
nor ( n239488 , n239486 , n239487 );
not ( n239489 , n239488 );
not ( n239490 , n29929 );
not ( n239491 , n32906 );
or ( n239492 , n239490 , n239491 );
not ( n239493 , n29929 );
nand ( n239494 , n239493 , n26475 );
nand ( n239495 , n239492 , n239494 );
and ( n239496 , n239495 , n204258 );
not ( n239497 , n239495 );
and ( n239498 , n239497 , n204259 );
nor ( n239499 , n239496 , n239498 );
not ( n239500 , n41736 );
not ( n239501 , n35275 );
or ( n239502 , n239500 , n239501 );
or ( n239503 , n35275 , n41736 );
nand ( n239504 , n239502 , n239503 );
xor ( n239505 , n239504 , n37820 );
nand ( n239506 , n239499 , n239505 );
not ( n239507 , n36813 );
buf ( n239508 , n36060 );
not ( n239509 , n239508 );
not ( n239510 , n36848 );
not ( n239511 , n239510 );
or ( n239512 , n239509 , n239511 );
not ( n239513 , n36848 );
or ( n239514 , n239513 , n239508 );
nand ( n239515 , n239512 , n239514 );
not ( n239516 , n239515 );
or ( n239517 , n239507 , n239516 );
or ( n239518 , n239515 , n36813 );
nand ( n239519 , n239517 , n239518 );
not ( n239520 , n239519 );
and ( n239521 , n239506 , n239520 );
not ( n239522 , n239506 );
and ( n239523 , n239522 , n239519 );
nor ( n239524 , n239521 , n239523 );
not ( n239525 , n239524 );
not ( n239526 , n239525 );
not ( n239527 , n26233 );
not ( n239528 , n42779 );
or ( n239529 , n239527 , n239528 );
or ( n239530 , n42779 , n26233 );
nand ( n239531 , n239529 , n239530 );
not ( n239532 , n43122 );
and ( n239533 , n239531 , n239532 );
not ( n239534 , n239531 );
and ( n239535 , n239534 , n43122 );
nor ( n239536 , n239533 , n239535 );
not ( n239537 , n34563 );
not ( n239538 , n42598 );
and ( n239539 , n239537 , n239538 );
and ( n239540 , n34563 , n42598 );
nor ( n239541 , n239539 , n239540 );
and ( n239542 , n239541 , n39411 );
not ( n239543 , n239541 );
and ( n239544 , n239543 , n51431 );
nor ( n239545 , n239542 , n239544 );
nand ( n239546 , n239536 , n239545 );
not ( n239547 , n239546 );
not ( n239548 , n204741 );
not ( n239549 , n42844 );
or ( n239550 , n239548 , n239549 );
not ( n239551 , n204741 );
nand ( n239552 , n239551 , n26370 );
nand ( n239553 , n239550 , n239552 );
and ( n239554 , n239553 , n234648 );
not ( n239555 , n239553 );
and ( n239556 , n239555 , n234773 );
nor ( n239557 , n239554 , n239556 );
buf ( n239558 , n239557 );
not ( n239559 , n239558 );
and ( n239560 , n239547 , n239559 );
not ( n239561 , n239545 );
not ( n239562 , n239561 );
nand ( n239563 , n239562 , n239536 );
and ( n239564 , n239563 , n239558 );
nor ( n239565 , n239560 , n239564 );
not ( n239566 , n239565 );
not ( n239567 , n239566 );
or ( n239568 , n239526 , n239567 );
nand ( n239569 , n239565 , n239524 );
nand ( n239570 , n239568 , n239569 );
xor ( n239571 , n28783 , n225270 );
xnor ( n239572 , n239571 , n34382 );
and ( n239573 , n31765 , n34303 );
not ( n239574 , n31765 );
and ( n239575 , n239574 , n34299 );
or ( n239576 , n239573 , n239575 );
not ( n239577 , n34263 );
buf ( n239578 , n239577 );
and ( n239579 , n239576 , n239578 );
not ( n239580 , n239576 );
and ( n239581 , n239580 , n34264 );
nor ( n239582 , n239579 , n239581 );
not ( n239583 , n239582 );
nand ( n239584 , n239572 , n239583 );
and ( n239585 , n31503 , n38689 );
not ( n239586 , n31503 );
and ( n239587 , n239586 , n37172 );
nor ( n239588 , n239585 , n239587 );
and ( n239589 , n239588 , n38795 );
not ( n239590 , n239588 );
and ( n239591 , n239590 , n37193 );
or ( n239592 , n239589 , n239591 );
and ( n239593 , n239584 , n239592 );
not ( n239594 , n239584 );
not ( n239595 , n239592 );
and ( n239596 , n239594 , n239595 );
nor ( n239597 , n239593 , n239596 );
and ( n239598 , n239570 , n239597 );
not ( n239599 , n239570 );
not ( n239600 , n239597 );
and ( n239601 , n239599 , n239600 );
nor ( n239602 , n239598 , n239601 );
not ( n239603 , n239602 );
and ( n239604 , n239489 , n239603 );
and ( n239605 , n239488 , n239602 );
nor ( n239606 , n239604 , n239605 );
not ( n239607 , n239606 );
not ( n239608 , n239607 );
or ( n239609 , n239425 , n239608 );
not ( n239610 , n239606 );
or ( n239611 , n239610 , n239424 );
nand ( n239612 , n239609 , n239611 );
not ( n239613 , n239612 );
not ( n239614 , n229255 );
nand ( n239615 , n36197 , n239614 );
not ( n239616 , n239615 );
not ( n239617 , n36249 );
and ( n239618 , n239616 , n239617 );
and ( n239619 , n239615 , n36249 );
nor ( n239620 , n239618 , n239619 );
not ( n239621 , n239620 );
not ( n239622 , n239621 );
not ( n239623 , n36259 );
not ( n239624 , n51525 );
nand ( n239625 , n239623 , n239624 );
and ( n239626 , n239625 , n36266 );
not ( n239627 , n239625 );
not ( n239628 , n36266 );
and ( n239629 , n239627 , n239628 );
nor ( n239630 , n239626 , n239629 );
not ( n239631 , n239630 );
not ( n239632 , n239631 );
or ( n239633 , n239622 , n239632 );
nand ( n239634 , n239630 , n239620 );
nand ( n239635 , n239633 , n239634 );
not ( n239636 , n35969 );
nand ( n239637 , n239636 , n51396 );
not ( n239638 , n239637 );
not ( n239639 , n35957 );
not ( n239640 , n239639 );
and ( n239641 , n239638 , n239640 );
and ( n239642 , n239637 , n239639 );
nor ( n239643 , n239641 , n239642 );
not ( n239644 , n239643 );
not ( n239645 , n35944 );
or ( n239646 , n239644 , n239645 );
or ( n239647 , n35944 , n239643 );
nand ( n239648 , n239646 , n239647 );
and ( n239649 , n239648 , n237743 );
not ( n239650 , n239648 );
and ( n239651 , n239650 , n237744 );
nor ( n239652 , n239649 , n239651 );
xor ( n239653 , n239635 , n239652 );
buf ( n239654 , n239653 );
not ( n239655 , n239654 );
and ( n239656 , n239613 , n239655 );
and ( n239657 , n239612 , n239654 );
nor ( n239658 , n239656 , n239657 );
not ( n239659 , n239658 );
nand ( n239660 , n236348 , n51875 );
and ( n239661 , n239660 , n236527 );
not ( n239662 , n239660 );
and ( n239663 , n239662 , n236526 );
nor ( n239664 , n239661 , n239663 );
not ( n239665 , n239664 );
not ( n239666 , n239665 );
not ( n239667 , n51781 );
not ( n239668 , n229532 );
nand ( n239669 , n236372 , n239668 );
not ( n239670 , n239669 );
or ( n239671 , n239667 , n239670 );
or ( n239672 , n239669 , n51781 );
nand ( n239673 , n239671 , n239672 );
not ( n239674 , n238939 );
nand ( n239675 , n239674 , n236281 );
and ( n239676 , n239675 , n238940 );
not ( n239677 , n239675 );
and ( n239678 , n239677 , n51928 );
nor ( n239679 , n239676 , n239678 );
not ( n239680 , n239679 );
not ( n239681 , n239680 );
nand ( n239682 , n238919 , n236304 );
and ( n239683 , n239682 , n51972 );
not ( n239684 , n239682 );
and ( n239685 , n239684 , n238921 );
nor ( n239686 , n239683 , n239685 );
not ( n239687 , n239686 );
not ( n239688 , n239687 );
or ( n239689 , n239681 , n239688 );
nand ( n239690 , n239686 , n239679 );
nand ( n239691 , n239689 , n239690 );
xor ( n239692 , n239673 , n239691 );
not ( n239693 , n238907 );
not ( n239694 , n239693 );
not ( n239695 , n238963 );
nand ( n239696 , n239695 , n236332 );
and ( n239697 , n239696 , n238964 );
not ( n239698 , n239696 );
and ( n239699 , n239698 , n51839 );
nor ( n239700 , n239697 , n239699 );
not ( n239701 , n239700 );
or ( n239702 , n239694 , n239701 );
or ( n239703 , n239700 , n239693 );
nand ( n239704 , n239702 , n239703 );
xnor ( n239705 , n239692 , n239704 );
not ( n239706 , n239705 );
or ( n239707 , n239666 , n239706 );
not ( n239708 , n239665 );
xor ( n239709 , n238907 , n239700 );
xnor ( n239710 , n239709 , n239673 );
not ( n239711 , n239691 );
and ( n239712 , n239710 , n239711 );
not ( n239713 , n239710 );
and ( n239714 , n239713 , n239691 );
nor ( n239715 , n239712 , n239714 );
nand ( n239716 , n239708 , n239715 );
nand ( n239717 , n239707 , n239716 );
not ( n239718 , n239084 );
nand ( n239719 , n239718 , n236252 );
and ( n239720 , n239719 , n52028 );
not ( n239721 , n239719 );
and ( n239722 , n239721 , n239072 );
nor ( n239723 , n239720 , n239722 );
not ( n239724 , n239723 );
not ( n239725 , n239724 );
not ( n239726 , n239060 );
nand ( n239727 , n239726 , n236233 );
not ( n239728 , n239727 );
not ( n239729 , n239044 );
not ( n239730 , n239729 );
and ( n239731 , n239728 , n239730 );
and ( n239732 , n239727 , n239729 );
nor ( n239733 , n239731 , n239732 );
not ( n239734 , n239733 );
not ( n239735 , n52113 );
nand ( n239736 , n236214 , n239036 );
not ( n239737 , n239736 );
or ( n239738 , n239735 , n239737 );
or ( n239739 , n239736 , n52113 );
nand ( n239740 , n239738 , n239739 );
not ( n239741 , n239740 );
or ( n239742 , n239734 , n239741 );
or ( n239743 , n239740 , n239733 );
nand ( n239744 , n239742 , n239743 );
not ( n239745 , n239744 );
not ( n239746 , n239745 );
or ( n239747 , n239725 , n239746 );
nand ( n239748 , n239744 , n239723 );
nand ( n239749 , n239747 , n239748 );
not ( n239750 , n229939 );
not ( n239751 , n239013 );
nand ( n239752 , n236176 , n239751 );
not ( n239753 , n239752 );
or ( n239754 , n239750 , n239753 );
not ( n239755 , n239013 );
nand ( n239756 , n239755 , n236176 );
or ( n239757 , n239756 , n229939 );
nand ( n239758 , n239754 , n239757 );
not ( n239759 , n239758 );
nand ( n239760 , n238997 , n236193 );
not ( n239761 , n239760 );
not ( n239762 , n52157 );
and ( n239763 , n239761 , n239762 );
and ( n239764 , n239760 , n52157 );
nor ( n239765 , n239763 , n239764 );
not ( n239766 , n239765 );
and ( n239767 , n239759 , n239766 );
and ( n239768 , n239758 , n239765 );
nor ( n239769 , n239767 , n239768 );
and ( n239770 , n239749 , n239769 );
not ( n239771 , n239749 );
not ( n239772 , n239769 );
and ( n239773 , n239771 , n239772 );
nor ( n239774 , n239770 , n239773 );
buf ( n239775 , n239774 );
not ( n239776 , n239775 );
and ( n239777 , n239717 , n239776 );
not ( n239778 , n239717 );
and ( n239779 , n239778 , n239775 );
nor ( n239780 , n239777 , n239779 );
not ( n239781 , n239780 );
nand ( n239782 , n239402 , n239659 , n239781 );
not ( n239783 , n239401 );
not ( n239784 , n239783 );
not ( n239785 , n239659 );
or ( n239786 , n239784 , n239785 );
nand ( n239787 , n239780 , n205649 );
not ( n239788 , n239787 );
nand ( n239789 , n239786 , n239788 );
nand ( n239790 , n31576 , n34145 );
nand ( n239791 , n239782 , n239789 , n239790 );
buf ( n239792 , n239791 );
not ( n239793 , RI1754b788_33);
or ( n239794 , n229127 , n239793 );
not ( n239795 , RI19aadb70_2470);
or ( n239796 , n226822 , n239795 );
nand ( n239797 , n239794 , n239796 );
buf ( n239798 , n239797 );
nand ( n239799 , n46052 , n46040 );
not ( n239800 , n239799 );
not ( n239801 , n46697 );
or ( n239802 , n239800 , n239801 );
or ( n239803 , n46697 , n239799 );
nand ( n239804 , n239802 , n239803 );
not ( n239805 , n239804 );
not ( n239806 , n46673 );
not ( n239807 , n239806 );
nand ( n239808 , n46658 , n223784 );
not ( n239809 , n239808 );
or ( n239810 , n239807 , n239809 );
not ( n239811 , n46022 );
nand ( n239812 , n239811 , n46658 );
or ( n239813 , n239812 , n239806 );
nand ( n239814 , n239810 , n239813 );
nand ( n239815 , n46696 , n46051 );
not ( n239816 , n239815 );
not ( n239817 , n46693 );
and ( n239818 , n239816 , n239817 );
and ( n239819 , n239815 , n46693 );
nor ( n239820 , n239818 , n239819 );
and ( n239821 , n239814 , n239820 );
not ( n239822 , n239814 );
not ( n239823 , n239820 );
and ( n239824 , n239822 , n239823 );
nor ( n239825 , n239821 , n239824 );
not ( n239826 , n239825 );
not ( n239827 , n45913 );
nand ( n239828 , n46541 , n239827 );
not ( n239829 , n239828 );
not ( n239830 , n46529 );
and ( n239831 , n239829 , n239830 );
nand ( n239832 , n46541 , n239827 );
and ( n239833 , n239832 , n46529 );
nor ( n239834 , n239831 , n239833 );
not ( n239835 , n239834 );
nand ( n239836 , n45984 , n46607 );
and ( n239837 , n239836 , n46598 );
not ( n239838 , n239836 );
not ( n239839 , n46598 );
and ( n239840 , n239838 , n239839 );
nor ( n239841 , n239837 , n239840 );
not ( n239842 , n239841 );
or ( n239843 , n239835 , n239842 );
or ( n239844 , n239841 , n239834 );
nand ( n239845 , n239843 , n239844 );
and ( n239846 , n239845 , n230006 );
not ( n239847 , n239845 );
and ( n239848 , n239847 , n230007 );
nor ( n239849 , n239846 , n239848 );
not ( n239850 , n239849 );
and ( n239851 , n239826 , n239850 );
and ( n239852 , n239825 , n239849 );
nor ( n239853 , n239851 , n239852 );
not ( n239854 , n239853 );
not ( n239855 , n239854 );
not ( n239856 , n239855 );
or ( n239857 , n239805 , n239856 );
buf ( n239858 , n239853 );
or ( n239859 , n239858 , n239804 );
nand ( n239860 , n239857 , n239859 );
not ( n239861 , n52273 );
not ( n239862 , n239861 );
not ( n239863 , n52262 );
nand ( n239864 , n239863 , n238747 );
not ( n239865 , n239864 );
or ( n239866 , n239862 , n239865 );
not ( n239867 , n52262 );
nand ( n239868 , n239867 , n238747 );
or ( n239869 , n239868 , n239861 );
nand ( n239870 , n239866 , n239869 );
not ( n239871 , n239870 );
not ( n239872 , n230064 );
nand ( n239873 , n239872 , n238779 );
not ( n239874 , n239873 );
not ( n239875 , n52294 );
not ( n239876 , n239875 );
and ( n239877 , n239874 , n239876 );
and ( n239878 , n239873 , n239875 );
nor ( n239879 , n239877 , n239878 );
not ( n239880 , n239879 );
and ( n239881 , n239871 , n239880 );
and ( n239882 , n239870 , n239879 );
nor ( n239883 , n239881 , n239882 );
not ( n239884 , n239883 );
not ( n239885 , n239884 );
not ( n239886 , n52371 );
not ( n239887 , n239886 );
not ( n239888 , n52378 );
not ( n239889 , n238665 );
nand ( n239890 , n239888 , n239889 );
not ( n239891 , n239890 );
or ( n239892 , n239887 , n239891 );
or ( n239893 , n239890 , n239886 );
nand ( n239894 , n239892 , n239893 );
not ( n239895 , n239894 );
nand ( n239896 , n230103 , n238720 );
not ( n239897 , n239896 );
buf ( n239898 , n230088 );
not ( n239899 , n239898 );
and ( n239900 , n239897 , n239899 );
and ( n239901 , n239896 , n239898 );
nor ( n239902 , n239900 , n239901 );
not ( n239903 , n239902 );
or ( n239904 , n239895 , n239903 );
or ( n239905 , n239902 , n239894 );
nand ( n239906 , n239904 , n239905 );
not ( n239907 , n52397 );
nand ( n239908 , n239907 , n238690 );
and ( n239909 , n239908 , n230168 );
not ( n239910 , n239908 );
and ( n239911 , n239910 , n230167 );
nor ( n239912 , n239909 , n239911 );
and ( n239913 , n239906 , n239912 );
not ( n239914 , n239906 );
not ( n239915 , n239912 );
and ( n239916 , n239914 , n239915 );
nor ( n239917 , n239913 , n239916 );
not ( n239918 , n239917 );
not ( n239919 , n239918 );
or ( n239920 , n239885 , n239919 );
nand ( n239921 , n239917 , n239883 );
nand ( n239922 , n239920 , n239921 );
not ( n239923 , n239922 );
not ( n239924 , n239923 );
and ( n239925 , n239860 , n239924 );
not ( n239926 , n239860 );
and ( n239927 , n239917 , n239883 );
not ( n239928 , n239917 );
and ( n239929 , n239928 , n239884 );
nor ( n239930 , n239927 , n239929 );
buf ( n239931 , n239930 );
and ( n239932 , n239926 , n239931 );
nor ( n239933 , n239925 , n239932 );
not ( n239934 , n226003 );
nand ( n239935 , n239933 , n239934 );
not ( n239936 , n55978 );
nand ( n239937 , n223397 , n45611 );
not ( n239938 , n239937 );
and ( n239939 , n239936 , n239938 );
and ( n239940 , n55978 , n239937 );
nor ( n239941 , n239939 , n239940 );
not ( n239942 , n239941 );
not ( n239943 , n55992 );
nand ( n239944 , n239943 , n223437 );
xor ( n239945 , n239944 , n233763 );
not ( n239946 , n239945 );
not ( n239947 , n239946 );
not ( n239948 , n56020 );
nand ( n239949 , n239948 , n45711 );
not ( n239950 , n239949 );
not ( n239951 , n233786 );
and ( n239952 , n239950 , n239951 );
and ( n239953 , n239949 , n233786 );
nor ( n239954 , n239952 , n239953 );
not ( n239955 , n239954 );
not ( n239956 , n239955 );
or ( n239957 , n239947 , n239956 );
nand ( n239958 , n239954 , n239945 );
nand ( n239959 , n239957 , n239958 );
nand ( n239960 , n55952 , n45545 );
not ( n239961 , n239960 );
not ( n239962 , n238159 );
and ( n239963 , n239961 , n239962 );
and ( n239964 , n239960 , n238159 );
nor ( n239965 , n239963 , n239964 );
not ( n239966 , n239965 );
not ( n239967 , n233686 );
nand ( n239968 , n239967 , n45593 );
not ( n239969 , n238166 );
and ( n239970 , n239968 , n239969 );
not ( n239971 , n239968 );
and ( n239972 , n239971 , n238166 );
nor ( n239973 , n239970 , n239972 );
not ( n239974 , n239973 );
or ( n239975 , n239966 , n239974 );
or ( n239976 , n239973 , n239965 );
nand ( n239977 , n239975 , n239976 );
not ( n239978 , n55978 );
nand ( n239979 , n239978 , n45637 );
not ( n239980 , n239979 );
not ( n239981 , n233736 );
and ( n239982 , n239980 , n239981 );
and ( n239983 , n239979 , n233736 );
nor ( n239984 , n239982 , n239983 );
and ( n239985 , n239977 , n239984 );
not ( n239986 , n239977 );
not ( n239987 , n239984 );
and ( n239988 , n239986 , n239987 );
nor ( n239989 , n239985 , n239988 );
not ( n239990 , n239989 );
and ( n239991 , n239959 , n239990 );
not ( n239992 , n239959 );
and ( n239993 , n239992 , n239989 );
nor ( n239994 , n239991 , n239993 );
not ( n239995 , n239994 );
or ( n239996 , n239942 , n239995 );
not ( n239997 , n239941 );
and ( n239998 , n239959 , n239989 );
not ( n239999 , n239959 );
and ( n240000 , n239999 , n239990 );
nor ( n240001 , n239998 , n240000 );
nand ( n240002 , n239997 , n240001 );
nand ( n240003 , n239996 , n240002 );
nand ( n240004 , n230301 , n52468 );
and ( n240005 , n240004 , n40080 );
not ( n240006 , n240004 );
and ( n240007 , n240006 , n235752 );
nor ( n240008 , n240005 , n240007 );
not ( n240009 , n240008 );
not ( n240010 , n240009 );
not ( n240011 , n39933 );
nand ( n240012 , n240011 , n52492 );
not ( n240013 , n240012 );
not ( n240014 , n235743 );
and ( n240015 , n240013 , n240014 );
and ( n240016 , n240012 , n235743 );
nor ( n240017 , n240015 , n240016 );
not ( n240018 , n240017 );
not ( n240019 , n240018 );
or ( n240020 , n240010 , n240019 );
nand ( n240021 , n240008 , n240017 );
nand ( n240022 , n240020 , n240021 );
not ( n240023 , n52514 );
nand ( n240024 , n40137 , n240023 );
and ( n240025 , n240024 , n235765 );
not ( n240026 , n240024 );
and ( n240027 , n240026 , n217935 );
nor ( n240028 , n240025 , n240027 );
and ( n240029 , n240022 , n240028 );
not ( n240030 , n240022 );
not ( n240031 , n240028 );
and ( n240032 , n240030 , n240031 );
nor ( n240033 , n240029 , n240032 );
not ( n240034 , n240033 );
not ( n240035 , n240034 );
not ( n240036 , n39858 );
nand ( n240037 , n240036 , n52589 );
not ( n240038 , n240037 );
not ( n240039 , n235792 );
or ( n240040 , n240038 , n240039 );
or ( n240041 , n235792 , n240037 );
nand ( n240042 , n240040 , n240041 );
not ( n240043 , n240042 );
not ( n240044 , n39822 );
or ( n240045 , n240043 , n240044 );
or ( n240046 , n39822 , n240042 );
nand ( n240047 , n240045 , n240046 );
not ( n240048 , n240047 );
not ( n240049 , n240048 );
or ( n240050 , n240035 , n240049 );
nand ( n240051 , n240033 , n240047 );
nand ( n240052 , n240050 , n240051 );
not ( n240053 , n240052 );
and ( n240054 , n240003 , n240053 );
not ( n240055 , n240003 );
buf ( n240056 , n240052 );
buf ( n240057 , n240056 );
and ( n240058 , n240055 , n240057 );
nor ( n240059 , n240054 , n240058 );
nand ( n240060 , n45051 , n45038 );
not ( n240061 , n240060 );
not ( n240062 , n54890 );
and ( n240063 , n240061 , n240062 );
and ( n240064 , n240060 , n54890 );
nor ( n240065 , n240063 , n240064 );
not ( n240066 , n240065 );
not ( n240067 , n240066 );
not ( n240068 , n54917 );
or ( n240069 , n240067 , n240068 );
not ( n240070 , n240066 );
nand ( n240071 , n240070 , n54926 );
nand ( n240072 , n240069 , n240071 );
not ( n240073 , n55068 );
and ( n240074 , n240072 , n240073 );
not ( n240075 , n240072 );
and ( n240076 , n240075 , n55068 );
nor ( n240077 , n240074 , n240076 );
nor ( n240078 , n240059 , n240077 );
or ( n240079 , n239935 , n240078 );
not ( n240080 , n226010 );
nor ( n240081 , n239933 , n240080 );
nand ( n240082 , n240081 , n240078 );
nand ( n240083 , n39766 , n53981 );
nand ( n240084 , n240079 , n240082 , n240083 );
buf ( n240085 , n240084 );
buf ( n240086 , n239179 );
not ( n240087 , n240086 );
nand ( n240088 , n226502 , n239194 );
not ( n240089 , n240088 );
buf ( n240090 , n48049 );
not ( n240091 , n240090 );
and ( n240092 , n240089 , n240091 );
and ( n240093 , n240088 , n240090 );
nor ( n240094 , n240092 , n240093 );
not ( n240095 , n240094 );
nand ( n240096 , n48759 , n239152 );
buf ( n240097 , n48076 );
xor ( n240098 , n240096 , n240097 );
not ( n240099 , n240098 );
or ( n240100 , n240095 , n240099 );
or ( n240101 , n240094 , n240098 );
nand ( n240102 , n240100 , n240101 );
not ( n240103 , n239134 );
nand ( n240104 , n240103 , n226544 );
not ( n240105 , n225888 );
and ( n240106 , n240104 , n240105 );
not ( n240107 , n240104 );
and ( n240108 , n240107 , n225888 );
nor ( n240109 , n240106 , n240108 );
and ( n240110 , n240102 , n240109 );
not ( n240111 , n240102 );
not ( n240112 , n240109 );
and ( n240113 , n240111 , n240112 );
nor ( n240114 , n240110 , n240113 );
not ( n240115 , n48217 );
not ( n240116 , n240115 );
not ( n240117 , n239210 );
nand ( n240118 , n240117 , n48719 );
not ( n240119 , n240118 );
or ( n240120 , n240116 , n240119 );
not ( n240121 , n239210 );
nand ( n240122 , n240121 , n48719 );
or ( n240123 , n240122 , n240115 );
nand ( n240124 , n240120 , n240123 );
not ( n240125 , n240124 );
nand ( n240126 , n239174 , n226463 );
not ( n240127 , n240126 );
buf ( n240128 , n48184 );
not ( n240129 , n240128 );
and ( n240130 , n240127 , n240129 );
and ( n240131 , n240126 , n240128 );
nor ( n240132 , n240130 , n240131 );
not ( n240133 , n240132 );
and ( n240134 , n240125 , n240133 );
and ( n240135 , n240124 , n240132 );
nor ( n240136 , n240134 , n240135 );
and ( n240137 , n240114 , n240136 );
not ( n240138 , n240114 );
not ( n240139 , n240136 );
and ( n240140 , n240138 , n240139 );
or ( n240141 , n240137 , n240140 );
not ( n240142 , n240141 );
or ( n240143 , n240087 , n240142 );
and ( n240144 , n240114 , n240136 );
not ( n240145 , n240114 );
and ( n240146 , n240145 , n240139 );
nor ( n240147 , n240144 , n240146 );
not ( n240148 , n240147 );
or ( n240149 , n240148 , n240086 );
nand ( n240150 , n240143 , n240149 );
not ( n240151 , n240150 );
not ( n240152 , n227174 );
not ( n240153 , n240152 );
not ( n240154 , n240153 );
and ( n240155 , n240151 , n240154 );
and ( n240156 , n240150 , n240153 );
nor ( n240157 , n240155 , n240156 );
nand ( n240158 , n240157 , n222532 );
not ( n240159 , n49573 );
buf ( n240160 , n204934 );
xor ( n240161 , n240160 , n49922 );
xnor ( n240162 , n240161 , n34004 );
nand ( n240163 , n240159 , n240162 );
and ( n240164 , n30161 , n30158 );
not ( n240165 , n30161 );
buf ( n240166 , RI1749b7a8_978);
and ( n240167 , n240165 , n240166 );
nor ( n240168 , n240164 , n240167 );
not ( n240169 , n240168 );
not ( n240170 , n41360 );
or ( n240171 , n240169 , n240170 );
not ( n240172 , n240168 );
nand ( n240173 , n240172 , n47262 );
nand ( n240174 , n240171 , n240173 );
and ( n240175 , n240174 , n52705 );
not ( n240176 , n240174 );
and ( n240177 , n240176 , n27716 );
nor ( n240178 , n240175 , n240177 );
not ( n240179 , n240178 );
and ( n240180 , n240163 , n240179 );
not ( n240181 , n240163 );
and ( n240182 , n240181 , n240178 );
nor ( n240183 , n240180 , n240182 );
not ( n240184 , n240183 );
not ( n240185 , n224642 );
not ( n240186 , n37939 );
not ( n240187 , n29213 );
or ( n240188 , n240186 , n240187 );
not ( n240189 , n37939 );
nand ( n240190 , n240189 , n29212 );
nand ( n240191 , n240188 , n240190 );
not ( n240192 , n240191 );
and ( n240193 , n240185 , n240192 );
and ( n240194 , n224642 , n240191 );
nor ( n240195 , n240193 , n240194 );
not ( n240196 , n40773 );
not ( n240197 , n41252 );
not ( n240198 , n33443 );
or ( n240199 , n240197 , n240198 );
not ( n240200 , n41252 );
not ( n240201 , n33443 );
nand ( n240202 , n240200 , n240201 );
nand ( n240203 , n240199 , n240202 );
not ( n240204 , n240203 );
or ( n240205 , n240196 , n240204 );
or ( n240206 , n240203 , n33474 );
nand ( n240207 , n240205 , n240206 );
nand ( n240208 , n240195 , n240207 );
not ( n240209 , n240208 );
not ( n240210 , n227203 );
and ( n240211 , n240209 , n240210 );
and ( n240212 , n240208 , n227203 );
nor ( n240213 , n240211 , n240212 );
buf ( n240214 , n36510 );
not ( n240215 , n240214 );
not ( n240216 , n40224 );
or ( n240217 , n240215 , n240216 );
not ( n240218 , n240214 );
nand ( n240219 , n240218 , n26204 );
nand ( n240220 , n240217 , n240219 );
not ( n240221 , n240220 );
not ( n240222 , n30534 );
and ( n240223 , n240221 , n240222 );
and ( n240224 , n240220 , n40231 );
nor ( n240225 , n240223 , n240224 );
not ( n240226 , n42207 );
buf ( n240227 , n40561 );
not ( n240228 , n240227 );
not ( n240229 , n34225 );
or ( n240230 , n240228 , n240229 );
not ( n240231 , n240227 );
nand ( n240232 , n240231 , n34218 );
nand ( n240233 , n240230 , n240232 );
not ( n240234 , n240233 );
not ( n240235 , n240234 );
or ( n240236 , n240226 , n240235 );
not ( n240237 , n42207 );
nand ( n240238 , n240237 , n240233 );
nand ( n240239 , n240236 , n240238 );
nand ( n240240 , n240225 , n240239 );
not ( n240241 , n240240 );
not ( n240242 , n49515 );
and ( n240243 , n240241 , n240242 );
and ( n240244 , n240240 , n49515 );
nor ( n240245 , n240243 , n240244 );
xor ( n240246 , n240213 , n240245 );
buf ( n240247 , n30484 );
not ( n240248 , n240247 );
not ( n240249 , n41449 );
or ( n240250 , n240248 , n240249 );
not ( n240251 , n240247 );
nand ( n240252 , n240251 , n41448 );
nand ( n240253 , n240250 , n240252 );
and ( n240254 , n240253 , n33229 );
not ( n240255 , n240253 );
and ( n240256 , n240255 , n33230 );
nor ( n240257 , n240254 , n240256 );
not ( n240258 , n240257 );
not ( n240259 , n31062 );
not ( n240260 , n52884 );
or ( n240261 , n240259 , n240260 );
or ( n240262 , n52884 , n31062 );
nand ( n240263 , n240261 , n240262 );
xor ( n240264 , n240263 , n223614 );
not ( n240265 , n240264 );
nand ( n240266 , n240258 , n240265 );
and ( n240267 , n240266 , n49478 );
not ( n240268 , n240266 );
and ( n240269 , n240268 , n227240 );
nor ( n240270 , n240267 , n240269 );
xnor ( n240271 , n240246 , n240270 );
buf ( n240272 , n33223 );
not ( n240273 , n240272 );
not ( n240274 , n25772 );
or ( n240275 , n240273 , n240274 );
or ( n240276 , n34328 , n240272 );
nand ( n240277 , n240275 , n240276 );
and ( n240278 , n240277 , n44352 );
not ( n240279 , n240277 );
and ( n240280 , n240279 , n44348 );
nor ( n240281 , n240278 , n240280 );
not ( n240282 , n240281 );
not ( n240283 , n30219 );
not ( n240284 , n37123 );
or ( n240285 , n240283 , n240284 );
not ( n240286 , n30219 );
nand ( n240287 , n240286 , n37128 );
nand ( n240288 , n240285 , n240287 );
and ( n240289 , n240288 , n44334 );
not ( n240290 , n240288 );
and ( n240291 , n240290 , n44338 );
nor ( n240292 , n240289 , n240291 );
not ( n240293 , n240292 );
nand ( n240294 , n240282 , n240293 );
not ( n240295 , n240294 );
not ( n240296 , n49590 );
and ( n240297 , n240295 , n240296 );
and ( n240298 , n240294 , n49590 );
nor ( n240299 , n240297 , n240298 );
not ( n240300 , n240299 );
not ( n240301 , n240162 );
nand ( n240302 , n240301 , n240179 );
and ( n240303 , n240302 , n49559 );
not ( n240304 , n240302 );
and ( n240305 , n240304 , n49560 );
nor ( n240306 , n240303 , n240305 );
not ( n240307 , n240306 );
or ( n240308 , n240300 , n240307 );
or ( n240309 , n240306 , n240299 );
nand ( n240310 , n240308 , n240309 );
xor ( n240311 , n240271 , n240310 );
buf ( n240312 , n240311 );
not ( n240313 , n240312 );
or ( n240314 , n240184 , n240313 );
not ( n240315 , n240183 );
not ( n240316 , n240311 );
nand ( n240317 , n240315 , n240316 );
nand ( n240318 , n240314 , n240317 );
not ( n240319 , n204608 );
not ( n240320 , n30137 );
or ( n240321 , n240319 , n240320 );
not ( n240322 , n204608 );
nand ( n240323 , n240322 , n43577 );
nand ( n240324 , n240321 , n240323 );
and ( n240325 , n240324 , n33954 );
not ( n240326 , n240324 );
and ( n240327 , n240326 , n33957 );
nor ( n240328 , n240325 , n240327 );
not ( n240329 , n240328 );
not ( n240330 , n37036 );
not ( n240331 , n46993 );
or ( n240332 , n240330 , n240331 );
or ( n240333 , n46993 , n37036 );
nand ( n240334 , n240332 , n240333 );
and ( n240335 , n240334 , n221462 );
not ( n240336 , n240334 );
and ( n240337 , n240336 , n29371 );
nor ( n240338 , n240335 , n240337 );
not ( n240339 , n36321 );
not ( n240340 , n31053 );
or ( n240341 , n240339 , n240340 );
nand ( n240342 , n31052 , n36317 );
nand ( n240343 , n240341 , n240342 );
not ( n240344 , n240343 );
not ( n240345 , n31075 );
or ( n240346 , n240344 , n240345 );
or ( n240347 , n31075 , n240343 );
nand ( n240348 , n240346 , n240347 );
and ( n240349 , n240348 , n41894 );
not ( n240350 , n240348 );
and ( n240351 , n240350 , n39798 );
nor ( n240352 , n240349 , n240351 );
not ( n240353 , n240352 );
nand ( n240354 , n240338 , n240353 );
not ( n240355 , n240354 );
or ( n240356 , n240329 , n240355 );
not ( n240357 , n240352 );
nand ( n240358 , n240357 , n240338 );
or ( n240359 , n240358 , n240328 );
nand ( n240360 , n240356 , n240359 );
not ( n240361 , n240360 );
not ( n240362 , n30415 );
not ( n240363 , n28969 );
or ( n240364 , n240362 , n240363 );
or ( n240365 , n28969 , n30415 );
nand ( n240366 , n240364 , n240365 );
and ( n240367 , n240366 , n39532 );
not ( n240368 , n240366 );
and ( n240369 , n240368 , n33002 );
nor ( n240370 , n240367 , n240369 );
not ( n240371 , n28108 );
not ( n240372 , n37222 );
or ( n240373 , n240371 , n240372 );
or ( n240374 , n37222 , n28108 );
nand ( n240375 , n240373 , n240374 );
and ( n240376 , n240375 , n28680 );
not ( n240377 , n240375 );
and ( n240378 , n240377 , n28677 );
nor ( n240379 , n240376 , n240378 );
not ( n240380 , n240379 );
nand ( n240381 , n240370 , n240380 );
not ( n240382 , n240381 );
not ( n240383 , n29409 );
not ( n240384 , n32356 );
and ( n240385 , n240383 , n240384 );
and ( n240386 , n29415 , n32356 );
nor ( n240387 , n240385 , n240386 );
xor ( n240388 , n240387 , n207216 );
buf ( n240389 , n240388 );
not ( n240390 , n240389 );
and ( n240391 , n240382 , n240390 );
and ( n240392 , n240381 , n240389 );
nor ( n240393 , n240391 , n240392 );
not ( n240394 , n240393 );
or ( n240395 , n240361 , n240394 );
or ( n240396 , n240393 , n240360 );
nand ( n240397 , n240395 , n240396 );
xor ( n240398 , n36205 , n222628 );
xnor ( n240399 , n240398 , n29991 );
not ( n240400 , n217056 );
not ( n240401 , n205033 );
or ( n240402 , n240400 , n240401 );
not ( n240403 , n217056 );
nand ( n240404 , n240403 , n205029 );
nand ( n240405 , n240402 , n240404 );
and ( n240406 , n240405 , n205074 );
not ( n240407 , n240405 );
and ( n240408 , n240407 , n205068 );
nor ( n240409 , n240406 , n240408 );
not ( n240410 , n240409 );
nand ( n240411 , n240399 , n240410 );
not ( n240412 , n240411 );
not ( n240413 , n32173 );
not ( n240414 , n33613 );
or ( n240415 , n240413 , n240414 );
not ( n240416 , n32173 );
nand ( n240417 , n240416 , n33618 );
nand ( n240418 , n240415 , n240417 );
not ( n240419 , n240418 );
not ( n240420 , n43787 );
and ( n240421 , n240419 , n240420 );
and ( n240422 , n240418 , n43787 );
nor ( n240423 , n240421 , n240422 );
not ( n240424 , n240423 );
not ( n240425 , n240424 );
and ( n240426 , n240412 , n240425 );
and ( n240427 , n240411 , n240424 );
nor ( n240428 , n240426 , n240427 );
and ( n240429 , n240397 , n240428 );
not ( n240430 , n240397 );
not ( n240431 , n240428 );
and ( n240432 , n240430 , n240431 );
nor ( n240433 , n240429 , n240432 );
not ( n240434 , n240433 );
buf ( n240435 , n25580 );
not ( n240436 , n240435 );
not ( n240437 , n224022 );
or ( n240438 , n240436 , n240437 );
not ( n240439 , n240435 );
nand ( n240440 , n240439 , n219538 );
nand ( n240441 , n240438 , n240440 );
and ( n240442 , n240441 , n44683 );
not ( n240443 , n240441 );
and ( n240444 , n240443 , n44686 );
nor ( n240445 , n240442 , n240444 );
not ( n240446 , n240445 );
not ( n240447 , n36572 );
not ( n240448 , n29059 );
and ( n240449 , n240447 , n240448 );
and ( n240450 , n36568 , n29059 );
nor ( n240451 , n240449 , n240450 );
and ( n240452 , n240451 , n32916 );
not ( n240453 , n240451 );
and ( n240454 , n240453 , n32915 );
nor ( n240455 , n240452 , n240454 );
not ( n240456 , n240455 );
not ( n240457 , n34352 );
not ( n240458 , n219430 );
or ( n240459 , n240457 , n240458 );
nand ( n240460 , n37023 , n34357 );
nand ( n240461 , n240459 , n240460 );
and ( n240462 , n240461 , n45773 );
not ( n240463 , n240461 );
and ( n240464 , n240463 , n45770 );
nor ( n240465 , n240462 , n240464 );
nand ( n240466 , n240456 , n240465 );
not ( n240467 , n240466 );
or ( n240468 , n240446 , n240467 );
nand ( n240469 , n240456 , n240465 );
or ( n240470 , n240469 , n240445 );
nand ( n240471 , n240468 , n240470 );
not ( n240472 , n240471 );
xor ( n240473 , n25640 , n221149 );
xor ( n240474 , n240473 , n47938 );
not ( n240475 , n35242 );
not ( n240476 , n36934 );
or ( n240477 , n240475 , n240476 );
or ( n240478 , n52070 , n35242 );
nand ( n240479 , n240477 , n240478 );
and ( n240480 , n240479 , n50335 );
not ( n240481 , n240479 );
and ( n240482 , n240481 , n231699 );
nor ( n240483 , n240480 , n240482 );
not ( n240484 , n240483 );
nand ( n240485 , n240474 , n240484 );
not ( n240486 , n240485 );
buf ( n240487 , n39234 );
xor ( n240488 , n240487 , n43262 );
xor ( n240489 , n240488 , n28405 );
not ( n240490 , n240489 );
and ( n240491 , n240486 , n240490 );
nand ( n240492 , n240474 , n240484 );
and ( n240493 , n240492 , n240489 );
nor ( n240494 , n240491 , n240493 );
not ( n240495 , n240494 );
or ( n240496 , n240472 , n240495 );
or ( n240497 , n240494 , n240471 );
nand ( n240498 , n240496 , n240497 );
not ( n240499 , n240498 );
and ( n240500 , n240434 , n240499 );
and ( n240501 , n240433 , n240498 );
nor ( n240502 , n240500 , n240501 );
not ( n240503 , n240502 );
not ( n240504 , n240503 );
not ( n240505 , n240504 );
and ( n240506 , n240318 , n240505 );
not ( n240507 , n240318 );
buf ( n240508 , n240502 );
and ( n240509 , n240507 , n240508 );
nor ( n240510 , n240506 , n240509 );
not ( n240511 , n49998 );
not ( n240512 , n240511 );
not ( n240513 , n48875 );
or ( n240514 , n240512 , n240513 );
not ( n240515 , n240511 );
nand ( n240516 , n240515 , n48883 );
nand ( n240517 , n240514 , n240516 );
and ( n240518 , n240517 , n226807 );
not ( n240519 , n240517 );
and ( n240520 , n240519 , n49043 );
nor ( n240521 , n240518 , n240520 );
not ( n240522 , n240521 );
nand ( n240523 , n240510 , n240522 );
or ( n240524 , n240158 , n240523 );
not ( n240525 , n240510 );
not ( n240526 , n240157 );
or ( n240527 , n240525 , n240526 );
nor ( n240528 , n240522 , n55104 );
nand ( n240529 , n240527 , n240528 );
nand ( n240530 , n234448 , n25787 );
nand ( n240531 , n240524 , n240529 , n240530 );
buf ( n240532 , n240531 );
buf ( n240533 , n30569 );
not ( n240534 , n240533 );
not ( n240535 , n27801 );
or ( n240536 , n240534 , n240535 );
or ( n240537 , n27801 , n240533 );
nand ( n240538 , n240536 , n240537 );
and ( n240539 , n240538 , n38775 );
not ( n240540 , n240538 );
and ( n240541 , n240540 , n38771 );
nor ( n240542 , n240539 , n240541 );
nand ( n240543 , n240542 , n240445 );
xor ( n240544 , n34679 , n40218 );
xnor ( n240545 , n240544 , n204892 );
and ( n240546 , n240543 , n240545 );
not ( n240547 , n240543 );
not ( n240548 , n240545 );
and ( n240549 , n240547 , n240548 );
nor ( n240550 , n240546 , n240549 );
not ( n240551 , n240550 );
not ( n240552 , n27758 );
not ( n240553 , n31827 );
and ( n240554 , n240552 , n240553 );
and ( n240555 , n27758 , n31827 );
nor ( n240556 , n240554 , n240555 );
xor ( n240557 , n34644 , n240556 );
not ( n240558 , n240557 );
not ( n240559 , n36500 );
not ( n240560 , n40224 );
or ( n240561 , n240559 , n240560 );
or ( n240562 , n40224 , n36500 );
nand ( n240563 , n240561 , n240562 );
and ( n240564 , n240563 , n30537 );
not ( n240565 , n240563 );
not ( n240566 , n40230 );
and ( n240567 , n240565 , n240566 );
nor ( n240568 , n240564 , n240567 );
nand ( n240569 , n240558 , n240568 );
and ( n240570 , n240569 , n240379 );
not ( n240571 , n240569 );
and ( n240572 , n240571 , n240380 );
nor ( n240573 , n240570 , n240572 );
xor ( n240574 , n25709 , n30582 );
xnor ( n240575 , n240574 , n41891 );
not ( n240576 , n32660 );
not ( n240577 , n45308 );
or ( n240578 , n240576 , n240577 );
not ( n240579 , n32660 );
nand ( n240580 , n240579 , n48312 );
nand ( n240581 , n240578 , n240580 );
and ( n240582 , n240581 , n54849 );
not ( n240583 , n240581 );
and ( n240584 , n240583 , n48317 );
nor ( n240585 , n240582 , n240584 );
not ( n240586 , n240585 );
nand ( n240587 , n240575 , n240586 );
not ( n240588 , n240338 );
and ( n240589 , n240587 , n240588 );
not ( n240590 , n240587 );
and ( n240591 , n240590 , n240338 );
nor ( n240592 , n240589 , n240591 );
xor ( n240593 , n240573 , n240592 );
not ( n240594 , n208100 );
not ( n240595 , n29334 );
or ( n240596 , n240594 , n240595 );
or ( n240597 , n46746 , n208100 );
nand ( n240598 , n240596 , n240597 );
and ( n240599 , n240598 , n41149 );
not ( n240600 , n240598 );
and ( n240601 , n240600 , n46753 );
nor ( n240602 , n240599 , n240601 );
not ( n240603 , n240602 );
not ( n240604 , n46585 );
not ( n240605 , n46915 );
not ( n240606 , n240605 );
or ( n240607 , n240604 , n240606 );
not ( n240608 , n46585 );
nand ( n240609 , n240608 , n46915 );
nand ( n240610 , n240607 , n240609 );
and ( n240611 , n240610 , n25766 );
not ( n240612 , n240610 );
and ( n240613 , n240612 , n224685 );
nor ( n240614 , n240611 , n240613 );
not ( n240615 , n240614 );
nand ( n240616 , n240603 , n240615 );
not ( n240617 , n240616 );
not ( n240618 , n240617 );
not ( n240619 , n240399 );
not ( n240620 , n240619 );
or ( n240621 , n240618 , n240620 );
nand ( n240622 , n240399 , n240616 );
nand ( n240623 , n240621 , n240622 );
xor ( n240624 , n240593 , n240623 );
not ( n240625 , n240624 );
not ( n240626 , n32258 );
not ( n240627 , n29563 );
or ( n240628 , n240626 , n240627 );
nand ( n240629 , n220400 , n32255 );
nand ( n240630 , n240628 , n240629 );
and ( n240631 , n240630 , n41971 );
not ( n240632 , n240630 );
and ( n240633 , n240632 , n215031 );
nor ( n240634 , n240631 , n240633 );
buf ( n240635 , RI1749baf0_977);
and ( n240636 , n25454 , n240635 );
not ( n240637 , n25454 );
and ( n240638 , n240637 , n25448 );
nor ( n240639 , n240636 , n240638 );
and ( n240640 , n240639 , n42057 );
not ( n240641 , n240639 );
and ( n240642 , n240641 , n41113 );
or ( n240643 , n240640 , n240642 );
buf ( n240644 , n37946 );
and ( n240645 , n240643 , n240644 );
not ( n240646 , n240643 );
not ( n240647 , n240644 );
and ( n240648 , n240646 , n240647 );
nor ( n240649 , n240645 , n240648 );
not ( n240650 , n240649 );
nand ( n240651 , n240634 , n240650 );
not ( n240652 , n240651 );
not ( n240653 , n240474 );
or ( n240654 , n240652 , n240653 );
or ( n240655 , n240474 , n240651 );
nand ( n240656 , n240654 , n240655 );
not ( n240657 , n240656 );
not ( n240658 , n240657 );
not ( n240659 , n240542 );
nand ( n240660 , n240545 , n240659 );
not ( n240661 , n240660 );
not ( n240662 , n240465 );
and ( n240663 , n240661 , n240662 );
nand ( n240664 , n240545 , n240659 );
and ( n240665 , n240664 , n240465 );
nor ( n240666 , n240663 , n240665 );
not ( n240667 , n240666 );
not ( n240668 , n240667 );
or ( n240669 , n240658 , n240668 );
nand ( n240670 , n240666 , n240656 );
nand ( n240671 , n240669 , n240670 );
and ( n240672 , n240625 , n240671 );
not ( n240673 , n240625 );
not ( n240674 , n240671 );
and ( n240675 , n240673 , n240674 );
nor ( n240676 , n240672 , n240675 );
not ( n240677 , n240676 );
or ( n240678 , n240551 , n240677 );
not ( n240679 , n240550 );
not ( n240680 , n240674 );
not ( n240681 , n240624 );
or ( n240682 , n240680 , n240681 );
nand ( n240683 , n240625 , n240671 );
nand ( n240684 , n240682 , n240683 );
nand ( n240685 , n240679 , n240684 );
nand ( n240686 , n240678 , n240685 );
nand ( n240687 , n36985 , n37025 );
not ( n240688 , n240687 );
buf ( n240689 , n30348 );
not ( n240690 , n240689 );
not ( n240691 , n29335 );
or ( n240692 , n240690 , n240691 );
or ( n240693 , n29335 , n240689 );
nand ( n240694 , n240692 , n240693 );
and ( n240695 , n240694 , n45108 );
not ( n240696 , n240694 );
and ( n240697 , n240696 , n222865 );
nor ( n240698 , n240695 , n240697 );
not ( n240699 , n240698 );
and ( n240700 , n240688 , n240699 );
and ( n240701 , n240687 , n240698 );
nor ( n240702 , n240700 , n240701 );
not ( n240703 , n240702 );
nand ( n240704 , n37273 , n36772 );
not ( n240705 , n40004 );
not ( n240706 , n28646 );
or ( n240707 , n240705 , n240706 );
not ( n240708 , n40004 );
nand ( n240709 , n240708 , n38747 );
nand ( n240710 , n240707 , n240709 );
and ( n240711 , n240710 , n32457 );
not ( n240712 , n240710 );
and ( n240713 , n240712 , n32454 );
nor ( n240714 , n240711 , n240713 );
and ( n240715 , n240704 , n240714 );
not ( n240716 , n240704 );
not ( n240717 , n240714 );
and ( n240718 , n240716 , n240717 );
nor ( n240719 , n240715 , n240718 );
not ( n240720 , n240719 );
or ( n240721 , n240703 , n240720 );
or ( n240722 , n240719 , n240702 );
nand ( n240723 , n240721 , n240722 );
nand ( n240724 , n36894 , n36857 );
not ( n240725 , n205345 );
not ( n240726 , n205348 );
or ( n240727 , n240725 , n240726 );
or ( n240728 , n205348 , n205345 );
nand ( n240729 , n240727 , n240728 );
not ( n240730 , n240729 );
not ( n240731 , n239075 );
or ( n240732 , n240730 , n240731 );
not ( n240733 , n240729 );
nand ( n240734 , n240733 , n31832 );
nand ( n240735 , n240732 , n240734 );
not ( n240736 , n240735 );
not ( n240737 , n38709 );
and ( n240738 , n240736 , n240737 );
and ( n240739 , n240735 , n38704 );
nor ( n240740 , n240738 , n240739 );
and ( n240741 , n240724 , n240740 );
not ( n240742 , n240724 );
not ( n240743 , n240740 );
and ( n240744 , n240742 , n240743 );
nor ( n240745 , n240741 , n240744 );
and ( n240746 , n240723 , n240745 );
not ( n240747 , n240723 );
not ( n240748 , n240745 );
and ( n240749 , n240747 , n240748 );
nor ( n240750 , n240746 , n240749 );
not ( n240751 , n37216 );
nand ( n240752 , n37231 , n240751 );
not ( n240753 , n240752 );
not ( n240754 , n27791 );
not ( n240755 , n49375 );
or ( n240756 , n240754 , n240755 );
or ( n240757 , n31253 , n27791 );
nand ( n240758 , n240756 , n240757 );
and ( n240759 , n240758 , n31264 );
not ( n240760 , n240758 );
and ( n240761 , n240760 , n31273 );
nor ( n240762 , n240759 , n240761 );
not ( n240763 , n240762 );
not ( n240764 , n240763 );
and ( n240765 , n240753 , n240764 );
and ( n240766 , n240752 , n240763 );
nor ( n240767 , n240765 , n240766 );
not ( n240768 , n240767 );
not ( n240769 , n240768 );
not ( n240770 , n37112 );
nand ( n240771 , n240770 , n55128 );
not ( n240772 , n221761 );
not ( n240773 , n37448 );
not ( n240774 , n31899 );
or ( n240775 , n240773 , n240774 );
not ( n240776 , n37448 );
nand ( n240777 , n240776 , n31905 );
nand ( n240778 , n240775 , n240777 );
not ( n240779 , n240778 );
and ( n240780 , n240772 , n240779 );
and ( n240781 , n221761 , n240778 );
nor ( n240782 , n240780 , n240781 );
not ( n240783 , n240782 );
buf ( n240784 , n240783 );
not ( n240785 , n240784 );
and ( n240786 , n240771 , n240785 );
not ( n240787 , n240771 );
and ( n240788 , n240787 , n240784 );
nor ( n240789 , n240786 , n240788 );
not ( n240790 , n240789 );
not ( n240791 , n240790 );
or ( n240792 , n240769 , n240791 );
nand ( n240793 , n240789 , n240767 );
nand ( n240794 , n240792 , n240793 );
not ( n240795 , n240794 );
and ( n240796 , n240750 , n240795 );
not ( n240797 , n240750 );
and ( n240798 , n240797 , n240794 );
nor ( n240799 , n240796 , n240798 );
not ( n240800 , n240799 );
not ( n240801 , n240800 );
and ( n240802 , n240686 , n240801 );
not ( n240803 , n240686 );
not ( n240804 , n240794 );
not ( n240805 , n240750 );
not ( n240806 , n240805 );
or ( n240807 , n240804 , n240806 );
not ( n240808 , n240794 );
nand ( n240809 , n240808 , n240750 );
nand ( n240810 , n240807 , n240809 );
buf ( n240811 , n240810 );
and ( n240812 , n240803 , n240811 );
nor ( n240813 , n240802 , n240812 );
not ( n240814 , n240813 );
nand ( n240815 , n240814 , n235051 );
buf ( n240816 , n40884 );
not ( n240817 , n240816 );
not ( n240818 , n42966 );
or ( n240819 , n240817 , n240818 );
or ( n240820 , n220726 , n240816 );
nand ( n240821 , n240819 , n240820 );
and ( n240822 , n240821 , n38662 );
not ( n240823 , n240821 );
and ( n240824 , n240823 , n38677 );
nor ( n240825 , n240822 , n240824 );
not ( n240826 , n42604 );
not ( n240827 , n34564 );
or ( n240828 , n240826 , n240827 );
nand ( n240829 , n34558 , n42600 );
nand ( n240830 , n240828 , n240829 );
and ( n240831 , n240830 , n42473 );
not ( n240832 , n240830 );
and ( n240833 , n240832 , n42472 );
nor ( n240834 , n240831 , n240833 );
nand ( n240835 , n240825 , n240834 );
not ( n240836 , n37460 );
and ( n240837 , n240835 , n240836 );
not ( n240838 , n240835 );
and ( n240839 , n240838 , n37460 );
nor ( n240840 , n240837 , n240839 );
not ( n240841 , n240840 );
not ( n240842 , n37670 );
buf ( n240843 , n33040 );
not ( n240844 , n240843 );
not ( n240845 , n213924 );
or ( n240846 , n240844 , n240845 );
or ( n240847 , n36168 , n240843 );
nand ( n240848 , n240846 , n240847 );
and ( n240849 , n240848 , n36189 );
not ( n240850 , n240848 );
and ( n240851 , n240850 , n36190 );
nor ( n240852 , n240849 , n240851 );
not ( n240853 , n240852 );
nand ( n240854 , n240842 , n240853 );
not ( n240855 , n240854 );
not ( n240856 , n37681 );
not ( n240857 , n240856 );
and ( n240858 , n240855 , n240857 );
and ( n240859 , n240854 , n240856 );
nor ( n240860 , n240858 , n240859 );
not ( n240861 , n240860 );
not ( n240862 , n240861 );
not ( n240863 , n37512 );
not ( n240864 , n29365 );
not ( n240865 , n31514 );
or ( n240866 , n240864 , n240865 );
not ( n240867 , n29365 );
nand ( n240868 , n240867 , n31527 );
nand ( n240869 , n240866 , n240868 );
and ( n240870 , n240869 , n33849 );
not ( n240871 , n240869 );
and ( n240872 , n240871 , n33853 );
nor ( n240873 , n240870 , n240872 );
not ( n240874 , n240873 );
nand ( n240875 , n240863 , n240874 );
not ( n240876 , n240875 );
not ( n240877 , n37522 );
not ( n240878 , n240877 );
and ( n240879 , n240876 , n240878 );
and ( n240880 , n240875 , n240877 );
nor ( n240881 , n240879 , n240880 );
not ( n240882 , n240881 );
not ( n240883 , n215416 );
buf ( n240884 , n32556 );
not ( n240885 , n240884 );
not ( n240886 , n28461 );
or ( n240887 , n240885 , n240886 );
or ( n240888 , n28461 , n240884 );
nand ( n240889 , n240887 , n240888 );
and ( n240890 , n240889 , n28502 );
not ( n240891 , n240889 );
and ( n240892 , n240891 , n206271 );
nor ( n240893 , n240890 , n240892 );
nor ( n240894 , n37594 , n240893 );
not ( n240895 , n240894 );
or ( n240896 , n240883 , n240895 );
or ( n240897 , n240894 , n215416 );
nand ( n240898 , n240896 , n240897 );
not ( n240899 , n240898 );
or ( n240900 , n240882 , n240899 );
or ( n240901 , n240898 , n240881 );
nand ( n240902 , n240900 , n240901 );
not ( n240903 , n240902 );
not ( n240904 , n240903 );
or ( n240905 , n240862 , n240904 );
nand ( n240906 , n240902 , n240860 );
nand ( n240907 , n240905 , n240906 );
not ( n240908 , n240825 );
nand ( n240909 , n240908 , n240836 );
not ( n240910 , n240909 );
not ( n240911 , n37409 );
not ( n240912 , n240911 );
and ( n240913 , n240910 , n240912 );
and ( n240914 , n240909 , n240911 );
nor ( n240915 , n240913 , n240914 );
not ( n240916 , n240915 );
not ( n240917 , n37311 );
not ( n240918 , n224859 );
buf ( n240919 , n205938 );
not ( n240920 , n240919 );
not ( n240921 , n40743 );
or ( n240922 , n240920 , n240921 );
or ( n240923 , n40743 , n240919 );
nand ( n240924 , n240922 , n240923 );
not ( n240925 , n240924 );
and ( n240926 , n240918 , n240925 );
and ( n240927 , n224859 , n240924 );
nor ( n240928 , n240926 , n240927 );
not ( n240929 , n240928 );
nand ( n240930 , n240917 , n240929 );
buf ( n240931 , n37299 );
xor ( n240932 , n240930 , n240931 );
not ( n240933 , n240932 );
and ( n240934 , n240916 , n240933 );
and ( n240935 , n240915 , n240932 );
nor ( n240936 , n240934 , n240935 );
and ( n240937 , n240907 , n240936 );
not ( n240938 , n240907 );
not ( n240939 , n240936 );
and ( n240940 , n240938 , n240939 );
nor ( n240941 , n240937 , n240940 );
not ( n240942 , n240941 );
or ( n240943 , n240841 , n240942 );
not ( n240944 , n240840 );
and ( n240945 , n240907 , n240939 );
not ( n240946 , n240907 );
and ( n240947 , n240946 , n240936 );
nor ( n240948 , n240945 , n240947 );
nand ( n240949 , n240944 , n240948 );
nand ( n240950 , n240943 , n240949 );
nand ( n240951 , n34816 , n34878 );
not ( n240952 , n240951 );
not ( n240953 , n54053 );
and ( n240954 , n240952 , n240953 );
and ( n240955 , n240951 , n54053 );
nor ( n240956 , n240954 , n240955 );
not ( n240957 , n240956 );
nand ( n240958 , n34765 , n34744 );
and ( n240959 , n240958 , n54071 );
not ( n240960 , n240958 );
and ( n240961 , n240960 , n237719 );
nor ( n240962 , n240959 , n240961 );
not ( n240963 , n240962 );
or ( n240964 , n240957 , n240963 );
or ( n240965 , n240956 , n240962 );
nand ( n240966 , n240964 , n240965 );
nand ( n240967 , n34931 , n34919 );
and ( n240968 , n240967 , n231855 );
not ( n240969 , n240967 );
not ( n240970 , n231855 );
and ( n240971 , n240969 , n240970 );
nor ( n240972 , n240968 , n240971 );
and ( n240973 , n240966 , n240972 );
not ( n240974 , n240966 );
not ( n240975 , n240972 );
and ( n240976 , n240974 , n240975 );
nor ( n240977 , n240973 , n240976 );
not ( n240978 , n34615 );
nand ( n240979 , n240978 , n34600 );
not ( n240980 , n240979 );
not ( n240981 , n39510 );
or ( n240982 , n240980 , n240981 );
not ( n240983 , n34615 );
nand ( n240984 , n240983 , n34600 );
or ( n240985 , n39510 , n240984 );
nand ( n240986 , n240982 , n240985 );
not ( n240987 , n240986 );
not ( n240988 , n54036 );
and ( n240989 , n240987 , n240988 );
and ( n240990 , n240986 , n54036 );
nor ( n240991 , n240989 , n240990 );
nand ( n240992 , n240977 , n240991 );
not ( n240993 , n240977 );
not ( n240994 , n240991 );
nand ( n240995 , n240993 , n240994 );
and ( n240996 , n240992 , n240995 );
not ( n240997 , n240996 );
xor ( n240998 , n240950 , n240997 );
not ( n240999 , n41310 );
nand ( n241000 , n232971 , n41235 );
not ( n241001 , n241000 );
or ( n241002 , n240999 , n241001 );
or ( n241003 , n241000 , n41310 );
nand ( n241004 , n241002 , n241003 );
not ( n241005 , n241004 );
not ( n241006 , n41368 );
nand ( n241007 , n239333 , n41400 );
and ( n241008 , n241007 , n41381 );
not ( n241009 , n241007 );
and ( n241010 , n241009 , n232998 );
nor ( n241011 , n241008 , n241010 );
not ( n241012 , n241011 );
or ( n241013 , n241006 , n241012 );
or ( n241014 , n41368 , n241011 );
nand ( n241015 , n241013 , n241014 );
not ( n241016 , n219219 );
nand ( n241017 , n241016 , n239315 );
and ( n241018 , n241017 , n55218 );
not ( n241019 , n241017 );
and ( n241020 , n241019 , n41475 );
nor ( n241021 , n241018 , n241020 );
and ( n241022 , n241015 , n241021 );
not ( n241023 , n241015 );
not ( n241024 , n241021 );
and ( n241025 , n241023 , n241024 );
nor ( n241026 , n241022 , n241025 );
not ( n241027 , n41606 );
nand ( n241028 , n241027 , n239353 );
not ( n241029 , n241028 );
not ( n241030 , n41589 );
and ( n241031 , n241029 , n241030 );
and ( n241032 , n241028 , n41589 );
nor ( n241033 , n241031 , n241032 );
not ( n241034 , n241033 );
buf ( n241035 , n41540 );
not ( n241036 , n241035 );
nand ( n241037 , n239371 , n241036 );
and ( n241038 , n241037 , n41530 );
not ( n241039 , n241037 );
and ( n241040 , n241039 , n55160 );
nor ( n241041 , n241038 , n241040 );
not ( n241042 , n241041 );
or ( n241043 , n241034 , n241042 );
or ( n241044 , n241041 , n241033 );
nand ( n241045 , n241043 , n241044 );
and ( n241046 , n241026 , n241045 );
not ( n241047 , n241026 );
not ( n241048 , n241045 );
and ( n241049 , n241047 , n241048 );
nor ( n241050 , n241046 , n241049 );
not ( n241051 , n241050 );
or ( n241052 , n241005 , n241051 );
not ( n241053 , n241004 );
not ( n241054 , n241050 );
nand ( n241055 , n241053 , n241054 );
nand ( n241056 , n241052 , n241055 );
buf ( n241057 , n234243 );
and ( n241058 , n241056 , n241057 );
not ( n241059 , n241056 );
buf ( n241060 , n234252 );
and ( n241061 , n241059 , n241060 );
nor ( n241062 , n241058 , n241061 );
nor ( n241063 , n240998 , n241062 );
or ( n241064 , n240815 , n241063 );
not ( n241065 , n222532 );
nor ( n241066 , n240814 , n241065 );
nand ( n241067 , n241066 , n241063 );
buf ( n241068 , n35431 );
nand ( n241069 , n241068 , n27972 );
nand ( n241070 , n241064 , n241067 , n241069 );
buf ( n241071 , n241070 );
not ( n241072 , n238506 );
not ( n241073 , n241072 );
nand ( n241074 , n235453 , n238553 );
not ( n241075 , n241074 );
not ( n241076 , n235442 );
not ( n241077 , n241076 );
and ( n241078 , n241075 , n241077 );
and ( n241079 , n241074 , n241076 );
nor ( n241080 , n241078 , n241079 );
not ( n241081 , n241080 );
not ( n241082 , n235417 );
or ( n241083 , n241081 , n241082 );
or ( n241084 , n235417 , n241080 );
nand ( n241085 , n241083 , n241084 );
not ( n241086 , n235476 );
nand ( n241087 , n241086 , n238496 );
and ( n241088 , n241087 , n235486 );
not ( n241089 , n241087 );
not ( n241090 , n235486 );
and ( n241091 , n241089 , n241090 );
nor ( n241092 , n241088 , n241091 );
and ( n241093 , n241085 , n241092 );
not ( n241094 , n241085 );
not ( n241095 , n241092 );
and ( n241096 , n241094 , n241095 );
nor ( n241097 , n241093 , n241096 );
not ( n241098 , n241097 );
not ( n241099 , n241098 );
not ( n241100 , n238570 );
nand ( n241101 , n235544 , n241100 );
and ( n241102 , n241101 , n235556 );
not ( n241103 , n241101 );
and ( n241104 , n241103 , n235555 );
nor ( n241105 , n241102 , n241104 );
not ( n241106 , n241105 );
not ( n241107 , n241106 );
not ( n241108 , n238592 );
nand ( n241109 , n241108 , n235528 );
and ( n241110 , n241109 , n235518 );
not ( n241111 , n241109 );
and ( n241112 , n241111 , n235517 );
nor ( n241113 , n241110 , n241112 );
not ( n241114 , n241113 );
or ( n241115 , n241107 , n241114 );
not ( n241116 , n241113 );
nand ( n241117 , n241116 , n241105 );
nand ( n241118 , n241115 , n241117 );
not ( n241119 , n241118 );
and ( n241120 , n241099 , n241119 );
and ( n241121 , n241098 , n241118 );
nor ( n241122 , n241120 , n241121 );
not ( n241123 , n241122 );
or ( n241124 , n241073 , n241123 );
not ( n241125 , n241072 );
not ( n241126 , n241097 );
not ( n241127 , n241118 );
not ( n241128 , n241127 );
or ( n241129 , n241126 , n241128 );
nand ( n241130 , n241098 , n241118 );
nand ( n241131 , n241129 , n241130 );
nand ( n241132 , n241125 , n241131 );
nand ( n241133 , n241124 , n241132 );
not ( n241134 , n236402 );
nand ( n241135 , n235617 , n228767 );
not ( n241136 , n241135 );
not ( n241137 , n238414 );
and ( n241138 , n241136 , n241137 );
nand ( n241139 , n235617 , n228767 );
and ( n241140 , n241139 , n238414 );
nor ( n241141 , n241138 , n241140 );
not ( n241142 , n241141 );
or ( n241143 , n241134 , n241142 );
or ( n241144 , n241141 , n236402 );
nand ( n241145 , n241143 , n241144 );
not ( n241146 , n235658 );
nand ( n241147 , n241146 , n51055 );
not ( n241148 , n241147 );
not ( n241149 , n235647 );
and ( n241150 , n241148 , n241149 );
and ( n241151 , n241147 , n235647 );
nor ( n241152 , n241150 , n241151 );
xor ( n241153 , n241145 , n241152 );
not ( n241154 , n51075 );
nand ( n241155 , n235692 , n241154 );
not ( n241156 , n241155 );
not ( n241157 , n238447 );
and ( n241158 , n241156 , n241157 );
and ( n241159 , n241155 , n238447 );
nor ( n241160 , n241158 , n241159 );
not ( n241161 , n241160 );
not ( n241162 , n241161 );
not ( n241163 , n51142 );
nand ( n241164 , n241163 , n235676 );
not ( n241165 , n241164 );
not ( n241166 , n238440 );
or ( n241167 , n241165 , n241166 );
or ( n241168 , n238440 , n241164 );
nand ( n241169 , n241167 , n241168 );
not ( n241170 , n241169 );
not ( n241171 , n241170 );
or ( n241172 , n241162 , n241171 );
nand ( n241173 , n241169 , n241160 );
nand ( n241174 , n241172 , n241173 );
and ( n241175 , n241153 , n241174 );
not ( n241176 , n241153 );
not ( n241177 , n241174 );
and ( n241178 , n241176 , n241177 );
nor ( n241179 , n241175 , n241178 );
buf ( n241180 , n241179 );
not ( n241181 , n241180 );
and ( n241182 , n241133 , n241181 );
not ( n241183 , n241133 );
and ( n241184 , n241183 , n241180 );
nor ( n241185 , n241182 , n241184 );
not ( n241186 , n56059 );
nand ( n241187 , n238881 , n241186 );
not ( n241188 , n241187 );
not ( n241189 , n43419 );
not ( n241190 , n241189 );
and ( n241191 , n241188 , n241190 );
and ( n241192 , n241187 , n241189 );
nor ( n241193 , n241191 , n241192 );
not ( n241194 , n241193 );
not ( n241195 , n241194 );
not ( n241196 , n236631 );
or ( n241197 , n241195 , n241196 );
not ( n241198 , n241194 );
nand ( n241199 , n241198 , n236637 );
nand ( n241200 , n241197 , n241199 );
xor ( n241201 , n241200 , n236766 );
nand ( n241202 , n241185 , n241201 );
not ( n241203 , n236198 );
not ( n241204 , n239013 );
not ( n241205 , n236176 );
nand ( n241206 , n241205 , n52208 );
not ( n241207 , n241206 );
or ( n241208 , n241204 , n241207 );
nand ( n241209 , n241205 , n52208 );
or ( n241210 , n241209 , n239013 );
nand ( n241211 , n241208 , n241210 );
not ( n241212 , n241211 );
nand ( n241213 , n229923 , n236194 );
not ( n241214 , n241213 );
not ( n241215 , n238998 );
and ( n241216 , n241214 , n241215 );
and ( n241217 , n241213 , n238998 );
nor ( n241218 , n241216 , n241217 );
not ( n241219 , n241218 );
or ( n241220 , n241212 , n241219 );
or ( n241221 , n241218 , n241211 );
nand ( n241222 , n241220 , n241221 );
not ( n241223 , n52015 );
nand ( n241224 , n241223 , n236253 );
not ( n241225 , n241224 );
not ( n241226 , n239084 );
and ( n241227 , n241225 , n241226 );
and ( n241228 , n241224 , n239084 );
nor ( n241229 , n241227 , n241228 );
not ( n241230 , n241229 );
not ( n241231 , n239060 );
not ( n241232 , n236233 );
nand ( n241233 , n241232 , n52084 );
not ( n241234 , n241233 );
or ( n241235 , n241231 , n241234 );
or ( n241236 , n241233 , n239060 );
nand ( n241237 , n241235 , n241236 );
not ( n241238 , n241237 );
nand ( n241239 , n236213 , n52125 );
not ( n241240 , n241239 );
not ( n241241 , n239036 );
not ( n241242 , n241241 );
and ( n241243 , n241240 , n241242 );
and ( n241244 , n241239 , n241241 );
nor ( n241245 , n241243 , n241244 );
not ( n241246 , n241245 );
or ( n241247 , n241238 , n241246 );
or ( n241248 , n241245 , n241237 );
nand ( n241249 , n241247 , n241248 );
not ( n241250 , n241249 );
or ( n241251 , n241230 , n241250 );
or ( n241252 , n241249 , n241229 );
nand ( n241253 , n241251 , n241252 );
xor ( n241254 , n241222 , n241253 );
buf ( n241255 , n241254 );
not ( n241256 , n241255 );
not ( n241257 , n241256 );
or ( n241258 , n241203 , n241257 );
not ( n241259 , n236198 );
nand ( n241260 , n241259 , n241255 );
nand ( n241261 , n241258 , n241260 );
not ( n241262 , n44473 );
not ( n241263 , n222229 );
nand ( n241264 , n241262 , n241263 );
not ( n241265 , n241264 );
not ( n241266 , n38411 );
not ( n241267 , n219850 );
or ( n241268 , n241266 , n241267 );
or ( n241269 , n52385 , n38411 );
nand ( n241270 , n241268 , n241269 );
not ( n241271 , n241270 );
not ( n241272 , n36168 );
or ( n241273 , n241271 , n241272 );
or ( n241274 , n238579 , n241270 );
nand ( n241275 , n241273 , n241274 );
buf ( n241276 , n241275 );
not ( n241277 , n241276 );
and ( n241278 , n241265 , n241277 );
nand ( n241279 , n241262 , n241263 );
and ( n241280 , n241279 , n241276 );
nor ( n241281 , n241278 , n241280 );
not ( n241282 , n241281 );
not ( n241283 , n44432 );
not ( n241284 , n222205 );
nand ( n241285 , n241283 , n241284 );
not ( n241286 , n241285 );
not ( n241287 , n29944 );
and ( n241288 , n210737 , n29908 );
not ( n241289 , n210737 );
and ( n241290 , n241289 , n228070 );
nor ( n241291 , n241288 , n241290 );
not ( n241292 , n241291 );
or ( n241293 , n241287 , n241292 );
or ( n241294 , n241291 , n207706 );
nand ( n241295 , n241293 , n241294 );
buf ( n241296 , n241295 );
not ( n241297 , n241296 );
and ( n241298 , n241286 , n241297 );
and ( n241299 , n241285 , n241296 );
nor ( n241300 , n241298 , n241299 );
not ( n241301 , n241300 );
not ( n241302 , n44402 );
not ( n241303 , n222147 );
nand ( n241304 , n241302 , n241303 );
not ( n241305 , n34971 );
not ( n241306 , n226397 );
or ( n241307 , n241305 , n241306 );
not ( n241308 , n34971 );
nand ( n241309 , n241308 , n31926 );
nand ( n241310 , n241307 , n241309 );
and ( n241311 , n241310 , n25550 );
not ( n241312 , n241310 );
and ( n241313 , n241312 , n35224 );
nor ( n241314 , n241311 , n241313 );
buf ( n241315 , n241314 );
xor ( n241316 , n241304 , n241315 );
not ( n241317 , n241316 );
or ( n241318 , n241301 , n241317 );
or ( n241319 , n241300 , n241316 );
nand ( n241320 , n241318 , n241319 );
not ( n241321 , n241320 );
and ( n241322 , n241282 , n241321 );
and ( n241323 , n241281 , n241320 );
nor ( n241324 , n241322 , n241323 );
not ( n241325 , n241324 );
not ( n241326 , n44500 );
nand ( n241327 , n241326 , n44512 );
not ( n241328 , n241327 );
xor ( n241329 , n28795 , n225270 );
xor ( n241330 , n241329 , n34381 );
not ( n241331 , n241330 );
and ( n241332 , n241328 , n241331 );
and ( n241333 , n241327 , n241330 );
nor ( n241334 , n241332 , n241333 );
not ( n241335 , n222281 );
nand ( n241336 , n241335 , n44359 );
not ( n241337 , n31592 );
not ( n241338 , n28680 );
or ( n241339 , n241337 , n241338 );
nand ( n241340 , n37229 , n31589 );
nand ( n241341 , n241339 , n241340 );
and ( n241342 , n241341 , n50950 );
not ( n241343 , n241341 );
and ( n241344 , n241343 , n205096 );
nor ( n241345 , n241342 , n241344 );
not ( n241346 , n241345 );
and ( n241347 , n241336 , n241346 );
not ( n241348 , n241336 );
and ( n241349 , n241348 , n241345 );
nor ( n241350 , n241347 , n241349 );
and ( n241351 , n241334 , n241350 );
not ( n241352 , n241334 );
not ( n241353 , n241350 );
and ( n241354 , n241352 , n241353 );
nor ( n241355 , n241351 , n241354 );
not ( n241356 , n241355 );
not ( n241357 , n241356 );
and ( n241358 , n241325 , n241357 );
and ( n241359 , n241356 , n241324 );
nor ( n241360 , n241358 , n241359 );
buf ( n241361 , n241360 );
and ( n241362 , n241261 , n241361 );
not ( n241363 , n241261 );
not ( n241364 , n241324 );
not ( n241365 , n241364 );
not ( n241366 , n241355 );
or ( n241367 , n241365 , n241366 );
nand ( n241368 , n241324 , n241356 );
nand ( n241369 , n241367 , n241368 );
buf ( n241370 , n241369 );
and ( n241371 , n241363 , n241370 );
nor ( n241372 , n241362 , n241371 );
buf ( n241373 , n222531 );
nand ( n241374 , n241372 , n241373 );
or ( n241375 , n241202 , n241374 );
nor ( n241376 , n241372 , n240080 );
nand ( n241377 , n241376 , n241202 );
buf ( n241378 , n35431 );
nand ( n241379 , n241378 , n205492 );
nand ( n241380 , n241375 , n241377 , n241379 );
buf ( n241381 , n241380 );
not ( n241382 , RI19a88208_2737);
or ( n241383 , n233507 , n241382 );
not ( n241384 , RI19acc5c0_2236);
or ( n241385 , n25335 , n241384 );
nand ( n241386 , n241383 , n241385 );
buf ( n241387 , n241386 );
nand ( n241388 , n47337 , n234320 );
not ( n241389 , n241388 );
not ( n241390 , n47354 );
and ( n241391 , n241389 , n241390 );
and ( n241392 , n241388 , n47354 );
nor ( n241393 , n241391 , n241392 );
not ( n241394 , n241393 );
not ( n241395 , n225128 );
nand ( n241396 , n241395 , n48319 );
not ( n241397 , n241396 );
not ( n241398 , n48255 );
and ( n241399 , n241397 , n241398 );
and ( n241400 , n241396 , n48255 );
nor ( n241401 , n241399 , n241400 );
not ( n241402 , n241401 );
not ( n241403 , n47407 );
nand ( n241404 , n241403 , n48298 );
buf ( n241405 , n225178 );
and ( n241406 , n241404 , n241405 );
not ( n241407 , n241404 );
not ( n241408 , n241405 );
and ( n241409 , n241407 , n241408 );
nor ( n241410 , n241406 , n241409 );
not ( n241411 , n241410 );
or ( n241412 , n241402 , n241411 );
or ( n241413 , n241410 , n241401 );
nand ( n241414 , n241412 , n241413 );
not ( n241415 , n47446 );
nand ( n241416 , n241415 , n226100 );
buf ( n241417 , n47459 );
and ( n241418 , n241416 , n241417 );
not ( n241419 , n241416 );
not ( n241420 , n241417 );
and ( n241421 , n241419 , n241420 );
nor ( n241422 , n241418 , n241421 );
not ( n241423 , n241422 );
and ( n241424 , n241414 , n241423 );
not ( n241425 , n241414 );
and ( n241426 , n241425 , n241422 );
nor ( n241427 , n241424 , n241426 );
not ( n241428 , n241427 );
not ( n241429 , n241428 );
not ( n241430 , n225257 );
nand ( n241431 , n241430 , n48370 );
not ( n241432 , n241431 );
not ( n241433 , n47506 );
not ( n241434 , n241433 );
and ( n241435 , n241432 , n241434 );
nand ( n241436 , n241430 , n48370 );
and ( n241437 , n241436 , n241433 );
nor ( n241438 , n241435 , n241437 );
not ( n241439 , n241438 );
not ( n241440 , n225119 );
or ( n241441 , n241439 , n241440 );
or ( n241442 , n225119 , n241438 );
nand ( n241443 , n241441 , n241442 );
not ( n241444 , n241443 );
not ( n241445 , n241444 );
or ( n241446 , n241429 , n241445 );
nand ( n241447 , n241443 , n241427 );
nand ( n241448 , n241446 , n241447 );
not ( n241449 , n241448 );
or ( n241450 , n241394 , n241449 );
or ( n241451 , n241448 , n241393 );
nand ( n241452 , n241450 , n241451 );
not ( n241453 , n236781 );
not ( n241454 , n241453 );
and ( n241455 , n241452 , n241454 );
not ( n241456 , n241452 );
and ( n241457 , n241456 , n241453 );
nor ( n241458 , n241455 , n241457 );
not ( n241459 , n236795 );
nand ( n241460 , n241458 , n241459 );
not ( n241461 , n34077 );
not ( n241462 , n48039 );
or ( n241463 , n241461 , n241462 );
not ( n241464 , n34077 );
nand ( n241465 , n241464 , n48038 );
nand ( n241466 , n241463 , n241465 );
and ( n241467 , n241466 , n55941 );
not ( n241468 , n241466 );
and ( n241469 , n241468 , n55938 );
nor ( n241470 , n241467 , n241469 );
not ( n241471 , n35047 );
not ( n241472 , n204671 );
or ( n241473 , n241471 , n241472 );
or ( n241474 , n204671 , n35047 );
nand ( n241475 , n241473 , n241474 );
and ( n241476 , n241475 , n26261 );
not ( n241477 , n241475 );
and ( n241478 , n241477 , n204681 );
nor ( n241479 , n241476 , n241478 );
nand ( n241480 , n241470 , n241479 );
not ( n241481 , n241480 );
not ( n241482 , n31144 );
not ( n241483 , n42284 );
or ( n241484 , n241482 , n241483 );
or ( n241485 , n42284 , n31144 );
nand ( n241486 , n241484 , n241485 );
nor ( n241487 , n29989 , n241486 );
not ( n241488 , n241487 );
nand ( n241489 , n241486 , n29990 );
nand ( n241490 , n241488 , n241489 );
not ( n241491 , n241490 );
and ( n241492 , n241481 , n241491 );
and ( n241493 , n241480 , n241490 );
nor ( n241494 , n241492 , n241493 );
not ( n241495 , n241494 );
not ( n241496 , n241495 );
not ( n241497 , n241490 );
not ( n241498 , n241479 );
nand ( n241499 , n241497 , n241498 );
not ( n241500 , n46560 );
not ( n241501 , n232877 );
or ( n241502 , n241500 , n241501 );
or ( n241503 , n35703 , n46560 );
nand ( n241504 , n241502 , n241503 );
and ( n241505 , n241504 , n25762 );
not ( n241506 , n241504 );
and ( n241507 , n241506 , n224685 );
nor ( n241508 , n241505 , n241507 );
and ( n241509 , n241499 , n241508 );
not ( n241510 , n241499 );
not ( n241511 , n241508 );
and ( n241512 , n241510 , n241511 );
nor ( n241513 , n241509 , n241512 );
not ( n241514 , n34736 );
not ( n241515 , n31105 );
not ( n241516 , n34177 );
or ( n241517 , n241515 , n241516 );
nand ( n241518 , n218085 , n31102 );
nand ( n241519 , n241517 , n241518 );
not ( n241520 , n241519 );
and ( n241521 , n241514 , n241520 );
and ( n241522 , n34736 , n241519 );
nor ( n241523 , n241521 , n241522 );
not ( n241524 , n241523 );
not ( n241525 , n25771 );
buf ( n241526 , RI173dc3a8_1682);
not ( n241527 , n241526 );
and ( n241528 , n241525 , n241527 );
and ( n241529 , n25722 , n241526 );
nor ( n241530 , n241528 , n241529 );
and ( n241531 , n241530 , n44347 );
not ( n241532 , n241530 );
and ( n241533 , n241532 , n44351 );
nor ( n241534 , n241531 , n241533 );
not ( n241535 , n241534 );
nand ( n241536 , n241524 , n241535 );
not ( n241537 , n241536 );
not ( n241538 , n37080 );
not ( n241539 , RI17411f58_1420);
xor ( n241540 , n241539 , n29363 );
xor ( n241541 , n241540 , n29370 );
not ( n241542 , n241541 );
or ( n241543 , n241538 , n241542 );
or ( n241544 , n241541 , n37080 );
nand ( n241545 , n241543 , n241544 );
and ( n241546 , n241545 , n29352 );
not ( n241547 , n241545 );
not ( n241548 , n29352 );
and ( n241549 , n241547 , n241548 );
nor ( n241550 , n241546 , n241549 );
not ( n241551 , n241550 );
not ( n241552 , n241551 );
and ( n241553 , n241537 , n241552 );
and ( n241554 , n241536 , n241551 );
nor ( n241555 , n241553 , n241554 );
xor ( n241556 , n241513 , n241555 );
xor ( n241557 , n38883 , n26205 );
xnor ( n241558 , n241557 , n35188 );
not ( n241559 , n241558 );
not ( n241560 , n31452 );
not ( n241561 , n207216 );
or ( n241562 , n241560 , n241561 );
nand ( n241563 , n29456 , n31449 );
nand ( n241564 , n241562 , n241563 );
and ( n241565 , n241564 , n218864 );
not ( n241566 , n241564 );
and ( n241567 , n241566 , n41100 );
nor ( n241568 , n241565 , n241567 );
nand ( n241569 , n241559 , n241568 );
not ( n241570 , n36171 );
not ( n241571 , n44886 );
or ( n241572 , n241570 , n241571 );
or ( n241573 , n28594 , n36171 );
nand ( n241574 , n241572 , n241573 );
and ( n241575 , n241574 , n222643 );
not ( n241576 , n241574 );
and ( n241577 , n241576 , n225104 );
nor ( n241578 , n241575 , n241577 );
buf ( n241579 , n241578 );
xor ( n241580 , n241569 , n241579 );
xnor ( n241581 , n241556 , n241580 );
not ( n241582 , n30856 );
not ( n241583 , n36457 );
or ( n241584 , n241582 , n241583 );
or ( n241585 , n36457 , n30856 );
nand ( n241586 , n241584 , n241585 );
and ( n241587 , n241586 , n39211 );
not ( n241588 , n241586 );
and ( n241589 , n241588 , n43014 );
nor ( n241590 , n241587 , n241589 );
not ( n241591 , n241590 );
not ( n241592 , n34496 );
not ( n241593 , n43636 );
or ( n241594 , n241592 , n241593 );
nand ( n241595 , n50335 , n34493 );
nand ( n241596 , n241594 , n241595 );
not ( n241597 , n241596 );
not ( n241598 , n47330 );
and ( n241599 , n241597 , n241598 );
and ( n241600 , n47330 , n241596 );
nor ( n241601 , n241599 , n241600 );
not ( n241602 , n241601 );
nand ( n241603 , n241591 , n241602 );
not ( n241604 , n241603 );
and ( n241605 , n205361 , n42113 );
not ( n241606 , n205361 );
and ( n241607 , n241606 , n38708 );
or ( n241608 , n241605 , n241607 );
and ( n241609 , n241608 , n219329 );
not ( n241610 , n241608 );
and ( n241611 , n241610 , n31637 );
nor ( n241612 , n241609 , n241611 );
not ( n241613 , n241612 );
not ( n241614 , n241613 );
not ( n241615 , n241614 );
and ( n241616 , n241604 , n241615 );
and ( n241617 , n241603 , n241614 );
nor ( n241618 , n241616 , n241617 );
not ( n241619 , n241618 );
xor ( n241620 , n41840 , n30943 );
xnor ( n241621 , n241620 , n41195 );
not ( n241622 , n25437 );
not ( n241623 , n42058 );
or ( n241624 , n241622 , n241623 );
or ( n241625 , n42058 , n25437 );
nand ( n241626 , n241624 , n241625 );
and ( n241627 , n241626 , n240647 );
not ( n241628 , n241626 );
and ( n241629 , n241628 , n240644 );
nor ( n241630 , n241627 , n241629 );
not ( n241631 , n241630 );
nand ( n241632 , n241621 , n241631 );
not ( n241633 , n41405 );
not ( n241634 , n25349 );
not ( n241635 , n30282 );
or ( n241636 , n241634 , n241635 );
or ( n241637 , n30282 , n25349 );
nand ( n241638 , n241636 , n241637 );
not ( n241639 , n241638 );
or ( n241640 , n241633 , n241639 );
or ( n241641 , n241638 , n41405 );
nand ( n241642 , n241640 , n241641 );
not ( n241643 , n241642 );
and ( n241644 , n241632 , n241643 );
not ( n241645 , n241632 );
and ( n241646 , n241645 , n241642 );
nor ( n241647 , n241644 , n241646 );
not ( n241648 , n241647 );
or ( n241649 , n241619 , n241648 );
or ( n241650 , n241647 , n241618 );
nand ( n241651 , n241649 , n241650 );
and ( n241652 , n241581 , n241651 );
not ( n241653 , n241581 );
not ( n241654 , n241651 );
and ( n241655 , n241653 , n241654 );
nor ( n241656 , n241652 , n241655 );
not ( n241657 , n241656 );
not ( n241658 , n241657 );
or ( n241659 , n241496 , n241658 );
nand ( n241660 , n241656 , n241494 );
nand ( n241661 , n241659 , n241660 );
buf ( n241662 , n49786 );
not ( n241663 , n241662 );
and ( n241664 , n241661 , n241663 );
not ( n241665 , n241661 );
and ( n241666 , n241665 , n241662 );
nor ( n241667 , n241664 , n241666 );
not ( n241668 , n220331 );
not ( n241669 , n241668 );
not ( n241670 , n237639 );
or ( n241671 , n241669 , n241670 );
not ( n241672 , n241668 );
nand ( n241673 , n241672 , n237647 );
nand ( n241674 , n241671 , n241673 );
and ( n241675 , n241674 , n237700 );
not ( n241676 , n241674 );
not ( n241677 , n237704 );
and ( n241678 , n241676 , n241677 );
nor ( n241679 , n241675 , n241678 );
not ( n241680 , n241679 );
nand ( n241681 , n241667 , n241680 );
or ( n241682 , n241460 , n241681 );
not ( n241683 , n241680 );
not ( n241684 , n241458 );
or ( n241685 , n241683 , n241684 );
nor ( n241686 , n241667 , n52445 );
nand ( n241687 , n241685 , n241686 );
nand ( n241688 , n239240 , n29515 );
nand ( n241689 , n241682 , n241687 , n241688 );
buf ( n241690 , n241689 );
not ( n241691 , n229338 );
not ( n241692 , n241691 );
not ( n241693 , n45877 );
or ( n241694 , n241692 , n241693 );
not ( n241695 , n45876 );
or ( n241696 , n241695 , n241691 );
nand ( n241697 , n241694 , n241696 );
and ( n241698 , n241697 , n223836 );
not ( n241699 , n241697 );
not ( n241700 , n223827 );
not ( n241701 , n241700 );
and ( n241702 , n241699 , n241701 );
nor ( n241703 , n241698 , n241702 );
not ( n241704 , n226003 );
nand ( n241705 , n241703 , n241704 );
nand ( n241706 , n237029 , n231176 );
not ( n241707 , n241706 );
not ( n241708 , n53420 );
not ( n241709 , n241708 );
and ( n241710 , n241707 , n241709 );
and ( n241711 , n241706 , n241708 );
nor ( n241712 , n241710 , n241711 );
not ( n241713 , n241712 );
not ( n241714 , n241713 );
not ( n241715 , n231211 );
not ( n241716 , n241715 );
or ( n241717 , n241714 , n241716 );
not ( n241718 , n241713 );
not ( n241719 , n231205 );
and ( n241720 , n241719 , n53448 );
not ( n241721 , n241719 );
and ( n241722 , n241721 , n231094 );
nor ( n241723 , n241720 , n241722 );
nand ( n241724 , n241718 , n241723 );
nand ( n241725 , n241717 , n241724 );
not ( n241726 , n237314 );
not ( n241727 , n28146 );
not ( n241728 , n36995 );
not ( n241729 , n41592 );
or ( n241730 , n241728 , n241729 );
or ( n241731 , n41592 , n36995 );
nand ( n241732 , n241730 , n241731 );
not ( n241733 , n241732 );
and ( n241734 , n241727 , n241733 );
and ( n241735 , n36093 , n241732 );
nor ( n241736 , n241734 , n241735 );
not ( n241737 , n241736 );
not ( n241738 , n31622 );
not ( n241739 , n26102 );
or ( n241740 , n241738 , n241739 );
not ( n241741 , n31622 );
nand ( n241742 , n241741 , n26109 );
nand ( n241743 , n241740 , n241742 );
and ( n241744 , n241743 , n26146 );
not ( n241745 , n241743 );
and ( n241746 , n241745 , n26149 );
nor ( n241747 , n241744 , n241746 );
nand ( n241748 , n241737 , n241747 );
not ( n241749 , n241748 );
or ( n241750 , n241726 , n241749 );
or ( n241751 , n241748 , n237314 );
nand ( n241752 , n241750 , n241751 );
not ( n241753 , n241752 );
not ( n241754 , n29827 );
not ( n241755 , n35548 );
or ( n241756 , n241754 , n241755 );
or ( n241757 , n35548 , n29827 );
nand ( n241758 , n241756 , n241757 );
and ( n241759 , n241758 , n40414 );
not ( n241760 , n241758 );
and ( n241761 , n241760 , n44238 );
nor ( n241762 , n241759 , n241761 );
not ( n241763 , n38056 );
not ( n241764 , n30034 );
or ( n241765 , n241763 , n241764 );
not ( n241766 , n236320 );
or ( n241767 , n241766 , n38056 );
nand ( n241768 , n241765 , n241767 );
and ( n241769 , n241768 , n42756 );
not ( n241770 , n241768 );
and ( n241771 , n241770 , n42760 );
nor ( n241772 , n241769 , n241771 );
nand ( n241773 , n241762 , n241772 );
not ( n241774 , n241773 );
not ( n241775 , n237286 );
and ( n241776 , n241774 , n241775 );
and ( n241777 , n241773 , n237286 );
nor ( n241778 , n241776 , n241777 );
not ( n241779 , n241778 );
or ( n241780 , n241753 , n241779 );
or ( n241781 , n241778 , n241752 );
nand ( n241782 , n241780 , n241781 );
not ( n241783 , n31838 );
not ( n241784 , n224642 );
or ( n241785 , n241783 , n241784 );
or ( n241786 , n224642 , n31838 );
nand ( n241787 , n241785 , n241786 );
buf ( n241788 , n205383 );
xnor ( n241789 , n241787 , n241788 );
not ( n241790 , n27716 );
not ( n241791 , n30147 );
not ( n241792 , n44109 );
or ( n241793 , n241791 , n241792 );
or ( n241794 , n47261 , n30147 );
nand ( n241795 , n241793 , n241794 );
not ( n241796 , n241795 );
or ( n241797 , n241790 , n241796 );
or ( n241798 , n241795 , n27716 );
nand ( n241799 , n241797 , n241798 );
not ( n241800 , n241799 );
nand ( n241801 , n241789 , n241800 );
not ( n241802 , n237172 );
xor ( n241803 , n241801 , n241802 );
not ( n241804 , n241803 );
and ( n241805 , n241782 , n241804 );
not ( n241806 , n241782 );
and ( n241807 , n241806 , n241803 );
nor ( n241808 , n241805 , n241807 );
not ( n241809 , n237230 );
not ( n241810 , n241809 );
not ( n241811 , n241810 );
not ( n241812 , n28973 );
not ( n241813 , n31263 );
or ( n241814 , n241812 , n241813 );
or ( n241815 , n31264 , n28973 );
nand ( n241816 , n241814 , n241815 );
and ( n241817 , n241816 , n30321 );
not ( n241818 , n241816 );
and ( n241819 , n241818 , n35169 );
nor ( n241820 , n241817 , n241819 );
not ( n241821 , n241820 );
not ( n241822 , n26177 );
not ( n241823 , n36626 );
or ( n241824 , n241822 , n241823 );
not ( n241825 , n26177 );
nand ( n241826 , n241825 , n36618 );
nand ( n241827 , n241824 , n241826 );
and ( n241828 , n241827 , n225683 );
not ( n241829 , n241827 );
and ( n241830 , n241829 , n48428 );
nor ( n241831 , n241828 , n241830 );
not ( n241832 , n241831 );
nand ( n241833 , n241821 , n241832 );
not ( n241834 , n241833 );
or ( n241835 , n241811 , n241834 );
not ( n241836 , n241831 );
nand ( n241837 , n241836 , n241821 );
or ( n241838 , n241837 , n241810 );
nand ( n241839 , n241835 , n241838 );
not ( n241840 , n241839 );
not ( n241841 , n33069 );
not ( n241842 , n36812 );
or ( n241843 , n241841 , n241842 );
or ( n241844 , n36812 , n33069 );
nand ( n241845 , n241843 , n241844 );
not ( n241846 , n241845 );
not ( n241847 , n39020 );
or ( n241848 , n241846 , n241847 );
or ( n241849 , n39020 , n241845 );
nand ( n241850 , n241848 , n241849 );
not ( n241851 , n241850 );
not ( n241852 , n30790 );
not ( n241853 , n45468 );
or ( n241854 , n241852 , n241853 );
nand ( n241855 , n51517 , n30786 );
nand ( n241856 , n241854 , n241855 );
and ( n241857 , n241856 , n229282 );
not ( n241858 , n241856 );
and ( n241859 , n241858 , n38912 );
nor ( n241860 , n241857 , n241859 );
not ( n241861 , n241860 );
nand ( n241862 , n241851 , n241861 );
not ( n241863 , n241862 );
buf ( n241864 , n237208 );
not ( n241865 , n241864 );
and ( n241866 , n241863 , n241865 );
and ( n241867 , n241862 , n241864 );
nor ( n241868 , n241866 , n241867 );
not ( n241869 , n241868 );
and ( n241870 , n241840 , n241869 );
and ( n241871 , n241839 , n241868 );
nor ( n241872 , n241870 , n241871 );
and ( n241873 , n241808 , n241872 );
not ( n241874 , n241808 );
not ( n241875 , n241872 );
and ( n241876 , n241874 , n241875 );
nor ( n241877 , n241873 , n241876 );
buf ( n241878 , n241877 );
and ( n241879 , n241725 , n241878 );
not ( n241880 , n241725 );
and ( n241881 , n241808 , n241875 );
not ( n241882 , n241808 );
and ( n241883 , n241882 , n241872 );
nor ( n241884 , n241881 , n241883 );
buf ( n241885 , n241884 );
and ( n241886 , n241880 , n241885 );
nor ( n241887 , n241879 , n241886 );
not ( n241888 , n241887 );
and ( n241889 , n55000 , n55062 );
not ( n241890 , n55000 );
and ( n241891 , n241890 , n55061 );
nor ( n241892 , n241889 , n241891 );
not ( n241893 , n241892 );
not ( n241894 , n54641 );
nand ( n241895 , n241894 , n54616 );
not ( n241896 , n241895 );
not ( n241897 , n55011 );
and ( n241898 , n241896 , n241897 );
not ( n241899 , n54641 );
nand ( n241900 , n241899 , n54616 );
and ( n241901 , n241900 , n55011 );
nor ( n241902 , n241898 , n241901 );
not ( n241903 , n241902 );
nor ( n241904 , n241893 , n241903 );
not ( n241905 , n241904 );
nand ( n241906 , n55067 , n241903 );
nand ( n241907 , n241905 , n241906 );
not ( n241908 , n54417 );
nand ( n241909 , n241908 , n237499 );
and ( n241910 , n241909 , n237489 );
not ( n241911 , n241909 );
not ( n241912 , n237489 );
and ( n241913 , n241911 , n241912 );
nor ( n241914 , n241910 , n241913 );
not ( n241915 , n241914 );
not ( n241916 , n237473 );
nand ( n241917 , n241916 , n54372 );
not ( n241918 , n241917 );
not ( n241919 , n237462 );
and ( n241920 , n241918 , n241919 );
not ( n241921 , n237473 );
nand ( n241922 , n241921 , n54372 );
and ( n241923 , n241922 , n237462 );
nor ( n241924 , n241920 , n241923 );
not ( n241925 , n241924 );
or ( n241926 , n241915 , n241925 );
or ( n241927 , n241924 , n241914 );
nand ( n241928 , n241926 , n241927 );
not ( n241929 , n237520 );
nand ( n241930 , n241929 , n54453 );
and ( n241931 , n241930 , n237510 );
not ( n241932 , n241930 );
not ( n241933 , n237510 );
and ( n241934 , n241932 , n241933 );
nor ( n241935 , n241931 , n241934 );
not ( n241936 , n241935 );
and ( n241937 , n241928 , n241936 );
not ( n241938 , n241928 );
and ( n241939 , n241938 , n241935 );
nor ( n241940 , n241937 , n241939 );
not ( n241941 , n241940 );
nand ( n241942 , n54492 , n237553 );
not ( n241943 , n241942 );
not ( n241944 , n237550 );
and ( n241945 , n241943 , n241944 );
and ( n241946 , n241942 , n237550 );
nor ( n241947 , n241945 , n241946 );
not ( n241948 , n241947 );
nand ( n241949 , n237564 , n54522 );
and ( n241950 , n241949 , n237574 );
not ( n241951 , n241949 );
and ( n241952 , n241951 , n237575 );
or ( n241953 , n241950 , n241952 );
not ( n241954 , n241953 );
or ( n241955 , n241948 , n241954 );
or ( n241956 , n241953 , n241947 );
nand ( n241957 , n241955 , n241956 );
not ( n241958 , n241957 );
and ( n241959 , n241941 , n241958 );
and ( n241960 , n241940 , n241957 );
nor ( n241961 , n241959 , n241960 );
buf ( n241962 , n241961 );
buf ( n241963 , n241962 );
and ( n241964 , n241907 , n241963 );
not ( n241965 , n241907 );
not ( n241966 , n241963 );
and ( n241967 , n241965 , n241966 );
nor ( n241968 , n241964 , n241967 );
nand ( n241969 , n241888 , n241968 );
or ( n241970 , n241705 , n241969 );
not ( n241971 , n241888 );
not ( n241972 , n241703 );
or ( n241973 , n241971 , n241972 );
nor ( n241974 , n241968 , n35816 );
nand ( n241975 , n241973 , n241974 );
buf ( n241976 , n35431 );
nand ( n241977 , n241976 , n30982 );
nand ( n241978 , n241970 , n241975 , n241977 );
buf ( n241979 , n241978 );
not ( n241980 , RI19ace618_2222);
or ( n241981 , n233507 , n241980 );
not ( n241982 , RI19ac5978_2287);
or ( n241983 , n226822 , n241982 );
nand ( n241984 , n241981 , n241983 );
buf ( n241985 , n241984 );
not ( n241986 , RI1754b878_31);
or ( n241987 , n229127 , n241986 );
or ( n241988 , n25335 , n233508 );
nand ( n241989 , n241987 , n241988 );
buf ( n241990 , n241989 );
not ( n241991 , n49048 );
xor ( n241992 , n39448 , n39875 );
xnor ( n241993 , n241992 , n37507 );
nand ( n241994 , n241993 , n241275 );
not ( n241995 , n241994 );
not ( n241996 , n44460 );
and ( n241997 , n241995 , n241996 );
and ( n241998 , n241994 , n44460 );
nor ( n241999 , n241997 , n241998 );
not ( n242000 , n38943 );
not ( n242001 , n204935 );
or ( n242002 , n242000 , n242001 );
or ( n242003 , n204935 , n38943 );
nand ( n242004 , n242002 , n242003 );
and ( n242005 , n242004 , n204977 );
not ( n242006 , n242004 );
and ( n242007 , n242006 , n204976 );
nor ( n242008 , n242005 , n242007 );
nand ( n242009 , n241296 , n242008 );
not ( n242010 , n44425 );
xor ( n242011 , n242009 , n242010 );
not ( n242012 , n242011 );
not ( n242013 , n242012 );
not ( n242014 , n44136 );
and ( n242015 , n34484 , n43635 );
not ( n242016 , n34484 );
and ( n242017 , n242016 , n227480 );
nor ( n242018 , n242015 , n242017 );
not ( n242019 , n242018 );
not ( n242020 , n242019 );
and ( n242021 , n242014 , n242020 );
and ( n242022 , n47330 , n242019 );
nor ( n242023 , n242021 , n242022 );
not ( n242024 , n241314 );
nand ( n242025 , n242023 , n242024 );
not ( n242026 , n242025 );
not ( n242027 , n222137 );
and ( n242028 , n242026 , n242027 );
and ( n242029 , n242025 , n222137 );
nor ( n242030 , n242028 , n242029 );
not ( n242031 , n242030 );
not ( n242032 , n242031 );
or ( n242033 , n242013 , n242032 );
nand ( n242034 , n242030 , n242011 );
nand ( n242035 , n242033 , n242034 );
xor ( n242036 , n241999 , n242035 );
nand ( n242037 , n241345 , n44340 );
and ( n242038 , n242037 , n44354 );
not ( n242039 , n242037 );
and ( n242040 , n242039 , n44522 );
nor ( n242041 , n242038 , n242040 );
not ( n242042 , n242041 );
not ( n242043 , n242042 );
buf ( n242044 , RI17407800_1471);
not ( n242045 , n242044 );
not ( n242046 , n40230 );
or ( n242047 , n242045 , n242046 );
nand ( n242048 , n30533 , n206411 );
nand ( n242049 , n242047 , n242048 );
and ( n242050 , n242049 , n208303 );
not ( n242051 , n242049 );
and ( n242052 , n242051 , n30543 );
nor ( n242053 , n242050 , n242052 );
not ( n242054 , n242053 );
nand ( n242055 , n242054 , n241330 );
not ( n242056 , n242055 );
not ( n242057 , n222252 );
and ( n242058 , n242056 , n242057 );
not ( n242059 , n242053 );
nand ( n242060 , n242059 , n241330 );
and ( n242061 , n242060 , n222252 );
nor ( n242062 , n242058 , n242061 );
not ( n242063 , n242062 );
not ( n242064 , n242063 );
or ( n242065 , n242043 , n242064 );
nand ( n242066 , n242062 , n242041 );
nand ( n242067 , n242065 , n242066 );
xor ( n242068 , n242036 , n242067 );
buf ( n242069 , n242068 );
not ( n242070 , n242069 );
not ( n242071 , n239740 );
not ( n242072 , n239107 );
or ( n242073 , n242071 , n242072 );
not ( n242074 , n239740 );
nand ( n242075 , n242074 , n239099 );
nand ( n242076 , n242073 , n242075 );
not ( n242077 , n242076 );
or ( n242078 , n242070 , n242077 );
not ( n242079 , n242068 );
not ( n242080 , n242079 );
or ( n242081 , n242080 , n242076 );
nand ( n242082 , n242078 , n242081 );
not ( n242083 , n242082 );
nand ( n242084 , n241991 , n242083 );
or ( n242085 , n48565 , n242084 );
not ( n242086 , n241991 );
not ( n242087 , n48564 );
or ( n242088 , n242086 , n242087 );
nor ( n242089 , n242083 , n55152 );
nand ( n242090 , n242088 , n242089 );
nand ( n242091 , n31577 , n26380 );
nand ( n242092 , n242085 , n242090 , n242091 );
buf ( n242093 , n242092 );
not ( n242094 , n204352 );
nand ( n242095 , n31348 , n31430 );
not ( n242096 , n242095 );
or ( n242097 , n242094 , n242096 );
or ( n242098 , n242095 , n204352 );
nand ( n242099 , n242097 , n242098 );
not ( n242100 , n242099 );
not ( n242101 , n25775 );
nand ( n242102 , n31276 , n242101 );
not ( n242103 , n242102 );
not ( n242104 , n228318 );
and ( n242105 , n242103 , n242104 );
and ( n242106 , n242102 , n228318 );
nor ( n242107 , n242105 , n242106 );
not ( n242108 , n242107 );
not ( n242109 , n242108 );
not ( n242110 , n204352 );
nand ( n242111 , n242110 , n31349 );
not ( n242112 , n242111 );
not ( n242113 , n204447 );
and ( n242114 , n242112 , n242113 );
and ( n242115 , n242111 , n204447 );
nor ( n242116 , n242114 , n242115 );
not ( n242117 , n242116 );
not ( n242118 , n25606 );
or ( n242119 , n242117 , n242118 );
or ( n242120 , n25606 , n242116 );
nand ( n242121 , n242119 , n242120 );
not ( n242122 , n242121 );
not ( n242123 , n242122 );
or ( n242124 , n242109 , n242123 );
nand ( n242125 , n242121 , n242107 );
nand ( n242126 , n242124 , n242125 );
nand ( n242127 , n31215 , n26321 );
not ( n242128 , n242127 );
not ( n242129 , n26223 );
and ( n242130 , n242128 , n242129 );
and ( n242131 , n242127 , n26223 );
nor ( n242132 , n242130 , n242131 );
not ( n242133 , n242132 );
not ( n242134 , n26057 );
nand ( n242135 , n208778 , n242134 );
and ( n242136 , n242135 , n26151 );
not ( n242137 , n242135 );
and ( n242138 , n242137 , n228332 );
nor ( n242139 , n242136 , n242138 );
not ( n242140 , n242139 );
and ( n242141 , n242133 , n242140 );
and ( n242142 , n242132 , n242139 );
nor ( n242143 , n242141 , n242142 );
and ( n242144 , n242126 , n242143 );
not ( n242145 , n242126 );
not ( n242146 , n242143 );
and ( n242147 , n242145 , n242146 );
nor ( n242148 , n242144 , n242147 );
not ( n242149 , n242148 );
or ( n242150 , n242100 , n242149 );
not ( n242151 , n242099 );
and ( n242152 , n242126 , n242146 );
not ( n242153 , n242126 );
and ( n242154 , n242153 , n242143 );
nor ( n242155 , n242152 , n242154 );
nand ( n242156 , n242151 , n242155 );
nand ( n242157 , n242150 , n242156 );
not ( n242158 , n35626 );
nand ( n242159 , n242158 , n205076 );
and ( n242160 , n242159 , n205146 );
not ( n242161 , n242159 );
and ( n242162 , n242161 , n205145 );
nor ( n242163 , n242160 , n242162 );
nand ( n242164 , n205245 , n35600 );
and ( n242165 , n242164 , n205328 );
not ( n242166 , n242164 );
and ( n242167 , n242166 , n205327 );
nor ( n242168 , n242165 , n242167 );
xor ( n242169 , n242163 , n242168 );
not ( n242170 , n27679 );
nand ( n242171 , n35467 , n27765 );
not ( n242172 , n242171 );
or ( n242173 , n242170 , n242172 );
or ( n242174 , n242171 , n27679 );
nand ( n242175 , n242173 , n242174 );
xnor ( n242176 , n242169 , n242175 );
not ( n242177 , n242176 );
nand ( n242178 , n204634 , n35749 );
not ( n242179 , n242178 );
not ( n242180 , n204685 );
and ( n242181 , n242179 , n242180 );
and ( n242182 , n242178 , n204685 );
nor ( n242183 , n242181 , n242182 );
not ( n242184 , n242183 );
not ( n242185 , n242184 );
not ( n242186 , n204897 );
nand ( n242187 , n242186 , n35730 );
and ( n242188 , n242187 , n204827 );
not ( n242189 , n242187 );
and ( n242190 , n242189 , n204826 );
nor ( n242191 , n242188 , n242190 );
not ( n242192 , n242191 );
not ( n242193 , n242192 );
or ( n242194 , n242185 , n242193 );
nand ( n242195 , n242191 , n242183 );
nand ( n242196 , n242194 , n242195 );
not ( n242197 , n242196 );
and ( n242198 , n242177 , n242197 );
and ( n242199 , n242176 , n242196 );
nor ( n242200 , n242198 , n242199 );
not ( n242201 , n242200 );
not ( n242202 , n242201 );
and ( n242203 , n242157 , n242202 );
not ( n242204 , n242157 );
not ( n242205 , n242200 );
buf ( n242206 , n242205 );
and ( n242207 , n242204 , n242206 );
nor ( n242208 , n242203 , n242207 );
nor ( n242209 , n242208 , n54208 );
not ( n242210 , n41813 );
not ( n242211 , n233090 );
or ( n242212 , n242210 , n242211 );
or ( n242213 , n233090 , n41813 );
nand ( n242214 , n242212 , n242213 );
not ( n242215 , n242214 );
not ( n242216 , n43648 );
nand ( n242217 , n242216 , n221303 );
and ( n242218 , n242217 , n220157 );
not ( n242219 , n242217 );
not ( n242220 , n220157 );
and ( n242221 , n242219 , n242220 );
nor ( n242222 , n242218 , n242221 );
not ( n242223 , n242222 );
not ( n242224 , n242223 );
not ( n242225 , n43596 );
nand ( n242226 , n242225 , n43581 );
not ( n242227 , n242226 );
not ( n242228 , n42334 );
and ( n242229 , n242227 , n242228 );
and ( n242230 , n242226 , n42334 );
nor ( n242231 , n242229 , n242230 );
not ( n242232 , n242231 );
not ( n242233 , n242232 );
or ( n242234 , n242224 , n242233 );
nand ( n242235 , n242231 , n242222 );
nand ( n242236 , n242234 , n242235 );
nand ( n242237 , n230864 , n55766 );
xnor ( n242238 , n242237 , n53105 );
not ( n242239 , n242238 );
and ( n242240 , n242236 , n242239 );
not ( n242241 , n242236 );
and ( n242242 , n242241 , n242238 );
nor ( n242243 , n242240 , n242242 );
not ( n242244 , n242243 );
not ( n242245 , n242244 );
nand ( n242246 , n234284 , n43681 );
not ( n242247 , n242246 );
not ( n242248 , n53113 );
and ( n242249 , n242247 , n242248 );
and ( n242250 , n242246 , n53113 );
nor ( n242251 , n242249 , n242250 );
not ( n242252 , n242251 );
not ( n242253 , n242252 );
not ( n242254 , n43691 );
nand ( n242255 , n242254 , n234273 );
not ( n242256 , n242255 );
not ( n242257 , n53124 );
not ( n242258 , n242257 );
and ( n242259 , n242256 , n242258 );
and ( n242260 , n242255 , n242257 );
nor ( n242261 , n242259 , n242260 );
not ( n242262 , n242261 );
or ( n242263 , n242253 , n242262 );
not ( n242264 , n242261 );
nand ( n242265 , n242264 , n242251 );
nand ( n242266 , n242263 , n242265 );
not ( n242267 , n242266 );
and ( n242268 , n242245 , n242267 );
and ( n242269 , n242244 , n242266 );
nor ( n242270 , n242268 , n242269 );
not ( n242271 , n242270 );
not ( n242272 , n242271 );
not ( n242273 , n242272 );
and ( n242274 , n242215 , n242273 );
and ( n242275 , n242214 , n242272 );
nor ( n242276 , n242274 , n242275 );
not ( n242277 , n242276 );
not ( n242278 , n54115 );
not ( n242279 , n234005 );
not ( n242280 , n237725 );
or ( n242281 , n242279 , n242280 );
or ( n242282 , n234005 , n237725 );
nand ( n242283 , n242281 , n242282 );
nand ( n242284 , n54096 , n240970 );
not ( n242285 , n242284 );
not ( n242286 , n34942 );
and ( n242287 , n242285 , n242286 );
and ( n242288 , n242284 , n34942 );
nor ( n242289 , n242287 , n242288 );
xor ( n242290 , n242283 , n242289 );
nand ( n242291 , n54032 , n231881 );
not ( n242292 , n242291 );
not ( n242293 , n34625 );
and ( n242294 , n242292 , n242293 );
and ( n242295 , n242291 , n34625 );
nor ( n242296 , n242294 , n242295 );
not ( n242297 , n242296 );
not ( n242298 , n242297 );
not ( n242299 , n39599 );
or ( n242300 , n242298 , n242299 );
nand ( n242301 , n39515 , n242296 );
nand ( n242302 , n242300 , n242301 );
and ( n242303 , n242290 , n242302 );
not ( n242304 , n242290 );
not ( n242305 , n242302 );
and ( n242306 , n242304 , n242305 );
nor ( n242307 , n242303 , n242306 );
not ( n242308 , n242307 );
or ( n242309 , n242278 , n242308 );
not ( n242310 , n54115 );
and ( n242311 , n242290 , n242302 );
not ( n242312 , n242290 );
and ( n242313 , n242312 , n242305 );
nor ( n242314 , n242311 , n242313 );
not ( n242315 , n242314 );
nand ( n242316 , n242310 , n242315 );
nand ( n242317 , n242309 , n242316 );
not ( n242318 , n35303 );
nand ( n242319 , n46176 , n54171 );
not ( n242320 , n242319 );
or ( n242321 , n242318 , n242320 );
or ( n242322 , n242319 , n35303 );
nand ( n242323 , n242321 , n242322 );
not ( n242324 , n242323 );
not ( n242325 , n242324 );
not ( n242326 , n217478 );
nand ( n242327 , n46157 , n242326 );
not ( n242328 , n242327 );
not ( n242329 , n35287 );
and ( n242330 , n242328 , n242329 );
and ( n242331 , n242327 , n35287 );
nor ( n242332 , n242330 , n242331 );
not ( n242333 , n242332 );
not ( n242334 , n242333 );
or ( n242335 , n242325 , n242334 );
nand ( n242336 , n242332 , n242323 );
nand ( n242337 , n242335 , n242336 );
not ( n242338 , n242337 );
not ( n242339 , n242338 );
not ( n242340 , n39643 );
nand ( n242341 , n242340 , n46100 );
not ( n242342 , n242341 );
not ( n242343 , n35119 );
and ( n242344 , n242342 , n242343 );
and ( n242345 , n242341 , n35119 );
nor ( n242346 , n242344 , n242345 );
not ( n242347 , n242346 );
nand ( n242348 , n223880 , n54148 );
and ( n242349 , n242348 , n35030 );
not ( n242350 , n242348 );
and ( n242351 , n242350 , n35031 );
nor ( n242352 , n242349 , n242351 );
not ( n242353 , n242352 );
or ( n242354 , n242347 , n242353 );
or ( n242355 , n242352 , n242346 );
nand ( n242356 , n242354 , n242355 );
not ( n242357 , n39681 );
nand ( n242358 , n242357 , n46134 );
not ( n242359 , n242358 );
not ( n242360 , n35193 );
and ( n242361 , n242359 , n242360 );
and ( n242362 , n242358 , n35193 );
nor ( n242363 , n242361 , n242362 );
and ( n242364 , n242356 , n242363 );
not ( n242365 , n242356 );
not ( n242366 , n242363 );
and ( n242367 , n242365 , n242366 );
nor ( n242368 , n242364 , n242367 );
not ( n242369 , n242368 );
not ( n242370 , n242369 );
or ( n242371 , n242339 , n242370 );
nand ( n242372 , n242368 , n242337 );
nand ( n242373 , n242371 , n242372 );
buf ( n242374 , n242373 );
and ( n242375 , n242317 , n242374 );
not ( n242376 , n242317 );
and ( n242377 , n242368 , n242337 );
not ( n242378 , n242368 );
and ( n242379 , n242378 , n242338 );
nor ( n242380 , n242377 , n242379 );
buf ( n242381 , n242380 );
and ( n242382 , n242376 , n242381 );
nor ( n242383 , n242375 , n242382 );
nor ( n242384 , n242277 , n242383 );
nand ( n242385 , n242209 , n242384 );
not ( n242386 , n242208 );
not ( n242387 , n242386 );
not ( n242388 , n242276 );
or ( n242389 , n242387 , n242388 );
not ( n242390 , n242383 );
not ( n242391 , n241373 );
nor ( n242392 , n242390 , n242391 );
nand ( n242393 , n242389 , n242392 );
nand ( n242394 , n238638 , n219094 );
nand ( n242395 , n242385 , n242393 , n242394 );
buf ( n242396 , n242395 );
not ( n242397 , n204356 );
not ( n242398 , n234823 );
or ( n242399 , n242397 , n242398 );
not ( n242400 , n55681 );
not ( n242401 , n242400 );
not ( n242402 , n235008 );
or ( n242403 , n242401 , n242402 );
not ( n242404 , n242400 );
nand ( n242405 , n242404 , n235016 );
nand ( n242406 , n242403 , n242405 );
and ( n242407 , n242406 , n235022 );
not ( n242408 , n242406 );
and ( n242409 , n242408 , n235019 );
nor ( n242410 , n242407 , n242409 );
not ( n242411 , n204853 );
not ( n242412 , n37464 );
or ( n242413 , n242411 , n242412 );
not ( n242414 , n204853 );
nand ( n242415 , n242414 , n28876 );
nand ( n242416 , n242413 , n242415 );
xnor ( n242417 , n242416 , n37472 );
buf ( n242418 , n215106 );
not ( n242419 , n242418 );
not ( n242420 , n41754 );
or ( n242421 , n242419 , n242420 );
or ( n242422 , n41754 , n242418 );
nand ( n242423 , n242421 , n242422 );
and ( n242424 , n242423 , n47112 );
not ( n242425 , n242423 );
and ( n242426 , n242425 , n228145 );
nor ( n242427 , n242424 , n242426 );
buf ( n242428 , n242427 );
nand ( n242429 , n242417 , n242428 );
not ( n242430 , n241568 );
and ( n242431 , n242429 , n242430 );
not ( n242432 , n242429 );
and ( n242433 , n242432 , n241568 );
nor ( n242434 , n242431 , n242433 );
not ( n242435 , n242434 );
not ( n242436 , n242435 );
not ( n242437 , n241494 );
buf ( n242438 , n32596 );
and ( n242439 , n242438 , n28508 );
not ( n242440 , n242438 );
and ( n242441 , n242440 , n28502 );
nor ( n242442 , n242439 , n242441 );
not ( n242443 , n242442 );
and ( n242444 , n44690 , n242443 );
not ( n242445 , n44690 );
and ( n242446 , n242445 , n242442 );
nor ( n242447 , n242444 , n242446 );
not ( n242448 , n242447 );
nand ( n242449 , n241523 , n242448 );
and ( n242450 , n242449 , n241535 );
not ( n242451 , n242449 );
and ( n242452 , n242451 , n241534 );
nor ( n242453 , n242450 , n242452 );
not ( n242454 , n242453 );
or ( n242455 , n242437 , n242454 );
or ( n242456 , n242453 , n241494 );
nand ( n242457 , n242455 , n242456 );
not ( n242458 , n241558 );
not ( n242459 , n242417 );
nand ( n242460 , n242459 , n242430 );
not ( n242461 , n242460 );
and ( n242462 , n242458 , n242461 );
and ( n242463 , n241558 , n242460 );
nor ( n242464 , n242462 , n242463 );
and ( n242465 , n242457 , n242464 );
not ( n242466 , n242457 );
not ( n242467 , n242464 );
and ( n242468 , n242466 , n242467 );
nor ( n242469 , n242465 , n242468 );
not ( n242470 , n241590 );
not ( n242471 , n55481 );
buf ( n242472 , n31341 );
buf ( n242473 , RI1749ffd8_956);
and ( n242474 , n242472 , n242473 );
not ( n242475 , n242472 );
and ( n242476 , n242475 , n31338 );
nor ( n242477 , n242474 , n242476 );
not ( n242478 , n242477 );
not ( n242479 , n31613 );
or ( n242480 , n242478 , n242479 );
or ( n242481 , n51033 , n242477 );
nand ( n242482 , n242480 , n242481 );
not ( n242483 , n242482 );
or ( n242484 , n242471 , n242483 );
or ( n242485 , n242482 , n50111 );
nand ( n242486 , n242484 , n242485 );
nand ( n242487 , n241601 , n242486 );
not ( n242488 , n242487 );
or ( n242489 , n242470 , n242488 );
or ( n242490 , n242487 , n241590 );
nand ( n242491 , n242489 , n242490 );
not ( n242492 , n242491 );
not ( n242493 , n241621 );
buf ( n242494 , n38557 );
not ( n242495 , n242494 );
not ( n242496 , n33473 );
or ( n242497 , n242495 , n242496 );
or ( n242498 , n40772 , n242494 );
nand ( n242499 , n242497 , n242498 );
not ( n242500 , n242499 );
not ( n242501 , n43696 );
or ( n242502 , n242500 , n242501 );
or ( n242503 , n52635 , n242499 );
nand ( n242504 , n242502 , n242503 );
nand ( n242505 , n242493 , n242504 );
and ( n242506 , n242505 , n241631 );
not ( n242507 , n242505 );
and ( n242508 , n242507 , n241630 );
nor ( n242509 , n242506 , n242508 );
not ( n242510 , n242509 );
not ( n242511 , n242510 );
or ( n242512 , n242492 , n242511 );
not ( n242513 , n242491 );
nand ( n242514 , n242513 , n242509 );
nand ( n242515 , n242512 , n242514 );
not ( n242516 , n242515 );
and ( n242517 , n242469 , n242516 );
not ( n242518 , n242469 );
and ( n242519 , n242518 , n242515 );
nor ( n242520 , n242517 , n242519 );
not ( n242521 , n242520 );
or ( n242522 , n242436 , n242521 );
not ( n242523 , n242435 );
and ( n242524 , n242469 , n242515 );
not ( n242525 , n242469 );
and ( n242526 , n242525 , n242516 );
nor ( n242527 , n242524 , n242526 );
nand ( n242528 , n242523 , n242527 );
nand ( n242529 , n242522 , n242528 );
nor ( n242530 , n49727 , n38914 );
not ( n242531 , n242530 );
not ( n242532 , n49714 );
and ( n242533 , n242531 , n242532 );
and ( n242534 , n242530 , n49714 );
nor ( n242535 , n242533 , n242534 );
not ( n242536 , n242535 );
not ( n242537 , n49645 );
or ( n242538 , n242536 , n242537 );
or ( n242539 , n49645 , n242535 );
nand ( n242540 , n242538 , n242539 );
not ( n242541 , n242540 );
nand ( n242542 , n49761 , n39038 );
not ( n242543 , n242542 );
not ( n242544 , n49757 );
and ( n242545 , n242543 , n242544 );
and ( n242546 , n242542 , n49757 );
nor ( n242547 , n242545 , n242546 );
not ( n242548 , n242547 );
and ( n242549 , n242541 , n242548 );
and ( n242550 , n242540 , n242547 );
nor ( n242551 , n242549 , n242550 );
not ( n242552 , n49687 );
not ( n242553 , n242552 );
not ( n242554 , n49697 );
nand ( n242555 , n38756 , n242554 );
not ( n242556 , n242555 );
or ( n242557 , n242553 , n242556 );
or ( n242558 , n242555 , n242552 );
nand ( n242559 , n242557 , n242558 );
not ( n242560 , n242559 );
not ( n242561 , n237372 );
or ( n242562 , n242560 , n242561 );
or ( n242563 , n237372 , n242559 );
nand ( n242564 , n242562 , n242563 );
and ( n242565 , n242551 , n242564 );
not ( n242566 , n242551 );
not ( n242567 , n242564 );
and ( n242568 , n242566 , n242567 );
nor ( n242569 , n242565 , n242568 );
buf ( n242570 , n242569 );
not ( n242571 , n242570 );
and ( n242572 , n242529 , n242571 );
not ( n242573 , n242529 );
not ( n242574 , n242569 );
not ( n242575 , n242574 );
and ( n242576 , n242573 , n242575 );
nor ( n242577 , n242572 , n242576 );
nand ( n242578 , n242410 , n242577 );
not ( n242579 , n236444 );
and ( n242580 , n32096 , n32468 );
not ( n242581 , n32096 );
not ( n242582 , n32468 );
and ( n242583 , n242581 , n242582 );
nor ( n242584 , n242580 , n242583 );
not ( n242585 , n242584 );
not ( n242586 , n242585 );
or ( n242587 , n242579 , n242586 );
or ( n242588 , n32473 , n236444 );
nand ( n242589 , n242587 , n242588 );
not ( n242590 , n242589 );
not ( n242591 , n33247 );
and ( n242592 , n242590 , n242591 );
and ( n242593 , n242589 , n33247 );
nor ( n242594 , n242592 , n242593 );
not ( n242595 , n242594 );
and ( n242596 , n242578 , n242595 );
not ( n242597 , n242578 );
and ( n242598 , n242597 , n242594 );
nor ( n242599 , n242596 , n242598 );
or ( n242600 , n242599 , n235052 );
nand ( n242601 , n242399 , n242600 );
buf ( n242602 , n242601 );
not ( n242603 , RI19a852b0_2758);
or ( n242604 , n233507 , n242603 );
not ( n242605 , RI19aca040_2255);
or ( n242606 , n25335 , n242605 );
nand ( n242607 , n242604 , n242606 );
buf ( n242608 , n242607 );
not ( n242609 , n234760 );
not ( n242610 , n242609 );
not ( n242611 , n234786 );
nand ( n242612 , n242611 , n234788 );
not ( n242613 , n242612 );
not ( n242614 , n34400 );
and ( n242615 , n242613 , n242614 );
and ( n242616 , n242612 , n34400 );
nor ( n242617 , n242615 , n242616 );
not ( n242618 , n242617 );
not ( n242619 , n242618 );
not ( n242620 , n234755 );
nand ( n242621 , n242620 , n234744 );
not ( n242622 , n242621 );
not ( n242623 , n34229 );
and ( n242624 , n242622 , n242623 );
not ( n242625 , n234755 );
nand ( n242626 , n242625 , n234744 );
and ( n242627 , n242626 , n34229 );
nor ( n242628 , n242624 , n242627 );
not ( n242629 , n242628 );
not ( n242630 , n234763 );
nand ( n242631 , n242630 , n234775 );
not ( n242632 , n33897 );
and ( n242633 , n242631 , n242632 );
not ( n242634 , n242631 );
and ( n242635 , n242634 , n33897 );
nor ( n242636 , n242633 , n242635 );
not ( n242637 , n242636 );
or ( n242638 , n242629 , n242637 );
or ( n242639 , n242636 , n242628 );
nand ( n242640 , n242638 , n242639 );
not ( n242641 , n242640 );
not ( n242642 , n242641 );
or ( n242643 , n242619 , n242642 );
nand ( n242644 , n242640 , n242617 );
nand ( n242645 , n242643 , n242644 );
not ( n242646 , n34349 );
not ( n242647 , n234727 );
not ( n242648 , n234714 );
nand ( n242649 , n242647 , n242648 );
not ( n242650 , n242649 );
or ( n242651 , n242646 , n242650 );
not ( n242652 , n234727 );
nand ( n242653 , n242652 , n242648 );
or ( n242654 , n242653 , n34349 );
nand ( n242655 , n242651 , n242654 );
not ( n242656 , n242655 );
not ( n242657 , n242656 );
nand ( n242658 , n234707 , n234702 );
not ( n242659 , n242658 );
buf ( n242660 , n34106 );
not ( n242661 , n242660 );
and ( n242662 , n242659 , n242661 );
and ( n242663 , n242658 , n242660 );
nor ( n242664 , n242662 , n242663 );
not ( n242665 , n242664 );
not ( n242666 , n242665 );
or ( n242667 , n242657 , n242666 );
nand ( n242668 , n242664 , n242655 );
nand ( n242669 , n242667 , n242668 );
not ( n242670 , n242669 );
and ( n242671 , n242645 , n242670 );
not ( n242672 , n242645 );
and ( n242673 , n242672 , n242669 );
nor ( n242674 , n242671 , n242673 );
not ( n242675 , n242674 );
not ( n242676 , n242675 );
or ( n242677 , n242610 , n242676 );
or ( n242678 , n242675 , n242609 );
nand ( n242679 , n242677 , n242678 );
buf ( n242680 , n28929 );
and ( n242681 , n242679 , n242680 );
not ( n242682 , n242679 );
buf ( n242683 , n28936 );
and ( n242684 , n242682 , n242683 );
nor ( n242685 , n242681 , n242684 );
not ( n242686 , n242685 );
nand ( n242687 , n242686 , n241704 );
nand ( n242688 , n236601 , n238850 );
and ( n242689 , n242688 , n43314 );
not ( n242690 , n242688 );
and ( n242691 , n242690 , n43315 );
nor ( n242692 , n242689 , n242691 );
not ( n242693 , n242692 );
not ( n242694 , n236631 );
or ( n242695 , n242693 , n242694 );
buf ( n242696 , n236631 );
or ( n242697 , n242696 , n242692 );
nand ( n242698 , n242695 , n242697 );
buf ( n242699 , n236762 );
and ( n242700 , n242698 , n242699 );
not ( n242701 , n242698 );
and ( n242702 , n242701 , n236763 );
nor ( n242703 , n242700 , n242702 );
buf ( n242704 , n37104 );
not ( n242705 , n242704 );
not ( n242706 , n241541 );
not ( n242707 , n242706 );
or ( n242708 , n242705 , n242707 );
or ( n242709 , n242706 , n242704 );
nand ( n242710 , n242708 , n242709 );
and ( n242711 , n242710 , n241548 );
not ( n242712 , n242710 );
and ( n242713 , n242712 , n29352 );
nor ( n242714 , n242711 , n242713 );
not ( n242715 , n242714 );
not ( n242716 , n52850 );
not ( n242717 , n52873 );
nand ( n242718 , n242716 , n242717 );
not ( n242719 , n242718 );
or ( n242720 , n242715 , n242719 );
or ( n242721 , n242718 , n242714 );
nand ( n242722 , n242720 , n242721 );
not ( n242723 , n242722 );
not ( n242724 , n242723 );
not ( n242725 , n33934 );
not ( n242726 , n204726 );
or ( n242727 , n242725 , n242726 );
or ( n242728 , n204726 , n33934 );
nand ( n242729 , n242727 , n242728 );
not ( n242730 , n242729 );
not ( n242731 , n31735 );
or ( n242732 , n242730 , n242731 );
or ( n242733 , n36702 , n242729 );
nand ( n242734 , n242732 , n242733 );
nor ( n242735 , n242734 , n52885 );
not ( n242736 , n242735 );
not ( n242737 , n52783 );
not ( n242738 , n242737 );
and ( n242739 , n242736 , n242738 );
and ( n242740 , n242735 , n242737 );
nor ( n242741 , n242739 , n242740 );
not ( n242742 , n38514 );
buf ( n242743 , n40167 );
not ( n242744 , n242743 );
not ( n242745 , n38558 );
or ( n242746 , n242744 , n242745 );
or ( n242747 , n38558 , n242743 );
nand ( n242748 , n242746 , n242747 );
not ( n242749 , n242748 );
and ( n242750 , n242742 , n242749 );
and ( n242751 , n38570 , n242748 );
nor ( n242752 , n242750 , n242751 );
nand ( n242753 , n242752 , n230594 );
not ( n242754 , n234718 );
not ( n242755 , n29034 );
and ( n242756 , n242754 , n242755 );
and ( n242757 , n28043 , n29034 );
nor ( n242758 , n242756 , n242757 );
not ( n242759 , n242758 );
xor ( n242760 , n36572 , n242759 );
and ( n242761 , n242753 , n242760 );
not ( n242762 , n242753 );
not ( n242763 , n242760 );
and ( n242764 , n242762 , n242763 );
nor ( n242765 , n242761 , n242764 );
xor ( n242766 , n242741 , n242765 );
not ( n242767 , n46810 );
not ( n242768 , n45789 );
not ( n242769 , n39001 );
or ( n242770 , n242768 , n242769 );
or ( n242771 , n39001 , n45789 );
nand ( n242772 , n242770 , n242771 );
not ( n242773 , n242772 );
or ( n242774 , n242767 , n242773 );
or ( n242775 , n242772 , n46810 );
nand ( n242776 , n242774 , n242775 );
not ( n242777 , n242776 );
not ( n242778 , n242714 );
nand ( n242779 , n242778 , n52850 );
not ( n242780 , n242779 );
or ( n242781 , n242777 , n242780 );
not ( n242782 , n242776 );
not ( n242783 , n242779 );
nand ( n242784 , n242782 , n242783 );
nand ( n242785 , n242781 , n242784 );
xor ( n242786 , n242766 , n242785 );
not ( n242787 , n242786 );
not ( n242788 , n33812 );
buf ( n242789 , n27950 );
not ( n242790 , n242789 );
not ( n242791 , n33853 );
or ( n242792 , n242790 , n242791 );
or ( n242793 , n33853 , n242789 );
nand ( n242794 , n242792 , n242793 );
not ( n242795 , n242794 );
and ( n242796 , n242788 , n242795 );
and ( n242797 , n33812 , n242794 );
nor ( n242798 , n242796 , n242797 );
nand ( n242799 , n242798 , n52936 );
not ( n242800 , n242799 );
xor ( n242801 , n205045 , n49504 );
xnor ( n242802 , n242801 , n209844 );
not ( n242803 , n242802 );
or ( n242804 , n242800 , n242803 );
or ( n242805 , n242802 , n242799 );
nand ( n242806 , n242804 , n242805 );
not ( n242807 , n242806 );
not ( n242808 , n242807 );
not ( n242809 , n207855 );
buf ( n242810 , n30097 );
not ( n242811 , n242810 );
or ( n242812 , n242809 , n242811 );
or ( n242813 , n242810 , n207855 );
nand ( n242814 , n242812 , n242813 );
not ( n242815 , n242814 );
not ( n242816 , n53417 );
or ( n242817 , n242815 , n242816 );
not ( n242818 , n242814 );
nand ( n242819 , n242818 , n40726 );
nand ( n242820 , n242817 , n242819 );
and ( n242821 , n242820 , n54509 );
not ( n242822 , n242820 );
and ( n242823 , n242822 , n42397 );
nor ( n242824 , n242821 , n242823 );
not ( n242825 , n242824 );
nand ( n242826 , n242825 , n52966 );
not ( n242827 , n242826 );
not ( n242828 , n45293 );
not ( n242829 , n34603 );
or ( n242830 , n242828 , n242829 );
or ( n242831 , n34603 , n45293 );
nand ( n242832 , n242830 , n242831 );
and ( n242833 , n242832 , n34141 );
not ( n242834 , n242832 );
and ( n242835 , n242834 , n30638 );
nor ( n242836 , n242833 , n242835 );
not ( n242837 , n242836 );
and ( n242838 , n242827 , n242837 );
not ( n242839 , n242824 );
nand ( n242840 , n242839 , n52966 );
and ( n242841 , n242840 , n242836 );
nor ( n242842 , n242838 , n242841 );
not ( n242843 , n242842 );
not ( n242844 , n242843 );
or ( n242845 , n242808 , n242844 );
nand ( n242846 , n242842 , n242806 );
nand ( n242847 , n242845 , n242846 );
not ( n242848 , n242847 );
and ( n242849 , n242787 , n242848 );
and ( n242850 , n242786 , n242847 );
nor ( n242851 , n242849 , n242850 );
not ( n242852 , n242851 );
not ( n242853 , n242852 );
or ( n242854 , n242724 , n242853 );
and ( n242855 , n242786 , n242847 );
not ( n242856 , n242786 );
not ( n242857 , n242847 );
and ( n242858 , n242856 , n242857 );
nor ( n242859 , n242855 , n242858 );
not ( n242860 , n242859 );
or ( n242861 , n242860 , n242723 );
nand ( n242862 , n242854 , n242861 );
not ( n242863 , n242862 );
not ( n242864 , n208725 );
and ( n242865 , n242863 , n242864 );
not ( n242866 , n208725 );
not ( n242867 , n242866 );
and ( n242868 , n242862 , n242867 );
nor ( n242869 , n242865 , n242868 );
nor ( n242870 , n242703 , n242869 );
or ( n242871 , n242687 , n242870 );
nor ( n242872 , n242686 , n226003 );
nand ( n242873 , n242872 , n242870 );
nand ( n242874 , n49054 , n31507 );
nand ( n242875 , n242871 , n242873 , n242874 );
buf ( n242876 , n242875 );
not ( n242877 , RI19ac4dc0_2293);
or ( n242878 , n25328 , n242877 );
not ( n242879 , RI19abc6c0_2364);
or ( n242880 , n25335 , n242879 );
nand ( n242881 , n242878 , n242880 );
buf ( n242882 , n242881 );
not ( n242883 , RI19a9d1a8_2590);
or ( n242884 , n25328 , n242883 );
not ( n242885 , RI19a92e10_2662);
or ( n242886 , n226822 , n242885 );
nand ( n242887 , n242884 , n242886 );
buf ( n242888 , n242887 );
buf ( n242889 , n34869 );
buf ( n242890 , n52221 );
not ( n242891 , n238970 );
not ( n242892 , n51998 );
not ( n242893 , n242892 );
or ( n242894 , n242891 , n242893 );
or ( n242895 , n242892 , n238970 );
nand ( n242896 , n242894 , n242895 );
xor ( n242897 , n242890 , n242896 );
not ( n242898 , n242897 );
not ( n242899 , n242898 );
not ( n242900 , n49860 );
nand ( n242901 , n242900 , n39101 );
and ( n242902 , n242901 , n227631 );
not ( n242903 , n242901 );
and ( n242904 , n242903 , n49869 );
nor ( n242905 , n242902 , n242904 );
not ( n242906 , n242905 );
not ( n242907 , n242906 );
not ( n242908 , n227707 );
or ( n242909 , n242907 , n242908 );
not ( n242910 , n242906 );
not ( n242911 , n227706 );
nand ( n242912 , n242910 , n242911 );
nand ( n242913 , n242909 , n242912 );
nand ( n242914 , n242737 , n242734 );
not ( n242915 , n242914 );
not ( n242916 , n52880 );
and ( n242917 , n242915 , n242916 );
nand ( n242918 , n242737 , n242734 );
and ( n242919 , n242918 , n52880 );
nor ( n242920 , n242917 , n242919 );
not ( n242921 , n242920 );
not ( n242922 , n242776 );
nand ( n242923 , n242922 , n242714 );
and ( n242924 , n242923 , n230623 );
not ( n242925 , n242923 );
and ( n242926 , n242925 , n230624 );
nor ( n242927 , n242924 , n242926 );
not ( n242928 , n242927 );
or ( n242929 , n242921 , n242928 );
or ( n242930 , n242927 , n242920 );
nand ( n242931 , n242929 , n242930 );
not ( n242932 , n242752 );
nand ( n242933 , n242760 , n242932 );
not ( n242934 , n242933 );
not ( n242935 , n230572 );
or ( n242936 , n242934 , n242935 );
or ( n242937 , n230572 , n242933 );
nand ( n242938 , n242936 , n242937 );
and ( n242939 , n242931 , n242938 );
not ( n242940 , n242931 );
not ( n242941 , n242938 );
and ( n242942 , n242940 , n242941 );
nor ( n242943 , n242939 , n242942 );
not ( n242944 , n242943 );
not ( n242945 , n242836 );
nand ( n242946 , n242945 , n242824 );
not ( n242947 , n242946 );
not ( n242948 , n52949 );
and ( n242949 , n242947 , n242948 );
and ( n242950 , n242946 , n52949 );
nor ( n242951 , n242949 , n242950 );
not ( n242952 , n242951 );
or ( n242953 , n242802 , n242798 );
buf ( n242954 , n52911 );
not ( n242955 , n242954 );
and ( n242956 , n242953 , n242955 );
not ( n242957 , n242953 );
and ( n242958 , n242957 , n242954 );
nor ( n242959 , n242956 , n242958 );
not ( n242960 , n242959 );
or ( n242961 , n242952 , n242960 );
or ( n242962 , n242959 , n242951 );
nand ( n242963 , n242961 , n242962 );
not ( n242964 , n242963 );
not ( n242965 , n242964 );
or ( n242966 , n242944 , n242965 );
not ( n242967 , n242943 );
nand ( n242968 , n242967 , n242963 );
nand ( n242969 , n242966 , n242968 );
buf ( n242970 , n242969 );
and ( n242971 , n242913 , n242970 );
not ( n242972 , n242913 );
not ( n242973 , n242964 );
not ( n242974 , n242943 );
and ( n242975 , n242973 , n242974 );
and ( n242976 , n242964 , n242943 );
nor ( n242977 , n242975 , n242976 );
buf ( n242978 , n242977 );
and ( n242979 , n242972 , n242978 );
nor ( n242980 , n242971 , n242979 );
not ( n242981 , n242980 );
not ( n242982 , n242981 );
or ( n242983 , n242899 , n242982 );
not ( n242984 , n229405 );
not ( n242985 , n40144 );
and ( n242986 , n242984 , n242985 );
and ( n242987 , n229405 , n40144 );
nor ( n242988 , n242986 , n242987 );
and ( n242989 , n242988 , n38570 );
not ( n242990 , n242988 );
and ( n242991 , n242990 , n38569 );
nor ( n242992 , n242989 , n242991 );
nand ( n242993 , n242992 , n46386 );
not ( n242994 , n242993 );
not ( n242995 , n46374 );
or ( n242996 , n242994 , n242995 );
or ( n242997 , n46374 , n242993 );
nand ( n242998 , n242996 , n242997 );
not ( n242999 , n242998 );
not ( n243000 , n46420 );
or ( n243001 , n242999 , n243000 );
not ( n243002 , n242998 );
not ( n243003 , n224094 );
not ( n243004 , n46414 );
or ( n243005 , n243003 , n243004 );
nand ( n243006 , n243005 , n224179 );
nand ( n243007 , n243002 , n243006 );
nand ( n243008 , n243001 , n243007 );
not ( n243009 , n28015 );
not ( n243010 , n37580 );
or ( n243011 , n243009 , n243010 );
or ( n243012 , n37580 , n28015 );
nand ( n243013 , n243011 , n243012 );
and ( n243014 , n243013 , n236302 );
not ( n243015 , n243013 );
and ( n243016 , n243015 , n204508 );
nor ( n243017 , n243014 , n243016 );
not ( n243018 , n32661 );
not ( n243019 , n48308 );
or ( n243020 , n243018 , n243019 );
or ( n243021 , n45308 , n32661 );
nand ( n243022 , n243020 , n243021 );
and ( n243023 , n243022 , n54849 );
not ( n243024 , n243022 );
and ( n243025 , n243024 , n48317 );
nor ( n243026 , n243023 , n243025 );
or ( n243027 , n243017 , n243026 );
not ( n243028 , n243027 );
not ( n243029 , n26112 );
not ( n243030 , n45042 );
or ( n243031 , n243029 , n243030 );
or ( n243032 , n45045 , n26112 );
nand ( n243033 , n243031 , n243032 );
and ( n243034 , n243033 , n40480 );
not ( n243035 , n243033 );
and ( n243036 , n243035 , n39569 );
nor ( n243037 , n243034 , n243036 );
not ( n243038 , n243037 );
not ( n243039 , n243038 );
and ( n243040 , n243028 , n243039 );
and ( n243041 , n243027 , n243038 );
nor ( n243042 , n243040 , n243041 );
not ( n243043 , n243042 );
not ( n243044 , n243043 );
and ( n243045 , n30512 , n46587 );
not ( n243046 , n30512 );
and ( n243047 , n243046 , n230227 );
or ( n243048 , n243045 , n243047 );
and ( n243049 , n243048 , n41448 );
not ( n243050 , n243048 );
and ( n243051 , n243050 , n236734 );
nor ( n243052 , n243049 , n243051 );
not ( n243053 , n243052 );
not ( n243054 , n40780 );
not ( n243055 , n31473 );
or ( n243056 , n243054 , n243055 );
or ( n243057 , n37297 , n40780 );
nand ( n243058 , n243056 , n243057 );
and ( n243059 , n243058 , n233632 );
not ( n243060 , n243058 );
and ( n243061 , n243060 , n31515 );
nor ( n243062 , n243059 , n243061 );
not ( n243063 , n243062 );
nand ( n243064 , n243053 , n243063 );
not ( n243065 , n34151 );
not ( n243066 , n47607 );
or ( n243067 , n243065 , n243066 );
nand ( n243068 , n49132 , n34147 );
nand ( n243069 , n243067 , n243068 );
and ( n243070 , n243069 , n204860 );
not ( n243071 , n243069 );
and ( n243072 , n243071 , n49137 );
nor ( n243073 , n243070 , n243072 );
and ( n243074 , n243064 , n243073 );
not ( n243075 , n243064 );
not ( n243076 , n243073 );
and ( n243077 , n243075 , n243076 );
nor ( n243078 , n243074 , n243077 );
not ( n243079 , n243078 );
not ( n243080 , n243079 );
or ( n243081 , n243044 , n243080 );
nand ( n243082 , n243078 , n243042 );
nand ( n243083 , n243081 , n243082 );
not ( n243084 , n243083 );
not ( n243085 , n243084 );
not ( n243086 , n230239 );
not ( n243087 , n29409 );
or ( n243088 , n243086 , n243087 );
or ( n243089 , n29409 , n230239 );
nand ( n243090 , n243088 , n243089 );
xor ( n243091 , n243090 , n29454 );
not ( n243092 , n243091 );
not ( n243093 , n224642 );
not ( n243094 , n37914 );
not ( n243095 , n29213 );
or ( n243096 , n243094 , n243095 );
nand ( n243097 , n29212 , n37910 );
nand ( n243098 , n243096 , n243097 );
not ( n243099 , n243098 );
and ( n243100 , n243093 , n243099 );
and ( n243101 , n224642 , n243098 );
nor ( n243102 , n243100 , n243101 );
nand ( n243103 , n243092 , n243102 );
not ( n243104 , n243103 );
not ( n243105 , n26019 );
not ( n243106 , n29174 );
or ( n243107 , n243105 , n243106 );
nand ( n243108 , n29161 , n26015 );
nand ( n243109 , n243107 , n243108 );
not ( n243110 , n243109 );
not ( n243111 , n33936 );
and ( n243112 , n243110 , n243111 );
and ( n243113 , n243109 , n41077 );
nor ( n243114 , n243112 , n243113 );
not ( n243115 , n243114 );
not ( n243116 , n243115 );
and ( n243117 , n243104 , n243116 );
and ( n243118 , n243103 , n243115 );
nor ( n243119 , n243117 , n243118 );
not ( n243120 , n243119 );
not ( n243121 , n35827 );
not ( n243122 , n33261 );
or ( n243123 , n243121 , n243122 );
not ( n243124 , n35827 );
nand ( n243125 , n243124 , n205142 );
nand ( n243126 , n243123 , n243125 );
xor ( n243127 , n243126 , n33303 );
not ( n243128 , n39621 );
not ( n243129 , n28829 );
or ( n243130 , n243128 , n243129 );
or ( n243131 , n206591 , n39621 );
nand ( n243132 , n243130 , n243131 );
not ( n243133 , n243132 );
not ( n243134 , n32219 );
or ( n243135 , n243133 , n243134 );
or ( n243136 , n32219 , n243132 );
nand ( n243137 , n243135 , n243136 );
nand ( n243138 , n243127 , n243137 );
not ( n243139 , n30232 );
not ( n243140 , n37211 );
or ( n243141 , n243139 , n243140 );
not ( n243142 , n30232 );
nand ( n243143 , n243142 , n44966 );
nand ( n243144 , n243141 , n243143 );
and ( n243145 , n243144 , n28466 );
not ( n243146 , n243144 );
and ( n243147 , n243146 , n218203 );
nor ( n243148 , n243145 , n243147 );
not ( n243149 , n243148 );
and ( n243150 , n243138 , n243149 );
not ( n243151 , n243138 );
and ( n243152 , n243151 , n243148 );
nor ( n243153 , n243150 , n243152 );
not ( n243154 , n243153 );
or ( n243155 , n243120 , n243154 );
or ( n243156 , n243153 , n243119 );
nand ( n243157 , n243155 , n243156 );
not ( n243158 , n32906 );
not ( n243159 , n29875 );
not ( n243160 , n32898 );
or ( n243161 , n243159 , n243160 );
or ( n243162 , n32898 , n29875 );
nand ( n243163 , n243161 , n243162 );
not ( n243164 , n243163 );
or ( n243165 , n243158 , n243164 );
or ( n243166 , n243163 , n32909 );
nand ( n243167 , n243165 , n243166 );
not ( n243168 , n243167 );
xor ( n243169 , n41128 , n51954 );
xnor ( n243170 , n243169 , n225948 );
not ( n243171 , n243170 );
nand ( n243172 , n243168 , n243171 );
not ( n243173 , n41710 );
not ( n243174 , n28146 );
or ( n243175 , n243173 , n243174 );
not ( n243176 , n41710 );
nand ( n243177 , n243176 , n44712 );
nand ( n243178 , n243175 , n243177 );
and ( n243179 , n243178 , n35275 );
not ( n243180 , n243178 );
and ( n243181 , n243180 , n44720 );
nor ( n243182 , n243179 , n243181 );
and ( n243183 , n243172 , n243182 );
not ( n243184 , n243172 );
not ( n243185 , n243182 );
and ( n243186 , n243184 , n243185 );
nor ( n243187 , n243183 , n243186 );
and ( n243188 , n243157 , n243187 );
not ( n243189 , n243157 );
not ( n243190 , n243187 );
and ( n243191 , n243189 , n243190 );
nor ( n243192 , n243188 , n243191 );
not ( n243193 , n243192 );
or ( n243194 , n243085 , n243193 );
not ( n243195 , n243192 );
nand ( n243196 , n243195 , n243083 );
nand ( n243197 , n243194 , n243196 );
buf ( n243198 , n243197 );
not ( n243199 , n243198 );
and ( n243200 , n243008 , n243199 );
not ( n243201 , n243008 );
and ( n243202 , n243201 , n243198 );
nor ( n243203 , n243200 , n243202 );
not ( n243204 , n226010 );
nor ( n243205 , n243203 , n243204 );
nand ( n243206 , n242983 , n243205 );
nor ( n243207 , n242897 , n243204 );
nand ( n243208 , n243203 , n243207 , n242981 );
nand ( n243209 , n39767 , n27918 );
nand ( n243210 , n243206 , n243208 , n243209 );
buf ( n243211 , n243210 );
buf ( n243212 , n32266 );
buf ( n243213 , n36614 );
not ( n243214 , n42837 );
not ( n243215 , n237699 );
not ( n243216 , n243215 );
or ( n243217 , n243214 , n243216 );
not ( n243218 , n42837 );
nand ( n243219 , n237695 , n237671 );
not ( n243220 , n237695 );
nand ( n243221 , n243220 , n237670 );
nand ( n243222 , n243219 , n243221 );
nand ( n243223 , n243218 , n243222 );
nand ( n243224 , n243217 , n243223 );
not ( n243225 , n48875 );
not ( n243226 , n243225 );
and ( n243227 , n243224 , n243226 );
not ( n243228 , n243224 );
not ( n243229 , n48883 );
not ( n243230 , n243229 );
and ( n243231 , n243228 , n243230 );
nor ( n243232 , n243227 , n243231 );
not ( n243233 , n47173 );
nand ( n243234 , n243232 , n243233 );
not ( n243235 , n243234 );
not ( n243236 , n241092 );
not ( n243237 , n235580 );
or ( n243238 , n243236 , n243237 );
nand ( n243239 , n235590 , n241095 );
nand ( n243240 , n243238 , n243239 );
and ( n243241 , n243240 , n235720 );
not ( n243242 , n243240 );
not ( n243243 , n235728 );
not ( n243244 , n243243 );
and ( n243245 , n243242 , n243244 );
nor ( n243246 , n243241 , n243245 );
not ( n243247 , n243246 );
and ( n243248 , n243235 , n243247 );
and ( n243249 , n31577 , n35877 );
nor ( n243250 , n243248 , n243249 );
nor ( n243251 , n243246 , n235732 );
nand ( n243252 , n229194 , n36081 );
and ( n243253 , n243252 , n35929 );
not ( n243254 , n243252 );
and ( n243255 , n243254 , n35928 );
nor ( n243256 , n243253 , n243255 );
not ( n243257 , n243256 );
not ( n243258 , n243257 );
not ( n243259 , n229300 );
or ( n243260 , n243258 , n243259 );
not ( n243261 , n243257 );
nand ( n243262 , n243261 , n51549 );
nand ( n243263 , n243260 , n243262 );
and ( n243264 , n243263 , n51598 );
not ( n243265 , n243263 );
and ( n243266 , n243265 , n51607 );
nor ( n243267 , n243264 , n243266 );
nand ( n243268 , n243251 , n243267 );
not ( n243269 , n243267 );
nor ( n243270 , n243232 , n33254 );
nand ( n243271 , n243269 , n243246 , n243270 );
nand ( n243272 , n243250 , n243268 , n243271 );
buf ( n243273 , n243272 );
not ( n243274 , n48583 );
not ( n243275 , n243274 );
not ( n243276 , n234420 );
or ( n243277 , n243275 , n243276 );
not ( n243278 , n243274 );
nand ( n243279 , n243278 , n239119 );
nand ( n243280 , n243277 , n243279 );
and ( n243281 , n243280 , n239229 );
not ( n243282 , n243280 );
and ( n243283 , n243282 , n239221 );
nor ( n243284 , n243281 , n243283 );
not ( n243285 , n241618 );
not ( n243286 , n243285 );
nand ( n243287 , n241490 , n241508 );
not ( n243288 , n243287 );
buf ( n243289 , n28635 );
not ( n243290 , n243289 );
not ( n243291 , n230437 );
or ( n243292 , n243290 , n243291 );
or ( n243293 , n230437 , n243289 );
nand ( n243294 , n243292 , n243293 );
not ( n243295 , n33756 );
and ( n243296 , n243294 , n243295 );
not ( n243297 , n243294 );
and ( n243298 , n243297 , n33760 );
nor ( n243299 , n243296 , n243298 );
not ( n243300 , n243299 );
and ( n243301 , n243288 , n243300 );
and ( n243302 , n243287 , n243299 );
nor ( n243303 , n243301 , n243302 );
not ( n243304 , n243303 );
nand ( n243305 , n241550 , n241534 );
not ( n243306 , n39303 );
not ( n243307 , n205033 );
not ( n243308 , n243307 );
or ( n243309 , n243306 , n243308 );
not ( n243310 , n39303 );
nand ( n243311 , n243310 , n205033 );
nand ( n243312 , n243309 , n243311 );
and ( n243313 , n243312 , n205074 );
not ( n243314 , n243312 );
and ( n243315 , n243314 , n221787 );
nor ( n243316 , n243313 , n243315 );
not ( n243317 , n243316 );
and ( n243318 , n243305 , n243317 );
not ( n243319 , n243305 );
and ( n243320 , n243319 , n243316 );
nor ( n243321 , n243318 , n243320 );
not ( n243322 , n243321 );
or ( n243323 , n243304 , n243322 );
or ( n243324 , n243321 , n243303 );
nand ( n243325 , n243323 , n243324 );
nand ( n243326 , n241558 , n241579 );
and ( n243327 , n243326 , n242428 );
not ( n243328 , n243326 );
not ( n243329 , n242428 );
and ( n243330 , n243328 , n243329 );
nor ( n243331 , n243327 , n243330 );
xnor ( n243332 , n243325 , n243331 );
not ( n243333 , n243332 );
not ( n243334 , n243333 );
buf ( n243335 , n27990 );
not ( n243336 , n243335 );
not ( n243337 , n41319 );
or ( n243338 , n243336 , n243337 );
or ( n243339 , n41319 , n243335 );
nand ( n243340 , n243338 , n243339 );
xor ( n243341 , n243340 , n41360 );
not ( n243342 , n243341 );
not ( n243343 , n243342 );
nand ( n243344 , n241630 , n241643 );
not ( n243345 , n243344 );
or ( n243346 , n243343 , n243345 );
or ( n243347 , n243344 , n243342 );
nand ( n243348 , n243346 , n243347 );
xor ( n243349 , n29517 , n43201 );
xnor ( n243350 , n243349 , n216225 );
not ( n243351 , n243350 );
not ( n243352 , n243351 );
nand ( n243353 , n241613 , n241590 );
not ( n243354 , n243353 );
and ( n243355 , n243352 , n243354 );
and ( n243356 , n243353 , n243351 );
nor ( n243357 , n243355 , n243356 );
xor ( n243358 , n243348 , n243357 );
not ( n243359 , n243358 );
not ( n243360 , n243359 );
and ( n243361 , n243334 , n243360 );
and ( n243362 , n243333 , n243359 );
nor ( n243363 , n243361 , n243362 );
not ( n243364 , n243363 );
or ( n243365 , n243286 , n243364 );
not ( n243366 , n243285 );
not ( n243367 , n243358 );
not ( n243368 , n243332 );
or ( n243369 , n243367 , n243368 );
not ( n243370 , n243358 );
nand ( n243371 , n243370 , n243333 );
nand ( n243372 , n243369 , n243371 );
nand ( n243373 , n243366 , n243372 );
nand ( n243374 , n243365 , n243373 );
not ( n243375 , n38791 );
nand ( n243376 , n243375 , n49657 );
not ( n243377 , n243376 );
not ( n243378 , n38777 );
and ( n243379 , n243377 , n243378 );
and ( n243380 , n243376 , n38777 );
nor ( n243381 , n243379 , n243380 );
not ( n243382 , n243381 );
not ( n243383 , n49714 );
nand ( n243384 , n243383 , n38850 );
and ( n243385 , n243384 , n38833 );
not ( n243386 , n243384 );
and ( n243387 , n243386 , n38832 );
nor ( n243388 , n243385 , n243387 );
not ( n243389 , n243388 );
or ( n243390 , n243382 , n243389 );
or ( n243391 , n243388 , n243381 );
nand ( n243392 , n243390 , n243391 );
nand ( n243393 , n242552 , n227460 );
and ( n243394 , n243393 , n38726 );
not ( n243395 , n243393 );
not ( n243396 , n38726 );
and ( n243397 , n243395 , n243396 );
or ( n243398 , n243394 , n243397 );
and ( n243399 , n243392 , n243398 );
not ( n243400 , n243392 );
not ( n243401 , n243398 );
and ( n243402 , n243400 , n243401 );
nor ( n243403 , n243399 , n243402 );
not ( n243404 , n234530 );
not ( n243405 , n38716 );
not ( n243406 , n243405 );
or ( n243407 , n243404 , n243406 );
not ( n243408 , n234530 );
nand ( n243409 , n243408 , n38716 );
nand ( n243410 , n243407 , n243409 );
and ( n243411 , n243403 , n243410 );
not ( n243412 , n243403 );
not ( n243413 , n243410 );
and ( n243414 , n243412 , n243413 );
nor ( n243415 , n243411 , n243414 );
buf ( n243416 , n243415 );
xor ( n243417 , n243374 , n243416 );
nand ( n243418 , n243284 , n243417 );
not ( n243419 , n243418 );
not ( n243420 , n38578 );
not ( n243421 , n234513 );
or ( n243422 , n243420 , n243421 );
not ( n243423 , n38578 );
nand ( n243424 , n243423 , n234521 );
nand ( n243425 , n243422 , n243424 );
not ( n243426 , n223266 );
not ( n243427 , n243426 );
and ( n243428 , n243425 , n243427 );
not ( n243429 , n243425 );
buf ( n243430 , n223266 );
not ( n243431 , n243430 );
and ( n243432 , n243429 , n243431 );
nor ( n243433 , n243428 , n243432 );
buf ( n243434 , n33252 );
nor ( n243435 , n243433 , n243434 );
not ( n243436 , n243435 );
or ( n243437 , n243419 , n243436 );
not ( n243438 , n233971 );
nand ( n243439 , n243433 , n243438 );
or ( n243440 , n243439 , n243418 );
nand ( n243441 , n239240 , n30372 );
nand ( n243442 , n243437 , n243440 , n243441 );
buf ( n243443 , n243442 );
not ( n243444 , n41558 );
not ( n243445 , n243444 );
not ( n243446 , n233026 );
or ( n243447 , n243445 , n243446 );
not ( n243448 , n243444 );
nand ( n243449 , n243448 , n233035 );
nand ( n243450 , n243447 , n243449 );
and ( n243451 , n243450 , n233084 );
not ( n243452 , n243450 );
and ( n243453 , n243452 , n233091 );
nor ( n243454 , n243451 , n243453 );
nand ( n243455 , n243454 , n239934 );
not ( n243456 , n238720 );
nand ( n243457 , n243456 , n238707 );
and ( n243458 , n243457 , n230103 );
not ( n243459 , n243457 );
and ( n243460 , n243459 , n52343 );
nor ( n243461 , n243458 , n243460 );
not ( n243462 , n243461 );
not ( n243463 , n239930 );
or ( n243464 , n243462 , n243463 );
not ( n243465 , n243461 );
nand ( n243466 , n243465 , n239922 );
nand ( n243467 , n243464 , n243466 );
not ( n243468 , n238810 );
not ( n243469 , n236576 );
nand ( n243470 , n243468 , n243469 );
not ( n243471 , n243470 );
not ( n243472 , n221107 );
and ( n243473 , n243471 , n243472 );
and ( n243474 , n243470 , n221107 );
nor ( n243475 , n243473 , n243474 );
not ( n243476 , n243475 );
not ( n243477 , n43266 );
nand ( n243478 , n243477 , n238827 );
buf ( n243479 , n43281 );
and ( n243480 , n243478 , n243479 );
not ( n243481 , n243478 );
not ( n243482 , n243479 );
and ( n243483 , n243481 , n243482 );
nor ( n243484 , n243480 , n243483 );
not ( n243485 , n243484 );
or ( n243486 , n243476 , n243485 );
or ( n243487 , n243484 , n243475 );
nand ( n243488 , n243486 , n243487 );
not ( n243489 , n242692 );
and ( n243490 , n243488 , n243489 );
not ( n243491 , n243488 );
and ( n243492 , n243491 , n242692 );
nor ( n243493 , n243490 , n243492 );
not ( n243494 , n236638 );
not ( n243495 , n241194 );
or ( n243496 , n243494 , n243495 );
nand ( n243497 , n241193 , n236567 );
nand ( n243498 , n243496 , n243497 );
not ( n243499 , n243498 );
and ( n243500 , n243493 , n243499 );
not ( n243501 , n243493 );
and ( n243502 , n243501 , n243498 );
nor ( n243503 , n243500 , n243502 );
buf ( n243504 , n243503 );
and ( n243505 , n243467 , n243504 );
not ( n243506 , n243467 );
and ( n243507 , n243493 , n243498 );
not ( n243508 , n243493 );
and ( n243509 , n243508 , n243499 );
nor ( n243510 , n243507 , n243509 );
buf ( n243511 , n243510 );
and ( n243512 , n243506 , n243511 );
nor ( n243513 , n243505 , n243512 );
not ( n243514 , n243513 );
not ( n243515 , n54164 );
not ( n243516 , n242380 );
or ( n243517 , n243515 , n243516 );
not ( n243518 , n54164 );
nand ( n243519 , n243518 , n242373 );
nand ( n243520 , n243517 , n243519 );
not ( n243521 , n32961 );
not ( n243522 , n28685 );
and ( n243523 , n243521 , n243522 );
and ( n243524 , n32961 , n28685 );
nor ( n243525 , n243523 , n243524 );
and ( n243526 , n243525 , n32989 );
not ( n243527 , n243525 );
and ( n243528 , n243527 , n54623 );
nor ( n243529 , n243526 , n243528 );
buf ( n243530 , n243529 );
not ( n243531 , n243530 );
xor ( n243532 , n28982 , n209033 );
xnor ( n243533 , n243532 , n35169 );
nand ( n243534 , n243533 , n223967 );
not ( n243535 , n243534 );
or ( n243536 , n243531 , n243535 );
or ( n243537 , n243534 , n243530 );
nand ( n243538 , n243536 , n243537 );
not ( n243539 , n243538 );
not ( n243540 , n41237 );
not ( n243541 , n33443 );
or ( n243542 , n243540 , n243541 );
or ( n243543 , n33443 , n41237 );
nand ( n243544 , n243542 , n243543 );
and ( n243545 , n243544 , n40776 );
not ( n243546 , n243544 );
and ( n243547 , n243546 , n33475 );
nor ( n243548 , n243545 , n243547 );
nand ( n243549 , n224024 , n243548 );
not ( n243550 , n243549 );
not ( n243551 , n36982 );
nand ( n243552 , n25963 , n41322 );
not ( n243553 , n243552 );
nor ( n243554 , n25963 , n41322 );
nor ( n243555 , n243553 , n243554 );
not ( n243556 , n243555 );
or ( n243557 , n243551 , n243556 );
or ( n243558 , n53925 , n243555 );
nand ( n243559 , n243557 , n243558 );
not ( n243560 , n243559 );
and ( n243561 , n243550 , n243560 );
not ( n243562 , n243548 );
not ( n243563 , n243562 );
nand ( n243564 , n243563 , n224024 );
and ( n243565 , n243564 , n243559 );
nor ( n243566 , n243561 , n243565 );
not ( n243567 , n243566 );
or ( n243568 , n243539 , n243567 );
or ( n243569 , n243566 , n243538 );
nand ( n243570 , n243568 , n243569 );
not ( n243571 , n45702 );
not ( n243572 , n34849 );
not ( n243573 , n55591 );
or ( n243574 , n243572 , n243573 );
or ( n243575 , n239577 , n34849 );
nand ( n243576 , n243574 , n243575 );
not ( n243577 , n243576 );
or ( n243578 , n243571 , n243577 );
or ( n243579 , n243576 , n41593 );
nand ( n243580 , n243578 , n243579 );
not ( n243581 , n243580 );
nand ( n243582 , n224085 , n243581 );
not ( n243583 , n32863 );
not ( n243584 , n206190 );
not ( n243585 , n34339 );
or ( n243586 , n243584 , n243585 );
or ( n243587 , n34339 , n206190 );
nand ( n243588 , n243586 , n243587 );
not ( n243589 , n243588 );
and ( n243590 , n243583 , n243589 );
and ( n243591 , n32863 , n243588 );
nor ( n243592 , n243590 , n243591 );
and ( n243593 , n243582 , n243592 );
not ( n243594 , n243582 );
not ( n243595 , n243592 );
and ( n243596 , n243594 , n243595 );
nor ( n243597 , n243593 , n243596 );
not ( n243598 , n243597 );
and ( n243599 , n243570 , n243598 );
not ( n243600 , n243570 );
and ( n243601 , n243600 , n243597 );
nor ( n243602 , n243599 , n243601 );
not ( n243603 , n242992 );
not ( n243604 , n28665 );
not ( n243605 , n29622 );
not ( n243606 , n43469 );
or ( n243607 , n243605 , n243606 );
or ( n243608 , n223166 , n29622 );
nand ( n243609 , n243607 , n243608 );
not ( n243610 , n243609 );
or ( n243611 , n243604 , n243610 );
or ( n243612 , n243609 , n28665 );
nand ( n243613 , n243611 , n243612 );
not ( n243614 , n243613 );
nand ( n243615 , n46404 , n243614 );
not ( n243616 , n243615 );
or ( n243617 , n243603 , n243616 );
or ( n243618 , n243615 , n242992 );
nand ( n243619 , n243617 , n243618 );
not ( n243620 , n243619 );
not ( n243621 , n33828 );
not ( n243622 , n38795 );
or ( n243623 , n243621 , n243622 );
not ( n243624 , n33828 );
nand ( n243625 , n243624 , n37193 );
nand ( n243626 , n243623 , n243625 );
and ( n243627 , n243626 , n237226 );
not ( n243628 , n243626 );
and ( n243629 , n243628 , n38801 );
nor ( n243630 , n243627 , n243629 );
not ( n243631 , n243630 );
nand ( n243632 , n46340 , n243631 );
not ( n243633 , n243632 );
buf ( n243634 , RI1740ac80_1455);
not ( n243635 , n243634 );
not ( n243636 , n44932 );
or ( n243637 , n243635 , n243636 );
or ( n243638 , n44932 , n243634 );
nand ( n243639 , n243637 , n243638 );
not ( n243640 , n243639 );
not ( n243641 , n222667 );
and ( n243642 , n243640 , n243641 );
and ( n243643 , n243639 , n222700 );
nor ( n243644 , n243642 , n243643 );
not ( n243645 , n243644 );
not ( n243646 , n243645 );
and ( n243647 , n243633 , n243646 );
and ( n243648 , n243632 , n243645 );
nor ( n243649 , n243647 , n243648 );
not ( n243650 , n243649 );
or ( n243651 , n243620 , n243650 );
or ( n243652 , n243649 , n243619 );
nand ( n243653 , n243651 , n243652 );
not ( n243654 , n243653 );
and ( n243655 , n243602 , n243654 );
not ( n243656 , n243602 );
and ( n243657 , n243656 , n243653 );
nor ( n243658 , n243655 , n243657 );
buf ( n243659 , n243658 );
not ( n243660 , n243659 );
and ( n243661 , n243520 , n243660 );
not ( n243662 , n243520 );
and ( n243663 , n243662 , n243659 );
nor ( n243664 , n243661 , n243663 );
nand ( n243665 , n243514 , n243664 );
or ( n243666 , n243455 , n243665 );
not ( n243667 , n243513 );
not ( n243668 , n243667 );
not ( n243669 , n243454 );
or ( n243670 , n243668 , n243669 );
nor ( n243671 , n243664 , n233972 );
nand ( n243672 , n243670 , n243671 );
nand ( n243673 , n35431 , n29764 );
nand ( n243674 , n243666 , n243672 , n243673 );
buf ( n243675 , n243674 );
nand ( n243676 , n48283 , n48297 );
not ( n243677 , n243676 );
not ( n243678 , n47407 );
and ( n243679 , n243677 , n243678 );
and ( n243680 , n243676 , n47407 );
nor ( n243681 , n243679 , n243680 );
not ( n243682 , n243681 );
not ( n243683 , n243682 );
not ( n243684 , n241428 );
not ( n243685 , n241444 );
or ( n243686 , n243684 , n243685 );
nand ( n243687 , n243686 , n241447 );
not ( n243688 , n243687 );
not ( n243689 , n243688 );
or ( n243690 , n243683 , n243689 );
not ( n243691 , n243682 );
nand ( n243692 , n243691 , n243687 );
nand ( n243693 , n243690 , n243692 );
and ( n243694 , n243693 , n241453 );
not ( n243695 , n243693 );
and ( n243696 , n243695 , n236781 );
nor ( n243697 , n243694 , n243696 );
not ( n243698 , n243697 );
not ( n243699 , n30235 );
not ( n243700 , n37212 );
or ( n243701 , n243699 , n243700 );
nand ( n243702 , n44966 , n30230 );
nand ( n243703 , n243701 , n243702 );
not ( n243704 , n243703 );
not ( n243705 , n218203 );
and ( n243706 , n243704 , n243705 );
and ( n243707 , n243703 , n218203 );
nor ( n243708 , n243706 , n243707 );
nand ( n243709 , n43205 , n243708 );
and ( n243710 , n243709 , n236745 );
not ( n243711 , n243709 );
and ( n243712 , n243711 , n236746 );
nor ( n243713 , n243710 , n243712 );
not ( n243714 , n243713 );
not ( n243715 , n29699 );
not ( n243716 , n34699 );
or ( n243717 , n243715 , n243716 );
or ( n243718 , n34699 , n29699 );
nand ( n243719 , n243717 , n243718 );
and ( n243720 , n243719 , n39845 );
not ( n243721 , n243719 );
and ( n243722 , n243721 , n44823 );
nor ( n243723 , n243720 , n243722 );
not ( n243724 , n243723 );
nand ( n243725 , n243724 , n236658 );
not ( n243726 , n243725 );
not ( n243727 , n43051 );
and ( n243728 , n243726 , n243727 );
and ( n243729 , n243725 , n43051 );
nor ( n243730 , n243728 , n243729 );
not ( n243731 , n243730 );
not ( n243732 , n236680 );
not ( n243733 , n28561 );
not ( n243734 , n43885 );
or ( n243735 , n243733 , n243734 );
or ( n243736 , n43885 , n28561 );
nand ( n243737 , n243735 , n243736 );
not ( n243738 , n243737 );
not ( n243739 , n243738 );
not ( n243740 , n30809 );
or ( n243741 , n243739 , n243740 );
nand ( n243742 , n30810 , n243737 );
nand ( n243743 , n243741 , n243742 );
nand ( n243744 , n243732 , n243743 );
and ( n243745 , n243744 , n236681 );
not ( n243746 , n243744 );
and ( n243747 , n243746 , n43086 );
nor ( n243748 , n243745 , n243747 );
not ( n243749 , n243748 );
or ( n243750 , n243731 , n243749 );
or ( n243751 , n243748 , n243730 );
nand ( n243752 , n243750 , n243751 );
not ( n243753 , n38097 );
not ( n243754 , n39417 );
or ( n243755 , n243753 , n243754 );
not ( n243756 , n38097 );
nand ( n243757 , n243756 , n32688 );
nand ( n243758 , n243755 , n243757 );
not ( n243759 , n243758 );
not ( n243760 , n47939 );
and ( n243761 , n243759 , n243760 );
and ( n243762 , n243758 , n47939 );
nor ( n243763 , n243761 , n243762 );
not ( n243764 , n243763 );
not ( n243765 , n236701 );
nand ( n243766 , n243764 , n243765 );
buf ( n243767 , n43119 );
not ( n243768 , n243767 );
and ( n243769 , n243766 , n243768 );
not ( n243770 , n243766 );
and ( n243771 , n243770 , n243767 );
nor ( n243772 , n243769 , n243771 );
xor ( n243773 , n243752 , n243772 );
not ( n243774 , n243773 );
not ( n243775 , n243774 );
not ( n243776 , n43187 );
not ( n243777 , n243708 );
nand ( n243778 , n236745 , n243777 );
not ( n243779 , n243778 );
and ( n243780 , n243776 , n243779 );
and ( n243781 , n43187 , n243778 );
nor ( n243782 , n243780 , n243781 );
not ( n243783 , n243782 );
not ( n243784 , n243783 );
xor ( n243785 , n26438 , n44471 );
xnor ( n243786 , n243785 , n31730 );
not ( n243787 , n243786 );
nand ( n243788 , n243787 , n236725 );
and ( n243789 , n243788 , n236715 );
not ( n243790 , n243788 );
and ( n243791 , n243790 , n43162 );
nor ( n243792 , n243789 , n243791 );
not ( n243793 , n243792 );
not ( n243794 , n243793 );
or ( n243795 , n243784 , n243794 );
nand ( n243796 , n243792 , n243782 );
nand ( n243797 , n243795 , n243796 );
not ( n243798 , n243797 );
and ( n243799 , n243775 , n243798 );
and ( n243800 , n243774 , n243797 );
nor ( n243801 , n243799 , n243800 );
not ( n243802 , n243801 );
or ( n243803 , n243714 , n243802 );
not ( n243804 , n243713 );
not ( n243805 , n243773 );
not ( n243806 , n243797 );
not ( n243807 , n243806 );
or ( n243808 , n243805 , n243807 );
nand ( n243809 , n243774 , n243797 );
nand ( n243810 , n243808 , n243809 );
nand ( n243811 , n243804 , n243810 );
nand ( n243812 , n243803 , n243811 );
not ( n243813 , n44800 );
not ( n243814 , n31248 );
not ( n243815 , n31251 );
or ( n243816 , n243814 , n243815 );
or ( n243817 , n31251 , n31248 );
nand ( n243818 , n243816 , n243817 );
not ( n243819 , n243818 );
nor ( n243820 , n243819 , n34820 );
not ( n243821 , n243820 );
not ( n243822 , n243818 );
nand ( n243823 , n243822 , n34820 );
nand ( n243824 , n243821 , n243823 );
and ( n243825 , n243824 , n47135 );
not ( n243826 , n243824 );
and ( n243827 , n243826 , n29336 );
nor ( n243828 , n243825 , n243827 );
nand ( n243829 , n243813 , n243828 );
not ( n243830 , n243829 );
buf ( n243831 , n44790 );
not ( n243832 , n243831 );
and ( n243833 , n243830 , n243832 );
and ( n243834 , n243829 , n243831 );
nor ( n243835 , n243833 , n243834 );
buf ( n243836 , n31206 );
not ( n243837 , n243836 );
not ( n243838 , n31425 );
or ( n243839 , n243837 , n243838 );
or ( n243840 , n31425 , n243836 );
nand ( n243841 , n243839 , n243840 );
not ( n243842 , n243841 );
not ( n243843 , n42285 );
and ( n243844 , n243842 , n243843 );
and ( n243845 , n243841 , n42285 );
nor ( n243846 , n243844 , n243845 );
not ( n243847 , n243846 );
nand ( n243848 , n237957 , n243847 );
and ( n243849 , n243848 , n44997 );
not ( n243850 , n243848 );
and ( n243851 , n243850 , n44998 );
nor ( n243852 , n243849 , n243851 );
and ( n243853 , n243835 , n243852 );
not ( n243854 , n243835 );
not ( n243855 , n243852 );
and ( n243856 , n243854 , n243855 );
nor ( n243857 , n243853 , n243856 );
not ( n243858 , n243857 );
not ( n243859 , n29006 );
buf ( n243860 , n35155 );
not ( n243861 , n243860 );
and ( n243862 , n243859 , n243861 );
and ( n243863 , n29006 , n243860 );
nor ( n243864 , n243862 , n243863 );
xor ( n243865 , n28968 , n243864 );
not ( n243866 , n243865 );
not ( n243867 , n26301 );
not ( n243868 , n38971 );
or ( n243869 , n243867 , n243868 );
not ( n243870 , n26301 );
nand ( n243871 , n243870 , n219976 );
nand ( n243872 , n243869 , n243871 );
and ( n243873 , n243872 , n39007 );
not ( n243874 , n243872 );
and ( n243875 , n243874 , n39002 );
nor ( n243876 , n243873 , n243875 );
nand ( n243877 , n243866 , n243876 );
not ( n243878 , n243877 );
not ( n243879 , n44879 );
and ( n243880 , n243878 , n243879 );
and ( n243881 , n243877 , n44879 );
nor ( n243882 , n243880 , n243881 );
not ( n243883 , n243882 );
not ( n243884 , n41043 );
not ( n243885 , n35722 );
or ( n243886 , n243884 , n243885 );
or ( n243887 , n35722 , n41043 );
nand ( n243888 , n243886 , n243887 );
and ( n243889 , n243888 , n34191 );
not ( n243890 , n243888 );
and ( n243891 , n243890 , n211419 );
nor ( n243892 , n243889 , n243891 );
not ( n243893 , n243892 );
not ( n243894 , n31213 );
buf ( n243895 , n40893 );
not ( n243896 , n243895 );
not ( n243897 , n220726 );
or ( n243898 , n243896 , n243897 );
or ( n243899 , n220726 , n243895 );
nand ( n243900 , n243898 , n243899 );
not ( n243901 , n243900 );
or ( n243902 , n243894 , n243901 );
or ( n243903 , n243900 , n31213 );
nand ( n243904 , n243902 , n243903 );
nand ( n243905 , n243893 , n243904 );
and ( n243906 , n243905 , n222599 );
not ( n243907 , n243905 );
and ( n243908 , n243907 , n222600 );
nor ( n243909 , n243906 , n243908 );
not ( n243910 , n243909 );
or ( n243911 , n243883 , n243910 );
or ( n243912 , n243909 , n243882 );
nand ( n243913 , n243911 , n243912 );
not ( n243914 , n204794 );
not ( n243915 , n205068 );
or ( n243916 , n243914 , n243915 );
not ( n243917 , n204794 );
nand ( n243918 , n243917 , n205072 );
nand ( n243919 , n243916 , n243918 );
and ( n243920 , n243919 , n43757 );
not ( n243921 , n243919 );
and ( n243922 , n243921 , n48461 );
nor ( n243923 , n243920 , n243922 );
not ( n243924 , n243923 );
buf ( n243925 , n204974 );
not ( n243926 , n243925 );
not ( n243927 , n213777 );
or ( n243928 , n243926 , n243927 );
not ( n243929 , n243925 );
nand ( n243930 , n243929 , n36024 );
nand ( n243931 , n243928 , n243930 );
and ( n243932 , n243931 , n221434 );
not ( n243933 , n243931 );
and ( n243934 , n243933 , n40862 );
nor ( n243935 , n243932 , n243934 );
not ( n243936 , n243935 );
nand ( n243937 , n243924 , n243936 );
not ( n243938 , n243937 );
not ( n243939 , n44947 );
or ( n243940 , n243938 , n243939 );
or ( n243941 , n44947 , n243937 );
nand ( n243942 , n243940 , n243941 );
and ( n243943 , n243913 , n243942 );
not ( n243944 , n243913 );
not ( n243945 , n243942 );
and ( n243946 , n243944 , n243945 );
nor ( n243947 , n243943 , n243946 );
not ( n243948 , n243947 );
or ( n243949 , n243858 , n243948 );
not ( n243950 , n243947 );
not ( n243951 , n243857 );
nand ( n243952 , n243950 , n243951 );
nand ( n243953 , n243949 , n243952 );
buf ( n243954 , n243953 );
and ( n243955 , n243812 , n243954 );
not ( n243956 , n243812 );
buf ( n243957 , n243947 );
buf ( n243958 , n243857 );
xor ( n243959 , n243957 , n243958 );
buf ( n243960 , n243959 );
and ( n243961 , n243956 , n243960 );
nor ( n243962 , n243955 , n243961 );
not ( n243963 , n243962 );
nor ( n243964 , n243698 , n243963 );
not ( n243965 , n243964 );
buf ( n243966 , n44901 );
not ( n243967 , n243966 );
not ( n243968 , n44869 );
nand ( n243969 , n243968 , n44896 );
buf ( n243970 , n243865 );
xor ( n243971 , n243969 , n243970 );
not ( n243972 , n243904 );
nand ( n243973 , n44848 , n222586 );
not ( n243974 , n243973 );
and ( n243975 , n243972 , n243974 );
and ( n243976 , n243904 , n243973 );
nor ( n243977 , n243975 , n243976 );
not ( n243978 , n243977 );
not ( n243979 , n243978 );
nand ( n243980 , n44958 , n44941 );
and ( n243981 , n243980 , n243935 );
not ( n243982 , n243980 );
and ( n243983 , n243982 , n243936 );
nor ( n243984 , n243981 , n243983 );
not ( n243985 , n243984 );
not ( n243986 , n243985 );
or ( n243987 , n243979 , n243986 );
nand ( n243988 , n243984 , n243977 );
nand ( n243989 , n243987 , n243988 );
xor ( n243990 , n243971 , n243989 );
not ( n243991 , n44809 );
nand ( n243992 , n243991 , n45008 );
not ( n243993 , n243992 );
not ( n243994 , n243828 );
and ( n243995 , n243993 , n243994 );
and ( n243996 , n243992 , n243828 );
nor ( n243997 , n243995 , n243996 );
not ( n243998 , n243997 );
nand ( n243999 , n222729 , n44981 );
and ( n244000 , n243999 , n243846 );
not ( n244001 , n243999 );
and ( n244002 , n244001 , n243847 );
nor ( n244003 , n244000 , n244002 );
not ( n244004 , n244003 );
or ( n244005 , n243998 , n244004 );
or ( n244006 , n244003 , n243997 );
nand ( n244007 , n244005 , n244006 );
xnor ( n244008 , n243990 , n244007 );
not ( n244009 , n244008 );
not ( n244010 , n244009 );
or ( n244011 , n243967 , n244010 );
or ( n244012 , n244009 , n243966 );
nand ( n244013 , n244011 , n244012 );
not ( n244014 , n244013 );
not ( n244015 , n237920 );
nand ( n244016 , n45141 , n45127 );
not ( n244017 , n244016 );
or ( n244018 , n244015 , n244017 );
or ( n244019 , n244016 , n237920 );
nand ( n244020 , n244018 , n244019 );
not ( n244021 , n244020 );
not ( n244022 , n222930 );
nand ( n244023 , n45175 , n244022 );
not ( n244024 , n244023 );
not ( n244025 , n232582 );
not ( n244026 , n244025 );
and ( n244027 , n244024 , n244026 );
and ( n244028 , n244023 , n244025 );
nor ( n244029 , n244027 , n244028 );
not ( n244030 , n244029 );
or ( n244031 , n244021 , n244030 );
or ( n244032 , n244029 , n244020 );
nand ( n244033 , n244031 , n244032 );
nand ( n244034 , n45241 , n222981 );
and ( n244035 , n244034 , n54854 );
not ( n244036 , n244034 );
and ( n244037 , n244036 , n54853 );
nor ( n244038 , n244035 , n244037 );
not ( n244039 , n244038 );
and ( n244040 , n244033 , n244039 );
not ( n244041 , n244033 );
and ( n244042 , n244041 , n244038 );
nor ( n244043 , n244040 , n244042 );
not ( n244044 , n244043 );
not ( n244045 , n240065 );
not ( n244046 , n232543 );
or ( n244047 , n244045 , n244046 );
or ( n244048 , n232543 , n240065 );
nand ( n244049 , n244047 , n244048 );
not ( n244050 , n244049 );
and ( n244051 , n244044 , n244050 );
not ( n244052 , n244044 );
and ( n244053 , n244052 , n244049 );
nor ( n244054 , n244051 , n244053 );
not ( n244055 , n244054 );
not ( n244056 , n244055 );
not ( n244057 , n244056 );
and ( n244058 , n244014 , n244057 );
and ( n244059 , n244013 , n244056 );
nor ( n244060 , n244058 , n244059 );
not ( n244061 , n244060 );
nor ( n244062 , n244061 , n238900 );
not ( n244063 , n244062 );
or ( n244064 , n243965 , n244063 );
nand ( n244065 , n244060 , n243962 );
and ( n244066 , n244065 , n243698 , n241704 );
and ( n244067 , n32386 , n35431 );
nor ( n244068 , n244066 , n244067 );
nand ( n244069 , n244064 , n244068 );
buf ( n244070 , n244069 );
buf ( n244071 , n38552 );
not ( n244072 , n31957 );
buf ( n244073 , n236798 );
not ( n244074 , n244073 );
or ( n244075 , n244072 , n244074 );
not ( n244076 , n236906 );
not ( n244077 , n239298 );
or ( n244078 , n244076 , n244077 );
not ( n244079 , n236906 );
nand ( n244080 , n244079 , n239297 );
nand ( n244081 , n244078 , n244080 );
and ( n244082 , n244081 , n239399 );
not ( n244083 , n244081 );
and ( n244084 , n244083 , n239391 );
nor ( n244085 , n244082 , n244084 );
not ( n244086 , n27737 );
not ( n244087 , n25501 );
or ( n244088 , n244086 , n244087 );
or ( n244089 , n25501 , n27737 );
nand ( n244090 , n244088 , n244089 );
and ( n244091 , n244090 , n43936 );
not ( n244092 , n244090 );
and ( n244093 , n244092 , n37450 );
nor ( n244094 , n244091 , n244093 );
not ( n244095 , n244094 );
nand ( n244096 , n239561 , n244095 );
not ( n244097 , n244096 );
not ( n244098 , n239536 );
not ( n244099 , n244098 );
and ( n244100 , n244097 , n244099 );
and ( n244101 , n244096 , n244098 );
nor ( n244102 , n244100 , n244101 );
not ( n244103 , n244102 );
not ( n244104 , n239607 );
or ( n244105 , n244103 , n244104 );
not ( n244106 , n244102 );
not ( n244107 , n239488 );
not ( n244108 , n244107 );
and ( n244109 , n239570 , n239600 );
not ( n244110 , n239570 );
and ( n244111 , n244110 , n239597 );
nor ( n244112 , n244109 , n244111 );
not ( n244113 , n244112 );
and ( n244114 , n244108 , n244113 );
and ( n244115 , n244107 , n244112 );
nor ( n244116 , n244114 , n244115 );
nand ( n244117 , n244106 , n244116 );
nand ( n244118 , n244105 , n244117 );
not ( n244119 , n239652 );
not ( n244120 , n244119 );
not ( n244121 , n239635 );
not ( n244122 , n244121 );
or ( n244123 , n244120 , n244122 );
nand ( n244124 , n239635 , n239652 );
nand ( n244125 , n244123 , n244124 );
not ( n244126 , n244125 );
not ( n244127 , n244126 );
and ( n244128 , n244118 , n244127 );
not ( n244129 , n244118 );
and ( n244130 , n244129 , n239654 );
nor ( n244131 , n244128 , n244130 );
nand ( n244132 , n244085 , n244131 );
not ( n244133 , n34125 );
not ( n244134 , n242630 );
not ( n244135 , n33959 );
nand ( n244136 , n33941 , n244135 );
not ( n244137 , n244136 );
and ( n244138 , n244134 , n244137 );
and ( n244139 , n244136 , n242630 );
nor ( n244140 , n244138 , n244139 );
not ( n244141 , n244140 );
not ( n244142 , n244141 );
not ( n244143 , n234702 );
not ( n244144 , n34006 );
nand ( n244145 , n34119 , n244144 );
not ( n244146 , n244145 );
or ( n244147 , n244143 , n244146 );
or ( n244148 , n244145 , n234702 );
nand ( n244149 , n244147 , n244148 );
not ( n244150 , n244149 );
not ( n244151 , n244150 );
or ( n244152 , n244142 , n244151 );
nand ( n244153 , n244149 , n244140 );
nand ( n244154 , n244152 , n244153 );
nand ( n244155 , n235029 , n34311 );
not ( n244156 , n242625 );
and ( n244157 , n244155 , n244156 );
not ( n244158 , n244155 );
and ( n244159 , n244158 , n242625 );
nor ( n244160 , n244157 , n244159 );
not ( n244161 , n244160 );
and ( n244162 , n244154 , n244161 );
not ( n244163 , n244154 );
and ( n244164 , n244163 , n244160 );
nor ( n244165 , n244162 , n244164 );
not ( n244166 , n242648 );
not ( n244167 , n34393 );
nand ( n244168 , n244167 , n34333 );
not ( n244169 , n244168 );
or ( n244170 , n244166 , n244169 );
or ( n244171 , n244168 , n242648 );
nand ( n244172 , n244170 , n244171 );
not ( n244173 , n244172 );
not ( n244174 , n244173 );
nand ( n244175 , n34425 , n33864 );
not ( n244176 , n244175 );
not ( n244177 , n242611 );
and ( n244178 , n244176 , n244177 );
and ( n244179 , n244175 , n242611 );
nor ( n244180 , n244178 , n244179 );
not ( n244181 , n244180 );
not ( n244182 , n244181 );
or ( n244183 , n244174 , n244182 );
nand ( n244184 , n244180 , n244172 );
nand ( n244185 , n244183 , n244184 );
and ( n244186 , n244165 , n244185 );
not ( n244187 , n244165 );
not ( n244188 , n244185 );
and ( n244189 , n244187 , n244188 );
nor ( n244190 , n244186 , n244189 );
not ( n244191 , n244190 );
or ( n244192 , n244133 , n244191 );
not ( n244193 , n34125 );
not ( n244194 , n244185 );
not ( n244195 , n244165 );
or ( n244196 , n244194 , n244195 );
not ( n244197 , n244165 );
nand ( n244198 , n244197 , n244188 );
nand ( n244199 , n244196 , n244198 );
nand ( n244200 , n244193 , n244199 );
nand ( n244201 , n244192 , n244200 );
xor ( n244202 , n233874 , n233868 );
xor ( n244203 , n244202 , n233898 );
buf ( n244204 , n244203 );
and ( n244205 , n244201 , n244204 );
not ( n244206 , n244201 );
not ( n244207 , n244203 );
buf ( n244208 , n244207 );
and ( n244209 , n244206 , n244208 );
nor ( n244210 , n244205 , n244209 );
not ( n244211 , n244210 );
and ( n244212 , n244132 , n244211 );
not ( n244213 , n244132 );
and ( n244214 , n244213 , n244210 );
nor ( n244215 , n244212 , n244214 );
not ( n244216 , n241373 );
buf ( n244217 , n244216 );
or ( n244218 , n244215 , n244217 );
nand ( n244219 , n244075 , n244218 );
buf ( n244220 , n244219 );
not ( n244221 , n233894 );
nand ( n244222 , n33689 , n28726 );
and ( n244223 , n244222 , n28682 );
not ( n244224 , n244222 );
not ( n244225 , n28682 );
and ( n244226 , n244224 , n244225 );
nor ( n244227 , n244223 , n244226 );
not ( n244228 , n244227 );
not ( n244229 , n244228 );
not ( n244230 , n238202 );
nand ( n244231 , n206185 , n33479 );
not ( n244232 , n244231 );
or ( n244233 , n244230 , n244232 );
or ( n244234 , n244231 , n238202 );
nand ( n244235 , n244233 , n244234 );
not ( n244236 , n244235 );
not ( n244237 , n244236 );
or ( n244238 , n244229 , n244237 );
nand ( n244239 , n244235 , n244227 );
nand ( n244240 , n244238 , n244239 );
not ( n244241 , n33621 );
nand ( n244242 , n244241 , n28880 );
not ( n244243 , n244242 );
not ( n244244 , n206593 );
and ( n244245 , n244243 , n244244 );
and ( n244246 , n244242 , n206593 );
nor ( n244247 , n244245 , n244246 );
and ( n244248 , n244240 , n244247 );
not ( n244249 , n244240 );
not ( n244250 , n244247 );
and ( n244251 , n244249 , n244250 );
nor ( n244252 , n244248 , n244251 );
not ( n244253 , n244252 );
not ( n244254 , n28129 );
not ( n244255 , n244254 );
not ( n244256 , n233859 );
nand ( n244257 , n33306 , n244256 );
not ( n244258 , n244257 );
not ( n244259 , n28196 );
not ( n244260 , n244259 );
and ( n244261 , n244258 , n244260 );
and ( n244262 , n244257 , n244259 );
nor ( n244263 , n244261 , n244262 );
not ( n244264 , n244263 );
not ( n244265 , n244264 );
or ( n244266 , n244255 , n244265 );
nand ( n244267 , n244263 , n28129 );
nand ( n244268 , n244266 , n244267 );
not ( n244269 , n244268 );
and ( n244270 , n244253 , n244269 );
not ( n244271 , n244253 );
and ( n244272 , n244271 , n244268 );
nor ( n244273 , n244270 , n244272 );
not ( n244274 , n244273 );
or ( n244275 , n244221 , n244274 );
not ( n244276 , n233894 );
not ( n244277 , n244269 );
not ( n244278 , n244252 );
not ( n244279 , n244278 );
or ( n244280 , n244277 , n244279 );
nand ( n244281 , n244252 , n244268 );
nand ( n244282 , n244280 , n244281 );
nand ( n244283 , n244276 , n244282 );
nand ( n244284 , n244275 , n244283 );
not ( n244285 , n29569 );
nand ( n244286 , n233160 , n29652 );
not ( n244287 , n244286 );
or ( n244288 , n244285 , n244287 );
or ( n244289 , n244286 , n29569 );
nand ( n244290 , n244288 , n244289 );
not ( n244291 , n244290 );
nand ( n244292 , n233120 , n29862 );
not ( n244293 , n244292 );
not ( n244294 , n29779 );
and ( n244295 , n244293 , n244294 );
not ( n244296 , n29863 );
nand ( n244297 , n244296 , n233120 );
and ( n244298 , n244297 , n29779 );
nor ( n244299 , n244295 , n244298 );
not ( n244300 , n244299 );
or ( n244301 , n244291 , n244300 );
or ( n244302 , n244299 , n244290 );
nand ( n244303 , n244301 , n244302 );
not ( n244304 , n244303 );
nor ( n244305 , n233186 , n29260 );
and ( n244306 , n244305 , n29178 );
not ( n244307 , n244305 );
and ( n244308 , n244307 , n29177 );
nor ( n244309 , n244306 , n244308 );
not ( n244310 , n244309 );
nand ( n244311 , n206779 , n55461 );
and ( n244312 , n244311 , n29093 );
not ( n244313 , n244311 );
and ( n244314 , n244313 , n29092 );
nor ( n244315 , n244312 , n244314 );
not ( n244316 , n244315 );
or ( n244317 , n244310 , n244316 );
or ( n244318 , n244315 , n244309 );
nand ( n244319 , n244317 , n244318 );
nand ( n244320 , n29373 , n55487 );
not ( n244321 , n244320 );
not ( n244322 , n29462 );
not ( n244323 , n244322 );
and ( n244324 , n244321 , n244323 );
and ( n244325 , n244320 , n244322 );
nor ( n244326 , n244324 , n244325 );
and ( n244327 , n244319 , n244326 );
not ( n244328 , n244319 );
not ( n244329 , n244326 );
and ( n244330 , n244328 , n244329 );
nor ( n244331 , n244327 , n244330 );
buf ( n244332 , n244331 );
not ( n244333 , n244332 );
and ( n244334 , n244304 , n244333 );
and ( n244335 , n244303 , n244332 );
nor ( n244336 , n244334 , n244335 );
buf ( n244337 , n244336 );
and ( n244338 , n244284 , n244337 );
not ( n244339 , n244284 );
not ( n244340 , n244331 );
not ( n244341 , n244340 );
not ( n244342 , n244303 );
not ( n244343 , n244342 );
or ( n244344 , n244341 , n244343 );
nand ( n244345 , n244331 , n244303 );
nand ( n244346 , n244344 , n244345 );
buf ( n244347 , n244346 );
and ( n244348 , n244339 , n244347 );
nor ( n244349 , n244338 , n244348 );
not ( n244350 , n224643 );
not ( n244351 , n37908 );
not ( n244352 , n29213 );
or ( n244353 , n244351 , n244352 );
or ( n244354 , n206976 , n37908 );
nand ( n244355 , n244353 , n244354 );
not ( n244356 , n244355 );
or ( n244357 , n244350 , n244356 );
or ( n244358 , n244355 , n224643 );
nand ( n244359 , n244357 , n244358 );
nand ( n244360 , n240928 , n244359 );
not ( n244361 , n244360 );
not ( n244362 , n37311 );
and ( n244363 , n244361 , n244362 );
and ( n244364 , n244360 , n37311 );
nor ( n244365 , n244363 , n244364 );
not ( n244366 , n244365 );
not ( n244367 , n244366 );
not ( n244368 , n240941 );
or ( n244369 , n244367 , n244368 );
not ( n244370 , n244366 );
nand ( n244371 , n244370 , n240948 );
nand ( n244372 , n244369 , n244371 );
not ( n244373 , n240996 );
not ( n244374 , n244373 );
and ( n244375 , n244372 , n244374 );
not ( n244376 , n244372 );
and ( n244377 , n244376 , n240997 );
nor ( n244378 , n244375 , n244377 );
nand ( n244379 , n244349 , n244378 );
not ( n244380 , n234385 );
not ( n244381 , n238106 );
or ( n244382 , n244380 , n244381 );
not ( n244383 , n234385 );
nand ( n244384 , n244383 , n238101 );
nand ( n244385 , n244382 , n244384 );
not ( n244386 , n240147 );
buf ( n244387 , n244386 );
and ( n244388 , n244385 , n244387 );
not ( n244389 , n244385 );
buf ( n244390 , n240147 );
and ( n244391 , n244389 , n244390 );
nor ( n244392 , n244388 , n244391 );
not ( n244393 , n234440 );
nand ( n244394 , n244392 , n244393 );
or ( n244395 , n244379 , n244394 );
not ( n244396 , n244392 );
not ( n244397 , n244349 );
or ( n244398 , n244396 , n244397 );
buf ( n244399 , n35427 );
nor ( n244400 , n244378 , n244399 );
nand ( n244401 , n244398 , n244400 );
nand ( n244402 , n50615 , n39990 );
nand ( n244403 , n244395 , n244401 , n244402 );
buf ( n244404 , n244403 );
not ( n244405 , n43056 );
not ( n244406 , n43024 );
nand ( n244407 , n244406 , n236662 );
not ( n244408 , n244407 );
not ( n244409 , n243724 );
and ( n244410 , n244408 , n244409 );
and ( n244411 , n244407 , n243724 );
nor ( n244412 , n244410 , n244411 );
not ( n244413 , n244412 );
not ( n244414 , n43098 );
nand ( n244415 , n236669 , n244414 );
not ( n244416 , n243743 );
and ( n244417 , n244415 , n244416 );
not ( n244418 , n244415 );
and ( n244419 , n244418 , n243743 );
nor ( n244420 , n244417 , n244419 );
not ( n244421 , n244420 );
or ( n244422 , n244413 , n244421 );
or ( n244423 , n244420 , n244412 );
nand ( n244424 , n244422 , n244423 );
not ( n244425 , n243764 );
nand ( n244426 , n236705 , n43140 );
not ( n244427 , n244426 );
and ( n244428 , n244425 , n244427 );
and ( n244429 , n243764 , n244426 );
nor ( n244430 , n244428 , n244429 );
and ( n244431 , n244424 , n244430 );
not ( n244432 , n244424 );
not ( n244433 , n244430 );
and ( n244434 , n244432 , n244433 );
nor ( n244435 , n244431 , n244434 );
nand ( n244436 , n43159 , n43176 );
and ( n244437 , n244436 , n243787 );
not ( n244438 , n244436 );
and ( n244439 , n244438 , n243786 );
nor ( n244440 , n244437 , n244439 );
not ( n244441 , n244440 );
nand ( n244442 , n43206 , n236750 );
xor ( n244443 , n244442 , n243708 );
not ( n244444 , n244443 );
or ( n244445 , n244441 , n244444 );
or ( n244446 , n244443 , n244440 );
nand ( n244447 , n244445 , n244446 );
and ( n244448 , n244435 , n244447 );
not ( n244449 , n244435 );
not ( n244450 , n244447 );
and ( n244451 , n244449 , n244450 );
nor ( n244452 , n244448 , n244451 );
buf ( n244453 , n244452 );
not ( n244454 , n244453 );
or ( n244455 , n244405 , n244454 );
or ( n244456 , n244453 , n43056 );
nand ( n244457 , n244455 , n244456 );
not ( n244458 , n244457 );
not ( n244459 , n244008 );
not ( n244460 , n244459 );
not ( n244461 , n244460 );
and ( n244462 , n244458 , n244461 );
and ( n244463 , n244457 , n244460 );
nor ( n244464 , n244462 , n244463 );
nor ( n244465 , n244464 , n43968 );
not ( n244466 , n233941 );
not ( n244467 , n244336 );
or ( n244468 , n244466 , n244467 );
not ( n244469 , n233941 );
nand ( n244470 , n244469 , n244346 );
nand ( n244471 , n244468 , n244470 );
buf ( n244472 , n241131 );
and ( n244473 , n244471 , n244472 );
not ( n244474 , n244471 );
buf ( n244475 , n241122 );
and ( n244476 , n244474 , n244475 );
nor ( n244477 , n244473 , n244476 );
nor ( n244478 , n244477 , n49955 );
nand ( n244479 , n244465 , n244478 );
not ( n244480 , n244464 );
nor ( n244481 , n244480 , n226955 );
nand ( n244482 , n244481 , n49955 );
nand ( n244483 , n226956 , n244477 );
buf ( n244484 , n35431 );
nand ( n244485 , n244484 , n29690 );
nand ( n244486 , n244479 , n244482 , n244483 , n244485 );
buf ( n244487 , n244486 );
not ( n244488 , RI19aab938_2485);
or ( n244489 , n25328 , n244488 );
not ( n244490 , RI19aa17f8_2556);
or ( n244491 , n25335 , n244490 );
nand ( n244492 , n244489 , n244491 );
buf ( n244493 , n244492 );
nand ( n244494 , n45946 , n46643 );
not ( n244495 , n244494 );
not ( n244496 , n223692 );
not ( n244497 , n244496 );
and ( n244498 , n244495 , n244497 );
and ( n244499 , n244494 , n244496 );
nor ( n244500 , n244498 , n244499 );
not ( n244501 , n244500 );
not ( n244502 , n244501 );
not ( n244503 , n223827 );
or ( n244504 , n244502 , n244503 );
not ( n244505 , n244501 );
nand ( n244506 , n244505 , n46074 );
nand ( n244507 , n244504 , n244506 );
buf ( n244508 , n238792 );
not ( n244509 , n244508 );
and ( n244510 , n244507 , n244509 );
not ( n244511 , n244507 );
and ( n244512 , n244511 , n244508 );
nor ( n244513 , n244510 , n244512 );
not ( n244514 , n244513 );
not ( n244515 , n234021 );
nand ( n244516 , n244514 , n244515 );
not ( n244517 , n47075 );
nand ( n244518 , n224865 , n244517 );
and ( n244519 , n244518 , n228578 );
not ( n244520 , n244518 );
and ( n244521 , n244520 , n228577 );
nor ( n244522 , n244519 , n244521 );
not ( n244523 , n244522 );
not ( n244524 , n50940 );
or ( n244525 , n244523 , n244524 );
not ( n244526 , n244522 );
nand ( n244527 , n244526 , n50930 );
nand ( n244528 , n244525 , n244527 );
buf ( n244529 , n225301 );
and ( n244530 , n244528 , n244529 );
not ( n244531 , n244528 );
buf ( n244532 , n47531 );
and ( n244533 , n244531 , n244532 );
nor ( n244534 , n244530 , n244533 );
not ( n244535 , n244534 );
not ( n244536 , n236288 );
not ( n244537 , n239665 );
nand ( n244538 , n51815 , n236329 );
not ( n244539 , n244538 );
not ( n244540 , n238963 );
or ( n244541 , n244539 , n244540 );
or ( n244542 , n238963 , n244538 );
nand ( n244543 , n244541 , n244542 );
not ( n244544 , n244543 );
not ( n244545 , n244544 );
or ( n244546 , n244537 , n244545 );
nand ( n244547 , n244543 , n239664 );
nand ( n244548 , n244546 , n244547 );
nand ( n244549 , n236371 , n51898 );
and ( n244550 , n244549 , n239668 );
not ( n244551 , n244549 );
and ( n244552 , n244551 , n229532 );
nor ( n244553 , n244550 , n244552 );
xor ( n244554 , n244548 , n244553 );
not ( n244555 , n238920 );
nand ( n244556 , n236307 , n51984 );
not ( n244557 , n244556 );
or ( n244558 , n244555 , n244557 );
or ( n244559 , n244556 , n238920 );
nand ( n244560 , n244558 , n244559 );
not ( n244561 , n236281 );
nand ( n244562 , n244561 , n229678 );
and ( n244563 , n244562 , n238939 );
not ( n244564 , n244562 );
and ( n244565 , n244564 , n239674 );
nor ( n244566 , n244563 , n244565 );
or ( n244567 , n244560 , n244566 );
nand ( n244568 , n244566 , n244560 );
nand ( n244569 , n244567 , n244568 );
not ( n244570 , n244569 );
and ( n244571 , n244554 , n244570 );
not ( n244572 , n244554 );
and ( n244573 , n244572 , n244569 );
nor ( n244574 , n244571 , n244573 );
not ( n244575 , n244574 );
or ( n244576 , n244536 , n244575 );
not ( n244577 , n236288 );
not ( n244578 , n244554 );
not ( n244579 , n244570 );
and ( n244580 , n244578 , n244579 );
and ( n244581 , n244554 , n244570 );
nor ( n244582 , n244580 , n244581 );
not ( n244583 , n244582 );
nand ( n244584 , n244577 , n244583 );
nand ( n244585 , n244576 , n244584 );
not ( n244586 , n241255 );
not ( n244587 , n244586 );
and ( n244588 , n244585 , n244587 );
not ( n244589 , n244585 );
buf ( n244590 , n241255 );
not ( n244591 , n244590 );
and ( n244592 , n244589 , n244591 );
nor ( n244593 , n244588 , n244592 );
not ( n244594 , n244593 );
nand ( n244595 , n244535 , n244594 );
or ( n244596 , n244516 , n244595 );
not ( n244597 , n244535 );
not ( n244598 , n244514 );
or ( n244599 , n244597 , n244598 );
nor ( n244600 , n244594 , n33254 );
nand ( n244601 , n244599 , n244600 );
nand ( n244602 , n239240 , n45190 );
nand ( n244603 , n244596 , n244601 , n244602 );
buf ( n244604 , n244603 );
not ( n244605 , n207153 );
not ( n244606 , n25335 );
not ( n244607 , n244606 );
or ( n244608 , n244605 , n244607 );
not ( n244609 , n51375 );
nand ( n244610 , n244609 , n51363 );
and ( n244611 , n51368 , n244610 );
not ( n244612 , RI1754c430_6);
or ( n244613 , n244611 , n244612 );
nand ( n244614 , n244608 , n244613 );
buf ( n244615 , n244614 );
not ( n244616 , RI19aa1438_2558);
or ( n244617 , n25328 , n244616 );
or ( n244618 , n25335 , n41949 );
nand ( n244619 , n244617 , n244618 );
buf ( n244620 , n244619 );
not ( n244621 , n222419 );
not ( n244622 , n237810 );
or ( n244623 , n244621 , n244622 );
or ( n244624 , n237810 , n222419 );
nand ( n244625 , n244623 , n244624 );
and ( n244626 , n244625 , n237868 );
not ( n244627 , n244625 );
and ( n244628 , n244627 , n237869 );
nor ( n244629 , n244626 , n244628 );
nand ( n244630 , n244629 , n244515 );
not ( n244631 , n225052 );
not ( n244632 , n47294 );
nand ( n244633 , n244632 , n40683 );
not ( n244634 , n244633 );
or ( n244635 , n244631 , n244634 );
not ( n244636 , n40683 );
not ( n244637 , n244636 );
nand ( n244638 , n244637 , n244632 );
or ( n244639 , n244638 , n225052 );
nand ( n244640 , n244635 , n244639 );
not ( n244641 , n244640 );
not ( n244642 , n47310 );
or ( n244643 , n244641 , n244642 );
not ( n244644 , n244640 );
nand ( n244645 , n244644 , n47319 );
nand ( n244646 , n244643 , n244645 );
and ( n244647 , n244646 , n225086 );
not ( n244648 , n244646 );
and ( n244649 , n244648 , n225083 );
nor ( n244650 , n244647 , n244649 );
not ( n244651 , n53373 );
not ( n244652 , n244651 );
nand ( n244653 , n237010 , n237044 );
not ( n244654 , n244653 );
or ( n244655 , n244652 , n244654 );
or ( n244656 , n244653 , n244651 );
nand ( n244657 , n244655 , n244656 );
not ( n244658 , n244657 );
nand ( n244659 , n237045 , n53373 );
and ( n244660 , n244659 , n237014 );
not ( n244661 , n244659 );
and ( n244662 , n244661 , n53385 );
nor ( n244663 , n244660 , n244662 );
not ( n244664 , n244663 );
not ( n244665 , n231120 );
nand ( n244666 , n244665 , n237070 );
and ( n244667 , n244666 , n53349 );
not ( n244668 , n244666 );
not ( n244669 , n53349 );
and ( n244670 , n244668 , n244669 );
nor ( n244671 , n244667 , n244670 );
not ( n244672 , n244671 );
or ( n244673 , n244664 , n244672 );
or ( n244674 , n244671 , n244663 );
nand ( n244675 , n244673 , n244674 );
and ( n244676 , n244675 , n241713 );
not ( n244677 , n244675 );
and ( n244678 , n244677 , n241712 );
nor ( n244679 , n244676 , n244678 );
nand ( n244680 , n53282 , n237102 );
not ( n244681 , n231053 );
and ( n244682 , n244680 , n244681 );
not ( n244683 , n244680 );
and ( n244684 , n244683 , n231053 );
nor ( n244685 , n244682 , n244684 );
not ( n244686 , n244685 );
not ( n244687 , n244686 );
not ( n244688 , n231061 );
nand ( n244689 , n244688 , n237126 );
and ( n244690 , n244689 , n53313 );
not ( n244691 , n244689 );
not ( n244692 , n53313 );
and ( n244693 , n244691 , n244692 );
nor ( n244694 , n244690 , n244693 );
not ( n244695 , n244694 );
not ( n244696 , n244695 );
or ( n244697 , n244687 , n244696 );
nand ( n244698 , n244694 , n244685 );
nand ( n244699 , n244697 , n244698 );
not ( n244700 , n244699 );
and ( n244701 , n244679 , n244700 );
not ( n244702 , n244679 );
and ( n244703 , n244702 , n244699 );
nor ( n244704 , n244701 , n244703 );
not ( n244705 , n244704 );
or ( n244706 , n244658 , n244705 );
not ( n244707 , n244657 );
and ( n244708 , n244679 , n244699 );
not ( n244709 , n244679 );
and ( n244710 , n244709 , n244700 );
nor ( n244711 , n244708 , n244710 );
nand ( n244712 , n244707 , n244711 );
nand ( n244713 , n244706 , n244712 );
nand ( n244714 , n237212 , n241860 );
not ( n244715 , n244714 );
not ( n244716 , n241850 );
and ( n244717 , n244715 , n244716 );
and ( n244718 , n244714 , n241850 );
nor ( n244719 , n244717 , n244718 );
not ( n244720 , n244719 );
not ( n244721 , n244720 );
nand ( n244722 , n241820 , n237252 );
and ( n244723 , n244722 , n241832 );
not ( n244724 , n244722 );
and ( n244725 , n244724 , n241831 );
nor ( n244726 , n244723 , n244725 );
not ( n244727 , n244726 );
not ( n244728 , n244727 );
or ( n244729 , n244721 , n244728 );
nand ( n244730 , n244726 , n244719 );
nand ( n244731 , n244729 , n244730 );
not ( n244732 , n244731 );
not ( n244733 , n244732 );
nand ( n244734 , n241736 , n237325 );
not ( n244735 , n244734 );
not ( n244736 , n241747 );
not ( n244737 , n244736 );
and ( n244738 , n244735 , n244737 );
and ( n244739 , n244734 , n244736 );
nor ( n244740 , n244738 , n244739 );
not ( n244741 , n244740 );
not ( n244742 , n241772 );
nand ( n244743 , n237263 , n244742 );
and ( n244744 , n244743 , n241762 );
not ( n244745 , n244743 );
not ( n244746 , n241762 );
and ( n244747 , n244745 , n244746 );
nor ( n244748 , n244744 , n244747 );
not ( n244749 , n244748 );
or ( n244750 , n244741 , n244749 );
or ( n244751 , n244748 , n244740 );
nand ( n244752 , n244750 , n244751 );
not ( n244753 , n241789 );
nand ( n244754 , n244753 , n237183 );
and ( n244755 , n244754 , n241800 );
not ( n244756 , n244754 );
and ( n244757 , n244756 , n241799 );
nor ( n244758 , n244755 , n244757 );
and ( n244759 , n244752 , n244758 );
not ( n244760 , n244752 );
not ( n244761 , n244758 );
and ( n244762 , n244760 , n244761 );
nor ( n244763 , n244759 , n244762 );
not ( n244764 , n244763 );
or ( n244765 , n244733 , n244764 );
not ( n244766 , n244763 );
nand ( n244767 , n244766 , n244731 );
nand ( n244768 , n244765 , n244767 );
buf ( n244769 , n244768 );
and ( n244770 , n244713 , n244769 );
not ( n244771 , n244713 );
and ( n244772 , n244766 , n244731 );
not ( n244773 , n244766 );
not ( n244774 , n244731 );
and ( n244775 , n244773 , n244774 );
nor ( n244776 , n244772 , n244775 );
not ( n244777 , n244776 );
not ( n244778 , n244777 );
and ( n244779 , n244771 , n244778 );
nor ( n244780 , n244770 , n244779 );
not ( n244781 , n244780 );
nand ( n244782 , n244650 , n244781 );
or ( n244783 , n244630 , n244782 );
not ( n244784 , n244629 );
not ( n244785 , n244650 );
or ( n244786 , n244784 , n244785 );
nor ( n244787 , n244781 , n241065 );
nand ( n244788 , n244786 , n244787 );
buf ( n244789 , n35431 );
nand ( n244790 , n244789 , n39387 );
nand ( n244791 , n244783 , n244788 , n244790 );
buf ( n244792 , n244791 );
buf ( n244793 , n30275 );
buf ( n244794 , n25662 );
buf ( n244795 , n30075 );
buf ( n244796 , n41145 );
not ( n244797 , n240915 );
not ( n244798 , n37708 );
or ( n244799 , n244797 , n244798 );
or ( n244800 , n37708 , n240915 );
nand ( n244801 , n244799 , n244800 );
buf ( n244802 , n54134 );
and ( n244803 , n244801 , n244802 );
not ( n244804 , n244801 );
not ( n244805 , n244802 );
and ( n244806 , n244804 , n244805 );
nor ( n244807 , n244803 , n244806 );
not ( n244808 , n244807 );
not ( n244809 , n243434 );
nand ( n244810 , n244808 , n244809 );
not ( n244811 , n237680 );
not ( n244812 , n244811 );
not ( n244813 , n44176 );
or ( n244814 , n244812 , n244813 );
or ( n244815 , n44176 , n244811 );
nand ( n244816 , n244814 , n244815 );
and ( n244817 , n244816 , n44325 );
not ( n244818 , n244816 );
and ( n244819 , n244818 , n44316 );
nor ( n244820 , n244817 , n244819 );
not ( n244821 , n242509 );
not ( n244822 , n241657 );
or ( n244823 , n244821 , n244822 );
nand ( n244824 , n241656 , n242510 );
nand ( n244825 , n244823 , n244824 );
buf ( n244826 , n227548 );
and ( n244827 , n244825 , n244826 );
not ( n244828 , n244825 );
and ( n244829 , n244828 , n241662 );
nor ( n244830 , n244827 , n244829 );
nand ( n244831 , n244820 , n244830 );
or ( n244832 , n244810 , n244831 );
not ( n244833 , n244820 );
not ( n244834 , n244807 );
not ( n244835 , n244834 );
or ( n244836 , n244833 , n244835 );
not ( n244837 , n222532 );
nor ( n244838 , n244830 , n244837 );
nand ( n244839 , n244836 , n244838 );
buf ( n244840 , n35431 );
nand ( n244841 , n244840 , n37371 );
nand ( n244842 , n244832 , n244839 , n244841 );
buf ( n244843 , n244842 );
nand ( n244844 , n234619 , n234622 );
and ( n244845 , n244844 , n53459 );
not ( n244846 , n244844 );
and ( n244847 , n244846 , n53458 );
nor ( n244848 , n244845 , n244847 );
not ( n244849 , n244848 );
not ( n244850 , n236815 );
not ( n244851 , n53516 );
nand ( n244852 , n244851 , n234570 );
and ( n244853 , n244852 , n53528 );
not ( n244854 , n244852 );
not ( n244855 , n53528 );
and ( n244856 , n244854 , n244855 );
nor ( n244857 , n244853 , n244856 );
not ( n244858 , n244857 );
or ( n244859 , n244850 , n244858 );
or ( n244860 , n244857 , n236815 );
nand ( n244861 , n244859 , n244860 );
and ( n244862 , n244861 , n231422 );
not ( n244863 , n244861 );
and ( n244864 , n244863 , n53486 );
nor ( n244865 , n244862 , n244864 );
not ( n244866 , n244865 );
not ( n244867 , n234667 );
not ( n244868 , n53647 );
nand ( n244869 , n244867 , n244868 );
not ( n244870 , n244869 );
not ( n244871 , n231391 );
buf ( n244872 , n244871 );
not ( n244873 , n244872 );
and ( n244874 , n244870 , n244873 );
and ( n244875 , n244869 , n244872 );
nor ( n244876 , n244874 , n244875 );
not ( n244877 , n53594 );
nand ( n244878 , n244877 , n234639 );
and ( n244879 , n244878 , n53584 );
not ( n244880 , n244878 );
and ( n244881 , n244880 , n234544 );
nor ( n244882 , n244879 , n244881 );
or ( n244883 , n244876 , n244882 );
nand ( n244884 , n244882 , n244876 );
nand ( n244885 , n244883 , n244884 );
not ( n244886 , n244885 );
and ( n244887 , n244866 , n244886 );
and ( n244888 , n244865 , n244885 );
nor ( n244889 , n244887 , n244888 );
not ( n244890 , n244889 );
or ( n244891 , n244849 , n244890 );
not ( n244892 , n244848 );
not ( n244893 , n244885 );
not ( n244894 , n244893 );
not ( n244895 , n244865 );
not ( n244896 , n244895 );
or ( n244897 , n244894 , n244896 );
nand ( n244898 , n244865 , n244885 );
nand ( n244899 , n244897 , n244898 );
nand ( n244900 , n244892 , n244899 );
nand ( n244901 , n244891 , n244900 );
not ( n244902 , n34106 );
nand ( n244903 , n244902 , n234708 );
not ( n244904 , n244903 );
not ( n244905 , n244144 );
and ( n244906 , n244904 , n244905 );
not ( n244907 , n34106 );
nand ( n244908 , n244907 , n234708 );
and ( n244909 , n244908 , n244144 );
nor ( n244910 , n244906 , n244909 );
nand ( n244911 , n242632 , n234776 );
not ( n244912 , n244911 );
buf ( n244913 , n33941 );
not ( n244914 , n244913 );
and ( n244915 , n244912 , n244914 );
and ( n244916 , n244911 , n244913 );
nor ( n244917 , n244915 , n244916 );
not ( n244918 , n244917 );
not ( n244919 , n244918 );
not ( n244920 , n235033 );
not ( n244921 , n244920 );
or ( n244922 , n244919 , n244921 );
nand ( n244923 , n235033 , n244917 );
nand ( n244924 , n244922 , n244923 );
xor ( n244925 , n244910 , n244924 );
nand ( n244926 , n34348 , n234727 );
not ( n244927 , n244926 );
not ( n244928 , n34333 );
and ( n244929 , n244927 , n244928 );
and ( n244930 , n244926 , n34333 );
nor ( n244931 , n244929 , n244930 );
not ( n244932 , n244931 );
not ( n244933 , n244932 );
not ( n244934 , n33866 );
not ( n244935 , n244934 );
or ( n244936 , n244933 , n244935 );
nand ( n244937 , n33866 , n244931 );
nand ( n244938 , n244936 , n244937 );
xor ( n244939 , n244925 , n244938 );
buf ( n244940 , n244939 );
and ( n244941 , n244901 , n244940 );
not ( n244942 , n244901 );
not ( n244943 , n244924 );
not ( n244944 , n244943 );
not ( n244945 , n244910 );
not ( n244946 , n244938 );
or ( n244947 , n244945 , n244946 );
or ( n244948 , n244938 , n244910 );
nand ( n244949 , n244947 , n244948 );
not ( n244950 , n244949 );
or ( n244951 , n244944 , n244950 );
not ( n244952 , n244949 );
nand ( n244953 , n244952 , n244924 );
nand ( n244954 , n244951 , n244953 );
buf ( n244955 , n244954 );
and ( n244956 , n244942 , n244955 );
nor ( n244957 , n244941 , n244956 );
nor ( n244958 , n244957 , n43968 );
not ( n244959 , n53454 );
not ( n244960 , n33053 );
not ( n244961 , n244960 );
not ( n244962 , n53248 );
or ( n244963 , n244961 , n244962 );
nand ( n244964 , n53257 , n33053 );
nand ( n244965 , n244963 , n244964 );
not ( n244966 , n244965 );
or ( n244967 , n244959 , n244966 );
or ( n244968 , n244965 , n53694 );
nand ( n244969 , n244967 , n244968 );
not ( n244970 , n51530 );
not ( n244971 , n239653 );
or ( n244972 , n244970 , n244971 );
not ( n244973 , n51530 );
nand ( n244974 , n244973 , n244125 );
nand ( n244975 , n244972 , n244974 );
and ( n244976 , n244975 , n241695 );
not ( n244977 , n244975 );
not ( n244978 , n45873 );
and ( n244979 , n244977 , n244978 );
nor ( n244980 , n244976 , n244979 );
nor ( n244981 , n244969 , n244980 );
nand ( n244982 , n244958 , n244981 );
not ( n244983 , n244957 );
not ( n244984 , n244980 );
nand ( n244985 , n244983 , n244984 );
nand ( n244986 , n244985 , n244969 , n241373 );
buf ( n244987 , n31577 );
nand ( n244988 , n244987 , n29020 );
nand ( n244989 , n244982 , n244986 , n244988 );
buf ( n244990 , n244989 );
buf ( n244991 , RI175373a0_595);
and ( n244992 , n27883 , n244991 );
buf ( n244993 , n244992 );
not ( n244994 , RI19abf0f0_2340);
or ( n244995 , n25328 , n244994 );
not ( n244996 , RI19ab5d48_2410);
or ( n244997 , n25335 , n244996 );
nand ( n244998 , n244995 , n244997 );
buf ( n244999 , n244998 );
buf ( n245000 , RI17539e48_588);
nor ( n245001 , n204514 , n35631 , n35632 , n245000 );
not ( n245002 , n245001 );
not ( n245003 , RI17536d88_596);
and ( n245004 , n35629 , n245003 , n204525 );
and ( n245005 , n245004 , n204516 );
nand ( n245006 , n245005 , n204524 , n204517 , n35627 );
xor ( n245007 , n245006 , n53874 );
not ( n245008 , n34227 );
buf ( n245009 , n40513 );
not ( n245010 , n245009 );
not ( n245011 , n34191 );
or ( n245012 , n245010 , n245011 );
or ( n245013 , n34191 , n245009 );
nand ( n245014 , n245012 , n245013 );
not ( n245015 , n245014 );
or ( n245016 , n245008 , n245015 );
or ( n245017 , n245014 , n34227 );
nand ( n245018 , n245016 , n245017 );
nor ( n245019 , n245018 , n238331 );
xor ( n245020 , n245007 , n245019 );
not ( n245021 , n245020 );
not ( n245022 , n245021 );
not ( n245023 , n34637 );
not ( n245024 , n37449 );
or ( n245025 , n245023 , n245024 );
or ( n245026 , n37449 , n34637 );
nand ( n245027 , n245025 , n245026 );
and ( n245028 , n245027 , n37458 );
not ( n245029 , n245027 );
and ( n245030 , n245029 , n37455 );
nor ( n245031 , n245028 , n245030 );
not ( n245032 , n245031 );
nand ( n245033 , n245032 , n53841 );
not ( n245034 , n245033 );
not ( n245035 , n231591 );
and ( n245036 , n245034 , n245035 );
not ( n245037 , n245031 );
nand ( n245038 , n245037 , n53841 );
and ( n245039 , n245038 , n231591 );
nor ( n245040 , n245036 , n245039 );
not ( n245041 , n245040 );
nand ( n245042 , n53874 , n245018 );
and ( n245043 , n245042 , n53864 );
not ( n245044 , n245042 );
and ( n245045 , n245044 , n53863 );
nor ( n245046 , n245043 , n245045 );
not ( n245047 , n245046 );
or ( n245048 , n245041 , n245047 );
or ( n245049 , n245046 , n245040 );
nand ( n245050 , n245048 , n245049 );
not ( n245051 , n231670 );
not ( n245052 , n31254 );
not ( n245053 , n27845 );
not ( n245054 , n33759 );
or ( n245055 , n245053 , n245054 );
or ( n245056 , n243295 , n27845 );
nand ( n245057 , n245055 , n245056 );
not ( n245058 , n245057 );
and ( n245059 , n245052 , n245058 );
and ( n245060 , n33768 , n245057 );
nor ( n245061 , n245059 , n245060 );
not ( n245062 , n245061 );
nand ( n245063 , n245051 , n245062 );
and ( n245064 , n245063 , n231658 );
not ( n245065 , n245063 );
and ( n245066 , n245065 , n238338 );
nor ( n245067 , n245064 , n245066 );
not ( n245068 , n245067 );
and ( n245069 , n245050 , n245068 );
not ( n245070 , n245050 );
and ( n245071 , n245070 , n245067 );
nor ( n245072 , n245069 , n245071 );
not ( n245073 , n53977 );
and ( n245074 , n25424 , n41405 );
not ( n245075 , n25424 );
and ( n245076 , n245075 , n30247 );
or ( n245077 , n245074 , n245076 );
and ( n245078 , n245077 , n41412 );
not ( n245079 , n245077 );
and ( n245080 , n245079 , n41416 );
nor ( n245081 , n245078 , n245080 );
nand ( n245082 , n245073 , n245081 );
not ( n245083 , n245082 );
not ( n245084 , n238375 );
and ( n245085 , n245083 , n245084 );
not ( n245086 , n53977 );
nand ( n245087 , n245086 , n245081 );
and ( n245088 , n245087 , n238375 );
nor ( n245089 , n245085 , n245088 );
not ( n245090 , n245089 );
not ( n245091 , n245090 );
xor ( n245092 , n25674 , n52185 );
xnor ( n245093 , n245092 , n40969 );
nand ( n245094 , n245093 , n231703 );
not ( n245095 , n245094 );
not ( n245096 , n231688 );
and ( n245097 , n245095 , n245096 );
nand ( n245098 , n245093 , n231703 );
and ( n245099 , n245098 , n231688 );
nor ( n245100 , n245097 , n245099 );
not ( n245101 , n245100 );
or ( n245102 , n245091 , n245101 );
not ( n245103 , n245100 );
nand ( n245104 , n245103 , n245089 );
nand ( n245105 , n245102 , n245104 );
and ( n245106 , n245072 , n245105 );
not ( n245107 , n245072 );
not ( n245108 , n245105 );
and ( n245109 , n245107 , n245108 );
nor ( n245110 , n245106 , n245109 );
not ( n245111 , n245110 );
or ( n245112 , n245022 , n245111 );
not ( n245113 , n245021 );
not ( n245114 , n245110 );
nand ( n245115 , n245113 , n245114 );
nand ( n245116 , n245112 , n245115 );
not ( n245117 , n40669 );
nand ( n245118 , n225052 , n245117 );
buf ( n245119 , n40659 );
and ( n245120 , n245118 , n245119 );
not ( n245121 , n245118 );
not ( n245122 , n245119 );
and ( n245123 , n245121 , n245122 );
nor ( n245124 , n245120 , n245123 );
not ( n245125 , n245124 );
not ( n245126 , n245125 );
not ( n245127 , n40818 );
nand ( n245128 , n245127 , n47263 );
not ( n245129 , n245128 );
not ( n245130 , n40770 );
not ( n245131 , n245130 );
and ( n245132 , n245129 , n245131 );
and ( n245133 , n245128 , n245130 );
nor ( n245134 , n245132 , n245133 );
not ( n245135 , n245134 );
not ( n245136 , n245135 );
or ( n245137 , n245126 , n245136 );
nand ( n245138 , n245134 , n245124 );
nand ( n245139 , n245137 , n245138 );
not ( n245140 , n245139 );
not ( n245141 , n40579 );
nand ( n245142 , n40625 , n47202 );
not ( n245143 , n245142 );
not ( n245144 , n40611 );
and ( n245145 , n245143 , n245144 );
and ( n245146 , n245142 , n40611 );
nor ( n245147 , n245145 , n245146 );
not ( n245148 , n245147 );
or ( n245149 , n245141 , n245148 );
or ( n245150 , n245147 , n40579 );
nand ( n245151 , n245149 , n245150 );
not ( n245152 , n40736 );
nand ( n245153 , n245152 , n47235 );
buf ( n245154 , n40699 );
not ( n245155 , n245154 );
and ( n245156 , n245153 , n245155 );
not ( n245157 , n245153 );
and ( n245158 , n245157 , n245154 );
nor ( n245159 , n245156 , n245158 );
not ( n245160 , n245159 );
and ( n245161 , n245151 , n245160 );
not ( n245162 , n245151 );
and ( n245163 , n245162 , n245159 );
nor ( n245164 , n245161 , n245163 );
not ( n245165 , n245164 );
not ( n245166 , n245165 );
or ( n245167 , n245140 , n245166 );
not ( n245168 , n245139 );
nand ( n245169 , n245168 , n245164 );
nand ( n245170 , n245167 , n245169 );
buf ( n245171 , n245170 );
and ( n245172 , n245116 , n245171 );
not ( n245173 , n245116 );
not ( n245174 , n245170 );
and ( n245175 , n245173 , n245174 );
nor ( n245176 , n245172 , n245175 );
not ( n245177 , n245176 );
or ( n245178 , n245002 , n245177 );
or ( n245179 , n245176 , n245001 );
nand ( n245180 , n245178 , n245179 );
not ( n245181 , n242079 );
buf ( n245182 , n239733 );
not ( n245183 , n245182 );
not ( n245184 , n239099 );
or ( n245185 , n245183 , n245184 );
or ( n245186 , n239099 , n245182 );
nand ( n245187 , n245185 , n245186 );
not ( n245188 , n245187 );
not ( n245189 , n245188 );
or ( n245190 , n245181 , n245189 );
nand ( n245191 , n242069 , n245187 );
nand ( n245192 , n245190 , n245191 );
not ( n245193 , n245192 );
not ( n245194 , n51946 );
not ( n245195 , n236381 );
not ( n245196 , n245195 );
not ( n245197 , n236313 );
not ( n245198 , n245197 );
or ( n245199 , n245196 , n245198 );
nand ( n245200 , n236381 , n236313 );
nand ( n245201 , n245199 , n245200 );
not ( n245202 , n245201 );
or ( n245203 , n245194 , n245202 );
or ( n245204 , n245201 , n51946 );
nand ( n245205 , n245203 , n245204 );
not ( n245206 , n245205 );
not ( n245207 , n236392 );
or ( n245208 , n245206 , n245207 );
not ( n245209 , n245205 );
xnor ( n245210 , n236204 , n236266 );
buf ( n245211 , n245210 );
nand ( n245212 , n245209 , n245211 );
nand ( n245213 , n245208 , n245212 );
nand ( n245214 , n245193 , n245213 );
and ( n245215 , n245180 , n245214 );
not ( n245216 , n245180 );
not ( n245217 , n245214 );
and ( n245218 , n245216 , n245217 );
nor ( n245219 , n245215 , n245218 );
or ( n245220 , n245219 , n234818 );
buf ( n245221 , n35431 );
nand ( n245222 , n245221 , n41686 );
nand ( n245223 , n245220 , n245222 );
buf ( n245224 , n245223 );
nand ( n245225 , n46884 , n46755 );
and ( n245226 , n245225 , n50750 );
not ( n245227 , n245225 );
and ( n245228 , n245227 , n50749 );
nor ( n245229 , n245226 , n245228 );
not ( n245230 , n245229 );
not ( n245231 , n245230 );
not ( n245232 , n50776 );
or ( n245233 , n245231 , n245232 );
or ( n245234 , n50776 , n245230 );
nand ( n245235 , n245233 , n245234 );
and ( n245236 , n245235 , n50931 );
not ( n245237 , n245235 );
and ( n245238 , n245237 , n50941 );
nor ( n245239 , n245236 , n245238 );
not ( n245240 , n245239 );
buf ( n245241 , n205649 );
nand ( n245242 , n245240 , n245241 );
nand ( n245243 , n40180 , n235767 );
not ( n245244 , n245243 );
not ( n245245 , n240023 );
and ( n245246 , n245244 , n245245 );
and ( n245247 , n245243 , n240023 );
nor ( n245248 , n245246 , n245247 );
buf ( n245249 , n245248 );
not ( n245250 , n245249 );
not ( n245251 , n245250 );
not ( n245252 , n230367 );
or ( n245253 , n245251 , n245252 );
not ( n245254 , n245250 );
nand ( n245255 , n245254 , n230374 );
nand ( n245256 , n245253 , n245255 );
and ( n245257 , n245256 , n52757 );
not ( n245258 , n245256 );
not ( n245259 , n230512 );
not ( n245260 , n230455 );
not ( n245261 , n245260 );
or ( n245262 , n245259 , n245261 );
nand ( n245263 , n230455 , n52752 );
nand ( n245264 , n245262 , n245263 );
buf ( n245265 , n245264 );
and ( n245266 , n245258 , n245265 );
nor ( n245267 , n245257 , n245266 );
not ( n245268 , n245267 );
not ( n245269 , n242053 );
not ( n245270 , n241330 );
nand ( n245271 , n245270 , n44513 );
not ( n245272 , n245271 );
or ( n245273 , n245269 , n245272 );
not ( n245274 , n44512 );
nand ( n245275 , n245274 , n245270 );
or ( n245276 , n245275 , n242053 );
nand ( n245277 , n245273 , n245276 );
not ( n245278 , n245277 );
nand ( n245279 , n222281 , n241346 );
not ( n245280 , n245279 );
not ( n245281 , n222102 );
and ( n245282 , n245280 , n245281 );
and ( n245283 , n245279 , n222102 );
nor ( n245284 , n245282 , n245283 );
not ( n245285 , n245284 );
or ( n245286 , n245278 , n245285 );
or ( n245287 , n245284 , n245277 );
nand ( n245288 , n245286 , n245287 );
not ( n245289 , n245288 );
not ( n245290 , n241275 );
nand ( n245291 , n245290 , n44473 );
not ( n245292 , n245291 );
not ( n245293 , n241993 );
not ( n245294 , n245293 );
and ( n245295 , n245292 , n245294 );
and ( n245296 , n245291 , n245293 );
nor ( n245297 , n245295 , n245296 );
not ( n245298 , n245297 );
not ( n245299 , n242008 );
not ( n245300 , n245299 );
not ( n245301 , n241295 );
nand ( n245302 , n245301 , n222205 );
not ( n245303 , n245302 );
or ( n245304 , n245300 , n245303 );
or ( n245305 , n245302 , n245299 );
nand ( n245306 , n245304 , n245305 );
not ( n245307 , n245306 );
nand ( n245308 , n44402 , n241314 );
not ( n245309 , n245308 );
not ( n245310 , n49725 );
not ( n245311 , n242018 );
or ( n245312 , n245310 , n245311 );
or ( n245313 , n225090 , n242018 );
nand ( n245314 , n245312 , n245313 );
not ( n245315 , n245314 );
and ( n245316 , n245309 , n245315 );
not ( n245317 , n242024 );
nand ( n245318 , n245317 , n44402 );
and ( n245319 , n245318 , n245314 );
nor ( n245320 , n245316 , n245319 );
not ( n245321 , n245320 );
or ( n245322 , n245307 , n245321 );
or ( n245323 , n245320 , n245306 );
nand ( n245324 , n245322 , n245323 );
not ( n245325 , n245324 );
and ( n245326 , n245298 , n245325 );
and ( n245327 , n245297 , n245324 );
nor ( n245328 , n245326 , n245327 );
not ( n245329 , n245328 );
or ( n245330 , n245289 , n245329 );
or ( n245331 , n245288 , n245328 );
nand ( n245332 , n245330 , n245331 );
not ( n245333 , n245332 );
not ( n245334 , n245333 );
not ( n245335 , n245334 );
not ( n245336 , n241334 );
and ( n245337 , n245335 , n245336 );
buf ( n245338 , n245332 );
and ( n245339 , n245338 , n241334 );
nor ( n245340 , n245337 , n245339 );
nor ( n245341 , n235254 , n44617 );
not ( n245342 , n245341 );
buf ( n245343 , n235264 );
not ( n245344 , n245343 );
and ( n245345 , n245342 , n245344 );
and ( n245346 , n245341 , n245343 );
nor ( n245347 , n245345 , n245346 );
not ( n245348 , n245347 );
not ( n245349 , n245348 );
nor ( n245350 , n44745 , n235293 );
not ( n245351 , n245350 );
not ( n245352 , n245351 );
not ( n245353 , n235282 );
or ( n245354 , n245352 , n245353 );
nand ( n245355 , n235283 , n245350 );
nand ( n245356 , n245354 , n245355 );
not ( n245357 , n245356 );
not ( n245358 , n245357 );
or ( n245359 , n245349 , n245358 );
nand ( n245360 , n245356 , n245347 );
nand ( n245361 , n245359 , n245360 );
not ( n245362 , n245361 );
nand ( n245363 , n235302 , n44673 );
not ( n245364 , n245363 );
not ( n245365 , n235314 );
not ( n245366 , n245365 );
and ( n245367 , n245364 , n245366 );
and ( n245368 , n245363 , n245365 );
nor ( n245369 , n245367 , n245368 );
not ( n245370 , n245369 );
and ( n245371 , n245362 , n245370 );
and ( n245372 , n245361 , n245369 );
nor ( n245373 , n245371 , n245372 );
not ( n245374 , n245373 );
not ( n245375 , n235242 );
not ( n245376 , n235341 );
nand ( n245377 , n245376 , n44556 );
not ( n245378 , n245377 );
not ( n245379 , n235330 );
not ( n245380 , n245379 );
or ( n245381 , n245378 , n245380 );
or ( n245382 , n245379 , n245377 );
nand ( n245383 , n245381 , n245382 );
not ( n245384 , n245383 );
not ( n245385 , n245384 );
or ( n245386 , n245375 , n245385 );
nand ( n245387 , n245383 , n235241 );
nand ( n245388 , n245386 , n245387 );
not ( n245389 , n245388 );
and ( n245390 , n245374 , n245389 );
and ( n245391 , n245373 , n245388 );
nor ( n245392 , n245390 , n245391 );
buf ( n245393 , n245392 );
and ( n245394 , n245340 , n245393 );
not ( n245395 , n245340 );
not ( n245396 , n245388 );
not ( n245397 , n245373 );
or ( n245398 , n245396 , n245397 );
not ( n245399 , n245373 );
not ( n245400 , n245388 );
nand ( n245401 , n245399 , n245400 );
nand ( n245402 , n245398 , n245401 );
buf ( n245403 , n245402 );
and ( n245404 , n245395 , n245403 );
nor ( n245405 , n245394 , n245404 );
not ( n245406 , n245405 );
nand ( n245407 , n245268 , n245406 );
or ( n245408 , n245242 , n245407 );
not ( n245409 , n245240 );
not ( n245410 , n245268 );
or ( n245411 , n245409 , n245410 );
nor ( n245412 , n245406 , n226003 );
nand ( n245413 , n245411 , n245412 );
buf ( n245414 , n35431 );
nand ( n245415 , n245414 , n25649 );
nand ( n245416 , n245408 , n245413 , n245415 );
buf ( n245417 , n245416 );
not ( n245418 , n237500 );
nand ( n245419 , n54417 , n54404 );
not ( n245420 , n245419 );
or ( n245421 , n245418 , n245420 );
or ( n245422 , n245419 , n237500 );
nand ( n245423 , n245421 , n245422 );
not ( n245424 , n245423 );
nand ( n245425 , n232134 , n232111 );
not ( n245426 , n245425 );
buf ( n245427 , n237473 );
not ( n245428 , n245427 );
and ( n245429 , n245426 , n245428 );
and ( n245430 , n245425 , n245427 );
nor ( n245431 , n245429 , n245430 );
not ( n245432 , n245431 );
or ( n245433 , n245424 , n245432 );
or ( n245434 , n245423 , n245431 );
nand ( n245435 , n245433 , n245434 );
not ( n245436 , n232191 );
nand ( n245437 , n245436 , n54452 );
and ( n245438 , n245437 , n241929 );
not ( n245439 , n245437 );
and ( n245440 , n245439 , n237520 );
nor ( n245441 , n245438 , n245440 );
and ( n245442 , n245435 , n245441 );
not ( n245443 , n245435 );
not ( n245444 , n245441 );
and ( n245445 , n245443 , n245444 );
nor ( n245446 , n245442 , n245445 );
not ( n245447 , n54522 );
not ( n245448 , n232272 );
nand ( n245449 , n245447 , n245448 );
not ( n245450 , n245449 );
not ( n245451 , n245450 );
not ( n245452 , n237564 );
or ( n245453 , n245451 , n245452 );
nand ( n245454 , n237565 , n245449 );
nand ( n245455 , n245453 , n245454 );
not ( n245456 , n232234 );
nand ( n245457 , n245456 , n232254 );
not ( n245458 , n245457 );
not ( n245459 , n237554 );
and ( n245460 , n245458 , n245459 );
and ( n245461 , n245457 , n237554 );
nor ( n245462 , n245460 , n245461 );
not ( n245463 , n245462 );
and ( n245464 , n245455 , n245463 );
not ( n245465 , n245455 );
and ( n245466 , n245465 , n245462 );
nor ( n245467 , n245464 , n245466 );
not ( n245468 , n245467 );
and ( n245469 , n245446 , n245468 );
not ( n245470 , n245446 );
and ( n245471 , n245470 , n245467 );
nor ( n245472 , n245469 , n245471 );
not ( n245473 , n245472 );
not ( n245474 , n245473 );
not ( n245475 , n245474 );
not ( n245476 , n232374 );
nand ( n245477 , n54596 , n232352 );
xnor ( n245478 , n245477 , n55040 );
not ( n245479 , n245478 );
not ( n245480 , n241902 );
or ( n245481 , n245479 , n245480 );
or ( n245482 , n241902 , n245478 );
nand ( n245483 , n245481 , n245482 );
not ( n245484 , n245483 );
nand ( n245485 , n232503 , n54572 );
not ( n245486 , n245485 );
not ( n245487 , n232698 );
and ( n245488 , n245486 , n245487 );
and ( n245489 , n245485 , n232698 );
nor ( n245490 , n245488 , n245489 );
not ( n245491 , n245490 );
nand ( n245492 , n54663 , n232445 );
and ( n245493 , n245492 , n232740 );
not ( n245494 , n245492 );
and ( n245495 , n245494 , n237407 );
nor ( n245496 , n245493 , n245495 );
not ( n245497 , n245496 );
or ( n245498 , n245491 , n245497 );
or ( n245499 , n245496 , n245490 );
nand ( n245500 , n245498 , n245499 );
not ( n245501 , n232462 );
nand ( n245502 , n245501 , n54725 );
not ( n245503 , n245502 );
not ( n245504 , n232720 );
and ( n245505 , n245503 , n245504 );
and ( n245506 , n245502 , n232720 );
nor ( n245507 , n245505 , n245506 );
and ( n245508 , n245500 , n245507 );
not ( n245509 , n245500 );
not ( n245510 , n245507 );
and ( n245511 , n245509 , n245510 );
nor ( n245512 , n245508 , n245511 );
not ( n245513 , n245512 );
or ( n245514 , n245484 , n245513 );
or ( n245515 , n245483 , n245512 );
nand ( n245516 , n245514 , n245515 );
buf ( n245517 , n245516 );
not ( n245518 , n245517 );
or ( n245519 , n245476 , n245518 );
or ( n245520 , n245517 , n232374 );
nand ( n245521 , n245519 , n245520 );
not ( n245522 , n245521 );
and ( n245523 , n245475 , n245522 );
not ( n245524 , n245473 );
and ( n245525 , n245524 , n245521 );
nor ( n245526 , n245523 , n245525 );
nor ( n245527 , n245526 , n47173 );
not ( n245528 , n30612 );
not ( n245529 , n54667 );
or ( n245530 , n245528 , n245529 );
not ( n245531 , n30612 );
nand ( n245532 , n245531 , n232427 );
nand ( n245533 , n245530 , n245532 );
not ( n245534 , n245533 );
not ( n245535 , n49132 );
not ( n245536 , n245535 );
and ( n245537 , n245534 , n245536 );
not ( n245538 , n225372 );
and ( n245539 , n245533 , n245538 );
nor ( n245540 , n245537 , n245539 );
nand ( n245541 , n240763 , n245540 );
and ( n245542 , n245541 , n37198 );
not ( n245543 , n245541 );
not ( n245544 , n37198 );
and ( n245545 , n245543 , n245544 );
nor ( n245546 , n245542 , n245545 );
not ( n245547 , n245546 );
not ( n245548 , n245547 );
xor ( n245549 , n34066 , n55941 );
xnor ( n245550 , n245549 , n41258 );
nand ( n245551 , n36971 , n245550 );
and ( n245552 , n245551 , n36986 );
not ( n245553 , n245551 );
and ( n245554 , n245553 , n36985 );
nor ( n245555 , n245552 , n245554 );
not ( n245556 , n245555 );
not ( n245557 , n245556 );
not ( n245558 , n33023 );
not ( n245559 , n213924 );
or ( n245560 , n245558 , n245559 );
or ( n245561 , n213924 , n33023 );
nand ( n245562 , n245560 , n245561 );
and ( n245563 , n245562 , n36190 );
not ( n245564 , n245562 );
and ( n245565 , n245564 , n36189 );
nor ( n245566 , n245563 , n245565 );
nand ( n245567 , n245566 , n36870 );
not ( n245568 , n245567 );
not ( n245569 , n36857 );
and ( n245570 , n245568 , n245569 );
and ( n245571 , n245567 , n36857 );
nor ( n245572 , n245570 , n245571 );
not ( n245573 , n245572 );
not ( n245574 , n245573 );
or ( n245575 , n245557 , n245574 );
nand ( n245576 , n245572 , n245555 );
nand ( n245577 , n245575 , n245576 );
not ( n245578 , n232894 );
not ( n245579 , n245540 );
nand ( n245580 , n245544 , n245579 );
not ( n245581 , n240751 );
and ( n245582 , n245580 , n245581 );
not ( n245583 , n245580 );
and ( n245584 , n245583 , n240751 );
nor ( n245585 , n245582 , n245584 );
not ( n245586 , n245585 );
not ( n245587 , n245586 );
or ( n245588 , n245578 , n245587 );
nand ( n245589 , n245585 , n232893 );
nand ( n245590 , n245588 , n245589 );
and ( n245591 , n245590 , n36777 );
not ( n245592 , n245590 );
and ( n245593 , n245592 , n37293 );
nor ( n245594 , n245591 , n245593 );
and ( n245595 , n245577 , n245594 );
not ( n245596 , n245577 );
and ( n245597 , n245590 , n37293 );
not ( n245598 , n245590 );
and ( n245599 , n245598 , n36777 );
nor ( n245600 , n245597 , n245599 );
and ( n245601 , n245596 , n245600 );
nor ( n245602 , n245595 , n245601 );
not ( n245603 , n245602 );
or ( n245604 , n245548 , n245603 );
not ( n245605 , n245547 );
not ( n245606 , n245600 );
not ( n245607 , n245577 );
not ( n245608 , n245607 );
or ( n245609 , n245606 , n245608 );
nand ( n245610 , n245577 , n245594 );
nand ( n245611 , n245609 , n245610 );
nand ( n245612 , n245605 , n245611 );
nand ( n245613 , n245604 , n245612 );
not ( n245614 , n240941 );
not ( n245615 , n245614 );
and ( n245616 , n245613 , n245615 );
not ( n245617 , n245613 );
buf ( n245618 , n240948 );
and ( n245619 , n245617 , n245618 );
nor ( n245620 , n245616 , n245619 );
not ( n245621 , n47000 );
nand ( n245622 , n245621 , n50888 );
and ( n245623 , n245622 , n47009 );
not ( n245624 , n245622 );
not ( n245625 , n47009 );
and ( n245626 , n245624 , n245625 );
nor ( n245627 , n245623 , n245626 );
buf ( n245628 , n245627 );
not ( n245629 , n245628 );
not ( n245630 , n224924 );
or ( n245631 , n245629 , n245630 );
not ( n245632 , n245628 );
nand ( n245633 , n245632 , n47156 );
nand ( n245634 , n245631 , n245633 );
not ( n245635 , n225257 );
nand ( n245636 , n226132 , n48380 );
not ( n245637 , n245636 );
or ( n245638 , n245635 , n245637 );
nand ( n245639 , n48380 , n226132 );
or ( n245640 , n245639 , n225257 );
nand ( n245641 , n245638 , n245640 );
not ( n245642 , n245641 );
not ( n245643 , n241393 );
or ( n245644 , n245642 , n245643 );
or ( n245645 , n241393 , n245641 );
nand ( n245646 , n245644 , n245645 );
not ( n245647 , n243681 );
not ( n245648 , n47446 );
not ( n245649 , n226110 );
nand ( n245650 , n245649 , n226099 );
not ( n245651 , n245650 );
or ( n245652 , n245648 , n245651 );
or ( n245653 , n245650 , n47446 );
nand ( n245654 , n245652 , n245653 );
not ( n245655 , n245654 );
or ( n245656 , n245647 , n245655 );
or ( n245657 , n245654 , n243681 );
nand ( n245658 , n245656 , n245657 );
not ( n245659 , n48319 );
nand ( n245660 , n245659 , n48267 );
not ( n245661 , n245660 );
buf ( n245662 , n225128 );
not ( n245663 , n245662 );
and ( n245664 , n245661 , n245663 );
and ( n245665 , n245660 , n245662 );
nor ( n245666 , n245664 , n245665 );
and ( n245667 , n245658 , n245666 );
not ( n245668 , n245658 );
not ( n245669 , n245666 );
and ( n245670 , n245668 , n245669 );
nor ( n245671 , n245667 , n245670 );
and ( n245672 , n245646 , n245671 );
not ( n245673 , n245646 );
not ( n245674 , n245671 );
and ( n245675 , n245673 , n245674 );
nor ( n245676 , n245672 , n245675 );
not ( n245677 , n245676 );
and ( n245678 , n245634 , n245677 );
not ( n245679 , n245634 );
not ( n245680 , n245677 );
and ( n245681 , n245679 , n245680 );
nor ( n245682 , n245678 , n245681 );
not ( n245683 , n245682 );
nand ( n245684 , n245527 , n245620 , n245683 );
not ( n245685 , n245526 );
not ( n245686 , n245685 );
not ( n245687 , n245683 );
or ( n245688 , n245686 , n245687 );
nor ( n245689 , n245620 , n37725 );
nand ( n245690 , n245688 , n245689 );
nand ( n245691 , n37728 , n214640 );
nand ( n245692 , n245684 , n245690 , n245691 );
buf ( n245693 , n245692 );
not ( n245694 , RI1754b800_32);
or ( n245695 , n229127 , n245694 );
not ( n245696 , RI19aac388_2481);
or ( n245697 , n25335 , n245696 );
nand ( n245698 , n245695 , n245697 );
buf ( n245699 , n245698 );
not ( n245700 , n41237 );
buf ( n245701 , n35431 );
buf ( n245702 , n245701 );
not ( n245703 , n245702 );
or ( n245704 , n245700 , n245703 );
not ( n245705 , n235759 );
nand ( n245706 , n52489 , n40012 );
not ( n245707 , n245706 );
not ( n245708 , n52492 );
and ( n245709 , n245707 , n245708 );
not ( n245710 , n40011 );
nand ( n245711 , n245710 , n52489 );
and ( n245712 , n245711 , n52492 );
nor ( n245713 , n245709 , n245712 );
or ( n245714 , n245713 , n52474 );
nand ( n245715 , n52474 , n245713 );
nand ( n245716 , n245714 , n245715 );
and ( n245717 , n245716 , n245250 );
not ( n245718 , n245716 );
and ( n245719 , n245718 , n245249 );
nor ( n245720 , n245717 , n245719 );
nand ( n245721 , n39880 , n52560 );
not ( n245722 , n245721 );
not ( n245723 , n39788 );
not ( n245724 , n245723 );
and ( n245725 , n245722 , n245724 );
and ( n245726 , n245721 , n245723 );
nor ( n245727 , n245725 , n245726 );
not ( n245728 , n245727 );
nand ( n245729 , n39862 , n52577 );
and ( n245730 , n245729 , n52590 );
not ( n245731 , n245729 );
and ( n245732 , n245731 , n52589 );
nor ( n245733 , n245730 , n245732 );
not ( n245734 , n245733 );
or ( n245735 , n245728 , n245734 );
or ( n245736 , n245733 , n245727 );
nand ( n245737 , n245735 , n245736 );
xnor ( n245738 , n245720 , n245737 );
not ( n245739 , n245738 );
or ( n245740 , n245705 , n245739 );
not ( n245741 , n235759 );
xor ( n245742 , n245248 , n245716 );
xnor ( n245743 , n245742 , n245737 );
nand ( n245744 , n245741 , n245743 );
nand ( n245745 , n245740 , n245744 );
nand ( n245746 , n40331 , n52637 );
not ( n245747 , n245746 );
not ( n245748 , n230387 );
and ( n245749 , n245747 , n245748 );
and ( n245750 , n245746 , n230387 );
nor ( n245751 , n245749 , n245750 );
not ( n245752 , n245751 );
nand ( n245753 , n217981 , n52660 );
and ( n245754 , n245753 , n52650 );
not ( n245755 , n245753 );
and ( n245756 , n245755 , n52649 );
nor ( n245757 , n245754 , n245756 );
not ( n245758 , n245757 );
or ( n245759 , n245752 , n245758 );
or ( n245760 , n245757 , n245751 );
nand ( n245761 , n245759 , n245760 );
not ( n245762 , n230434 );
nand ( n245763 , n245762 , n40290 );
not ( n245764 , n245763 );
not ( n245765 , n230444 );
not ( n245766 , n245765 );
and ( n245767 , n245764 , n245766 );
and ( n245768 , n245763 , n245765 );
nor ( n245769 , n245767 , n245768 );
not ( n245770 , n245769 );
and ( n245771 , n245761 , n245770 );
not ( n245772 , n245761 );
and ( n245773 , n245772 , n245769 );
nor ( n245774 , n245771 , n245773 );
nand ( n245775 , n52738 , n40446 );
not ( n245776 , n245775 );
not ( n245777 , n230488 );
and ( n245778 , n245776 , n245777 );
and ( n245779 , n245775 , n230488 );
nor ( n245780 , n245778 , n245779 );
nand ( n245781 , n230458 , n40374 );
and ( n245782 , n245781 , n52710 );
not ( n245783 , n245781 );
and ( n245784 , n245783 , n52709 );
nor ( n245785 , n245782 , n245784 );
xor ( n245786 , n245780 , n245785 );
and ( n245787 , n245774 , n245786 );
not ( n245788 , n245774 );
not ( n245789 , n245786 );
and ( n245790 , n245788 , n245789 );
nor ( n245791 , n245787 , n245790 );
not ( n245792 , n245791 );
not ( n245793 , n245792 );
not ( n245794 , n245793 );
and ( n245795 , n245745 , n245794 );
not ( n245796 , n245745 );
not ( n245797 , n245791 );
buf ( n245798 , n245797 );
not ( n245799 , n245798 );
and ( n245800 , n245796 , n245799 );
nor ( n245801 , n245795 , n245800 );
not ( n245802 , n245801 );
nand ( n245803 , n48248 , n245802 );
not ( n245804 , n49876 );
nand ( n245805 , n49872 , n49869 );
not ( n245806 , n245805 );
not ( n245807 , n39088 );
not ( n245808 , n245807 );
and ( n245809 , n245806 , n245808 );
and ( n245810 , n245805 , n245807 );
nor ( n245811 , n245809 , n245810 );
not ( n245812 , n245811 );
not ( n245813 , n39276 );
not ( n245814 , n245813 );
nand ( n245815 , n49892 , n39288 );
not ( n245816 , n245815 );
or ( n245817 , n245814 , n245816 );
or ( n245818 , n245813 , n245815 );
nand ( n245819 , n245817 , n245818 );
not ( n245820 , n245819 );
or ( n245821 , n245812 , n245820 );
or ( n245822 , n245819 , n245811 );
nand ( n245823 , n245821 , n245822 );
not ( n245824 , n39363 );
not ( n245825 , n227681 );
nand ( n245826 , n245824 , n245825 );
not ( n245827 , n245826 );
not ( n245828 , n39406 );
not ( n245829 , n245828 );
and ( n245830 , n245827 , n245829 );
and ( n245831 , n245826 , n245828 );
nor ( n245832 , n245830 , n245831 );
and ( n245833 , n245823 , n245832 );
not ( n245834 , n245823 );
not ( n245835 , n245832 );
and ( n245836 , n245834 , n245835 );
nor ( n245837 , n245833 , n245836 );
not ( n245838 , n245837 );
not ( n245839 , RI17537fd0_593);
and ( n245840 , n52537 , n245839 );
and ( n245841 , n245005 , n245840 , n204523 );
xor ( n245842 , n245841 , n39169 );
nor ( n245843 , n39180 , n227611 );
xnor ( n245844 , n245842 , n245843 );
not ( n245845 , n245844 );
not ( n245846 , n227568 );
nand ( n245847 , n245846 , n39147 );
not ( n245848 , n245847 );
buf ( n245849 , n39136 );
not ( n245850 , n245849 );
and ( n245851 , n245848 , n245850 );
and ( n245852 , n245847 , n245849 );
nor ( n245853 , n245851 , n245852 );
not ( n245854 , n245853 );
and ( n245855 , n245845 , n245854 );
and ( n245856 , n245844 , n245853 );
nor ( n245857 , n245855 , n245856 );
and ( n245858 , n245838 , n245857 );
not ( n245859 , n245838 );
not ( n245860 , n245857 );
and ( n245861 , n245859 , n245860 );
nor ( n245862 , n245858 , n245861 );
not ( n245863 , n245862 );
or ( n245864 , n245804 , n245863 );
not ( n245865 , n49876 );
not ( n245866 , n245857 );
not ( n245867 , n245837 );
not ( n245868 , n245867 );
or ( n245869 , n245866 , n245868 );
not ( n245870 , n245857 );
nand ( n245871 , n245870 , n245837 );
nand ( n245872 , n245869 , n245871 );
nand ( n245873 , n245865 , n245872 );
nand ( n245874 , n245864 , n245873 );
nand ( n245875 , n242836 , n52948 );
not ( n245876 , n245875 );
not ( n245877 , n52961 );
not ( n245878 , n245877 );
and ( n245879 , n245876 , n245878 );
and ( n245880 , n245875 , n245877 );
nor ( n245881 , n245879 , n245880 );
not ( n245882 , n245881 );
not ( n245883 , n52911 );
nand ( n245884 , n245883 , n242802 );
and ( n245885 , n245884 , n52922 );
not ( n245886 , n245884 );
and ( n245887 , n245886 , n52921 );
nor ( n245888 , n245885 , n245887 );
not ( n245889 , n245888 );
or ( n245890 , n245882 , n245889 );
or ( n245891 , n245888 , n245881 );
nand ( n245892 , n245890 , n245891 );
not ( n245893 , n245892 );
nand ( n245894 , n230571 , n242763 );
and ( n245895 , n245894 , n230582 );
not ( n245896 , n245894 );
and ( n245897 , n245896 , n52820 );
nor ( n245898 , n245895 , n245897 );
not ( n245899 , n245898 );
not ( n245900 , n245899 );
nand ( n245901 , n230623 , n242776 );
not ( n245902 , n245901 );
not ( n245903 , n242717 );
and ( n245904 , n245902 , n245903 );
and ( n245905 , n245901 , n242717 );
nor ( n245906 , n245904 , n245905 );
nor ( n245907 , n52798 , n245906 );
not ( n245908 , n245907 );
nand ( n245909 , n52798 , n245906 );
nand ( n245910 , n245908 , n245909 );
not ( n245911 , n245910 );
and ( n245912 , n245900 , n245911 );
and ( n245913 , n245899 , n245910 );
nor ( n245914 , n245912 , n245913 );
not ( n245915 , n245914 );
and ( n245916 , n245893 , n245915 );
and ( n245917 , n245892 , n245914 );
nor ( n245918 , n245916 , n245917 );
not ( n245919 , n245918 );
not ( n245920 , n245919 );
and ( n245921 , n245874 , n245920 );
not ( n245922 , n245874 );
not ( n245923 , n245914 );
not ( n245924 , n245923 );
not ( n245925 , n245892 );
not ( n245926 , n245925 );
or ( n245927 , n245924 , n245926 );
nand ( n245928 , n245914 , n245892 );
nand ( n245929 , n245927 , n245928 );
buf ( n245930 , n245929 );
and ( n245931 , n245922 , n245930 );
nor ( n245932 , n245921 , n245931 );
not ( n245933 , n245932 );
and ( n245934 , n245803 , n245933 );
not ( n245935 , n245803 );
and ( n245936 , n245935 , n245932 );
nor ( n245937 , n245934 , n245936 );
buf ( n245938 , n244216 );
or ( n245939 , n245937 , n245938 );
nand ( n245940 , n245704 , n245939 );
buf ( n245941 , n245940 );
not ( n245942 , n32306 );
buf ( n245943 , n239240 );
not ( n245944 , n245943 );
or ( n245945 , n245942 , n245944 );
and ( n245946 , n245005 , n204518 );
not ( n245947 , n245946 );
xor ( n245948 , n48355 , n226087 );
xnor ( n245949 , n245948 , n226169 );
not ( n245950 , n245949 );
not ( n245951 , n245950 );
not ( n245952 , n224801 );
nand ( n245953 , n245952 , n50917 );
not ( n245954 , n245953 );
not ( n245955 , n47052 );
and ( n245956 , n245954 , n245955 );
and ( n245957 , n245953 , n47052 );
nor ( n245958 , n245956 , n245957 );
not ( n245959 , n245958 );
not ( n245960 , n245627 );
or ( n245961 , n245959 , n245960 );
or ( n245962 , n245627 , n245958 );
nand ( n245963 , n245961 , n245962 );
not ( n245964 , n224723 );
nand ( n245965 , n245964 , n50863 );
not ( n245966 , n245965 );
not ( n245967 , n224736 );
not ( n245968 , n245967 );
and ( n245969 , n245966 , n245968 );
and ( n245970 , n245965 , n245967 );
nor ( n245971 , n245969 , n245970 );
and ( n245972 , n245963 , n245971 );
not ( n245973 , n245963 );
not ( n245974 , n245971 );
and ( n245975 , n245973 , n245974 );
nor ( n245976 , n245972 , n245975 );
nand ( n245977 , n224903 , n50789 );
not ( n245978 , n224875 );
xor ( n245979 , n245977 , n245978 );
not ( n245980 , n245979 );
nand ( n245981 , n50829 , n224851 );
and ( n245982 , n245981 , n47075 );
not ( n245983 , n245981 );
and ( n245984 , n245983 , n244517 );
nor ( n245985 , n245982 , n245984 );
not ( n245986 , n245985 );
or ( n245987 , n245980 , n245986 );
or ( n245988 , n245985 , n245979 );
nand ( n245989 , n245987 , n245988 );
and ( n245990 , n245976 , n245989 );
not ( n245991 , n245976 );
not ( n245992 , n245989 );
and ( n245993 , n245991 , n245992 );
nor ( n245994 , n245990 , n245993 );
not ( n245995 , n245994 );
not ( n245996 , n245995 );
nand ( n245997 , n50862 , n50849 );
nand ( n245998 , n204519 , n204522 );
not ( n245999 , n245998 );
and ( n246000 , n245997 , n245999 );
not ( n246001 , n245997 );
and ( n246002 , n246001 , n245998 );
nor ( n246003 , n246000 , n246002 );
and ( n246004 , n246003 , n224723 );
not ( n246005 , n246003 );
and ( n246006 , n246005 , n245964 );
nor ( n246007 , n246004 , n246006 );
not ( n246008 , n246007 );
not ( n246009 , n246008 );
and ( n246010 , n245996 , n246009 );
not ( n246011 , n245994 );
and ( n246012 , n246011 , n246008 );
nor ( n246013 , n246010 , n246012 );
not ( n246014 , n246013 );
or ( n246015 , n245951 , n246014 );
not ( n246016 , n246013 );
buf ( n246017 , n245949 );
nand ( n246018 , n246016 , n246017 );
nand ( n246019 , n246015 , n246018 );
not ( n246020 , n246019 );
or ( n246021 , n245947 , n246020 );
or ( n246022 , n246019 , n245946 );
nand ( n246023 , n246021 , n246022 );
not ( n246024 , n246023 );
and ( n246025 , n236760 , n236713 );
not ( n246026 , n236760 );
and ( n246027 , n246026 , n236712 );
nor ( n246028 , n246025 , n246027 );
nor ( n246029 , n246028 , n243730 );
not ( n246030 , n246029 );
nand ( n246031 , n243730 , n246028 );
nand ( n246032 , n246030 , n246031 );
not ( n246033 , n246032 );
not ( n246034 , n243876 );
nand ( n246035 , n246034 , n44878 );
not ( n246036 , n246035 );
not ( n246037 , n243968 );
and ( n246038 , n246036 , n246037 );
and ( n246039 , n246035 , n243968 );
nor ( n246040 , n246038 , n246039 );
not ( n246041 , n246040 );
nand ( n246042 , n222599 , n243892 );
and ( n246043 , n246042 , n44849 );
not ( n246044 , n246042 );
and ( n246045 , n246044 , n44848 );
nor ( n246046 , n246043 , n246045 );
not ( n246047 , n246046 );
or ( n246048 , n246041 , n246047 );
or ( n246049 , n246040 , n246046 );
nand ( n246050 , n246048 , n246049 );
nand ( n246051 , n44946 , n243923 );
not ( n246052 , n246051 );
not ( n246053 , n44942 );
and ( n246054 , n246052 , n246053 );
and ( n246055 , n246051 , n44942 );
nor ( n246056 , n246054 , n246055 );
and ( n246057 , n246050 , n246056 );
not ( n246058 , n246050 );
not ( n246059 , n246056 );
and ( n246060 , n246058 , n246059 );
nor ( n246061 , n246057 , n246060 );
xor ( n246062 , n44814 , n237963 );
not ( n246063 , n246062 );
xor ( n246064 , n246061 , n246063 );
buf ( n246065 , n246064 );
not ( n246066 , n246065 );
and ( n246067 , n246033 , n246066 );
and ( n246068 , n246032 , n246065 );
nor ( n246069 , n246067 , n246068 );
not ( n246070 , n43487 );
not ( n246071 , n238894 );
or ( n246072 , n246070 , n246071 );
not ( n246073 , n43487 );
and ( n246074 , n238859 , n238889 );
not ( n246075 , n238859 );
and ( n246076 , n246075 , n238890 );
nor ( n246077 , n246074 , n246076 );
nand ( n246078 , n246073 , n246077 );
nand ( n246079 , n246072 , n246078 );
and ( n246080 , n246079 , n244453 );
not ( n246081 , n246079 );
not ( n246082 , n244453 );
and ( n246083 , n246081 , n246082 );
nor ( n246084 , n246080 , n246083 );
not ( n246085 , n246084 );
nand ( n246086 , n246069 , n246085 );
not ( n246087 , n246086 );
and ( n246088 , n246024 , n246087 );
and ( n246089 , n246086 , n246023 );
nor ( n246090 , n246088 , n246089 );
not ( n246091 , n222532 );
or ( n246092 , n246090 , n246091 );
nand ( n246093 , n245945 , n246092 );
buf ( n246094 , n246093 );
not ( n246095 , RI19aa9f70_2496);
or ( n246096 , n233507 , n246095 );
not ( n246097 , RI19aa0358_2567);
or ( n246098 , n25336 , n246097 );
nand ( n246099 , n246096 , n246098 );
buf ( n246100 , n246099 );
not ( n246101 , n240474 );
not ( n246102 , n240634 );
nand ( n246103 , n246101 , n246102 );
and ( n246104 , n246103 , n240484 );
not ( n246105 , n246103 );
and ( n246106 , n246105 , n240483 );
nor ( n246107 , n246104 , n246106 );
buf ( n246108 , n246107 );
not ( n246109 , n246108 );
not ( n246110 , n240508 );
or ( n246111 , n246109 , n246110 );
or ( n246112 , n240508 , n246108 );
nand ( n246113 , n246111 , n246112 );
not ( n246114 , n36972 );
not ( n246115 , n245550 );
nand ( n246116 , n246115 , n240698 );
not ( n246117 , n246116 );
or ( n246118 , n246114 , n246117 );
not ( n246119 , n240698 );
not ( n246120 , n246119 );
nand ( n246121 , n246120 , n246115 );
or ( n246122 , n246121 , n36972 );
nand ( n246123 , n246118 , n246122 );
not ( n246124 , n246123 );
not ( n246125 , n245566 );
nand ( n246126 , n246125 , n240743 );
not ( n246127 , n246126 );
not ( n246128 , n36871 );
and ( n246129 , n246127 , n246128 );
not ( n246130 , n240740 );
nand ( n246131 , n246130 , n246125 );
and ( n246132 , n246131 , n36871 );
nor ( n246133 , n246129 , n246132 );
not ( n246134 , n246133 );
or ( n246135 , n246124 , n246134 );
or ( n246136 , n246123 , n246133 );
nand ( n246137 , n246135 , n246136 );
not ( n246138 , n246137 );
nand ( n246139 , n240783 , n55124 );
and ( n246140 , n246139 , n37139 );
not ( n246141 , n246139 );
and ( n246142 , n246141 , n37140 );
nor ( n246143 , n246140 , n246142 );
not ( n246144 , n246143 );
not ( n246145 , n246144 );
not ( n246146 , n245546 );
not ( n246147 , n246146 );
or ( n246148 , n246145 , n246147 );
nand ( n246149 , n245546 , n246143 );
nand ( n246150 , n246148 , n246149 );
nand ( n246151 , n36760 , n240717 );
not ( n246152 , n246151 );
not ( n246153 , n36744 );
and ( n246154 , n246152 , n246153 );
and ( n246155 , n246151 , n36744 );
nor ( n246156 , n246154 , n246155 );
and ( n246157 , n246150 , n246156 );
not ( n246158 , n246150 );
not ( n246159 , n246156 );
and ( n246160 , n246158 , n246159 );
nor ( n246161 , n246157 , n246160 );
not ( n246162 , n246161 );
and ( n246163 , n246138 , n246162 );
and ( n246164 , n246137 , n246161 );
nor ( n246165 , n246163 , n246164 );
buf ( n246166 , n246165 );
buf ( n246167 , n246166 );
not ( n246168 , n246167 );
and ( n246169 , n246113 , n246168 );
not ( n246170 , n246113 );
not ( n246171 , n246165 );
buf ( n246172 , n246171 );
not ( n246173 , n246172 );
and ( n246174 , n246170 , n246173 );
nor ( n246175 , n246169 , n246174 );
not ( n246176 , n246175 );
not ( n246177 , n49959 );
nand ( n246178 , n246176 , n246177 );
not ( n246179 , n54440 );
nand ( n246180 , n246179 , n241933 );
and ( n246181 , n246180 , n232191 );
not ( n246182 , n246180 );
and ( n246183 , n246182 , n245436 );
nor ( n246184 , n246181 , n246183 );
not ( n246185 , n246184 );
not ( n246186 , n246185 );
xor ( n246187 , n54457 , n54427 );
xnor ( n246188 , n246187 , n54531 );
not ( n246189 , n246188 );
or ( n246190 , n246186 , n246189 );
or ( n246191 , n246188 , n246185 );
nand ( n246192 , n246190 , n246191 );
buf ( n246193 , n244899 );
and ( n246194 , n246192 , n246193 );
not ( n246195 , n246192 );
buf ( n246196 , n244889 );
and ( n246197 , n246195 , n246196 );
nor ( n246198 , n246194 , n246197 );
not ( n246199 , n234862 );
not ( n246200 , n225525 );
or ( n246201 , n246199 , n246200 );
not ( n246202 , n234862 );
nand ( n246203 , n246202 , n47773 );
nand ( n246204 , n246201 , n246203 );
and ( n246205 , n246204 , n234437 );
not ( n246206 , n246204 );
buf ( n246207 , n239119 );
and ( n246208 , n246206 , n246207 );
nor ( n246209 , n246205 , n246208 );
nand ( n246210 , n246198 , n246209 );
or ( n246211 , n246178 , n246210 );
not ( n246212 , n246176 );
not ( n246213 , n246198 );
or ( n246214 , n246212 , n246213 );
nor ( n246215 , n246209 , n38637 );
nand ( n246216 , n246214 , n246215 );
buf ( n246217 , n35431 );
nand ( n246218 , n246217 , n26013 );
nand ( n246219 , n246211 , n246216 , n246218 );
buf ( n246220 , n246219 );
not ( n246221 , RI19ab36d8_2428);
or ( n246222 , n25328 , n246221 );
not ( n246223 , RI19aa9bb0_2498);
or ( n246224 , n25335 , n246223 );
nand ( n246225 , n246222 , n246224 );
buf ( n246226 , n246225 );
not ( n246227 , n240898 );
not ( n246228 , n37714 );
or ( n246229 , n246227 , n246228 );
not ( n246230 , n240898 );
nand ( n246231 , n246230 , n37708 );
nand ( n246232 , n246229 , n246231 );
not ( n246233 , n54134 );
and ( n246234 , n246232 , n246233 );
not ( n246235 , n246232 );
and ( n246236 , n246235 , n244802 );
nor ( n246237 , n246234 , n246236 );
nor ( n246238 , n246237 , n54208 );
not ( n246239 , n35899 );
not ( n246240 , n30853 );
or ( n246241 , n246239 , n246240 );
or ( n246242 , n30850 , n35899 );
nand ( n246243 , n246241 , n246242 );
and ( n246244 , n246243 , n30890 );
not ( n246245 , n246243 );
and ( n246246 , n246245 , n30893 );
nor ( n246247 , n246244 , n246246 );
buf ( n246248 , n31897 );
not ( n246249 , n246248 );
not ( n246250 , n205383 );
or ( n246251 , n246249 , n246250 );
not ( n246252 , n246248 );
nand ( n246253 , n246252 , n205384 );
nand ( n246254 , n246251 , n246253 );
and ( n246255 , n246254 , n30771 );
not ( n246256 , n246254 );
and ( n246257 , n246256 , n30757 );
nor ( n246258 , n246255 , n246257 );
nand ( n246259 , n246247 , n246258 );
not ( n246260 , n239572 );
and ( n246261 , n246259 , n246260 );
not ( n246262 , n246259 );
and ( n246263 , n246262 , n239572 );
nor ( n246264 , n246261 , n246263 );
not ( n246265 , n246264 );
not ( n246266 , n239466 );
xor ( n246267 , n39390 , n28721 );
xnor ( n246268 , n246267 , n30100 );
not ( n246269 , n246268 );
nand ( n246270 , n246266 , n246269 );
not ( n246271 , n246270 );
buf ( n246272 , n239455 );
not ( n246273 , n246272 );
and ( n246274 , n246271 , n246273 );
and ( n246275 , n246270 , n246272 );
nor ( n246276 , n246274 , n246275 );
not ( n246277 , n246276 );
not ( n246278 , n246277 );
not ( n246279 , n239424 );
or ( n246280 , n246278 , n246279 );
not ( n246281 , n239424 );
nand ( n246282 , n246281 , n246276 );
nand ( n246283 , n246280 , n246282 );
not ( n246284 , n246283 );
not ( n246285 , n244102 );
not ( n246286 , n239499 );
not ( n246287 , n55434 );
not ( n246288 , n37211 );
or ( n246289 , n246287 , n246288 );
or ( n246290 , n55434 , n35527 );
nand ( n246291 , n246289 , n246290 );
and ( n246292 , n246291 , n28463 );
not ( n246293 , n246291 );
and ( n246294 , n246293 , n28466 );
nor ( n246295 , n246292 , n246294 );
not ( n246296 , n246295 );
nand ( n246297 , n246286 , n246296 );
and ( n246298 , n246297 , n239505 );
not ( n246299 , n246297 );
not ( n246300 , n239505 );
and ( n246301 , n246299 , n246300 );
nor ( n246302 , n246298 , n246301 );
not ( n246303 , n246302 );
or ( n246304 , n246285 , n246303 );
or ( n246305 , n246302 , n244102 );
nand ( n246306 , n246304 , n246305 );
not ( n246307 , n246247 );
nand ( n246308 , n246260 , n246307 );
and ( n246309 , n246308 , n239583 );
not ( n246310 , n246308 );
and ( n246311 , n246310 , n239582 );
nor ( n246312 , n246309 , n246311 );
not ( n246313 , n246312 );
and ( n246314 , n246306 , n246313 );
not ( n246315 , n246306 );
and ( n246316 , n246315 , n246312 );
nor ( n246317 , n246314 , n246316 );
not ( n246318 , n246317 );
and ( n246319 , n246284 , n246318 );
and ( n246320 , n246283 , n246317 );
nor ( n246321 , n246319 , n246320 );
not ( n246322 , n246321 );
or ( n246323 , n246265 , n246322 );
or ( n246324 , n246317 , n246283 );
nand ( n246325 , n246283 , n246317 );
nand ( n246326 , n246324 , n246325 );
not ( n246327 , n246264 );
nand ( n246328 , n246326 , n246327 );
nand ( n246329 , n246323 , n246328 );
not ( n246330 , n246329 );
buf ( n246331 , n229300 );
not ( n246332 , n246331 );
and ( n246333 , n246330 , n246332 );
and ( n246334 , n246329 , n246331 );
nor ( n246335 , n246333 , n246334 );
not ( n246336 , n242041 );
not ( n246337 , n241303 );
nand ( n246338 , n245314 , n222136 );
not ( n246339 , n246338 );
or ( n246340 , n246337 , n246339 );
or ( n246341 , n246338 , n241303 );
nand ( n246342 , n246340 , n246341 );
not ( n246343 , n246342 );
nand ( n246344 , n242010 , n245299 );
not ( n246345 , n246344 );
not ( n246346 , n44432 );
not ( n246347 , n246346 );
and ( n246348 , n246345 , n246347 );
not ( n246349 , n242008 );
nand ( n246350 , n246349 , n242010 );
and ( n246351 , n246350 , n246346 );
nor ( n246352 , n246348 , n246351 );
not ( n246353 , n246352 );
or ( n246354 , n246343 , n246353 );
or ( n246355 , n246352 , n246342 );
nand ( n246356 , n246354 , n246355 );
not ( n246357 , n44460 );
nand ( n246358 , n246357 , n245293 );
and ( n246359 , n246358 , n241263 );
not ( n246360 , n246358 );
and ( n246361 , n246360 , n222229 );
nor ( n246362 , n246359 , n246361 );
and ( n246363 , n246356 , n246362 );
not ( n246364 , n246356 );
not ( n246365 , n246362 );
and ( n246366 , n246364 , n246365 );
nor ( n246367 , n246363 , n246366 );
not ( n246368 , n222252 );
nand ( n246369 , n246368 , n242053 );
not ( n246370 , n246369 );
not ( n246371 , n241326 );
and ( n246372 , n246370 , n246371 );
and ( n246373 , n246369 , n241326 );
nor ( n246374 , n246372 , n246373 );
not ( n246375 , n246374 );
not ( n246376 , n44363 );
or ( n246377 , n246375 , n246376 );
or ( n246378 , n44363 , n246374 );
nand ( n246379 , n246377 , n246378 );
not ( n246380 , n246379 );
and ( n246381 , n246367 , n246380 );
not ( n246382 , n246367 );
and ( n246383 , n246382 , n246379 );
nor ( n246384 , n246381 , n246383 );
not ( n246385 , n246384 );
not ( n246386 , n246385 );
or ( n246387 , n246336 , n246386 );
not ( n246388 , n242041 );
not ( n246389 , n246385 );
nand ( n246390 , n246388 , n246389 );
nand ( n246391 , n246387 , n246390 );
or ( n246392 , n245343 , n44604 );
xor ( n246393 , n246392 , n237793 );
not ( n246394 , n246393 );
not ( n246395 , n44644 );
nand ( n246396 , n44630 , n235237 );
not ( n246397 , n246396 );
or ( n246398 , n246395 , n246397 );
not ( n246399 , n246396 );
nand ( n246400 , n246399 , n44645 );
nand ( n246401 , n246398 , n246400 );
not ( n246402 , n246401 );
or ( n246403 , n246394 , n246402 );
or ( n246404 , n246401 , n246393 );
nand ( n246405 , n246403 , n246404 );
not ( n246406 , n246405 );
not ( n246407 , n44688 );
nand ( n246408 , n44700 , n235313 );
not ( n246409 , n246408 );
or ( n246410 , n246407 , n246409 );
or ( n246411 , n246408 , n44688 );
nand ( n246412 , n246410 , n246411 );
nand ( n246413 , n235282 , n44722 );
xor ( n246414 , n246413 , n44734 );
not ( n246415 , n246414 );
and ( n246416 , n246412 , n246415 );
not ( n246417 , n246412 );
and ( n246418 , n246417 , n246414 );
nor ( n246419 , n246416 , n246418 );
not ( n246420 , n246419 );
nand ( n246421 , n245379 , n235343 );
and ( n246422 , n246421 , n44568 );
not ( n246423 , n246421 );
and ( n246424 , n246423 , n222328 );
nor ( n246425 , n246422 , n246424 );
not ( n246426 , n246425 );
and ( n246427 , n246420 , n246426 );
and ( n246428 , n246419 , n246425 );
nor ( n246429 , n246427 , n246428 );
not ( n246430 , n246429 );
or ( n246431 , n246406 , n246430 );
not ( n246432 , n246429 );
not ( n246433 , n246401 );
not ( n246434 , n246393 );
and ( n246435 , n246433 , n246434 );
and ( n246436 , n246401 , n246393 );
nor ( n246437 , n246435 , n246436 );
nand ( n246438 , n246432 , n246437 );
nand ( n246439 , n246431 , n246438 );
not ( n246440 , n246439 );
not ( n246441 , n246440 );
and ( n246442 , n246391 , n246441 );
not ( n246443 , n246391 );
not ( n246444 , n246429 );
and ( n246445 , n246444 , n246437 );
not ( n246446 , n246444 );
and ( n246447 , n246446 , n246405 );
nor ( n246448 , n246445 , n246447 );
buf ( n246449 , n246448 );
and ( n246450 , n246443 , n246449 );
nor ( n246451 , n246442 , n246450 );
not ( n246452 , n246451 );
nand ( n246453 , n246238 , n246335 , n246452 );
not ( n246454 , n246237 );
not ( n246455 , n246454 );
not ( n246456 , n246335 );
or ( n246457 , n246455 , n246456 );
nor ( n246458 , n246452 , n53680 );
nand ( n246459 , n246457 , n246458 );
buf ( n246460 , n35431 );
nand ( n246461 , n246460 , n204995 );
nand ( n246462 , n246453 , n246459 , n246461 );
buf ( n246463 , n246462 );
not ( n246464 , RI19aa2e78_2546);
or ( n246465 , n25328 , n246464 );
not ( n246466 , RI19a99440_2617);
or ( n246467 , n226822 , n246466 );
nand ( n246468 , n246465 , n246467 );
buf ( n246469 , n246468 );
not ( n246470 , n49043 );
not ( n246471 , n50016 );
not ( n246472 , n48875 );
or ( n246473 , n246471 , n246472 );
nand ( n246474 , n48883 , n50019 );
nand ( n246475 , n246473 , n246474 );
not ( n246476 , n246475 );
or ( n246477 , n246470 , n246476 );
not ( n246478 , n49043 );
not ( n246479 , n246478 );
or ( n246480 , n246475 , n246479 );
nand ( n246481 , n246477 , n246480 );
not ( n246482 , n246481 );
not ( n246483 , n31909 );
nand ( n246484 , n246483 , n51182 );
not ( n246485 , n246484 );
not ( n246486 , n236461 );
and ( n246487 , n246485 , n246486 );
not ( n246488 , n31909 );
nand ( n246489 , n246488 , n51182 );
and ( n246490 , n246489 , n236461 );
nor ( n246491 , n246487 , n246490 );
not ( n246492 , n246491 );
not ( n246493 , n246492 );
not ( n246494 , n236461 );
nand ( n246495 , n246494 , n228944 );
not ( n246496 , n246495 );
not ( n246497 , n31789 );
and ( n246498 , n246496 , n246497 );
not ( n246499 , n236461 );
nand ( n246500 , n246499 , n228944 );
and ( n246501 , n246500 , n31789 );
nor ( n246502 , n246498 , n246501 );
not ( n246503 , n246502 );
not ( n246504 , n246503 );
not ( n246505 , n31615 );
nand ( n246506 , n246505 , n51200 );
and ( n246507 , n246506 , n31683 );
not ( n246508 , n246506 );
and ( n246509 , n246508 , n31682 );
nor ( n246510 , n246507 , n246509 );
not ( n246511 , n246510 );
not ( n246512 , n246511 );
or ( n246513 , n246504 , n246512 );
nand ( n246514 , n246510 , n246502 );
nand ( n246515 , n246513 , n246514 );
not ( n246516 , n51208 );
not ( n246517 , n236481 );
nand ( n246518 , n246516 , n246517 );
not ( n246519 , n246518 );
not ( n246520 , n32014 );
and ( n246521 , n246519 , n246520 );
and ( n246522 , n246518 , n32014 );
nor ( n246523 , n246521 , n246522 );
not ( n246524 , n246523 );
and ( n246525 , n246515 , n246524 );
not ( n246526 , n246515 );
and ( n246527 , n246526 , n246523 );
nor ( n246528 , n246525 , n246527 );
not ( n246529 , n236422 );
nand ( n246530 , n246529 , n51236 );
not ( n246531 , n246530 );
not ( n246532 , n32459 );
and ( n246533 , n246531 , n246532 );
and ( n246534 , n246530 , n32459 );
nor ( n246535 , n246533 , n246534 );
nand ( n246536 , n236437 , n51257 );
not ( n246537 , n246536 );
not ( n246538 , n32329 );
and ( n246539 , n246537 , n246538 );
and ( n246540 , n246536 , n32329 );
nor ( n246541 , n246539 , n246540 );
not ( n246542 , n246541 );
and ( n246543 , n246535 , n246542 );
not ( n246544 , n246535 );
and ( n246545 , n246544 , n246541 );
nor ( n246546 , n246543 , n246545 );
buf ( n246547 , n246546 );
xor ( n246548 , n246528 , n246547 );
not ( n246549 , n246548 );
or ( n246550 , n246493 , n246549 );
not ( n246551 , n246492 );
xor ( n246552 , n246523 , n246515 );
xor ( n246553 , n246552 , n246546 );
nand ( n246554 , n246551 , n246553 );
nand ( n246555 , n246550 , n246554 );
not ( n246556 , n33612 );
not ( n246557 , n44239 );
or ( n246558 , n246556 , n246557 );
not ( n246559 , n33612 );
nand ( n246560 , n246559 , n222159 );
nand ( n246561 , n246558 , n246560 );
and ( n246562 , n246561 , n210046 );
not ( n246563 , n246561 );
and ( n246564 , n246563 , n32280 );
nor ( n246565 , n246562 , n246564 );
not ( n246566 , n246565 );
nand ( n246567 , n246566 , n53217 );
buf ( n246568 , n32990 );
xor ( n246569 , n246567 , n246568 );
xor ( n246570 , n29452 , n25827 );
xnor ( n246571 , n246570 , n33404 );
not ( n246572 , n246571 );
nand ( n246573 , n246572 , n53233 );
not ( n246574 , n246573 );
not ( n246575 , n33145 );
and ( n246576 , n246574 , n246575 );
and ( n246577 , n246573 , n33145 );
nor ( n246578 , n246576 , n246577 );
and ( n246579 , n246569 , n246578 );
not ( n246580 , n246569 );
not ( n246581 , n246578 );
and ( n246582 , n246580 , n246581 );
nor ( n246583 , n246579 , n246582 );
not ( n246584 , n246583 );
not ( n246585 , n29991 );
buf ( n246586 , n208936 );
and ( n246587 , n246586 , n42285 );
not ( n246588 , n246586 );
and ( n246589 , n246588 , n220896 );
nor ( n246590 , n246587 , n246589 );
not ( n246591 , n246590 );
or ( n246592 , n246585 , n246591 );
or ( n246593 , n246590 , n29991 );
nand ( n246594 , n246592 , n246593 );
not ( n246595 , n246594 );
nand ( n246596 , n246595 , n230953 );
not ( n246597 , n246596 );
not ( n246598 , n32865 );
and ( n246599 , n246597 , n246598 );
and ( n246600 , n246596 , n32865 );
nor ( n246601 , n246599 , n246600 );
not ( n246602 , n246601 );
not ( n246603 , n32530 );
buf ( n246604 , n205382 );
not ( n246605 , n246604 );
not ( n246606 , n42113 );
or ( n246607 , n246605 , n246606 );
not ( n246608 , n246604 );
nand ( n246609 , n246608 , n31672 );
nand ( n246610 , n246607 , n246609 );
and ( n246611 , n246610 , n31637 );
not ( n246612 , n246610 );
and ( n246613 , n246612 , n219329 );
nor ( n246614 , n246611 , n246613 );
nand ( n246615 , n230920 , n246614 );
not ( n246616 , n246615 );
or ( n246617 , n246603 , n246616 );
or ( n246618 , n246615 , n32530 );
nand ( n246619 , n246617 , n246618 );
not ( n246620 , n246619 );
not ( n246621 , n33879 );
not ( n246622 , n205219 );
or ( n246623 , n246621 , n246622 );
not ( n246624 , n33879 );
nand ( n246625 , n246624 , n205214 );
nand ( n246626 , n246623 , n246625 );
and ( n246627 , n246626 , n43913 );
not ( n246628 , n246626 );
and ( n246629 , n246628 , n35200 );
nor ( n246630 , n246627 , n246629 );
not ( n246631 , n246630 );
nand ( n246632 , n246631 , n230941 );
not ( n246633 , n246632 );
not ( n246634 , n32692 );
and ( n246635 , n246633 , n246634 );
not ( n246636 , n246630 );
nand ( n246637 , n246636 , n230941 );
and ( n246638 , n246637 , n32692 );
nor ( n246639 , n246635 , n246638 );
not ( n246640 , n246639 );
or ( n246641 , n246620 , n246640 );
or ( n246642 , n246639 , n246619 );
nand ( n246643 , n246641 , n246642 );
not ( n246644 , n246643 );
or ( n246645 , n246602 , n246644 );
or ( n246646 , n246601 , n246643 );
nand ( n246647 , n246645 , n246646 );
not ( n246648 , n246647 );
or ( n246649 , n246584 , n246648 );
not ( n246650 , n246647 );
not ( n246651 , n246583 );
nand ( n246652 , n246650 , n246651 );
nand ( n246653 , n246649 , n246652 );
buf ( n246654 , n246653 );
and ( n246655 , n246555 , n246654 );
not ( n246656 , n246555 );
and ( n246657 , n246647 , n246583 );
not ( n246658 , n246647 );
and ( n246659 , n246658 , n246651 );
nor ( n246660 , n246657 , n246659 );
buf ( n246661 , n246660 );
and ( n246662 , n246656 , n246661 );
nor ( n246663 , n246655 , n246662 );
nand ( n246664 , n246482 , n246663 );
not ( n246665 , n43445 );
not ( n246666 , n238894 );
or ( n246667 , n246665 , n246666 );
not ( n246668 , n43445 );
nand ( n246669 , n246668 , n246077 );
nand ( n246670 , n246667 , n246669 );
not ( n246671 , n244453 );
and ( n246672 , n246670 , n246671 );
not ( n246673 , n246670 );
and ( n246674 , n246673 , n244453 );
nor ( n246675 , n246672 , n246674 );
nor ( n246676 , n246675 , n31571 );
not ( n246677 , n246676 );
or ( n246678 , n246664 , n246677 );
not ( n246679 , n246675 );
buf ( n246680 , n233971 );
nor ( n246681 , n246679 , n246680 );
nand ( n246682 , n246664 , n246681 );
nand ( n246683 , n234448 , n37036 );
nand ( n246684 , n246678 , n246682 , n246683 );
buf ( n246685 , n246684 );
not ( n246686 , n241555 );
not ( n246687 , n243372 );
or ( n246688 , n246686 , n246687 );
or ( n246689 , n243372 , n241555 );
nand ( n246690 , n246688 , n246689 );
and ( n246691 , n246690 , n243416 );
not ( n246692 , n246690 );
not ( n246693 , n243415 );
buf ( n246694 , n246693 );
and ( n246695 , n246692 , n246694 );
nor ( n246696 , n246691 , n246695 );
not ( n246697 , n52445 );
nand ( n246698 , n246696 , n246697 );
not ( n246699 , n243855 );
not ( n246700 , n246062 );
not ( n246701 , n246061 );
not ( n246702 , n246701 );
or ( n246703 , n246700 , n246702 );
nand ( n246704 , n246061 , n246063 );
nand ( n246705 , n246703 , n246704 );
not ( n246706 , n246705 );
or ( n246707 , n246699 , n246706 );
or ( n246708 , n246705 , n243855 );
nand ( n246709 , n246707 , n246708 );
not ( n246710 , n232528 );
not ( n246711 , n45080 );
nand ( n246712 , n246711 , n232664 );
not ( n246713 , n246712 );
or ( n246714 , n246710 , n246713 );
not ( n246715 , n45080 );
nand ( n246716 , n246715 , n232664 );
or ( n246717 , n246716 , n232528 );
nand ( n246718 , n246714 , n246717 );
not ( n246719 , n246718 );
not ( n246720 , n45063 );
nand ( n246721 , n246720 , n232640 );
not ( n246722 , n246721 );
not ( n246723 , n45051 );
and ( n246724 , n246722 , n246723 );
not ( n246725 , n45063 );
nand ( n246726 , n246725 , n232640 );
and ( n246727 , n246726 , n45051 );
nor ( n246728 , n246724 , n246727 );
not ( n246729 , n246728 );
and ( n246730 , n246719 , n246729 );
and ( n246731 , n246718 , n246728 );
nor ( n246732 , n246730 , n246731 );
not ( n246733 , n246732 );
nand ( n246734 , n222877 , n232555 );
not ( n246735 , n246734 );
not ( n246736 , n45127 );
and ( n246737 , n246735 , n246736 );
and ( n246738 , n246734 , n45127 );
nor ( n246739 , n246737 , n246738 );
not ( n246740 , n222981 );
nand ( n246741 , n222996 , n54868 );
not ( n246742 , n246741 );
or ( n246743 , n246740 , n246742 );
or ( n246744 , n246741 , n222981 );
nand ( n246745 , n246743 , n246744 );
xor ( n246746 , n246739 , n246745 );
not ( n246747 , n45159 );
nand ( n246748 , n246747 , n232594 );
and ( n246749 , n246748 , n222930 );
not ( n246750 , n246748 );
and ( n246751 , n246750 , n244022 );
nor ( n246752 , n246749 , n246751 );
xnor ( n246753 , n246746 , n246752 );
not ( n246754 , n246753 );
or ( n246755 , n246733 , n246754 );
not ( n246756 , n246753 );
not ( n246757 , n246732 );
nand ( n246758 , n246756 , n246757 );
nand ( n246759 , n246755 , n246758 );
buf ( n246760 , n246759 );
and ( n246761 , n246709 , n246760 );
not ( n246762 , n246709 );
and ( n246763 , n246756 , n246757 );
not ( n246764 , n246756 );
not ( n246765 , n246757 );
and ( n246766 , n246764 , n246765 );
nor ( n246767 , n246763 , n246766 );
buf ( n246768 , n246767 );
and ( n246769 , n246762 , n246768 );
nor ( n246770 , n246761 , n246769 );
not ( n246771 , n246770 );
not ( n246772 , n39426 );
not ( n246773 , n246772 );
nand ( n246774 , n39116 , n39136 );
not ( n246775 , n246774 );
not ( n246776 , n227577 );
and ( n246777 , n246775 , n246776 );
nand ( n246778 , n39116 , n245849 );
and ( n246779 , n246778 , n227577 );
nor ( n246780 , n246777 , n246779 );
not ( n246781 , n246780 );
not ( n246782 , n39253 );
nand ( n246783 , n246782 , n39169 );
and ( n246784 , n246783 , n227595 );
not ( n246785 , n246783 );
and ( n246786 , n246785 , n227596 );
nor ( n246787 , n246784 , n246786 );
not ( n246788 , n246787 );
or ( n246789 , n246781 , n246788 );
or ( n246790 , n246787 , n246780 );
nand ( n246791 , n246789 , n246790 );
not ( n246792 , n39101 );
nand ( n246793 , n246792 , n245807 );
and ( n246794 , n246793 , n242900 );
not ( n246795 , n246793 );
and ( n246796 , n246795 , n49860 );
nor ( n246797 , n246794 , n246796 );
not ( n246798 , n246797 );
and ( n246799 , n246791 , n246798 );
not ( n246800 , n246791 );
and ( n246801 , n246800 , n246797 );
nor ( n246802 , n246799 , n246801 );
not ( n246803 , n246802 );
not ( n246804 , n49931 );
not ( n246805 , n39419 );
nand ( n246806 , n246805 , n39422 );
not ( n246807 , n246806 );
or ( n246808 , n246804 , n246807 );
or ( n246809 , n49931 , n246806 );
nand ( n246810 , n246808 , n246809 );
nand ( n246811 , n39329 , n245813 );
not ( n246812 , n246811 );
not ( n246813 , n49903 );
and ( n246814 , n246812 , n246813 );
and ( n246815 , n246811 , n49903 );
nor ( n246816 , n246814 , n246815 );
and ( n246817 , n246810 , n246816 );
not ( n246818 , n246810 );
not ( n246819 , n246816 );
and ( n246820 , n246818 , n246819 );
nor ( n246821 , n246817 , n246820 );
not ( n246822 , n246821 );
not ( n246823 , n246822 );
and ( n246824 , n246803 , n246823 );
and ( n246825 , n246822 , n246802 );
nor ( n246826 , n246824 , n246825 );
not ( n246827 , n246826 );
or ( n246828 , n246773 , n246827 );
not ( n246829 , n246772 );
not ( n246830 , n246822 );
not ( n246831 , n246802 );
or ( n246832 , n246830 , n246831 );
not ( n246833 , n246802 );
nand ( n246834 , n246833 , n246821 );
nand ( n246835 , n246832 , n246834 );
nand ( n246836 , n246829 , n246835 );
nand ( n246837 , n246828 , n246836 );
nand ( n246838 , n230595 , n52820 );
not ( n246839 , n246838 );
not ( n246840 , n242932 );
and ( n246841 , n246839 , n246840 );
and ( n246842 , n246838 , n242932 );
nor ( n246843 , n246841 , n246842 );
not ( n246844 , n246843 );
nand ( n246845 , n52921 , n52935 );
xor ( n246846 , n242798 , n246845 );
not ( n246847 , n246846 );
or ( n246848 , n246844 , n246847 );
or ( n246849 , n246846 , n246843 );
nand ( n246850 , n246848 , n246849 );
nand ( n246851 , n52969 , n245877 );
buf ( n246852 , n242824 );
not ( n246853 , n246852 );
and ( n246854 , n246851 , n246853 );
not ( n246855 , n246851 );
and ( n246856 , n246855 , n246852 );
nor ( n246857 , n246854 , n246856 );
and ( n246858 , n246850 , n246857 );
not ( n246859 , n246850 );
not ( n246860 , n246857 );
and ( n246861 , n246859 , n246860 );
nor ( n246862 , n246858 , n246861 );
not ( n246863 , n246862 );
not ( n246864 , n246863 );
not ( n246865 , n52886 );
nand ( n246866 , n246865 , n230533 );
not ( n246867 , n246866 );
buf ( n246868 , n242734 );
not ( n246869 , n246868 );
and ( n246870 , n246867 , n246869 );
and ( n246871 , n246866 , n246868 );
nor ( n246872 , n246870 , n246871 );
not ( n246873 , n246872 );
not ( n246874 , n242722 );
and ( n246875 , n246873 , n246874 );
and ( n246876 , n246872 , n242722 );
nor ( n246877 , n246875 , n246876 );
not ( n246878 , n246877 );
not ( n246879 , n246878 );
and ( n246880 , n246864 , n246879 );
and ( n246881 , n246863 , n246878 );
nor ( n246882 , n246880 , n246881 );
buf ( n246883 , n246882 );
and ( n246884 , n246837 , n246883 );
not ( n246885 , n246837 );
not ( n246886 , n246877 );
not ( n246887 , n246862 );
or ( n246888 , n246886 , n246887 );
not ( n246889 , n246877 );
nand ( n246890 , n246889 , n246863 );
nand ( n246891 , n246888 , n246890 );
buf ( n246892 , n246891 );
and ( n246893 , n246885 , n246892 );
nor ( n246894 , n246884 , n246893 );
not ( n246895 , n246894 );
nand ( n246896 , n246771 , n246895 );
or ( n246897 , n246698 , n246896 );
nor ( n246898 , n246696 , n40465 );
nand ( n246899 , n246898 , n246896 );
nand ( n246900 , n241378 , n34605 );
nand ( n246901 , n246897 , n246899 , n246900 );
buf ( n246902 , n246901 );
not ( n246903 , n30703 );
not ( n246904 , n246903 );
not ( n246905 , n30811 );
not ( n246906 , n30895 );
nand ( n246907 , n246905 , n246906 );
not ( n246908 , n246907 );
buf ( n246909 , n229472 );
not ( n246910 , n246909 );
and ( n246911 , n246908 , n246910 );
and ( n246912 , n246907 , n246909 );
nor ( n246913 , n246911 , n246912 );
not ( n246914 , n246913 );
not ( n246915 , n30209 );
nand ( n246916 , n246915 , n207903 );
not ( n246917 , n246916 );
not ( n246918 , n229422 );
and ( n246919 , n246917 , n246918 );
and ( n246920 , n246916 , n229422 );
nor ( n246921 , n246919 , n246920 );
not ( n246922 , n246921 );
nand ( n246923 , n245004 , n245840 , n35627 );
not ( n246924 , n246923 );
and ( n246925 , n229394 , n246924 );
not ( n246926 , n229394 );
and ( n246927 , n246926 , n246923 );
nor ( n246928 , n246925 , n246927 );
not ( n246929 , n30452 );
not ( n246930 , n30369 );
nand ( n246931 , n246929 , n246930 );
and ( n246932 , n246928 , n246931 );
not ( n246933 , n246928 );
nor ( n246934 , n30452 , n30369 );
and ( n246935 , n246933 , n246934 );
nor ( n246936 , n246932 , n246935 );
not ( n246937 , n246936 );
and ( n246938 , n246922 , n246937 );
and ( n246939 , n246921 , n246936 );
nor ( n246940 , n246938 , n246939 );
not ( n246941 , n246940 );
xor ( n246942 , n246914 , n246941 );
nand ( n246943 , n30696 , n30545 );
not ( n246944 , n246943 );
not ( n246945 , n51687 );
not ( n246946 , n246945 );
and ( n246947 , n246944 , n246946 );
and ( n246948 , n246943 , n246945 );
nor ( n246949 , n246947 , n246948 );
not ( n246950 , n246949 );
not ( n246951 , n246950 );
nand ( n246952 , n30104 , n30773 );
not ( n246953 , n51730 );
and ( n246954 , n246952 , n246953 );
not ( n246955 , n246952 );
and ( n246956 , n246955 , n51730 );
nor ( n246957 , n246954 , n246956 );
not ( n246958 , n246957 );
not ( n246959 , n246958 );
or ( n246960 , n246951 , n246959 );
nand ( n246961 , n246957 , n246949 );
nand ( n246962 , n246960 , n246961 );
xnor ( n246963 , n246942 , n246962 );
not ( n246964 , n246963 );
or ( n246965 , n246904 , n246964 );
not ( n246966 , n246903 );
xor ( n246967 , n246913 , n246962 );
xor ( n246968 , n246967 , n246940 );
nand ( n246969 , n246966 , n246968 );
nand ( n246970 , n246965 , n246969 );
nand ( n246971 , n31530 , n25600 );
not ( n246972 , n246971 );
not ( n246973 , n26426 );
and ( n246974 , n246972 , n246973 );
and ( n246975 , n246971 , n26426 );
nor ( n246976 , n246974 , n246975 );
not ( n246977 , n246976 );
not ( n246978 , n242099 );
or ( n246979 , n246977 , n246978 );
or ( n246980 , n242099 , n246976 );
nand ( n246981 , n246979 , n246980 );
not ( n246982 , n246981 );
nand ( n246983 , n31275 , n50559 );
xnor ( n246984 , n246983 , n242101 );
not ( n246985 , n246984 );
or ( n246986 , n246982 , n246985 );
or ( n246987 , n246984 , n246981 );
nand ( n246988 , n246986 , n246987 );
not ( n246989 , n246988 );
not ( n246990 , n208778 );
nand ( n246991 , n246990 , n31083 );
not ( n246992 , n246991 );
not ( n246993 , n26057 );
and ( n246994 , n246992 , n246993 );
not ( n246995 , n242134 );
and ( n246996 , n246991 , n246995 );
nor ( n246997 , n246994 , n246996 );
not ( n246998 , n246997 );
nand ( n246999 , n31214 , n31139 );
and ( n247000 , n246999 , n26321 );
not ( n247001 , n246999 );
and ( n247002 , n247001 , n26322 );
nor ( n247003 , n247000 , n247002 );
not ( n247004 , n247003 );
or ( n247005 , n246998 , n247004 );
or ( n247006 , n246997 , n247003 );
nand ( n247007 , n247005 , n247006 );
not ( n247008 , n247007 );
not ( n247009 , n247008 );
or ( n247010 , n246989 , n247009 );
not ( n247011 , n246988 );
nand ( n247012 , n247011 , n247007 );
nand ( n247013 , n247010 , n247012 );
buf ( n247014 , n247013 );
and ( n247015 , n246970 , n247014 );
not ( n247016 , n246970 );
buf ( n247017 , n246988 );
xor ( n247018 , n247017 , n247008 );
buf ( n247019 , n247018 );
and ( n247020 , n247016 , n247019 );
nor ( n247021 , n247015 , n247020 );
not ( n247022 , n247021 );
not ( n247023 , n227002 );
not ( n247024 , n49232 );
nand ( n247025 , n247024 , n49218 );
not ( n247026 , n42207 );
and ( n247027 , n34218 , n40541 );
not ( n247028 , n34218 );
and ( n247029 , n247028 , n40538 );
nor ( n247030 , n247027 , n247029 );
not ( n247031 , n247030 );
and ( n247032 , n247026 , n247031 );
and ( n247033 , n42207 , n247030 );
nor ( n247034 , n247032 , n247033 );
and ( n247035 , n247025 , n247034 );
not ( n247036 , n247025 );
not ( n247037 , n247034 );
and ( n247038 , n247036 , n247037 );
nor ( n247039 , n247035 , n247038 );
not ( n247040 , n247039 );
not ( n247041 , n247040 );
not ( n247042 , n49261 );
nand ( n247043 , n247042 , n227005 );
not ( n247044 , n247043 );
xor ( n247045 , n47601 , n28877 );
xnor ( n247046 , n247045 , n25683 );
not ( n247047 , n247046 );
not ( n247048 , n247047 );
and ( n247049 , n247044 , n247048 );
not ( n247050 , n49261 );
nand ( n247051 , n247050 , n227005 );
and ( n247052 , n247051 , n247047 );
nor ( n247053 , n247049 , n247052 );
not ( n247054 , n247053 );
not ( n247055 , n247054 );
or ( n247056 , n247041 , n247055 );
nand ( n247057 , n247053 , n247039 );
nand ( n247058 , n247056 , n247057 );
nand ( n247059 , n227130 , n227159 );
not ( n247060 , n247059 );
not ( n247061 , n32418 );
not ( n247062 , n233666 );
or ( n247063 , n247061 , n247062 );
not ( n247064 , n233665 );
or ( n247065 , n247064 , n32418 );
nand ( n247066 , n247063 , n247065 );
and ( n247067 , n247066 , n48780 );
not ( n247068 , n247066 );
and ( n247069 , n247068 , n33565 );
nor ( n247070 , n247067 , n247069 );
not ( n247071 , n247070 );
and ( n247072 , n247060 , n247071 );
buf ( n247073 , n247070 );
and ( n247074 , n247059 , n247073 );
nor ( n247075 , n247072 , n247074 );
not ( n247076 , n247075 );
nand ( n247077 , n49347 , n227081 );
not ( n247078 , n33095 );
not ( n247079 , n44121 );
and ( n247080 , n247078 , n247079 );
and ( n247081 , n33095 , n44121 );
nor ( n247082 , n247080 , n247081 );
and ( n247083 , n247082 , n41063 );
not ( n247084 , n247082 );
and ( n247085 , n247084 , n33141 );
nor ( n247086 , n247083 , n247085 );
not ( n247087 , n247086 );
and ( n247088 , n247077 , n247087 );
not ( n247089 , n247077 );
and ( n247090 , n247089 , n247086 );
nor ( n247091 , n247088 , n247090 );
not ( n247092 , n247091 );
or ( n247093 , n247076 , n247092 );
or ( n247094 , n247075 , n247091 );
nand ( n247095 , n247093 , n247094 );
not ( n247096 , n49282 );
nand ( n247097 , n247096 , n49302 );
buf ( n247098 , RI17453e80_1327);
not ( n247099 , n247098 );
not ( n247100 , n25771 );
or ( n247101 , n247099 , n247100 );
not ( n247102 , n247098 );
nand ( n247103 , n247102 , n25772 );
nand ( n247104 , n247101 , n247103 );
and ( n247105 , n247104 , n44352 );
not ( n247106 , n247104 );
and ( n247107 , n247106 , n44348 );
nor ( n247108 , n247105 , n247107 );
xnor ( n247109 , n247097 , n247108 );
not ( n247110 , n247109 );
and ( n247111 , n247095 , n247110 );
not ( n247112 , n247095 );
and ( n247113 , n247112 , n247109 );
nor ( n247114 , n247111 , n247113 );
and ( n247115 , n247058 , n247114 );
not ( n247116 , n247058 );
not ( n247117 , n247114 );
and ( n247118 , n247116 , n247117 );
nor ( n247119 , n247115 , n247118 );
not ( n247120 , n247119 );
or ( n247121 , n247023 , n247120 );
not ( n247122 , n227002 );
and ( n247123 , n247058 , n247117 );
not ( n247124 , n247058 );
and ( n247125 , n247124 , n247114 );
nor ( n247126 , n247123 , n247125 );
nand ( n247127 , n247122 , n247126 );
nand ( n247128 , n247121 , n247127 );
not ( n247129 , n240292 );
not ( n247130 , n247129 );
not ( n247131 , n49603 );
not ( n247132 , n227360 );
nand ( n247133 , n247131 , n247132 );
not ( n247134 , n247133 );
or ( n247135 , n247130 , n247134 );
nand ( n247136 , n247131 , n247132 );
or ( n247137 , n247136 , n247129 );
nand ( n247138 , n247135 , n247137 );
not ( n247139 , n247138 );
nand ( n247140 , n49549 , n49573 );
and ( n247141 , n247140 , n240301 );
not ( n247142 , n247140 );
and ( n247143 , n247142 , n240162 );
nor ( n247144 , n247141 , n247143 );
not ( n247145 , n247144 );
and ( n247146 , n247139 , n247145 );
and ( n247147 , n247138 , n247144 );
nor ( n247148 , n247146 , n247147 );
not ( n247149 , n247148 );
not ( n247150 , n240265 );
nand ( n247151 , n49466 , n49493 );
not ( n247152 , n247151 );
or ( n247153 , n247150 , n247152 );
or ( n247154 , n247151 , n240265 );
nand ( n247155 , n247153 , n247154 );
not ( n247156 , n247155 );
not ( n247157 , n49432 );
nand ( n247158 , n49449 , n247157 );
not ( n247159 , n247158 );
not ( n247160 , n240207 );
and ( n247161 , n247159 , n247160 );
and ( n247162 , n247158 , n240207 );
nor ( n247163 , n247161 , n247162 );
not ( n247164 , n247163 );
or ( n247165 , n247156 , n247164 );
or ( n247166 , n247163 , n247155 );
nand ( n247167 , n247165 , n247166 );
not ( n247168 , n49506 );
nand ( n247169 , n247168 , n49527 );
not ( n247170 , n247169 );
not ( n247171 , n240239 );
and ( n247172 , n247170 , n247171 );
not ( n247173 , n49528 );
nand ( n247174 , n247173 , n247168 );
and ( n247175 , n247174 , n240239 );
nor ( n247176 , n247172 , n247175 );
not ( n247177 , n247176 );
and ( n247178 , n247167 , n247177 );
not ( n247179 , n247167 );
and ( n247180 , n247179 , n247176 );
nor ( n247181 , n247178 , n247180 );
not ( n247182 , n247181 );
or ( n247183 , n247149 , n247182 );
not ( n247184 , n247181 );
not ( n247185 , n247148 );
nand ( n247186 , n247184 , n247185 );
nand ( n247187 , n247183 , n247186 );
buf ( n247188 , n247187 );
and ( n247189 , n247128 , n247188 );
not ( n247190 , n247128 );
not ( n247191 , n247181 );
and ( n247192 , n247191 , n247185 );
not ( n247193 , n247191 );
and ( n247194 , n247193 , n247148 );
nor ( n247195 , n247192 , n247194 );
buf ( n247196 , n247195 );
and ( n247197 , n247190 , n247196 );
nor ( n247198 , n247189 , n247197 );
not ( n247199 , n247198 );
not ( n247200 , n247199 );
or ( n247201 , n247022 , n247200 );
not ( n247202 , n47950 );
not ( n247203 , n48676 );
or ( n247204 , n247202 , n247203 );
not ( n247205 , n47950 );
nand ( n247206 , n247205 , n48686 );
nand ( n247207 , n247204 , n247206 );
and ( n247208 , n247207 , n48797 );
not ( n247209 , n247207 );
and ( n247210 , n247209 , n48806 );
nor ( n247211 , n247208 , n247210 );
not ( n247212 , n226010 );
nor ( n247213 , n247211 , n247212 );
nand ( n247214 , n247201 , n247213 );
nor ( n247215 , n247198 , n33254 );
not ( n247216 , n247211 );
not ( n247217 , n247021 );
nor ( n247218 , n247216 , n247217 );
nand ( n247219 , n247215 , n247218 );
nand ( n247220 , n224937 , n31475 );
nand ( n247221 , n247214 , n247219 , n247220 );
buf ( n247222 , n247221 );
not ( n247223 , RI19aa62f8_2521);
or ( n247224 , n226819 , n247223 );
not ( n247225 , RI19a9ca28_2593);
or ( n247226 , n226822 , n247225 );
nand ( n247227 , n247224 , n247226 );
buf ( n247228 , n247227 );
buf ( n247229 , n233572 );
not ( n247230 , n247229 );
not ( n247231 , n49190 );
or ( n247232 , n247230 , n247231 );
or ( n247233 , n49190 , n247229 );
nand ( n247234 , n247232 , n247233 );
and ( n247235 , n247234 , n238186 );
not ( n247236 , n247234 );
and ( n247237 , n247236 , n238183 );
nor ( n247238 , n247235 , n247237 );
not ( n247239 , n247238 );
nand ( n247240 , n247239 , n222532 );
not ( n247241 , n227030 );
not ( n247242 , n247119 );
or ( n247243 , n247241 , n247242 );
not ( n247244 , n227030 );
nand ( n247245 , n247244 , n247126 );
nand ( n247246 , n247243 , n247245 );
and ( n247247 , n247246 , n247196 );
not ( n247248 , n247246 );
not ( n247249 , n247187 );
not ( n247250 , n247249 );
and ( n247251 , n247248 , n247250 );
nor ( n247252 , n247247 , n247251 );
not ( n247253 , n54616 );
not ( n247254 , n54627 );
nand ( n247255 , n247254 , n232785 );
not ( n247256 , n247255 );
or ( n247257 , n247253 , n247256 );
or ( n247258 , n247255 , n54616 );
nand ( n247259 , n247257 , n247258 );
not ( n247260 , n247259 );
not ( n247261 , n247260 );
not ( n247262 , n232514 );
or ( n247263 , n247261 , n247262 );
not ( n247264 , n247260 );
nand ( n247265 , n247264 , n232520 );
nand ( n247266 , n247263 , n247265 );
and ( n247267 , n247266 , n232299 );
not ( n247268 , n247266 );
buf ( n247269 , n246188 );
and ( n247270 , n247268 , n247269 );
nor ( n247271 , n247267 , n247270 );
not ( n247272 , n247271 );
nand ( n247273 , n247252 , n247272 );
or ( n247274 , n247240 , n247273 );
buf ( n247275 , n239934 );
not ( n247276 , n247275 );
nor ( n247277 , n247239 , n247276 );
nand ( n247278 , n247277 , n247273 );
nand ( n247279 , n39767 , n33508 );
nand ( n247280 , n247274 , n247278 , n247279 );
buf ( n247281 , n247280 );
not ( n247282 , n236438 );
nand ( n247283 , n32185 , n229015 );
not ( n247284 , n247283 );
or ( n247285 , n247282 , n247284 );
or ( n247286 , n236438 , n247283 );
nand ( n247287 , n247285 , n247286 );
not ( n247288 , n247287 );
not ( n247289 , n246548 );
or ( n247290 , n247288 , n247289 );
not ( n247291 , n247287 );
nand ( n247292 , n247291 , n246553 );
nand ( n247293 , n247290 , n247292 );
and ( n247294 , n247293 , n246661 );
not ( n247295 , n247293 );
and ( n247296 , n247295 , n246654 );
nor ( n247297 , n247294 , n247296 );
not ( n247298 , n55125 );
nand ( n247299 , n240782 , n37111 );
not ( n247300 , n247299 );
or ( n247301 , n247298 , n247300 );
or ( n247302 , n247299 , n55125 );
nand ( n247303 , n247301 , n247302 );
not ( n247304 , n247303 );
nand ( n247305 , n240762 , n37232 );
not ( n247306 , n247305 );
not ( n247307 , n245579 );
and ( n247308 , n247306 , n247307 );
not ( n247309 , n37231 );
nand ( n247310 , n247309 , n240762 );
and ( n247311 , n247310 , n245579 );
nor ( n247312 , n247308 , n247311 );
not ( n247313 , n247312 );
or ( n247314 , n247304 , n247313 );
or ( n247315 , n247312 , n247303 );
nand ( n247316 , n247314 , n247315 );
nand ( n247317 , n240714 , n37274 );
not ( n247318 , n247317 );
not ( n247319 , n36761 );
and ( n247320 , n247318 , n247319 );
and ( n247321 , n247317 , n36761 );
nor ( n247322 , n247320 , n247321 );
and ( n247323 , n247316 , n247322 );
not ( n247324 , n247316 );
not ( n247325 , n247322 );
and ( n247326 , n247324 , n247325 );
nor ( n247327 , n247323 , n247326 );
nand ( n247328 , n36895 , n240740 );
and ( n247329 , n247328 , n245566 );
not ( n247330 , n247328 );
and ( n247331 , n247330 , n246125 );
nor ( n247332 , n247329 , n247331 );
not ( n247333 , n247332 );
nand ( n247334 , n246119 , n37028 );
not ( n247335 , n247334 );
not ( n247336 , n245550 );
or ( n247337 , n247335 , n247336 );
or ( n247338 , n245550 , n247334 );
nand ( n247339 , n247337 , n247338 );
not ( n247340 , n247339 );
and ( n247341 , n247333 , n247340 );
and ( n247342 , n247332 , n247339 );
nor ( n247343 , n247341 , n247342 );
not ( n247344 , n247343 );
and ( n247345 , n247327 , n247344 );
not ( n247346 , n247327 );
and ( n247347 , n247346 , n247343 );
nor ( n247348 , n247345 , n247347 );
buf ( n247349 , n247348 );
not ( n247350 , n247349 );
not ( n247351 , n240573 );
not ( n247352 , n240370 );
not ( n247353 , n247352 );
not ( n247354 , n240568 );
nand ( n247355 , n247354 , n240379 );
not ( n247356 , n247355 );
and ( n247357 , n247353 , n247356 );
and ( n247358 , n247352 , n247355 );
nor ( n247359 , n247357 , n247358 );
not ( n247360 , n247359 );
nand ( n247361 , n240588 , n240585 );
and ( n247362 , n247361 , n240353 );
not ( n247363 , n247361 );
and ( n247364 , n247363 , n240352 );
nor ( n247365 , n247362 , n247364 );
not ( n247366 , n247365 );
or ( n247367 , n247360 , n247366 );
or ( n247368 , n247365 , n247359 );
nand ( n247369 , n247367 , n247368 );
nand ( n247370 , n240619 , n240602 );
and ( n247371 , n247370 , n240410 );
not ( n247372 , n247370 );
and ( n247373 , n247372 , n240409 );
nor ( n247374 , n247371 , n247373 );
not ( n247375 , n247374 );
and ( n247376 , n247369 , n247375 );
not ( n247377 , n247369 );
and ( n247378 , n247377 , n247374 );
nor ( n247379 , n247376 , n247378 );
not ( n247380 , n240465 );
nand ( n247381 , n247380 , n240548 );
and ( n247382 , n247381 , n240456 );
not ( n247383 , n247381 );
and ( n247384 , n247383 , n240455 );
nor ( n247385 , n247382 , n247384 );
not ( n247386 , n247385 );
not ( n247387 , n247386 );
not ( n247388 , n246107 );
or ( n247389 , n247387 , n247388 );
not ( n247390 , n246107 );
nand ( n247391 , n247390 , n247385 );
nand ( n247392 , n247389 , n247391 );
xor ( n247393 , n247379 , n247392 );
not ( n247394 , n247393 );
or ( n247395 , n247351 , n247394 );
not ( n247396 , n240573 );
or ( n247397 , n247379 , n247392 );
nand ( n247398 , n247379 , n247392 );
nand ( n247399 , n247397 , n247398 );
nand ( n247400 , n247396 , n247399 );
nand ( n247401 , n247395 , n247400 );
not ( n247402 , n247401 );
or ( n247403 , n247350 , n247402 );
or ( n247404 , n247401 , n247349 );
nand ( n247405 , n247403 , n247404 );
not ( n247406 , n247405 );
nand ( n247407 , n247297 , n247406 );
and ( n247408 , n244695 , n241723 );
not ( n247409 , n244695 );
and ( n247410 , n247409 , n241715 );
or ( n247411 , n247408 , n247410 );
and ( n247412 , n247411 , n241878 );
not ( n247413 , n247411 );
and ( n247414 , n247413 , n241885 );
nor ( n247415 , n247412 , n247414 );
nand ( n247416 , n247415 , n33255 );
or ( n247417 , n247407 , n247416 );
not ( n247418 , n247415 );
not ( n247419 , n247297 );
or ( n247420 , n247418 , n247419 );
nor ( n247421 , n247406 , n47173 );
nand ( n247422 , n247420 , n247421 );
buf ( n247423 , n35431 );
nand ( n247424 , n247423 , n42500 );
nand ( n247425 , n247417 , n247422 , n247424 );
buf ( n247426 , n247425 );
not ( n247427 , n50653 );
not ( n247428 , n46780 );
nand ( n247429 , n247428 , n46791 );
not ( n247430 , n247429 );
or ( n247431 , n247427 , n247430 );
or ( n247432 , n247429 , n50653 );
nand ( n247433 , n247431 , n247432 );
not ( n247434 , n247433 );
not ( n247435 , n228527 );
or ( n247436 , n247434 , n247435 );
not ( n247437 , n247433 );
nand ( n247438 , n247437 , n50776 );
nand ( n247439 , n247436 , n247438 );
and ( n247440 , n247439 , n50931 );
not ( n247441 , n247439 );
and ( n247442 , n247441 , n50941 );
nor ( n247443 , n247440 , n247442 );
not ( n247444 , n33253 );
nand ( n247445 , n247443 , n247444 );
not ( n247446 , n247445 );
not ( n247447 , n238813 );
nand ( n247448 , n43373 , n238811 );
buf ( n247449 , n236576 );
xor ( n247450 , n247448 , n247449 );
not ( n247451 , n247450 );
not ( n247452 , n247451 );
nand ( n247453 , n238828 , n221154 );
and ( n247454 , n247453 , n243477 );
not ( n247455 , n247453 );
and ( n247456 , n247455 , n43266 );
nor ( n247457 , n247454 , n247456 );
not ( n247458 , n247457 );
not ( n247459 , n247458 );
or ( n247460 , n247452 , n247459 );
nand ( n247461 , n247457 , n247450 );
nand ( n247462 , n247460 , n247461 );
not ( n247463 , n247462 );
nand ( n247464 , n43479 , n236560 );
and ( n247465 , n247464 , n236553 );
not ( n247466 , n247464 );
and ( n247467 , n247466 , n236618 );
nor ( n247468 , n247465 , n247467 );
not ( n247469 , n247468 );
not ( n247470 , n247469 );
nor ( n247471 , n238850 , n43328 );
not ( n247472 , n247471 );
not ( n247473 , n236601 );
and ( n247474 , n247472 , n247473 );
and ( n247475 , n247471 , n236601 );
nor ( n247476 , n247474 , n247475 );
not ( n247477 , n247476 );
not ( n247478 , n247477 );
or ( n247479 , n247470 , n247478 );
nand ( n247480 , n247476 , n247468 );
nand ( n247481 , n247479 , n247480 );
nand ( n247482 , n238878 , n43440 );
not ( n247483 , n247482 );
not ( n247484 , n56059 );
and ( n247485 , n247483 , n247484 );
not ( n247486 , n241186 );
and ( n247487 , n247482 , n247486 );
nor ( n247488 , n247485 , n247487 );
and ( n247489 , n247481 , n247488 );
not ( n247490 , n247481 );
not ( n247491 , n247488 );
and ( n247492 , n247490 , n247491 );
nor ( n247493 , n247489 , n247492 );
not ( n247494 , n247493 );
or ( n247495 , n247463 , n247494 );
not ( n247496 , n247493 );
not ( n247497 , n247462 );
nand ( n247498 , n247496 , n247497 );
nand ( n247499 , n247495 , n247498 );
not ( n247500 , n247499 );
not ( n247501 , n247500 );
or ( n247502 , n247447 , n247501 );
not ( n247503 , n238813 );
nand ( n247504 , n247503 , n247499 );
nand ( n247505 , n247502 , n247504 );
nand ( n247506 , n243723 , n43024 );
not ( n247507 , n247506 );
not ( n247508 , n236659 );
and ( n247509 , n247507 , n247508 );
and ( n247510 , n247506 , n236659 );
nor ( n247511 , n247509 , n247510 );
not ( n247512 , n247511 );
not ( n247513 , n243743 );
nand ( n247514 , n247513 , n43098 );
not ( n247515 , n236680 );
and ( n247516 , n247514 , n247515 );
not ( n247517 , n247514 );
and ( n247518 , n247517 , n236680 );
nor ( n247519 , n247516 , n247518 );
not ( n247520 , n247519 );
or ( n247521 , n247512 , n247520 );
or ( n247522 , n247519 , n247511 );
nand ( n247523 , n247521 , n247522 );
nand ( n247524 , n243763 , n43139 );
and ( n247525 , n247524 , n243765 );
not ( n247526 , n247524 );
and ( n247527 , n247526 , n236701 );
nor ( n247528 , n247525 , n247527 );
and ( n247529 , n247523 , n247528 );
not ( n247530 , n247523 );
not ( n247531 , n247528 );
and ( n247532 , n247530 , n247531 );
nor ( n247533 , n247529 , n247532 );
not ( n247534 , n247533 );
not ( n247535 , n247534 );
nand ( n247536 , n243786 , n43175 );
not ( n247537 , n247536 );
not ( n247538 , n236726 );
and ( n247539 , n247537 , n247538 );
nand ( n247540 , n243786 , n43175 );
and ( n247541 , n247540 , n236726 );
nor ( n247542 , n247539 , n247541 );
not ( n247543 , n247542 );
not ( n247544 , n243713 );
nand ( n247545 , n247543 , n247544 );
nand ( n247546 , n247542 , n243713 );
nand ( n247547 , n247545 , n247546 );
not ( n247548 , n247547 );
and ( n247549 , n247535 , n247548 );
and ( n247550 , n247534 , n247547 );
nor ( n247551 , n247549 , n247550 );
not ( n247552 , n247551 );
not ( n247553 , n247552 );
and ( n247554 , n247505 , n247553 );
not ( n247555 , n247505 );
not ( n247556 , n247533 );
not ( n247557 , n247547 );
not ( n247558 , n247557 );
or ( n247559 , n247556 , n247558 );
nand ( n247560 , n247534 , n247547 );
nand ( n247561 , n247559 , n247560 );
not ( n247562 , n247561 );
not ( n247563 , n247562 );
and ( n247564 , n247555 , n247563 );
nor ( n247565 , n247554 , n247564 );
not ( n247566 , n247565 );
not ( n247567 , n247566 );
not ( n247568 , n239870 );
not ( n247569 , n230199 );
not ( n247570 , n247569 );
or ( n247571 , n247568 , n247570 );
not ( n247572 , n230199 );
or ( n247573 , n247572 , n239870 );
nand ( n247574 , n247571 , n247573 );
buf ( n247575 , n236637 );
and ( n247576 , n247574 , n247575 );
not ( n247577 , n247574 );
and ( n247578 , n247577 , n242696 );
nor ( n247579 , n247576 , n247578 );
nand ( n247580 , n247567 , n247579 );
nand ( n247581 , n247446 , n247580 );
nor ( n247582 , n247566 , n33254 );
not ( n247583 , n247443 );
nand ( n247584 , n247582 , n247579 , n247583 );
buf ( n247585 , n35431 );
nand ( n247586 , n247585 , n41006 );
nand ( n247587 , n247581 , n247584 , n247586 );
buf ( n247588 , n247587 );
nand ( n247589 , n239151 , n48076 );
not ( n247590 , n247589 );
not ( n247591 , n226512 );
and ( n247592 , n247590 , n247591 );
and ( n247593 , n247589 , n226512 );
nor ( n247594 , n247592 , n247593 );
not ( n247595 , n247594 );
not ( n247596 , n225796 );
nor ( n247597 , n48049 , n239194 );
not ( n247598 , n247597 );
or ( n247599 , n247596 , n247598 );
or ( n247600 , n247597 , n225796 );
nand ( n247601 , n247599 , n247600 );
not ( n247602 , n247601 );
or ( n247603 , n247595 , n247602 );
or ( n247604 , n247594 , n247601 );
nand ( n247605 , n247603 , n247604 );
nand ( n247606 , n240105 , n239134 );
buf ( n247607 , n48137 );
and ( n247608 , n247606 , n247607 );
not ( n247609 , n247606 );
not ( n247610 , n247607 );
and ( n247611 , n247609 , n247610 );
nor ( n247612 , n247608 , n247611 );
not ( n247613 , n247612 );
and ( n247614 , n247605 , n247613 );
not ( n247615 , n247605 );
and ( n247616 , n247615 , n247612 );
nor ( n247617 , n247614 , n247616 );
not ( n247618 , n247617 );
not ( n247619 , n247618 );
nand ( n247620 , n239210 , n48217 );
not ( n247621 , n48207 );
and ( n247622 , n247620 , n247621 );
not ( n247623 , n247620 );
and ( n247624 , n247623 , n48207 );
nor ( n247625 , n247622 , n247624 );
not ( n247626 , n247625 );
not ( n247627 , n247626 );
not ( n247628 , n48184 );
nand ( n247629 , n239173 , n247628 );
not ( n247630 , n247629 );
not ( n247631 , n48689 );
and ( n247632 , n247630 , n247631 );
and ( n247633 , n247629 , n48689 );
nor ( n247634 , n247632 , n247633 );
not ( n247635 , n247634 );
not ( n247636 , n247635 );
or ( n247637 , n247627 , n247636 );
nand ( n247638 , n247634 , n247625 );
nand ( n247639 , n247637 , n247638 );
not ( n247640 , n247639 );
not ( n247641 , n247640 );
or ( n247642 , n247619 , n247641 );
nand ( n247643 , n247617 , n247639 );
nand ( n247644 , n247642 , n247643 );
buf ( n247645 , n247644 );
not ( n247646 , n247645 );
not ( n247647 , n247646 );
not ( n247648 , n55092 );
not ( n247649 , n47841 );
nand ( n247650 , n247649 , n234381 );
and ( n247651 , n247650 , n225581 );
not ( n247652 , n247650 );
and ( n247653 , n247652 , n226328 );
nor ( n247654 , n247651 , n247653 );
not ( n247655 , n247654 );
or ( n247656 , n247648 , n247655 );
or ( n247657 , n55092 , n247654 );
nand ( n247658 , n247656 , n247657 );
nand ( n247659 , n225674 , n234397 );
not ( n247660 , n247659 );
not ( n247661 , n48633 );
and ( n247662 , n247660 , n247661 );
and ( n247663 , n247659 , n48633 );
nor ( n247664 , n247662 , n247663 );
and ( n247665 , n247658 , n247664 );
not ( n247666 , n247658 );
not ( n247667 , n247664 );
and ( n247668 , n247666 , n247667 );
nor ( n247669 , n247665 , n247668 );
not ( n247670 , n247669 );
not ( n247671 , n247670 );
not ( n247672 , n47968 );
nand ( n247673 , n247672 , n234357 );
not ( n247674 , n247673 );
not ( n247675 , n48607 );
or ( n247676 , n247674 , n247675 );
or ( n247677 , n48607 , n247673 );
nand ( n247678 , n247676 , n247677 );
not ( n247679 , n247678 );
not ( n247680 , n47807 );
or ( n247681 , n247679 , n247680 );
not ( n247682 , n247678 );
nand ( n247683 , n247682 , n47806 );
nand ( n247684 , n247681 , n247683 );
not ( n247685 , n247684 );
not ( n247686 , n247685 );
or ( n247687 , n247671 , n247686 );
nand ( n247688 , n247684 , n247669 );
nand ( n247689 , n247687 , n247688 );
and ( n247690 , n247689 , n238048 );
not ( n247691 , n247689 );
and ( n247692 , n247691 , n238047 );
or ( n247693 , n247690 , n247692 );
not ( n247694 , n247693 );
or ( n247695 , n247647 , n247694 );
or ( n247696 , n247693 , n247646 );
nand ( n247697 , n247695 , n247696 );
buf ( n247698 , n31571 );
nor ( n247699 , n247697 , n247698 );
not ( n247700 , n226284 );
nand ( n247701 , n247700 , n237977 );
not ( n247702 , n247701 );
not ( n247703 , n225423 );
and ( n247704 , n247702 , n247703 );
and ( n247705 , n247701 , n225423 );
nor ( n247706 , n247704 , n247705 );
not ( n247707 , n247706 );
not ( n247708 , n236781 );
or ( n247709 , n247707 , n247708 );
or ( n247710 , n236781 , n247706 );
nand ( n247711 , n247709 , n247710 );
and ( n247712 , n247711 , n236789 );
not ( n247713 , n247711 );
and ( n247714 , n247713 , n234889 );
nor ( n247715 , n247712 , n247714 );
not ( n247716 , n247715 );
not ( n247717 , n238173 );
not ( n247718 , n247717 );
not ( n247719 , n45727 );
or ( n247720 , n247718 , n247719 );
not ( n247721 , n247717 );
not ( n247722 , n45722 );
not ( n247723 , n223407 );
or ( n247724 , n247722 , n247723 );
not ( n247725 , n223407 );
nand ( n247726 , n247725 , n223486 );
nand ( n247727 , n247724 , n247726 );
nand ( n247728 , n247721 , n247727 );
nand ( n247729 , n247720 , n247728 );
buf ( n247730 , n245743 );
and ( n247731 , n247729 , n247730 );
not ( n247732 , n247729 );
buf ( n247733 , n245738 );
and ( n247734 , n247732 , n247733 );
nor ( n247735 , n247731 , n247734 );
not ( n247736 , n247735 );
nand ( n247737 , n247699 , n247716 , n247736 );
not ( n247738 , n247697 );
not ( n247739 , n247738 );
not ( n247740 , n247716 );
or ( n247741 , n247739 , n247740 );
nor ( n247742 , n247736 , n31572 );
nand ( n247743 , n247741 , n247742 );
buf ( n247744 , n35431 );
nand ( n247745 , n247744 , n223314 );
nand ( n247746 , n247737 , n247743 , n247745 );
buf ( n247747 , n247746 );
buf ( n247748 , n40883 );
buf ( n247749 , n205902 );
not ( n247750 , n29053 );
not ( n247751 , n31577 );
or ( n247752 , n247750 , n247751 );
not ( n247753 , n239700 );
not ( n247754 , n238975 );
or ( n247755 , n247753 , n247754 );
not ( n247756 , n239700 );
nand ( n247757 , n247756 , n238985 );
nand ( n247758 , n247755 , n247757 );
and ( n247759 , n247758 , n239108 );
not ( n247760 , n247758 );
and ( n247761 , n247760 , n239100 );
nor ( n247762 , n247759 , n247761 );
not ( n247763 , n247762 );
not ( n247764 , n40187 );
not ( n247765 , n235807 );
or ( n247766 , n247764 , n247765 );
not ( n247767 , n40187 );
nand ( n247768 , n247767 , n235815 );
nand ( n247769 , n247766 , n247768 );
and ( n247770 , n247769 , n235879 );
not ( n247771 , n247769 );
and ( n247772 , n247771 , n235888 );
nor ( n247773 , n247770 , n247772 );
nand ( n247774 , n247763 , n247773 );
not ( n247775 , n237426 );
nand ( n247776 , n54956 , n54711 );
not ( n247777 , n247776 );
not ( n247778 , n245501 );
and ( n247779 , n247777 , n247778 );
and ( n247780 , n247776 , n245501 );
nor ( n247781 , n247779 , n247780 );
not ( n247782 , n247781 );
not ( n247783 , n232338 );
or ( n247784 , n247782 , n247783 );
or ( n247785 , n232338 , n247781 );
nand ( n247786 , n247784 , n247785 );
not ( n247787 , n237410 );
nand ( n247788 , n247787 , n54991 );
xor ( n247789 , n247788 , n54664 );
and ( n247790 , n247786 , n247789 );
not ( n247791 , n247786 );
not ( n247792 , n247789 );
and ( n247793 , n247791 , n247792 );
nor ( n247794 , n247790 , n247793 );
not ( n247795 , n247794 );
not ( n247796 , n247795 );
nand ( n247797 , n232367 , n232815 );
not ( n247798 , n247797 );
not ( n247799 , n54597 );
not ( n247800 , n247799 );
and ( n247801 , n247798 , n247800 );
and ( n247802 , n247797 , n247799 );
nor ( n247803 , n247801 , n247802 );
not ( n247804 , n247803 );
not ( n247805 , n247804 );
not ( n247806 , n247260 );
or ( n247807 , n247805 , n247806 );
nand ( n247808 , n247803 , n247259 );
nand ( n247809 , n247807 , n247808 );
not ( n247810 , n247809 );
and ( n247811 , n247796 , n247810 );
and ( n247812 , n247795 , n247809 );
nor ( n247813 , n247811 , n247812 );
not ( n247814 , n247813 );
or ( n247815 , n247775 , n247814 );
not ( n247816 , n237426 );
not ( n247817 , n247809 );
not ( n247818 , n247817 );
not ( n247819 , n247794 );
or ( n247820 , n247818 , n247819 );
nand ( n247821 , n247795 , n247809 );
nand ( n247822 , n247820 , n247821 );
nand ( n247823 , n247816 , n247822 );
nand ( n247824 , n247815 , n247823 );
not ( n247825 , n232111 );
nand ( n247826 , n237462 , n232122 );
not ( n247827 , n247826 );
or ( n247828 , n247825 , n247827 );
or ( n247829 , n247826 , n232111 );
nand ( n247830 , n247828 , n247829 );
not ( n247831 , n247830 );
nand ( n247832 , n241912 , n232152 );
not ( n247833 , n247832 );
not ( n247834 , n54405 );
not ( n247835 , n247834 );
and ( n247836 , n247833 , n247835 );
nand ( n247837 , n232152 , n241912 );
and ( n247838 , n247837 , n247834 );
nor ( n247839 , n247836 , n247838 );
not ( n247840 , n247839 );
or ( n247841 , n247831 , n247840 );
or ( n247842 , n247839 , n247830 );
nand ( n247843 , n247841 , n247842 );
and ( n247844 , n247843 , n246185 );
not ( n247845 , n247843 );
and ( n247846 , n247845 , n246184 );
nor ( n247847 , n247844 , n247846 );
nand ( n247848 , n237533 , n237550 );
not ( n247849 , n247848 );
not ( n247850 , n245456 );
and ( n247851 , n247849 , n247850 );
and ( n247852 , n247848 , n245456 );
nor ( n247853 , n247851 , n247852 );
not ( n247854 , n247853 );
not ( n247855 , n232261 );
nand ( n247856 , n247855 , n237574 );
not ( n247857 , n245448 );
and ( n247858 , n247856 , n247857 );
not ( n247859 , n247856 );
and ( n247860 , n247859 , n245448 );
nor ( n247861 , n247858 , n247860 );
not ( n247862 , n247861 );
or ( n247863 , n247854 , n247862 );
or ( n247864 , n247861 , n247853 );
nand ( n247865 , n247863 , n247864 );
and ( n247866 , n247847 , n247865 );
not ( n247867 , n247847 );
not ( n247868 , n247865 );
and ( n247869 , n247867 , n247868 );
nor ( n247870 , n247866 , n247869 );
buf ( n247871 , n247870 );
buf ( n247872 , n247871 );
not ( n247873 , n247872 );
and ( n247874 , n247824 , n247873 );
not ( n247875 , n247824 );
and ( n247876 , n247875 , n247872 );
nor ( n247877 , n247874 , n247876 );
and ( n247878 , n247774 , n247877 );
not ( n247879 , n247774 );
not ( n247880 , n247877 );
and ( n247881 , n247879 , n247880 );
nor ( n247882 , n247878 , n247881 );
or ( n247883 , n247882 , n237358 );
nand ( n247884 , n247752 , n247883 );
buf ( n247885 , n247884 );
not ( n247886 , n29503 );
not ( n247887 , n245943 );
or ( n247888 , n247886 , n247887 );
not ( n247889 , n223817 );
nand ( n247890 , n45888 , n45913 );
not ( n247891 , n247890 );
not ( n247892 , n46542 );
and ( n247893 , n247891 , n247892 );
and ( n247894 , n247890 , n46542 );
nor ( n247895 , n247893 , n247894 );
not ( n247896 , n247895 );
not ( n247897 , n45984 );
nand ( n247898 , n247897 , n45973 );
and ( n247899 , n247898 , n46607 );
not ( n247900 , n247898 );
and ( n247901 , n247900 , n224369 );
nor ( n247902 , n247899 , n247901 );
not ( n247903 , n247902 );
or ( n247904 , n247896 , n247903 );
or ( n247905 , n247902 , n247895 );
nand ( n247906 , n247904 , n247905 );
not ( n247907 , n45952 );
nand ( n247908 , n247907 , n244496 );
and ( n247909 , n247908 , n46630 );
not ( n247910 , n247908 );
and ( n247911 , n247910 , n46631 );
nor ( n247912 , n247909 , n247911 );
not ( n247913 , n247912 );
and ( n247914 , n247906 , n247913 );
not ( n247915 , n247906 );
and ( n247916 , n247915 , n247912 );
nor ( n247917 , n247914 , n247916 );
not ( n247918 , n46659 );
nand ( n247919 , n46022 , n46010 );
not ( n247920 , n247919 );
and ( n247921 , n247918 , n247920 );
and ( n247922 , n46659 , n247919 );
nor ( n247923 , n247921 , n247922 );
not ( n247924 , n247923 );
not ( n247925 , n247924 );
not ( n247926 , n239804 );
not ( n247927 , n247926 );
or ( n247928 , n247925 , n247927 );
nand ( n247929 , n239804 , n247923 );
nand ( n247930 , n247928 , n247929 );
xor ( n247931 , n247917 , n247930 );
not ( n247932 , n247931 );
or ( n247933 , n247889 , n247932 );
not ( n247934 , n247931 );
nand ( n247935 , n247934 , n46060 );
nand ( n247936 , n247933 , n247935 );
not ( n247937 , n230064 );
not ( n247938 , n238779 );
not ( n247939 , n238766 );
not ( n247940 , n247939 );
nand ( n247941 , n247938 , n247940 );
not ( n247942 , n247941 );
or ( n247943 , n247937 , n247942 );
or ( n247944 , n247941 , n230064 );
nand ( n247945 , n247943 , n247944 );
not ( n247946 , n247945 );
not ( n247947 , n247946 );
not ( n247948 , n238747 );
nand ( n247949 , n247948 , n238794 );
not ( n247950 , n247949 );
buf ( n247951 , n52262 );
not ( n247952 , n247951 );
and ( n247953 , n247950 , n247952 );
nand ( n247954 , n247948 , n238794 );
and ( n247955 , n247954 , n247951 );
nor ( n247956 , n247953 , n247955 );
not ( n247957 , n247956 );
not ( n247958 , n247957 );
or ( n247959 , n247947 , n247958 );
nand ( n247960 , n247956 , n247945 );
nand ( n247961 , n247959 , n247960 );
nand ( n247962 , n238665 , n238652 );
not ( n247963 , n247962 );
not ( n247964 , n52378 );
not ( n247965 , n247964 );
not ( n247966 , n247965 );
and ( n247967 , n247963 , n247966 );
and ( n247968 , n247962 , n247965 );
nor ( n247969 , n247967 , n247968 );
not ( n247970 , n247969 );
not ( n247971 , n243461 );
or ( n247972 , n247970 , n247971 );
or ( n247973 , n243461 , n247969 );
nand ( n247974 , n247972 , n247973 );
not ( n247975 , n238677 );
nand ( n247976 , n238687 , n247975 );
not ( n247977 , n247976 );
not ( n247978 , n52397 );
or ( n247979 , n247977 , n247978 );
or ( n247980 , n52397 , n247976 );
nand ( n247981 , n247979 , n247980 );
not ( n247982 , n247981 );
and ( n247983 , n247974 , n247982 );
not ( n247984 , n247974 );
and ( n247985 , n247984 , n247981 );
nor ( n247986 , n247983 , n247985 );
not ( n247987 , n247986 );
and ( n247988 , n247961 , n247987 );
not ( n247989 , n247961 );
and ( n247990 , n247989 , n247986 );
or ( n247991 , n247988 , n247990 );
and ( n247992 , n247936 , n247991 );
not ( n247993 , n247936 );
not ( n247994 , n247961 );
not ( n247995 , n247994 );
not ( n247996 , n247987 );
or ( n247997 , n247995 , n247996 );
nand ( n247998 , n247986 , n247961 );
nand ( n247999 , n247997 , n247998 );
buf ( n248000 , n247999 );
and ( n248001 , n247993 , n248000 );
nor ( n248002 , n247992 , n248001 );
not ( n248003 , n248002 );
buf ( n248004 , n230152 );
not ( n248005 , n248004 );
not ( n248006 , n238795 );
not ( n248007 , n52421 );
nand ( n248008 , n248007 , n230167 );
and ( n248009 , n248008 , n238677 );
not ( n248010 , n248008 );
and ( n248011 , n248010 , n247975 );
nor ( n248012 , n248009 , n248011 );
not ( n248013 , n248012 );
or ( n248014 , n248006 , n248013 );
or ( n248015 , n238795 , n248012 );
nand ( n248016 , n248014 , n248015 );
not ( n248017 , n248016 );
not ( n248018 , n52307 );
nand ( n248019 , n248018 , n239875 );
not ( n248020 , n248019 );
not ( n248021 , n247940 );
and ( n248022 , n248020 , n248021 );
not ( n248023 , n52294 );
nand ( n248024 , n248023 , n248018 );
and ( n248025 , n248024 , n247940 );
nor ( n248026 , n248022 , n248025 );
not ( n248027 , n248026 );
and ( n248028 , n248017 , n248027 );
and ( n248029 , n248016 , n248026 );
nor ( n248030 , n248028 , n248029 );
not ( n248031 , n52356 );
nand ( n248032 , n248031 , n239898 );
not ( n248033 , n248032 );
not ( n248034 , n238707 );
and ( n248035 , n248033 , n248034 );
and ( n248036 , n248032 , n238707 );
nor ( n248037 , n248035 , n248036 );
not ( n248038 , n248037 );
buf ( n248039 , n238652 );
not ( n248040 , n248039 );
nand ( n248041 , n239886 , n52390 );
not ( n248042 , n248041 );
or ( n248043 , n248040 , n248042 );
or ( n248044 , n248041 , n248039 );
nand ( n248045 , n248043 , n248044 );
not ( n248046 , n248045 );
or ( n248047 , n248038 , n248046 );
or ( n248048 , n248045 , n248037 );
nand ( n248049 , n248047 , n248048 );
and ( n248050 , n248030 , n248049 );
not ( n248051 , n248030 );
not ( n248052 , n248049 );
and ( n248053 , n248051 , n248052 );
nor ( n248054 , n248050 , n248053 );
not ( n248055 , n248054 );
not ( n248056 , n248055 );
not ( n248057 , n248056 );
or ( n248058 , n248005 , n248057 );
not ( n248059 , n248004 );
nand ( n248060 , n248059 , n248055 );
nand ( n248061 , n248058 , n248060 );
not ( n248062 , n43496 );
buf ( n248063 , n248062 );
and ( n248064 , n248061 , n248063 );
not ( n248065 , n248061 );
not ( n248066 , n43497 );
buf ( n248067 , n248066 );
and ( n248068 , n248065 , n248067 );
nor ( n248069 , n248064 , n248068 );
nand ( n248070 , n248003 , n248069 );
not ( n248071 , n245383 );
not ( n248072 , n235357 );
or ( n248073 , n248071 , n248072 );
not ( n248074 , n245383 );
nand ( n248075 , n248074 , n235366 );
nand ( n248076 , n248073 , n248075 );
and ( n248077 , n248076 , n235372 );
not ( n248078 , n248076 );
and ( n248079 , n248078 , n235369 );
nor ( n248080 , n248077 , n248079 );
and ( n248081 , n248070 , n248080 );
not ( n248082 , n248070 );
not ( n248083 , n248080 );
and ( n248084 , n248082 , n248083 );
nor ( n248085 , n248081 , n248084 );
or ( n248086 , n248085 , n244217 );
nand ( n248087 , n247888 , n248086 );
buf ( n248088 , n248087 );
not ( n248089 , n34010 );
not ( n248090 , n50615 );
or ( n248091 , n248089 , n248090 );
not ( n248092 , n235439 );
nand ( n248093 , n235433 , n235411 );
not ( n248094 , n248093 );
not ( n248095 , n238519 );
and ( n248096 , n248094 , n248095 );
nand ( n248097 , n235433 , n235411 );
and ( n248098 , n248097 , n238519 );
nor ( n248099 , n248096 , n248098 );
nand ( n248100 , n241076 , n235464 );
buf ( n248101 , n238536 );
xor ( n248102 , n248100 , n248101 );
xor ( n248103 , n248099 , n248102 );
not ( n248104 , n238500 );
not ( n248105 , n248104 );
nor ( n248106 , n235494 , n235486 );
not ( n248107 , n248106 );
and ( n248108 , n248105 , n248107 );
and ( n248109 , n248104 , n248106 );
nor ( n248110 , n248108 , n248109 );
xnor ( n248111 , n248103 , n248110 );
not ( n248112 , n238582 );
nand ( n248113 , n235555 , n235567 );
not ( n248114 , n248113 );
or ( n248115 , n248112 , n248114 );
or ( n248116 , n248113 , n238582 );
nand ( n248117 , n248115 , n248116 );
not ( n248118 , n248117 );
not ( n248119 , n235514 );
nand ( n248120 , n248119 , n235517 );
and ( n248121 , n248120 , n238602 );
not ( n248122 , n248120 );
and ( n248123 , n248122 , n238603 );
nor ( n248124 , n248121 , n248123 );
not ( n248125 , n248124 );
not ( n248126 , n248125 );
or ( n248127 , n248118 , n248126 );
not ( n248128 , n248117 );
nand ( n248129 , n248128 , n248124 );
nand ( n248130 , n248127 , n248129 );
and ( n248131 , n248111 , n248130 );
not ( n248132 , n248111 );
not ( n248133 , n248130 );
and ( n248134 , n248132 , n248133 );
nor ( n248135 , n248131 , n248134 );
not ( n248136 , n248135 );
or ( n248137 , n248092 , n248136 );
not ( n248138 , n235439 );
not ( n248139 , n248111 );
and ( n248140 , n248139 , n248130 );
not ( n248141 , n248139 );
and ( n248142 , n248141 , n248133 );
nor ( n248143 , n248140 , n248142 );
nand ( n248144 , n248138 , n248143 );
nand ( n248145 , n248137 , n248144 );
buf ( n248146 , n238461 );
and ( n248147 , n248145 , n248146 );
not ( n248148 , n248145 );
buf ( n248149 , n238470 );
and ( n248150 , n248148 , n248149 );
nor ( n248151 , n248147 , n248150 );
not ( n248152 , n248151 );
not ( n248153 , n45498 );
not ( n248154 , n234184 );
not ( n248155 , n248154 );
or ( n248156 , n248153 , n248155 );
not ( n248157 , n45498 );
and ( n248158 , n234149 , n234179 );
not ( n248159 , n234149 );
and ( n248160 , n248159 , n234182 );
nor ( n248161 , n248158 , n248160 );
nand ( n248162 , n248157 , n248161 );
nand ( n248163 , n248156 , n248162 );
nand ( n248164 , n45710 , n45688 );
not ( n248165 , n248164 );
not ( n248166 , n239948 );
not ( n248167 , n248166 );
or ( n248168 , n248165 , n248167 );
or ( n248169 , n248166 , n248164 );
nand ( n248170 , n248168 , n248169 );
not ( n248171 , n248170 );
not ( n248172 , n248171 );
not ( n248173 , n55992 );
nand ( n248174 , n45673 , n45666 );
not ( n248175 , n248174 );
or ( n248176 , n248173 , n248175 );
or ( n248177 , n248174 , n55992 );
nand ( n248178 , n248176 , n248177 );
not ( n248179 , n248178 );
or ( n248180 , n248172 , n248179 );
not ( n248181 , n248178 );
nand ( n248182 , n248181 , n248170 );
nand ( n248183 , n248180 , n248182 );
not ( n248184 , n45545 );
nand ( n248185 , n248184 , n238157 );
not ( n248186 , n248185 );
not ( n248187 , n55953 );
and ( n248188 , n248186 , n248187 );
and ( n248189 , n248185 , n55953 );
nor ( n248190 , n248188 , n248189 );
not ( n248191 , n248190 );
nand ( n248192 , n238169 , n45590 );
and ( n248193 , n248192 , n239967 );
not ( n248194 , n248192 );
and ( n248195 , n248194 , n233686 );
nor ( n248196 , n248193 , n248195 );
not ( n248197 , n248196 );
or ( n248198 , n248191 , n248197 );
or ( n248199 , n248196 , n248190 );
nand ( n248200 , n248198 , n248199 );
and ( n248201 , n248200 , n239941 );
not ( n248202 , n248200 );
not ( n248203 , n239941 );
and ( n248204 , n248202 , n248203 );
nor ( n248205 , n248201 , n248204 );
and ( n248206 , n248183 , n248205 );
not ( n248207 , n248183 );
not ( n248208 , n248205 );
and ( n248209 , n248207 , n248208 );
nor ( n248210 , n248206 , n248209 );
buf ( n248211 , n248210 );
and ( n248212 , n248163 , n248211 );
not ( n248213 , n248163 );
not ( n248214 , n248183 );
not ( n248215 , n248205 );
or ( n248216 , n248214 , n248215 );
not ( n248217 , n248183 );
nand ( n248218 , n248217 , n248208 );
nand ( n248219 , n248216 , n248218 );
buf ( n248220 , n248219 );
and ( n248221 , n248213 , n248220 );
nor ( n248222 , n248212 , n248221 );
nand ( n248223 , n248152 , n248222 );
not ( n248224 , n247144 );
nor ( n248225 , n240239 , n49527 );
not ( n248226 , n248225 );
not ( n248227 , n240225 );
and ( n248228 , n248226 , n248227 );
and ( n248229 , n248225 , n240225 );
nor ( n248230 , n248228 , n248229 );
not ( n248231 , n248230 );
not ( n248232 , n248231 );
not ( n248233 , n49493 );
nand ( n248234 , n248233 , n240264 );
not ( n248235 , n248234 );
not ( n248236 , n240257 );
or ( n248237 , n248235 , n248236 );
or ( n248238 , n240257 , n248234 );
nand ( n248239 , n248237 , n248238 );
not ( n248240 , n248239 );
not ( n248241 , n248240 );
or ( n248242 , n248232 , n248241 );
nand ( n248243 , n248239 , n248230 );
nand ( n248244 , n248242 , n248243 );
not ( n248245 , n240207 );
nand ( n248246 , n248245 , n227211 );
buf ( n248247 , n240195 );
xor ( n248248 , n248246 , n248247 );
and ( n248249 , n248244 , n248248 );
not ( n248250 , n248244 );
not ( n248251 , n248248 );
and ( n248252 , n248250 , n248251 );
nor ( n248253 , n248249 , n248252 );
not ( n248254 , n248253 );
not ( n248255 , n240183 );
nand ( n248256 , n49603 , n240292 );
not ( n248257 , n248256 );
not ( n248258 , n240281 );
and ( n248259 , n248257 , n248258 );
not ( n248260 , n240293 );
nand ( n248261 , n248260 , n49603 );
not ( n248262 , n240282 );
and ( n248263 , n248261 , n248262 );
nor ( n248264 , n248259 , n248263 );
not ( n248265 , n248264 );
or ( n248266 , n248255 , n248265 );
not ( n248267 , n248264 );
not ( n248268 , n240183 );
nand ( n248269 , n248267 , n248268 );
nand ( n248270 , n248266 , n248269 );
not ( n248271 , n248270 );
not ( n248272 , n248271 );
or ( n248273 , n248254 , n248272 );
not ( n248274 , n248253 );
nand ( n248275 , n248274 , n248270 );
nand ( n248276 , n248273 , n248275 );
not ( n248277 , n248276 );
or ( n248278 , n248224 , n248277 );
or ( n248279 , n248276 , n247144 );
nand ( n248280 , n248278 , n248279 );
buf ( n248281 , n247399 );
and ( n248282 , n248280 , n248281 );
not ( n248283 , n248280 );
buf ( n248284 , n247393 );
and ( n248285 , n248283 , n248284 );
nor ( n248286 , n248282 , n248285 );
and ( n248287 , n248223 , n248286 );
not ( n248288 , n248223 );
not ( n248289 , n248286 );
and ( n248290 , n248288 , n248289 );
nor ( n248291 , n248287 , n248290 );
or ( n248292 , n248291 , n245938 );
nand ( n248293 , n248091 , n248292 );
buf ( n248294 , n248293 );
buf ( n248295 , n38087 );
not ( n248296 , n248295 );
not ( n248297 , n30034 );
or ( n248298 , n248296 , n248297 );
not ( n248299 , n248295 );
nand ( n248300 , n248299 , n236320 );
nand ( n248301 , n248298 , n248300 );
and ( n248302 , n248301 , n42760 );
not ( n248303 , n248301 );
and ( n248304 , n248303 , n50452 );
nor ( n248305 , n248302 , n248304 );
not ( n248306 , n248305 );
nand ( n248307 , n246268 , n248306 );
not ( n248308 , n248307 );
not ( n248309 , n239466 );
and ( n248310 , n248308 , n248309 );
and ( n248311 , n248307 , n239466 );
nor ( n248312 , n248310 , n248311 );
not ( n248313 , n248312 );
not ( n248314 , n248313 );
not ( n248315 , n239404 );
xor ( n248316 , n36185 , n36182 );
not ( n248317 , n248316 );
not ( n248318 , n28597 );
or ( n248319 , n248317 , n248318 );
or ( n248320 , n44887 , n248316 );
nand ( n248321 , n248319 , n248320 );
not ( n248322 , n248321 );
not ( n248323 , n28603 );
and ( n248324 , n248322 , n248323 );
and ( n248325 , n248321 , n28557 );
nor ( n248326 , n248324 , n248325 );
not ( n248327 , n248326 );
nand ( n248328 , n239407 , n248327 );
not ( n248329 , n248328 );
or ( n248330 , n248315 , n248329 );
not ( n248331 , n248326 );
nand ( n248332 , n248331 , n239407 );
or ( n248333 , n248332 , n239404 );
nand ( n248334 , n248330 , n248333 );
not ( n248335 , n248334 );
not ( n248336 , n248335 );
or ( n248337 , n248314 , n248336 );
nand ( n248338 , n248334 , n248312 );
nand ( n248339 , n248337 , n248338 );
not ( n248340 , n26222 );
not ( n248341 , n32441 );
not ( n248342 , n38876 );
and ( n248343 , n248341 , n248342 );
and ( n248344 , n32441 , n38876 );
nor ( n248345 , n248343 , n248344 );
not ( n248346 , n248345 );
not ( n248347 , n248346 );
or ( n248348 , n248340 , n248347 );
nand ( n248349 , n222589 , n248345 );
nand ( n248350 , n248348 , n248349 );
nand ( n248351 , n248350 , n244094 );
not ( n248352 , n248351 );
not ( n248353 , n239545 );
and ( n248354 , n248352 , n248353 );
and ( n248355 , n248351 , n239545 );
nor ( n248356 , n248354 , n248355 );
not ( n248357 , n248356 );
buf ( n248358 , n39469 );
not ( n248359 , n248358 );
not ( n248360 , n41681 );
or ( n248361 , n248359 , n248360 );
or ( n248362 , n37506 , n248358 );
nand ( n248363 , n248361 , n248362 );
and ( n248364 , n248363 , n38090 );
not ( n248365 , n248363 );
and ( n248366 , n248365 , n39875 );
nor ( n248367 , n248364 , n248366 );
nand ( n248368 , n248367 , n246295 );
and ( n248369 , n248368 , n246286 );
not ( n248370 , n248368 );
and ( n248371 , n248370 , n239499 );
nor ( n248372 , n248369 , n248371 );
not ( n248373 , n248372 );
or ( n248374 , n248357 , n248373 );
or ( n248375 , n248372 , n248356 );
nand ( n248376 , n248374 , n248375 );
and ( n248377 , n248376 , n246327 );
not ( n248378 , n248376 );
and ( n248379 , n248378 , n246264 );
nor ( n248380 , n248377 , n248379 );
and ( n248381 , n248339 , n248380 );
not ( n248382 , n248339 );
not ( n248383 , n248380 );
and ( n248384 , n248382 , n248383 );
nor ( n248385 , n248381 , n248384 );
buf ( n248386 , n248385 );
not ( n248387 , n248386 );
not ( n248388 , n235094 );
not ( n248389 , n248388 );
not ( n248390 , n235116 );
nand ( n248391 , n43869 , n248390 );
not ( n248392 , n248391 );
not ( n248393 , n43879 );
and ( n248394 , n248392 , n248393 );
and ( n248395 , n248391 , n43879 );
nor ( n248396 , n248394 , n248395 );
not ( n248397 , n248396 );
not ( n248398 , n248397 );
not ( n248399 , n235133 );
not ( n248400 , n43845 );
nand ( n248401 , n248399 , n248400 );
and ( n248402 , n248401 , n43828 );
not ( n248403 , n248401 );
and ( n248404 , n248403 , n43827 );
nor ( n248405 , n248402 , n248404 );
not ( n248406 , n248405 );
not ( n248407 , n248406 );
or ( n248408 , n248398 , n248407 );
nand ( n248409 , n248405 , n248396 );
nand ( n248410 , n248408 , n248409 );
not ( n248411 , n235085 );
nand ( n248412 , n248411 , n43916 );
and ( n248413 , n248412 , n43928 );
not ( n248414 , n248412 );
not ( n248415 , n43928 );
and ( n248416 , n248414 , n248415 );
nor ( n248417 , n248413 , n248416 );
not ( n248418 , n248417 );
and ( n248419 , n248410 , n248418 );
not ( n248420 , n248410 );
and ( n248421 , n248420 , n248417 );
nor ( n248422 , n248419 , n248421 );
nand ( n248423 , n43791 , n235189 );
not ( n248424 , n248423 );
not ( n248425 , n43779 );
and ( n248426 , n248424 , n248425 );
and ( n248427 , n248423 , n43779 );
nor ( n248428 , n248426 , n248427 );
not ( n248429 , n248428 );
not ( n248430 , n248429 );
not ( n248431 , n235160 );
nand ( n248432 , n248431 , n43762 );
and ( n248433 , n248432 , n43749 );
not ( n248434 , n248432 );
and ( n248435 , n248434 , n43748 );
nor ( n248436 , n248433 , n248435 );
not ( n248437 , n248436 );
not ( n248438 , n248437 );
or ( n248439 , n248430 , n248438 );
nand ( n248440 , n248436 , n248428 );
nand ( n248441 , n248439 , n248440 );
and ( n248442 , n248422 , n248441 );
not ( n248443 , n248422 );
not ( n248444 , n248441 );
and ( n248445 , n248443 , n248444 );
nor ( n248446 , n248442 , n248445 );
not ( n248447 , n248446 );
or ( n248448 , n248389 , n248447 );
not ( n248449 , n248388 );
not ( n248450 , n248444 );
not ( n248451 , n248422 );
not ( n248452 , n248451 );
or ( n248453 , n248450 , n248452 );
nand ( n248454 , n248422 , n248441 );
nand ( n248455 , n248453 , n248454 );
nand ( n248456 , n248449 , n248455 );
nand ( n248457 , n248448 , n248456 );
not ( n248458 , n248457 );
or ( n248459 , n248387 , n248458 );
or ( n248460 , n248457 , n248386 );
nand ( n248461 , n248459 , n248460 );
not ( n248462 , n38616 );
not ( n248463 , n234521 );
or ( n248464 , n248462 , n248463 );
or ( n248465 , n234521 , n38616 );
nand ( n248466 , n248464 , n248465 );
and ( n248467 , n248466 , n243427 );
not ( n248468 , n248466 );
and ( n248469 , n248468 , n243431 );
nor ( n248470 , n248467 , n248469 );
nand ( n248471 , n248461 , n248470 );
not ( n248472 , n247468 );
not ( n248473 , n243510 );
or ( n248474 , n248472 , n248473 );
not ( n248475 , n247468 );
nand ( n248476 , n248475 , n243503 );
nand ( n248477 , n248474 , n248476 );
buf ( n248478 , n243810 );
and ( n248479 , n248477 , n248478 );
not ( n248480 , n248477 );
buf ( n248481 , n243801 );
and ( n248482 , n248480 , n248481 );
nor ( n248483 , n248479 , n248482 );
nor ( n248484 , n248483 , n234021 );
not ( n248485 , n248484 );
or ( n248486 , n248471 , n248485 );
not ( n248487 , n248483 );
nor ( n248488 , n248487 , n236795 );
nand ( n248489 , n248471 , n248488 );
nand ( n248490 , n39767 , n41384 );
nand ( n248491 , n248486 , n248489 , n248490 );
buf ( n248492 , n248491 );
not ( n248493 , n224011 );
not ( n248494 , n248493 );
not ( n248495 , n223967 );
not ( n248496 , n46228 );
nand ( n248497 , n248495 , n248496 );
and ( n248498 , n248497 , n243533 );
not ( n248499 , n248497 );
not ( n248500 , n243533 );
and ( n248501 , n248499 , n248500 );
nor ( n248502 , n248498 , n248501 );
not ( n248503 , n248502 );
not ( n248504 , n248503 );
not ( n248505 , n224024 );
not ( n248506 , n46289 );
nand ( n248507 , n248505 , n248506 );
not ( n248508 , n248507 );
not ( n248509 , n243562 );
and ( n248510 , n248508 , n248509 );
and ( n248511 , n248507 , n243562 );
nor ( n248512 , n248510 , n248511 );
not ( n248513 , n248512 );
not ( n248514 , n248513 );
or ( n248515 , n248504 , n248514 );
nand ( n248516 , n248512 , n248502 );
nand ( n248517 , n248515 , n248516 );
not ( n248518 , n224085 );
nand ( n248519 , n248518 , n224068 );
and ( n248520 , n248519 , n243581 );
not ( n248521 , n248519 );
and ( n248522 , n248521 , n243580 );
nor ( n248523 , n248520 , n248522 );
not ( n248524 , n248523 );
and ( n248525 , n248517 , n248524 );
not ( n248526 , n248517 );
and ( n248527 , n248526 , n248523 );
nor ( n248528 , n248525 , n248527 );
not ( n248529 , n248528 );
not ( n248530 , n46340 );
nand ( n248531 , n248530 , n46353 );
not ( n248532 , n248531 );
not ( n248533 , n243631 );
not ( n248534 , n248533 );
and ( n248535 , n248532 , n248534 );
and ( n248536 , n248531 , n248533 );
nor ( n248537 , n248535 , n248536 );
not ( n248538 , n248537 );
not ( n248539 , n46404 );
nand ( n248540 , n248539 , n46374 );
not ( n248541 , n248540 );
not ( n248542 , n243614 );
not ( n248543 , n248542 );
and ( n248544 , n248541 , n248543 );
and ( n248545 , n248540 , n248542 );
nor ( n248546 , n248544 , n248545 );
not ( n248547 , n248546 );
not ( n248548 , n248547 );
or ( n248549 , n248538 , n248548 );
not ( n248550 , n248537 );
nand ( n248551 , n248550 , n248546 );
nand ( n248552 , n248549 , n248551 );
not ( n248553 , n248552 );
and ( n248554 , n248529 , n248553 );
not ( n248555 , n248529 );
and ( n248556 , n248555 , n248552 );
nor ( n248557 , n248554 , n248556 );
not ( n248558 , n248557 );
or ( n248559 , n248494 , n248558 );
not ( n248560 , n248493 );
not ( n248561 , n248553 );
not ( n248562 , n248529 );
or ( n248563 , n248561 , n248562 );
nand ( n248564 , n248528 , n248552 );
nand ( n248565 , n248563 , n248564 );
nand ( n248566 , n248560 , n248565 );
nand ( n248567 , n248559 , n248566 );
nand ( n248568 , n243037 , n243026 );
not ( n248569 , n36811 );
not ( n248570 , n248569 );
not ( n248571 , n42624 );
or ( n248572 , n248570 , n248571 );
or ( n248573 , n42624 , n248569 );
nand ( n248574 , n248572 , n248573 );
and ( n248575 , n248574 , n45817 );
not ( n248576 , n248574 );
and ( n248577 , n248576 , n45818 );
nor ( n248578 , n248575 , n248577 );
and ( n248579 , n248568 , n248578 );
not ( n248580 , n248568 );
not ( n248581 , n248578 );
and ( n248582 , n248580 , n248581 );
nor ( n248583 , n248579 , n248582 );
not ( n248584 , n248583 );
not ( n248585 , n248584 );
nand ( n248586 , n243073 , n243062 );
not ( n248587 , n248586 );
not ( n248588 , n31036 );
not ( n248589 , n48070 );
and ( n248590 , n248588 , n248589 );
and ( n248591 , n33186 , n48070 );
nor ( n248592 , n248590 , n248591 );
and ( n248593 , n248592 , n31078 );
not ( n248594 , n248592 );
and ( n248595 , n248594 , n31081 );
nor ( n248596 , n248593 , n248595 );
not ( n248597 , n248596 );
and ( n248598 , n248587 , n248597 );
and ( n248599 , n248586 , n248596 );
nor ( n248600 , n248598 , n248599 );
not ( n248601 , n248600 );
not ( n248602 , n248601 );
or ( n248603 , n248585 , n248602 );
nand ( n248604 , n248600 , n248583 );
nand ( n248605 , n248603 , n248604 );
not ( n248606 , n248605 );
not ( n248607 , n248606 );
not ( n248608 , n28716 );
not ( n248609 , n32961 );
or ( n248610 , n248608 , n248609 );
not ( n248611 , n28716 );
not ( n248612 , n32961 );
nand ( n248613 , n248611 , n248612 );
nand ( n248614 , n248610 , n248613 );
and ( n248615 , n248614 , n32989 );
not ( n248616 , n248614 );
and ( n248617 , n248616 , n54623 );
nor ( n248618 , n248615 , n248617 );
not ( n248619 , n248618 );
not ( n248620 , n248619 );
not ( n248621 , n243102 );
nand ( n248622 , n248621 , n243114 );
not ( n248623 , n248622 );
or ( n248624 , n248620 , n248623 );
nand ( n248625 , n248621 , n243114 );
or ( n248626 , n248625 , n248619 );
nand ( n248627 , n248624 , n248626 );
not ( n248628 , n248627 );
nand ( n248629 , n243182 , n243167 );
not ( n248630 , n248629 );
not ( n248631 , n207918 );
not ( n248632 , n219116 );
or ( n248633 , n248631 , n248632 );
not ( n248634 , n207918 );
nand ( n248635 , n248634 , n219115 );
nand ( n248636 , n248633 , n248635 );
and ( n248637 , n248636 , n52705 );
not ( n248638 , n248636 );
and ( n248639 , n248638 , n27716 );
nor ( n248640 , n248637 , n248639 );
not ( n248641 , n248640 );
and ( n248642 , n248630 , n248641 );
and ( n248643 , n248629 , n248640 );
nor ( n248644 , n248642 , n248643 );
not ( n248645 , n248644 );
or ( n248646 , n248628 , n248645 );
or ( n248647 , n248644 , n248627 );
nand ( n248648 , n248646 , n248647 );
not ( n248649 , n243127 );
nand ( n248650 , n248649 , n243149 );
not ( n248651 , n248650 );
not ( n248652 , n28665 );
buf ( n248653 , n29635 );
not ( n248654 , n248653 );
not ( n248655 , n45404 );
or ( n248656 , n248654 , n248655 );
or ( n248657 , n45404 , n248653 );
nand ( n248658 , n248656 , n248657 );
not ( n248659 , n248658 );
and ( n248660 , n248652 , n248659 );
and ( n248661 , n28665 , n248658 );
nor ( n248662 , n248660 , n248661 );
not ( n248663 , n248662 );
not ( n248664 , n248663 );
and ( n248665 , n248651 , n248664 );
and ( n248666 , n248650 , n248663 );
nor ( n248667 , n248665 , n248666 );
not ( n248668 , n248667 );
and ( n248669 , n248648 , n248668 );
not ( n248670 , n248648 );
and ( n248671 , n248670 , n248667 );
nor ( n248672 , n248669 , n248671 );
not ( n248673 , n248672 );
or ( n248674 , n248607 , n248673 );
not ( n248675 , n248672 );
nand ( n248676 , n248675 , n248605 );
nand ( n248677 , n248674 , n248676 );
buf ( n248678 , n248677 );
not ( n248679 , n248678 );
and ( n248680 , n248567 , n248679 );
not ( n248681 , n248567 );
and ( n248682 , n248681 , n248678 );
nor ( n248683 , n248680 , n248682 );
nor ( n248684 , n248683 , n35427 );
not ( n248685 , n47899 );
not ( n248686 , n48676 );
or ( n248687 , n248685 , n248686 );
not ( n248688 , n47899 );
nand ( n248689 , n248688 , n48686 );
nand ( n248690 , n248687 , n248689 );
and ( n248691 , n248690 , n48797 );
not ( n248692 , n248690 );
and ( n248693 , n248692 , n48806 );
nor ( n248694 , n248691 , n248693 );
not ( n248695 , n242175 );
not ( n248696 , n27876 );
or ( n248697 , n248695 , n248696 );
not ( n248698 , n242175 );
nand ( n248699 , n248698 , n27869 );
nand ( n248700 , n248697 , n248699 );
not ( n248701 , n55574 );
nand ( n248702 , n55586 , n236920 );
not ( n248703 , n248702 );
or ( n248704 , n248701 , n248703 );
or ( n248705 , n248702 , n55574 );
nand ( n248706 , n248704 , n248705 );
not ( n248707 , n248706 );
not ( n248708 , n55543 );
nand ( n248709 , n248708 , n236900 );
not ( n248710 , n248709 );
not ( n248711 , n233319 );
and ( n248712 , n248710 , n248711 );
not ( n248713 , n236899 );
nand ( n248714 , n248713 , n248708 );
and ( n248715 , n248714 , n233319 );
nor ( n248716 , n248712 , n248715 );
not ( n248717 , n248716 );
or ( n248718 , n248707 , n248717 );
or ( n248719 , n248716 , n248706 );
nand ( n248720 , n248718 , n248719 );
nand ( n248721 , n236943 , n239282 );
buf ( n248722 , n233386 );
and ( n248723 , n248721 , n248722 );
not ( n248724 , n248721 );
not ( n248725 , n248722 );
and ( n248726 , n248724 , n248725 );
nor ( n248727 , n248723 , n248726 );
not ( n248728 , n248727 );
and ( n248729 , n248720 , n248728 );
not ( n248730 , n248720 );
and ( n248731 , n248730 , n248727 );
nor ( n248732 , n248729 , n248731 );
and ( n248733 , n236967 , n55701 );
and ( n248734 , n248733 , n55692 );
not ( n248735 , n248733 );
and ( n248736 , n248735 , n234984 );
nor ( n248737 , n248734 , n248736 );
not ( n248738 , n248737 );
not ( n248739 , n248738 );
not ( n248740 , n55666 );
nand ( n248741 , n248740 , n236978 );
and ( n248742 , n248741 , n55652 );
not ( n248743 , n248741 );
and ( n248744 , n248743 , n234965 );
nor ( n248745 , n248742 , n248744 );
not ( n248746 , n248745 );
not ( n248747 , n248746 );
or ( n248748 , n248739 , n248747 );
nand ( n248749 , n248745 , n248737 );
nand ( n248750 , n248748 , n248749 );
and ( n248751 , n248732 , n248750 );
not ( n248752 , n248732 );
not ( n248753 , n248750 );
and ( n248754 , n248752 , n248753 );
nor ( n248755 , n248751 , n248754 );
buf ( n248756 , n248755 );
and ( n248757 , n248700 , n248756 );
not ( n248758 , n248700 );
and ( n248759 , n248732 , n248753 );
not ( n248760 , n248732 );
and ( n248761 , n248760 , n248750 );
nor ( n248762 , n248759 , n248761 );
buf ( n248763 , n248762 );
and ( n248764 , n248758 , n248763 );
nor ( n248765 , n248757 , n248764 );
nand ( n248766 , n248684 , n248694 , n248765 );
not ( n248767 , n248683 );
not ( n248768 , n248767 );
not ( n248769 , n248694 );
or ( n248770 , n248768 , n248769 );
nor ( n248771 , n248765 , n40465 );
nand ( n248772 , n248770 , n248771 );
nand ( n248773 , n31577 , n204636 );
nand ( n248774 , n248766 , n248772 , n248773 );
buf ( n248775 , n248774 );
not ( n248776 , n42690 );
not ( n248777 , n237647 );
or ( n248778 , n248776 , n248777 );
not ( n248779 , n42689 );
or ( n248780 , n237647 , n248779 );
nand ( n248781 , n248778 , n248780 );
not ( n248782 , n248781 );
not ( n248783 , n237701 );
and ( n248784 , n248782 , n248783 );
and ( n248785 , n248781 , n241677 );
nor ( n248786 , n248784 , n248785 );
nand ( n248787 , n248786 , n243233 );
buf ( n248788 , n245811 );
not ( n248789 , n248788 );
not ( n248790 , n39444 );
or ( n248791 , n248789 , n248790 );
or ( n248792 , n39444 , n248788 );
nand ( n248793 , n248791 , n248792 );
not ( n248794 , n248793 );
buf ( n248795 , n52982 );
not ( n248796 , n248795 );
and ( n248797 , n248794 , n248796 );
and ( n248798 , n248793 , n248795 );
nor ( n248799 , n248797 , n248798 );
not ( n248800 , n248799 );
not ( n248801 , n42139 );
not ( n248802 , n234243 );
or ( n248803 , n248801 , n248802 );
not ( n248804 , n42139 );
nand ( n248805 , n248804 , n234252 );
nand ( n248806 , n248803 , n248805 );
and ( n248807 , n248806 , n234299 );
not ( n248808 , n248806 );
and ( n248809 , n248808 , n234306 );
nor ( n248810 , n248807 , n248809 );
not ( n248811 , n248810 );
nand ( n248812 , n248800 , n248811 );
or ( n248813 , n248787 , n248812 );
not ( n248814 , n248800 );
not ( n248815 , n248786 );
or ( n248816 , n248814 , n248815 );
nor ( n248817 , n248811 , n35427 );
nand ( n248818 , n248816 , n248817 );
nand ( n248819 , n237714 , n41122 );
nand ( n248820 , n248813 , n248818 , n248819 );
buf ( n248821 , n248820 );
buf ( n248822 , n25494 );
not ( n248823 , RI19ab8958_2391);
or ( n248824 , n25328 , n248823 );
not ( n248825 , RI19aaeb60_2463);
or ( n248826 , n25336 , n248825 );
nand ( n248827 , n248824 , n248826 );
buf ( n248828 , n248827 );
not ( n248829 , RI19ab4bf0_2418);
or ( n248830 , n233507 , n248829 );
not ( n248831 , RI19aaad80_2489);
or ( n248832 , n25335 , n248831 );
nand ( n248833 , n248830 , n248832 );
buf ( n248834 , n248833 );
buf ( n248835 , n33654 );
not ( n248836 , n241778 );
not ( n248837 , n248836 );
nand ( n248838 , n241802 , n241799 );
and ( n248839 , n248838 , n237162 );
not ( n248840 , n248838 );
not ( n248841 , n237162 );
and ( n248842 , n248840 , n248841 );
nor ( n248843 , n248839 , n248842 );
not ( n248844 , n248843 );
not ( n248845 , n248844 );
not ( n248846 , n237208 );
nand ( n248847 , n241850 , n248846 );
not ( n248848 , n237198 );
and ( n248849 , n248847 , n248848 );
not ( n248850 , n248847 );
and ( n248851 , n248850 , n237198 );
nor ( n248852 , n248849 , n248851 );
not ( n248853 , n248852 );
not ( n248854 , n248853 );
or ( n248855 , n248845 , n248854 );
nand ( n248856 , n248852 , n248843 );
nand ( n248857 , n248855 , n248856 );
nand ( n248858 , n241809 , n241831 );
not ( n248859 , n248858 );
not ( n248860 , n237239 );
not ( n248861 , n248860 );
and ( n248862 , n248859 , n248861 );
and ( n248863 , n248858 , n248860 );
nor ( n248864 , n248862 , n248863 );
not ( n248865 , n248864 );
and ( n248866 , n248857 , n248865 );
not ( n248867 , n248857 );
and ( n248868 , n248867 , n248864 );
nor ( n248869 , n248866 , n248868 );
not ( n248870 , n237276 );
not ( n248871 , n248870 );
nand ( n248872 , n244746 , n237285 );
not ( n248873 , n248872 );
or ( n248874 , n248871 , n248873 );
or ( n248875 , n248872 , n248870 );
nand ( n248876 , n248874 , n248875 );
not ( n248877 , n248876 );
nand ( n248878 , n237313 , n244736 );
not ( n248879 , n248878 );
not ( n248880 , n237302 );
and ( n248881 , n248879 , n248880 );
and ( n248882 , n248878 , n237302 );
nor ( n248883 , n248881 , n248882 );
not ( n248884 , n248883 );
and ( n248885 , n248877 , n248884 );
and ( n248886 , n248876 , n248883 );
nor ( n248887 , n248885 , n248886 );
and ( n248888 , n248869 , n248887 );
not ( n248889 , n248869 );
not ( n248890 , n248887 );
and ( n248891 , n248889 , n248890 );
nor ( n248892 , n248888 , n248891 );
not ( n248893 , n248892 );
or ( n248894 , n248837 , n248893 );
not ( n248895 , n248836 );
not ( n248896 , n248887 );
not ( n248897 , n248869 );
or ( n248898 , n248896 , n248897 );
not ( n248899 , n248869 );
nand ( n248900 , n248899 , n248890 );
nand ( n248901 , n248898 , n248900 );
nand ( n248902 , n248895 , n248901 );
nand ( n248903 , n248894 , n248902 );
buf ( n248904 , n229763 );
and ( n248905 , n248903 , n248904 );
not ( n248906 , n248903 );
not ( n248907 , n229763 );
and ( n248908 , n248906 , n248907 );
nor ( n248909 , n248905 , n248908 );
not ( n248910 , n248909 );
not ( n248911 , n248910 );
not ( n248912 , n50089 );
not ( n248913 , n235984 );
not ( n248914 , n227845 );
nand ( n248915 , n248914 , n227810 );
not ( n248916 , n248915 );
or ( n248917 , n248913 , n248916 );
not ( n248918 , n227809 );
nand ( n248919 , n248918 , n248914 );
or ( n248920 , n248919 , n235984 );
nand ( n248921 , n248917 , n248920 );
not ( n248922 , n248921 );
nand ( n248923 , n50170 , n50146 );
and ( n248924 , n248923 , n236010 );
not ( n248925 , n248923 );
and ( n248926 , n248925 , n236009 );
nor ( n248927 , n248924 , n248926 );
not ( n248928 , n248927 );
and ( n248929 , n248922 , n248928 );
and ( n248930 , n248921 , n248927 );
nor ( n248931 , n248929 , n248930 );
not ( n248932 , n248931 );
not ( n248933 , n235944 );
nand ( n248934 , n50218 , n50202 );
not ( n248935 , n248934 );
or ( n248936 , n248933 , n248935 );
or ( n248937 , n248934 , n235944 );
nand ( n248938 , n248936 , n248937 );
not ( n248939 , n248938 );
nand ( n248940 , n227862 , n50125 );
not ( n248941 , n248940 );
not ( n248942 , n236040 );
and ( n248943 , n248941 , n248942 );
and ( n248944 , n248940 , n236040 );
nor ( n248945 , n248943 , n248944 );
not ( n248946 , n248945 );
or ( n248947 , n248939 , n248946 );
or ( n248948 , n248945 , n248938 );
nand ( n248949 , n248947 , n248948 );
not ( n248950 , n50231 );
not ( n248951 , n50259 );
nand ( n248952 , n248950 , n248951 );
and ( n248953 , n248952 , n235970 );
not ( n248954 , n248952 );
and ( n248955 , n248954 , n235971 );
nor ( n248956 , n248953 , n248955 );
not ( n248957 , n248956 );
and ( n248958 , n248949 , n248957 );
not ( n248959 , n248949 );
and ( n248960 , n248959 , n248956 );
nor ( n248961 , n248958 , n248960 );
not ( n248962 , n248961 );
not ( n248963 , n248962 );
or ( n248964 , n248932 , n248963 );
not ( n248965 , n248931 );
nand ( n248966 , n248961 , n248965 );
nand ( n248967 , n248964 , n248966 );
not ( n248968 , n248967 );
or ( n248969 , n248912 , n248968 );
or ( n248970 , n248967 , n50089 );
nand ( n248971 , n248969 , n248970 );
buf ( n248972 , n53820 );
and ( n248973 , n248971 , n248972 );
not ( n248974 , n248971 );
buf ( n248975 , n53811 );
and ( n248976 , n248974 , n248975 );
nor ( n248977 , n248973 , n248976 );
not ( n248978 , n248977 );
not ( n248979 , n248978 );
or ( n248980 , n248911 , n248979 );
not ( n248981 , n235732 );
nand ( n248982 , n248980 , n248981 );
not ( n248983 , n39105 );
not ( n248984 , n246826 );
or ( n248985 , n248983 , n248984 );
not ( n248986 , n39105 );
nand ( n248987 , n248986 , n246835 );
nand ( n248988 , n248985 , n248987 );
and ( n248989 , n248988 , n246883 );
not ( n248990 , n248988 );
and ( n248991 , n248990 , n246892 );
nor ( n248992 , n248989 , n248991 );
or ( n248993 , n248982 , n248992 );
nor ( n248994 , n248909 , n243434 );
nand ( n248995 , n248978 , n248994 , n248992 );
nand ( n248996 , n31577 , n28738 );
nand ( n248997 , n248993 , n248995 , n248996 );
buf ( n248998 , n248997 );
buf ( n248999 , n36182 );
nand ( n249000 , n242447 , n243316 );
not ( n249001 , n249000 );
not ( n249002 , n241524 );
and ( n249003 , n249001 , n249002 );
and ( n249004 , n249000 , n241524 );
nor ( n249005 , n249003 , n249004 );
not ( n249006 , n242569 );
xor ( n249007 , n249005 , n249006 );
xor ( n249008 , n249007 , n242520 );
not ( n249009 , n234021 );
nand ( n249010 , n249008 , n249009 );
not ( n249011 , n244378 );
not ( n249012 , n55194 );
not ( n249013 , n239398 );
or ( n249014 , n249012 , n249013 );
not ( n249015 , n55194 );
nand ( n249016 , n249015 , n239390 );
nand ( n249017 , n249014 , n249016 );
buf ( n249018 , n53081 );
and ( n249019 , n249017 , n249018 );
not ( n249020 , n249017 );
buf ( n249021 , n53080 );
and ( n249022 , n249020 , n249021 );
nor ( n249023 , n249019 , n249022 );
not ( n249024 , n249023 );
nand ( n249025 , n249011 , n249024 );
or ( n249026 , n249010 , n249025 );
not ( n249027 , n249011 );
not ( n249028 , n249008 );
or ( n249029 , n249027 , n249028 );
not ( n249030 , n205649 );
nor ( n249031 , n249024 , n249030 );
nand ( n249032 , n249029 , n249031 );
nand ( n249033 , n39766 , n30491 );
nand ( n249034 , n249026 , n249032 , n249033 );
buf ( n249035 , n249034 );
buf ( n249036 , n33437 );
buf ( n249037 , n32043 );
not ( n249038 , RI19ac04a0_2329);
or ( n249039 , n25328 , n249038 );
not ( n249040 , RI19ab7530_2399);
or ( n249041 , n226822 , n249040 );
nand ( n249042 , n249039 , n249041 );
buf ( n249043 , n249042 );
buf ( n249044 , n33218 );
buf ( n249045 , n25535 );
buf ( n249046 , n33780 );
nand ( n249047 , n237264 , n248870 );
and ( n249048 , n249047 , n244742 );
not ( n249049 , n249047 );
and ( n249050 , n249049 , n241772 );
nor ( n249051 , n249048 , n249050 );
not ( n249052 , n249051 );
not ( n249053 , n249052 );
not ( n249054 , n244768 );
or ( n249055 , n249053 , n249054 );
or ( n249056 , n244768 , n249052 );
nand ( n249057 , n249055 , n249056 );
not ( n249058 , n249057 );
buf ( n249059 , n239705 );
not ( n249060 , n249059 );
and ( n249061 , n249058 , n249060 );
and ( n249062 , n249057 , n249059 );
nor ( n249063 , n249061 , n249062 );
not ( n249064 , n249063 );
nor ( n249065 , n249064 , n31572 );
not ( n249066 , n49291 );
not ( n249067 , n31397 );
not ( n249068 , n39501 );
not ( n249069 , n249068 );
or ( n249070 , n249067 , n249069 );
or ( n249071 , n39320 , n31397 );
nand ( n249072 , n249070 , n249071 );
and ( n249073 , n249072 , n39327 );
not ( n249074 , n249072 );
and ( n249075 , n249074 , n204825 );
nor ( n249076 , n249073 , n249075 );
nand ( n249077 , n249066 , n249076 );
not ( n249078 , n249077 );
not ( n249079 , n247096 );
and ( n249080 , n249078 , n249079 );
not ( n249081 , n49291 );
nand ( n249082 , n249081 , n249076 );
and ( n249083 , n249082 , n247096 );
nor ( n249084 , n249080 , n249083 );
not ( n249085 , n249084 );
not ( n249086 , n249085 );
not ( n249087 , n227174 );
or ( n249088 , n249086 , n249087 );
not ( n249089 , n249085 );
nand ( n249090 , n249089 , n49420 );
nand ( n249091 , n249088 , n249090 );
and ( n249092 , n249091 , n49618 );
not ( n249093 , n249091 );
and ( n249094 , n249093 , n49627 );
nor ( n249095 , n249092 , n249094 );
not ( n249096 , n249095 );
nand ( n249097 , n249065 , n249096 );
nor ( n249098 , n249063 , n55146 );
not ( n249099 , n225178 );
nand ( n249100 , n225185 , n249099 );
and ( n249101 , n249100 , n48284 );
not ( n249102 , n249100 );
not ( n249103 , n48284 );
and ( n249104 , n249102 , n249103 );
nor ( n249105 , n249101 , n249104 );
not ( n249106 , n249105 );
not ( n249107 , n245949 );
or ( n249108 , n249106 , n249107 );
not ( n249109 , n249105 );
nand ( n249110 , n249109 , n48414 );
nand ( n249111 , n249108 , n249110 );
and ( n249112 , n249111 , n226320 );
not ( n249113 , n249111 );
and ( n249114 , n249113 , n226319 );
nor ( n249115 , n249112 , n249114 );
nor ( n249116 , n249096 , n249115 );
nand ( n249117 , n249098 , n249116 );
nor ( n249118 , n249095 , n40465 );
nand ( n249119 , n249118 , n249115 );
nand ( n249120 , n233501 , n47872 );
nand ( n249121 , n249097 , n249117 , n249119 , n249120 );
buf ( n249122 , n249121 );
nand ( n249123 , n229128 , RI1754a6a8_69);
not ( n249124 , RI1754a720_68);
nand ( n249125 , n51363 , n249124 );
and ( n249126 , n249123 , n249125 );
nand ( n249127 , n51363 , RI1754a6a8_69 , RI1754a5b8_71);
and ( n249128 , n249126 , n249127 );
not ( n249129 , RI1754b530_38);
or ( n249130 , n249128 , n249129 );
not ( n249131 , n25335 );
nand ( n249132 , n249131 , n29917 );
nand ( n249133 , n249130 , n249132 );
buf ( n249134 , n249133 );
not ( n249135 , n247678 );
not ( n249136 , n48019 );
or ( n249137 , n249135 , n249136 );
or ( n249138 , n48019 , n247678 );
nand ( n249139 , n249137 , n249138 );
not ( n249140 , n249139 );
not ( n249141 , n48233 );
and ( n249142 , n249140 , n249141 );
and ( n249143 , n249139 , n48238 );
nor ( n249144 , n249142 , n249143 );
not ( n249145 , n237331 );
nand ( n249146 , n237251 , n248860 );
not ( n249147 , n249146 );
not ( n249148 , n241821 );
and ( n249149 , n249147 , n249148 );
and ( n249150 , n249146 , n241821 );
nor ( n249151 , n249149 , n249150 );
not ( n249152 , n249151 );
not ( n249153 , n237212 );
nand ( n249154 , n249153 , n248848 );
and ( n249155 , n249154 , n241860 );
not ( n249156 , n249154 );
and ( n249157 , n249156 , n241861 );
nor ( n249158 , n249155 , n249157 );
not ( n249159 , n249158 );
or ( n249160 , n249152 , n249159 );
or ( n249161 , n249158 , n249151 );
nand ( n249162 , n249160 , n249161 );
not ( n249163 , n249162 );
not ( n249164 , n249163 );
not ( n249165 , n237183 );
nand ( n249166 , n249165 , n248841 );
not ( n249167 , n249166 );
not ( n249168 , n241789 );
and ( n249169 , n249167 , n249168 );
not ( n249170 , n237183 );
nand ( n249171 , n249170 , n248841 );
and ( n249172 , n249171 , n241789 );
nor ( n249173 , n249169 , n249172 );
not ( n249174 , n249173 );
not ( n249175 , n249174 );
not ( n249176 , n237325 );
nand ( n249177 , n237302 , n249176 );
and ( n249178 , n249177 , n241736 );
not ( n249179 , n249177 );
and ( n249180 , n249179 , n241737 );
nor ( n249181 , n249178 , n249180 );
not ( n249182 , n249181 );
not ( n249183 , n249182 );
or ( n249184 , n249175 , n249183 );
nand ( n249185 , n249173 , n249181 );
nand ( n249186 , n249184 , n249185 );
and ( n249187 , n249186 , n249051 );
not ( n249188 , n249186 );
and ( n249189 , n249188 , n249052 );
nor ( n249190 , n249187 , n249189 );
not ( n249191 , n249190 );
or ( n249192 , n249164 , n249191 );
or ( n249193 , n249190 , n249163 );
nand ( n249194 , n249192 , n249193 );
not ( n249195 , n249194 );
not ( n249196 , n249195 );
or ( n249197 , n249145 , n249196 );
not ( n249198 , n237331 );
not ( n249199 , n249162 );
not ( n249200 , n249190 );
not ( n249201 , n249200 );
or ( n249202 , n249199 , n249201 );
nand ( n249203 , n249190 , n249163 );
nand ( n249204 , n249202 , n249203 );
nand ( n249205 , n249198 , n249204 );
nand ( n249206 , n249197 , n249205 );
buf ( n249207 , n244574 );
not ( n249208 , n249207 );
and ( n249209 , n249206 , n249208 );
not ( n249210 , n249206 );
and ( n249211 , n249210 , n249207 );
nor ( n249212 , n249209 , n249211 );
not ( n249213 , n249212 );
nand ( n249214 , n249144 , n249213 );
or ( n249215 , n239935 , n249214 );
not ( n249216 , n249144 );
not ( n249217 , n239933 );
or ( n249218 , n249216 , n249217 );
nor ( n249219 , n249213 , n53680 );
nand ( n249220 , n249218 , n249219 );
nand ( n249221 , n244484 , n28006 );
nand ( n249222 , n249215 , n249220 , n249221 );
buf ( n249223 , n249222 );
not ( n249224 , n234654 );
nand ( n249225 , n234667 , n249224 );
and ( n249226 , n249225 , n244868 );
not ( n249227 , n249225 );
and ( n249228 , n249227 , n53647 );
nor ( n249229 , n249226 , n249228 );
not ( n249230 , n249229 );
nand ( n249231 , n234638 , n234552 );
not ( n249232 , n249231 );
not ( n249233 , n53594 );
and ( n249234 , n249232 , n249233 );
and ( n249235 , n249231 , n53594 );
nor ( n249236 , n249234 , n249235 );
not ( n249237 , n249236 );
or ( n249238 , n249230 , n249237 );
not ( n249239 , n249229 );
not ( n249240 , n249236 );
nand ( n249241 , n249239 , n249240 );
nand ( n249242 , n249238 , n249241 );
not ( n249243 , n249242 );
not ( n249244 , n249243 );
not ( n249245 , n53516 );
nand ( n249246 , n234569 , n234580 );
not ( n249247 , n249246 );
or ( n249248 , n249245 , n249247 );
or ( n249249 , n249246 , n53516 );
nand ( n249250 , n249248 , n249249 );
not ( n249251 , n249250 );
nand ( n249252 , n234596 , n234608 );
not ( n249253 , n249252 );
buf ( n249254 , n53556 );
not ( n249255 , n249254 );
and ( n249256 , n249253 , n249255 );
not ( n249257 , n234609 );
nand ( n249258 , n249257 , n234596 );
and ( n249259 , n249258 , n249254 );
nor ( n249260 , n249256 , n249259 );
not ( n249261 , n249260 );
or ( n249262 , n249251 , n249261 );
or ( n249263 , n249260 , n249250 );
nand ( n249264 , n249262 , n249263 );
and ( n249265 , n249264 , n244848 );
not ( n249266 , n249264 );
not ( n249267 , n244848 );
and ( n249268 , n249266 , n249267 );
nor ( n249269 , n249265 , n249268 );
not ( n249270 , n249269 );
or ( n249271 , n249244 , n249270 );
or ( n249272 , n249269 , n249243 );
nand ( n249273 , n249271 , n249272 );
buf ( n249274 , n249273 );
not ( n249275 , n249274 );
not ( n249276 , n247870 );
and ( n249277 , n237504 , n249276 );
not ( n249278 , n237504 );
and ( n249279 , n249278 , n247870 );
nor ( n249280 , n249277 , n249279 );
not ( n249281 , n249280 );
or ( n249282 , n249275 , n249281 );
not ( n249283 , n249280 );
not ( n249284 , n249273 );
buf ( n249285 , n249284 );
nand ( n249286 , n249283 , n249285 );
nand ( n249287 , n249282 , n249286 );
not ( n249288 , n54208 );
nand ( n249289 , n249287 , n249288 );
not ( n249290 , n242261 );
not ( n249291 , n230899 );
not ( n249292 , n53112 );
not ( n249293 , n249292 );
or ( n249294 , n249291 , n249293 );
not ( n249295 , n249292 );
not ( n249296 , n230899 );
nand ( n249297 , n249295 , n249296 );
nand ( n249298 , n249294 , n249297 );
not ( n249299 , n249298 );
or ( n249300 , n249290 , n249299 );
not ( n249301 , n242261 );
nand ( n249302 , n249301 , n53140 );
nand ( n249303 , n249300 , n249302 );
or ( n249304 , n221652 , n235107 );
and ( n249305 , n249304 , n248390 );
not ( n249306 , n249304 );
and ( n249307 , n249306 , n235116 );
nor ( n249308 , n249305 , n249307 );
not ( n249309 , n249308 );
not ( n249310 , n249309 );
not ( n249311 , n235143 );
nand ( n249312 , n43859 , n249311 );
and ( n249313 , n249312 , n235133 );
not ( n249314 , n249312 );
and ( n249315 , n249314 , n248399 );
nor ( n249316 , n249313 , n249315 );
not ( n249317 , n249316 );
not ( n249318 , n249317 );
or ( n249319 , n249310 , n249318 );
nand ( n249320 , n249316 , n249308 );
nand ( n249321 , n249319 , n249320 );
nand ( n249322 , n221702 , n235082 );
and ( n249323 , n249322 , n248411 );
not ( n249324 , n249322 );
and ( n249325 , n249324 , n235085 );
nor ( n249326 , n249323 , n249325 );
and ( n249327 , n249321 , n249326 );
not ( n249328 , n249321 );
not ( n249329 , n249326 );
and ( n249330 , n249328 , n249329 );
nor ( n249331 , n249327 , n249330 );
not ( n249332 , n249331 );
not ( n249333 , n249332 );
not ( n249334 , n235184 );
not ( n249335 , n249334 );
not ( n249336 , n235176 );
nand ( n249337 , n249336 , n221567 );
not ( n249338 , n249337 );
or ( n249339 , n249335 , n249338 );
not ( n249340 , n221566 );
nand ( n249341 , n249340 , n249336 );
or ( n249342 , n249341 , n249334 );
nand ( n249343 , n249339 , n249342 );
not ( n249344 , n249343 );
not ( n249345 , n235168 );
nand ( n249346 , n43737 , n249345 );
not ( n249347 , n249346 );
not ( n249348 , n248431 );
and ( n249349 , n249347 , n249348 );
not ( n249350 , n235168 );
nand ( n249351 , n249350 , n43737 );
and ( n249352 , n249351 , n248431 );
nor ( n249353 , n249349 , n249352 );
not ( n249354 , n249353 );
or ( n249355 , n249344 , n249354 );
or ( n249356 , n249353 , n249343 );
nand ( n249357 , n249355 , n249356 );
not ( n249358 , n249357 );
not ( n249359 , n249358 );
or ( n249360 , n249333 , n249359 );
nand ( n249361 , n249331 , n249357 );
nand ( n249362 , n249360 , n249361 );
buf ( n249363 , n249362 );
and ( n249364 , n249303 , n249363 );
not ( n249365 , n249303 );
not ( n249366 , n249363 );
and ( n249367 , n249365 , n249366 );
nor ( n249368 , n249364 , n249367 );
not ( n249369 , n249368 );
xor ( n249370 , n37761 , n205215 );
xnor ( n249371 , n249370 , n39532 );
not ( n249372 , n243137 );
nand ( n249373 , n249371 , n249372 );
not ( n249374 , n249373 );
not ( n249375 , n248649 );
and ( n249376 , n249374 , n249375 );
and ( n249377 , n249373 , n248649 );
nor ( n249378 , n249376 , n249377 );
not ( n249379 , n249378 );
not ( n249380 , n249379 );
not ( n249381 , n243197 );
not ( n249382 , n249381 );
or ( n249383 , n249380 , n249382 );
not ( n249384 , n249379 );
and ( n249385 , n243192 , n243083 );
not ( n249386 , n243192 );
and ( n249387 , n249386 , n243084 );
nor ( n249388 , n249385 , n249387 );
nand ( n249389 , n249384 , n249388 );
nand ( n249390 , n249383 , n249389 );
and ( n249391 , n248961 , n248965 );
not ( n249392 , n248961 );
and ( n249393 , n249392 , n248931 );
nor ( n249394 , n249391 , n249393 );
buf ( n249395 , n249394 );
and ( n249396 , n249390 , n249395 );
not ( n249397 , n249390 );
buf ( n249398 , n248967 );
and ( n249399 , n249397 , n249398 );
nor ( n249400 , n249396 , n249399 );
nand ( n249401 , n249369 , n249400 );
or ( n249402 , n249289 , n249401 );
not ( n249403 , n249287 );
not ( n249404 , n249400 );
or ( n249405 , n249403 , n249404 );
nor ( n249406 , n249369 , n49051 );
nand ( n249407 , n249405 , n249406 );
nand ( n249408 , n233501 , n45284 );
nand ( n249409 , n249402 , n249407 , n249408 );
buf ( n249410 , n249409 );
not ( n249411 , n44205 );
not ( n249412 , n234097 );
or ( n249413 , n249411 , n249412 );
not ( n249414 , n44205 );
nand ( n249415 , n249414 , n234106 );
nand ( n249416 , n249413 , n249415 );
not ( n249417 , n38261 );
nand ( n249418 , n249417 , n226690 );
xor ( n249419 , n249418 , n234487 );
not ( n249420 , n249419 );
not ( n249421 , n38313 );
nand ( n249422 , n249421 , n48911 );
and ( n249423 , n249422 , n38358 );
not ( n249424 , n249422 );
and ( n249425 , n249424 , n234494 );
nor ( n249426 , n249423 , n249425 );
not ( n249427 , n249426 );
or ( n249428 , n249420 , n249427 );
or ( n249429 , n249426 , n249419 );
nand ( n249430 , n249428 , n249429 );
not ( n249431 , n249430 );
not ( n249432 , n249431 );
not ( n249433 , n49075 );
or ( n249434 , n249432 , n249433 );
nand ( n249435 , n226835 , n249430 );
nand ( n249436 , n249434 , n249435 );
not ( n249437 , n216261 );
nand ( n249438 , n249437 , n48998 );
not ( n249439 , n249438 );
not ( n249440 , n38511 );
not ( n249441 , n249440 );
and ( n249442 , n249439 , n249441 );
not ( n249443 , n216261 );
nand ( n249444 , n249443 , n48998 );
and ( n249445 , n249444 , n249440 );
nor ( n249446 , n249442 , n249445 );
not ( n249447 , n249446 );
not ( n249448 , n234114 );
nand ( n249449 , n38609 , n49029 );
not ( n249450 , n249449 );
or ( n249451 , n249448 , n249450 );
or ( n249452 , n249449 , n234114 );
nand ( n249453 , n249451 , n249452 );
not ( n249454 , n249453 );
and ( n249455 , n249447 , n249454 );
and ( n249456 , n249446 , n249453 );
nor ( n249457 , n249455 , n249456 );
and ( n249458 , n249436 , n249457 );
not ( n249459 , n249436 );
not ( n249460 , n249457 );
and ( n249461 , n249459 , n249460 );
nor ( n249462 , n249458 , n249461 );
buf ( n249463 , n249462 );
and ( n249464 , n249416 , n249463 );
not ( n249465 , n249416 );
and ( n249466 , n249436 , n249460 );
not ( n249467 , n249436 );
and ( n249468 , n249467 , n249457 );
nor ( n249469 , n249466 , n249468 );
buf ( n249470 , n249469 );
and ( n249471 , n249465 , n249470 );
nor ( n249472 , n249464 , n249471 );
nand ( n249473 , n249472 , n247444 );
not ( n249474 , n249473 );
not ( n249475 , n45827 );
not ( n249476 , n36729 );
or ( n249477 , n249475 , n249476 );
not ( n249478 , n45827 );
and ( n249479 , n36566 , n36727 );
not ( n249480 , n36566 );
and ( n249481 , n249480 , n36724 );
nor ( n249482 , n249479 , n249481 );
nand ( n249483 , n249478 , n249482 );
nand ( n249484 , n249477 , n249483 );
not ( n249485 , n247917 );
not ( n249486 , n247930 );
and ( n249487 , n249485 , n249486 );
and ( n249488 , n247917 , n247930 );
nor ( n249489 , n249487 , n249488 );
buf ( n249490 , n249489 );
not ( n249491 , n249490 );
and ( n249492 , n249484 , n249491 );
not ( n249493 , n249484 );
not ( n249494 , n249489 );
not ( n249495 , n249494 );
and ( n249496 , n249493 , n249495 );
nor ( n249497 , n249492 , n249496 );
not ( n249498 , n249497 );
not ( n249499 , n229086 );
not ( n249500 , n43005 );
or ( n249501 , n249499 , n249500 );
not ( n249502 , n229086 );
nand ( n249503 , n249502 , n43010 );
nand ( n249504 , n249501 , n249503 );
and ( n249505 , n249504 , n50028 );
not ( n249506 , n249504 );
and ( n249507 , n249506 , n227796 );
nor ( n249508 , n249505 , n249507 );
nand ( n249509 , n249474 , n249498 , n249508 );
nand ( n249510 , n249508 , n249472 );
nand ( n249511 , n249510 , n249497 , n249288 );
nand ( n249512 , n35431 , n30836 );
nand ( n249513 , n249509 , n249511 , n249512 );
buf ( n249514 , n249513 );
not ( n249515 , n234643 );
not ( n249516 , n249284 );
or ( n249517 , n249515 , n249516 );
not ( n249518 , n234643 );
and ( n249519 , n249269 , n249242 );
not ( n249520 , n249269 );
and ( n249521 , n249520 , n249243 );
nor ( n249522 , n249519 , n249521 );
nand ( n249523 , n249518 , n249522 );
nand ( n249524 , n249517 , n249523 );
buf ( n249525 , n242675 );
and ( n249526 , n249524 , n249525 );
not ( n249527 , n249524 );
buf ( n249528 , n242674 );
and ( n249529 , n249527 , n249528 );
nor ( n249530 , n249526 , n249529 );
buf ( n249531 , n226003 );
nor ( n249532 , n249530 , n249531 );
not ( n249533 , n249532 );
nand ( n249534 , n238437 , n51142 );
not ( n249535 , n249534 );
not ( n249536 , n235677 );
and ( n249537 , n249535 , n249536 );
and ( n249538 , n249534 , n235677 );
nor ( n249539 , n249537 , n249538 );
not ( n249540 , n249539 );
not ( n249541 , n241179 );
not ( n249542 , n249541 );
or ( n249543 , n249540 , n249542 );
or ( n249544 , n249541 , n249539 );
nand ( n249545 , n249543 , n249544 );
buf ( n249546 , n246553 );
and ( n249547 , n249545 , n249546 );
not ( n249548 , n249545 );
buf ( n249549 , n246548 );
and ( n249550 , n249548 , n249549 );
nor ( n249551 , n249547 , n249550 );
not ( n249552 , n39648 );
not ( n249553 , n35409 );
or ( n249554 , n249552 , n249553 );
not ( n249555 , n39648 );
nand ( n249556 , n249555 , n35417 );
nand ( n249557 , n249554 , n249556 );
nand ( n249558 , n46364 , n243645 );
not ( n249559 , n249558 );
not ( n249560 , n46353 );
and ( n249561 , n249559 , n249560 );
and ( n249562 , n249558 , n46353 );
nor ( n249563 , n249561 , n249562 );
not ( n249564 , n249563 );
not ( n249565 , n249564 );
not ( n249566 , n242998 );
not ( n249567 , n249566 );
or ( n249568 , n249565 , n249567 );
nand ( n249569 , n242998 , n249563 );
nand ( n249570 , n249568 , n249569 );
nand ( n249571 , n243559 , n46278 );
and ( n249572 , n249571 , n46289 );
not ( n249573 , n249571 );
and ( n249574 , n249573 , n248506 );
nor ( n249575 , n249572 , n249574 );
not ( n249576 , n249575 );
not ( n249577 , n249576 );
nand ( n249578 , n243529 , n46244 );
not ( n249579 , n249578 );
not ( n249580 , n248496 );
and ( n249581 , n249579 , n249580 );
and ( n249582 , n249578 , n248496 );
nor ( n249583 , n249581 , n249582 );
not ( n249584 , n249583 );
not ( n249585 , n249584 );
or ( n249586 , n249577 , n249585 );
nand ( n249587 , n249575 , n249583 );
nand ( n249588 , n249586 , n249587 );
nand ( n249589 , n46318 , n243595 );
not ( n249590 , n249589 );
not ( n249591 , n224068 );
and ( n249592 , n249590 , n249591 );
and ( n249593 , n249589 , n224068 );
nor ( n249594 , n249592 , n249593 );
and ( n249595 , n249588 , n249594 );
not ( n249596 , n249588 );
not ( n249597 , n249594 );
and ( n249598 , n249596 , n249597 );
nor ( n249599 , n249595 , n249598 );
xor ( n249600 , n249570 , n249599 );
buf ( n249601 , n249600 );
and ( n249602 , n249557 , n249601 );
not ( n249603 , n249557 );
not ( n249604 , n249599 );
not ( n249605 , n249604 );
not ( n249606 , n249570 );
not ( n249607 , n249606 );
or ( n249608 , n249605 , n249607 );
nand ( n249609 , n249599 , n249570 );
nand ( n249610 , n249608 , n249609 );
buf ( n249611 , n249610 );
and ( n249612 , n249603 , n249611 );
nor ( n249613 , n249602 , n249612 );
nand ( n249614 , n249551 , n249613 );
or ( n249615 , n249533 , n249614 );
not ( n249616 , n249551 );
not ( n249617 , n249530 );
not ( n249618 , n249617 );
or ( n249619 , n249616 , n249618 );
nor ( n249620 , n249613 , n238900 );
nand ( n249621 , n249619 , n249620 );
buf ( n249622 , n35431 );
nand ( n249623 , n249622 , n38056 );
nand ( n249624 , n249615 , n249621 , n249623 );
buf ( n249625 , n249624 );
not ( n249626 , RI19acb648_2244);
or ( n249627 , n25328 , n249626 );
not ( n249628 , RI19ac25e8_2311);
or ( n249629 , n25335 , n249628 );
nand ( n249630 , n249627 , n249629 );
buf ( n249631 , n249630 );
not ( n249632 , n246696 );
nand ( n249633 , n249632 , n235051 );
nand ( n249634 , n239582 , n239592 );
not ( n249635 , n249634 );
not ( n249636 , n246258 );
and ( n249637 , n249635 , n249636 );
and ( n249638 , n249634 , n246258 );
nor ( n249639 , n249637 , n249638 );
not ( n249640 , n249639 );
not ( n249641 , n249640 );
not ( n249642 , n248350 );
nand ( n249643 , n249642 , n239557 );
not ( n249644 , n249643 );
not ( n249645 , n244095 );
and ( n249646 , n249644 , n249645 );
and ( n249647 , n249643 , n244095 );
nor ( n249648 , n249646 , n249647 );
not ( n249649 , n249648 );
not ( n249650 , n248367 );
nand ( n249651 , n249650 , n239519 );
and ( n249652 , n249651 , n246295 );
not ( n249653 , n249651 );
and ( n249654 , n249653 , n246296 );
nor ( n249655 , n249652 , n249654 );
not ( n249656 , n249655 );
or ( n249657 , n249649 , n249656 );
or ( n249658 , n249655 , n249648 );
nand ( n249659 , n249657 , n249658 );
not ( n249660 , n246258 );
nand ( n249661 , n249660 , n239595 );
and ( n249662 , n249661 , n246247 );
not ( n249663 , n249661 );
and ( n249664 , n249663 , n246307 );
nor ( n249665 , n249662 , n249664 );
xnor ( n249666 , n249659 , n249665 );
nand ( n249667 , n248305 , n239480 );
not ( n249668 , n249667 );
not ( n249669 , n246269 );
or ( n249670 , n249668 , n249669 );
or ( n249671 , n246269 , n249667 );
nand ( n249672 , n249670 , n249671 );
not ( n249673 , n249672 );
not ( n249674 , n249673 );
nand ( n249675 , n239435 , n248326 );
and ( n249676 , n249675 , n239408 );
not ( n249677 , n249675 );
and ( n249678 , n249677 , n239407 );
nor ( n249679 , n249676 , n249678 );
not ( n249680 , n249679 );
not ( n249681 , n249680 );
or ( n249682 , n249674 , n249681 );
nand ( n249683 , n249679 , n249672 );
nand ( n249684 , n249682 , n249683 );
and ( n249685 , n249666 , n249684 );
not ( n249686 , n249666 );
not ( n249687 , n249684 );
and ( n249688 , n249686 , n249687 );
nor ( n249689 , n249685 , n249688 );
not ( n249690 , n249689 );
or ( n249691 , n249641 , n249690 );
not ( n249692 , n249640 );
not ( n249693 , n249689 );
nand ( n249694 , n249692 , n249693 );
nand ( n249695 , n249691 , n249694 );
not ( n249696 , n51434 );
nand ( n249697 , n35942 , n36080 );
not ( n249698 , n249697 );
or ( n249699 , n249696 , n249698 );
or ( n249700 , n249697 , n51434 );
nand ( n249701 , n249699 , n249700 );
not ( n249702 , n249701 );
nand ( n249703 , n36027 , n239639 );
not ( n249704 , n249703 );
not ( n249705 , n51406 );
and ( n249706 , n249704 , n249705 );
not ( n249707 , n35957 );
nand ( n249708 , n249707 , n36027 );
and ( n249709 , n249708 , n51406 );
nor ( n249710 , n249706 , n249709 );
not ( n249711 , n249710 );
or ( n249712 , n249702 , n249711 );
or ( n249713 , n249710 , n249701 );
nand ( n249714 , n249712 , n249713 );
nand ( n249715 , n237739 , n36115 );
not ( n249716 , n249715 );
not ( n249717 , n51460 );
and ( n249718 , n249716 , n249717 );
and ( n249719 , n249715 , n51460 );
nor ( n249720 , n249718 , n249719 );
and ( n249721 , n249714 , n249720 );
not ( n249722 , n249714 );
not ( n249723 , n249720 );
and ( n249724 , n249722 , n249723 );
nor ( n249725 , n249721 , n249724 );
not ( n249726 , n249725 );
not ( n249727 , n249726 );
not ( n249728 , n51511 );
nand ( n249729 , n239628 , n36354 );
not ( n249730 , n249729 );
or ( n249731 , n249728 , n249730 );
not ( n249732 , n36355 );
nand ( n249733 , n249732 , n239628 );
or ( n249734 , n249733 , n51511 );
nand ( n249735 , n249731 , n249734 );
not ( n249736 , n36194 );
nand ( n249737 , n249736 , n36249 );
not ( n249738 , n249737 );
buf ( n249739 , n51482 );
not ( n249740 , n249739 );
and ( n249741 , n249738 , n249740 );
and ( n249742 , n249737 , n249739 );
nor ( n249743 , n249741 , n249742 );
xor ( n249744 , n249735 , n249743 );
not ( n249745 , n249744 );
or ( n249746 , n249727 , n249745 );
not ( n249747 , n249744 );
nand ( n249748 , n249747 , n249725 );
nand ( n249749 , n249746 , n249748 );
buf ( n249750 , n249749 );
and ( n249751 , n249695 , n249750 );
not ( n249752 , n249695 );
not ( n249753 , n249747 );
not ( n249754 , n249725 );
and ( n249755 , n249753 , n249754 );
and ( n249756 , n249747 , n249725 );
nor ( n249757 , n249755 , n249756 );
not ( n249758 , n249757 );
not ( n249759 , n249758 );
and ( n249760 , n249752 , n249759 );
nor ( n249761 , n249751 , n249760 );
not ( n249762 , n249761 );
not ( n249763 , n38379 );
not ( n249764 , n234513 );
or ( n249765 , n249763 , n249764 );
not ( n249766 , n38379 );
nand ( n249767 , n249766 , n234521 );
nand ( n249768 , n249765 , n249767 );
and ( n249769 , n249768 , n45507 );
not ( n249770 , n249768 );
and ( n249771 , n249770 , n243431 );
nor ( n249772 , n249769 , n249771 );
nand ( n249773 , n249762 , n249772 );
or ( n249774 , n249633 , n249773 );
not ( n249775 , n249772 );
not ( n249776 , n249632 );
or ( n249777 , n249775 , n249776 );
nor ( n249778 , n249762 , n37725 );
nand ( n249779 , n249777 , n249778 );
nand ( n249780 , n237361 , n37869 );
nand ( n249781 , n249774 , n249779 , n249780 );
buf ( n249782 , n249781 );
buf ( n249783 , n43141 );
not ( n249784 , n249783 );
not ( n249785 , n244453 );
or ( n249786 , n249784 , n249785 );
or ( n249787 , n244453 , n249783 );
nand ( n249788 , n249786 , n249787 );
not ( n249789 , n244460 );
and ( n249790 , n249788 , n249789 );
not ( n249791 , n249788 );
not ( n249792 , n244459 );
and ( n249793 , n249791 , n249792 );
nor ( n249794 , n249790 , n249793 );
nor ( n249795 , n249794 , n247698 );
not ( n249796 , n249795 );
not ( n249797 , n242148 );
not ( n249798 , n246936 );
not ( n249799 , n249798 );
nand ( n249800 , n246953 , n208535 );
and ( n249801 , n249800 , n29993 );
not ( n249802 , n249800 );
and ( n249803 , n249802 , n29992 );
nor ( n249804 , n249801 , n249803 );
not ( n249805 , n249804 );
not ( n249806 , n249805 );
not ( n249807 , n229472 );
nand ( n249808 , n30811 , n249807 );
and ( n249809 , n249808 , n229463 );
not ( n249810 , n249808 );
not ( n249811 , n229463 );
and ( n249812 , n249810 , n249811 );
nor ( n249813 , n249809 , n249812 );
not ( n249814 , n249813 );
not ( n249815 , n249814 );
or ( n249816 , n249806 , n249815 );
nand ( n249817 , n249813 , n249804 );
nand ( n249818 , n249816 , n249817 );
not ( n249819 , n249818 );
nor ( n249820 , n229422 , n207903 );
not ( n249821 , n249820 );
not ( n249822 , n51652 );
or ( n249823 , n249821 , n249822 );
not ( n249824 , n249820 );
not ( n249825 , n51652 );
nand ( n249826 , n249824 , n249825 );
nand ( n249827 , n249823 , n249826 );
xor ( n249828 , n229391 , n249827 );
nand ( n249829 , n30697 , n51687 );
not ( n249830 , n249829 );
not ( n249831 , n229437 );
and ( n249832 , n249830 , n249831 );
and ( n249833 , n249829 , n229437 );
nor ( n249834 , n249832 , n249833 );
xor ( n249835 , n249828 , n249834 );
not ( n249836 , n249835 );
not ( n249837 , n249836 );
or ( n249838 , n249819 , n249837 );
not ( n249839 , n249818 );
nand ( n249840 , n249835 , n249839 );
nand ( n249841 , n249838 , n249840 );
not ( n249842 , n249841 );
or ( n249843 , n249799 , n249842 );
or ( n249844 , n249841 , n249798 );
nand ( n249845 , n249843 , n249844 );
not ( n249846 , n249845 );
or ( n249847 , n249797 , n249846 );
not ( n249848 , n242148 );
not ( n249849 , n249848 );
or ( n249850 , n249845 , n249849 );
nand ( n249851 , n249847 , n249850 );
buf ( n249852 , n240956 );
not ( n249853 , n249852 );
not ( n249854 , n54105 );
not ( n249855 , n231893 );
or ( n249856 , n249854 , n249855 );
nand ( n249857 , n54129 , n54106 );
nand ( n249858 , n249856 , n249857 );
not ( n249859 , n249858 );
or ( n249860 , n249853 , n249859 );
or ( n249861 , n249858 , n249852 );
nand ( n249862 , n249860 , n249861 );
not ( n249863 , n249862 );
not ( n249864 , n54192 );
and ( n249865 , n249863 , n249864 );
and ( n249866 , n249862 , n231957 );
nor ( n249867 , n249865 , n249866 );
or ( n249868 , n249851 , n249867 );
or ( n249869 , n249796 , n249868 );
not ( n249870 , n249794 );
nor ( n249871 , n249870 , n247698 );
nand ( n249872 , n249871 , n249868 );
nand ( n249873 , n247423 , n37187 );
nand ( n249874 , n249869 , n249872 , n249873 );
buf ( n249875 , n249874 );
not ( n249876 , n49931 );
nand ( n249877 , n249876 , n39419 );
not ( n249878 , n249877 );
not ( n249879 , n245825 );
and ( n249880 , n249878 , n249879 );
and ( n249881 , n249877 , n245825 );
nor ( n249882 , n249880 , n249881 );
not ( n249883 , n249882 );
not ( n249884 , n249883 );
not ( n249885 , n49903 );
nand ( n249886 , n249885 , n39330 );
not ( n249887 , n249886 );
not ( n249888 , n49892 );
and ( n249889 , n249887 , n249888 );
and ( n249890 , n249886 , n49892 );
nor ( n249891 , n249889 , n249890 );
not ( n249892 , n249891 );
or ( n249893 , n249884 , n249892 );
not ( n249894 , n249891 );
nand ( n249895 , n249894 , n249882 );
nand ( n249896 , n249893 , n249895 );
not ( n249897 , n245846 );
not ( n249898 , n39116 );
not ( n249899 , n227577 );
nand ( n249900 , n249898 , n249899 );
not ( n249901 , n249900 );
or ( n249902 , n249897 , n249901 );
not ( n249903 , n227577 );
nand ( n249904 , n249903 , n249898 );
or ( n249905 , n249904 , n245846 );
nand ( n249906 , n249902 , n249905 );
not ( n249907 , n249906 );
nand ( n249908 , n227595 , n39253 );
not ( n249909 , n249908 );
not ( n249910 , n227611 );
not ( n249911 , n249910 );
and ( n249912 , n249909 , n249911 );
and ( n249913 , n249908 , n249910 );
nor ( n249914 , n249912 , n249913 );
not ( n249915 , n249914 );
or ( n249916 , n249907 , n249915 );
or ( n249917 , n249914 , n249906 );
nand ( n249918 , n249916 , n249917 );
and ( n249919 , n249918 , n242905 );
not ( n249920 , n249918 );
and ( n249921 , n249920 , n242906 );
nor ( n249922 , n249919 , n249921 );
not ( n249923 , n249922 );
and ( n249924 , n249896 , n249923 );
not ( n249925 , n249896 );
and ( n249926 , n249925 , n249922 );
nor ( n249927 , n249924 , n249926 );
not ( n249928 , n249927 );
not ( n249929 , n249928 );
not ( n249930 , n249929 );
nand ( n249931 , n38810 , n38777 );
not ( n249932 , n249931 );
not ( n249933 , n49668 );
and ( n249934 , n249932 , n249933 );
and ( n249935 , n249931 , n49668 );
nor ( n249936 , n249934 , n249935 );
buf ( n249937 , n249936 );
not ( n249938 , n249937 );
not ( n249939 , n242569 );
not ( n249940 , n249939 );
or ( n249941 , n249938 , n249940 );
or ( n249942 , n242574 , n249937 );
nand ( n249943 , n249941 , n249942 );
not ( n249944 , n249943 );
and ( n249945 , n249930 , n249944 );
and ( n249946 , n249929 , n249943 );
nor ( n249947 , n249945 , n249946 );
not ( n249948 , n249947 );
not ( n249949 , n249948 );
not ( n249950 , n54729 );
not ( n249951 , n249950 );
not ( n249952 , n245517 );
or ( n249953 , n249951 , n249952 );
or ( n249954 , n245517 , n249950 );
nand ( n249955 , n249953 , n249954 );
and ( n249956 , n245474 , n249955 );
not ( n249957 , n245474 );
not ( n249958 , n249955 );
and ( n249959 , n249957 , n249958 );
nor ( n249960 , n249956 , n249959 );
not ( n249961 , n249960 );
or ( n249962 , n249949 , n249961 );
not ( n249963 , n245334 );
not ( n249964 , n241281 );
and ( n249965 , n249963 , n249964 );
and ( n249966 , n245334 , n241281 );
nor ( n249967 , n249965 , n249966 );
and ( n249968 , n249967 , n245393 );
not ( n249969 , n249967 );
and ( n249970 , n249969 , n245403 );
nor ( n249971 , n249968 , n249970 );
not ( n249972 , n249971 );
nor ( n249973 , n249972 , n55104 );
nand ( n249974 , n249962 , n249973 );
nor ( n249975 , n249947 , n43517 );
nand ( n249976 , n249975 , n249972 , n249960 );
nand ( n249977 , n241068 , n32074 );
nand ( n249978 , n249974 , n249976 , n249977 );
buf ( n249979 , n249978 );
not ( n249980 , n47601 );
not ( n249981 , n51381 );
or ( n249982 , n249980 , n249981 );
not ( n249983 , n235298 );
not ( n249984 , n246448 );
or ( n249985 , n249983 , n249984 );
not ( n249986 , n235298 );
nand ( n249987 , n249986 , n246439 );
nand ( n249988 , n249985 , n249987 );
not ( n249989 , n46927 );
nand ( n249990 , n249989 , n224659 );
not ( n249991 , n249990 );
not ( n249992 , n237850 );
and ( n249993 , n249991 , n249992 );
and ( n249994 , n249990 , n237850 );
nor ( n249995 , n249993 , n249994 );
not ( n249996 , n249995 );
not ( n249997 , n249996 );
not ( n249998 , n245229 );
not ( n249999 , n249998 );
or ( n250000 , n249997 , n249999 );
nand ( n250001 , n245229 , n249995 );
nand ( n250002 , n250000 , n250001 );
not ( n250003 , n247433 );
nand ( n250004 , n224626 , n46850 );
not ( n250005 , n250004 );
not ( n250006 , n50693 );
and ( n250007 , n250005 , n250006 );
and ( n250008 , n250004 , n50693 );
nor ( n250009 , n250007 , n250008 );
not ( n250010 , n250009 );
or ( n250011 , n250003 , n250010 );
or ( n250012 , n250009 , n247433 );
nand ( n250013 , n250011 , n250012 );
not ( n250014 , n228398 );
and ( n250015 , n250013 , n250014 );
not ( n250016 , n250013 );
and ( n250017 , n250016 , n228398 );
nor ( n250018 , n250015 , n250017 );
xor ( n250019 , n250002 , n250018 );
not ( n250020 , n250019 );
not ( n250021 , n250020 );
and ( n250022 , n249988 , n250021 );
not ( n250023 , n249988 );
not ( n250024 , n250018 );
and ( n250025 , n250002 , n250024 );
not ( n250026 , n250002 );
and ( n250027 , n250026 , n250018 );
nor ( n250028 , n250025 , n250027 );
not ( n250029 , n250028 );
not ( n250030 , n250029 );
and ( n250031 , n250023 , n250030 );
nor ( n250032 , n250022 , n250031 );
not ( n250033 , n250032 );
not ( n250034 , n236006 );
nand ( n250035 , n236009 , n50169 );
not ( n250036 , n250035 );
or ( n250037 , n250034 , n250036 );
nand ( n250038 , n236009 , n50169 );
or ( n250039 , n250038 , n236006 );
nand ( n250040 , n250037 , n250039 );
not ( n250041 , n250040 );
not ( n250042 , n236056 );
or ( n250043 , n250041 , n250042 );
not ( n250044 , n250040 );
nand ( n250045 , n250044 , n236063 );
nand ( n250046 , n250043 , n250045 );
and ( n250047 , n250046 , n236171 );
not ( n250048 , n250046 );
and ( n250049 , n250048 , n236167 );
nor ( n250050 , n250047 , n250049 );
not ( n250051 , n250050 );
nand ( n250052 , n250033 , n250051 );
not ( n250053 , n249426 );
not ( n250054 , n38633 );
or ( n250055 , n250053 , n250054 );
not ( n250056 , n249426 );
nand ( n250057 , n250056 , n38625 );
nand ( n250058 , n250055 , n250057 );
and ( n250059 , n250058 , n49182 );
not ( n250060 , n250058 );
and ( n250061 , n250060 , n49191 );
nor ( n250062 , n250059 , n250061 );
not ( n250063 , n250062 );
and ( n250064 , n250052 , n250063 );
not ( n250065 , n250052 );
and ( n250066 , n250065 , n250062 );
nor ( n250067 , n250064 , n250066 );
not ( n250068 , n234111 );
or ( n250069 , n250067 , n250068 );
nand ( n250070 , n249982 , n250069 );
buf ( n250071 , n250070 );
not ( n250072 , n248957 );
nand ( n250073 , n235983 , n227845 );
and ( n250074 , n250073 , n235985 );
not ( n250075 , n250073 );
and ( n250076 , n250075 , n227821 );
nor ( n250077 , n250074 , n250076 );
nand ( n250078 , n235970 , n50259 );
and ( n250079 , n250078 , n235960 );
not ( n250080 , n250078 );
not ( n250081 , n235960 );
and ( n250082 , n250080 , n250081 );
nor ( n250083 , n250079 , n250082 );
not ( n250084 , n250083 );
not ( n250085 , n250084 );
not ( n250086 , n235941 );
or ( n250087 , n250085 , n250086 );
nand ( n250088 , n235940 , n250083 );
nand ( n250089 , n250087 , n250088 );
xor ( n250090 , n250077 , n250089 );
not ( n250091 , n250040 );
nand ( n250092 , n236039 , n50126 );
xor ( n250093 , n250092 , n236028 );
not ( n250094 , n250093 );
and ( n250095 , n250091 , n250094 );
and ( n250096 , n250040 , n250093 );
nor ( n250097 , n250095 , n250096 );
xor ( n250098 , n250090 , n250097 );
not ( n250099 , n250098 );
not ( n250100 , n250099 );
or ( n250101 , n250072 , n250100 );
not ( n250102 , n250098 );
or ( n250103 , n250102 , n248957 );
nand ( n250104 , n250101 , n250103 );
buf ( n250105 , n238297 );
and ( n250106 , n250104 , n250105 );
not ( n250107 , n250104 );
buf ( n250108 , n238288 );
and ( n250109 , n250107 , n250108 );
nor ( n250110 , n250106 , n250109 );
not ( n250111 , n31571 );
nand ( n250112 , n250110 , n250111 );
not ( n250113 , n236886 );
not ( n250114 , n250113 );
not ( n250115 , n31089 );
not ( n250116 , n247018 );
or ( n250117 , n250115 , n250116 );
not ( n250118 , n31089 );
nand ( n250119 , n250118 , n247013 );
nand ( n250120 , n250117 , n250119 );
not ( n250121 , n250120 );
or ( n250122 , n250114 , n250121 );
not ( n250123 , n236886 );
or ( n250124 , n250120 , n250123 );
nand ( n250125 , n250122 , n250124 );
not ( n250126 , n250125 );
not ( n250127 , n243530 );
nand ( n250128 , n250127 , n248500 );
and ( n250129 , n250128 , n46244 );
not ( n250130 , n250128 );
and ( n250131 , n250130 , n46245 );
nor ( n250132 , n250129 , n250131 );
buf ( n250133 , n250132 );
not ( n250134 , n250133 );
not ( n250135 , n249600 );
or ( n250136 , n250134 , n250135 );
or ( n250137 , n249600 , n250133 );
nand ( n250138 , n250136 , n250137 );
not ( n250139 , n250138 );
not ( n250140 , n33986 );
buf ( n250141 , n216050 );
not ( n250142 , n250141 );
not ( n250143 , n30889 );
or ( n250144 , n250142 , n250143 );
or ( n250145 , n30889 , n250141 );
nand ( n250146 , n250144 , n250145 );
and ( n250147 , n250140 , n250146 );
not ( n250148 , n250140 );
not ( n250149 , n250146 );
and ( n250150 , n250148 , n250149 );
nor ( n250151 , n250147 , n250150 );
nand ( n250152 , n250151 , n243170 );
not ( n250153 , n250152 );
not ( n250154 , n243167 );
and ( n250155 , n250153 , n250154 );
and ( n250156 , n250152 , n243167 );
nor ( n250157 , n250155 , n250156 );
not ( n250158 , n250157 );
not ( n250159 , n205269 );
not ( n250160 , n31777 );
or ( n250161 , n250159 , n250160 );
not ( n250162 , n205269 );
nand ( n250163 , n250162 , n33684 );
nand ( n250164 , n250161 , n250163 );
and ( n250165 , n250164 , n221323 );
not ( n250166 , n250164 );
and ( n250167 , n250166 , n46656 );
nor ( n250168 , n250165 , n250167 );
nand ( n250169 , n250168 , n243091 );
and ( n250170 , n250169 , n243102 );
not ( n250171 , n250169 );
and ( n250172 , n250171 , n248621 );
nor ( n250173 , n250170 , n250172 );
not ( n250174 , n250173 );
or ( n250175 , n250158 , n250174 );
or ( n250176 , n250173 , n250157 );
nand ( n250177 , n250175 , n250176 );
and ( n250178 , n250177 , n249378 );
not ( n250179 , n250177 );
and ( n250180 , n250179 , n249379 );
nor ( n250181 , n250178 , n250180 );
buf ( n250182 , n212623 );
not ( n250183 , n250182 );
not ( n250184 , n34264 );
or ( n250185 , n250183 , n250184 );
not ( n250186 , n239577 );
or ( n250187 , n250186 , n250182 );
nand ( n250188 , n250185 , n250187 );
and ( n250189 , n250188 , n28188 );
not ( n250190 , n250188 );
and ( n250191 , n250190 , n41594 );
nor ( n250192 , n250189 , n250191 );
nand ( n250193 , n243017 , n250192 );
not ( n250194 , n250193 );
not ( n250195 , n243026 );
and ( n250196 , n250194 , n250195 );
and ( n250197 , n250193 , n243026 );
nor ( n250198 , n250196 , n250197 );
not ( n250199 , n250198 );
not ( n250200 , RI1749d1e8_970);
and ( n250201 , n35060 , n250200 );
not ( n250202 , n35060 );
and ( n250203 , n250202 , n35057 );
nor ( n250204 , n250201 , n250203 );
not ( n250205 , n250204 );
not ( n250206 , n204671 );
or ( n250207 , n250205 , n250206 );
not ( n250208 , n250204 );
nand ( n250209 , n238663 , n250208 );
nand ( n250210 , n250207 , n250209 );
and ( n250211 , n250210 , n26261 );
not ( n250212 , n250210 );
and ( n250213 , n250212 , n204681 );
nor ( n250214 , n250211 , n250213 );
not ( n250215 , n250214 );
nand ( n250216 , n243052 , n250215 );
and ( n250217 , n250216 , n243063 );
not ( n250218 , n250216 );
and ( n250219 , n250218 , n243062 );
nor ( n250220 , n250217 , n250219 );
not ( n250221 , n250220 );
or ( n250222 , n250199 , n250221 );
or ( n250223 , n250220 , n250198 );
nand ( n250224 , n250222 , n250223 );
and ( n250225 , n250181 , n250224 );
not ( n250226 , n250181 );
not ( n250227 , n250224 );
and ( n250228 , n250226 , n250227 );
nor ( n250229 , n250225 , n250228 );
not ( n250230 , n250229 );
not ( n250231 , n250230 );
not ( n250232 , n250231 );
and ( n250233 , n250139 , n250232 );
buf ( n250234 , n250229 );
and ( n250235 , n250234 , n250138 );
nor ( n250236 , n250233 , n250235 );
nand ( n250237 , n250126 , n250236 );
or ( n250238 , n250112 , n250237 );
not ( n250239 , n250126 );
not ( n250240 , n250110 );
or ( n250241 , n250239 , n250240 );
nor ( n250242 , n250236 , n37725 );
nand ( n250243 , n250241 , n250242 );
nand ( n250244 , n246217 , n28619 );
nand ( n250245 , n250238 , n250243 , n250244 );
buf ( n250246 , n250245 );
not ( n250247 , n245819 );
not ( n250248 , n39434 );
or ( n250249 , n250247 , n250248 );
not ( n250250 , n245819 );
nand ( n250251 , n250250 , n39444 );
nand ( n250252 , n250249 , n250251 );
and ( n250253 , n250252 , n248795 );
not ( n250254 , n250252 );
buf ( n250255 , n52989 );
and ( n250256 , n250254 , n250255 );
nor ( n250257 , n250253 , n250256 );
not ( n250258 , n250257 );
nor ( n250259 , n250258 , n238635 );
not ( n250260 , n246034 );
nand ( n250261 , n243865 , n222656 );
not ( n250262 , n250261 );
or ( n250263 , n250260 , n250262 );
or ( n250264 , n250261 , n246034 );
nand ( n250265 , n250263 , n250264 );
not ( n250266 , n250265 );
not ( n250267 , n243959 );
or ( n250268 , n250266 , n250267 );
not ( n250269 , n250265 );
nand ( n250270 , n250269 , n243953 );
nand ( n250271 , n250268 , n250270 );
buf ( n250272 , n237936 );
and ( n250273 , n250271 , n250272 );
not ( n250274 , n250271 );
buf ( n250275 , n237944 );
and ( n250276 , n250274 , n250275 );
nor ( n250277 , n250273 , n250276 );
nand ( n250278 , n250259 , n248286 , n250277 );
not ( n250279 , n250257 );
not ( n250280 , n248286 );
or ( n250281 , n250279 , n250280 );
nor ( n250282 , n250277 , n55146 );
nand ( n250283 , n250281 , n250282 );
nand ( n250284 , n236798 , n207477 );
nand ( n250285 , n250278 , n250283 , n250284 );
buf ( n250286 , n250285 );
not ( n250287 , RI19a9ad18_2606);
or ( n250288 , n226819 , n250287 );
not ( n250289 , RI19a90cc8_2677);
or ( n250290 , n25335 , n250289 );
nand ( n250291 , n250288 , n250290 );
buf ( n250292 , n250291 );
not ( n250293 , n47625 );
not ( n250294 , n238033 );
or ( n250295 , n250293 , n250294 );
not ( n250296 , n47625 );
nand ( n250297 , n250296 , n238040 );
nand ( n250298 , n250295 , n250297 );
and ( n250299 , n250298 , n238102 );
not ( n250300 , n250298 );
and ( n250301 , n250300 , n238107 );
nor ( n250302 , n250299 , n250301 );
nor ( n250303 , n250302 , n39763 );
not ( n250304 , n250303 );
not ( n250305 , n53402 );
not ( n250306 , n250305 );
not ( n250307 , n237021 );
not ( n250308 , n231097 );
nand ( n250309 , n250308 , n244669 );
not ( n250310 , n250309 );
buf ( n250311 , n237058 );
not ( n250312 , n250311 );
and ( n250313 , n250310 , n250312 );
and ( n250314 , n250309 , n250311 );
nor ( n250315 , n250313 , n250314 );
not ( n250316 , n250315 );
or ( n250317 , n250307 , n250316 );
or ( n250318 , n250315 , n237021 );
nand ( n250319 , n250317 , n250318 );
not ( n250320 , n53434 );
nand ( n250321 , n250320 , n241708 );
not ( n250322 , n250321 );
not ( n250323 , n237024 );
not ( n250324 , n250323 );
and ( n250325 , n250322 , n250324 );
and ( n250326 , n250321 , n250323 );
nor ( n250327 , n250325 , n250326 );
not ( n250328 , n250327 );
and ( n250329 , n250319 , n250328 );
not ( n250330 , n250319 );
and ( n250331 , n250330 , n250327 );
nor ( n250332 , n250329 , n250331 );
not ( n250333 , n53324 );
nand ( n250334 , n250333 , n244692 );
and ( n250335 , n250334 , n237114 );
not ( n250336 , n250334 );
not ( n250337 , n237114 );
and ( n250338 , n250336 , n250337 );
nor ( n250339 , n250335 , n250338 );
not ( n250340 , n250339 );
not ( n250341 , n250340 );
not ( n250342 , n53268 );
nand ( n250343 , n250342 , n244681 );
not ( n250344 , n250343 );
not ( n250345 , n237089 );
not ( n250346 , n250345 );
and ( n250347 , n250344 , n250346 );
and ( n250348 , n250343 , n250345 );
nor ( n250349 , n250347 , n250348 );
not ( n250350 , n250349 );
not ( n250351 , n250350 );
or ( n250352 , n250341 , n250351 );
nand ( n250353 , n250349 , n250339 );
nand ( n250354 , n250352 , n250353 );
not ( n250355 , n250354 );
and ( n250356 , n250332 , n250355 );
not ( n250357 , n250332 );
and ( n250358 , n250357 , n250354 );
nor ( n250359 , n250356 , n250358 );
not ( n250360 , n250359 );
or ( n250361 , n250306 , n250360 );
not ( n250362 , n250305 );
and ( n250363 , n250332 , n250354 );
not ( n250364 , n250332 );
and ( n250365 , n250364 , n250355 );
nor ( n250366 , n250363 , n250365 );
nand ( n250367 , n250362 , n250366 );
nand ( n250368 , n250361 , n250367 );
not ( n250369 , n248901 );
not ( n250370 , n250369 );
buf ( n250371 , n250370 );
and ( n250372 , n250368 , n250371 );
not ( n250373 , n250368 );
buf ( n250374 , n248892 );
and ( n250375 , n250373 , n250374 );
nor ( n250376 , n250372 , n250375 );
not ( n250377 , n250376 );
nand ( n250378 , n250377 , n45729 );
or ( n250379 , n250304 , n250378 );
not ( n250380 , n250302 );
not ( n250381 , n250380 );
not ( n250382 , n250377 );
or ( n250383 , n250381 , n250382 );
nor ( n250384 , n45729 , n54208 );
nand ( n250385 , n250383 , n250384 );
nand ( n250386 , n234024 , n45367 );
nand ( n250387 , n250379 , n250385 , n250386 );
buf ( n250388 , n250387 );
not ( n250389 , n244149 );
not ( n250390 , n234810 );
or ( n250391 , n250389 , n250390 );
not ( n250392 , n244149 );
nand ( n250393 , n250392 , n234803 );
nand ( n250394 , n250391 , n250393 );
buf ( n250395 , n244282 );
and ( n250396 , n250394 , n250395 );
not ( n250397 , n250394 );
buf ( n250398 , n244273 );
and ( n250399 , n250397 , n250398 );
nor ( n250400 , n250396 , n250399 );
nand ( n250401 , n250400 , n245241 );
not ( n250402 , n250339 );
not ( n250403 , n237135 );
or ( n250404 , n250402 , n250403 );
not ( n250405 , n250339 );
nand ( n250406 , n250405 , n237148 );
nand ( n250407 , n250404 , n250406 );
buf ( n250408 , n237340 );
and ( n250409 , n250407 , n250408 );
not ( n250410 , n250407 );
not ( n250411 , n237350 );
not ( n250412 , n250411 );
and ( n250413 , n250410 , n250412 );
nor ( n250414 , n250409 , n250413 );
not ( n250415 , n50465 );
not ( n250416 , n250415 );
not ( n250417 , n53811 );
or ( n250418 , n250416 , n250417 );
not ( n250419 , n250415 );
nand ( n250420 , n250419 , n53820 );
nand ( n250421 , n250418 , n250420 );
and ( n250422 , n250421 , n231776 );
not ( n250423 , n250421 );
and ( n250424 , n250423 , n231769 );
nor ( n250425 , n250422 , n250424 );
nand ( n250426 , n250414 , n250425 );
or ( n250427 , n250401 , n250426 );
not ( n250428 , n250400 );
not ( n250429 , n250414 );
or ( n250430 , n250428 , n250429 );
not ( n250431 , n226010 );
nor ( n250432 , n250425 , n250431 );
nand ( n250433 , n250430 , n250432 );
nand ( n250434 , n41945 , n31895 );
nand ( n250435 , n250427 , n250433 , n250434 );
buf ( n250436 , n250435 );
buf ( n250437 , n245431 );
not ( n250438 , n250437 );
not ( n250439 , n241962 );
not ( n250440 , n250439 );
or ( n250441 , n250438 , n250440 );
not ( n250442 , n241962 );
or ( n250443 , n250442 , n250437 );
nand ( n250444 , n250441 , n250443 );
not ( n250445 , n250444 );
not ( n250446 , n234596 );
nand ( n250447 , n231335 , n236810 );
not ( n250448 , n250447 );
or ( n250449 , n250446 , n250448 );
not ( n250450 , n234597 );
or ( n250451 , n250447 , n250450 );
nand ( n250452 , n250449 , n250451 );
not ( n250453 , n250452 );
not ( n250454 , n250453 );
not ( n250455 , n53541 );
nand ( n250456 , n250455 , n244855 );
not ( n250457 , n250456 );
not ( n250458 , n234580 );
and ( n250459 , n250457 , n250458 );
and ( n250460 , n250456 , n234580 );
nor ( n250461 , n250459 , n250460 );
not ( n250462 , n250461 );
not ( n250463 , n250462 );
or ( n250464 , n250454 , n250463 );
nand ( n250465 , n250452 , n250461 );
nand ( n250466 , n250464 , n250465 );
nand ( n250467 , n53490 , n231245 );
and ( n250468 , n250467 , n234620 );
not ( n250469 , n250467 );
and ( n250470 , n250469 , n234619 );
nor ( n250471 , n250468 , n250470 );
and ( n250472 , n250466 , n250471 );
not ( n250473 , n250466 );
not ( n250474 , n250471 );
and ( n250475 , n250473 , n250474 );
nor ( n250476 , n250472 , n250475 );
not ( n250477 , n250476 );
not ( n250478 , n249224 );
not ( n250479 , n53620 );
nand ( n250480 , n250479 , n244871 );
not ( n250481 , n250480 );
or ( n250482 , n250478 , n250481 );
or ( n250483 , n250480 , n249224 );
nand ( n250484 , n250482 , n250483 );
not ( n250485 , n250484 );
not ( n250486 , n250485 );
not ( n250487 , n234556 );
not ( n250488 , n250487 );
or ( n250489 , n250486 , n250488 );
nand ( n250490 , n234556 , n250484 );
nand ( n250491 , n250489 , n250490 );
not ( n250492 , n250491 );
not ( n250493 , n250492 );
and ( n250494 , n250477 , n250493 );
and ( n250495 , n250476 , n250492 );
nor ( n250496 , n250494 , n250495 );
not ( n250497 , n250496 );
not ( n250498 , n250497 );
not ( n250499 , n250498 );
and ( n250500 , n250445 , n250499 );
buf ( n250501 , n250496 );
and ( n250502 , n250444 , n250501 );
nor ( n250503 , n250500 , n250502 );
nor ( n250504 , n250503 , n52445 );
not ( n250505 , n250504 );
not ( n250506 , n48749 );
not ( n250507 , n239220 );
or ( n250508 , n250506 , n250507 );
not ( n250509 , n48749 );
nand ( n250510 , n250509 , n239228 );
nand ( n250511 , n250508 , n250510 );
not ( n250512 , n49370 );
not ( n250513 , n34913 );
not ( n250514 , n31044 );
and ( n250515 , n250513 , n250514 );
and ( n250516 , n34913 , n31044 );
nor ( n250517 , n250515 , n250516 );
and ( n250518 , n250517 , n223614 );
not ( n250519 , n250517 );
and ( n250520 , n250519 , n45850 );
nor ( n250521 , n250518 , n250520 );
nand ( n250522 , n227145 , n250521 );
not ( n250523 , n250522 );
or ( n250524 , n250512 , n250523 );
or ( n250525 , n250522 , n49370 );
nand ( n250526 , n250524 , n250525 );
not ( n250527 , n250526 );
and ( n250528 , n33411 , n39844 );
not ( n250529 , n33411 );
and ( n250530 , n250529 , n41797 );
nor ( n250531 , n250528 , n250530 );
not ( n250532 , n250531 );
not ( n250533 , n250532 );
not ( n250534 , n32362 );
or ( n250535 , n250533 , n250534 );
nand ( n250536 , n227439 , n250531 );
nand ( n250537 , n250535 , n250536 );
nand ( n250538 , n49331 , n250537 );
not ( n250539 , n250538 );
not ( n250540 , n227081 );
and ( n250541 , n250539 , n250540 );
and ( n250542 , n250538 , n227081 );
nor ( n250543 , n250541 , n250542 );
not ( n250544 , n250543 );
or ( n250545 , n250527 , n250544 );
or ( n250546 , n250543 , n250526 );
nand ( n250547 , n250545 , n250546 );
and ( n250548 , n250547 , n249085 );
not ( n250549 , n250547 );
and ( n250550 , n250549 , n249084 );
nor ( n250551 , n250548 , n250550 );
not ( n250552 , n250551 );
not ( n250553 , n227005 );
not ( n250554 , n31771 );
not ( n250555 , n44333 );
or ( n250556 , n250554 , n250555 );
nand ( n250557 , n227881 , n209528 );
nand ( n250558 , n250556 , n250557 );
xor ( n250559 , n250558 , n239578 );
not ( n250560 , n250559 );
nand ( n250561 , n227008 , n250560 );
not ( n250562 , n250561 );
or ( n250563 , n250553 , n250562 );
nand ( n250564 , n227008 , n250560 );
or ( n250565 , n250564 , n227005 );
nand ( n250566 , n250563 , n250565 );
not ( n250567 , n250566 );
not ( n250568 , n226983 );
and ( n250569 , n250567 , n250568 );
and ( n250570 , n250566 , n226983 );
nor ( n250571 , n250569 , n250570 );
not ( n250572 , n250571 );
or ( n250573 , n250552 , n250572 );
or ( n250574 , n250571 , n250551 );
nand ( n250575 , n250573 , n250574 );
buf ( n250576 , n250575 );
not ( n250577 , n250576 );
and ( n250578 , n250511 , n250577 );
not ( n250579 , n250511 );
buf ( n250580 , n250576 );
and ( n250581 , n250579 , n250580 );
nor ( n250582 , n250578 , n250581 );
not ( n250583 , n42543 );
not ( n250584 , n237639 );
or ( n250585 , n250583 , n250584 );
not ( n250586 , n42543 );
nand ( n250587 , n250586 , n237647 );
nand ( n250588 , n250585 , n250587 );
and ( n250589 , n250588 , n237704 );
not ( n250590 , n250588 );
and ( n250591 , n250590 , n241677 );
nor ( n250592 , n250589 , n250591 );
not ( n250593 , n250592 );
nand ( n250594 , n250582 , n250593 );
or ( n250595 , n250505 , n250594 );
not ( n250596 , n250582 );
not ( n250597 , n250503 );
not ( n250598 , n250597 );
or ( n250599 , n250596 , n250598 );
nor ( n250600 , n250593 , n226003 );
nand ( n250601 , n250599 , n250600 );
nand ( n250602 , n51381 , n35377 );
nand ( n250603 , n250595 , n250601 , n250602 );
buf ( n250604 , n250603 );
not ( n250605 , n247312 );
not ( n250606 , n246171 );
or ( n250607 , n250605 , n250606 );
not ( n250608 , n247312 );
nand ( n250609 , n250608 , n246166 );
nand ( n250610 , n250607 , n250609 );
not ( n250611 , n37594 );
not ( n250612 , n31290 );
not ( n250613 , n28117 );
or ( n250614 , n250612 , n250613 );
nand ( n250615 , n205877 , n209047 );
nand ( n250616 , n250614 , n250615 );
not ( n250617 , n250616 );
not ( n250618 , n28106 );
not ( n250619 , n250618 );
or ( n250620 , n250617 , n250619 );
or ( n250621 , n250618 , n250616 );
nand ( n250622 , n250620 , n250621 );
and ( n250623 , n250622 , n51033 );
not ( n250624 , n250622 );
and ( n250625 , n250624 , n44988 );
nor ( n250626 , n250623 , n250625 );
nand ( n250627 , n240893 , n250626 );
not ( n250628 , n250627 );
and ( n250629 , n250611 , n250628 );
and ( n250630 , n250627 , n37594 );
nor ( n250631 , n250629 , n250630 );
not ( n250632 , n25520 );
not ( n250633 , n33885 );
or ( n250634 , n250632 , n250633 );
or ( n250635 , n33885 , n25520 );
nand ( n250636 , n250634 , n250635 );
and ( n250637 , n250636 , n219538 );
not ( n250638 , n250636 );
and ( n250639 , n250638 , n224022 );
nor ( n250640 , n250637 , n250639 );
nand ( n250641 , n250640 , n240873 );
and ( n250642 , n250641 , n240863 );
not ( n250643 , n250641 );
and ( n250644 , n250643 , n37512 );
nor ( n250645 , n250642 , n250644 );
xor ( n250646 , n250631 , n250645 );
not ( n250647 , n250646 );
not ( n250648 , n250647 );
not ( n250649 , n37670 );
not ( n250650 , n29979 );
not ( n250651 , n204792 );
or ( n250652 , n250650 , n250651 );
or ( n250653 , n204792 , n29979 );
nand ( n250654 , n250652 , n250653 );
and ( n250655 , n250654 , n223510 );
not ( n250656 , n250654 );
and ( n250657 , n250656 , n45750 );
nor ( n250658 , n250655 , n250657 );
not ( n250659 , n250658 );
nand ( n250660 , n240852 , n250659 );
not ( n250661 , n250660 );
or ( n250662 , n250649 , n250661 );
not ( n250663 , n250658 );
nand ( n250664 , n250663 , n240852 );
or ( n250665 , n250664 , n37670 );
nand ( n250666 , n250662 , n250665 );
not ( n250667 , n250666 );
not ( n250668 , n250667 );
or ( n250669 , n250648 , n250668 );
nand ( n250670 , n250646 , n250666 );
nand ( n250671 , n250669 , n250670 );
not ( n250672 , n244365 );
not ( n250673 , n240840 );
or ( n250674 , n250672 , n250673 );
or ( n250675 , n240840 , n244365 );
nand ( n250676 , n250674 , n250675 );
not ( n250677 , n250676 );
and ( n250678 , n250671 , n250677 );
not ( n250679 , n250671 );
and ( n250680 , n250679 , n250676 );
nor ( n250681 , n250678 , n250680 );
buf ( n250682 , n250681 );
and ( n250683 , n250610 , n250682 );
not ( n250684 , n250610 );
buf ( n250685 , n250671 );
buf ( n250686 , n250676 );
and ( n250687 , n250685 , n250686 );
not ( n250688 , n250685 );
not ( n250689 , n250686 );
and ( n250690 , n250688 , n250689 );
nor ( n250691 , n250687 , n250690 );
buf ( n250692 , n250691 );
and ( n250693 , n250684 , n250692 );
nor ( n250694 , n250683 , n250693 );
nor ( n250695 , n250694 , n235895 );
not ( n250696 , n241211 );
not ( n250697 , n250696 );
and ( n250698 , n239749 , n239769 );
not ( n250699 , n239749 );
and ( n250700 , n250699 , n239772 );
nor ( n250701 , n250698 , n250700 );
not ( n250702 , n250701 );
not ( n250703 , n250702 );
or ( n250704 , n250697 , n250703 );
not ( n250705 , n239774 );
or ( n250706 , n250705 , n250696 );
nand ( n250707 , n250704 , n250706 );
not ( n250708 , n245333 );
not ( n250709 , n250708 );
and ( n250710 , n250707 , n250709 );
not ( n250711 , n250707 );
buf ( n250712 , n250708 );
and ( n250713 , n250711 , n250712 );
nor ( n250714 , n250710 , n250713 );
not ( n250715 , n249329 );
not ( n250716 , n235202 );
or ( n250717 , n250715 , n250716 );
nand ( n250718 , n235211 , n249326 );
nand ( n250719 , n250717 , n250718 );
not ( n250720 , n250719 );
buf ( n250721 , n249689 );
not ( n250722 , n250721 );
and ( n250723 , n250720 , n250722 );
and ( n250724 , n250719 , n250721 );
nor ( n250725 , n250723 , n250724 );
nand ( n250726 , n250695 , n250714 , n250725 );
not ( n250727 , n250694 );
not ( n250728 , n250727 );
not ( n250729 , n250725 );
or ( n250730 , n250728 , n250729 );
nor ( n250731 , n250714 , n52445 );
nand ( n250732 , n250730 , n250731 );
nand ( n250733 , n237714 , n209114 );
nand ( n250734 , n250726 , n250732 , n250733 );
buf ( n250735 , n250734 );
buf ( n250736 , n31939 );
not ( n250737 , n250736 );
not ( n250738 , n51269 );
not ( n250739 , n250738 );
or ( n250740 , n250737 , n250739 );
not ( n250741 , n250736 );
nand ( n250742 , n250741 , n51269 );
nand ( n250743 , n250740 , n250742 );
not ( n250744 , n250743 );
not ( n250745 , n53248 );
not ( n250746 , n250745 );
not ( n250747 , n250746 );
and ( n250748 , n250744 , n250747 );
and ( n250749 , n250743 , n250746 );
nor ( n250750 , n250748 , n250749 );
nor ( n250751 , n250750 , n40465 );
not ( n250752 , n250751 );
not ( n250753 , n235848 );
not ( n250754 , n245797 );
not ( n250755 , n250754 );
or ( n250756 , n250753 , n250755 );
nand ( n250757 , n245792 , n235851 );
nand ( n250758 , n250756 , n250757 );
nand ( n250759 , n241612 , n243350 );
not ( n250760 , n250759 );
not ( n250761 , n242486 );
and ( n250762 , n250760 , n250761 );
and ( n250763 , n250759 , n242486 );
nor ( n250764 , n250762 , n250763 );
not ( n250765 , n250764 );
nor ( n250766 , n242427 , n241578 );
not ( n250767 , n250766 );
not ( n250768 , n242417 );
and ( n250769 , n250767 , n250768 );
and ( n250770 , n250766 , n242417 );
nor ( n250771 , n250769 , n250770 );
not ( n250772 , n250771 );
not ( n250773 , n242504 );
nand ( n250774 , n241642 , n243341 );
not ( n250775 , n250774 );
or ( n250776 , n250773 , n250775 );
or ( n250777 , n242504 , n250774 );
nand ( n250778 , n250776 , n250777 );
not ( n250779 , n250778 );
or ( n250780 , n250772 , n250779 );
or ( n250781 , n250771 , n250778 );
nand ( n250782 , n250780 , n250781 );
not ( n250783 , n250782 );
and ( n250784 , n250765 , n250783 );
and ( n250785 , n250764 , n250782 );
nor ( n250786 , n250784 , n250785 );
not ( n250787 , n243299 );
nand ( n250788 , n250787 , n241511 );
buf ( n250789 , n241470 );
xor ( n250790 , n250788 , n250789 );
not ( n250791 , n250790 );
nand ( n250792 , n241551 , n243317 );
and ( n250793 , n250792 , n242447 );
not ( n250794 , n250792 );
and ( n250795 , n250794 , n242448 );
nor ( n250796 , n250793 , n250795 );
not ( n250797 , n250796 );
or ( n250798 , n250791 , n250797 );
or ( n250799 , n250796 , n250790 );
nand ( n250800 , n250798 , n250799 );
and ( n250801 , n250786 , n250800 );
not ( n250802 , n250786 );
not ( n250803 , n250800 );
and ( n250804 , n250802 , n250803 );
nor ( n250805 , n250801 , n250804 );
not ( n250806 , n250805 );
not ( n250807 , n250806 );
buf ( n250808 , n250807 );
and ( n250809 , n250758 , n250808 );
not ( n250810 , n250758 );
not ( n250811 , n250805 );
not ( n250812 , n250811 );
not ( n250813 , n250812 );
and ( n250814 , n250810 , n250813 );
nor ( n250815 , n250809 , n250814 );
not ( n250816 , n39664 );
not ( n250817 , n250816 );
not ( n250818 , n35409 );
or ( n250819 , n250817 , n250818 );
not ( n250820 , n250816 );
nand ( n250821 , n250820 , n35417 );
nand ( n250822 , n250819 , n250821 );
and ( n250823 , n250822 , n249601 );
not ( n250824 , n250822 );
and ( n250825 , n250824 , n249611 );
nor ( n250826 , n250823 , n250825 );
nand ( n250827 , n250815 , n250826 );
or ( n250828 , n250752 , n250827 );
not ( n250829 , n250826 );
not ( n250830 , n250750 );
not ( n250831 , n250830 );
or ( n250832 , n250829 , n250831 );
nor ( n250833 , n250815 , n43968 );
nand ( n250834 , n250832 , n250833 );
nand ( n250835 , n246217 , n34980 );
nand ( n250836 , n250828 , n250834 , n250835 );
buf ( n250837 , n250836 );
not ( n250838 , n244250 );
not ( n250839 , n28929 );
or ( n250840 , n250838 , n250839 );
not ( n250841 , n244250 );
nand ( n250842 , n250841 , n28936 );
nand ( n250843 , n250840 , n250842 );
and ( n250844 , n250843 , n29962 );
not ( n250845 , n250843 );
and ( n250846 , n250845 , n29965 );
nor ( n250847 , n250844 , n250846 );
not ( n250848 , n250847 );
not ( n250849 , n244882 );
not ( n250850 , n250849 );
not ( n250851 , n231421 );
or ( n250852 , n250850 , n250851 );
or ( n250853 , n231421 , n250849 );
nand ( n250854 , n250852 , n250853 );
and ( n250855 , n250854 , n236821 );
not ( n250856 , n250854 );
and ( n250857 , n250856 , n53665 );
nor ( n250858 , n250855 , n250857 );
nand ( n250859 , n250848 , n250858 );
buf ( n250860 , n225155 );
not ( n250861 , n250860 );
not ( n250862 , n47459 );
nand ( n250863 , n250862 , n225223 );
not ( n250864 , n250863 );
not ( n250865 , n48350 );
not ( n250866 , n250865 );
and ( n250867 , n250864 , n250866 );
and ( n250868 , n250863 , n250865 );
nor ( n250869 , n250867 , n250868 );
not ( n250870 , n250869 );
not ( n250871 , n226032 );
not ( n250872 , n249105 );
or ( n250873 , n250871 , n250872 );
or ( n250874 , n249105 , n226032 );
nand ( n250875 , n250873 , n250874 );
not ( n250876 , n250875 );
or ( n250877 , n250870 , n250876 );
or ( n250878 , n250875 , n250869 );
nand ( n250879 , n250877 , n250878 );
not ( n250880 , n234329 );
nand ( n250881 , n241433 , n47517 );
not ( n250882 , n250881 );
not ( n250883 , n48380 );
and ( n250884 , n250882 , n250883 );
and ( n250885 , n250881 , n48380 );
nor ( n250886 , n250884 , n250885 );
not ( n250887 , n250886 );
and ( n250888 , n250880 , n250887 );
and ( n250889 , n234329 , n250886 );
nor ( n250890 , n250888 , n250889 );
and ( n250891 , n250879 , n250890 );
not ( n250892 , n250879 );
not ( n250893 , n250890 );
and ( n250894 , n250892 , n250893 );
nor ( n250895 , n250891 , n250894 );
not ( n250896 , n250895 );
not ( n250897 , n250896 );
or ( n250898 , n250861 , n250897 );
buf ( n250899 , n250895 );
not ( n250900 , n250899 );
or ( n250901 , n250900 , n250860 );
nand ( n250902 , n250898 , n250901 );
buf ( n250903 , n238040 );
and ( n250904 , n250902 , n250903 );
not ( n250905 , n250902 );
buf ( n250906 , n238033 );
and ( n250907 , n250905 , n250906 );
nor ( n250908 , n250904 , n250907 );
buf ( n250909 , n43517 );
nor ( n250910 , n250908 , n250909 );
not ( n250911 , n250910 );
or ( n250912 , n250859 , n250911 );
not ( n250913 , n250908 );
nor ( n250914 , n250913 , n49051 );
nand ( n250915 , n250914 , n250859 );
buf ( n250916 , n35431 );
nand ( n250917 , n250916 , n36746 );
nand ( n250918 , n250912 , n250915 , n250917 );
buf ( n250919 , n250918 );
not ( n250920 , n247981 );
not ( n250921 , n239930 );
or ( n250922 , n250920 , n250921 );
or ( n250923 , n239930 , n247981 );
nand ( n250924 , n250922 , n250923 );
and ( n250925 , n250924 , n243511 );
not ( n250926 , n250924 );
and ( n250927 , n250926 , n243504 );
nor ( n250928 , n250925 , n250927 );
not ( n250929 , n55146 );
nand ( n250930 , n250928 , n250929 );
not ( n250931 , n250168 );
nand ( n250932 , n250931 , n248619 );
buf ( n250933 , n243091 );
xor ( n250934 , n250932 , n250933 );
not ( n250935 , n250934 );
not ( n250936 , n250234 );
or ( n250937 , n250935 , n250936 );
not ( n250938 , n250934 );
nand ( n250939 , n250938 , n250230 );
nand ( n250940 , n250937 , n250939 );
not ( n250941 , n250940 );
buf ( n250942 , n50274 );
not ( n250943 , n250942 );
and ( n250944 , n250941 , n250943 );
and ( n250945 , n250940 , n250942 );
nor ( n250946 , n250944 , n250945 );
nand ( n250947 , n223191 , n55804 );
not ( n250948 , n250947 );
buf ( n250949 , n226849 );
not ( n250950 , n250949 );
not ( n250951 , n250950 );
and ( n250952 , n250948 , n250951 );
and ( n250953 , n250947 , n250950 );
nor ( n250954 , n250952 , n250953 );
not ( n250955 , n250954 );
not ( n250956 , n250955 );
not ( n250957 , n55889 );
or ( n250958 , n250956 , n250957 );
not ( n250959 , n250955 );
nand ( n250960 , n250959 , n233660 );
nand ( n250961 , n250958 , n250960 );
and ( n250962 , n250961 , n233805 );
not ( n250963 , n250961 );
not ( n250964 , n56040 );
and ( n250965 , n250963 , n250964 );
nor ( n250966 , n250962 , n250965 );
not ( n250967 , n250966 );
nand ( n250968 , n250946 , n250967 );
or ( n250969 , n250930 , n250968 );
nor ( n250970 , n250928 , n237384 );
nand ( n250971 , n250968 , n250970 );
nand ( n250972 , n247423 , n204559 );
nand ( n250973 , n250969 , n250971 , n250972 );
buf ( n250974 , n250973 );
not ( n250975 , RI19ab63d8_2407);
or ( n250976 , n25328 , n250975 );
not ( n250977 , RI19aaca18_2478);
or ( n250978 , n226822 , n250977 );
nand ( n250979 , n250976 , n250978 );
buf ( n250980 , n250979 );
nor ( n250981 , n244060 , n226003 );
not ( n250982 , n250981 );
not ( n250983 , n238386 );
not ( n250984 , n245081 );
nand ( n250985 , n250983 , n250984 );
not ( n250986 , n250985 );
not ( n250987 , n53978 );
and ( n250988 , n250986 , n250987 );
nand ( n250989 , n250984 , n238387 );
and ( n250990 , n250989 , n53978 );
nor ( n250991 , n250988 , n250990 );
not ( n250992 , n250991 );
not ( n250993 , n245093 );
nand ( n250994 , n250993 , n238367 );
and ( n250995 , n250994 , n231703 );
not ( n250996 , n250994 );
and ( n250997 , n250996 , n53943 );
nor ( n250998 , n250995 , n250997 );
not ( n250999 , n250998 );
or ( n251000 , n250992 , n250999 );
or ( n251001 , n250998 , n250991 );
nand ( n251002 , n251000 , n251001 );
not ( n251003 , n251002 );
not ( n251004 , n231670 );
nand ( n251005 , n245061 , n238351 );
not ( n251006 , n251005 );
or ( n251007 , n251004 , n251006 );
or ( n251008 , n251005 , n231670 );
nand ( n251009 , n251007 , n251008 );
not ( n251010 , n251009 );
nand ( n251011 , n238312 , n245031 );
not ( n251012 , n251011 );
not ( n251013 , n231603 );
and ( n251014 , n251012 , n251013 );
and ( n251015 , n251011 , n231603 );
nor ( n251016 , n251014 , n251015 );
not ( n251017 , n251016 );
or ( n251018 , n251010 , n251017 );
or ( n251019 , n251016 , n251009 );
nand ( n251020 , n251018 , n251019 );
and ( n251021 , n251020 , n245020 );
not ( n251022 , n251020 );
and ( n251023 , n251022 , n245021 );
nor ( n251024 , n251021 , n251023 );
not ( n251025 , n251024 );
and ( n251026 , n251003 , n251025 );
and ( n251027 , n251002 , n251024 );
nor ( n251028 , n251026 , n251027 );
buf ( n251029 , n251028 );
not ( n251030 , n251029 );
not ( n251031 , n236114 );
nand ( n251032 , n238271 , n50427 );
not ( n251033 , n251032 );
not ( n251034 , n53783 );
and ( n251035 , n251033 , n251034 );
and ( n251036 , n251032 , n53783 );
nor ( n251037 , n251035 , n251036 );
not ( n251038 , n236131 );
nand ( n251039 , n50436 , n251038 );
and ( n251040 , n251039 , n228208 );
not ( n251041 , n251039 );
and ( n251042 , n251041 , n53762 );
nor ( n251043 , n251040 , n251042 );
and ( n251044 , n251037 , n251043 );
not ( n251045 , n251037 );
not ( n251046 , n251043 );
and ( n251047 , n251045 , n251046 );
nor ( n251048 , n251044 , n251047 );
not ( n251049 , n251048 );
not ( n251050 , n251049 );
nand ( n251051 , n50337 , n236110 );
not ( n251052 , n251051 );
not ( n251053 , n53721 );
or ( n251054 , n251052 , n251053 );
or ( n251055 , n53721 , n251051 );
nand ( n251056 , n251054 , n251055 );
not ( n251057 , n251056 );
nand ( n251058 , n236090 , n228139 );
not ( n251059 , n251058 );
not ( n251060 , n50367 );
and ( n251061 , n251059 , n251060 );
and ( n251062 , n251058 , n50367 );
nor ( n251063 , n251061 , n251062 );
not ( n251064 , n251063 );
or ( n251065 , n251057 , n251064 );
or ( n251066 , n251063 , n251056 );
nand ( n251067 , n251065 , n251066 );
nand ( n251068 , n238237 , n50294 );
and ( n251069 , n251068 , n50305 );
not ( n251070 , n251068 );
and ( n251071 , n251070 , n53701 );
nor ( n251072 , n251069 , n251071 );
and ( n251073 , n251067 , n251072 );
not ( n251074 , n251067 );
not ( n251075 , n251072 );
and ( n251076 , n251074 , n251075 );
nor ( n251077 , n251073 , n251076 );
not ( n251078 , n251077 );
not ( n251079 , n251078 );
or ( n251080 , n251050 , n251079 );
nand ( n251081 , n251077 , n251048 );
nand ( n251082 , n251080 , n251081 );
not ( n251083 , n251082 );
or ( n251084 , n251031 , n251083 );
or ( n251085 , n251082 , n236114 );
nand ( n251086 , n251084 , n251085 );
not ( n251087 , n251086 );
and ( n251088 , n251030 , n251087 );
and ( n251089 , n251029 , n251086 );
nor ( n251090 , n251088 , n251089 );
nand ( n251091 , n243697 , n251090 );
nor ( n251092 , n250982 , n251091 );
nor ( n251093 , n251090 , n40465 );
not ( n251094 , n251093 );
nor ( n251095 , n251094 , n243697 );
nor ( n251096 , n251092 , n251095 );
not ( n251097 , n251090 );
nand ( n251098 , n244062 , n251097 );
nand ( n251099 , n244987 , n36182 );
nand ( n251100 , n251096 , n251098 , n251099 );
buf ( n251101 , n251100 );
not ( n251102 , RI19aa9868_2499);
or ( n251103 , n226819 , n251102 );
not ( n251104 , RI19a9fae8_2571);
or ( n251105 , n25335 , n251104 );
nand ( n251106 , n251103 , n251105 );
buf ( n251107 , n251106 );
not ( n251108 , n245751 );
not ( n251109 , n251108 );
not ( n251110 , n52756 );
or ( n251111 , n251109 , n251110 );
nand ( n251112 , n245264 , n245751 );
nand ( n251113 , n251111 , n251112 );
not ( n251114 , n251113 );
not ( n251115 , n249005 );
not ( n251116 , n251115 );
not ( n251117 , n241470 );
nand ( n251118 , n251117 , n243299 );
buf ( n251119 , n241479 );
xor ( n251120 , n251118 , n251119 );
not ( n251121 , n251120 );
not ( n251122 , n251121 );
or ( n251123 , n251116 , n251122 );
nand ( n251124 , n251120 , n249005 );
nand ( n251125 , n251123 , n251124 );
and ( n251126 , n251125 , n242434 );
not ( n251127 , n251125 );
and ( n251128 , n251127 , n242435 );
nor ( n251129 , n251126 , n251128 );
not ( n251130 , n251129 );
not ( n251131 , n242486 );
nand ( n251132 , n251131 , n243351 );
not ( n251133 , n251132 );
not ( n251134 , n241602 );
and ( n251135 , n251133 , n251134 );
and ( n251136 , n251132 , n241602 );
nor ( n251137 , n251135 , n251136 );
not ( n251138 , n251137 );
not ( n251139 , n242504 );
nand ( n251140 , n251139 , n243342 );
not ( n251141 , n251140 );
not ( n251142 , n241621 );
or ( n251143 , n251141 , n251142 );
or ( n251144 , n241621 , n251140 );
nand ( n251145 , n251143 , n251144 );
not ( n251146 , n251145 );
and ( n251147 , n251138 , n251146 );
and ( n251148 , n251137 , n251145 );
nor ( n251149 , n251147 , n251148 );
not ( n251150 , n251149 );
and ( n251151 , n251130 , n251150 );
not ( n251152 , n251130 );
and ( n251153 , n251152 , n251149 );
nor ( n251154 , n251151 , n251153 );
not ( n251155 , n251154 );
not ( n251156 , n251155 );
not ( n251157 , n251156 );
and ( n251158 , n251114 , n251157 );
and ( n251159 , n251113 , n251156 );
nor ( n251160 , n251158 , n251159 );
not ( n251161 , n54497 );
buf ( n251162 , n245472 );
not ( n251163 , n251162 );
or ( n251164 , n251161 , n251163 );
not ( n251165 , n54497 );
nand ( n251166 , n251165 , n245473 );
nand ( n251167 , n251164 , n251166 );
buf ( n251168 , n53657 );
and ( n251169 , n251167 , n251168 );
not ( n251170 , n251167 );
not ( n251171 , n251168 );
and ( n251172 , n251170 , n251171 );
nor ( n251173 , n251169 , n251172 );
nand ( n251174 , n251160 , n251173 );
not ( n251175 , n52132 );
not ( n251176 , n236267 );
or ( n251177 , n251175 , n251176 );
not ( n251178 , n52132 );
nand ( n251179 , n251178 , n245210 );
nand ( n251180 , n251177 , n251179 );
not ( n251181 , n44539 );
xor ( n251182 , n251180 , n251181 );
nor ( n251183 , n251182 , n226955 );
not ( n251184 , n251183 );
or ( n251185 , n251174 , n251184 );
not ( n251186 , n251182 );
not ( n251187 , n251186 );
not ( n251188 , n251160 );
or ( n251189 , n251187 , n251188 );
buf ( n251190 , n233971 );
nor ( n251191 , n251173 , n251190 );
nand ( n251192 , n251189 , n251191 );
nand ( n251193 , n237361 , n41322 );
nand ( n251194 , n251185 , n251192 , n251193 );
buf ( n251195 , n251194 );
not ( n251196 , n45293 );
not ( n251197 , n234453 );
or ( n251198 , n251196 , n251197 );
not ( n251199 , n51292 );
not ( n251200 , n43005 );
or ( n251201 , n251199 , n251200 );
nand ( n251202 , n43010 , n51293 );
nand ( n251203 , n251201 , n251202 );
and ( n251204 , n251203 , n50027 );
not ( n251205 , n251203 );
and ( n251206 , n251205 , n227796 );
nor ( n251207 , n251204 , n251206 );
not ( n251208 , n55983 );
not ( n251209 , n238156 );
not ( n251210 , n238177 );
and ( n251211 , n251209 , n251210 );
and ( n251212 , n238156 , n238177 );
nor ( n251213 , n251211 , n251212 );
not ( n251214 , n251213 );
or ( n251215 , n251208 , n251214 );
not ( n251216 , n55983 );
not ( n251217 , n251213 );
nand ( n251218 , n251216 , n251217 );
nand ( n251219 , n251215 , n251218 );
buf ( n251220 , n235807 );
and ( n251221 , n251219 , n251220 );
not ( n251222 , n251219 );
not ( n251223 , n235815 );
not ( n251224 , n251223 );
and ( n251225 , n251222 , n251224 );
nor ( n251226 , n251221 , n251225 );
nand ( n251227 , n251207 , n251226 );
not ( n251228 , n245369 );
not ( n251229 , n251228 );
not ( n251230 , n235357 );
or ( n251231 , n251229 , n251230 );
not ( n251232 , n251228 );
nand ( n251233 , n251232 , n235366 );
nand ( n251234 , n251231 , n251233 );
and ( n251235 , n251234 , n235369 );
not ( n251236 , n251234 );
and ( n251237 , n251236 , n235372 );
nor ( n251238 , n251235 , n251237 );
not ( n251239 , n251238 );
and ( n251240 , n251227 , n251239 );
not ( n251241 , n251227 );
and ( n251242 , n251241 , n251238 );
nor ( n251243 , n251240 , n251242 );
or ( n251244 , n251243 , n240080 );
nand ( n251245 , n251198 , n251244 );
buf ( n251246 , n251245 );
buf ( n251247 , n250764 );
not ( n251248 , n251247 );
not ( n251249 , n251149 );
not ( n251250 , n251129 );
or ( n251251 , n251249 , n251250 );
nand ( n251252 , n251130 , n251150 );
nand ( n251253 , n251251 , n251252 );
not ( n251254 , n251253 );
or ( n251255 , n251248 , n251254 );
or ( n251256 , n251253 , n251247 );
nand ( n251257 , n251255 , n251256 );
not ( n251258 , n38936 );
nand ( n251259 , n251258 , n38711 );
not ( n251260 , n251259 );
not ( n251261 , n49771 );
and ( n251262 , n251260 , n251261 );
and ( n251263 , n251259 , n49771 );
nor ( n251264 , n251262 , n251263 );
not ( n251265 , n251264 );
not ( n251266 , n39038 );
nand ( n251267 , n251266 , n39011 );
not ( n251268 , n251267 );
not ( n251269 , n227523 );
and ( n251270 , n251268 , n251269 );
and ( n251271 , n251267 , n227523 );
nor ( n251272 , n251270 , n251271 );
not ( n251273 , n251272 );
not ( n251274 , n251273 );
or ( n251275 , n251265 , n251274 );
not ( n251276 , n251264 );
nand ( n251277 , n251276 , n251272 );
nand ( n251278 , n251275 , n251277 );
xor ( n251279 , n249936 , n251278 );
nand ( n251280 , n38755 , n243396 );
and ( n251281 , n251280 , n242554 );
not ( n251282 , n251280 );
and ( n251283 , n251282 , n49697 );
nor ( n251284 , n251281 , n251283 );
not ( n251285 , n251284 );
not ( n251286 , n251285 );
nand ( n251287 , n38832 , n38915 );
not ( n251288 , n251287 );
not ( n251289 , n227489 );
and ( n251290 , n251288 , n251289 );
and ( n251291 , n251287 , n227489 );
nor ( n251292 , n251290 , n251291 );
not ( n251293 , n251292 );
not ( n251294 , n251293 );
or ( n251295 , n251286 , n251294 );
nand ( n251296 , n251292 , n251284 );
nand ( n251297 , n251295 , n251296 );
xor ( n251298 , n251279 , n251297 );
buf ( n251299 , n251298 );
and ( n251300 , n251257 , n251299 );
not ( n251301 , n251257 );
not ( n251302 , n251278 );
not ( n251303 , n251302 );
not ( n251304 , n249936 );
and ( n251305 , n251297 , n251304 );
not ( n251306 , n251297 );
and ( n251307 , n251306 , n249936 );
nor ( n251308 , n251305 , n251307 );
not ( n251309 , n251308 );
or ( n251310 , n251303 , n251309 );
not ( n251311 , n251308 );
nand ( n251312 , n251311 , n251278 );
nand ( n251313 , n251310 , n251312 );
buf ( n251314 , n251313 );
and ( n251315 , n251301 , n251314 );
nor ( n251316 , n251300 , n251315 );
nor ( n251317 , n251316 , n250909 );
not ( n251318 , n51563 );
nand ( n251319 , n36528 , n36552 );
not ( n251320 , n251319 );
or ( n251321 , n251318 , n251320 );
nand ( n251322 , n36528 , n36552 );
or ( n251323 , n251322 , n51563 );
nand ( n251324 , n251321 , n251323 );
not ( n251325 , n251324 );
not ( n251326 , n46506 );
or ( n251327 , n251325 , n251326 );
not ( n251328 , n251324 );
nand ( n251329 , n251328 , n46514 );
nand ( n251330 , n251327 , n251329 );
and ( n251331 , n251330 , n224478 );
not ( n251332 , n251330 );
buf ( n251333 , n46708 );
and ( n251334 , n251332 , n251333 );
nor ( n251335 , n251331 , n251334 );
not ( n251336 , n240042 );
not ( n251337 , n40194 );
or ( n251338 , n251336 , n251337 );
not ( n251339 , n240042 );
nand ( n251340 , n251339 , n40203 );
nand ( n251341 , n251338 , n251340 );
and ( n251342 , n40340 , n40455 );
not ( n251343 , n40340 );
and ( n251344 , n251343 , n40456 );
nor ( n251345 , n251342 , n251344 );
buf ( n251346 , n251345 );
and ( n251347 , n251341 , n251346 );
not ( n251348 , n251341 );
not ( n251349 , n40460 );
not ( n251350 , n251349 );
and ( n251351 , n251348 , n251350 );
nor ( n251352 , n251347 , n251351 );
nor ( n251353 , n251335 , n251352 );
nand ( n251354 , n251317 , n251353 );
not ( n251355 , n251352 );
not ( n251356 , n251355 );
not ( n251357 , n251316 );
not ( n251358 , n251357 );
or ( n251359 , n251356 , n251358 );
not ( n251360 , n251335 );
buf ( n251361 , n31571 );
nor ( n251362 , n251360 , n251361 );
nand ( n251363 , n251359 , n251362 );
nand ( n251364 , n231444 , n28319 );
nand ( n251365 , n251354 , n251363 , n251364 );
buf ( n251366 , n251365 );
buf ( n251367 , n25482 );
buf ( n251368 , n247303 );
not ( n251369 , n251368 );
not ( n251370 , n246166 );
or ( n251371 , n251369 , n251370 );
not ( n251372 , n246171 );
or ( n251373 , n251372 , n251368 );
nand ( n251374 , n251371 , n251373 );
not ( n251375 , n251374 );
not ( n251376 , n250682 );
and ( n251377 , n251375 , n251376 );
and ( n251378 , n251374 , n250682 );
nor ( n251379 , n251377 , n251378 );
nor ( n251380 , n251379 , n35428 );
not ( n251381 , n250471 );
not ( n251382 , n234682 );
or ( n251383 , n251381 , n251382 );
nand ( n251384 , n234691 , n250474 );
nand ( n251385 , n251383 , n251384 );
and ( n251386 , n251385 , n234804 );
not ( n251387 , n251385 );
and ( n251388 , n251387 , n234811 );
nor ( n251389 , n251386 , n251388 );
not ( n251390 , n231648 );
not ( n251391 , n238400 );
or ( n251392 , n251390 , n251391 );
not ( n251393 , n231648 );
nand ( n251394 , n251393 , n238408 );
nand ( n251395 , n251392 , n251394 );
not ( n251396 , n40595 );
nand ( n251397 , n251396 , n40478 );
buf ( n251398 , n47217 );
xor ( n251399 , n251397 , n251398 );
not ( n251400 , n251399 );
not ( n251401 , n251400 );
nand ( n251402 , n40638 , n40611 );
buf ( n251403 , n224950 );
xor ( n251404 , n251402 , n251403 );
not ( n251405 , n251404 );
not ( n251406 , n251405 );
or ( n251407 , n251401 , n251406 );
nand ( n251408 , n251399 , n251404 );
nand ( n251409 , n251407 , n251408 );
not ( n251410 , n218511 );
nand ( n251411 , n251410 , n245155 );
buf ( n251412 , n47245 );
xnor ( n251413 , n251411 , n251412 );
not ( n251414 , n251413 );
and ( n251415 , n251409 , n251414 );
not ( n251416 , n251409 );
and ( n251417 , n251416 , n251413 );
nor ( n251418 , n251415 , n251417 );
nand ( n251419 , n244636 , n245122 );
not ( n251420 , n251419 );
not ( n251421 , n47294 );
or ( n251422 , n251420 , n251421 );
or ( n251423 , n47294 , n251419 );
nand ( n251424 , n251422 , n251423 );
not ( n251425 , n251424 );
not ( n251426 , n251425 );
not ( n251427 , n40900 );
nand ( n251428 , n251427 , n245130 );
not ( n251429 , n251428 );
not ( n251430 , n47275 );
and ( n251431 , n251429 , n251430 );
and ( n251432 , n251428 , n47275 );
nor ( n251433 , n251431 , n251432 );
not ( n251434 , n251433 );
not ( n251435 , n251434 );
or ( n251436 , n251426 , n251435 );
nand ( n251437 , n251433 , n251424 );
nand ( n251438 , n251436 , n251437 );
not ( n251439 , n251438 );
and ( n251440 , n251418 , n251439 );
not ( n251441 , n251418 );
and ( n251442 , n251441 , n251438 );
nor ( n251443 , n251440 , n251442 );
buf ( n251444 , n251443 );
and ( n251445 , n251395 , n251444 );
not ( n251446 , n251395 );
and ( n251447 , n251418 , n251438 );
not ( n251448 , n251418 );
and ( n251449 , n251448 , n251439 );
nor ( n251450 , n251447 , n251449 );
buf ( n251451 , n251450 );
and ( n251452 , n251446 , n251451 );
nor ( n251453 , n251445 , n251452 );
nor ( n251454 , n251389 , n251453 );
nand ( n251455 , n251380 , n251454 );
not ( n251456 , n251453 );
not ( n251457 , n251456 );
not ( n251458 , n251379 );
not ( n251459 , n251458 );
or ( n251460 , n251457 , n251459 );
not ( n251461 , n251389 );
not ( n251462 , n205649 );
nor ( n251463 , n251461 , n251462 );
nand ( n251464 , n251460 , n251463 );
buf ( n251465 , n31577 );
nand ( n251466 , n251465 , n30240 );
nand ( n251467 , n251455 , n251464 , n251466 );
buf ( n251468 , n251467 );
not ( n251469 , n33386 );
not ( n251470 , n39766 );
or ( n251471 , n251469 , n251470 );
not ( n251472 , n241513 );
not ( n251473 , n243363 );
or ( n251474 , n251472 , n251473 );
not ( n251475 , n241513 );
nand ( n251476 , n251475 , n243372 );
nand ( n251477 , n251474 , n251476 );
and ( n251478 , n251477 , n243416 );
not ( n251479 , n251477 );
and ( n251480 , n251479 , n246694 );
nor ( n251481 , n251478 , n251480 );
not ( n251482 , n54282 );
not ( n251483 , n51342 );
or ( n251484 , n251482 , n251483 );
not ( n251485 , n54282 );
nand ( n251486 , n251485 , n51343 );
nand ( n251487 , n251484 , n251486 );
buf ( n251488 , n38232 );
and ( n251489 , n251487 , n251488 );
not ( n251490 , n251487 );
and ( n251491 , n251490 , n51349 );
nor ( n251492 , n251489 , n251491 );
nand ( n251493 , n251481 , n251492 );
and ( n251494 , n251493 , n247021 );
not ( n251495 , n251493 );
and ( n251496 , n251495 , n247217 );
nor ( n251497 , n251494 , n251496 );
buf ( n251498 , n249531 );
or ( n251499 , n251497 , n251498 );
nand ( n251500 , n251471 , n251499 );
buf ( n251501 , n251500 );
buf ( n251502 , n234289 );
not ( n251503 , n251502 );
not ( n251504 , n43725 );
not ( n251505 , n251504 );
or ( n251506 , n251503 , n251505 );
or ( n251507 , n43726 , n251502 );
nand ( n251508 , n251506 , n251507 );
and ( n251509 , n251508 , n43956 );
not ( n251510 , n251508 );
and ( n251511 , n251510 , n43964 );
nor ( n251512 , n251509 , n251511 );
nor ( n251513 , n251512 , n244399 );
not ( n251514 , n239435 );
nand ( n251515 , n251514 , n239420 );
and ( n251516 , n251515 , n248326 );
not ( n251517 , n251515 );
and ( n251518 , n251517 , n248327 );
nor ( n251519 , n251516 , n251518 );
not ( n251520 , n251519 );
not ( n251521 , n251520 );
and ( n251522 , n249666 , n249684 );
not ( n251523 , n249666 );
and ( n251524 , n251523 , n249687 );
nor ( n251525 , n251522 , n251524 );
not ( n251526 , n251525 );
not ( n251527 , n251526 );
or ( n251528 , n251521 , n251527 );
or ( n251529 , n249693 , n251520 );
nand ( n251530 , n251528 , n251529 );
not ( n251531 , n251530 );
buf ( n251532 , n249757 );
not ( n251533 , n251532 );
and ( n251534 , n251531 , n251533 );
and ( n251535 , n251530 , n251532 );
nor ( n251536 , n251534 , n251535 );
not ( n251537 , n244475 );
buf ( n251538 , n233932 );
not ( n251539 , n251538 );
not ( n251540 , n244346 );
or ( n251541 , n251539 , n251540 );
or ( n251542 , n244346 , n251538 );
nand ( n251543 , n251541 , n251542 );
not ( n251544 , n251543 );
or ( n251545 , n251537 , n251544 );
or ( n251546 , n251543 , n244475 );
nand ( n251547 , n251545 , n251546 );
nor ( n251548 , n251536 , n251547 );
nand ( n251549 , n251513 , n251548 );
not ( n251550 , n251536 );
not ( n251551 , n251550 );
not ( n251552 , n251512 );
not ( n251553 , n251552 );
or ( n251554 , n251551 , n251553 );
not ( n251555 , n251547 );
nor ( n251556 , n251555 , n234440 );
nand ( n251557 , n251554 , n251556 );
nand ( n251558 , n247585 , n32119 );
nand ( n251559 , n251549 , n251557 , n251558 );
buf ( n251560 , n251559 );
buf ( n251561 , RI19a822e0_2779);
buf ( n251562 , n25361 );
and ( n251563 , n251561 , n251562 , n25326 );
buf ( n251564 , n251563 );
not ( n251565 , RI19ac63c8_2283);
or ( n251566 , n25328 , n251565 );
not ( n251567 , RI19abd890_2354);
or ( n251568 , n25336 , n251567 );
nand ( n251569 , n251566 , n251568 );
buf ( n251570 , n251569 );
buf ( n251571 , n32000 );
not ( n251572 , n240001 );
not ( n251573 , n251572 );
not ( n251574 , n251573 );
not ( n251575 , n234163 );
not ( n251576 , n251575 );
not ( n251577 , n233558 );
not ( n251578 , n251577 );
nand ( n251579 , n55833 , n223252 );
and ( n251580 , n251579 , n223077 );
not ( n251581 , n251579 );
and ( n251582 , n251581 , n55835 );
nor ( n251583 , n251580 , n251582 );
not ( n251584 , n251583 );
not ( n251585 , n251584 );
or ( n251586 , n251578 , n251585 );
nand ( n251587 , n251583 , n233558 );
nand ( n251588 , n251586 , n251587 );
and ( n251589 , n251588 , n250954 );
not ( n251590 , n251588 );
and ( n251591 , n251590 , n250955 );
nor ( n251592 , n251589 , n251591 );
not ( n251593 , n251592 );
not ( n251594 , n251593 );
not ( n251595 , n233636 );
nand ( n251596 , n45386 , n251595 );
buf ( n251597 , n226900 );
and ( n251598 , n251596 , n251597 );
not ( n251599 , n251596 );
not ( n251600 , n251597 );
and ( n251601 , n251599 , n251600 );
nor ( n251602 , n251598 , n251601 );
not ( n251603 , n251602 );
not ( n251604 , n251603 );
nand ( n251605 , n55856 , n45361 );
and ( n251606 , n251605 , n226928 );
not ( n251607 , n251605 );
and ( n251608 , n251607 , n233619 );
nor ( n251609 , n251606 , n251608 );
not ( n251610 , n251609 );
not ( n251611 , n251610 );
or ( n251612 , n251604 , n251611 );
nand ( n251613 , n251609 , n251602 );
nand ( n251614 , n251612 , n251613 );
not ( n251615 , n251614 );
not ( n251616 , n251615 );
and ( n251617 , n251594 , n251616 );
and ( n251618 , n251593 , n251615 );
nor ( n251619 , n251617 , n251618 );
not ( n251620 , n251619 );
or ( n251621 , n251576 , n251620 );
not ( n251622 , n251575 );
not ( n251623 , n251615 );
not ( n251624 , n251593 );
or ( n251625 , n251623 , n251624 );
nand ( n251626 , n251592 , n251614 );
nand ( n251627 , n251625 , n251626 );
nand ( n251628 , n251622 , n251627 );
nand ( n251629 , n251621 , n251628 );
not ( n251630 , n251629 );
or ( n251631 , n251574 , n251630 );
or ( n251632 , n251629 , n251573 );
nand ( n251633 , n251631 , n251632 );
not ( n251634 , n251633 );
nand ( n251635 , n251634 , n223839 );
buf ( n251636 , n237862 );
not ( n251637 , n251636 );
not ( n251638 , n224660 );
not ( n251639 , n251638 );
not ( n251640 , n46909 );
nand ( n251641 , n251640 , n228493 );
not ( n251642 , n251641 );
or ( n251643 , n251639 , n251642 );
not ( n251644 , n46909 );
nand ( n251645 , n251644 , n228493 );
or ( n251646 , n251645 , n251638 );
nand ( n251647 , n251643 , n251646 );
not ( n251648 , n251647 );
not ( n251649 , n224520 );
and ( n251650 , n251648 , n251649 );
and ( n251651 , n251647 , n224520 );
nor ( n251652 , n251650 , n251651 );
not ( n251653 , n251652 );
nand ( n251654 , n50674 , n46818 );
and ( n251655 , n251654 , n46806 );
not ( n251656 , n251654 );
and ( n251657 , n251656 , n50620 );
nor ( n251658 , n251655 , n251657 );
nand ( n251659 , n237829 , n50650 );
not ( n251660 , n251659 );
not ( n251661 , n247428 );
and ( n251662 , n251660 , n251661 );
and ( n251663 , n251659 , n247428 );
nor ( n251664 , n251662 , n251663 );
or ( n251665 , n251658 , n251664 );
nand ( n251666 , n251664 , n251658 );
nand ( n251667 , n251665 , n251666 );
nand ( n251668 , n46853 , n228469 );
not ( n251669 , n251668 );
not ( n251670 , n46850 );
and ( n251671 , n251669 , n251670 );
and ( n251672 , n251668 , n46850 );
nor ( n251673 , n251671 , n251672 );
not ( n251674 , n251673 );
and ( n251675 , n251667 , n251674 );
not ( n251676 , n251667 );
and ( n251677 , n251676 , n251673 );
nor ( n251678 , n251675 , n251677 );
not ( n251679 , n251678 );
or ( n251680 , n251653 , n251679 );
not ( n251681 , n251678 );
not ( n251682 , n251652 );
nand ( n251683 , n251681 , n251682 );
nand ( n251684 , n251680 , n251683 );
not ( n251685 , n251684 );
or ( n251686 , n251637 , n251685 );
or ( n251687 , n251684 , n251636 );
nand ( n251688 , n251686 , n251687 );
not ( n251689 , n245994 );
and ( n251690 , n251688 , n251689 );
not ( n251691 , n251688 );
buf ( n251692 , n251689 );
not ( n251693 , n251692 );
and ( n251694 , n251691 , n251693 );
nor ( n251695 , n251690 , n251694 );
not ( n251696 , n249446 );
not ( n251697 , n251696 );
not ( n251698 , n38633 );
or ( n251699 , n251697 , n251698 );
not ( n251700 , n251696 );
nand ( n251701 , n251700 , n38625 );
nand ( n251702 , n251699 , n251701 );
and ( n251703 , n251702 , n49182 );
not ( n251704 , n251702 );
and ( n251705 , n251704 , n49191 );
nor ( n251706 , n251703 , n251705 );
nand ( n251707 , n251695 , n251706 );
or ( n251708 , n251635 , n251707 );
nand ( n251709 , n251633 , n226010 );
not ( n251710 , n251709 );
nand ( n251711 , n251710 , n251707 );
buf ( n251712 , n35431 );
nand ( n251713 , n251712 , n38968 );
nand ( n251714 , n251708 , n251711 , n251713 );
buf ( n251715 , n251714 );
not ( n251716 , n220690 );
buf ( n251717 , n35431 );
not ( n251718 , n251717 );
or ( n251719 , n251716 , n251718 );
not ( n251720 , n40194 );
not ( n251721 , n251720 );
not ( n251722 , n251721 );
not ( n251723 , n239945 );
not ( n251724 , n56040 );
or ( n251725 , n251723 , n251724 );
nand ( n251726 , n250964 , n239946 );
nand ( n251727 , n251725 , n251726 );
not ( n251728 , n251727 );
or ( n251729 , n251722 , n251728 );
buf ( n251730 , n40194 );
or ( n251731 , n251727 , n251730 );
nand ( n251732 , n251729 , n251731 );
not ( n251733 , n251732 );
not ( n251734 , n47522 );
not ( n251735 , n250899 );
or ( n251736 , n251734 , n251735 );
not ( n251737 , n47522 );
nand ( n251738 , n251737 , n250896 );
nand ( n251739 , n251736 , n251738 );
and ( n251740 , n251739 , n250906 );
not ( n251741 , n251739 );
and ( n251742 , n251741 , n250903 );
nor ( n251743 , n251740 , n251742 );
not ( n251744 , n249207 );
not ( n251745 , n237188 );
not ( n251746 , n249195 );
or ( n251747 , n251745 , n251746 );
nand ( n251748 , n249204 , n237187 );
nand ( n251749 , n251747 , n251748 );
not ( n251750 , n251749 );
or ( n251751 , n251744 , n251750 );
or ( n251752 , n251749 , n249207 );
nand ( n251753 , n251751 , n251752 );
nand ( n251754 , n251743 , n251753 );
not ( n251755 , n251754 );
and ( n251756 , n251733 , n251755 );
and ( n251757 , n251732 , n251754 );
nor ( n251758 , n251756 , n251757 );
or ( n251759 , n251758 , n31572 );
nand ( n251760 , n251719 , n251759 );
buf ( n251761 , n251760 );
not ( n251762 , n251583 );
not ( n251763 , n251762 );
not ( n251764 , n55889 );
or ( n251765 , n251763 , n251764 );
not ( n251766 , n251762 );
nand ( n251767 , n251766 , n233660 );
nand ( n251768 , n251765 , n251767 );
and ( n251769 , n251768 , n250964 );
not ( n251770 , n251768 );
not ( n251771 , n56041 );
and ( n251772 , n251770 , n251771 );
nor ( n251773 , n251769 , n251772 );
not ( n251774 , n251773 );
not ( n251775 , n250543 );
not ( n251776 , n251775 );
not ( n251777 , n227174 );
or ( n251778 , n251776 , n251777 );
not ( n251779 , n251775 );
nand ( n251780 , n251779 , n49420 );
nand ( n251781 , n251778 , n251780 );
and ( n251782 , n251781 , n49618 );
not ( n251783 , n251781 );
and ( n251784 , n251783 , n49627 );
nor ( n251785 , n251782 , n251784 );
not ( n251786 , n251785 );
nand ( n251787 , n251774 , n251786 );
not ( n251788 , n248546 );
not ( n251789 , n243659 );
or ( n251790 , n251788 , n251789 );
or ( n251791 , n243659 , n248546 );
nand ( n251792 , n251790 , n251791 );
nand ( n251793 , n243115 , n248618 );
not ( n251794 , n251793 );
not ( n251795 , n250168 );
and ( n251796 , n251794 , n251795 );
nand ( n251797 , n243115 , n248618 );
and ( n251798 , n251797 , n250168 );
nor ( n251799 , n251796 , n251798 );
not ( n251800 , n251799 );
not ( n251801 , n251800 );
nand ( n251802 , n248662 , n243148 );
not ( n251803 , n251802 );
not ( n251804 , n249371 );
or ( n251805 , n251803 , n251804 );
or ( n251806 , n249371 , n251802 );
nand ( n251807 , n251805 , n251806 );
not ( n251808 , n251807 );
not ( n251809 , n251808 );
or ( n251810 , n251801 , n251809 );
nand ( n251811 , n251807 , n251799 );
nand ( n251812 , n251810 , n251811 );
not ( n251813 , n248640 );
nand ( n251814 , n251813 , n243185 );
not ( n251815 , n251814 );
not ( n251816 , n250151 );
and ( n251817 , n251815 , n251816 );
and ( n251818 , n251814 , n250151 );
nor ( n251819 , n251817 , n251818 );
not ( n251820 , n251819 );
and ( n251821 , n251812 , n251820 );
not ( n251822 , n251812 );
and ( n251823 , n251822 , n251819 );
nor ( n251824 , n251821 , n251823 );
buf ( n251825 , n251824 );
not ( n251826 , n248596 );
nand ( n251827 , n251826 , n243076 );
not ( n251828 , n251827 );
not ( n251829 , n250215 );
and ( n251830 , n251828 , n251829 );
and ( n251831 , n251827 , n250215 );
nor ( n251832 , n251830 , n251831 );
not ( n251833 , n251832 );
nand ( n251834 , n243038 , n248578 );
not ( n251835 , n250192 );
and ( n251836 , n251834 , n251835 );
not ( n251837 , n251834 );
and ( n251838 , n251837 , n250192 );
nor ( n251839 , n251836 , n251838 );
not ( n251840 , n251839 );
and ( n251841 , n251833 , n251840 );
and ( n251842 , n251832 , n251839 );
nor ( n251843 , n251841 , n251842 );
buf ( n251844 , n251843 );
xor ( n251845 , n251825 , n251844 );
buf ( n251846 , n251845 );
and ( n251847 , n251792 , n251846 );
not ( n251848 , n251792 );
not ( n251849 , n251843 );
not ( n251850 , n251824 );
or ( n251851 , n251849 , n251850 );
not ( n251852 , n251824 );
not ( n251853 , n251843 );
nand ( n251854 , n251852 , n251853 );
nand ( n251855 , n251851 , n251854 );
buf ( n251856 , n251855 );
and ( n251857 , n251848 , n251856 );
nor ( n251858 , n251847 , n251857 );
not ( n251859 , n238635 );
nand ( n251860 , n251858 , n251859 );
or ( n251861 , n251787 , n251860 );
not ( n251862 , n222532 );
nor ( n251863 , n251858 , n251862 );
nand ( n251864 , n251863 , n251787 );
nand ( n251865 , n35431 , n207380 );
nand ( n251866 , n251861 , n251864 , n251865 );
buf ( n251867 , n251866 );
not ( n251868 , n48465 );
nand ( n251869 , n251868 , n48451 );
and ( n251870 , n251869 , n47584 );
not ( n251871 , n251869 );
not ( n251872 , n47584 );
and ( n251873 , n251871 , n251872 );
nor ( n251874 , n251870 , n251873 );
and ( n251875 , n251874 , n236781 );
not ( n251876 , n251874 );
and ( n251877 , n251876 , n234881 );
or ( n251878 , n251875 , n251877 );
and ( n251879 , n251878 , n234889 );
not ( n251880 , n251878 );
and ( n251881 , n251880 , n236789 );
nor ( n251882 , n251879 , n251881 );
nor ( n251883 , n251882 , n234021 );
not ( n251884 , n50130 );
not ( n251885 , n248967 );
or ( n251886 , n251884 , n251885 );
not ( n251887 , n50130 );
nand ( n251888 , n251887 , n249394 );
nand ( n251889 , n251886 , n251888 );
and ( n251890 , n251889 , n248972 );
not ( n251891 , n251889 );
and ( n251892 , n251891 , n248975 );
nor ( n251893 , n251890 , n251892 );
nand ( n251894 , n251883 , n251893 );
not ( n251895 , n251882 );
nor ( n251896 , n251895 , n250909 );
not ( n251897 , n246342 );
not ( n251898 , n251897 );
not ( n251899 , n44539 );
or ( n251900 , n251898 , n251899 );
or ( n251901 , n44539 , n251897 );
nand ( n251902 , n251900 , n251901 );
and ( n251903 , n251902 , n222525 );
not ( n251904 , n251902 );
and ( n251905 , n251904 , n44761 );
nor ( n251906 , n251903 , n251905 );
nor ( n251907 , n251893 , n251906 );
nand ( n251908 , n251896 , n251907 );
not ( n251909 , n251893 );
nor ( n251910 , n251909 , n54208 );
nand ( n251911 , n251910 , n251906 );
nand ( n251912 , n50615 , n26486 );
nand ( n251913 , n251894 , n251908 , n251911 , n251912 );
buf ( n251914 , n251913 );
buf ( n251915 , n38171 );
not ( n251916 , RI19aaf628_2458);
or ( n251917 , n25328 , n251916 );
not ( n251918 , RI19aa5218_2529);
or ( n251919 , n25335 , n251918 );
nand ( n251920 , n251917 , n251919 );
buf ( n251921 , n251920 );
not ( n251922 , n228567 );
not ( n251923 , n47126 );
nand ( n251924 , n228561 , n50788 );
not ( n251925 , n251924 );
or ( n251926 , n251923 , n251925 );
or ( n251927 , n251924 , n47126 );
nand ( n251928 , n251926 , n251927 );
not ( n251929 , n251928 );
not ( n251930 , n50917 );
nand ( n251931 , n251930 , n228665 );
not ( n251932 , n251931 );
not ( n251933 , n47041 );
and ( n251934 , n251932 , n251933 );
and ( n251935 , n251931 , n47041 );
nor ( n251936 , n251934 , n251935 );
not ( n251937 , n251936 );
or ( n251938 , n251929 , n251937 );
or ( n251939 , n251936 , n251928 );
nand ( n251940 , n251938 , n251939 );
nand ( n251941 , n50830 , n228577 );
and ( n251942 , n251941 , n47091 );
not ( n251943 , n251941 );
and ( n251944 , n251943 , n224851 );
nor ( n251945 , n251942 , n251944 );
not ( n251946 , n251945 );
and ( n251947 , n251940 , n251946 );
not ( n251948 , n251940 );
and ( n251949 , n251948 , n251945 );
nor ( n251950 , n251947 , n251949 );
not ( n251951 , n251950 );
not ( n251952 , n246008 );
not ( n251953 , n228638 );
nand ( n251954 , n251953 , n50889 );
not ( n251955 , n251954 );
buf ( n251956 , n47000 );
not ( n251957 , n251956 );
and ( n251958 , n251955 , n251957 );
and ( n251959 , n251954 , n251956 );
nor ( n251960 , n251958 , n251959 );
not ( n251961 , n251960 );
not ( n251962 , n251961 );
or ( n251963 , n251952 , n251962 );
nand ( n251964 , n246007 , n251960 );
nand ( n251965 , n251963 , n251964 );
not ( n251966 , n251965 );
not ( n251967 , n251966 );
and ( n251968 , n251951 , n251967 );
and ( n251969 , n251950 , n251966 );
nor ( n251970 , n251968 , n251969 );
not ( n251971 , n251970 );
or ( n251972 , n251922 , n251971 );
or ( n251973 , n228567 , n251970 );
nand ( n251974 , n251972 , n251973 );
not ( n251975 , n250899 );
and ( n251976 , n251974 , n251975 );
not ( n251977 , n251974 );
and ( n251978 , n251977 , n250899 );
nor ( n251979 , n251976 , n251978 );
not ( n251980 , n251979 );
not ( n251981 , n251980 );
not ( n251982 , n250576 );
not ( n251983 , n49236 );
not ( n251984 , n226975 );
nand ( n251985 , n251984 , n247037 );
not ( n251986 , n251985 );
or ( n251987 , n251983 , n251986 );
or ( n251988 , n251985 , n49236 );
nand ( n251989 , n251987 , n251988 );
not ( n251990 , n251989 );
not ( n251991 , n251990 );
and ( n251992 , n251982 , n251991 );
and ( n251993 , n250576 , n251990 );
nor ( n251994 , n251992 , n251993 );
nor ( n251995 , n49515 , n240225 );
and ( n251996 , n251995 , n49506 );
not ( n251997 , n251995 );
and ( n251998 , n251997 , n247168 );
nor ( n251999 , n251996 , n251998 );
not ( n252000 , n251999 );
not ( n252001 , n247132 );
nand ( n252002 , n49589 , n240281 );
not ( n252003 , n252002 );
or ( n252004 , n252001 , n252003 );
or ( n252005 , n252002 , n247132 );
nand ( n252006 , n252004 , n252005 );
not ( n252007 , n252006 );
not ( n252008 , n252007 );
nand ( n252009 , n49559 , n240178 );
not ( n252010 , n252009 );
not ( n252011 , n49549 );
and ( n252012 , n252010 , n252011 );
and ( n252013 , n252009 , n49549 );
nor ( n252014 , n252012 , n252013 );
not ( n252015 , n252014 );
not ( n252016 , n252015 );
or ( n252017 , n252008 , n252016 );
nand ( n252018 , n252014 , n252006 );
nand ( n252019 , n252017 , n252018 );
xor ( n252020 , n252000 , n252019 );
not ( n252021 , n240195 );
nand ( n252022 , n252021 , n49441 );
not ( n252023 , n252022 );
not ( n252024 , n247157 );
and ( n252025 , n252023 , n252024 );
and ( n252026 , n252022 , n247157 );
nor ( n252027 , n252025 , n252026 );
nand ( n252028 , n240257 , n49478 );
and ( n252029 , n252028 , n49467 );
not ( n252030 , n252028 );
and ( n252031 , n252030 , n49466 );
nor ( n252032 , n252029 , n252031 );
or ( n252033 , n252027 , n252032 );
nand ( n252034 , n252032 , n252027 );
nand ( n252035 , n252033 , n252034 );
xnor ( n252036 , n252020 , n252035 );
buf ( n252037 , n252036 );
and ( n252038 , n251994 , n252037 );
not ( n252039 , n251994 );
not ( n252040 , n252019 );
not ( n252041 , n252040 );
and ( n252042 , n252035 , n252000 );
not ( n252043 , n252035 );
and ( n252044 , n252043 , n251999 );
nor ( n252045 , n252042 , n252044 );
not ( n252046 , n252045 );
or ( n252047 , n252041 , n252046 );
not ( n252048 , n252045 );
not ( n252049 , n252040 );
nand ( n252050 , n252048 , n252049 );
nand ( n252051 , n252047 , n252050 );
buf ( n252052 , n252051 );
and ( n252053 , n252039 , n252052 );
nor ( n252054 , n252038 , n252053 );
not ( n252055 , n252054 );
or ( n252056 , n251981 , n252055 );
not ( n252057 , n250796 );
not ( n252058 , n251154 );
or ( n252059 , n252057 , n252058 );
not ( n252060 , n250796 );
nand ( n252061 , n252060 , n251253 );
nand ( n252062 , n252059 , n252061 );
and ( n252063 , n252062 , n251313 );
not ( n252064 , n252062 );
and ( n252065 , n252064 , n251299 );
nor ( n252066 , n252063 , n252065 );
not ( n252067 , n252066 );
nor ( n252068 , n252067 , n50944 );
nand ( n252069 , n252056 , n252068 );
buf ( n252070 , n35427 );
nor ( n252071 , n251979 , n252070 );
nand ( n252072 , n252054 , n252071 , n252067 );
nand ( n252073 , n31577 , n32849 );
nand ( n252074 , n252069 , n252072 , n252073 );
buf ( n252075 , n252074 );
buf ( n252076 , n31822 );
buf ( n252077 , n55601 );
not ( n252078 , n252077 );
not ( n252079 , n235016 );
or ( n252080 , n252078 , n252079 );
not ( n252081 , n235016 );
not ( n252082 , n252081 );
or ( n252083 , n252082 , n252077 );
nand ( n252084 , n252080 , n252083 );
and ( n252085 , n252084 , n235022 );
not ( n252086 , n252084 );
and ( n252087 , n252086 , n235019 );
nor ( n252088 , n252085 , n252087 );
nand ( n252089 , n252088 , n250929 );
not ( n252090 , n237693 );
not ( n252091 , n233997 );
or ( n252092 , n252090 , n252091 );
not ( n252093 , n237693 );
nand ( n252094 , n252093 , n44176 );
nand ( n252095 , n252092 , n252094 );
and ( n252096 , n252095 , n44316 );
not ( n252097 , n252095 );
and ( n252098 , n252097 , n44325 );
nor ( n252099 , n252096 , n252098 );
not ( n252100 , n252099 );
not ( n252101 , n251425 );
not ( n252102 , n224967 );
nand ( n252103 , n47217 , n40595 );
and ( n252104 , n252103 , n224980 );
not ( n252105 , n252103 );
and ( n252106 , n252105 , n40491 );
nor ( n252107 , n252104 , n252106 );
not ( n252108 , n252107 );
or ( n252109 , n252102 , n252108 );
or ( n252110 , n252107 , n224967 );
nand ( n252111 , n252109 , n252110 );
not ( n252112 , n47245 );
nand ( n252113 , n252112 , n218511 );
buf ( n252114 , n47235 );
xnor ( n252115 , n252113 , n252114 );
xnor ( n252116 , n252111 , n252115 );
not ( n252117 , n244640 );
nand ( n252118 , n47274 , n40900 );
not ( n252119 , n252118 );
not ( n252120 , n47263 );
and ( n252121 , n252119 , n252120 );
and ( n252122 , n252118 , n47263 );
nor ( n252123 , n252121 , n252122 );
not ( n252124 , n252123 );
and ( n252125 , n252117 , n252124 );
and ( n252126 , n244640 , n252123 );
nor ( n252127 , n252125 , n252126 );
and ( n252128 , n252116 , n252127 );
not ( n252129 , n252116 );
not ( n252130 , n252127 );
and ( n252131 , n252129 , n252130 );
nor ( n252132 , n252128 , n252131 );
not ( n252133 , n252132 );
or ( n252134 , n252101 , n252133 );
not ( n252135 , n251425 );
and ( n252136 , n252116 , n252130 );
not ( n252137 , n252116 );
and ( n252138 , n252137 , n252127 );
nor ( n252139 , n252136 , n252138 );
nand ( n252140 , n252135 , n252139 );
nand ( n252141 , n252134 , n252140 );
not ( n252142 , n42482 );
not ( n252143 , n42664 );
nand ( n252144 , n252143 , n41106 );
and ( n252145 , n252144 , n42684 );
not ( n252146 , n252144 );
and ( n252147 , n252146 , n42683 );
nor ( n252148 , n252145 , n252147 );
not ( n252149 , n252148 );
not ( n252150 , n252149 );
or ( n252151 , n252142 , n252150 );
nand ( n252152 , n252148 , n42481 );
nand ( n252153 , n252151 , n252152 );
not ( n252154 , n252153 );
nand ( n252155 , n40952 , n42641 );
and ( n252156 , n252155 , n42630 );
not ( n252157 , n252155 );
and ( n252158 , n252157 , n42629 );
nor ( n252159 , n252156 , n252158 );
nand ( n252160 , n54231 , n41084 );
not ( n252161 , n252160 );
not ( n252162 , n42523 );
and ( n252163 , n252161 , n252162 );
and ( n252164 , n252160 , n42523 );
nor ( n252165 , n252163 , n252164 );
or ( n252166 , n252159 , n252165 );
nand ( n252167 , n252165 , n252159 );
nand ( n252168 , n252166 , n252167 );
nand ( n252169 , n40974 , n54220 );
not ( n252170 , n252169 );
not ( n252171 , n237599 );
and ( n252172 , n252170 , n252171 );
and ( n252173 , n252169 , n237599 );
nor ( n252174 , n252172 , n252173 );
and ( n252175 , n252168 , n252174 );
not ( n252176 , n252168 );
not ( n252177 , n252174 );
and ( n252178 , n252176 , n252177 );
nor ( n252179 , n252175 , n252178 );
not ( n252180 , n252179 );
or ( n252181 , n252154 , n252180 );
not ( n252182 , n252153 );
not ( n252183 , n252179 );
nand ( n252184 , n252182 , n252183 );
nand ( n252185 , n252181 , n252184 );
buf ( n252186 , n252185 );
and ( n252187 , n252141 , n252186 );
not ( n252188 , n252141 );
and ( n252189 , n252153 , n252179 );
not ( n252190 , n252153 );
and ( n252191 , n252190 , n252183 );
nor ( n252192 , n252189 , n252191 );
not ( n252193 , n252192 );
not ( n252194 , n252193 );
and ( n252195 , n252188 , n252194 );
nor ( n252196 , n252187 , n252195 );
not ( n252197 , n252196 );
nand ( n252198 , n252100 , n252197 );
or ( n252199 , n252089 , n252198 );
not ( n252200 , n239934 );
nor ( n252201 , n252088 , n252200 );
nand ( n252202 , n252201 , n252198 );
nand ( n252203 , n247744 , n36386 );
nand ( n252204 , n252199 , n252202 , n252203 );
buf ( n252205 , n252204 );
not ( n252206 , RI19ac3290_2305);
or ( n252207 , n226819 , n252206 );
not ( n252208 , RI19abaa28_2376);
or ( n252209 , n226822 , n252208 );
nand ( n252210 , n252207 , n252209 );
buf ( n252211 , n252210 );
buf ( n252212 , n26086 );
buf ( n252213 , RI19ad0700_2208);
buf ( n252214 , n252213 );
not ( n252215 , n235661 );
not ( n252216 , n238461 );
or ( n252217 , n252215 , n252216 );
not ( n252218 , n235661 );
nand ( n252219 , n252218 , n238470 );
nand ( n252220 , n252217 , n252219 );
and ( n252221 , n252220 , n238473 );
not ( n252222 , n252220 );
and ( n252223 , n252222 , n238476 );
nor ( n252224 , n252221 , n252223 );
not ( n252225 , n252224 );
not ( n252226 , n245277 );
not ( n252227 , n242068 );
or ( n252228 , n252226 , n252227 );
not ( n252229 , n245277 );
and ( n252230 , n242035 , n241999 );
not ( n252231 , n242035 );
not ( n252232 , n241999 );
and ( n252233 , n252231 , n252232 );
nor ( n252234 , n252230 , n252233 );
xor ( n252235 , n242067 , n252234 );
not ( n252236 , n252235 );
nand ( n252237 , n252229 , n252236 );
nand ( n252238 , n252228 , n252237 );
buf ( n252239 , n235366 );
and ( n252240 , n252238 , n252239 );
not ( n252241 , n252238 );
buf ( n252242 , n235357 );
and ( n252243 , n252241 , n252242 );
nor ( n252244 , n252240 , n252243 );
not ( n252245 , n252244 );
nand ( n252246 , n252225 , n252245 );
not ( n252247 , n220944 );
not ( n252248 , n252247 );
not ( n252249 , n244453 );
or ( n252250 , n252248 , n252249 );
or ( n252251 , n244453 , n252247 );
nand ( n252252 , n252250 , n252251 );
and ( n252253 , n252252 , n249789 );
not ( n252254 , n252252 );
and ( n252255 , n252254 , n249792 );
nor ( n252256 , n252253 , n252255 );
not ( n252257 , n252256 );
buf ( n252258 , n233971 );
not ( n252259 , n252258 );
nand ( n252260 , n252257 , n252259 );
or ( n252261 , n252246 , n252260 );
not ( n252262 , n252257 );
not ( n252263 , n252225 );
or ( n252264 , n252262 , n252263 );
nor ( n252265 , n252245 , n234440 );
nand ( n252266 , n252264 , n252265 );
nand ( n252267 , n49054 , n31881 );
nand ( n252268 , n252261 , n252266 , n252267 );
buf ( n252269 , n252268 );
not ( n252270 , n243984 );
not ( n252271 , n252270 );
not ( n252272 , n250265 );
nand ( n252273 , n44955 , n243935 );
not ( n252274 , n252273 );
not ( n252275 , n243923 );
and ( n252276 , n252274 , n252275 );
and ( n252277 , n252273 , n243923 );
nor ( n252278 , n252276 , n252277 );
not ( n252279 , n252278 );
or ( n252280 , n252272 , n252279 );
or ( n252281 , n250265 , n252278 );
nand ( n252282 , n252280 , n252281 );
not ( n252283 , n243904 );
nand ( n252284 , n252283 , n44826 );
not ( n252285 , n252284 );
buf ( n252286 , n243892 );
not ( n252287 , n252286 );
and ( n252288 , n252285 , n252287 );
and ( n252289 , n252284 , n252286 );
nor ( n252290 , n252288 , n252289 );
and ( n252291 , n252282 , n252290 );
not ( n252292 , n252282 );
not ( n252293 , n252290 );
and ( n252294 , n252292 , n252293 );
nor ( n252295 , n252291 , n252294 );
not ( n252296 , n252295 );
not ( n252297 , n243828 );
nand ( n252298 , n45011 , n252297 );
xor ( n252299 , n252298 , n44800 );
not ( n252300 , n252299 );
not ( n252301 , n237958 );
nand ( n252302 , n44969 , n243846 );
not ( n252303 , n252302 );
or ( n252304 , n252301 , n252303 );
not ( n252305 , n243847 );
nand ( n252306 , n252305 , n44969 );
or ( n252307 , n252306 , n237958 );
nand ( n252308 , n252304 , n252307 );
not ( n252309 , n252308 );
or ( n252310 , n252300 , n252309 );
or ( n252311 , n252308 , n252299 );
nand ( n252312 , n252310 , n252311 );
not ( n252313 , n252312 );
and ( n252314 , n252296 , n252313 );
and ( n252315 , n252295 , n252312 );
nor ( n252316 , n252314 , n252315 );
buf ( n252317 , n252316 );
not ( n252318 , n252317 );
not ( n252319 , n252318 );
or ( n252320 , n252271 , n252319 );
not ( n252321 , n252317 );
or ( n252322 , n252321 , n252270 );
nand ( n252323 , n252320 , n252322 );
buf ( n252324 , n54926 );
and ( n252325 , n252323 , n252324 );
not ( n252326 , n252323 );
buf ( n252327 , n54917 );
and ( n252328 , n252326 , n252327 );
nor ( n252329 , n252325 , n252328 );
not ( n252330 , n233921 );
not ( n252331 , n244336 );
or ( n252332 , n252330 , n252331 );
not ( n252333 , n233921 );
nand ( n252334 , n252333 , n244346 );
nand ( n252335 , n252332 , n252334 );
and ( n252336 , n252335 , n244472 );
not ( n252337 , n252335 );
and ( n252338 , n252337 , n244475 );
nor ( n252339 , n252336 , n252338 );
not ( n252340 , n252339 );
nand ( n252341 , n252329 , n252340 );
not ( n252342 , n230807 );
not ( n252343 , n42149 );
or ( n252344 , n252342 , n252343 );
nand ( n252345 , n42156 , n53042 );
nand ( n252346 , n252344 , n252345 );
not ( n252347 , n252346 );
not ( n252348 , n42436 );
not ( n252349 , n252348 );
and ( n252350 , n252347 , n252349 );
and ( n252351 , n252346 , n220201 );
nor ( n252352 , n252350 , n252351 );
nand ( n252353 , n252352 , n241459 );
or ( n252354 , n252341 , n252353 );
not ( n252355 , n252352 );
not ( n252356 , n252329 );
or ( n252357 , n252355 , n252356 );
buf ( n252358 , n233971 );
nor ( n252359 , n252340 , n252358 );
nand ( n252360 , n252357 , n252359 );
nand ( n252361 , n46083 , n40150 );
nand ( n252362 , n252354 , n252360 , n252361 );
buf ( n252363 , n252362 );
not ( n252364 , RI19a82f88_2773);
or ( n252365 , n226819 , n252364 );
not ( n252366 , RI19ac81c8_2269);
or ( n252367 , n25336 , n252366 );
nand ( n252368 , n252365 , n252367 );
buf ( n252369 , n252368 );
not ( n252370 , n207202 );
not ( n252371 , n234453 );
or ( n252372 , n252370 , n252371 );
not ( n252373 , n247385 );
not ( n252374 , n240508 );
or ( n252375 , n252373 , n252374 );
not ( n252376 , n247385 );
nand ( n252377 , n252376 , n240503 );
nand ( n252378 , n252375 , n252377 );
and ( n252379 , n252378 , n246173 );
not ( n252380 , n252378 );
and ( n252381 , n252380 , n246168 );
nor ( n252382 , n252379 , n252381 );
not ( n252383 , n252382 );
buf ( n252384 , n37145 );
not ( n252385 , n252384 );
not ( n252386 , n240799 );
or ( n252387 , n252385 , n252386 );
or ( n252388 , n240799 , n252384 );
nand ( n252389 , n252387 , n252388 );
nand ( n252390 , n240877 , n37541 );
not ( n252391 , n250640 );
and ( n252392 , n252390 , n252391 );
not ( n252393 , n252390 );
and ( n252394 , n252393 , n250640 );
nor ( n252395 , n252392 , n252394 );
not ( n252396 , n252395 );
nand ( n252397 , n37585 , n37654 );
not ( n252398 , n252397 );
not ( n252399 , n250626 );
and ( n252400 , n252398 , n252399 );
and ( n252401 , n252397 , n250626 );
nor ( n252402 , n252400 , n252401 );
not ( n252403 , n252402 );
and ( n252404 , n252396 , n252403 );
and ( n252405 , n252395 , n252402 );
nor ( n252406 , n252404 , n252405 );
not ( n252407 , n252406 );
not ( n252408 , n252407 );
nand ( n252409 , n37692 , n240856 );
and ( n252410 , n252409 , n250658 );
not ( n252411 , n252409 );
and ( n252412 , n252411 , n250659 );
nor ( n252413 , n252410 , n252412 );
not ( n252414 , n252413 );
not ( n252415 , n252414 );
or ( n252416 , n252408 , n252415 );
nand ( n252417 , n252406 , n252413 );
nand ( n252418 , n252416 , n252417 );
nand ( n252419 , n240911 , n37474 );
not ( n252420 , n252419 );
not ( n252421 , n240834 );
and ( n252422 , n252420 , n252421 );
and ( n252423 , n252419 , n240834 );
nor ( n252424 , n252422 , n252423 );
not ( n252425 , n252424 );
not ( n252426 , n37299 );
nand ( n252427 , n252426 , n37358 );
not ( n252428 , n244359 );
and ( n252429 , n252427 , n252428 );
not ( n252430 , n252427 );
and ( n252431 , n252430 , n244359 );
nor ( n252432 , n252429 , n252431 );
not ( n252433 , n252432 );
or ( n252434 , n252425 , n252433 );
not ( n252435 , n252424 );
not ( n252436 , n252432 );
nand ( n252437 , n252435 , n252436 );
nand ( n252438 , n252434 , n252437 );
and ( n252439 , n252418 , n252438 );
not ( n252440 , n252418 );
not ( n252441 , n252438 );
and ( n252442 , n252440 , n252441 );
nor ( n252443 , n252439 , n252442 );
not ( n252444 , n252443 );
and ( n252445 , n252389 , n252444 );
not ( n252446 , n252389 );
not ( n252447 , n252444 );
and ( n252448 , n252446 , n252447 );
nor ( n252449 , n252445 , n252448 );
nand ( n252450 , n252383 , n252449 );
and ( n252451 , n204519 , n245840 , n245003 );
not ( n252452 , n252451 );
not ( n252453 , n245844 );
not ( n252454 , n39434 );
or ( n252455 , n252453 , n252454 );
not ( n252456 , n245844 );
nand ( n252457 , n252456 , n39444 );
nand ( n252458 , n252455 , n252457 );
and ( n252459 , n252458 , n250255 );
not ( n252460 , n252458 );
and ( n252461 , n252460 , n248795 );
nor ( n252462 , n252459 , n252461 );
not ( n252463 , n252462 );
or ( n252464 , n252452 , n252463 );
or ( n252465 , n252462 , n252451 );
nand ( n252466 , n252464 , n252465 );
and ( n252467 , n252450 , n252466 );
not ( n252468 , n252450 );
not ( n252469 , n252466 );
and ( n252470 , n252468 , n252469 );
nor ( n252471 , n252467 , n252470 );
or ( n252472 , n252471 , n52445 );
nand ( n252473 , n252372 , n252472 );
buf ( n252474 , n252473 );
not ( n252475 , n240575 );
nand ( n252476 , n252475 , n240328 );
not ( n252477 , n252476 );
buf ( n252478 , n240585 );
not ( n252479 , n252478 );
and ( n252480 , n252477 , n252479 );
and ( n252481 , n252476 , n252478 );
nor ( n252482 , n252480 , n252481 );
not ( n252483 , n252482 );
not ( n252484 , n240684 );
or ( n252485 , n252483 , n252484 );
not ( n252486 , n252482 );
nand ( n252487 , n252486 , n240676 );
nand ( n252488 , n252485 , n252487 );
and ( n252489 , n252488 , n240801 );
not ( n252490 , n252488 );
and ( n252491 , n252490 , n240811 );
nor ( n252492 , n252489 , n252491 );
not ( n252493 , n252492 );
not ( n252494 , n43568 );
not ( n252495 , n242270 );
or ( n252496 , n252494 , n252495 );
not ( n252497 , n43568 );
not ( n252498 , n242243 );
not ( n252499 , n242266 );
not ( n252500 , n252499 );
or ( n252501 , n252498 , n252500 );
nand ( n252502 , n242244 , n242266 );
nand ( n252503 , n252501 , n252502 );
nand ( n252504 , n252497 , n252503 );
nand ( n252505 , n252496 , n252504 );
nand ( n252506 , n221652 , n43879 );
not ( n252507 , n252506 );
not ( n252508 , n235107 );
and ( n252509 , n252507 , n252508 );
and ( n252510 , n252506 , n235107 );
nor ( n252511 , n252509 , n252510 );
not ( n252512 , n252511 );
nand ( n252513 , n43860 , n43827 );
and ( n252514 , n252513 , n249311 );
not ( n252515 , n252513 );
and ( n252516 , n252515 , n235143 );
nor ( n252517 , n252514 , n252516 );
not ( n252518 , n252517 );
or ( n252519 , n252512 , n252518 );
or ( n252520 , n252517 , n252511 );
nand ( n252521 , n252519 , n252520 );
not ( n252522 , n221702 );
nand ( n252523 , n252522 , n248415 );
and ( n252524 , n252523 , n235082 );
not ( n252525 , n252523 );
and ( n252526 , n252525 , n235091 );
nor ( n252527 , n252524 , n252526 );
and ( n252528 , n252521 , n252527 );
not ( n252529 , n252521 );
not ( n252530 , n252527 );
and ( n252531 , n252529 , n252530 );
nor ( n252532 , n252528 , n252531 );
nand ( n252533 , n43736 , n43748 );
and ( n252534 , n252533 , n249345 );
not ( n252535 , n252533 );
and ( n252536 , n252535 , n235168 );
nor ( n252537 , n252534 , n252536 );
not ( n252538 , n252537 );
and ( n252539 , n43779 , n221566 );
and ( n252540 , n252539 , n249336 );
not ( n252541 , n252539 );
and ( n252542 , n252541 , n235176 );
nor ( n252543 , n252540 , n252542 );
not ( n252544 , n252543 );
and ( n252545 , n252538 , n252544 );
and ( n252546 , n252537 , n252543 );
nor ( n252547 , n252545 , n252546 );
and ( n252548 , n252532 , n252547 );
not ( n252549 , n252532 );
not ( n252550 , n252547 );
and ( n252551 , n252549 , n252550 );
nor ( n252552 , n252548 , n252551 );
buf ( n252553 , n252552 );
and ( n252554 , n252505 , n252553 );
not ( n252555 , n252505 );
not ( n252556 , n252547 );
not ( n252557 , n252532 );
or ( n252558 , n252556 , n252557 );
not ( n252559 , n252532 );
nand ( n252560 , n252559 , n252550 );
nand ( n252561 , n252558 , n252560 );
buf ( n252562 , n252561 );
and ( n252563 , n252555 , n252562 );
nor ( n252564 , n252554 , n252563 );
nand ( n252565 , n252493 , n252564 );
not ( n252566 , n51989 );
not ( n252567 , n245201 );
not ( n252568 , n252567 );
or ( n252569 , n252566 , n252568 );
nand ( n252570 , n236385 , n229749 );
nand ( n252571 , n252569 , n252570 );
and ( n252572 , n245211 , n252571 );
not ( n252573 , n245211 );
not ( n252574 , n252571 );
and ( n252575 , n252573 , n252574 );
nor ( n252576 , n252572 , n252575 );
nor ( n252577 , n252576 , n55146 );
not ( n252578 , n252577 );
or ( n252579 , n252565 , n252578 );
not ( n252580 , n252576 );
nor ( n252581 , n252580 , n31572 );
nand ( n252582 , n252565 , n252581 );
nand ( n252583 , n35431 , n40828 );
nand ( n252584 , n252579 , n252582 , n252583 );
buf ( n252585 , n252584 );
not ( n252586 , n208229 );
not ( n252587 , n245943 );
or ( n252588 , n252586 , n252587 );
not ( n252589 , n240360 );
nand ( n252590 , n240423 , n240409 );
and ( n252591 , n252590 , n240615 );
not ( n252592 , n252590 );
and ( n252593 , n252592 , n240614 );
nor ( n252594 , n252591 , n252593 );
buf ( n252595 , n252594 );
not ( n252596 , n252595 );
not ( n252597 , n240388 );
nand ( n252598 , n252597 , n247352 );
and ( n252599 , n252598 , n240558 );
not ( n252600 , n252598 );
and ( n252601 , n252600 , n240557 );
nor ( n252602 , n252599 , n252601 );
not ( n252603 , n252602 );
not ( n252604 , n252603 );
or ( n252605 , n252596 , n252604 );
not ( n252606 , n252594 );
nand ( n252607 , n252606 , n252602 );
nand ( n252608 , n252605 , n252607 );
not ( n252609 , n240445 );
nand ( n252610 , n252609 , n240455 );
not ( n252611 , n252610 );
not ( n252612 , n240659 );
and ( n252613 , n252611 , n252612 );
and ( n252614 , n252610 , n240659 );
nor ( n252615 , n252613 , n252614 );
buf ( n252616 , n252615 );
not ( n252617 , n252616 );
and ( n252618 , n252608 , n252617 );
not ( n252619 , n252608 );
and ( n252620 , n252619 , n252616 );
nor ( n252621 , n252618 , n252620 );
not ( n252622 , n252475 );
nor ( n252623 , n240328 , n240353 );
not ( n252624 , n252623 );
and ( n252625 , n252622 , n252624 );
and ( n252626 , n252475 , n252623 );
nor ( n252627 , n252625 , n252626 );
not ( n252628 , n252627 );
not ( n252629 , n240489 );
nand ( n252630 , n252629 , n240483 );
and ( n252631 , n252630 , n240649 );
not ( n252632 , n252630 );
and ( n252633 , n252632 , n240650 );
nor ( n252634 , n252631 , n252633 );
not ( n252635 , n252634 );
or ( n252636 , n252628 , n252635 );
or ( n252637 , n252634 , n252627 );
nand ( n252638 , n252636 , n252637 );
buf ( n252639 , n252638 );
not ( n252640 , n252639 );
and ( n252641 , n252621 , n252640 );
not ( n252642 , n252621 );
and ( n252643 , n252642 , n252639 );
nor ( n252644 , n252641 , n252643 );
not ( n252645 , n252644 );
or ( n252646 , n252589 , n252645 );
not ( n252647 , n240360 );
xor ( n252648 , n252615 , n252608 );
xnor ( n252649 , n252648 , n252638 );
nand ( n252650 , n252647 , n252649 );
nand ( n252651 , n252646 , n252650 );
buf ( n252652 , n245602 );
and ( n252653 , n252651 , n252652 );
not ( n252654 , n252651 );
not ( n252655 , n245611 );
not ( n252656 , n252655 );
and ( n252657 , n252654 , n252656 );
nor ( n252658 , n252653 , n252657 );
not ( n252659 , n252658 );
nand ( n252660 , n250125 , n250236 );
and ( n252661 , n252659 , n252660 );
not ( n252662 , n252659 );
not ( n252663 , n252660 );
and ( n252664 , n252662 , n252663 );
nor ( n252665 , n252661 , n252664 );
or ( n252666 , n252665 , n240080 );
nand ( n252667 , n252588 , n252666 );
buf ( n252668 , n252667 );
not ( n252669 , n47487 );
not ( n252670 , n250896 );
or ( n252671 , n252669 , n252670 );
or ( n252672 , n251975 , n47487 );
nand ( n252673 , n252671 , n252672 );
and ( n252674 , n252673 , n250903 );
not ( n252675 , n252673 );
and ( n252676 , n252675 , n250906 );
nor ( n252677 , n252674 , n252676 );
not ( n252678 , n252677 );
not ( n252679 , n205649 );
nor ( n252680 , n252678 , n252679 );
not ( n252681 , n252680 );
not ( n252682 , n247895 );
not ( n252683 , n252682 );
not ( n252684 , n239853 );
or ( n252685 , n252683 , n252684 );
not ( n252686 , n239853 );
nand ( n252687 , n252686 , n247895 );
nand ( n252688 , n252685 , n252687 );
and ( n252689 , n252688 , n239930 );
not ( n252690 , n252688 );
and ( n252691 , n252690 , n239922 );
nor ( n252692 , n252689 , n252691 );
not ( n252693 , n244020 );
not ( n252694 , n54917 );
or ( n252695 , n252693 , n252694 );
not ( n252696 , n244020 );
nand ( n252697 , n252696 , n54926 );
nand ( n252698 , n252695 , n252697 );
and ( n252699 , n252698 , n240073 );
not ( n252700 , n252698 );
and ( n252701 , n252700 , n55068 );
nor ( n252702 , n252699 , n252701 );
not ( n252703 , n252702 );
nand ( n252704 , n252692 , n252703 );
or ( n252705 , n252681 , n252704 );
not ( n252706 , n252703 );
not ( n252707 , n252677 );
or ( n252708 , n252706 , n252707 );
nor ( n252709 , n252692 , n40465 );
nand ( n252710 , n252708 , n252709 );
buf ( n252711 , n35431 );
nand ( n252712 , n252711 , n30822 );
nand ( n252713 , n252705 , n252710 , n252712 );
buf ( n252714 , n252713 );
not ( n252715 , n247332 );
not ( n252716 , n252715 );
not ( n252717 , n251372 );
or ( n252718 , n252716 , n252717 );
or ( n252719 , n251372 , n252715 );
nand ( n252720 , n252718 , n252719 );
not ( n252721 , n252720 );
not ( n252722 , n250682 );
and ( n252723 , n252721 , n252722 );
and ( n252724 , n252720 , n250682 );
nor ( n252725 , n252723 , n252724 );
nand ( n252726 , n252725 , n252259 );
not ( n252727 , n245785 );
not ( n252728 , n52756 );
or ( n252729 , n252727 , n252728 );
not ( n252730 , n245785 );
nand ( n252731 , n252730 , n245264 );
nand ( n252732 , n252729 , n252731 );
buf ( n252733 , n251253 );
and ( n252734 , n252732 , n252733 );
not ( n252735 , n252732 );
and ( n252736 , n252735 , n251156 );
nor ( n252737 , n252734 , n252736 );
not ( n252738 , n252737 );
not ( n252739 , n252165 );
not ( n252740 , n252739 );
not ( n252741 , n220460 );
or ( n252742 , n252740 , n252741 );
not ( n252743 , n252739 );
nand ( n252744 , n252743 , n220467 );
nand ( n252745 , n252742 , n252744 );
and ( n252746 , n252745 , n43006 );
not ( n252747 , n252745 );
and ( n252748 , n252747 , n43011 );
nor ( n252749 , n252746 , n252748 );
nand ( n252750 , n252738 , n252749 );
or ( n252751 , n252726 , n252750 );
not ( n252752 , n252749 );
not ( n252753 , n252725 );
or ( n252754 , n252752 , n252753 );
nor ( n252755 , n252738 , n234440 );
nand ( n252756 , n252754 , n252755 );
nand ( n252757 , n252711 , n36129 );
nand ( n252758 , n252751 , n252756 , n252757 );
buf ( n252759 , n252758 );
not ( n252760 , n204972 );
not ( n252761 , n245221 );
or ( n252762 , n252760 , n252761 );
not ( n252763 , n53440 );
not ( n252764 , n252763 );
not ( n252765 , n250359 );
or ( n252766 , n252764 , n252765 );
not ( n252767 , n252763 );
nand ( n252768 , n252767 , n250366 );
nand ( n252769 , n252766 , n252768 );
and ( n252770 , n252769 , n250374 );
not ( n252771 , n252769 );
and ( n252772 , n252771 , n250371 );
nor ( n252773 , n252770 , n252772 );
not ( n252774 , n252773 );
not ( n252775 , n47108 );
not ( n252776 , n251953 );
nand ( n252777 , n245625 , n47021 );
not ( n252778 , n252777 );
or ( n252779 , n252776 , n252778 );
or ( n252780 , n252777 , n251953 );
nand ( n252781 , n252779 , n252780 );
not ( n252782 , n252781 );
not ( n252783 , n46983 );
nand ( n252784 , n252783 , n245967 );
not ( n252785 , n252784 );
not ( n252786 , n228611 );
not ( n252787 , n252786 );
and ( n252788 , n252785 , n252787 );
and ( n252789 , n252784 , n252786 );
nor ( n252790 , n252788 , n252789 );
not ( n252791 , n252790 );
or ( n252792 , n252782 , n252791 );
or ( n252793 , n252790 , n252781 );
nand ( n252794 , n252792 , n252793 );
nand ( n252795 , n47057 , n47052 );
and ( n252796 , n252795 , n228666 );
not ( n252797 , n252795 );
and ( n252798 , n252797 , n228665 );
nor ( n252799 , n252796 , n252798 );
and ( n252800 , n252794 , n252799 );
not ( n252801 , n252794 );
not ( n252802 , n252799 );
and ( n252803 , n252801 , n252802 );
nor ( n252804 , n252800 , n252803 );
not ( n252805 , n252804 );
not ( n252806 , n47139 );
nand ( n252807 , n252806 , n245978 );
not ( n252808 , n252807 );
not ( n252809 , n228561 );
and ( n252810 , n252808 , n252809 );
and ( n252811 , n252807 , n228561 );
nor ( n252812 , n252810 , n252811 );
and ( n252813 , n244522 , n252812 );
not ( n252814 , n244522 );
not ( n252815 , n252812 );
and ( n252816 , n252814 , n252815 );
nor ( n252817 , n252813 , n252816 );
not ( n252818 , n252817 );
and ( n252819 , n252805 , n252818 );
not ( n252820 , n252805 );
not ( n252821 , n252818 );
and ( n252822 , n252820 , n252821 );
nor ( n252823 , n252819 , n252822 );
not ( n252824 , n252823 );
or ( n252825 , n252775 , n252824 );
not ( n252826 , n47108 );
not ( n252827 , n252817 );
not ( n252828 , n252804 );
or ( n252829 , n252827 , n252828 );
nand ( n252830 , n252805 , n252818 );
nand ( n252831 , n252829 , n252830 );
nand ( n252832 , n252826 , n252831 );
nand ( n252833 , n252825 , n252832 );
buf ( n252834 , n241448 );
and ( n252835 , n252833 , n252834 );
not ( n252836 , n252833 );
not ( n252837 , n252834 );
and ( n252838 , n252836 , n252837 );
nor ( n252839 , n252835 , n252838 );
not ( n252840 , n252839 );
nand ( n252841 , n252774 , n252840 );
not ( n252842 , n223152 );
not ( n252843 , n248161 );
not ( n252844 , n252843 );
or ( n252845 , n252842 , n252844 );
not ( n252846 , n223152 );
nand ( n252847 , n252846 , n248161 );
nand ( n252848 , n252845 , n252847 );
and ( n252849 , n252848 , n248211 );
not ( n252850 , n252848 );
and ( n252851 , n252850 , n248220 );
nor ( n252852 , n252849 , n252851 );
not ( n252853 , n252852 );
and ( n252854 , n252841 , n252853 );
not ( n252855 , n252841 );
and ( n252856 , n252855 , n252852 );
nor ( n252857 , n252854 , n252856 );
not ( n252858 , n237358 );
not ( n252859 , n252858 );
or ( n252860 , n252857 , n252859 );
nand ( n252861 , n252762 , n252860 );
buf ( n252862 , n252861 );
not ( n252863 , n244173 );
not ( n252864 , n234803 );
or ( n252865 , n252863 , n252864 );
or ( n252866 , n234803 , n244173 );
nand ( n252867 , n252865 , n252866 );
and ( n252868 , n252867 , n250398 );
not ( n252869 , n252867 );
and ( n252870 , n252869 , n250395 );
nor ( n252871 , n252868 , n252870 );
buf ( n252872 , n236795 );
not ( n252873 , n252872 );
nand ( n252874 , n252871 , n252873 );
not ( n252875 , n239249 );
not ( n252876 , n248755 );
or ( n252877 , n252875 , n252876 );
not ( n252878 , n239249 );
nand ( n252879 , n252878 , n248762 );
nand ( n252880 , n252877 , n252879 );
nand ( n252881 , n55249 , n239330 );
not ( n252882 , n252881 );
not ( n252883 , n41401 );
and ( n252884 , n252882 , n252883 );
and ( n252885 , n252881 , n41401 );
nor ( n252886 , n252884 , n252885 );
not ( n252887 , n252886 );
not ( n252888 , n252887 );
nand ( n252889 , n239314 , n55230 );
and ( n252890 , n252889 , n241016 );
not ( n252891 , n252889 );
and ( n252892 , n252891 , n219219 );
nor ( n252893 , n252890 , n252892 );
not ( n252894 , n252893 );
not ( n252895 , n252894 );
or ( n252896 , n252888 , n252895 );
nand ( n252897 , n252893 , n252886 );
nand ( n252898 , n252896 , n252897 );
xor ( n252899 , n241004 , n252898 );
not ( n252900 , n239353 );
nand ( n252901 , n252900 , n232953 );
not ( n252902 , n252901 );
not ( n252903 , n41606 );
and ( n252904 , n252902 , n252903 );
and ( n252905 , n252901 , n41606 );
nor ( n252906 , n252904 , n252905 );
not ( n252907 , n252906 );
nand ( n252908 , n239368 , n55172 );
and ( n252909 , n252908 , n241036 );
not ( n252910 , n252908 );
and ( n252911 , n252910 , n241035 );
nor ( n252912 , n252909 , n252911 );
not ( n252913 , n252912 );
or ( n252914 , n252907 , n252913 );
or ( n252915 , n252912 , n252906 );
nand ( n252916 , n252914 , n252915 );
xnor ( n252917 , n252899 , n252916 );
buf ( n252918 , n252917 );
not ( n252919 , n252918 );
and ( n252920 , n252880 , n252919 );
not ( n252921 , n252880 );
not ( n252922 , n252917 );
buf ( n252923 , n252922 );
not ( n252924 , n252923 );
and ( n252925 , n252921 , n252924 );
nor ( n252926 , n252920 , n252925 );
not ( n252927 , n249181 );
not ( n252928 , n244776 );
or ( n252929 , n252927 , n252928 );
not ( n252930 , n249181 );
nand ( n252931 , n252930 , n244768 );
nand ( n252932 , n252929 , n252931 );
not ( n252933 , n239715 );
not ( n252934 , n252933 );
and ( n252935 , n252932 , n252934 );
not ( n252936 , n252932 );
and ( n252937 , n252936 , n249059 );
nor ( n252938 , n252935 , n252937 );
not ( n252939 , n252938 );
nand ( n252940 , n252926 , n252939 );
or ( n252941 , n252874 , n252940 );
not ( n252942 , n252926 );
not ( n252943 , n252871 );
or ( n252944 , n252942 , n252943 );
nor ( n252945 , n252939 , n55146 );
nand ( n252946 , n252944 , n252945 );
nand ( n252947 , n245701 , n33833 );
nand ( n252948 , n252941 , n252946 , n252947 );
buf ( n252949 , n252948 );
not ( n252950 , n29952 );
not ( n252951 , n252950 );
not ( n252952 , n233907 );
nand ( n252953 , n29737 , n29569 );
not ( n252954 , n252953 );
or ( n252955 , n252952 , n252954 );
or ( n252956 , n252953 , n233907 );
nand ( n252957 , n252955 , n252956 );
not ( n252958 , n252957 );
nand ( n252959 , n29779 , n29950 );
not ( n252960 , n252959 );
not ( n252961 , n233133 );
and ( n252962 , n252960 , n252961 );
and ( n252963 , n252959 , n233133 );
nor ( n252964 , n252962 , n252963 );
not ( n252965 , n252964 );
or ( n252966 , n252958 , n252965 );
or ( n252967 , n252964 , n252957 );
nand ( n252968 , n252966 , n252967 );
not ( n252969 , n252968 );
nand ( n252970 , n29092 , n28948 );
not ( n252971 , n252970 );
not ( n252972 , n55448 );
and ( n252973 , n252971 , n252972 );
and ( n252974 , n252970 , n55448 );
nor ( n252975 , n252973 , n252974 );
not ( n252976 , n252975 );
not ( n252977 , n252976 );
not ( n252978 , n55412 );
nand ( n252979 , n29177 , n29341 );
not ( n252980 , n252979 );
or ( n252981 , n252978 , n252980 );
not ( n252982 , n55414 );
nand ( n252983 , n252982 , n29177 );
not ( n252984 , n55413 );
or ( n252985 , n252983 , n252984 );
nand ( n252986 , n252981 , n252985 );
not ( n252987 , n252986 );
not ( n252988 , n252987 );
or ( n252989 , n252977 , n252988 );
nand ( n252990 , n252986 , n252975 );
nand ( n252991 , n252989 , n252990 );
not ( n252992 , n55474 );
nor ( n252993 , n29473 , n29462 );
not ( n252994 , n252993 );
and ( n252995 , n252992 , n252994 );
nor ( n252996 , n29473 , n29462 );
and ( n252997 , n55474 , n252996 );
nor ( n252998 , n252995 , n252997 );
and ( n252999 , n252991 , n252998 );
not ( n253000 , n252991 );
not ( n253001 , n252998 );
and ( n253002 , n253000 , n253001 );
nor ( n253003 , n252999 , n253002 );
not ( n253004 , n253003 );
or ( n253005 , n252969 , n253004 );
not ( n253006 , n252968 );
not ( n253007 , n253003 );
nand ( n253008 , n253006 , n253007 );
nand ( n253009 , n253005 , n253008 );
not ( n253010 , n253009 );
or ( n253011 , n252951 , n253010 );
or ( n253012 , n253009 , n252950 );
nand ( n253013 , n253011 , n253012 );
not ( n253014 , n253013 );
buf ( n253015 , n248135 );
not ( n253016 , n253015 );
and ( n253017 , n253014 , n253016 );
and ( n253018 , n253013 , n253015 );
nor ( n253019 , n253017 , n253018 );
nand ( n253020 , n253019 , n247275 );
not ( n253021 , n227936 );
not ( n253022 , n248967 );
or ( n253023 , n253021 , n253022 );
not ( n253024 , n227936 );
nand ( n253025 , n253024 , n249394 );
nand ( n253026 , n253023 , n253025 );
and ( n253027 , n253026 , n248972 );
not ( n253028 , n253026 );
and ( n253029 , n253028 , n248975 );
nor ( n253030 , n253027 , n253029 );
not ( n253031 , n253030 );
not ( n253032 , n237130 );
not ( n253033 , n253032 );
not ( n253034 , n244657 );
nand ( n253035 , n237067 , n237058 );
not ( n253036 , n253035 );
not ( n253037 , n231120 );
and ( n253038 , n253036 , n253037 );
nand ( n253039 , n237067 , n237058 );
and ( n253040 , n253039 , n231120 );
nor ( n253041 , n253038 , n253040 );
not ( n253042 , n253041 );
or ( n253043 , n253034 , n253042 );
or ( n253044 , n253041 , n244657 );
nand ( n253045 , n253043 , n253044 );
nand ( n253046 , n250323 , n237028 );
and ( n253047 , n253046 , n231176 );
not ( n253048 , n253046 );
and ( n253049 , n253048 , n231198 );
nor ( n253050 , n253047 , n253049 );
xor ( n253051 , n253045 , n253050 );
nand ( n253052 , n237099 , n250345 );
and ( n253053 , n253052 , n53282 );
not ( n253054 , n253052 );
and ( n253055 , n253054 , n53283 );
nor ( n253056 , n253053 , n253055 );
not ( n253057 , n253056 );
nand ( n253058 , n237125 , n250337 );
not ( n253059 , n253058 );
not ( n253060 , n231061 );
and ( n253061 , n253059 , n253060 );
and ( n253062 , n253058 , n231061 );
nor ( n253063 , n253061 , n253062 );
not ( n253064 , n253063 );
or ( n253065 , n253057 , n253064 );
or ( n253066 , n253063 , n253056 );
nand ( n253067 , n253065 , n253066 );
not ( n253068 , n253067 );
and ( n253069 , n253051 , n253068 );
not ( n253070 , n253051 );
and ( n253071 , n253070 , n253067 );
nor ( n253072 , n253069 , n253071 );
not ( n253073 , n253072 );
not ( n253074 , n253073 );
not ( n253075 , n253074 );
or ( n253076 , n253033 , n253075 );
not ( n253077 , n253032 );
nand ( n253078 , n253077 , n253073 );
nand ( n253079 , n253076 , n253078 );
buf ( n253080 , n249194 );
buf ( n253081 , n253080 );
xor ( n253082 , n253079 , n253081 );
nand ( n253083 , n253031 , n253082 );
or ( n253084 , n253020 , n253083 );
not ( n253085 , n253082 );
not ( n253086 , n253019 );
or ( n253087 , n253085 , n253086 );
nor ( n253088 , n253031 , n251361 );
nand ( n253089 , n253087 , n253088 );
nand ( n253090 , n48251 , n38943 );
nand ( n253091 , n253084 , n253089 , n253090 );
buf ( n253092 , n253091 );
buf ( n253093 , n32336 );
not ( n253094 , n253093 );
not ( n253095 , n51269 );
or ( n253096 , n253094 , n253095 );
or ( n253097 , n51269 , n253093 );
nand ( n253098 , n253096 , n253097 );
not ( n253099 , n253098 );
not ( n253100 , n250746 );
and ( n253101 , n253099 , n253100 );
and ( n253102 , n253098 , n250746 );
nor ( n253103 , n253101 , n253102 );
nand ( n253104 , n253103 , n244515 );
not ( n253105 , n250714 );
buf ( n253106 , n54263 );
not ( n253107 , n253106 );
not ( n253108 , n218404 );
not ( n253109 , n253108 );
not ( n253110 , n251450 );
or ( n253111 , n253109 , n253110 );
nand ( n253112 , n251443 , n218404 );
nand ( n253113 , n253111 , n253112 );
not ( n253114 , n253113 );
or ( n253115 , n253107 , n253114 );
or ( n253116 , n253113 , n253106 );
nand ( n253117 , n253115 , n253116 );
not ( n253118 , n253117 );
nand ( n253119 , n253105 , n253118 );
or ( n253120 , n253104 , n253119 );
not ( n253121 , n253105 );
not ( n253122 , n253103 );
or ( n253123 , n253121 , n253122 );
nor ( n253124 , n253118 , n40465 );
nand ( n253125 , n253123 , n253124 );
nand ( n253126 , n31577 , n30902 );
nand ( n253127 , n253120 , n253125 , n253126 );
buf ( n253128 , n253127 );
buf ( n253129 , n247902 );
not ( n253130 , n253129 );
not ( n253131 , n239858 );
or ( n253132 , n253130 , n253131 );
or ( n253133 , n239858 , n253129 );
nand ( n253134 , n253132 , n253133 );
and ( n253135 , n253134 , n239924 );
not ( n253136 , n253134 );
and ( n253137 , n253136 , n239931 );
nor ( n253138 , n253135 , n253137 );
nand ( n253139 , n253138 , n205649 );
not ( n253140 , n224246 );
not ( n253141 , n51606 );
or ( n253142 , n253140 , n253141 );
not ( n253143 , n224246 );
nand ( n253144 , n253143 , n51597 );
nand ( n253145 , n253142 , n253144 );
not ( n253146 , n46001 );
nand ( n253147 , n253146 , n239806 );
and ( n253148 , n253147 , n46011 );
not ( n253149 , n253147 );
and ( n253150 , n253149 , n46010 );
nor ( n253151 , n253148 , n253150 );
nand ( n253152 , n223804 , n46693 );
not ( n253153 , n253152 );
buf ( n253154 , n46040 );
not ( n253155 , n253154 );
and ( n253156 , n253153 , n253155 );
and ( n253157 , n253152 , n253154 );
nor ( n253158 , n253156 , n253157 );
and ( n253159 , n253151 , n253158 );
not ( n253160 , n253151 );
not ( n253161 , n253158 );
and ( n253162 , n253160 , n253161 );
nor ( n253163 , n253159 , n253162 );
not ( n253164 , n253163 );
not ( n253165 , n244500 );
not ( n253166 , n45902 );
nand ( n253167 , n46529 , n253166 );
and ( n253168 , n253167 , n223650 );
not ( n253169 , n253167 );
and ( n253170 , n253169 , n45888 );
nor ( n253171 , n253168 , n253170 );
not ( n253172 , n253171 );
or ( n253173 , n253165 , n253172 );
or ( n253174 , n253171 , n244500 );
nand ( n253175 , n253173 , n253174 );
not ( n253176 , n45963 );
nand ( n253177 , n253176 , n239839 );
and ( n253178 , n253177 , n45974 );
not ( n253179 , n253177 );
and ( n253180 , n253179 , n45973 );
nor ( n253181 , n253178 , n253180 );
xor ( n253182 , n253175 , n253181 );
not ( n253183 , n253182 );
or ( n253184 , n253164 , n253183 );
not ( n253185 , n253182 );
not ( n253186 , n253163 );
nand ( n253187 , n253185 , n253186 );
nand ( n253188 , n253184 , n253187 );
buf ( n253189 , n253188 );
and ( n253190 , n253145 , n253189 );
not ( n253191 , n253145 );
not ( n253192 , n253185 );
not ( n253193 , n253186 );
and ( n253194 , n253192 , n253193 );
and ( n253195 , n253185 , n253186 );
nor ( n253196 , n253194 , n253195 );
buf ( n253197 , n253196 );
and ( n253198 , n253191 , n253197 );
nor ( n253199 , n253190 , n253198 );
not ( n253200 , n237630 );
not ( n253201 , n253200 );
not ( n253202 , n41216 );
or ( n253203 , n253201 , n253202 );
nand ( n253204 , n233987 , n237630 );
nand ( n253205 , n253203 , n253204 );
buf ( n253206 , n233997 );
and ( n253207 , n253205 , n253206 );
not ( n253208 , n253205 );
and ( n253209 , n253208 , n233990 );
nor ( n253210 , n253207 , n253209 );
nor ( n253211 , n253199 , n253210 );
or ( n253212 , n253139 , n253211 );
buf ( n253213 , n40465 );
nor ( n253214 , n253138 , n253213 );
nand ( n253215 , n253214 , n253211 );
nand ( n253216 , n48251 , n32124 );
nand ( n253217 , n253212 , n253215 , n253216 );
buf ( n253218 , n253217 );
not ( n253219 , RI19ab54d8_2414);
or ( n253220 , n25328 , n253219 );
not ( n253221 , RI19a83438_2771);
or ( n253222 , n25335 , n253221 );
nand ( n253223 , n253220 , n253222 );
buf ( n253224 , n253223 );
not ( n253225 , n252027 );
not ( n253226 , n253225 );
not ( n253227 , n49617 );
or ( n253228 , n253226 , n253227 );
not ( n253229 , n253225 );
nand ( n253230 , n253229 , n49626 );
nand ( n253231 , n253228 , n253230 );
nand ( n253232 , n240557 , n240388 );
not ( n253233 , n253232 );
not ( n253234 , n247354 );
and ( n253235 , n253233 , n253234 );
and ( n253236 , n253232 , n247354 );
nor ( n253237 , n253235 , n253236 );
nand ( n253238 , n240424 , n240614 );
not ( n253239 , n253238 );
not ( n253240 , n240602 );
and ( n253241 , n253239 , n253240 );
and ( n253242 , n253238 , n240602 );
nor ( n253243 , n253241 , n253242 );
xor ( n253244 , n253237 , n253243 );
xnor ( n253245 , n253244 , n252482 );
not ( n253246 , n253245 );
not ( n253247 , n240550 );
nand ( n253248 , n240489 , n240649 );
not ( n253249 , n253248 );
not ( n253250 , n246102 );
and ( n253251 , n253249 , n253250 );
and ( n253252 , n253248 , n246102 );
nor ( n253253 , n253251 , n253252 );
not ( n253254 , n253253 );
or ( n253255 , n253247 , n253254 );
not ( n253256 , n240550 );
not ( n253257 , n253253 );
nand ( n253258 , n253256 , n253257 );
nand ( n253259 , n253255 , n253258 );
and ( n253260 , n253246 , n253259 );
not ( n253261 , n253246 );
not ( n253262 , n253259 );
and ( n253263 , n253261 , n253262 );
nor ( n253264 , n253260 , n253263 );
buf ( n253265 , n253264 );
and ( n253266 , n253231 , n253265 );
not ( n253267 , n253231 );
and ( n253268 , n253245 , n253259 );
not ( n253269 , n253245 );
and ( n253270 , n253269 , n253262 );
nor ( n253271 , n253268 , n253270 );
buf ( n253272 , n253271 );
and ( n253273 , n253267 , n253272 );
nor ( n253274 , n253266 , n253273 );
nor ( n253275 , n253274 , n234110 );
not ( n253276 , n245159 );
not ( n253277 , n40914 );
or ( n253278 , n253276 , n253277 );
or ( n253279 , n40918 , n245159 );
nand ( n253280 , n253278 , n253279 );
not ( n253281 , n253280 );
not ( n253282 , n41217 );
and ( n253283 , n253281 , n253282 );
and ( n253284 , n253280 , n218982 );
nor ( n253285 , n253283 , n253284 );
not ( n253286 , n253285 );
buf ( n253287 , n250098 );
not ( n253288 , n253287 );
not ( n253289 , n253288 );
and ( n253290 , n248672 , n248605 );
not ( n253291 , n248672 );
and ( n253292 , n253291 , n248606 );
nor ( n253293 , n253290 , n253292 );
not ( n253294 , n253293 );
buf ( n253295 , n243119 );
not ( n253296 , n253295 );
and ( n253297 , n253294 , n253296 );
and ( n253298 , n248677 , n253295 );
nor ( n253299 , n253297 , n253298 );
not ( n253300 , n253299 );
or ( n253301 , n253289 , n253300 );
not ( n253302 , n253299 );
nand ( n253303 , n253302 , n253287 );
nand ( n253304 , n253301 , n253303 );
nor ( n253305 , n253286 , n253304 );
nand ( n253306 , n253275 , n253305 );
not ( n253307 , n253304 );
not ( n253308 , n253307 );
not ( n253309 , n253274 );
not ( n253310 , n253309 );
or ( n253311 , n253308 , n253310 );
nor ( n253312 , n253285 , n43968 );
nand ( n253313 , n253311 , n253312 );
nand ( n253314 , n55760 , n47408 );
nand ( n253315 , n253306 , n253313 , n253314 );
buf ( n253316 , n253315 );
not ( n253317 , n25840 );
not ( n253318 , n39766 );
or ( n253319 , n253317 , n253318 );
not ( n253320 , n249914 );
not ( n253321 , n227707 );
or ( n253322 , n253320 , n253321 );
or ( n253323 , n227707 , n249914 );
nand ( n253324 , n253322 , n253323 );
and ( n253325 , n253324 , n242978 );
not ( n253326 , n253324 );
and ( n253327 , n253326 , n242970 );
nor ( n253328 , n253325 , n253327 );
not ( n253329 , n253328 );
not ( n253330 , n228270 );
not ( n253331 , n35804 );
or ( n253332 , n253330 , n253331 );
nand ( n253333 , n35811 , n50506 );
nand ( n253334 , n253332 , n253333 );
not ( n253335 , n253334 );
buf ( n253336 , n235008 );
not ( n253337 , n253336 );
and ( n253338 , n253335 , n253337 );
and ( n253339 , n253334 , n253336 );
nor ( n253340 , n253338 , n253339 );
nand ( n253341 , n253329 , n253340 );
not ( n253342 , n252634 );
not ( n253343 , n253264 );
or ( n253344 , n253342 , n253343 );
not ( n253345 , n252634 );
nand ( n253346 , n253345 , n253271 );
nand ( n253347 , n253344 , n253346 );
not ( n253348 , n232900 );
and ( n253349 , n253347 , n253348 );
not ( n253350 , n253347 );
and ( n253351 , n253350 , n55135 );
nor ( n253352 , n253349 , n253351 );
and ( n253353 , n253341 , n253352 );
not ( n253354 , n253341 );
not ( n253355 , n253352 );
and ( n253356 , n253354 , n253355 );
nor ( n253357 , n253353 , n253356 );
not ( n253358 , n205649 );
or ( n253359 , n253357 , n253358 );
nand ( n253360 , n253319 , n253359 );
buf ( n253361 , n253360 );
not ( n253362 , n245392 );
not ( n253363 , n253362 );
not ( n253364 , n253363 );
not ( n253365 , n241316 );
not ( n253366 , n245333 );
or ( n253367 , n253365 , n253366 );
not ( n253368 , n241316 );
nand ( n253369 , n253368 , n245338 );
nand ( n253370 , n253367 , n253369 );
not ( n253371 , n253370 );
or ( n253372 , n253364 , n253371 );
or ( n253373 , n253370 , n253363 );
nand ( n253374 , n253372 , n253373 );
not ( n253375 , n253374 );
xor ( n253376 , n242467 , n227548 );
buf ( n253377 , n241656 );
not ( n253378 , n253377 );
xnor ( n253379 , n253376 , n253378 );
not ( n253380 , n253379 );
or ( n253381 , n253375 , n253380 );
not ( n253382 , n250485 );
not ( n253383 , n234691 );
or ( n253384 , n253382 , n253383 );
not ( n253385 , n234691 );
not ( n253386 , n253385 );
or ( n253387 , n253386 , n250485 );
nand ( n253388 , n253384 , n253387 );
and ( n253389 , n253388 , n234804 );
not ( n253390 , n253388 );
and ( n253391 , n253390 , n234811 );
nor ( n253392 , n253389 , n253391 );
not ( n253393 , n219702 );
nand ( n253394 , n253392 , n253393 );
not ( n253395 , n253394 );
nand ( n253396 , n253381 , n253395 );
not ( n253397 , n55152 );
nand ( n253398 , n253379 , n253397 );
not ( n253399 , n253398 );
not ( n253400 , n253374 );
nor ( n253401 , n253392 , n253400 );
nand ( n253402 , n253399 , n253401 );
nand ( n253403 , n245702 , n37914 );
nand ( n253404 , n253396 , n253402 , n253403 );
buf ( n253405 , n253404 );
nor ( n253406 , n253352 , n253340 );
not ( n253407 , n247054 );
not ( n253408 , n226975 );
nand ( n253409 , n49232 , n247034 );
not ( n253410 , n253409 );
or ( n253411 , n253408 , n253410 );
or ( n253412 , n253409 , n226975 );
nand ( n253413 , n253411 , n253412 );
not ( n253414 , n253413 );
nand ( n253415 , n247046 , n49261 );
not ( n253416 , n253415 );
not ( n253417 , n250560 );
and ( n253418 , n253416 , n253417 );
and ( n253419 , n253415 , n250560 );
nor ( n253420 , n253418 , n253419 );
not ( n253421 , n253420 );
or ( n253422 , n253414 , n253421 );
or ( n253423 , n253420 , n253413 );
nand ( n253424 , n253422 , n253423 );
not ( n253425 , n253424 );
not ( n253426 , n253425 );
not ( n253427 , n247070 );
nand ( n253428 , n253427 , n227160 );
not ( n253429 , n253428 );
not ( n253430 , n250521 );
and ( n253431 , n253429 , n253430 );
not ( n253432 , n250521 );
not ( n253433 , n253432 );
and ( n253434 , n253428 , n253433 );
nor ( n253435 , n253431 , n253434 );
not ( n253436 , n253435 );
nand ( n253437 , n49348 , n247087 );
not ( n253438 , n250537 );
and ( n253439 , n253437 , n253438 );
not ( n253440 , n253437 );
and ( n253441 , n253440 , n250537 );
nor ( n253442 , n253439 , n253441 );
not ( n253443 , n253442 );
or ( n253444 , n253436 , n253443 );
or ( n253445 , n253435 , n253442 );
nand ( n253446 , n253444 , n253445 );
not ( n253447 , n249076 );
not ( n253448 , n253447 );
nor ( n253449 , n247108 , n49302 );
not ( n253450 , n253449 );
and ( n253451 , n253448 , n253450 );
and ( n253452 , n253447 , n253449 );
nor ( n253453 , n253451 , n253452 );
not ( n253454 , n253453 );
and ( n253455 , n253446 , n253454 );
not ( n253456 , n253446 );
and ( n253457 , n253456 , n253453 );
nor ( n253458 , n253455 , n253457 );
not ( n253459 , n253458 );
or ( n253460 , n253426 , n253459 );
not ( n253461 , n253458 );
nand ( n253462 , n253461 , n253424 );
nand ( n253463 , n253460 , n253462 );
not ( n253464 , n253463 );
not ( n253465 , n253464 );
or ( n253466 , n253407 , n253465 );
or ( n253467 , n253464 , n247054 );
nand ( n253468 , n253466 , n253467 );
not ( n253469 , n248253 );
not ( n253470 , n253469 );
not ( n253471 , n248270 );
and ( n253472 , n253470 , n253471 );
and ( n253473 , n253469 , n248270 );
nor ( n253474 , n253472 , n253473 );
buf ( n253475 , n253474 );
and ( n253476 , n253468 , n253475 );
not ( n253477 , n253468 );
buf ( n253478 , n248276 );
and ( n253479 , n253477 , n253478 );
nor ( n253480 , n253476 , n253479 );
not ( n253481 , n253480 );
nand ( n253482 , n253481 , n237385 );
or ( n253483 , n253406 , n253482 );
nor ( n253484 , n253481 , n219702 );
nand ( n253485 , n253484 , n253406 );
buf ( n253486 , n35431 );
nand ( n253487 , n253486 , n37549 );
nand ( n253488 , n253483 , n253485 , n253487 );
buf ( n253489 , n253488 );
not ( n253490 , n204764 );
not ( n253491 , n245702 );
or ( n253492 , n253490 , n253491 );
not ( n253493 , n234586 );
not ( n253494 , n249284 );
or ( n253495 , n253493 , n253494 );
not ( n253496 , n234586 );
nand ( n253497 , n253496 , n249522 );
nand ( n253498 , n253495 , n253497 );
and ( n253499 , n253498 , n249525 );
not ( n253500 , n253498 );
and ( n253501 , n253500 , n249528 );
nor ( n253502 , n253499 , n253501 );
not ( n253503 , n47711 );
not ( n253504 , n253503 );
not ( n253505 , n238033 );
or ( n253506 , n253504 , n253505 );
not ( n253507 , n253503 );
nand ( n253508 , n253507 , n238040 );
nand ( n253509 , n253506 , n253508 );
and ( n253510 , n253509 , n238102 );
not ( n253511 , n253509 );
and ( n253512 , n253511 , n238107 );
nor ( n253513 , n253510 , n253512 );
nand ( n253514 , n253502 , n253513 );
not ( n253515 , n53223 );
nand ( n253516 , n246571 , n33144 );
not ( n253517 , n253516 );
or ( n253518 , n253515 , n253517 );
or ( n253519 , n253516 , n53223 );
nand ( n253520 , n253518 , n253519 );
not ( n253521 , n253520 );
not ( n253522 , n33246 );
or ( n253523 , n253521 , n253522 );
not ( n253524 , n253520 );
not ( n253525 , n33240 );
not ( n253526 , n32927 );
or ( n253527 , n253525 , n253526 );
not ( n253528 , n32927 );
nand ( n253529 , n253528 , n33241 );
nand ( n253530 , n253527 , n253529 );
nand ( n253531 , n253524 , n253530 );
nand ( n253532 , n253523 , n253531 );
buf ( n253533 , n244704 );
and ( n253534 , n253532 , n253533 );
not ( n253535 , n253532 );
buf ( n253536 , n244711 );
and ( n253537 , n253535 , n253536 );
nor ( n253538 , n253534 , n253537 );
not ( n253539 , n253538 );
and ( n253540 , n253514 , n253539 );
not ( n253541 , n253514 );
and ( n253542 , n253541 , n253538 );
nor ( n253543 , n253540 , n253542 );
not ( n253544 , n205649 );
or ( n253545 , n253543 , n253544 );
nand ( n253546 , n253492 , n253545 );
buf ( n253547 , n253546 );
not ( n253548 , n45068 );
not ( n253549 , n244054 );
or ( n253550 , n253548 , n253549 );
not ( n253551 , n45068 );
not ( n253552 , n244050 );
not ( n253553 , n244043 );
not ( n253554 , n253553 );
or ( n253555 , n253552 , n253554 );
nand ( n253556 , n244043 , n244049 );
nand ( n253557 , n253555 , n253556 );
nand ( n253558 , n253551 , n253557 );
nand ( n253559 , n253550 , n253558 );
not ( n253560 , n245517 );
and ( n253561 , n253559 , n253560 );
not ( n253562 , n253559 );
and ( n253563 , n253562 , n245517 );
nor ( n253564 , n253561 , n253563 );
not ( n253565 , n247698 );
nand ( n253566 , n253564 , n253565 );
not ( n253567 , n244978 );
not ( n253568 , n229231 );
not ( n253569 , n253568 );
not ( n253570 , n239653 );
or ( n253571 , n253569 , n253570 );
nand ( n253572 , n244125 , n229231 );
nand ( n253573 , n253571 , n253572 );
not ( n253574 , n253573 );
or ( n253575 , n253567 , n253574 );
or ( n253576 , n253573 , n244978 );
nand ( n253577 , n253575 , n253576 );
not ( n253578 , n253463 );
buf ( n253579 , n253578 );
not ( n253580 , n253579 );
not ( n253581 , n247635 );
not ( n253582 , n48233 );
or ( n253583 , n253581 , n253582 );
not ( n253584 , n247635 );
nand ( n253585 , n253584 , n48232 );
nand ( n253586 , n253583 , n253585 );
not ( n253587 , n253586 );
or ( n253588 , n253580 , n253587 );
or ( n253589 , n253579 , n253586 );
nand ( n253590 , n253588 , n253589 );
not ( n253591 , n253590 );
nand ( n253592 , n253577 , n253591 );
or ( n253593 , n253566 , n253592 );
not ( n253594 , n253577 );
not ( n253595 , n253564 );
or ( n253596 , n253594 , n253595 );
nor ( n253597 , n253591 , n52445 );
nand ( n253598 , n253596 , n253597 );
nand ( n253599 , n50615 , n41284 );
nand ( n253600 , n253593 , n253598 , n253599 );
buf ( n253601 , n253600 );
not ( n253602 , n248196 );
not ( n253603 , n240001 );
or ( n253604 , n253602 , n253603 );
not ( n253605 , n248196 );
nand ( n253606 , n253605 , n239994 );
nand ( n253607 , n253604 , n253606 );
and ( n253608 , n253607 , n240053 );
not ( n253609 , n253607 );
and ( n253610 , n253609 , n240057 );
nor ( n253611 , n253608 , n253610 );
nor ( n253612 , n253611 , n221279 );
not ( n253613 , n253612 );
not ( n253614 , n53197 );
nand ( n253615 , n230940 , n32786 );
not ( n253616 , n253615 );
buf ( n253617 , n246630 );
not ( n253618 , n253617 );
and ( n253619 , n253616 , n253618 );
nand ( n253620 , n230940 , n32786 );
and ( n253621 , n253620 , n253617 );
nor ( n253622 , n253619 , n253621 );
not ( n253623 , n230920 );
nand ( n253624 , n32496 , n253623 );
and ( n253625 , n253624 , n246614 );
not ( n253626 , n253624 );
not ( n253627 , n246614 );
and ( n253628 , n253626 , n253627 );
nor ( n253629 , n253625 , n253628 );
or ( n253630 , n253622 , n253629 );
nand ( n253631 , n253629 , n253622 );
nand ( n253632 , n253630 , n253631 );
nand ( n253633 , n53193 , n32917 );
not ( n253634 , n253633 );
buf ( n253635 , n246594 );
not ( n253636 , n253635 );
and ( n253637 , n253634 , n253636 );
and ( n253638 , n253633 , n253635 );
nor ( n253639 , n253637 , n253638 );
and ( n253640 , n253632 , n253639 );
not ( n253641 , n253632 );
not ( n253642 , n253639 );
and ( n253643 , n253641 , n253642 );
nor ( n253644 , n253640 , n253643 );
not ( n253645 , n253644 );
not ( n253646 , n53216 );
nand ( n253647 , n253646 , n33049 );
not ( n253648 , n253647 );
not ( n253649 , n246565 );
and ( n253650 , n253648 , n253649 );
not ( n253651 , n53217 );
nand ( n253652 , n253651 , n33049 );
and ( n253653 , n253652 , n246565 );
nor ( n253654 , n253650 , n253653 );
not ( n253655 , n253654 );
nand ( n253656 , n33232 , n230995 );
and ( n253657 , n253656 , n246572 );
not ( n253658 , n253656 );
and ( n253659 , n253658 , n246571 );
nor ( n253660 , n253657 , n253659 );
not ( n253661 , n253660 );
or ( n253662 , n253655 , n253661 );
or ( n253663 , n253654 , n253660 );
nand ( n253664 , n253662 , n253663 );
not ( n253665 , n253664 );
and ( n253666 , n253645 , n253665 );
and ( n253667 , n253644 , n253664 );
nor ( n253668 , n253666 , n253667 );
buf ( n253669 , n253668 );
not ( n253670 , n253669 );
or ( n253671 , n253614 , n253670 );
not ( n253672 , n53197 );
not ( n253673 , n253668 );
nand ( n253674 , n253672 , n253673 );
nand ( n253675 , n253671 , n253674 );
buf ( n253676 , n250359 );
and ( n253677 , n253675 , n253676 );
not ( n253678 , n253675 );
buf ( n253679 , n250366 );
and ( n253680 , n253678 , n253679 );
nor ( n253681 , n253677 , n253680 );
buf ( n253682 , n51559 );
not ( n253683 , n253682 );
not ( n253684 , n45877 );
or ( n253685 , n253683 , n253684 );
or ( n253686 , n241695 , n253682 );
nand ( n253687 , n253685 , n253686 );
not ( n253688 , n253687 );
not ( n253689 , n46067 );
and ( n253690 , n253688 , n253689 );
and ( n253691 , n253687 , n241701 );
nor ( n253692 , n253690 , n253691 );
nand ( n253693 , n253681 , n253692 );
or ( n253694 , n253613 , n253693 );
not ( n253695 , n253611 );
not ( n253696 , n253695 );
not ( n253697 , n253681 );
or ( n253698 , n253696 , n253697 );
nor ( n253699 , n253692 , n55104 );
nand ( n253700 , n253698 , n253699 );
nand ( n253701 , n245414 , n29922 );
nand ( n253702 , n253694 , n253700 , n253701 );
buf ( n253703 , n253702 );
not ( n253704 , n33009 );
not ( n253705 , n253704 );
nand ( n253706 , n32990 , n246565 );
not ( n253707 , n253706 );
and ( n253708 , n253705 , n253707 );
and ( n253709 , n253704 , n253706 );
nor ( n253710 , n253708 , n253709 );
not ( n253711 , n253710 );
not ( n253712 , n253530 );
or ( n253713 , n253711 , n253712 );
or ( n253714 , n253530 , n253710 );
nand ( n253715 , n253713 , n253714 );
and ( n253716 , n253715 , n253533 );
not ( n253717 , n253715 );
and ( n253718 , n253717 , n253536 );
nor ( n253719 , n253716 , n253718 );
nor ( n253720 , n253719 , n243434 );
not ( n253721 , n253720 );
not ( n253722 , n228085 );
not ( n253723 , n253722 );
not ( n253724 , n53811 );
or ( n253725 , n253723 , n253724 );
not ( n253726 , n253722 );
nand ( n253727 , n253726 , n53820 );
nand ( n253728 , n253725 , n253727 );
not ( n253729 , n231768 );
not ( n253730 , n253729 );
and ( n253731 , n253728 , n253730 );
not ( n253732 , n253728 );
and ( n253733 , n253732 , n231776 );
nor ( n253734 , n253731 , n253733 );
not ( n253735 , n253734 );
not ( n253736 , n245615 );
buf ( n253737 , n246143 );
not ( n253738 , n253737 );
not ( n253739 , n245602 );
or ( n253740 , n253738 , n253739 );
not ( n253741 , n253737 );
nand ( n253742 , n253741 , n245611 );
nand ( n253743 , n253740 , n253742 );
not ( n253744 , n253743 );
or ( n253745 , n253736 , n253744 );
buf ( n253746 , n240941 );
or ( n253747 , n253743 , n253746 );
nand ( n253748 , n253745 , n253747 );
not ( n253749 , n253748 );
nand ( n253750 , n253735 , n253749 );
or ( n253751 , n253721 , n253750 );
not ( n253752 , n253749 );
not ( n253753 , n253719 );
not ( n253754 , n253753 );
or ( n253755 , n253752 , n253754 );
nor ( n253756 , n253735 , n221279 );
nand ( n253757 , n253755 , n253756 );
nand ( n253758 , n234453 , n36913 );
nand ( n253759 , n253751 , n253757 , n253758 );
buf ( n253760 , n253759 );
buf ( n253761 , n253453 );
not ( n253762 , n253761 );
nand ( n253763 , n247047 , n250559 );
and ( n253764 , n253763 , n49248 );
not ( n253765 , n253763 );
and ( n253766 , n253765 , n227008 );
nor ( n253767 , n253764 , n253766 );
not ( n253768 , n253767 );
not ( n253769 , n251989 );
and ( n253770 , n253768 , n253769 );
and ( n253771 , n253767 , n251989 );
nor ( n253772 , n253770 , n253771 );
not ( n253773 , n253772 );
not ( n253774 , n227146 );
nand ( n253775 , n253432 , n247070 );
not ( n253776 , n253775 );
or ( n253777 , n253774 , n253776 );
nand ( n253778 , n253432 , n247073 );
or ( n253779 , n253778 , n227146 );
nand ( n253780 , n253777 , n253779 );
not ( n253781 , n253780 );
nand ( n253782 , n253438 , n247086 );
not ( n253783 , n253782 );
not ( n253784 , n49332 );
and ( n253785 , n253783 , n253784 );
and ( n253786 , n253782 , n49332 );
nor ( n253787 , n253785 , n253786 );
not ( n253788 , n253787 );
or ( n253789 , n253781 , n253788 );
or ( n253790 , n253787 , n253780 );
nand ( n253791 , n253789 , n253790 );
not ( n253792 , n253791 );
nand ( n253793 , n253447 , n247108 );
not ( n253794 , n253793 );
not ( n253795 , n49291 );
and ( n253796 , n253794 , n253795 );
and ( n253797 , n253793 , n49291 );
nor ( n253798 , n253796 , n253797 );
not ( n253799 , n253798 );
or ( n253800 , n253792 , n253799 );
or ( n253801 , n253798 , n253791 );
nand ( n253802 , n253800 , n253801 );
not ( n253803 , n253802 );
or ( n253804 , n253773 , n253803 );
or ( n253805 , n253802 , n253772 );
nand ( n253806 , n253804 , n253805 );
buf ( n253807 , n253806 );
not ( n253808 , n253807 );
or ( n253809 , n253762 , n253808 );
or ( n253810 , n253807 , n253761 );
nand ( n253811 , n253809 , n253810 );
not ( n253812 , n253811 );
not ( n253813 , n240316 );
not ( n253814 , n253813 );
and ( n253815 , n253812 , n253814 );
and ( n253816 , n253811 , n253813 );
nor ( n253817 , n253815 , n253816 );
nand ( n253818 , n253817 , n235051 );
not ( n253819 , n239858 );
not ( n253820 , n36485 );
not ( n253821 , n251324 );
nand ( n253822 , n36458 , n36417 );
not ( n253823 , n253822 );
not ( n253824 , n46461 );
and ( n253825 , n253823 , n253824 );
and ( n253826 , n253822 , n46461 );
nor ( n253827 , n253825 , n253826 );
not ( n253828 , n253827 );
or ( n253829 , n253821 , n253828 );
or ( n253830 , n253827 , n251324 );
nand ( n253831 , n253829 , n253830 );
not ( n253832 , n253831 );
not ( n253833 , n224197 );
and ( n253834 , n253832 , n253833 );
and ( n253835 , n253831 , n224197 );
nor ( n253836 , n253834 , n253835 );
not ( n253837 , n253836 );
nand ( n253838 , n36580 , n36628 );
not ( n253839 , n253838 );
not ( n253840 , n224248 );
and ( n253841 , n253839 , n253840 );
and ( n253842 , n253838 , n224248 );
nor ( n253843 , n253841 , n253842 );
not ( n253844 , n253843 );
nand ( n253845 , n36715 , n45836 );
and ( n253846 , n253845 , n46478 );
not ( n253847 , n253845 );
and ( n253848 , n253847 , n45754 );
nor ( n253849 , n253846 , n253848 );
not ( n253850 , n253849 );
or ( n253851 , n253844 , n253850 );
or ( n253852 , n253849 , n253843 );
nand ( n253853 , n253851 , n253852 );
not ( n253854 , n253853 );
xor ( n253855 , n253837 , n253854 );
not ( n253856 , n253855 );
or ( n253857 , n253820 , n253856 );
not ( n253858 , n36485 );
not ( n253859 , n253853 );
not ( n253860 , n253836 );
or ( n253861 , n253859 , n253860 );
nand ( n253862 , n253837 , n253854 );
nand ( n253863 , n253861 , n253862 );
nand ( n253864 , n253858 , n253863 );
nand ( n253865 , n253857 , n253864 );
not ( n253866 , n253865 );
or ( n253867 , n253819 , n253866 );
or ( n253868 , n253865 , n239855 );
nand ( n253869 , n253867 , n253868 );
not ( n253870 , n249882 );
not ( n253871 , n227707 );
or ( n253872 , n253870 , n253871 );
or ( n253873 , n227707 , n249882 );
nand ( n253874 , n253872 , n253873 );
and ( n253875 , n253874 , n242978 );
not ( n253876 , n253874 );
and ( n253877 , n253876 , n242970 );
nor ( n253878 , n253875 , n253877 );
nand ( n253879 , n253869 , n253878 );
or ( n253880 , n253818 , n253879 );
not ( n253881 , n253869 );
not ( n253882 , n253817 );
or ( n253883 , n253881 , n253882 );
nor ( n253884 , n253878 , n239237 );
nand ( n253885 , n253883 , n253884 );
nand ( n253886 , n238114 , n32487 );
nand ( n253887 , n253880 , n253885 , n253886 );
buf ( n253888 , n253887 );
not ( n253889 , n250826 );
nand ( n253890 , n250815 , n253889 );
not ( n253891 , n242191 );
not ( n253892 , n27876 );
or ( n253893 , n253891 , n253892 );
not ( n253894 , n242191 );
nand ( n253895 , n253894 , n27869 );
nand ( n253896 , n253893 , n253895 );
and ( n253897 , n253896 , n248756 );
not ( n253898 , n253896 );
and ( n253899 , n253898 , n248763 );
nor ( n253900 , n253897 , n253899 );
not ( n253901 , n253900 );
not ( n253902 , n226004 );
nand ( n253903 , n253890 , n253901 , n253902 );
buf ( n253904 , n233971 );
nor ( n253905 , n250826 , n253904 );
nand ( n253906 , n253900 , n253905 , n250815 );
nand ( n253907 , n37728 , n204329 );
nand ( n253908 , n253903 , n253906 , n253907 );
buf ( n253909 , n253908 );
buf ( n253910 , n31669 );
or ( n253911 , n233507 , n49062 );
not ( n253912 , RI19ac6bc0_2279);
or ( n253913 , n25335 , n253912 );
nand ( n253914 , n253911 , n253913 );
buf ( n253915 , n253914 );
buf ( n253916 , n210076 );
not ( n253917 , n52757 );
not ( n253918 , n245733 );
not ( n253919 , n230367 );
or ( n253920 , n253918 , n253919 );
not ( n253921 , n245733 );
nand ( n253922 , n253921 , n230374 );
nand ( n253923 , n253920 , n253922 );
not ( n253924 , n253923 );
or ( n253925 , n253917 , n253924 );
or ( n253926 , n253923 , n52757 );
nand ( n253927 , n253925 , n253926 );
not ( n253928 , n246680 );
nand ( n253929 , n253927 , n253928 );
not ( n253930 , n253929 );
not ( n253931 , n34398 );
not ( n253932 , n244190 );
or ( n253933 , n253931 , n253932 );
not ( n253934 , n34398 );
nand ( n253935 , n253934 , n244199 );
nand ( n253936 , n253933 , n253935 );
and ( n253937 , n253936 , n244208 );
not ( n253938 , n253936 );
and ( n253939 , n253938 , n244204 );
nor ( n253940 , n253937 , n253939 );
not ( n253941 , n253940 );
not ( n253942 , n46551 );
not ( n253943 , n253196 );
or ( n253944 , n253942 , n253943 );
not ( n253945 , n46551 );
nand ( n253946 , n253945 , n253188 );
nand ( n253947 , n253944 , n253946 );
buf ( n253948 , n248055 );
not ( n253949 , n253948 );
and ( n253950 , n253947 , n253949 );
not ( n253951 , n253947 );
and ( n253952 , n253951 , n253948 );
nor ( n253953 , n253950 , n253952 );
nand ( n253954 , n253941 , n253953 );
not ( n253955 , n253954 );
and ( n253956 , n253930 , n253955 );
and ( n253957 , n39766 , n34231 );
nor ( n253958 , n253956 , n253957 );
nor ( n253959 , n253927 , n252358 );
not ( n253960 , n253953 );
nand ( n253961 , n253959 , n253960 );
nor ( n253962 , n253953 , n219702 );
nand ( n253963 , n253962 , n253940 );
nand ( n253964 , n253958 , n253961 , n253963 );
buf ( n253965 , n253964 );
not ( n253966 , n242139 );
not ( n253967 , n204544 );
or ( n253968 , n253966 , n253967 );
not ( n253969 , n242139 );
nand ( n253970 , n253969 , n204553 );
nand ( n253971 , n253968 , n253970 );
not ( n253972 , n253971 );
not ( n253973 , n27878 );
and ( n253974 , n253972 , n253973 );
and ( n253975 , n253971 , n27878 );
nor ( n253976 , n253974 , n253975 );
not ( n253977 , n253976 );
nor ( n253978 , n253977 , n221279 );
nand ( n253979 , n253978 , n249287 );
not ( n253980 , n249287 );
nor ( n253981 , n253980 , n33254 );
not ( n253982 , n244671 );
not ( n253983 , n241715 );
or ( n253984 , n253982 , n253983 );
not ( n253985 , n244671 );
nand ( n253986 , n253985 , n241723 );
nand ( n253987 , n253984 , n253986 );
and ( n253988 , n253987 , n241878 );
not ( n253989 , n253987 );
and ( n253990 , n253989 , n241885 );
nor ( n253991 , n253988 , n253990 );
nand ( n253992 , n253981 , n253991 );
nor ( n253993 , n249287 , n253991 );
nor ( n253994 , n253976 , n46425 );
nand ( n253995 , n253993 , n253994 );
nand ( n253996 , n46083 , n38097 );
nand ( n253997 , n253979 , n253992 , n253995 , n253996 );
buf ( n253998 , n253997 );
buf ( n253999 , n35543 );
buf ( n254000 , n204880 );
not ( n254001 , n237891 );
not ( n254002 , n246759 );
or ( n254003 , n254001 , n254002 );
or ( n254004 , n246759 , n237891 );
nand ( n254005 , n254003 , n254004 );
buf ( n254006 , n247822 );
and ( n254007 , n254005 , n254006 );
not ( n254008 , n254005 );
not ( n254009 , n247813 );
not ( n254010 , n254009 );
and ( n254011 , n254008 , n254010 );
nor ( n254012 , n254007 , n254011 );
not ( n254013 , n252070 );
nand ( n254014 , n254012 , n254013 );
not ( n254015 , n43210 );
not ( n254016 , n244453 );
or ( n254017 , n254015 , n254016 );
or ( n254018 , n244453 , n43210 );
nand ( n254019 , n254017 , n254018 );
and ( n254020 , n254019 , n249789 );
not ( n254021 , n254019 );
and ( n254022 , n254021 , n249792 );
nor ( n254023 , n254020 , n254022 );
not ( n254024 , n254023 );
not ( n254025 , n236239 );
not ( n254026 , n254025 );
not ( n254027 , n241256 );
or ( n254028 , n254026 , n254027 );
not ( n254029 , n254025 );
nand ( n254030 , n254029 , n241255 );
nand ( n254031 , n254028 , n254030 );
and ( n254032 , n254031 , n241360 );
not ( n254033 , n254031 );
and ( n254034 , n254033 , n241370 );
nor ( n254035 , n254032 , n254034 );
nand ( n254036 , n254024 , n254035 );
or ( n254037 , n254014 , n254036 );
not ( n254038 , n254024 );
not ( n254039 , n254012 );
or ( n254040 , n254038 , n254039 );
nor ( n254041 , n254035 , n243204 );
nand ( n254042 , n254040 , n254041 );
nand ( n254043 , n251465 , n35684 );
nand ( n254044 , n254037 , n254042 , n254043 );
buf ( n254045 , n254044 );
not ( n254046 , RI19aa3c88_2539);
or ( n254047 , n25328 , n254046 );
not ( n254048 , RI19a9a610_2609);
or ( n254049 , n25335 , n254048 );
nand ( n254050 , n254047 , n254049 );
buf ( n254051 , n254050 );
buf ( n254052 , n204809 );
buf ( n254053 , n205168 );
not ( n254054 , n242785 );
not ( n254055 , n242977 );
or ( n254056 , n254054 , n254055 );
not ( n254057 , n242785 );
nand ( n254058 , n254057 , n242969 );
nand ( n254059 , n254056 , n254058 );
buf ( n254060 , n246963 );
and ( n254061 , n254059 , n254060 );
not ( n254062 , n254059 );
buf ( n254063 , n246968 );
and ( n254064 , n254062 , n254063 );
nor ( n254065 , n254061 , n254064 );
nor ( n254066 , n254065 , n40465 );
not ( n254067 , n47281 );
not ( n254068 , n245170 );
or ( n254069 , n254067 , n254068 );
not ( n254070 , n47281 );
not ( n254071 , n245139 );
not ( n254072 , n254071 );
not ( n254073 , n245164 );
or ( n254074 , n254072 , n254073 );
nand ( n254075 , n245165 , n245139 );
nand ( n254076 , n254074 , n254075 );
not ( n254077 , n254076 );
nand ( n254078 , n254070 , n254077 );
nand ( n254079 , n254069 , n254078 );
buf ( n254080 , n237647 );
and ( n254081 , n254079 , n254080 );
not ( n254082 , n254079 );
buf ( n254083 , n237639 );
and ( n254084 , n254082 , n254083 );
nor ( n254085 , n254081 , n254084 );
not ( n254086 , n249174 );
not ( n254087 , n244776 );
or ( n254088 , n254086 , n254087 );
not ( n254089 , n249174 );
nand ( n254090 , n254089 , n244768 );
nand ( n254091 , n254088 , n254090 );
and ( n254092 , n254091 , n252934 );
not ( n254093 , n254091 );
and ( n254094 , n254093 , n249059 );
nor ( n254095 , n254092 , n254094 );
nor ( n254096 , n254085 , n254095 );
nand ( n254097 , n254066 , n254096 );
not ( n254098 , n254095 );
not ( n254099 , n254098 );
not ( n254100 , n254065 );
not ( n254101 , n254100 );
or ( n254102 , n254099 , n254101 );
not ( n254103 , n254085 );
nor ( n254104 , n254103 , n235050 );
nand ( n254105 , n254102 , n254104 );
nand ( n254106 , n55760 , n38854 );
nand ( n254107 , n254097 , n254105 , n254106 );
buf ( n254108 , n254107 );
buf ( n254109 , n32514 );
nor ( n254110 , n252352 , n31571 );
buf ( n254111 , n234930 );
not ( n254112 , n254111 );
not ( n254113 , n236988 );
not ( n254114 , n236954 );
or ( n254115 , n254113 , n254114 );
nand ( n254116 , n236987 , n236955 );
nand ( n254117 , n254115 , n254116 );
not ( n254118 , n254117 );
or ( n254119 , n254112 , n254118 );
or ( n254120 , n254117 , n254111 );
nand ( n254121 , n254119 , n254120 );
buf ( n254122 , n233035 );
and ( n254123 , n254121 , n254122 );
not ( n254124 , n254121 );
buf ( n254125 , n233026 );
and ( n254126 , n254124 , n254125 );
nor ( n254127 , n254123 , n254126 );
nor ( n254128 , n252339 , n254127 );
nand ( n254129 , n254110 , n254128 );
not ( n254130 , n252352 );
not ( n254131 , n254130 );
not ( n254132 , n252340 );
or ( n254133 , n254131 , n254132 );
not ( n254134 , n254127 );
nor ( n254135 , n254134 , n252070 );
nand ( n254136 , n254133 , n254135 );
nand ( n254137 , n246217 , n38526 );
nand ( n254138 , n254129 , n254136 , n254137 );
buf ( n254139 , n254138 );
not ( n254140 , n240471 );
not ( n254141 , n252644 );
or ( n254142 , n254140 , n254141 );
not ( n254143 , n240471 );
nand ( n254144 , n254143 , n252649 );
nand ( n254145 , n254142 , n254144 );
and ( n254146 , n254145 , n252652 );
not ( n254147 , n254145 );
and ( n254148 , n254147 , n252656 );
nor ( n254149 , n254146 , n254148 );
not ( n254150 , n222532 );
nor ( n254151 , n254149 , n254150 );
not ( n254152 , n254151 );
not ( n254153 , n239276 );
not ( n254154 , n248755 );
or ( n254155 , n254153 , n254154 );
not ( n254156 , n239276 );
nand ( n254157 , n254156 , n248762 );
nand ( n254158 , n254155 , n254157 );
and ( n254159 , n254158 , n252923 );
not ( n254160 , n254158 );
and ( n254161 , n254160 , n252924 );
nor ( n254162 , n254159 , n254161 );
not ( n254163 , n254162 );
not ( n254164 , n240008 );
not ( n254165 , n40194 );
or ( n254166 , n254164 , n254165 );
not ( n254167 , n240008 );
nand ( n254168 , n254167 , n40203 );
nand ( n254169 , n254166 , n254168 );
and ( n254170 , n254169 , n251350 );
not ( n254171 , n254169 );
and ( n254172 , n254171 , n251346 );
nor ( n254173 , n254170 , n254172 );
nand ( n254174 , n254163 , n254173 );
or ( n254175 , n254152 , n254174 );
not ( n254176 , n254163 );
not ( n254177 , n254149 );
not ( n254178 , n254177 );
or ( n254179 , n254176 , n254178 );
nor ( n254180 , n254173 , n241065 );
nand ( n254181 , n254179 , n254180 );
nand ( n254182 , n239240 , n29821 );
nand ( n254183 , n254175 , n254181 , n254182 );
buf ( n254184 , n254183 );
not ( n254185 , RI19acadd8_2249);
or ( n254186 , n25328 , n254185 );
not ( n254187 , RI19ac1850_2318);
or ( n254188 , n226822 , n254187 );
nand ( n254189 , n254186 , n254188 );
buf ( n254190 , n254189 );
not ( n254191 , n239758 );
not ( n254192 , n239107 );
or ( n254193 , n254191 , n254192 );
not ( n254194 , n239758 );
nand ( n254195 , n254194 , n239099 );
nand ( n254196 , n254193 , n254195 );
and ( n254197 , n254196 , n242069 );
not ( n254198 , n254196 );
not ( n254199 , n242069 );
and ( n254200 , n254198 , n254199 );
nor ( n254201 , n254197 , n254200 );
not ( n254202 , n254201 );
not ( n254203 , n43013 );
nand ( n254204 , n254202 , n254203 );
not ( n254205 , n42444 );
or ( n254206 , n254204 , n254205 );
nor ( n254207 , n43513 , n221279 );
nand ( n254208 , n254204 , n254207 );
nand ( n254209 , n234024 , n39626 );
nand ( n254210 , n254206 , n254208 , n254209 );
buf ( n254211 , n254210 );
buf ( n254212 , n28181 );
buf ( n254213 , n33606 );
not ( n254214 , n240270 );
not ( n254215 , n254214 );
not ( n254216 , n252051 );
or ( n254217 , n254215 , n254216 );
not ( n254218 , n254214 );
nand ( n254219 , n254218 , n252036 );
nand ( n254220 , n254217 , n254219 );
and ( n254221 , n254220 , n252649 );
not ( n254222 , n254220 );
buf ( n254223 , n252644 );
and ( n254224 , n254222 , n254223 );
nor ( n254225 , n254221 , n254224 );
buf ( n254226 , n233971 );
not ( n254227 , n254226 );
nand ( n254228 , n254225 , n254227 );
not ( n254229 , n244727 );
not ( n254230 , n241877 );
or ( n254231 , n254229 , n254230 );
not ( n254232 , n244727 );
nand ( n254233 , n254232 , n241884 );
nand ( n254234 , n254231 , n254233 );
buf ( n254235 , n238975 );
and ( n254236 , n254234 , n254235 );
not ( n254237 , n254234 );
buf ( n254238 , n238985 );
and ( n254239 , n254237 , n254238 );
nor ( n254240 , n254236 , n254239 );
not ( n254241 , n42071 );
not ( n254242 , n234243 );
or ( n254243 , n254241 , n254242 );
not ( n254244 , n42071 );
nand ( n254245 , n254244 , n234252 );
nand ( n254246 , n254243 , n254245 );
and ( n254247 , n254246 , n234306 );
not ( n254248 , n254246 );
and ( n254249 , n254248 , n234299 );
nor ( n254250 , n254247 , n254249 );
nand ( n254251 , n254240 , n254250 );
or ( n254252 , n254228 , n254251 );
not ( n254253 , n254250 );
not ( n254254 , n254225 );
or ( n254255 , n254253 , n254254 );
nor ( n254256 , n254240 , n37725 );
nand ( n254257 , n254255 , n254256 );
nand ( n254258 , n49054 , n38978 );
nand ( n254259 , n254252 , n254257 , n254258 );
buf ( n254260 , n254259 );
not ( n254261 , n236354 );
not ( n254262 , n244582 );
or ( n254263 , n254261 , n254262 );
nand ( n254264 , n244583 , n236353 );
nand ( n254265 , n254263 , n254264 );
and ( n254266 , n254265 , n241255 );
not ( n254267 , n254265 );
and ( n254268 , n254267 , n244586 );
nor ( n254269 , n254266 , n254268 );
not ( n254270 , n254269 );
nand ( n254271 , n254270 , n241373 );
not ( n254272 , n236162 );
not ( n254273 , n236119 );
or ( n254274 , n254272 , n254273 );
nand ( n254275 , n254274 , n236165 );
and ( n254276 , n238241 , n254275 );
not ( n254277 , n238241 );
not ( n254278 , n254275 );
and ( n254279 , n254277 , n254278 );
nor ( n254280 , n254276 , n254279 );
nand ( n254281 , n53882 , n238331 );
not ( n254282 , n254281 );
not ( n254283 , n245018 );
and ( n254284 , n254282 , n254283 );
and ( n254285 , n254281 , n245018 );
nor ( n254286 , n254284 , n254285 );
not ( n254287 , n254286 );
not ( n254288 , n231615 );
nand ( n254289 , n238311 , n254288 );
buf ( n254290 , n245031 );
and ( n254291 , n254289 , n254290 );
not ( n254292 , n254289 );
not ( n254293 , n254290 );
and ( n254294 , n254292 , n254293 );
nor ( n254295 , n254291 , n254294 );
not ( n254296 , n254295 );
or ( n254297 , n254287 , n254296 );
or ( n254298 , n254295 , n254286 );
nand ( n254299 , n254297 , n254298 );
not ( n254300 , n238352 );
nand ( n254301 , n254300 , n231675 );
not ( n254302 , n254301 );
not ( n254303 , n245062 );
and ( n254304 , n254302 , n254303 );
and ( n254305 , n254301 , n245062 );
nor ( n254306 , n254304 , n254305 );
and ( n254307 , n254299 , n254306 );
not ( n254308 , n254299 );
not ( n254309 , n254306 );
and ( n254310 , n254308 , n254309 );
nor ( n254311 , n254307 , n254310 );
not ( n254312 , n254311 );
nand ( n254313 , n53992 , n238386 );
and ( n254314 , n254313 , n250984 );
not ( n254315 , n254313 );
and ( n254316 , n254315 , n245081 );
nor ( n254317 , n254314 , n254316 );
not ( n254318 , n254317 );
not ( n254319 , n238367 );
nand ( n254320 , n254319 , n53922 );
not ( n254321 , n254320 );
not ( n254322 , n245093 );
and ( n254323 , n254321 , n254322 );
not ( n254324 , n238367 );
nand ( n254325 , n254324 , n53922 );
and ( n254326 , n254325 , n245093 );
nor ( n254327 , n254323 , n254326 );
not ( n254328 , n254327 );
or ( n254329 , n254318 , n254328 );
or ( n254330 , n254327 , n254317 );
nand ( n254331 , n254329 , n254330 );
not ( n254332 , n254331 );
or ( n254333 , n254312 , n254332 );
not ( n254334 , n254331 );
not ( n254335 , n254311 );
nand ( n254336 , n254334 , n254335 );
nand ( n254337 , n254333 , n254336 );
and ( n254338 , n254280 , n254337 );
not ( n254339 , n254280 );
not ( n254340 , n254334 );
not ( n254341 , n254335 );
and ( n254342 , n254340 , n254341 );
and ( n254343 , n254334 , n254335 );
nor ( n254344 , n254342 , n254343 );
and ( n254345 , n254339 , n254344 );
nor ( n254346 , n254338 , n254345 );
not ( n254347 , n244719 );
not ( n254348 , n241877 );
or ( n254349 , n254347 , n254348 );
not ( n254350 , n244719 );
nand ( n254351 , n254350 , n241884 );
nand ( n254352 , n254349 , n254351 );
and ( n254353 , n254352 , n254238 );
not ( n254354 , n254352 );
and ( n254355 , n254354 , n254235 );
nor ( n254356 , n254353 , n254355 );
nand ( n254357 , n254346 , n254356 );
or ( n254358 , n254271 , n254357 );
not ( n254359 , n254270 );
not ( n254360 , n254356 );
or ( n254361 , n254359 , n254360 );
nor ( n254362 , n254346 , n251361 );
nand ( n254363 , n254361 , n254362 );
nand ( n254364 , n234024 , n28810 );
nand ( n254365 , n254358 , n254363 , n254364 );
buf ( n254366 , n254365 );
not ( n254367 , n249316 );
not ( n254368 , n235202 );
or ( n254369 , n254367 , n254368 );
not ( n254370 , n249316 );
nand ( n254371 , n254370 , n235211 );
nand ( n254372 , n254369 , n254371 );
and ( n254373 , n254372 , n250721 );
not ( n254374 , n254372 );
not ( n254375 , n250721 );
and ( n254376 , n254374 , n254375 );
nor ( n254377 , n254373 , n254376 );
not ( n254378 , n254377 );
not ( n254379 , n242741 );
not ( n254380 , n254379 );
not ( n254381 , n242977 );
or ( n254382 , n254380 , n254381 );
nand ( n254383 , n242969 , n242741 );
nand ( n254384 , n254382 , n254383 );
not ( n254385 , n254384 );
not ( n254386 , n254060 );
and ( n254387 , n254385 , n254386 );
and ( n254388 , n254384 , n254060 );
nor ( n254389 , n254387 , n254388 );
not ( n254390 , n254389 );
not ( n254391 , n254390 );
or ( n254392 , n254378 , n254391 );
not ( n254393 , n49532 );
not ( n254394 , n247187 );
or ( n254395 , n254393 , n254394 );
not ( n254396 , n49532 );
nand ( n254397 , n254396 , n247195 );
nand ( n254398 , n254395 , n254397 );
not ( n254399 , n240684 );
not ( n254400 , n254399 );
and ( n254401 , n254398 , n254400 );
not ( n254402 , n254398 );
buf ( n254403 , n240676 );
and ( n254404 , n254402 , n254403 );
nor ( n254405 , n254401 , n254404 );
not ( n254406 , n254405 );
nor ( n254407 , n254406 , n226003 );
nand ( n254408 , n254392 , n254407 );
nor ( n254409 , n254389 , n234440 );
not ( n254410 , n254377 );
nor ( n254411 , n254405 , n254410 );
nand ( n254412 , n254409 , n254411 );
nand ( n254413 , n251465 , n238538 );
nand ( n254414 , n254408 , n254412 , n254413 );
buf ( n254415 , n254414 );
not ( n254416 , RI19a946e8_2651);
or ( n254417 , n25328 , n254416 );
not ( n254418 , RI19a8a878_2721);
or ( n254419 , n25335 , n254418 );
nand ( n254420 , n254417 , n254419 );
buf ( n254421 , n254420 );
not ( n254422 , RI19ac9de8_2256);
or ( n254423 , n25328 , n254422 );
not ( n254424 , RI19ac0ba8_2325);
or ( n254425 , n25336 , n254424 );
nand ( n254426 , n254423 , n254425 );
buf ( n254427 , n254426 );
not ( n254428 , RI19aa8080_2509);
or ( n254429 , n226819 , n254428 );
not ( n254430 , RI19a9e8a0_2580);
or ( n254431 , n25336 , n254430 );
nand ( n254432 , n254429 , n254431 );
buf ( n254433 , n254432 );
not ( n254434 , RI19ac4f28_2292);
or ( n254435 , n25328 , n254434 );
not ( n254436 , RI19a85058_2759);
or ( n254437 , n25335 , n254436 );
nand ( n254438 , n254435 , n254437 );
buf ( n254439 , n254438 );
not ( n254440 , n26011 );
buf ( n254441 , n35431 );
not ( n254442 , n254441 );
or ( n254443 , n254440 , n254442 );
not ( n254444 , n54101 );
not ( n254445 , n242315 );
or ( n254446 , n254444 , n254445 );
or ( n254447 , n242315 , n54101 );
nand ( n254448 , n254446 , n254447 );
and ( n254449 , n254448 , n242380 );
not ( n254450 , n254448 );
and ( n254451 , n254450 , n242374 );
nor ( n254452 , n254449 , n254451 );
nand ( n254453 , n244780 , n254452 );
not ( n254454 , n245985 );
not ( n254455 , n224924 );
or ( n254456 , n254454 , n254455 );
not ( n254457 , n245985 );
nand ( n254458 , n254457 , n47156 );
nand ( n254459 , n254456 , n254458 );
and ( n254460 , n254459 , n245680 );
not ( n254461 , n254459 );
buf ( n254462 , n245677 );
and ( n254463 , n254461 , n254462 );
nor ( n254464 , n254460 , n254463 );
not ( n254465 , n254464 );
and ( n254466 , n254453 , n254465 );
not ( n254467 , n254453 );
and ( n254468 , n254467 , n254464 );
nor ( n254469 , n254466 , n254468 );
buf ( n254470 , n251862 );
or ( n254471 , n254469 , n254470 );
nand ( n254472 , n254443 , n254471 );
buf ( n254473 , n254472 );
not ( n254474 , n219510 );
not ( n254475 , n55760 );
or ( n254476 , n254474 , n254475 );
not ( n254477 , n248334 );
not ( n254478 , n246321 );
or ( n254479 , n254477 , n254478 );
not ( n254480 , n248334 );
nand ( n254481 , n254480 , n246326 );
nand ( n254482 , n254479 , n254481 );
buf ( n254483 , n51549 );
and ( n254484 , n254482 , n254483 );
not ( n254485 , n254482 );
and ( n254486 , n254485 , n246331 );
nor ( n254487 , n254484 , n254486 );
not ( n254488 , n254487 );
not ( n254489 , n228325 );
not ( n254490 , n31560 );
or ( n254491 , n254489 , n254490 );
not ( n254492 , n228325 );
nand ( n254493 , n254492 , n209312 );
nand ( n254494 , n254491 , n254493 );
and ( n254495 , n254494 , n35813 );
not ( n254496 , n254494 );
and ( n254497 , n254496 , n35805 );
nor ( n254498 , n254495 , n254497 );
nand ( n254499 , n254488 , n254498 );
buf ( n254500 , n241218 );
not ( n254501 , n254500 );
not ( n254502 , n250705 );
or ( n254503 , n254501 , n254502 );
or ( n254504 , n250705 , n254500 );
nand ( n254505 , n254503 , n254504 );
and ( n254506 , n254505 , n250709 );
not ( n254507 , n254505 );
and ( n254508 , n254507 , n250712 );
nor ( n254509 , n254506 , n254508 );
not ( n254510 , n254509 );
and ( n254511 , n254499 , n254510 );
not ( n254512 , n254499 );
and ( n254513 , n254512 , n254509 );
nor ( n254514 , n254511 , n254513 );
buf ( n254515 , n40465 );
or ( n254516 , n254514 , n254515 );
nand ( n254517 , n254476 , n254516 );
buf ( n254518 , n254517 );
not ( n254519 , n48708 );
not ( n254520 , n239228 );
or ( n254521 , n254519 , n254520 );
or ( n254522 , n239228 , n48708 );
nand ( n254523 , n254521 , n254522 );
and ( n254524 , n254523 , n250577 );
not ( n254525 , n254523 );
and ( n254526 , n254525 , n250580 );
nor ( n254527 , n254524 , n254526 );
not ( n254528 , n37725 );
nand ( n254529 , n254527 , n254528 );
not ( n254530 , n54896 );
not ( n254531 , n237936 );
or ( n254532 , n254530 , n254531 );
not ( n254533 , n54896 );
nand ( n254534 , n254533 , n237944 );
nand ( n254535 , n254532 , n254534 );
and ( n254536 , n254535 , n237948 );
not ( n254537 , n254535 );
and ( n254538 , n254537 , n237947 );
nor ( n254539 , n254536 , n254538 );
nand ( n254540 , n49028 , n49015 );
and ( n254541 , n254540 , n38609 );
not ( n254542 , n254540 );
and ( n254543 , n254542 , n38610 );
nor ( n254544 , n254541 , n254543 );
not ( n254545 , n254544 );
nand ( n254546 , n226689 , n226701 );
not ( n254547 , n254546 );
not ( n254548 , n249417 );
not ( n254549 , n254548 );
and ( n254550 , n254547 , n254549 );
and ( n254551 , n254546 , n254548 );
nor ( n254552 , n254550 , n254551 );
not ( n254553 , n254552 );
and ( n254554 , n254545 , n254553 );
and ( n254555 , n254544 , n254552 );
nor ( n254556 , n254554 , n254555 );
not ( n254557 , n48998 );
nand ( n254558 , n254557 , n48993 );
buf ( n254559 , n216261 );
not ( n254560 , n254559 );
and ( n254561 , n254558 , n254560 );
not ( n254562 , n254558 );
and ( n254563 , n254562 , n254559 );
nor ( n254564 , n254561 , n254563 );
not ( n254565 , n254564 );
and ( n254566 , n254556 , n254565 );
not ( n254567 , n254556 );
and ( n254568 , n254567 , n254564 );
nor ( n254569 , n254566 , n254568 );
nand ( n254570 , n226730 , n234461 );
not ( n254571 , n254570 );
not ( n254572 , n216226 );
or ( n254573 , n254571 , n254572 );
or ( n254574 , n216226 , n254570 );
nand ( n254575 , n254573 , n254574 );
not ( n254576 , n254575 );
not ( n254577 , n254576 );
nand ( n254578 , n48896 , n48914 );
not ( n254579 , n254578 );
buf ( n254580 , n38313 );
not ( n254581 , n254580 );
and ( n254582 , n254579 , n254581 );
and ( n254583 , n254578 , n254580 );
nor ( n254584 , n254582 , n254583 );
not ( n254585 , n254584 );
not ( n254586 , n254585 );
or ( n254587 , n254577 , n254586 );
nand ( n254588 , n254584 , n254575 );
nand ( n254589 , n254587 , n254588 );
and ( n254590 , n254569 , n254589 );
not ( n254591 , n254569 );
not ( n254592 , n254589 );
and ( n254593 , n254591 , n254592 );
nor ( n254594 , n254590 , n254593 );
and ( n254595 , n226708 , n254594 );
not ( n254596 , n226708 );
not ( n254597 , n254589 );
not ( n254598 , n254569 );
not ( n254599 , n254598 );
or ( n254600 , n254597 , n254599 );
nand ( n254601 , n254569 , n254592 );
nand ( n254602 , n254600 , n254601 );
not ( n254603 , n254602 );
and ( n254604 , n254596 , n254603 );
or ( n254605 , n254595 , n254604 );
not ( n254606 , n254605 );
not ( n254607 , n251619 );
not ( n254608 , n254607 );
not ( n254609 , n254608 );
and ( n254610 , n254606 , n254609 );
not ( n254611 , n254607 );
and ( n254612 , n254605 , n254611 );
nor ( n254613 , n254610 , n254612 );
nand ( n254614 , n254539 , n254613 );
or ( n254615 , n254529 , n254614 );
not ( n254616 , n254539 );
not ( n254617 , n254527 );
or ( n254618 , n254616 , n254617 );
nor ( n254619 , n254613 , n49051 );
nand ( n254620 , n254618 , n254619 );
nand ( n254621 , n234024 , n38365 );
nand ( n254622 , n254615 , n254620 , n254621 );
buf ( n254623 , n254622 );
not ( n254624 , n248756 );
not ( n254625 , n242168 );
not ( n254626 , n27876 );
or ( n254627 , n254625 , n254626 );
not ( n254628 , n242168 );
nand ( n254629 , n254628 , n27869 );
nand ( n254630 , n254627 , n254629 );
not ( n254631 , n254630 );
or ( n254632 , n254624 , n254631 );
or ( n254633 , n254630 , n248756 );
nand ( n254634 , n254632 , n254633 );
not ( n254635 , n254634 );
nor ( n254636 , n254635 , n252070 );
not ( n254637 , n254636 );
not ( n254638 , n36086 );
not ( n254639 , n249757 );
or ( n254640 , n254638 , n254639 );
not ( n254641 , n36086 );
nand ( n254642 , n254641 , n249749 );
nand ( n254643 , n254640 , n254642 );
buf ( n254644 , n253863 );
and ( n254645 , n254643 , n254644 );
not ( n254646 , n254643 );
buf ( n254647 , n253855 );
and ( n254648 , n254646 , n254647 );
nor ( n254649 , n254645 , n254648 );
not ( n254650 , n254649 );
not ( n254651 , n238855 );
not ( n254652 , n247500 );
or ( n254653 , n254651 , n254652 );
not ( n254654 , n238855 );
nand ( n254655 , n254654 , n247499 );
nand ( n254656 , n254653 , n254655 );
and ( n254657 , n254656 , n247563 );
not ( n254658 , n254656 );
and ( n254659 , n254658 , n247553 );
nor ( n254660 , n254657 , n254659 );
not ( n254661 , n254660 );
nand ( n254662 , n254650 , n254661 );
or ( n254663 , n254637 , n254662 );
not ( n254664 , n254634 );
not ( n254665 , n254650 );
or ( n254666 , n254664 , n254665 );
nor ( n254667 , n254661 , n250431 );
nand ( n254668 , n254666 , n254667 );
nand ( n254669 , n55760 , n38728 );
nand ( n254670 , n254663 , n254668 , n254669 );
buf ( n254671 , n254670 );
buf ( n254672 , n38085 );
buf ( n254673 , n32751 );
buf ( n254674 , n35851 );
not ( n254675 , n242352 );
not ( n254676 , n254675 );
not ( n254677 , n39749 );
or ( n254678 , n254676 , n254677 );
or ( n254679 , n217515 , n254675 );
nand ( n254680 , n254678 , n254679 );
not ( n254681 , n254680 );
nand ( n254682 , n243630 , n243644 );
not ( n254683 , n254682 );
not ( n254684 , n46365 );
and ( n254685 , n254683 , n254684 );
and ( n254686 , n254682 , n46365 );
nor ( n254687 , n254685 , n254686 );
not ( n254688 , n254687 );
not ( n254689 , n242992 );
nand ( n254690 , n254689 , n243613 );
and ( n254691 , n254690 , n46386 );
not ( n254692 , n254690 );
and ( n254693 , n254692 , n224148 );
nor ( n254694 , n254691 , n254693 );
not ( n254695 , n254694 );
or ( n254696 , n254688 , n254695 );
or ( n254697 , n254687 , n254694 );
nand ( n254698 , n254696 , n254697 );
not ( n254699 , n254698 );
not ( n254700 , n254699 );
nor ( n254701 , n243559 , n243548 );
not ( n254702 , n254701 );
not ( n254703 , n46278 );
and ( n254704 , n254702 , n254703 );
and ( n254705 , n254701 , n46278 );
nor ( n254706 , n254704 , n254705 );
not ( n254707 , n254706 );
not ( n254708 , n254707 );
nand ( n254709 , n243592 , n243580 );
and ( n254710 , n254709 , n46318 );
not ( n254711 , n254709 );
and ( n254712 , n254711 , n46319 );
nor ( n254713 , n254710 , n254712 );
not ( n254714 , n254713 );
not ( n254715 , n254714 );
or ( n254716 , n254708 , n254715 );
nand ( n254717 , n254713 , n254706 );
nand ( n254718 , n254716 , n254717 );
and ( n254719 , n254718 , n250132 );
not ( n254720 , n254718 );
not ( n254721 , n250132 );
and ( n254722 , n254720 , n254721 );
nor ( n254723 , n254719 , n254722 );
not ( n254724 , n254723 );
or ( n254725 , n254700 , n254724 );
not ( n254726 , n254723 );
nand ( n254727 , n254726 , n254698 );
nand ( n254728 , n254725 , n254727 );
buf ( n254729 , n254728 );
not ( n254730 , n254729 );
not ( n254731 , n254730 );
and ( n254732 , n254681 , n254731 );
and ( n254733 , n254680 , n254730 );
nor ( n254734 , n254732 , n254733 );
nor ( n254735 , n248800 , n254734 );
nor ( n254736 , n248786 , n235050 );
not ( n254737 , n254736 );
or ( n254738 , n254735 , n254737 );
not ( n254739 , n248786 );
not ( n254740 , n250111 );
nor ( n254741 , n254739 , n254740 );
nand ( n254742 , n254741 , n254735 );
nand ( n254743 , n241378 , n30294 );
nand ( n254744 , n254738 , n254742 , n254743 );
buf ( n254745 , n254744 );
not ( n254746 , n241080 );
not ( n254747 , n254746 );
not ( n254748 , n235580 );
or ( n254749 , n254747 , n254748 );
not ( n254750 , n254746 );
nand ( n254751 , n254750 , n235590 );
nand ( n254752 , n254749 , n254751 );
not ( n254753 , n254752 );
not ( n254754 , n235720 );
and ( n254755 , n254753 , n254754 );
and ( n254756 , n254752 , n235720 );
nor ( n254757 , n254755 , n254756 );
nor ( n254758 , n254757 , n249030 );
not ( n254759 , n254758 );
not ( n254760 , n245320 );
not ( n254761 , n242068 );
not ( n254762 , n254761 );
or ( n254763 , n254760 , n254762 );
or ( n254764 , n254761 , n245320 );
nand ( n254765 , n254763 , n254764 );
and ( n254766 , n254765 , n252239 );
not ( n254767 , n254765 );
and ( n254768 , n254767 , n252242 );
nor ( n254769 , n254766 , n254768 );
not ( n254770 , n254769 );
not ( n254771 , n31561 );
nand ( n254772 , n51666 , n229437 );
not ( n254773 , n254772 );
buf ( n254774 , n30545 );
not ( n254775 , n254774 );
and ( n254776 , n254773 , n254775 );
and ( n254777 , n254772 , n254774 );
nor ( n254778 , n254776 , n254777 );
not ( n254779 , n254778 );
not ( n254780 , n254779 );
not ( n254781 , n208725 );
or ( n254782 , n254780 , n254781 );
nand ( n254783 , n30968 , n254778 );
nand ( n254784 , n254782 , n254783 );
not ( n254785 , n254784 );
or ( n254786 , n254771 , n254785 );
or ( n254787 , n254784 , n31561 );
nand ( n254788 , n254786 , n254787 );
not ( n254789 , n254788 );
nand ( n254790 , n254770 , n254789 );
or ( n254791 , n254759 , n254790 );
not ( n254792 , n254770 );
not ( n254793 , n254757 );
not ( n254794 , n254793 );
or ( n254795 , n254792 , n254794 );
nor ( n254796 , n254789 , n49051 );
nand ( n254797 , n254795 , n254796 );
buf ( n254798 , n41944 );
nand ( n254799 , n254798 , n207918 );
nand ( n254800 , n254791 , n254797 , n254799 );
buf ( n254801 , n254800 );
not ( n254802 , n31796 );
not ( n254803 , n245701 );
or ( n254804 , n254802 , n254803 );
not ( n254805 , n235347 );
not ( n254806 , n246448 );
or ( n254807 , n254805 , n254806 );
not ( n254808 , n235347 );
nand ( n254809 , n254808 , n246439 );
nand ( n254810 , n254807 , n254809 );
buf ( n254811 , n250019 );
and ( n254812 , n254810 , n254811 );
not ( n254813 , n254810 );
and ( n254814 , n254813 , n250030 );
nor ( n254815 , n254812 , n254814 );
not ( n254816 , n254815 );
buf ( n254817 , n243388 );
not ( n254818 , n254817 );
not ( n254819 , n39052 );
or ( n254820 , n254818 , n254819 );
not ( n254821 , n254817 );
nand ( n254822 , n254821 , n39059 );
nand ( n254823 , n254820 , n254822 );
and ( n254824 , n254823 , n39435 );
not ( n254825 , n254823 );
and ( n254826 , n254825 , n39445 );
nor ( n254827 , n254824 , n254826 );
nand ( n254828 , n254816 , n254827 );
not ( n254829 , n242628 );
not ( n254830 , n254829 );
not ( n254831 , n244939 );
or ( n254832 , n254830 , n254831 );
not ( n254833 , n254829 );
nand ( n254834 , n254833 , n244954 );
nand ( n254835 , n254832 , n254834 );
nand ( n254836 , n244259 , n28292 );
not ( n254837 , n254836 );
not ( n254838 , n233856 );
and ( n254839 , n254837 , n254838 );
and ( n254840 , n254836 , n233856 );
nor ( n254841 , n254839 , n254840 );
nand ( n254842 , n28127 , n206369 );
not ( n254843 , n254842 );
not ( n254844 , n233848 );
and ( n254845 , n254843 , n254844 );
and ( n254846 , n254842 , n233848 );
nor ( n254847 , n254845 , n254846 );
xor ( n254848 , n254841 , n254847 );
xor ( n254849 , n254848 , n238207 );
nand ( n254850 , n28914 , n206593 );
and ( n254851 , n254850 , n33572 );
not ( n254852 , n254850 );
and ( n254853 , n254852 , n33571 );
nor ( n254854 , n254851 , n254853 );
not ( n254855 , n254854 );
not ( n254856 , n254855 );
not ( n254857 , n55340 );
not ( n254858 , n254857 );
or ( n254859 , n254856 , n254858 );
nand ( n254860 , n55340 , n254854 );
nand ( n254861 , n254859 , n254860 );
and ( n254862 , n254849 , n254861 );
not ( n254863 , n254849 );
not ( n254864 , n254861 );
and ( n254865 , n254863 , n254864 );
nor ( n254866 , n254862 , n254865 );
buf ( n254867 , n254866 );
and ( n254868 , n254835 , n254867 );
not ( n254869 , n254835 );
and ( n254870 , n254849 , n254864 );
not ( n254871 , n254849 );
and ( n254872 , n254871 , n254861 );
nor ( n254873 , n254870 , n254872 );
buf ( n254874 , n254873 );
and ( n254875 , n254869 , n254874 );
nor ( n254876 , n254868 , n254875 );
not ( n254877 , n254876 );
and ( n254878 , n254828 , n254877 );
not ( n254879 , n254828 );
and ( n254880 , n254879 , n254876 );
nor ( n254881 , n254878 , n254880 );
not ( n254882 , n205649 );
or ( n254883 , n254881 , n254882 );
nand ( n254884 , n254804 , n254883 );
buf ( n254885 , n254884 );
not ( n254886 , n49499 );
not ( n254887 , n254886 );
not ( n254888 , n247187 );
or ( n254889 , n254887 , n254888 );
not ( n254890 , n254886 );
nand ( n254891 , n254890 , n247195 );
nand ( n254892 , n254889 , n254891 );
and ( n254893 , n254892 , n254400 );
not ( n254894 , n254892 );
and ( n254895 , n254894 , n254403 );
nor ( n254896 , n254893 , n254895 );
not ( n254897 , n254896 );
not ( n254898 , n245478 );
not ( n254899 , n55067 );
or ( n254900 , n254898 , n254899 );
or ( n254901 , n55067 , n245478 );
nand ( n254902 , n254900 , n254901 );
not ( n254903 , n254902 );
not ( n254904 , n254903 );
not ( n254905 , n241966 );
or ( n254906 , n254904 , n254905 );
nand ( n254907 , n241963 , n254902 );
nand ( n254908 , n254906 , n254907 );
nand ( n254909 , n254897 , n254908 );
not ( n254910 , n237826 );
not ( n254911 , n254910 );
not ( n254912 , n251678 );
not ( n254913 , n251652 );
and ( n254914 , n254912 , n254913 );
and ( n254915 , n251652 , n251678 );
nor ( n254916 , n254914 , n254915 );
not ( n254917 , n254916 );
or ( n254918 , n254911 , n254917 );
not ( n254919 , n254910 );
nand ( n254920 , n254919 , n251684 );
nand ( n254921 , n254918 , n254920 );
xnor ( n254922 , n254921 , n251692 );
nand ( n254923 , n254922 , n205649 );
or ( n254924 , n254909 , n254923 );
not ( n254925 , n254908 );
not ( n254926 , n254922 );
or ( n254927 , n254925 , n254926 );
nand ( n254928 , n254927 , n235051 );
or ( n254929 , n254928 , n254897 );
nand ( n254930 , n252711 , n27781 );
nand ( n254931 , n254924 , n254929 , n254930 );
buf ( n254932 , n254931 );
buf ( n254933 , n225013 );
not ( n254934 , n254933 );
not ( n254935 , n254934 );
not ( n254936 , n245170 );
or ( n254937 , n254935 , n254936 );
nand ( n254938 , n254077 , n254933 );
nand ( n254939 , n254937 , n254938 );
and ( n254940 , n254939 , n254080 );
not ( n254941 , n254939 );
and ( n254942 , n254941 , n254083 );
nor ( n254943 , n254940 , n254942 );
nand ( n254944 , n254943 , n247275 );
not ( n254945 , n226147 );
not ( n254946 , n245676 );
not ( n254947 , n254946 );
not ( n254948 , n254947 );
or ( n254949 , n254945 , n254948 );
nand ( n254950 , n254946 , n48385 );
nand ( n254951 , n254949 , n254950 );
not ( n254952 , n254951 );
not ( n254953 , n251874 );
not ( n254954 , n254953 );
not ( n254955 , n236778 );
not ( n254956 , n254955 );
or ( n254957 , n254954 , n254956 );
nand ( n254958 , n236778 , n251874 );
nand ( n254959 , n254957 , n254958 );
xor ( n254960 , n234831 , n254959 );
not ( n254961 , n47733 );
not ( n254962 , n48483 );
nand ( n254963 , n254962 , n238015 );
not ( n254964 , n254963 );
or ( n254965 , n254961 , n254964 );
or ( n254966 , n254963 , n47733 );
nand ( n254967 , n254965 , n254966 );
not ( n254968 , n254967 );
not ( n254969 , n247706 );
or ( n254970 , n254968 , n254969 );
or ( n254971 , n247706 , n254967 );
nand ( n254972 , n254970 , n254971 );
xor ( n254973 , n254960 , n254972 );
buf ( n254974 , n254973 );
not ( n254975 , n254974 );
and ( n254976 , n254952 , n254975 );
and ( n254977 , n254951 , n254974 );
nor ( n254978 , n254976 , n254977 );
not ( n254979 , n238147 );
not ( n254980 , n45727 );
or ( n254981 , n254979 , n254980 );
not ( n254982 , n238147 );
nand ( n254983 , n254982 , n247727 );
nand ( n254984 , n254981 , n254983 );
and ( n254985 , n254984 , n247733 );
not ( n254986 , n254984 );
and ( n254987 , n254986 , n247730 );
nor ( n254988 , n254985 , n254987 );
nand ( n254989 , n254978 , n254988 );
or ( n254990 , n254944 , n254989 );
not ( n254991 , n254943 );
not ( n254992 , n254978 );
or ( n254993 , n254991 , n254992 );
nor ( n254994 , n254988 , n33253 );
nand ( n254995 , n254993 , n254994 );
nand ( n254996 , n41945 , n32636 );
nand ( n254997 , n254990 , n254995 , n254996 );
buf ( n254998 , n254997 );
not ( n254999 , n44327 );
buf ( n255000 , n244420 );
not ( n255001 , n255000 );
not ( n255002 , n247551 );
or ( n255003 , n255001 , n255002 );
or ( n255004 , n247551 , n255000 );
nand ( n255005 , n255003 , n255004 );
buf ( n255006 , n252317 );
xnor ( n255007 , n255005 , n255006 );
not ( n255008 , n255007 );
nand ( n255009 , n254999 , n255008 );
or ( n255010 , n43970 , n255009 );
not ( n255011 , n254999 );
not ( n255012 , n43967 );
or ( n255013 , n255011 , n255012 );
not ( n255014 , n205649 );
nor ( n255015 , n255008 , n255014 );
nand ( n255016 , n255013 , n255015 );
nand ( n255017 , n50615 , n41698 );
nand ( n255018 , n255010 , n255016 , n255017 );
buf ( n255019 , n255018 );
not ( n255020 , RI19aa90e8_2502);
or ( n255021 , n25328 , n255020 );
not ( n255022 , RI19a9f548_2574);
or ( n255023 , n25335 , n255022 );
nand ( n255024 , n255021 , n255023 );
buf ( n255025 , n255024 );
not ( n255026 , n247091 );
not ( n255027 , n253578 );
or ( n255028 , n255026 , n255027 );
not ( n255029 , n247091 );
nand ( n255030 , n255029 , n253463 );
nand ( n255031 , n255028 , n255030 );
and ( n255032 , n255031 , n253475 );
not ( n255033 , n255031 );
and ( n255034 , n255033 , n253478 );
nor ( n255035 , n255032 , n255034 );
not ( n255036 , n255035 );
not ( n255037 , n255036 );
not ( n255038 , n55213 );
not ( n255039 , n239390 );
or ( n255040 , n255038 , n255039 );
or ( n255041 , n239390 , n55213 );
nand ( n255042 , n255040 , n255041 );
and ( n255043 , n255042 , n249021 );
not ( n255044 , n255042 );
and ( n255045 , n255044 , n249018 );
nor ( n255046 , n255043 , n255045 );
not ( n255047 , n255046 );
or ( n255048 , n255037 , n255047 );
not ( n255049 , n253082 );
nor ( n255050 , n255049 , n250431 );
nand ( n255051 , n255048 , n255050 );
nor ( n255052 , n255035 , n55146 );
nand ( n255053 , n255052 , n255046 , n255049 );
nand ( n255054 , n241068 , n38306 );
nand ( n255055 , n255051 , n255053 , n255054 );
buf ( n255056 , n255055 );
not ( n255057 , n233910 );
not ( n255058 , n244336 );
or ( n255059 , n255057 , n255058 );
not ( n255060 , n233910 );
nand ( n255061 , n255060 , n244346 );
nand ( n255062 , n255059 , n255061 );
and ( n255063 , n255062 , n244472 );
not ( n255064 , n255062 );
and ( n255065 , n255064 , n244475 );
nor ( n255066 , n255063 , n255065 );
nand ( n255067 , n255066 , n33255 );
and ( n255068 , n46146 , n46186 );
not ( n255069 , n46146 );
and ( n255070 , n255069 , n46185 );
nor ( n255071 , n255068 , n255070 );
not ( n255072 , n255071 );
not ( n255073 , n255072 );
not ( n255074 , n255073 );
not ( n255075 , n34662 );
not ( n255076 , n240993 );
not ( n255077 , n240994 );
and ( n255078 , n255076 , n255077 );
and ( n255079 , n240993 , n240994 );
nor ( n255080 , n255078 , n255079 );
not ( n255081 , n255080 );
or ( n255082 , n255075 , n255081 );
not ( n255083 , n34661 );
or ( n255084 , n240996 , n255083 );
nand ( n255085 , n255082 , n255084 );
not ( n255086 , n255085 );
or ( n255087 , n255074 , n255086 );
not ( n255088 , n255071 );
not ( n255089 , n255088 );
or ( n255090 , n255089 , n255085 );
nand ( n255091 , n255087 , n255090 );
not ( n255092 , n255091 );
buf ( n255093 , n242346 );
not ( n255094 , n255093 );
not ( n255095 , n217514 );
or ( n255096 , n255094 , n255095 );
or ( n255097 , n39749 , n255093 );
nand ( n255098 , n255096 , n255097 );
not ( n255099 , n255098 );
not ( n255100 , n254728 );
not ( n255101 , n255100 );
and ( n255102 , n255099 , n255101 );
and ( n255103 , n255098 , n255100 );
nor ( n255104 , n255102 , n255103 );
nand ( n255105 , n255092 , n255104 );
or ( n255106 , n255067 , n255105 );
not ( n255107 , n255092 );
not ( n255108 , n255066 );
or ( n255109 , n255107 , n255108 );
nor ( n255110 , n255104 , n235895 );
nand ( n255111 , n255109 , n255110 );
nand ( n255112 , n31577 , n29043 );
nand ( n255113 , n255106 , n255111 , n255112 );
buf ( n255114 , n255113 );
not ( n255115 , n28760 );
buf ( n255116 , n41944 );
not ( n255117 , n255116 );
or ( n255118 , n255115 , n255117 );
nand ( n255119 , n243664 , n243513 );
not ( n255120 , n236309 );
not ( n255121 , n244574 );
not ( n255122 , n255121 );
or ( n255123 , n255120 , n255122 );
or ( n255124 , n255121 , n236309 );
nand ( n255125 , n255123 , n255124 );
and ( n255126 , n255125 , n244587 );
not ( n255127 , n255125 );
and ( n255128 , n255127 , n244591 );
nor ( n255129 , n255126 , n255128 );
and ( n255130 , n255119 , n255129 );
not ( n255131 , n255119 );
not ( n255132 , n255129 );
and ( n255133 , n255131 , n255132 );
nor ( n255134 , n255130 , n255133 );
buf ( n255135 , n254150 );
or ( n255136 , n255134 , n255135 );
nand ( n255137 , n255118 , n255136 );
buf ( n255138 , n255137 );
not ( n255139 , n237788 );
not ( n255140 , n255139 );
not ( n255141 , n245392 );
or ( n255142 , n255140 , n255141 );
not ( n255143 , n255139 );
nand ( n255144 , n255143 , n245402 );
nand ( n255145 , n255142 , n255144 );
buf ( n255146 , n254916 );
and ( n255147 , n255145 , n255146 );
not ( n255148 , n255145 );
buf ( n255149 , n251684 );
and ( n255150 , n255148 , n255149 );
nor ( n255151 , n255147 , n255150 );
not ( n255152 , n35427 );
nand ( n255153 , n255151 , n255152 );
not ( n255154 , n242201 );
buf ( n255155 , n236870 );
not ( n255156 , n255155 );
and ( n255157 , n255154 , n255156 );
and ( n255158 , n242205 , n255155 );
nor ( n255159 , n255157 , n255158 );
buf ( n255160 , n239298 );
and ( n255161 , n255159 , n255160 );
not ( n255162 , n255159 );
buf ( n255163 , n239297 );
and ( n255164 , n255162 , n255163 );
nor ( n255165 , n255161 , n255164 );
not ( n255166 , n255165 );
nor ( n255167 , n255153 , n255166 );
not ( n255168 , n255167 );
nor ( n255169 , n255151 , n46425 );
not ( n255170 , n43011 );
not ( n255171 , n252159 );
not ( n255172 , n220460 );
or ( n255173 , n255171 , n255172 );
not ( n255174 , n252159 );
nand ( n255175 , n255174 , n220467 );
nand ( n255176 , n255173 , n255175 );
not ( n255177 , n255176 );
or ( n255178 , n255170 , n255177 );
or ( n255179 , n255176 , n43011 );
nand ( n255180 , n255178 , n255179 );
not ( n255181 , n255180 );
nand ( n255182 , n255169 , n255181 , n255166 );
not ( n255183 , n255165 );
nor ( n255184 , n255183 , n226003 );
nand ( n255185 , n255184 , n255180 );
nand ( n255186 , n251465 , n228982 );
nand ( n255187 , n255168 , n255182 , n255185 , n255186 );
buf ( n255188 , n255187 );
not ( n255189 , RI19ab9df8_2381);
or ( n255190 , n25328 , n255189 );
not ( n255191 , RI19a83d20_2767);
or ( n255192 , n25336 , n255191 );
nand ( n255193 , n255190 , n255192 );
buf ( n255194 , n255193 );
not ( n255195 , n245958 );
not ( n255196 , n255195 );
not ( n255197 , n224924 );
or ( n255198 , n255196 , n255197 );
not ( n255199 , n255195 );
nand ( n255200 , n255199 , n47156 );
nand ( n255201 , n255198 , n255200 );
and ( n255202 , n255201 , n245680 );
not ( n255203 , n255201 );
and ( n255204 , n255203 , n254462 );
nor ( n255205 , n255202 , n255204 );
nor ( n255206 , n255205 , n235050 );
not ( n255207 , n34429 );
not ( n255208 , n244190 );
or ( n255209 , n255207 , n255208 );
not ( n255210 , n34429 );
nand ( n255211 , n255210 , n244199 );
nand ( n255212 , n255209 , n255211 );
not ( n255213 , n244204 );
and ( n255214 , n255212 , n255213 );
not ( n255215 , n255212 );
and ( n255216 , n255215 , n244204 );
nor ( n255217 , n255214 , n255216 );
nand ( n255218 , n255206 , n255217 );
not ( n255219 , n205649 );
not ( n255220 , n30227 );
not ( n255221 , n246963 );
or ( n255222 , n255220 , n255221 );
not ( n255223 , n30227 );
nand ( n255224 , n255223 , n246968 );
nand ( n255225 , n255222 , n255224 );
and ( n255226 , n255225 , n247014 );
not ( n255227 , n255225 );
and ( n255228 , n255227 , n247019 );
nor ( n255229 , n255226 , n255228 );
nor ( n255230 , n255219 , n255229 );
not ( n255231 , n255205 );
nand ( n255232 , n255230 , n255231 );
not ( n255233 , n255229 );
nor ( n255234 , n255233 , n221279 );
not ( n255235 , n255217 );
nand ( n255236 , n255234 , n255235 , n255205 );
nand ( n255237 , n48251 , n204575 );
nand ( n255238 , n255218 , n255232 , n255236 , n255237 );
buf ( n255239 , n255238 );
not ( n255240 , n246728 );
not ( n255241 , n45253 );
or ( n255242 , n255240 , n255241 );
or ( n255243 , n45253 , n246728 );
nand ( n255244 , n255242 , n255243 );
buf ( n255245 , n232514 );
and ( n255246 , n255244 , n255245 );
not ( n255247 , n255244 );
buf ( n255248 , n232520 );
and ( n255249 , n255247 , n255248 );
nor ( n255250 , n255246 , n255249 );
nand ( n255251 , n255250 , n43969 );
not ( n255252 , n237855 );
not ( n255253 , n255146 );
or ( n255254 , n255252 , n255253 );
not ( n255255 , n237855 );
nand ( n255256 , n255255 , n251684 );
nand ( n255257 , n255254 , n255256 );
and ( n255258 , n255257 , n251689 );
not ( n255259 , n255257 );
and ( n255260 , n255259 , n251693 );
nor ( n255261 , n255258 , n255260 );
not ( n255262 , n255261 );
not ( n255263 , n247511 );
not ( n255264 , n255263 );
not ( n255265 , n243801 );
or ( n255266 , n255264 , n255265 );
not ( n255267 , n255263 );
nand ( n255268 , n255267 , n243810 );
nand ( n255269 , n255266 , n255268 );
and ( n255270 , n255269 , n243960 );
not ( n255271 , n255269 );
and ( n255272 , n255271 , n243954 );
nor ( n255273 , n255270 , n255272 );
nand ( n255274 , n255262 , n255273 );
or ( n255275 , n255251 , n255274 );
not ( n255276 , n255262 );
not ( n255277 , n255250 );
or ( n255278 , n255276 , n255277 );
nor ( n255279 , n255273 , n31572 );
nand ( n255280 , n255278 , n255279 );
nand ( n255281 , n46083 , n35777 );
nand ( n255282 , n255275 , n255280 , n255281 );
buf ( n255283 , n255282 );
not ( n255284 , n32671 );
not ( n255285 , n31577 );
or ( n255286 , n255284 , n255285 );
not ( n255287 , n53545 );
not ( n255288 , n250496 );
or ( n255289 , n255287 , n255288 );
xor ( n255290 , n250471 , n250491 );
xor ( n255291 , n255290 , n250466 );
nand ( n255292 , n255291 , n53546 );
nand ( n255293 , n255289 , n255292 );
not ( n255294 , n244190 );
not ( n255295 , n255294 );
xor ( n255296 , n255293 , n255295 );
not ( n255297 , n46614 );
not ( n255298 , n253196 );
or ( n255299 , n255297 , n255298 );
not ( n255300 , n46614 );
nand ( n255301 , n255300 , n253188 );
nand ( n255302 , n255299 , n255301 );
buf ( n255303 , n248056 );
and ( n255304 , n255302 , n255303 );
not ( n255305 , n255302 );
and ( n255306 , n255305 , n253948 );
nor ( n255307 , n255304 , n255306 );
not ( n255308 , n255307 );
nand ( n255309 , n255296 , n255308 );
not ( n255310 , n41090 );
not ( n255311 , n54263 );
or ( n255312 , n255310 , n255311 );
not ( n255313 , n41090 );
nand ( n255314 , n255313 , n54273 );
nand ( n255315 , n255312 , n255314 );
not ( n255316 , n232084 );
not ( n255317 , n54300 );
or ( n255318 , n255316 , n255317 );
nand ( n255319 , n54301 , n54320 );
nand ( n255320 , n255318 , n255319 );
buf ( n255321 , n255320 );
and ( n255322 , n255315 , n255321 );
not ( n255323 , n255315 );
buf ( n255324 , n54325 );
and ( n255325 , n255323 , n255324 );
nor ( n255326 , n255322 , n255325 );
and ( n255327 , n255309 , n255326 );
not ( n255328 , n255309 );
not ( n255329 , n255326 );
and ( n255330 , n255328 , n255329 );
nor ( n255331 , n255327 , n255330 );
or ( n255332 , n255331 , n238223 );
nand ( n255333 , n255286 , n255332 );
buf ( n255334 , n255333 );
not ( n255335 , n38267 );
not ( n255336 , n51381 );
or ( n255337 , n255335 , n255336 );
not ( n255338 , n233399 );
not ( n255339 , n235008 );
or ( n255340 , n255338 , n255339 );
not ( n255341 , n233399 );
nand ( n255342 , n255341 , n235016 );
nand ( n255343 , n255340 , n255342 );
and ( n255344 , n255343 , n235022 );
not ( n255345 , n255343 );
and ( n255346 , n255345 , n235019 );
nor ( n255347 , n255344 , n255346 );
not ( n255348 , n240141 );
not ( n255349 , n239199 );
and ( n255350 , n255348 , n255349 );
and ( n255351 , n240141 , n239199 );
nor ( n255352 , n255350 , n255351 );
buf ( n255353 , n227174 );
and ( n255354 , n255352 , n255353 );
not ( n255355 , n255352 );
buf ( n255356 , n49420 );
and ( n255357 , n255355 , n255356 );
nor ( n255358 , n255354 , n255357 );
nand ( n255359 , n255347 , n255358 );
not ( n255360 , n230999 );
not ( n255361 , n253669 );
or ( n255362 , n255360 , n255361 );
not ( n255363 , n230999 );
nand ( n255364 , n255363 , n253673 );
nand ( n255365 , n255362 , n255364 );
and ( n255366 , n255365 , n253676 );
not ( n255367 , n255365 );
and ( n255368 , n255367 , n253679 );
nor ( n255369 , n255366 , n255368 );
not ( n255370 , n255369 );
and ( n255371 , n255359 , n255370 );
not ( n255372 , n255359 );
and ( n255373 , n255372 , n255369 );
nor ( n255374 , n255371 , n255373 );
or ( n255375 , n255374 , n31572 );
nand ( n255376 , n255337 , n255375 );
buf ( n255377 , n255376 );
not ( n255378 , n32244 );
not ( n255379 , n254441 );
or ( n255380 , n255378 , n255379 );
not ( n255381 , n230903 );
not ( n255382 , n55316 );
not ( n255383 , n53080 );
or ( n255384 , n255382 , n255383 );
not ( n255385 , n53076 );
nand ( n255386 , n255385 , n55315 );
nand ( n255387 , n255384 , n255386 );
not ( n255388 , n255387 );
or ( n255389 , n255381 , n255388 );
or ( n255390 , n255387 , n230906 );
nand ( n255391 , n255389 , n255390 );
not ( n255392 , n251121 );
not ( n255393 , n242520 );
or ( n255394 , n255392 , n255393 );
not ( n255395 , n251121 );
nand ( n255396 , n255395 , n242527 );
nand ( n255397 , n255394 , n255396 );
and ( n255398 , n255397 , n242571 );
not ( n255399 , n255397 );
and ( n255400 , n255399 , n242575 );
nor ( n255401 , n255398 , n255400 );
not ( n255402 , n255401 );
nand ( n255403 , n255391 , n255402 );
not ( n255404 , n246523 );
not ( n255405 , n236449 );
not ( n255406 , n236498 );
or ( n255407 , n255405 , n255406 );
nand ( n255408 , n255407 , n236501 );
not ( n255409 , n255408 );
or ( n255410 , n255404 , n255409 );
or ( n255411 , n236502 , n246523 );
nand ( n255412 , n255410 , n255411 );
not ( n255413 , n53167 );
nand ( n255414 , n32691 , n246630 );
not ( n255415 , n255414 );
or ( n255416 , n255413 , n255415 );
or ( n255417 , n255414 , n53167 );
nand ( n255418 , n255416 , n255417 );
not ( n255419 , n255418 );
not ( n255420 , n32530 );
nand ( n255421 , n255420 , n253627 );
not ( n255422 , n255421 );
buf ( n255423 , n32507 );
not ( n255424 , n255423 );
and ( n255425 , n255422 , n255424 );
not ( n255426 , n246614 );
nand ( n255427 , n255426 , n255420 );
and ( n255428 , n255427 , n255423 );
nor ( n255429 , n255425 , n255428 );
not ( n255430 , n255429 );
or ( n255431 , n255419 , n255430 );
or ( n255432 , n255429 , n255418 );
nand ( n255433 , n255431 , n255432 );
nand ( n255434 , n32864 , n246594 );
not ( n255435 , n255434 );
not ( n255436 , n53189 );
and ( n255437 , n255435 , n255436 );
and ( n255438 , n255434 , n53189 );
nor ( n255439 , n255437 , n255438 );
not ( n255440 , n255439 );
and ( n255441 , n255433 , n255440 );
not ( n255442 , n255433 );
and ( n255443 , n255442 , n255439 );
nor ( n255444 , n255441 , n255443 );
not ( n255445 , n255444 );
not ( n255446 , n253520 );
not ( n255447 , n253710 );
and ( n255448 , n255446 , n255447 );
and ( n255449 , n253520 , n253710 );
nor ( n255450 , n255448 , n255449 );
not ( n255451 , n255450 );
and ( n255452 , n255445 , n255451 );
not ( n255453 , n255445 );
and ( n255454 , n255453 , n255450 );
nor ( n255455 , n255452 , n255454 );
not ( n255456 , n255455 );
not ( n255457 , n255456 );
and ( n255458 , n255412 , n255457 );
not ( n255459 , n255412 );
not ( n255460 , n255450 );
not ( n255461 , n255444 );
or ( n255462 , n255460 , n255461 );
nand ( n255463 , n255445 , n255451 );
nand ( n255464 , n255462 , n255463 );
buf ( n255465 , n255464 );
and ( n255466 , n255459 , n255465 );
nor ( n255467 , n255458 , n255466 );
not ( n255468 , n255467 );
and ( n255469 , n255403 , n255468 );
not ( n255470 , n255403 );
and ( n255471 , n255470 , n255467 );
nor ( n255472 , n255469 , n255471 );
or ( n255473 , n255472 , n251498 );
nand ( n255474 , n255380 , n255473 );
buf ( n255475 , n255474 );
or ( n255476 , n233507 , n235064 );
not ( n255477 , RI19a9efa8_2577);
or ( n255478 , n25336 , n255477 );
nand ( n255479 , n255476 , n255478 );
buf ( n255480 , n255479 );
not ( n255481 , n37417 );
not ( n255482 , n51381 );
or ( n255483 , n255481 , n255482 );
not ( n255484 , n246797 );
not ( n255485 , n249927 );
or ( n255486 , n255484 , n255485 );
not ( n255487 , n246797 );
not ( n255488 , n249923 );
not ( n255489 , n249896 );
or ( n255490 , n255488 , n255489 );
not ( n255491 , n249896 );
nand ( n255492 , n255491 , n249922 );
nand ( n255493 , n255490 , n255492 );
nand ( n255494 , n255487 , n255493 );
nand ( n255495 , n255486 , n255494 );
not ( n255496 , n242859 );
not ( n255497 , n255496 );
and ( n255498 , n255495 , n255497 );
not ( n255499 , n255495 );
buf ( n255500 , n242860 );
and ( n255501 , n255499 , n255500 );
nor ( n255502 , n255498 , n255501 );
xor ( n255503 , n237848 , n237866 );
not ( n255504 , n255503 );
not ( n255505 , n50661 );
not ( n255506 , n255505 );
and ( n255507 , n255504 , n255506 );
not ( n255508 , n237867 );
and ( n255509 , n255508 , n255505 );
nor ( n255510 , n255507 , n255509 );
and ( n255511 , n251950 , n251966 );
not ( n255512 , n251950 );
and ( n255513 , n255512 , n251965 );
nor ( n255514 , n255511 , n255513 );
buf ( n255515 , n255514 );
xor ( n255516 , n255510 , n255515 );
nand ( n255517 , n255502 , n255516 );
not ( n255518 , n233968 );
not ( n255519 , n33622 );
not ( n255520 , n233904 );
or ( n255521 , n255519 , n255520 );
or ( n255522 , n244207 , n33622 );
nand ( n255523 , n255521 , n255522 );
not ( n255524 , n255523 );
or ( n255525 , n255518 , n255524 );
or ( n255526 , n255523 , n233968 );
nand ( n255527 , n255525 , n255526 );
not ( n255528 , n255527 );
and ( n255529 , n255517 , n255528 );
not ( n255530 , n255517 );
and ( n255531 , n255530 , n255527 );
or ( n255532 , n255529 , n255531 );
not ( n255533 , n222532 );
or ( n255534 , n255532 , n255533 );
nand ( n255535 , n255483 , n255534 );
buf ( n255536 , n255535 );
not ( n255537 , n248110 );
nand ( n255538 , n238581 , n235568 );
not ( n255539 , n255538 );
not ( n255540 , n241100 );
and ( n255541 , n255539 , n255540 );
and ( n255542 , n255538 , n241100 );
nor ( n255543 , n255541 , n255542 );
not ( n255544 , n255543 );
not ( n255545 , n255544 );
nand ( n255546 , n238602 , n235514 );
not ( n255547 , n255546 );
not ( n255548 , n241108 );
or ( n255549 , n255547 , n255548 );
or ( n255550 , n241108 , n255546 );
nand ( n255551 , n255549 , n255550 );
not ( n255552 , n255551 );
not ( n255553 , n255552 );
or ( n255554 , n255545 , n255553 );
nand ( n255555 , n255551 , n255543 );
nand ( n255556 , n255554 , n255555 );
not ( n255557 , n255556 );
not ( n255558 , n235400 );
nand ( n255559 , n235432 , n238518 );
not ( n255560 , n255559 );
or ( n255561 , n255558 , n255560 );
or ( n255562 , n255559 , n235400 );
nand ( n255563 , n255561 , n255562 );
nand ( n255564 , n238536 , n235467 );
not ( n255565 , n255564 );
not ( n255566 , n238553 );
and ( n255567 , n255565 , n255566 );
not ( n255568 , n235464 );
nand ( n255569 , n255568 , n238536 );
and ( n255570 , n255569 , n238553 );
nor ( n255571 , n255567 , n255570 );
and ( n255572 , n255563 , n255571 );
not ( n255573 , n255563 );
not ( n255574 , n255571 );
and ( n255575 , n255573 , n255574 );
nor ( n255576 , n255572 , n255575 );
not ( n255577 , n255576 );
nand ( n255578 , n248104 , n235494 );
xnor ( n255579 , n255578 , n238496 );
not ( n255580 , n255579 );
or ( n255581 , n255577 , n255580 );
or ( n255582 , n255579 , n255576 );
nand ( n255583 , n255581 , n255582 );
not ( n255584 , n255583 );
not ( n255585 , n255584 );
or ( n255586 , n255557 , n255585 );
not ( n255587 , n255556 );
nand ( n255588 , n255587 , n255583 );
nand ( n255589 , n255586 , n255588 );
not ( n255590 , n255589 );
or ( n255591 , n255537 , n255590 );
not ( n255592 , n248110 );
not ( n255593 , n255589 );
nand ( n255594 , n255592 , n255593 );
nand ( n255595 , n255591 , n255594 );
buf ( n255596 , n228918 );
and ( n255597 , n255595 , n255596 );
not ( n255598 , n255595 );
buf ( n255599 , n51167 );
and ( n255600 , n255598 , n255599 );
nor ( n255601 , n255597 , n255600 );
not ( n255602 , n255601 );
not ( n255603 , n248437 );
not ( n255604 , n221715 );
or ( n255605 , n255603 , n255604 );
not ( n255606 , n248437 );
nand ( n255607 , n255606 , n43962 );
nand ( n255608 , n255605 , n255607 );
buf ( n255609 , n246321 );
and ( n255610 , n255608 , n255609 );
not ( n255611 , n255608 );
buf ( n255612 , n246326 );
and ( n255613 , n255611 , n255612 );
nor ( n255614 , n255610 , n255613 );
nand ( n255615 , n255602 , n255614 );
not ( n255616 , n244566 );
not ( n255617 , n255616 );
not ( n255618 , n239705 );
or ( n255619 , n255617 , n255618 );
not ( n255620 , n255616 );
nand ( n255621 , n255620 , n239715 );
nand ( n255622 , n255619 , n255621 );
and ( n255623 , n255622 , n239775 );
not ( n255624 , n255622 );
buf ( n255625 , n250705 );
and ( n255626 , n255624 , n255625 );
nor ( n255627 , n255623 , n255626 );
nand ( n255628 , n255627 , n235051 );
or ( n255629 , n255615 , n255628 );
nor ( n255630 , n255627 , n243204 );
nand ( n255631 , n255615 , n255630 );
nand ( n255632 , n31576 , n26043 );
nand ( n255633 , n255629 , n255631 , n255632 );
buf ( n255634 , n255633 );
not ( n255635 , n35341 );
not ( n255636 , n51381 );
or ( n255637 , n255635 , n255636 );
not ( n255638 , n251414 );
not ( n255639 , n252132 );
or ( n255640 , n255638 , n255639 );
not ( n255641 , n251414 );
nand ( n255642 , n255641 , n252139 );
nand ( n255643 , n255640 , n255642 );
and ( n255644 , n255643 , n252186 );
not ( n255645 , n255643 );
and ( n255646 , n255645 , n252194 );
nor ( n255647 , n255644 , n255646 );
nand ( n255648 , n235890 , n255647 );
and ( n255649 , n255648 , n55069 );
not ( n255650 , n255648 );
not ( n255651 , n55069 );
and ( n255652 , n255650 , n255651 );
nor ( n255653 , n255649 , n255652 );
or ( n255654 , n255653 , n250068 );
nand ( n255655 , n255637 , n255654 );
buf ( n255656 , n255655 );
not ( n255657 , RI19a9fcc8_2570);
or ( n255658 , n25328 , n255657 );
not ( n255659 , RI19acf1d0_2217);
or ( n255660 , n25336 , n255659 );
nand ( n255661 , n255658 , n255660 );
buf ( n255662 , n255661 );
not ( n255663 , n32369 );
not ( n255664 , n46083 );
or ( n255665 , n255663 , n255664 );
not ( n255666 , n221658 );
not ( n255667 , n255666 );
not ( n255668 , n252552 );
or ( n255669 , n255667 , n255668 );
not ( n255670 , n255666 );
nand ( n255671 , n255670 , n252561 );
nand ( n255672 , n255669 , n255671 );
buf ( n255673 , n239607 );
and ( n255674 , n255672 , n255673 );
not ( n255675 , n255672 );
not ( n255676 , n255673 );
and ( n255677 , n255675 , n255676 );
nor ( n255678 , n255674 , n255677 );
not ( n255679 , n255678 );
not ( n255680 , n254730 );
not ( n255681 , n242333 );
not ( n255682 , n217511 );
or ( n255683 , n255681 , n255682 );
not ( n255684 , n242333 );
nand ( n255685 , n255684 , n39749 );
nand ( n255686 , n255683 , n255685 );
not ( n255687 , n255686 );
or ( n255688 , n255680 , n255687 );
or ( n255689 , n255686 , n254730 );
nand ( n255690 , n255688 , n255689 );
nand ( n255691 , n255679 , n255690 );
not ( n255692 , n39261 );
not ( n255693 , n246826 );
or ( n255694 , n255692 , n255693 );
not ( n255695 , n39261 );
nand ( n255696 , n255695 , n246835 );
nand ( n255697 , n255694 , n255696 );
and ( n255698 , n255697 , n246883 );
not ( n255699 , n255697 );
and ( n255700 , n255699 , n246892 );
nor ( n255701 , n255698 , n255700 );
not ( n255702 , n255701 );
and ( n255703 , n255691 , n255702 );
not ( n255704 , n255691 );
and ( n255705 , n255704 , n255701 );
nor ( n255706 , n255703 , n255705 );
buf ( n255707 , n55152 );
or ( n255708 , n255706 , n255707 );
nand ( n255709 , n255665 , n255708 );
buf ( n255710 , n255709 );
not ( n255711 , RI19ab0e10_2447);
or ( n255712 , n25328 , n255711 );
not ( n255713 , RI19aa6b68_2518);
or ( n255714 , n25336 , n255713 );
nand ( n255715 , n255712 , n255714 );
buf ( n255716 , n255715 );
nand ( n255717 , n51086 , n51075 );
not ( n255718 , n255717 );
not ( n255719 , n235693 );
and ( n255720 , n255718 , n255719 );
not ( n255721 , n241154 );
nand ( n255722 , n255721 , n51086 );
and ( n255723 , n255722 , n235693 );
nor ( n255724 , n255720 , n255723 );
not ( n255725 , n255724 );
and ( n255726 , n249539 , n255725 );
not ( n255727 , n249539 );
and ( n255728 , n255727 , n255724 );
nor ( n255729 , n255726 , n255728 );
not ( n255730 , n255729 );
not ( n255731 , n235658 );
nand ( n255732 , n51054 , n51045 );
not ( n255733 , n255732 );
or ( n255734 , n255731 , n255733 );
or ( n255735 , n255732 , n235658 );
nand ( n255736 , n255734 , n255735 );
not ( n255737 , n255736 );
nand ( n255738 , n228784 , n50979 );
not ( n255739 , n255738 );
not ( n255740 , n235602 );
and ( n255741 , n255739 , n255740 );
and ( n255742 , n255738 , n235602 );
nor ( n255743 , n255741 , n255742 );
not ( n255744 , n255743 );
or ( n255745 , n255737 , n255744 );
or ( n255746 , n255743 , n255736 );
nand ( n255747 , n255745 , n255746 );
not ( n255748 , n228767 );
nand ( n255749 , n255748 , n238417 );
buf ( n255750 , n235617 );
xor ( n255751 , n255749 , n255750 );
and ( n255752 , n255747 , n255751 );
not ( n255753 , n255747 );
not ( n255754 , n255751 );
and ( n255755 , n255753 , n255754 );
nor ( n255756 , n255752 , n255755 );
not ( n255757 , n255756 );
or ( n255758 , n255730 , n255757 );
not ( n255759 , n255756 );
not ( n255760 , n255729 );
nand ( n255761 , n255759 , n255760 );
nand ( n255762 , n255758 , n255761 );
not ( n255763 , n255762 );
buf ( n255764 , n51010 );
not ( n255765 , n255764 );
and ( n255766 , n255763 , n255765 );
and ( n255767 , n255762 , n255764 );
nor ( n255768 , n255766 , n255767 );
not ( n255769 , n31615 );
nand ( n255770 , n51199 , n31934 );
not ( n255771 , n255770 );
or ( n255772 , n255769 , n255771 );
or ( n255773 , n255770 , n31615 );
nand ( n255774 , n255772 , n255773 );
not ( n255775 , n255774 );
not ( n255776 , n246491 );
or ( n255777 , n255775 , n255776 );
or ( n255778 , n246491 , n255774 );
nand ( n255779 , n255777 , n255778 );
nand ( n255780 , n51208 , n32087 );
not ( n255781 , n255780 );
not ( n255782 , n246517 );
not ( n255783 , n255782 );
and ( n255784 , n255781 , n255783 );
and ( n255785 , n255780 , n255782 );
nor ( n255786 , n255784 , n255785 );
and ( n255787 , n255779 , n255786 );
not ( n255788 , n255779 );
not ( n255789 , n255786 );
and ( n255790 , n255788 , n255789 );
nor ( n255791 , n255787 , n255790 );
not ( n255792 , n247287 );
not ( n255793 , n255792 );
nand ( n255794 , n32365 , n228996 );
and ( n255795 , n255794 , n246529 );
not ( n255796 , n255794 );
and ( n255797 , n255796 , n236422 );
nor ( n255798 , n255795 , n255797 );
not ( n255799 , n255798 );
or ( n255800 , n255793 , n255799 );
not ( n255801 , n255798 );
nand ( n255802 , n255801 , n247287 );
nand ( n255803 , n255800 , n255802 );
and ( n255804 , n255791 , n255803 );
not ( n255805 , n255791 );
not ( n255806 , n255803 );
and ( n255807 , n255805 , n255806 );
nor ( n255808 , n255804 , n255807 );
not ( n255809 , n255808 );
not ( n255810 , n255809 );
and ( n255811 , n255768 , n255810 );
not ( n255812 , n255768 );
not ( n255813 , n255808 );
not ( n255814 , n255813 );
not ( n255815 , n255814 );
and ( n255816 , n255812 , n255815 );
nor ( n255817 , n255811 , n255816 );
nor ( n255818 , n255817 , n252258 );
not ( n255819 , n242030 );
not ( n255820 , n246389 );
or ( n255821 , n255819 , n255820 );
buf ( n255822 , n246384 );
or ( n255823 , n255822 , n242030 );
nand ( n255824 , n255821 , n255823 );
and ( n255825 , n255824 , n246441 );
not ( n255826 , n255824 );
and ( n255827 , n255826 , n246449 );
nor ( n255828 , n255825 , n255827 );
not ( n255829 , n249673 );
not ( n255830 , n248385 );
not ( n255831 , n255830 );
or ( n255832 , n255829 , n255831 );
not ( n255833 , n249673 );
nand ( n255834 , n255833 , n248385 );
nand ( n255835 , n255832 , n255834 );
not ( n255836 , n243256 );
not ( n255837 , n229175 );
or ( n255838 , n255836 , n255837 );
or ( n255839 , n229175 , n243256 );
nand ( n255840 , n255838 , n255839 );
not ( n255841 , n255840 );
not ( n255842 , n51460 );
nand ( n255843 , n255842 , n36116 );
not ( n255844 , n255843 );
not ( n255845 , n229218 );
and ( n255846 , n255844 , n255845 );
and ( n255847 , n255843 , n229218 );
nor ( n255848 , n255846 , n255847 );
not ( n255849 , n255848 );
or ( n255850 , n255841 , n255849 );
or ( n255851 , n255848 , n255840 );
nand ( n255852 , n255850 , n255851 );
not ( n255853 , n255852 );
not ( n255854 , n239614 );
not ( n255855 , n51482 );
nand ( n255856 , n255855 , n36194 );
not ( n255857 , n255856 );
or ( n255858 , n255854 , n255857 );
not ( n255859 , n51482 );
nand ( n255860 , n255859 , n36194 );
or ( n255861 , n255860 , n239614 );
nand ( n255862 , n255858 , n255861 );
not ( n255863 , n255862 );
not ( n255864 , n36354 );
nand ( n255865 , n255864 , n51510 );
not ( n255866 , n255865 );
not ( n255867 , n239624 );
and ( n255868 , n255866 , n255867 );
and ( n255869 , n255865 , n239624 );
nor ( n255870 , n255868 , n255869 );
not ( n255871 , n255870 );
and ( n255872 , n255863 , n255871 );
and ( n255873 , n255862 , n255870 );
nor ( n255874 , n255872 , n255873 );
not ( n255875 , n255874 );
and ( n255876 , n255853 , n255875 );
and ( n255877 , n255874 , n255852 );
nor ( n255878 , n255876 , n255877 );
not ( n255879 , n255878 );
not ( n255880 , n255879 );
not ( n255881 , n255880 );
and ( n255882 , n255835 , n255881 );
not ( n255883 , n255835 );
buf ( n255884 , n255878 );
buf ( n255885 , n255884 );
and ( n255886 , n255883 , n255885 );
nor ( n255887 , n255882 , n255886 );
not ( n255888 , n255887 );
nor ( n255889 , n255828 , n255888 );
nand ( n255890 , n255818 , n255889 );
not ( n255891 , n255887 );
not ( n255892 , n255817 );
not ( n255893 , n255892 );
or ( n255894 , n255891 , n255893 );
not ( n255895 , n255828 );
buf ( n255896 , n238635 );
nor ( n255897 , n255895 , n255896 );
nand ( n255898 , n255894 , n255897 );
nand ( n255899 , n255116 , n41001 );
nand ( n255900 , n255890 , n255898 , n255899 );
buf ( n255901 , n255900 );
not ( n255902 , n231622 );
not ( n255903 , n238408 );
or ( n255904 , n255902 , n255903 );
or ( n255905 , n238408 , n231622 );
nand ( n255906 , n255904 , n255905 );
not ( n255907 , n255906 );
not ( n255908 , n251451 );
and ( n255909 , n255907 , n255908 );
and ( n255910 , n255906 , n251451 );
nor ( n255911 , n255909 , n255910 );
nand ( n255912 , n255911 , n241459 );
nor ( n255913 , n47156 , n245979 );
not ( n255914 , n255913 );
nand ( n255915 , n47156 , n245979 );
nand ( n255916 , n255914 , n255915 );
not ( n255917 , n254462 );
and ( n255918 , n255916 , n255917 );
not ( n255919 , n255916 );
and ( n255920 , n255919 , n254462 );
nor ( n255921 , n255918 , n255920 );
not ( n255922 , n255921 );
not ( n255923 , n251721 );
not ( n255924 , n239973 );
not ( n255925 , n255924 );
buf ( n255926 , n56039 );
not ( n255927 , n255926 );
or ( n255928 , n255925 , n255927 );
or ( n255929 , n56041 , n255924 );
nand ( n255930 , n255928 , n255929 );
not ( n255931 , n255930 );
or ( n255932 , n255923 , n255931 );
or ( n255933 , n255930 , n251730 );
nand ( n255934 , n255932 , n255933 );
not ( n255935 , n255934 );
nand ( n255936 , n255922 , n255935 );
or ( n255937 , n255912 , n255936 );
not ( n255938 , n255922 );
not ( n255939 , n255911 );
or ( n255940 , n255938 , n255939 );
nor ( n255941 , n255935 , n40465 );
nand ( n255942 , n255940 , n255941 );
nand ( n255943 , n31577 , n34679 );
nand ( n255944 , n255937 , n255942 , n255943 );
buf ( n255945 , n255944 );
not ( n255946 , n204638 );
not ( n255947 , n234453 );
or ( n255948 , n255946 , n255947 );
not ( n255949 , n248694 );
nand ( n255950 , n255949 , n248765 );
not ( n255951 , n236427 );
not ( n255952 , n32472 );
or ( n255953 , n255951 , n255952 );
not ( n255954 , n236427 );
nand ( n255955 , n255954 , n242585 );
nand ( n255956 , n255953 , n255955 );
not ( n255957 , n255956 );
not ( n255958 , n33247 );
and ( n255959 , n255957 , n255958 );
and ( n255960 , n255956 , n33247 );
nor ( n255961 , n255959 , n255960 );
not ( n255962 , n255961 );
and ( n255963 , n255950 , n255962 );
not ( n255964 , n255950 );
and ( n255965 , n255964 , n255961 );
nor ( n255966 , n255963 , n255965 );
not ( n255967 , n230207 );
or ( n255968 , n255966 , n255967 );
nand ( n255969 , n255948 , n255968 );
buf ( n255970 , n255969 );
or ( n255971 , n226819 , n235905 );
not ( n255972 , RI19aaeea8_2462);
or ( n255973 , n25335 , n255972 );
nand ( n255974 , n255971 , n255973 );
buf ( n255975 , n255974 );
nand ( n255976 , n229128 , RI1754a5b8_71);
and ( n255977 , n255976 , n229127 );
not ( n255978 , RI1754bcb0_22);
or ( n255979 , n255977 , n255978 );
nand ( n255980 , n244606 , n204337 );
nand ( n255981 , n255979 , n255980 );
buf ( n255982 , n255981 );
buf ( n255983 , n31507 );
not ( n255984 , n247126 );
not ( n255985 , n240112 );
and ( n255986 , n247617 , n247640 );
not ( n255987 , n247617 );
and ( n255988 , n255987 , n247639 );
nor ( n255989 , n255986 , n255988 );
not ( n255990 , n255989 );
or ( n255991 , n255985 , n255990 );
not ( n255992 , n255989 );
nand ( n255993 , n255992 , n240109 );
nand ( n255994 , n255991 , n255993 );
not ( n255995 , n255994 );
not ( n255996 , n255995 );
or ( n255997 , n255984 , n255996 );
buf ( n255998 , n247119 );
nand ( n255999 , n255998 , n255994 );
nand ( n256000 , n255997 , n255999 );
not ( n256001 , n256000 );
not ( n256002 , n39043 );
not ( n256003 , n251298 );
or ( n256004 , n256002 , n256003 );
not ( n256005 , n39043 );
nand ( n256006 , n256005 , n251313 );
nand ( n256007 , n256004 , n256006 );
buf ( n256008 , n246826 );
and ( n256009 , n256007 , n256008 );
not ( n256010 , n256007 );
not ( n256011 , n246835 );
not ( n256012 , n256011 );
and ( n256013 , n256010 , n256012 );
nor ( n256014 , n256009 , n256013 );
not ( n256015 , n256014 );
or ( n256016 , n256001 , n256015 );
not ( n256017 , n234143 );
not ( n256018 , n251627 );
or ( n256019 , n256017 , n256018 );
or ( n256020 , n251627 , n234143 );
nand ( n256021 , n256019 , n256020 );
not ( n256022 , n256021 );
not ( n256023 , n251573 );
and ( n256024 , n256022 , n256023 );
and ( n256025 , n256021 , n251573 );
nor ( n256026 , n256024 , n256025 );
nor ( n256027 , n256026 , n226003 );
nand ( n256028 , n256016 , n256027 );
not ( n256029 , n256000 );
nor ( n256030 , n256029 , n247212 );
nand ( n256031 , n256030 , n256026 , n256014 );
nand ( n256032 , n234024 , n204381 );
nand ( n256033 , n256028 , n256031 , n256032 );
buf ( n256034 , n256033 );
buf ( n256035 , n204972 );
not ( n256036 , n54875 );
not ( n256037 , n237936 );
or ( n256038 , n256036 , n256037 );
not ( n256039 , n54875 );
nand ( n256040 , n256039 , n237944 );
nand ( n256041 , n256038 , n256040 );
not ( n256042 , n237444 );
and ( n256043 , n256041 , n256042 );
not ( n256044 , n256041 );
and ( n256045 , n256044 , n237948 );
nor ( n256046 , n256043 , n256045 );
not ( n256047 , n256046 );
nand ( n256048 , n234190 , n256047 );
or ( n256049 , n256048 , n234112 );
nor ( n256050 , n234109 , n238900 );
nand ( n256051 , n256050 , n256048 );
nand ( n256052 , n247744 , n42948 );
nand ( n256053 , n256049 , n256051 , n256052 );
buf ( n256054 , n256053 );
not ( n256055 , RI19a23678_2793);
or ( n256056 , n25328 , n256055 );
not ( n256057 , RI19a85c10_2754);
or ( n256058 , n25336 , n256057 );
nand ( n256059 , n256056 , n256058 );
buf ( n256060 , n256059 );
not ( n256061 , n236825 );
nand ( n256062 , n256061 , n226010 );
not ( n256063 , n241580 );
not ( n256064 , n243363 );
or ( n256065 , n256063 , n256064 );
not ( n256066 , n241580 );
nand ( n256067 , n256066 , n243372 );
nand ( n256068 , n256065 , n256067 );
not ( n256069 , n246693 );
and ( n256070 , n256068 , n256069 );
not ( n256071 , n256068 );
and ( n256072 , n256071 , n246694 );
nor ( n256073 , n256070 , n256072 );
nand ( n256074 , n237352 , n256073 );
or ( n256075 , n256062 , n256074 );
not ( n256076 , n237352 );
not ( n256077 , n256061 );
or ( n256078 , n256076 , n256077 );
nor ( n256079 , n256073 , n47173 );
nand ( n256080 , n256078 , n256079 );
nand ( n256081 , n244987 , n29365 );
nand ( n256082 , n256075 , n256080 , n256081 );
buf ( n256083 , n256082 );
buf ( n256084 , n43628 );
not ( n256085 , RI19a9d658_2588);
or ( n256086 , n25328 , n256085 );
not ( n256087 , RI19a932c0_2660);
or ( n256088 , n25336 , n256087 );
nand ( n256089 , n256086 , n256088 );
buf ( n256090 , n256089 );
buf ( n256091 , n204496 );
not ( n256092 , n247646 );
not ( n256093 , n238057 );
not ( n256094 , n247689 );
not ( n256095 , n256094 );
or ( n256096 , n256093 , n256095 );
nand ( n256097 , n247689 , n238056 );
nand ( n256098 , n256096 , n256097 );
not ( n256099 , n256098 );
or ( n256100 , n256092 , n256099 );
or ( n256101 , n256098 , n247646 );
nand ( n256102 , n256100 , n256101 );
nor ( n256103 , n38636 , n256102 );
not ( n256104 , n256103 );
not ( n256105 , n232914 );
or ( n256106 , n256104 , n256105 );
nand ( n256107 , n252711 , n208545 );
nand ( n256108 , n256106 , n256107 );
not ( n256109 , n256108 );
not ( n256110 , n55148 );
nand ( n256111 , n256110 , n38636 );
not ( n256112 , n38639 );
nand ( n256113 , n256112 , n256102 );
nand ( n256114 , n256109 , n256111 , n256113 );
buf ( n256115 , n256114 );
not ( n256116 , n50577 );
not ( n256117 , n209312 );
or ( n256118 , n256116 , n256117 );
or ( n256119 , n209312 , n50577 );
nand ( n256120 , n256118 , n256119 );
and ( n256121 , n256120 , n35805 );
not ( n256122 , n256120 );
and ( n256123 , n256122 , n35813 );
nor ( n256124 , n256121 , n256123 );
nor ( n256125 , n256124 , n226955 );
not ( n256126 , n255743 );
and ( n256127 , n241153 , n241174 );
not ( n256128 , n241153 );
and ( n256129 , n256128 , n241177 );
nor ( n256130 , n256127 , n256129 );
not ( n256131 , n256130 );
not ( n256132 , n256131 );
or ( n256133 , n256126 , n256132 );
not ( n256134 , n255743 );
nand ( n256135 , n256134 , n256130 );
nand ( n256136 , n256133 , n256135 );
and ( n256137 , n256136 , n249549 );
not ( n256138 , n256136 );
and ( n256139 , n256138 , n249546 );
nor ( n256140 , n256137 , n256139 );
not ( n256141 , n256140 );
buf ( n256142 , n54944 );
not ( n256143 , n256142 );
not ( n256144 , n237444 );
or ( n256145 , n256143 , n256144 );
or ( n256146 , n237444 , n256142 );
nand ( n256147 , n256145 , n256146 );
not ( n256148 , n256147 );
not ( n256149 , n256148 );
not ( n256150 , n237590 );
or ( n256151 , n256149 , n256150 );
not ( n256152 , n237590 );
buf ( n256153 , n256152 );
nand ( n256154 , n256153 , n256147 );
nand ( n256155 , n256151 , n256154 );
nor ( n256156 , n256141 , n256155 );
nand ( n256157 , n256125 , n256156 );
not ( n256158 , n256155 );
not ( n256159 , n256158 );
not ( n256160 , n256124 );
not ( n256161 , n256160 );
or ( n256162 , n256159 , n256161 );
nor ( n256163 , n256140 , n238635 );
nand ( n256164 , n256162 , n256163 );
nand ( n256165 , n255116 , n39390 );
nand ( n256166 , n256157 , n256164 , n256165 );
buf ( n256167 , n256166 );
not ( n256168 , n215255 );
not ( n256169 , n51381 );
or ( n256170 , n256168 , n256169 );
not ( n256171 , n242231 );
not ( n256172 , n249298 );
or ( n256173 , n256171 , n256172 );
not ( n256174 , n242231 );
nand ( n256175 , n256174 , n53140 );
nand ( n256176 , n256173 , n256175 );
and ( n256177 , n256176 , n249366 );
not ( n256178 , n256176 );
and ( n256179 , n256178 , n249363 );
nor ( n256180 , n256177 , n256179 );
not ( n256181 , n242920 );
not ( n256182 , n245929 );
or ( n256183 , n256181 , n256182 );
not ( n256184 , n242920 );
nand ( n256185 , n256184 , n245918 );
nand ( n256186 , n256183 , n256185 );
and ( n256187 , n249835 , n249818 );
not ( n256188 , n249835 );
and ( n256189 , n256188 , n249839 );
nor ( n256190 , n256187 , n256189 );
not ( n256191 , n256190 );
buf ( n256192 , n256191 );
and ( n256193 , n256186 , n256192 );
not ( n256194 , n256186 );
not ( n256195 , n256192 );
and ( n256196 , n256194 , n256195 );
nor ( n256197 , n256193 , n256196 );
not ( n256198 , n256197 );
nand ( n256199 , n256180 , n256198 );
not ( n256200 , n51589 );
not ( n256201 , n241695 );
or ( n256202 , n256200 , n256201 );
or ( n256203 , n241695 , n51589 );
nand ( n256204 , n256202 , n256203 );
and ( n256205 , n256204 , n46067 );
not ( n256206 , n256204 );
and ( n256207 , n256206 , n223836 );
nor ( n256208 , n256205 , n256207 );
not ( n256209 , n256208 );
and ( n256210 , n256199 , n256209 );
not ( n256211 , n256199 );
and ( n256212 , n256211 , n256208 );
nor ( n256213 , n256210 , n256212 );
buf ( n256214 , n226003 );
or ( n256215 , n256213 , n256214 );
nand ( n256216 , n256170 , n256215 );
buf ( n256217 , n256216 );
buf ( n256218 , n30929 );
buf ( n256219 , n38317 );
not ( n256220 , n240213 );
not ( n256221 , n252051 );
or ( n256222 , n256220 , n256221 );
or ( n256223 , n252051 , n240213 );
nand ( n256224 , n256222 , n256223 );
and ( n256225 , n256224 , n252644 );
not ( n256226 , n256224 );
buf ( n256227 , n252649 );
and ( n256228 , n256226 , n256227 );
nor ( n256229 , n256225 , n256228 );
not ( n256230 , n256229 );
nand ( n256231 , n256230 , n241459 );
not ( n256232 , n237415 );
not ( n256233 , n247813 );
or ( n256234 , n256232 , n256233 );
not ( n256235 , n237415 );
nand ( n256236 , n256235 , n247822 );
nand ( n256237 , n256234 , n256236 );
and ( n256238 , n256237 , n247872 );
not ( n256239 , n256237 );
and ( n256240 , n256239 , n247873 );
nor ( n256241 , n256238 , n256240 );
not ( n256242 , n250077 );
not ( n256243 , n236056 );
or ( n256244 , n256242 , n256243 );
not ( n256245 , n250077 );
nand ( n256246 , n256245 , n236055 );
nand ( n256247 , n256244 , n256246 );
and ( n256248 , n256247 , n236168 );
not ( n256249 , n256247 );
and ( n256250 , n256249 , n236172 );
nor ( n256251 , n256248 , n256250 );
not ( n256252 , n256251 );
nand ( n256253 , n256241 , n256252 );
or ( n256254 , n256231 , n256253 );
not ( n256255 , n256252 );
not ( n256256 , n256230 );
or ( n256257 , n256255 , n256256 );
nor ( n256258 , n256241 , n253904 );
nand ( n256259 , n256257 , n256258 );
nand ( n256260 , n31577 , n204570 );
nand ( n256261 , n256254 , n256259 , n256260 );
buf ( n256262 , n256261 );
nand ( n256263 , n253734 , n253393 );
not ( n256264 , n42872 );
not ( n256265 , n237700 );
or ( n256266 , n256264 , n256265 );
or ( n256267 , n237700 , n42872 );
nand ( n256268 , n256266 , n256267 );
and ( n256269 , n256268 , n243226 );
not ( n256270 , n256268 );
and ( n256271 , n256270 , n243230 );
nor ( n256272 , n256269 , n256271 );
not ( n256273 , n248865 );
not ( n256274 , n237340 );
or ( n256275 , n256273 , n256274 );
not ( n256276 , n248865 );
nand ( n256277 , n256276 , n237350 );
nand ( n256278 , n256275 , n256277 );
buf ( n256279 , n245201 );
not ( n256280 , n256279 );
and ( n256281 , n256278 , n256280 );
not ( n256282 , n256278 );
and ( n256283 , n256282 , n256279 );
nor ( n256284 , n256281 , n256283 );
nand ( n256285 , n256272 , n256284 );
or ( n256286 , n256263 , n256285 );
not ( n256287 , n256272 );
not ( n256288 , n253734 );
or ( n256289 , n256287 , n256288 );
nor ( n256290 , n256284 , n251361 );
nand ( n256291 , n256289 , n256290 );
buf ( n256292 , n35431 );
nand ( n256293 , n256292 , n37326 );
nand ( n256294 , n256286 , n256291 , n256293 );
buf ( n256295 , n256294 );
not ( n256296 , RI19ac7700_2274);
or ( n256297 , n25328 , n256296 );
not ( n256298 , RI19abe808_2345);
or ( n256299 , n25335 , n256298 );
nand ( n256300 , n256297 , n256299 );
buf ( n256301 , n256300 );
not ( n256302 , RI19abef88_2341);
or ( n256303 , n25328 , n256302 );
not ( n256304 , RI19ab5a00_2411);
or ( n256305 , n25335 , n256304 );
nand ( n256306 , n256303 , n256305 );
buf ( n256307 , n256306 );
not ( n256308 , n251226 );
not ( n256309 , n256308 );
not ( n256310 , n251238 );
or ( n256311 , n256309 , n256310 );
nand ( n256312 , n256311 , n241459 );
not ( n256313 , n52166 );
not ( n256314 , n236267 );
or ( n256315 , n256313 , n256314 );
not ( n256316 , n52166 );
nand ( n256317 , n256316 , n245210 );
nand ( n256318 , n256315 , n256317 );
and ( n256319 , n256318 , n251181 );
not ( n256320 , n256318 );
and ( n256321 , n256320 , n44539 );
nor ( n256322 , n256319 , n256321 );
or ( n256323 , n256312 , n256322 );
nor ( n256324 , n251226 , n238635 );
nand ( n256325 , n256324 , n251238 , n256322 );
nand ( n256326 , n245701 , n30661 );
nand ( n256327 , n256323 , n256325 , n256326 );
buf ( n256328 , n256327 );
or ( n256329 , n25328 , n55749 );
or ( n256330 , n226822 , n256296 );
nand ( n256331 , n256329 , n256330 );
buf ( n256332 , n256331 );
not ( n256333 , n30724 );
not ( n256334 , n237714 );
or ( n256335 , n256333 , n256334 );
not ( n256336 , n242941 );
not ( n256337 , n245929 );
or ( n256338 , n256336 , n256337 );
not ( n256339 , n242941 );
nand ( n256340 , n256339 , n245918 );
nand ( n256341 , n256338 , n256340 );
and ( n256342 , n256341 , n256192 );
not ( n256343 , n256341 );
and ( n256344 , n256343 , n256195 );
nor ( n256345 , n256342 , n256344 );
not ( n256346 , n245974 );
not ( n256347 , n224924 );
or ( n256348 , n256346 , n256347 );
not ( n256349 , n245974 );
nand ( n256350 , n256349 , n47156 );
nand ( n256351 , n256348 , n256350 );
and ( n256352 , n256351 , n245677 );
not ( n256353 , n256351 );
and ( n256354 , n256353 , n245680 );
nor ( n256355 , n256352 , n256354 );
nand ( n256356 , n256345 , n256355 );
not ( n256357 , n256356 );
not ( n256358 , n244290 );
not ( n256359 , n29962 );
or ( n256360 , n256358 , n256359 );
not ( n256361 , n244290 );
not ( n256362 , n29961 );
nand ( n256363 , n256361 , n256362 );
nand ( n256364 , n256360 , n256363 );
not ( n256365 , n256364 );
buf ( n256366 , n235580 );
not ( n256367 , n256366 );
and ( n256368 , n256365 , n256367 );
and ( n256369 , n256364 , n256366 );
nor ( n256370 , n256368 , n256369 );
not ( n256371 , n256370 );
not ( n256372 , n256371 );
and ( n256373 , n256357 , n256372 );
and ( n256374 , n256371 , n256356 );
nor ( n256375 , n256373 , n256374 );
not ( n256376 , n205649 );
or ( n256377 , n256375 , n256376 );
nand ( n256378 , n256335 , n256377 );
buf ( n256379 , n256378 );
not ( n256380 , RI19aa0f10_2561);
or ( n256381 , n25328 , n256380 );
not ( n256382 , RI19a97460_2631);
or ( n256383 , n25335 , n256382 );
nand ( n256384 , n256381 , n256383 );
buf ( n256385 , n256384 );
nor ( n256386 , n252257 , n241065 );
not ( n256387 , n256386 );
not ( n256388 , n239894 );
not ( n256389 , n247569 );
or ( n256390 , n256388 , n256389 );
not ( n256391 , n239894 );
nand ( n256392 , n256391 , n230199 );
nand ( n256393 , n256390 , n256392 );
and ( n256394 , n256393 , n242696 );
not ( n256395 , n256393 );
and ( n256396 , n256395 , n247575 );
nor ( n256397 , n256394 , n256396 );
nand ( n256398 , n252245 , n256397 );
or ( n256399 , n256387 , n256398 );
not ( n256400 , n252245 );
not ( n256401 , n252256 );
or ( n256402 , n256400 , n256401 );
nor ( n256403 , n256397 , n54208 );
nand ( n256404 , n256402 , n256403 );
nand ( n256405 , n50615 , n205361 );
nand ( n256406 , n256399 , n256404 , n256405 );
buf ( n256407 , n256406 );
not ( n256408 , n56046 );
nand ( n256409 , n234441 , n234339 , n256408 );
not ( n256410 , n234444 );
not ( n256411 , n234339 );
or ( n256412 , n256410 , n256411 );
not ( n256413 , n241373 );
nor ( n256414 , n256408 , n256413 );
nand ( n256415 , n256412 , n256414 );
nand ( n256416 , n35431 , n37969 );
nand ( n256417 , n256409 , n256415 , n256416 );
buf ( n256418 , n256417 );
not ( n256419 , RI19acbc60_2241);
or ( n256420 , n25328 , n256419 );
not ( n256421 , RI19ac2cf0_2308);
or ( n256422 , n25336 , n256421 );
nand ( n256423 , n256420 , n256422 );
buf ( n256424 , n256423 );
not ( n256425 , n38303 );
not ( n256426 , n256425 );
not ( n256427 , n234513 );
or ( n256428 , n256426 , n256427 );
nand ( n256429 , n234521 , n38303 );
nand ( n256430 , n256428 , n256429 );
not ( n256431 , n256430 );
not ( n256432 , n45507 );
and ( n256433 , n256431 , n256432 );
and ( n256434 , n256430 , n243427 );
nor ( n256435 , n256433 , n256434 );
not ( n256436 , n256435 );
nor ( n256437 , n256436 , n50944 );
not ( n256438 , n230199 );
not ( n256439 , n256438 );
buf ( n256440 , n239834 );
not ( n256441 , n256440 );
not ( n256442 , n256441 );
not ( n256443 , n46708 );
or ( n256444 , n256442 , n256443 );
nand ( n256445 , n46716 , n256440 );
nand ( n256446 , n256444 , n256445 );
not ( n256447 , n256446 );
or ( n256448 , n256439 , n256447 );
or ( n256449 , n256446 , n230201 );
nand ( n256450 , n256448 , n256449 );
not ( n256451 , n256450 );
not ( n256452 , n48865 );
not ( n256453 , n44315 );
or ( n256454 , n256452 , n256453 );
not ( n256455 , n48865 );
nand ( n256456 , n256455 , n44324 );
nand ( n256457 , n256454 , n256456 );
and ( n256458 , n256457 , n254603 );
not ( n256459 , n256457 );
buf ( n256460 , n254602 );
and ( n256461 , n256459 , n256460 );
nor ( n256462 , n256458 , n256461 );
not ( n256463 , n256462 );
nand ( n256464 , n256437 , n256451 , n256463 );
nand ( n256465 , n256463 , n256435 );
nand ( n256466 , n256465 , n256450 , n241459 );
nand ( n256467 , n254798 , n26248 );
nand ( n256468 , n256464 , n256466 , n256467 );
buf ( n256469 , n256468 );
not ( n256470 , n40755 );
not ( n256471 , n251450 );
or ( n256472 , n256470 , n256471 );
nand ( n256473 , n251443 , n40754 );
nand ( n256474 , n256472 , n256473 );
not ( n256475 , n256474 );
not ( n256476 , n253106 );
and ( n256477 , n256475 , n256476 );
and ( n256478 , n256474 , n253106 );
nor ( n256479 , n256477 , n256478 );
not ( n256480 , n256479 );
not ( n256481 , n205649 );
nor ( n256482 , n256480 , n256481 );
not ( n256483 , n253253 );
not ( n256484 , n240684 );
or ( n256485 , n256483 , n256484 );
not ( n256486 , n253253 );
nand ( n256487 , n256486 , n240676 );
nand ( n256488 , n256485 , n256487 );
and ( n256489 , n256488 , n240811 );
not ( n256490 , n256488 );
and ( n256491 , n256490 , n240801 );
nor ( n256492 , n256489 , n256491 );
not ( n256493 , n50867 );
not ( n256494 , n255514 );
not ( n256495 , n256494 );
or ( n256496 , n256493 , n256495 );
not ( n256497 , n255514 );
or ( n256498 , n256497 , n50867 );
nand ( n256499 , n256496 , n256498 );
not ( n256500 , n250900 );
and ( n256501 , n256499 , n256500 );
not ( n256502 , n256499 );
and ( n256503 , n256502 , n251975 );
nor ( n256504 , n256501 , n256503 );
nor ( n256505 , n256492 , n256504 );
nand ( n256506 , n256482 , n256505 );
not ( n256507 , n256504 );
not ( n256508 , n256507 );
not ( n256509 , n256479 );
or ( n256510 , n256508 , n256509 );
not ( n256511 , n256492 );
nor ( n256512 , n256511 , n31572 );
nand ( n256513 , n256510 , n256512 );
nand ( n256514 , n246460 , n32246 );
nand ( n256515 , n256506 , n256513 , n256514 );
buf ( n256516 , n256515 );
not ( n256517 , n40559 );
not ( n256518 , n237361 );
or ( n256519 , n256517 , n256518 );
not ( n256520 , n245757 );
not ( n256521 , n52756 );
or ( n256522 , n256520 , n256521 );
not ( n256523 , n245757 );
nand ( n256524 , n256523 , n245264 );
nand ( n256525 , n256522 , n256524 );
and ( n256526 , n256525 , n251156 );
not ( n256527 , n256525 );
and ( n256528 , n256527 , n252733 );
nor ( n256529 , n256526 , n256528 );
not ( n256530 , n256529 );
not ( n256531 , n244761 );
not ( n256532 , n241877 );
or ( n256533 , n256531 , n256532 );
not ( n256534 , n244761 );
nand ( n256535 , n256534 , n241884 );
nand ( n256536 , n256533 , n256535 );
and ( n256537 , n256536 , n254238 );
not ( n256538 , n256536 );
and ( n256539 , n256538 , n254235 );
nor ( n256540 , n256537 , n256539 );
not ( n256541 , n256540 );
nand ( n256542 , n256530 , n256541 );
not ( n256543 , n230073 );
not ( n256544 , n256543 );
not ( n256545 , n248055 );
or ( n256546 , n256544 , n256545 );
not ( n256547 , n248054 );
or ( n256548 , n256547 , n256543 );
nand ( n256549 , n256546 , n256548 );
and ( n256550 , n256549 , n248063 );
not ( n256551 , n256549 );
and ( n256552 , n256551 , n248067 );
nor ( n256553 , n256550 , n256552 );
not ( n256554 , n256553 );
and ( n256555 , n256542 , n256554 );
not ( n256556 , n256542 );
and ( n256557 , n256556 , n256553 );
nor ( n256558 , n256555 , n256557 );
or ( n256559 , n256558 , n244217 );
nand ( n256560 , n256519 , n256559 );
buf ( n256561 , n256560 );
not ( n256562 , RI19a841d0_2765);
or ( n256563 , n25328 , n256562 );
not ( n256564 , RI19ac90c8_2262);
or ( n256565 , n25335 , n256564 );
nand ( n256566 , n256563 , n256565 );
buf ( n256567 , n256566 );
not ( n256568 , RI19ab01e0_2453);
or ( n256569 , n25328 , n256568 );
not ( n256570 , RI19aa5fb0_2523);
or ( n256571 , n25336 , n256570 );
nand ( n256572 , n256569 , n256571 );
buf ( n256573 , n256572 );
not ( n256574 , RI19a93d88_2655);
or ( n256575 , n25328 , n256574 );
not ( n256576 , RI19a89bd0_2726);
or ( n256577 , n25335 , n256576 );
nand ( n256578 , n256575 , n256577 );
buf ( n256579 , n256578 );
xor ( n256580 , n238609 , n256131 );
xor ( n256581 , n256580 , n244472 );
not ( n256582 , n256581 );
nand ( n256583 , n256582 , n256252 );
not ( n256584 , n250909 );
nand ( n256585 , n256229 , n256584 );
or ( n256586 , n256583 , n256585 );
not ( n256587 , n256229 );
not ( n256588 , n256581 );
not ( n256589 , n256588 );
or ( n256590 , n256587 , n256589 );
nor ( n256591 , n256252 , n39763 );
nand ( n256592 , n256590 , n256591 );
nand ( n256593 , n247585 , n34906 );
nand ( n256594 , n256586 , n256592 , n256593 );
buf ( n256595 , n256594 );
not ( n256596 , n245125 );
not ( n256597 , n40914 );
or ( n256598 , n256596 , n256597 );
or ( n256599 , n40918 , n245125 );
nand ( n256600 , n256598 , n256599 );
not ( n256601 , n256600 );
not ( n256602 , n41217 );
and ( n256603 , n256601 , n256602 );
and ( n256604 , n256600 , n41217 );
nor ( n256605 , n256603 , n256604 );
not ( n256606 , n256605 );
nor ( n256607 , n256606 , n251190 );
not ( n256608 , n45365 );
not ( n256609 , n256608 );
not ( n256610 , n252843 );
or ( n256611 , n256609 , n256610 );
or ( n256612 , n248154 , n256608 );
nand ( n256613 , n256611 , n256612 );
and ( n256614 , n256613 , n248211 );
not ( n256615 , n256613 );
and ( n256616 , n256615 , n248220 );
nor ( n256617 , n256614 , n256616 );
not ( n256618 , n256617 );
not ( n256619 , n247451 );
not ( n256620 , n243510 );
or ( n256621 , n256619 , n256620 );
not ( n256622 , n247451 );
nand ( n256623 , n256622 , n243503 );
nand ( n256624 , n256621 , n256623 );
and ( n256625 , n256624 , n248478 );
not ( n256626 , n256624 );
and ( n256627 , n256626 , n248481 );
nor ( n256628 , n256625 , n256627 );
not ( n256629 , n256628 );
nand ( n256630 , n256607 , n256618 , n256629 );
not ( n256631 , n256605 );
not ( n256632 , n256617 );
not ( n256633 , n256632 );
or ( n256634 , n256631 , n256633 );
nor ( n256635 , n256629 , n239237 );
nand ( n256636 , n256634 , n256635 );
nand ( n256637 , n246460 , n241526 );
nand ( n256638 , n256630 , n256636 , n256637 );
buf ( n256639 , n256638 );
buf ( n256640 , n238391 );
not ( n256641 , n256640 );
not ( n256642 , n254337 );
or ( n256643 , n256641 , n256642 );
or ( n256644 , n254337 , n256640 );
nand ( n256645 , n256643 , n256644 );
buf ( n256646 , n252132 );
and ( n256647 , n256645 , n256646 );
not ( n256648 , n256645 );
buf ( n256649 , n252139 );
and ( n256650 , n256648 , n256649 );
nor ( n256651 , n256647 , n256650 );
not ( n256652 , n256651 );
nand ( n256653 , n256652 , n252873 );
not ( n256654 , n250328 );
not ( n256655 , n237135 );
or ( n256656 , n256654 , n256655 );
not ( n256657 , n250328 );
nand ( n256658 , n256657 , n237148 );
nand ( n256659 , n256656 , n256658 );
and ( n256660 , n256659 , n237342 );
not ( n256661 , n256659 );
and ( n256662 , n256661 , n250412 );
nor ( n256663 , n256660 , n256662 );
not ( n256664 , n256663 );
not ( n256665 , n255690 );
nand ( n256666 , n256664 , n256665 );
or ( n256667 , n256653 , n256666 );
not ( n256668 , n256664 );
not ( n256669 , n256652 );
or ( n256670 , n256668 , n256669 );
nor ( n256671 , n256665 , n234818 );
nand ( n256672 , n256670 , n256671 );
buf ( n256673 , n35431 );
nand ( n256674 , n256673 , n37365 );
nand ( n256675 , n256667 , n256672 , n256674 );
buf ( n256676 , n256675 );
not ( n256677 , RI19aa4a98_2532);
or ( n256678 , n25328 , n256677 );
not ( n256679 , RI19a9b1c8_2604);
or ( n256680 , n226822 , n256679 );
nand ( n256681 , n256678 , n256680 );
buf ( n256682 , n256681 );
not ( n256683 , n250453 );
not ( n256684 , n234691 );
or ( n256685 , n256683 , n256684 );
or ( n256686 , n253386 , n250453 );
nand ( n256687 , n256685 , n256686 );
and ( n256688 , n256687 , n234804 );
not ( n256689 , n256687 );
and ( n256690 , n256689 , n234811 );
nor ( n256691 , n256688 , n256690 );
nand ( n256692 , n256691 , n40466 );
not ( n256693 , n240132 );
not ( n256694 , n256693 );
not ( n256695 , n247644 );
not ( n256696 , n256695 );
or ( n256697 , n256694 , n256696 );
or ( n256698 , n256695 , n256693 );
nand ( n256699 , n256697 , n256698 );
and ( n256700 , n256699 , n255998 );
not ( n256701 , n256699 );
and ( n256702 , n256701 , n247126 );
nor ( n256703 , n256700 , n256702 );
not ( n256704 , n256703 );
not ( n256705 , n28918 );
not ( n256706 , n254866 );
or ( n256707 , n256705 , n256706 );
not ( n256708 , n28918 );
nand ( n256709 , n256708 , n254873 );
nand ( n256710 , n256707 , n256709 );
xnor ( n256711 , n253007 , n252968 );
buf ( n256712 , n256711 );
and ( n256713 , n256710 , n256712 );
not ( n256714 , n256710 );
not ( n256715 , n253009 );
not ( n256716 , n256715 );
and ( n256717 , n256714 , n256716 );
nor ( n256718 , n256713 , n256717 );
nor ( n256719 , n256704 , n256718 );
or ( n256720 , n256692 , n256719 );
not ( n256721 , n39766 );
not ( n256722 , n256721 );
not ( n256723 , n35999 );
and ( n256724 , n256722 , n256723 );
not ( n256725 , n43517 );
nand ( n256726 , n256725 , n256703 );
nor ( n256727 , n256726 , n256718 );
not ( n256728 , n256691 );
and ( n256729 , n256727 , n256728 );
nor ( n256730 , n256724 , n256729 );
nand ( n256731 , n256720 , n256730 );
buf ( n256732 , n256731 );
buf ( n256733 , n246414 );
not ( n256734 , n256733 );
and ( n256735 , n44663 , n44755 );
not ( n256736 , n44663 );
and ( n256737 , n256736 , n44758 );
nor ( n256738 , n256735 , n256737 );
not ( n256739 , n256738 );
not ( n256740 , n256739 );
or ( n256741 , n256734 , n256740 );
not ( n256742 , n44760 );
or ( n256743 , n256742 , n256733 );
nand ( n256744 , n256741 , n256743 );
not ( n256745 , n256744 );
not ( n256746 , n228527 );
and ( n256747 , n256745 , n256746 );
buf ( n256748 , n228527 );
and ( n256749 , n256744 , n256748 );
nor ( n256750 , n256747 , n256749 );
not ( n256751 , n49051 );
nand ( n256752 , n256750 , n256751 );
not ( n256753 , n51216 );
not ( n256754 , n255808 );
or ( n256755 , n256753 , n256754 );
not ( n256756 , n51216 );
not ( n256757 , n255791 );
not ( n256758 , n255803 );
and ( n256759 , n256757 , n256758 );
and ( n256760 , n255791 , n255803 );
nor ( n256761 , n256759 , n256760 );
not ( n256762 , n256761 );
nand ( n256763 , n256756 , n256762 );
nand ( n256764 , n256755 , n256763 );
not ( n256765 , n253673 );
and ( n256766 , n256764 , n256765 );
not ( n256767 , n256764 );
not ( n256768 , n253669 );
and ( n256769 , n256767 , n256768 );
nor ( n256770 , n256766 , n256769 );
not ( n256771 , n256770 );
buf ( n256772 , n252299 );
not ( n256773 , n256772 );
not ( n256774 , n243953 );
or ( n256775 , n256773 , n256774 );
or ( n256776 , n243953 , n256772 );
nand ( n256777 , n256775 , n256776 );
and ( n256778 , n256777 , n250272 );
not ( n256779 , n256777 );
and ( n256780 , n256779 , n250275 );
nor ( n256781 , n256778 , n256780 );
nand ( n256782 , n256771 , n256781 );
or ( n256783 , n256752 , n256782 );
nor ( n256784 , n256750 , n250431 );
nand ( n256785 , n256784 , n256782 );
nand ( n256786 , n231444 , n31622 );
nand ( n256787 , n256783 , n256785 , n256786 );
buf ( n256788 , n256787 );
not ( n256789 , n252926 );
not ( n256790 , n242324 );
not ( n256791 , n39749 );
or ( n256792 , n256790 , n256791 );
or ( n256793 , n217515 , n242324 );
nand ( n256794 , n256792 , n256793 );
not ( n256795 , n256794 );
not ( n256796 , n254730 );
and ( n256797 , n256795 , n256796 );
and ( n256798 , n256794 , n254730 );
nor ( n256799 , n256797 , n256798 );
nand ( n256800 , n256789 , n256799 );
not ( n256801 , n38920 );
not ( n256802 , n251298 );
or ( n256803 , n256801 , n256802 );
not ( n256804 , n38920 );
nand ( n256805 , n256804 , n251313 );
nand ( n256806 , n256803 , n256805 );
and ( n256807 , n256806 , n256012 );
not ( n256808 , n256806 );
and ( n256809 , n256808 , n256008 );
nor ( n256810 , n256807 , n256809 );
not ( n256811 , n40465 );
nand ( n256812 , n256810 , n256811 );
or ( n256813 , n256800 , n256812 );
nand ( n256814 , n256810 , n256799 );
nand ( n256815 , n256814 , n252926 , n254227 );
nand ( n256816 , n31577 , n37552 );
nand ( n256817 , n256813 , n256815 , n256816 );
buf ( n256818 , n256817 );
not ( n256819 , n26118 );
not ( n256820 , n234453 );
or ( n256821 , n256819 , n256820 );
not ( n256822 , n51692 );
not ( n256823 , n256822 );
not ( n256824 , n30287 );
nand ( n256825 , n256824 , n229387 );
not ( n256826 , n256825 );
not ( n256827 , n246930 );
and ( n256828 , n256826 , n256827 );
and ( n256829 , n256825 , n246930 );
nor ( n256830 , n256828 , n256829 );
not ( n256831 , n256830 );
not ( n256832 , n30222 );
nand ( n256833 , n256832 , n249825 );
and ( n256834 , n256833 , n30209 );
not ( n256835 , n256833 );
and ( n256836 , n256835 , n246915 );
nor ( n256837 , n256834 , n256836 );
not ( n256838 , n256837 );
or ( n256839 , n256831 , n256838 );
or ( n256840 , n256837 , n256830 );
nand ( n256841 , n256839 , n256840 );
and ( n256842 , n256841 , n254778 );
not ( n256843 , n256841 );
and ( n256844 , n256843 , n254779 );
nor ( n256845 , n256842 , n256844 );
not ( n256846 , n256845 );
nand ( n256847 , n249811 , n51715 );
and ( n256848 , n256847 , n30895 );
not ( n256849 , n256847 );
and ( n256850 , n256849 , n246906 );
nor ( n256851 , n256848 , n256850 );
not ( n256852 , n256851 );
not ( n256853 , n256852 );
not ( n256854 , n30109 );
or ( n256855 , n256853 , n256854 );
not ( n256856 , n30109 );
nand ( n256857 , n256856 , n256851 );
nand ( n256858 , n256855 , n256857 );
not ( n256859 , n256858 );
and ( n256860 , n256846 , n256859 );
and ( n256861 , n256845 , n256858 );
nor ( n256862 , n256860 , n256861 );
not ( n256863 , n256862 );
or ( n256864 , n256823 , n256863 );
not ( n256865 , n256822 );
not ( n256866 , n256858 );
and ( n256867 , n256845 , n256866 );
not ( n256868 , n256845 );
and ( n256869 , n256868 , n256858 );
nor ( n256870 , n256867 , n256869 );
nand ( n256871 , n256865 , n256870 );
nand ( n256872 , n256864 , n256871 );
and ( n256873 , n50568 , n228351 );
not ( n256874 , n50568 );
and ( n256875 , n256874 , n50589 );
nor ( n256876 , n256873 , n256875 );
not ( n256877 , n256876 );
buf ( n256878 , n256877 );
not ( n256879 , n256878 );
and ( n256880 , n256872 , n256879 );
not ( n256881 , n256872 );
and ( n256882 , n256881 , n256878 );
nor ( n256883 , n256880 , n256882 );
not ( n256884 , n241410 );
not ( n256885 , n47531 );
or ( n256886 , n256884 , n256885 );
not ( n256887 , n241410 );
nand ( n256888 , n256887 , n225301 );
nand ( n256889 , n256886 , n256888 );
and ( n256890 , n256889 , n225536 );
not ( n256891 , n256889 );
buf ( n256892 , n225525 );
and ( n256893 , n256891 , n256892 );
nor ( n256894 , n256890 , n256893 );
nand ( n256895 , n256883 , n256894 );
not ( n256896 , n248117 );
not ( n256897 , n256896 );
not ( n256898 , n255556 );
not ( n256899 , n255584 );
or ( n256900 , n256898 , n256899 );
nand ( n256901 , n256900 , n255588 );
not ( n256902 , n256901 );
or ( n256903 , n256897 , n256902 );
nand ( n256904 , n255593 , n248117 );
nand ( n256905 , n256903 , n256904 );
not ( n256906 , n256905 );
not ( n256907 , n255596 );
and ( n256908 , n256906 , n256907 );
and ( n256909 , n256905 , n255596 );
nor ( n256910 , n256908 , n256909 );
not ( n256911 , n256910 );
and ( n256912 , n256895 , n256911 );
not ( n256913 , n256895 );
and ( n256914 , n256913 , n256910 );
nor ( n256915 , n256912 , n256914 );
or ( n256916 , n256915 , n35816 );
nand ( n256917 , n256821 , n256916 );
buf ( n256918 , n256917 );
buf ( n256919 , n41284 );
buf ( n256920 , n30715 );
buf ( n256921 , n40410 );
not ( n256922 , n42427 );
not ( n256923 , n234305 );
or ( n256924 , n256922 , n256923 );
not ( n256925 , n42427 );
nand ( n256926 , n256925 , n234298 );
nand ( n256927 , n256924 , n256926 );
buf ( n256928 , n248455 );
and ( n256929 , n256927 , n256928 );
not ( n256930 , n256927 );
not ( n256931 , n248446 );
not ( n256932 , n256931 );
and ( n256933 , n256930 , n256932 );
nor ( n256934 , n256929 , n256933 );
not ( n256935 , n256934 );
nand ( n256936 , n54017 , n256935 );
or ( n256937 , n54201 , n256936 );
not ( n256938 , n54199 );
not ( n256939 , n54017 );
or ( n256940 , n256938 , n256939 );
nor ( n256941 , n256935 , n235050 );
nand ( n256942 , n256940 , n256941 );
nand ( n256943 , n252711 , n38328 );
nand ( n256944 , n256937 , n256942 , n256943 );
buf ( n256945 , n256944 );
not ( n256946 , n236136 );
not ( n256947 , n251049 );
not ( n256948 , n251078 );
or ( n256949 , n256947 , n256948 );
nand ( n256950 , n256949 , n251081 );
not ( n256951 , n256950 );
or ( n256952 , n256946 , n256951 );
or ( n256953 , n256950 , n236136 );
nand ( n256954 , n256952 , n256953 );
xnor ( n256955 , n256954 , n251029 );
not ( n256956 , n256955 );
not ( n256957 , n37724 );
nand ( n256958 , n256956 , n256957 );
not ( n256959 , n40908 );
not ( n256960 , n251450 );
or ( n256961 , n256959 , n256960 );
not ( n256962 , n40908 );
nand ( n256963 , n256962 , n251443 );
nand ( n256964 , n256961 , n256963 );
buf ( n256965 , n54273 );
and ( n256966 , n256964 , n256965 );
not ( n256967 , n256964 );
and ( n256968 , n256967 , n253106 );
nor ( n256969 , n256966 , n256968 );
not ( n256970 , n31536 );
not ( n256971 , n256970 );
not ( n256972 , n247018 );
or ( n256973 , n256971 , n256972 );
nand ( n256974 , n247013 , n31536 );
nand ( n256975 , n256973 , n256974 );
not ( n256976 , n256975 );
not ( n256977 , n250113 );
and ( n256978 , n256976 , n256977 );
and ( n256979 , n256975 , n250113 );
nor ( n256980 , n256978 , n256979 );
nand ( n256981 , n256969 , n256980 );
or ( n256982 , n256958 , n256981 );
not ( n256983 , n256956 );
not ( n256984 , n256969 );
or ( n256985 , n256983 , n256984 );
nor ( n256986 , n256980 , n42443 );
nand ( n256987 , n256985 , n256986 );
nand ( n256988 , n237361 , n35899 );
nand ( n256989 , n256982 , n256987 , n256988 );
buf ( n256990 , n256989 );
buf ( n256991 , n240393 );
not ( n256992 , n256991 );
not ( n256993 , n252649 );
or ( n256994 , n256992 , n256993 );
or ( n256995 , n252649 , n256991 );
nand ( n256996 , n256994 , n256995 );
and ( n256997 , n256996 , n252652 );
not ( n256998 , n256996 );
and ( n256999 , n256998 , n252656 );
nor ( n257000 , n256997 , n256999 );
nand ( n257001 , n257000 , n254227 );
not ( n257002 , n227369 );
not ( n257003 , n247187 );
or ( n257004 , n257002 , n257003 );
not ( n257005 , n227369 );
nand ( n257006 , n257005 , n247195 );
nand ( n257007 , n257004 , n257006 );
and ( n257008 , n257007 , n254400 );
not ( n257009 , n257007 );
and ( n257010 , n257009 , n254403 );
nor ( n257011 , n257008 , n257010 );
not ( n257012 , n257011 );
not ( n257013 , n247853 );
not ( n257014 , n246188 );
or ( n257015 , n257013 , n257014 );
or ( n257016 , n246188 , n247853 );
nand ( n257017 , n257015 , n257016 );
and ( n257018 , n257017 , n246196 );
not ( n257019 , n257017 );
and ( n257020 , n257019 , n246193 );
nor ( n257021 , n257018 , n257020 );
not ( n257022 , n257021 );
nand ( n257023 , n257012 , n257022 );
or ( n257024 , n257001 , n257023 );
not ( n257025 , n257000 );
nand ( n257026 , n257025 , n253397 );
not ( n257027 , n257026 );
nand ( n257028 , n257027 , n257023 );
nand ( n257029 , n251465 , n38552 );
nand ( n257030 , n257024 , n257028 , n257029 );
buf ( n257031 , n257030 );
buf ( n257032 , n236925 );
xor ( n257033 , n257032 , n239298 );
and ( n257034 , n257033 , n239399 );
not ( n257035 , n257033 );
and ( n257036 , n257035 , n239391 );
nor ( n257037 , n257034 , n257036 );
nor ( n257038 , n257037 , n252070 );
not ( n257039 , n257038 );
not ( n257040 , n257039 );
not ( n257041 , n47857 );
not ( n257042 , n257041 );
not ( n257043 , n48676 );
or ( n257044 , n257042 , n257043 );
not ( n257045 , n257041 );
nand ( n257046 , n257045 , n48686 );
nand ( n257047 , n257044 , n257046 );
and ( n257048 , n257047 , n48806 );
not ( n257049 , n257047 );
and ( n257050 , n257049 , n48797 );
nor ( n257051 , n257048 , n257050 );
not ( n257052 , n257051 );
not ( n257053 , n238525 );
not ( n257054 , n241122 );
or ( n257055 , n257053 , n257054 );
not ( n257056 , n238525 );
nand ( n257057 , n257056 , n241131 );
nand ( n257058 , n257055 , n257057 );
and ( n257059 , n257058 , n241181 );
not ( n257060 , n257058 );
and ( n257061 , n257060 , n241180 );
nor ( n257062 , n257059 , n257061 );
not ( n257063 , n257062 );
nand ( n257064 , n257052 , n257063 );
not ( n257065 , n257064 );
and ( n257066 , n257040 , n257065 );
and ( n257067 , n41945 , n242473 );
nor ( n257068 , n257066 , n257067 );
nand ( n257069 , n257037 , n253393 );
not ( n257070 , n257069 );
nand ( n257071 , n257070 , n257051 );
nand ( n257072 , n257051 , n253393 );
not ( n257073 , n257072 );
nand ( n257074 , n257073 , n257062 );
nand ( n257075 , n257068 , n257071 , n257074 );
buf ( n257076 , n257075 );
nor ( n257077 , n254922 , n234818 );
not ( n257078 , n240975 );
not ( n257079 , n54134 );
or ( n257080 , n257078 , n257079 );
not ( n257081 , n240975 );
not ( n257082 , n249858 );
nand ( n257083 , n257081 , n257082 );
nand ( n257084 , n257080 , n257083 );
not ( n257085 , n257084 );
not ( n257086 , n54192 );
and ( n257087 , n257085 , n257086 );
and ( n257088 , n257084 , n231957 );
nor ( n257089 , n257087 , n257088 );
nand ( n257090 , n257077 , n254897 , n257089 );
not ( n257091 , n231444 );
not ( n257092 , n257091 );
not ( n257093 , n227134 );
and ( n257094 , n257092 , n257093 );
nor ( n257095 , n257089 , n42443 );
and ( n257096 , n257095 , n254896 );
nor ( n257097 , n257094 , n257096 );
not ( n257098 , n254922 );
nor ( n257099 , n257098 , n243204 );
not ( n257100 , n257089 );
nand ( n257101 , n257099 , n257100 );
nand ( n257102 , n257090 , n257097 , n257101 );
buf ( n257103 , n257102 );
not ( n257104 , n30976 );
not ( n257105 , n251465 );
or ( n257106 , n257104 , n257105 );
not ( n257107 , n238023 );
not ( n257108 , n226319 );
or ( n257109 , n257107 , n257108 );
not ( n257110 , n48557 );
nand ( n257111 , n257110 , n238024 );
nand ( n257112 , n257109 , n257111 );
not ( n257113 , n247689 );
and ( n257114 , n257112 , n257113 );
not ( n257115 , n257112 );
buf ( n257116 , n247689 );
and ( n257117 , n257115 , n257116 );
nor ( n257118 , n257114 , n257117 );
not ( n257119 , n257118 );
not ( n257120 , n31280 );
not ( n257121 , n247013 );
or ( n257122 , n257120 , n257121 );
or ( n257123 , n247013 , n31280 );
nand ( n257124 , n257122 , n257123 );
not ( n257125 , n257124 );
not ( n257126 , n250113 );
and ( n257127 , n257125 , n257126 );
not ( n257128 , n236886 );
and ( n257129 , n257124 , n257128 );
nor ( n257130 , n257127 , n257129 );
nand ( n257131 , n257119 , n257130 );
and ( n257132 , n257131 , n249551 );
not ( n257133 , n257131 );
not ( n257134 , n249551 );
and ( n257135 , n257133 , n257134 );
nor ( n257136 , n257132 , n257135 );
or ( n257137 , n257136 , n244837 );
nand ( n257138 , n257106 , n257137 );
buf ( n257139 , n257138 );
not ( n257140 , n25952 );
not ( n257141 , n46083 );
or ( n257142 , n257140 , n257141 );
nand ( n257143 , n250081 , n50241 );
and ( n257144 , n257143 , n248950 );
not ( n257145 , n257143 );
and ( n257146 , n257145 , n50231 );
nor ( n257147 , n257144 , n257146 );
not ( n257148 , n257147 );
not ( n257149 , n257148 );
not ( n257150 , n50274 );
or ( n257151 , n257149 , n257150 );
not ( n257152 , n257148 );
nand ( n257153 , n257152 , n228042 );
nand ( n257154 , n257151 , n257153 );
xor ( n257155 , n257154 , n50475 );
nand ( n257156 , n257155 , n254788 );
not ( n257157 , n42237 );
not ( n257158 , n234298 );
or ( n257159 , n257157 , n257158 );
not ( n257160 , n42236 );
or ( n257161 , n234298 , n257160 );
nand ( n257162 , n257159 , n257161 );
not ( n257163 , n257162 );
buf ( n257164 , n248446 );
not ( n257165 , n257164 );
and ( n257166 , n257163 , n257165 );
and ( n257167 , n257162 , n257164 );
nor ( n257168 , n257166 , n257167 );
not ( n257169 , n257168 );
and ( n257170 , n257156 , n257169 );
not ( n257171 , n257156 );
and ( n257172 , n257171 , n257168 );
nor ( n257173 , n257170 , n257172 );
buf ( n257174 , n238900 );
or ( n257175 , n257173 , n257174 );
nand ( n257176 , n257142 , n257175 );
buf ( n257177 , n257176 );
not ( n257178 , n255579 );
not ( n257179 , n238628 );
or ( n257180 , n257178 , n257179 );
not ( n257181 , n255579 );
nand ( n257182 , n257181 , n238620 );
nand ( n257183 , n257180 , n257182 );
xnor ( n257184 , n255756 , n255760 );
buf ( n257185 , n257184 );
and ( n257186 , n257183 , n257185 );
not ( n257187 , n257183 );
buf ( n257188 , n255762 );
and ( n257189 , n257187 , n257188 );
nor ( n257190 , n257186 , n257189 );
not ( n257191 , n257190 );
not ( n257192 , n245835 );
not ( n257193 , n39434 );
or ( n257194 , n257192 , n257193 );
not ( n257195 , n245835 );
nand ( n257196 , n257195 , n39444 );
nand ( n257197 , n257194 , n257196 );
and ( n257198 , n257197 , n248795 );
not ( n257199 , n257197 );
and ( n257200 , n257199 , n250255 );
nor ( n257201 , n257198 , n257200 );
not ( n257202 , n257201 );
nor ( n257203 , n257202 , n251190 );
not ( n257204 , n242570 );
not ( n257205 , n251145 );
not ( n257206 , n257205 );
not ( n257207 , n242520 );
or ( n257208 , n257206 , n257207 );
nand ( n257209 , n242527 , n251145 );
nand ( n257210 , n257208 , n257209 );
not ( n257211 , n257210 );
or ( n257212 , n257204 , n257211 );
or ( n257213 , n257210 , n242575 );
nand ( n257214 , n257212 , n257213 );
not ( n257215 , n257214 );
nand ( n257216 , n257191 , n257203 , n257215 );
not ( n257217 , n257201 );
not ( n257218 , n257190 );
not ( n257219 , n257218 );
or ( n257220 , n257217 , n257219 );
nor ( n257221 , n257215 , n46425 );
nand ( n257222 , n257220 , n257221 );
nand ( n257223 , n239240 , n30258 );
nand ( n257224 , n257216 , n257222 , n257223 );
buf ( n257225 , n257224 );
nand ( n257226 , n256124 , n249009 );
not ( n257227 , n239259 );
not ( n257228 , n248755 );
or ( n257229 , n257227 , n257228 );
not ( n257230 , n239259 );
nand ( n257231 , n257230 , n248762 );
nand ( n257232 , n257229 , n257231 );
and ( n257233 , n257232 , n252918 );
not ( n257234 , n257232 );
and ( n257235 , n257234 , n252923 );
nor ( n257236 , n257233 , n257235 );
not ( n257237 , n241804 );
not ( n257238 , n248901 );
or ( n257239 , n257237 , n257238 );
or ( n257240 , n250370 , n241804 );
nand ( n257241 , n257239 , n257240 );
and ( n257242 , n257241 , n248904 );
not ( n257243 , n257241 );
and ( n257244 , n257243 , n248907 );
nor ( n257245 , n257242 , n257244 );
not ( n257246 , n257245 );
nand ( n257247 , n257236 , n257246 );
or ( n257248 , n257226 , n257247 );
nand ( n257249 , n256125 , n257247 );
nand ( n257250 , n31577 , n26022 );
nand ( n257251 , n257248 , n257249 , n257250 );
buf ( n257252 , n257251 );
not ( n257253 , n43866 );
not ( n257254 , n252552 );
or ( n257255 , n257253 , n257254 );
not ( n257256 , n43866 );
nand ( n257257 , n257256 , n252561 );
nand ( n257258 , n257255 , n257257 );
and ( n257259 , n257258 , n255673 );
not ( n257260 , n257258 );
and ( n257261 , n257260 , n255676 );
nor ( n257262 , n257259 , n257261 );
not ( n257263 , n28518 );
not ( n257264 , n254866 );
or ( n257265 , n257263 , n257264 );
not ( n257266 , n28518 );
nand ( n257267 , n257266 , n254873 );
nand ( n257268 , n257265 , n257267 );
and ( n257269 , n257268 , n256716 );
not ( n257270 , n257268 );
and ( n257271 , n257270 , n256712 );
nor ( n257272 , n257269 , n257271 );
not ( n257273 , n257272 );
nand ( n257274 , n257262 , n257273 );
not ( n257275 , n249151 );
not ( n257276 , n257275 );
not ( n257277 , n244776 );
or ( n257278 , n257276 , n257277 );
not ( n257279 , n257275 );
nand ( n257280 , n257279 , n244768 );
nand ( n257281 , n257278 , n257280 );
and ( n257282 , n257281 , n252934 );
not ( n257283 , n257281 );
and ( n257284 , n257283 , n249059 );
nor ( n257285 , n257282 , n257284 );
nor ( n257286 , n257285 , n226003 );
not ( n257287 , n257286 );
or ( n257288 , n257274 , n257287 );
not ( n257289 , n257285 );
nor ( n257290 , n257289 , n233972 );
nand ( n257291 , n257274 , n257290 );
nand ( n257292 , n35431 , n30741 );
nand ( n257293 , n257288 , n257291 , n257292 );
buf ( n257294 , n257293 );
buf ( n257295 , n27949 );
buf ( n257296 , n27786 );
not ( n257297 , n251928 );
not ( n257298 , n245994 );
not ( n257299 , n257298 );
not ( n257300 , n257299 );
or ( n257301 , n257297 , n257300 );
not ( n257302 , n251928 );
nand ( n257303 , n257302 , n246011 );
nand ( n257304 , n257301 , n257303 );
and ( n257305 , n257304 , n246017 );
not ( n257306 , n257304 );
not ( n257307 , n245950 );
not ( n257308 , n257307 );
and ( n257309 , n257306 , n257308 );
nor ( n257310 , n257305 , n257309 );
nand ( n257311 , n256553 , n257310 );
nand ( n257312 , n256540 , n244393 );
or ( n257313 , n257311 , n257312 );
not ( n257314 , n256540 );
not ( n257315 , n256553 );
or ( n257316 , n257314 , n257315 );
nor ( n257317 , n257310 , n252070 );
nand ( n257318 , n257316 , n257317 );
nand ( n257319 , n35431 , n32100 );
nand ( n257320 , n257313 , n257318 , n257319 );
buf ( n257321 , n257320 );
not ( n257322 , n244399 );
nand ( n257323 , n257322 , n251512 );
not ( n257324 , n236385 );
not ( n257325 , n51845 );
and ( n257326 , n257324 , n257325 );
and ( n257327 , n245201 , n51845 );
nor ( n257328 , n257326 , n257327 );
not ( n257329 , n257328 );
not ( n257330 , n245211 );
or ( n257331 , n257329 , n257330 );
or ( n257332 , n245211 , n257328 );
nand ( n257333 , n257331 , n257332 );
not ( n257334 , n257333 );
nand ( n257335 , n251555 , n257334 );
or ( n257336 , n257323 , n257335 );
not ( n257337 , n251555 );
not ( n257338 , n251512 );
or ( n257339 , n257337 , n257338 );
nor ( n257340 , n257334 , n39763 );
nand ( n257341 , n257339 , n257340 );
nand ( n257342 , n253486 , n207591 );
nand ( n257343 , n257336 , n257341 , n257342 );
buf ( n257344 , n257343 );
buf ( n257345 , RI19a24ed8_2782);
not ( n257346 , n257345 );
nor ( n257347 , n25335 , n251562 );
not ( n257348 , n257347 );
or ( n257349 , n257346 , n257348 );
or ( n257350 , n25328 , n251562 );
not ( n257351 , n257350 );
buf ( n257352 , RI19a250b8_2781);
nand ( n257353 , n257351 , n257352 );
nand ( n257354 , n257349 , n257353 );
buf ( n257355 , n257354 );
buf ( n257356 , n37860 );
not ( n257357 , n204869 );
not ( n257358 , n46083 );
or ( n257359 , n257357 , n257358 );
not ( n257360 , n242205 );
not ( n257361 , n257360 );
not ( n257362 , n246976 );
not ( n257363 , n257362 );
not ( n257364 , n242148 );
or ( n257365 , n257363 , n257364 );
nand ( n257366 , n242155 , n246976 );
nand ( n257367 , n257365 , n257366 );
not ( n257368 , n257367 );
or ( n257369 , n257361 , n257368 );
or ( n257370 , n257367 , n242202 );
nand ( n257371 , n257369 , n257370 );
not ( n257372 , n243303 );
not ( n257373 , n257372 );
not ( n257374 , n250805 );
or ( n257375 , n257373 , n257374 );
nand ( n257376 , n250806 , n243303 );
nand ( n257377 , n257375 , n257376 );
not ( n257378 , n39052 );
not ( n257379 , n257378 );
and ( n257380 , n257377 , n257379 );
not ( n257381 , n257377 );
buf ( n257382 , n39059 );
and ( n257383 , n257381 , n257382 );
nor ( n257384 , n257380 , n257383 );
nand ( n257385 , n257371 , n257384 );
not ( n257386 , n247477 );
not ( n257387 , n243510 );
or ( n257388 , n257386 , n257387 );
not ( n257389 , n247477 );
nand ( n257390 , n257389 , n243503 );
nand ( n257391 , n257388 , n257390 );
and ( n257392 , n257391 , n248481 );
not ( n257393 , n257391 );
and ( n257394 , n257393 , n248478 );
nor ( n257395 , n257392 , n257394 );
not ( n257396 , n257395 );
and ( n257397 , n257385 , n257396 );
not ( n257398 , n257385 );
and ( n257399 , n257398 , n257395 );
nor ( n257400 , n257397 , n257399 );
or ( n257401 , n257400 , n238223 );
nand ( n257402 , n257359 , n257401 );
buf ( n257403 , n257402 );
buf ( n257404 , n204655 );
buf ( n257405 , n40115 );
not ( n257406 , RI19acdf10_2225);
or ( n257407 , n25328 , n257406 );
not ( n257408 , RI19ac52e8_2290);
or ( n257409 , n25335 , n257408 );
nand ( n257410 , n257407 , n257409 );
buf ( n257411 , n257410 );
not ( n257412 , n248503 );
not ( n257413 , n243659 );
or ( n257414 , n257412 , n257413 );
or ( n257415 , n243659 , n248503 );
nand ( n257416 , n257414 , n257415 );
and ( n257417 , n257416 , n251856 );
not ( n257418 , n257416 );
and ( n257419 , n257418 , n251846 );
nor ( n257420 , n257417 , n257419 );
not ( n257421 , n257420 );
not ( n257422 , n257421 );
not ( n257423 , n255627 );
not ( n257424 , n257423 );
or ( n257425 , n257422 , n257424 );
not ( n257426 , n50005 );
not ( n257427 , n48875 );
or ( n257428 , n257426 , n257427 );
not ( n257429 , n50005 );
nand ( n257430 , n257429 , n48883 );
nand ( n257431 , n257428 , n257430 );
and ( n257432 , n257431 , n246478 );
not ( n257433 , n257431 );
and ( n257434 , n257433 , n246479 );
nor ( n257435 , n257432 , n257434 );
not ( n257436 , n257435 );
nor ( n257437 , n257436 , n235050 );
nand ( n257438 , n257425 , n257437 );
nor ( n257439 , n257435 , n257420 );
nand ( n257440 , n255630 , n257439 );
nand ( n257441 , n241976 , n38029 );
nand ( n257442 , n257438 , n257440 , n257441 );
buf ( n257443 , n257442 );
nor ( n257444 , n254012 , n39763 );
not ( n257445 , n257444 );
not ( n257446 , n240431 );
not ( n257447 , n252644 );
or ( n257448 , n257446 , n257447 );
not ( n257449 , n240431 );
nand ( n257450 , n257449 , n252649 );
nand ( n257451 , n257448 , n257450 );
and ( n257452 , n257451 , n252656 );
not ( n257453 , n257451 );
and ( n257454 , n257453 , n252652 );
nor ( n257455 , n257452 , n257454 );
nand ( n257456 , n257455 , n254024 );
or ( n257457 , n257445 , n257456 );
not ( n257458 , n257455 );
not ( n257459 , n254012 );
not ( n257460 , n257459 );
or ( n257461 , n257458 , n257460 );
nand ( n257462 , n254023 , n235051 );
not ( n257463 , n257462 );
nand ( n257464 , n257461 , n257463 );
nand ( n257465 , n237714 , n46566 );
nand ( n257466 , n257457 , n257464 , n257465 );
buf ( n257467 , n257466 );
or ( n257468 , n25328 , n25337 );
not ( n257469 , RI19aca4f0_2253);
or ( n257470 , n25335 , n257469 );
nand ( n257471 , n257468 , n257470 );
buf ( n257472 , n257471 );
not ( n257473 , RI19acda60_2227);
or ( n257474 , n25328 , n257473 );
or ( n257475 , n25335 , n242877 );
nand ( n257476 , n257474 , n257475 );
buf ( n257477 , n257476 );
or ( n257478 , n233507 , n249628 );
not ( n257479 , RI19ab9a38_2383);
or ( n257480 , n25335 , n257479 );
nand ( n257481 , n257478 , n257480 );
buf ( n257482 , n257481 );
not ( n257483 , n206058 );
not ( n257484 , n257483 );
not ( n257485 , n254866 );
or ( n257486 , n257484 , n257485 );
not ( n257487 , n257483 );
nand ( n257488 , n257487 , n254873 );
nand ( n257489 , n257486 , n257488 );
and ( n257490 , n257489 , n256716 );
not ( n257491 , n257489 );
and ( n257492 , n257491 , n256711 );
nor ( n257493 , n257490 , n257492 );
not ( n257494 , n257493 );
nand ( n257495 , n257494 , n254013 );
not ( n257496 , n241011 );
not ( n257497 , n257496 );
not ( n257498 , n41632 );
or ( n257499 , n257497 , n257498 );
or ( n257500 , n219397 , n257496 );
nand ( n257501 , n257499 , n257500 );
and ( n257502 , n257501 , n41930 );
not ( n257503 , n257501 );
and ( n257504 , n257503 , n41935 );
nor ( n257505 , n257502 , n257504 );
nand ( n257506 , n257505 , n242897 );
or ( n257507 , n257495 , n257506 );
not ( n257508 , n257505 );
not ( n257509 , n257493 );
not ( n257510 , n257509 );
or ( n257511 , n257508 , n257510 );
nand ( n257512 , n257511 , n243207 );
nand ( n257513 , n31576 , n28027 );
nand ( n257514 , n257507 , n257512 , n257513 );
buf ( n257515 , n257514 );
not ( n257516 , n43688 );
not ( n257517 , n257516 );
not ( n257518 , n242270 );
or ( n257519 , n257517 , n257518 );
not ( n257520 , n257516 );
nand ( n257521 , n257520 , n252503 );
nand ( n257522 , n257519 , n257521 );
and ( n257523 , n257522 , n252562 );
not ( n257524 , n257522 );
and ( n257525 , n257524 , n252553 );
nor ( n257526 , n257523 , n257525 );
not ( n257527 , n238635 );
nand ( n257528 , n257526 , n257527 );
buf ( n257529 , n47214 );
not ( n257530 , n257529 );
not ( n257531 , n254076 );
or ( n257532 , n257530 , n257531 );
or ( n257533 , n245170 , n257529 );
nand ( n257534 , n257532 , n257533 );
and ( n257535 , n257534 , n254080 );
not ( n257536 , n257534 );
and ( n257537 , n257536 , n254083 );
nor ( n257538 , n257535 , n257537 );
not ( n257539 , n257538 );
not ( n257540 , n249575 );
not ( n257541 , n224180 );
not ( n257542 , n257541 );
or ( n257543 , n257540 , n257542 );
not ( n257544 , n249575 );
nand ( n257545 , n257544 , n243006 );
nand ( n257546 , n257543 , n257545 );
and ( n257547 , n257546 , n243199 );
not ( n257548 , n257546 );
and ( n257549 , n257548 , n243198 );
nor ( n257550 , n257547 , n257549 );
nand ( n257551 , n257539 , n257550 );
or ( n257552 , n257528 , n257551 );
not ( n257553 , n257526 );
not ( n257554 , n257539 );
or ( n257555 , n257553 , n257554 );
nor ( n257556 , n257550 , n53680 );
nand ( n257557 , n257555 , n257556 );
nand ( n257558 , n39766 , n204408 );
nand ( n257559 , n257552 , n257557 , n257558 );
buf ( n257560 , n257559 );
not ( n257561 , n205007 );
not ( n257562 , n31577 );
or ( n257563 , n257561 , n257562 );
not ( n257564 , n245441 );
not ( n257565 , n241962 );
or ( n257566 , n257564 , n257565 );
not ( n257567 , n245441 );
nand ( n257568 , n257567 , n250442 );
nand ( n257569 , n257566 , n257568 );
and ( n257570 , n257569 , n250498 );
not ( n257571 , n257569 );
buf ( n257572 , n255291 );
and ( n257573 , n257571 , n257572 );
nor ( n257574 , n257570 , n257573 );
not ( n257575 , n247519 );
not ( n257576 , n243801 );
or ( n257577 , n257575 , n257576 );
not ( n257578 , n247519 );
nand ( n257579 , n257578 , n243810 );
nand ( n257580 , n257577 , n257579 );
and ( n257581 , n257580 , n243960 );
not ( n257582 , n257580 );
and ( n257583 , n257582 , n243954 );
nor ( n257584 , n257581 , n257583 );
not ( n257585 , n257584 );
nand ( n257586 , n257574 , n257585 );
not ( n257587 , n247733 );
not ( n257588 , n238133 );
not ( n257589 , n247727 );
or ( n257590 , n257588 , n257589 );
or ( n257591 , n247727 , n238133 );
nand ( n257592 , n257590 , n257591 );
not ( n257593 , n257592 );
or ( n257594 , n257587 , n257593 );
or ( n257595 , n257592 , n247733 );
nand ( n257596 , n257594 , n257595 );
and ( n257597 , n257586 , n257596 );
not ( n257598 , n257586 );
not ( n257599 , n257596 );
and ( n257600 , n257598 , n257599 );
nor ( n257601 , n257597 , n257600 );
or ( n257602 , n257601 , n237358 );
nand ( n257603 , n257563 , n257602 );
buf ( n257604 , n257603 );
not ( n257605 , RI19a952a0_2646);
or ( n257606 , n25328 , n257605 );
not ( n257607 , RI19a8af08_2718);
or ( n257608 , n226822 , n257607 );
nand ( n257609 , n257606 , n257608 );
buf ( n257610 , n257609 );
buf ( n257611 , n215590 );
not ( n257612 , n257611 );
not ( n257613 , n50027 );
or ( n257614 , n257612 , n257613 );
or ( n257615 , n50027 , n257611 );
nand ( n257616 , n257614 , n257615 );
not ( n257617 , n257616 );
not ( n257618 , n234514 );
and ( n257619 , n257617 , n257618 );
and ( n257620 , n257616 , n234514 );
nor ( n257621 , n257619 , n257620 );
nand ( n257622 , n257621 , n244809 );
not ( n257623 , n222774 );
not ( n257624 , n244009 );
or ( n257625 , n257623 , n257624 );
or ( n257626 , n244459 , n222774 );
nand ( n257627 , n257625 , n257626 );
and ( n257628 , n257627 , n244056 );
not ( n257629 , n257627 );
buf ( n257630 , n253557 );
and ( n257631 , n257629 , n257630 );
nor ( n257632 , n257628 , n257631 );
not ( n257633 , n257632 );
not ( n257634 , n247664 );
not ( n257635 , n48015 );
or ( n257636 , n257634 , n257635 );
not ( n257637 , n247664 );
nand ( n257638 , n257637 , n48019 );
nand ( n257639 , n257636 , n257638 );
and ( n257640 , n257639 , n48238 );
not ( n257641 , n257639 );
and ( n257642 , n257641 , n48234 );
nor ( n257643 , n257640 , n257642 );
nand ( n257644 , n257633 , n257643 );
or ( n257645 , n257622 , n257644 );
nor ( n257646 , n257621 , n50944 );
nand ( n257647 , n257646 , n257644 );
nand ( n257648 , n39766 , n37890 );
nand ( n257649 , n257645 , n257647 , n257648 );
buf ( n257650 , n257649 );
not ( n257651 , n248909 );
not ( n257652 , n237104 );
not ( n257653 , n253074 );
or ( n257654 , n257652 , n257653 );
not ( n257655 , n237104 );
nand ( n257656 , n257655 , n253073 );
nand ( n257657 , n257654 , n257656 );
not ( n257658 , n249195 );
not ( n257659 , n257658 );
and ( n257660 , n257657 , n257659 );
not ( n257661 , n257657 );
and ( n257662 , n257661 , n257658 );
nor ( n257663 , n257660 , n257662 );
not ( n257664 , n257663 );
not ( n257665 , n257664 );
or ( n257666 , n257651 , n257665 );
nor ( n257667 , n248978 , n243204 );
nand ( n257668 , n257666 , n257667 );
nand ( n257669 , n248909 , n237385 );
not ( n257670 , n257669 );
nand ( n257671 , n257670 , n248978 , n257664 );
nand ( n257672 , n48251 , n34251 );
nand ( n257673 , n257668 , n257671 , n257672 );
buf ( n257674 , n257673 );
not ( n257675 , n242842 );
not ( n257676 , n242969 );
or ( n257677 , n257675 , n257676 );
nand ( n257678 , n242977 , n242843 );
nand ( n257679 , n257677 , n257678 );
not ( n257680 , n257679 );
not ( n257681 , n246963 );
and ( n257682 , n257680 , n257681 );
and ( n257683 , n257679 , n254060 );
nor ( n257684 , n257682 , n257683 );
nor ( n257685 , n257684 , n31572 );
not ( n257686 , n257685 );
not ( n257687 , n38814 );
not ( n257688 , n251298 );
or ( n257689 , n257687 , n257688 );
not ( n257690 , n38814 );
nand ( n257691 , n257690 , n251313 );
nand ( n257692 , n257689 , n257691 );
and ( n257693 , n257692 , n256008 );
not ( n257694 , n257692 );
and ( n257695 , n257694 , n256012 );
nor ( n257696 , n257693 , n257695 );
not ( n257697 , n222860 );
not ( n257698 , n244054 );
or ( n257699 , n257697 , n257698 );
not ( n257700 , n222860 );
nand ( n257701 , n257700 , n253557 );
nand ( n257702 , n257699 , n257701 );
not ( n257703 , n245517 );
and ( n257704 , n257702 , n257703 );
not ( n257705 , n257702 );
not ( n257706 , n253560 );
and ( n257707 , n257705 , n257706 );
nor ( n257708 , n257704 , n257707 );
nand ( n257709 , n257696 , n257708 );
or ( n257710 , n257686 , n257709 );
not ( n257711 , n257708 );
not ( n257712 , n257684 );
not ( n257713 , n257712 );
or ( n257714 , n257711 , n257713 );
nor ( n257715 , n257696 , n46425 );
nand ( n257716 , n257714 , n257715 );
nand ( n257717 , n49054 , n37837 );
nand ( n257718 , n257710 , n257716 , n257717 );
buf ( n257719 , n257718 );
not ( n257720 , n37479 );
and ( n257721 , n252418 , n252438 );
not ( n257722 , n252418 );
and ( n257723 , n257722 , n252441 );
nor ( n257724 , n257721 , n257723 );
not ( n257725 , n257724 );
or ( n257726 , n257720 , n257725 );
or ( n257727 , n257724 , n37479 );
nand ( n257728 , n257726 , n257727 );
buf ( n257729 , n242307 );
and ( n257730 , n257728 , n257729 );
not ( n257731 , n257728 );
not ( n257732 , n257729 );
and ( n257733 , n257731 , n257732 );
nor ( n257734 , n257730 , n257733 );
not ( n257735 , n257734 );
not ( n257736 , n246997 );
not ( n257737 , n257736 );
not ( n257738 , n242148 );
or ( n257739 , n257737 , n257738 );
not ( n257740 , n257736 );
nand ( n257741 , n257740 , n242155 );
nand ( n257742 , n257739 , n257741 );
and ( n257743 , n257742 , n242206 );
not ( n257744 , n257742 );
and ( n257745 , n257744 , n257360 );
nor ( n257746 , n257743 , n257745 );
not ( n257747 , n257746 );
nand ( n257748 , n257735 , n257747 );
not ( n257749 , n228259 );
not ( n257750 , n35804 );
or ( n257751 , n257749 , n257750 );
not ( n257752 , n228259 );
nand ( n257753 , n257752 , n35811 );
nand ( n257754 , n257751 , n257753 );
and ( n257755 , n257754 , n253336 );
not ( n257756 , n257754 );
not ( n257757 , n252081 );
and ( n257758 , n257756 , n257757 );
nor ( n257759 , n257755 , n257758 );
nand ( n257760 , n257759 , n241459 );
or ( n257761 , n257748 , n257760 );
nor ( n257762 , n257759 , n254226 );
nand ( n257763 , n257748 , n257762 );
buf ( n257764 , n35431 );
nand ( n257765 , n257764 , n28091 );
nand ( n257766 , n257761 , n257763 , n257765 );
buf ( n257767 , n257766 );
not ( n257768 , n243433 );
not ( n257769 , n205649 );
nor ( n257770 , n257768 , n257769 );
not ( n257771 , n243417 );
not ( n257772 , n54744 );
not ( n257773 , n245517 );
or ( n257774 , n257772 , n257773 );
or ( n257775 , n245517 , n54744 );
nand ( n257776 , n257774 , n257775 );
not ( n257777 , n257776 );
not ( n257778 , n245524 );
and ( n257779 , n257777 , n257778 );
and ( n257780 , n251162 , n257776 );
nor ( n257781 , n257779 , n257780 );
nand ( n257782 , n257770 , n257771 , n257781 );
not ( n257783 , n257771 );
not ( n257784 , n243433 );
or ( n257785 , n257783 , n257784 );
nor ( n257786 , n257781 , n234021 );
nand ( n257787 , n257785 , n257786 );
nand ( n257788 , n50615 , n205151 );
nand ( n257789 , n257782 , n257787 , n257788 );
buf ( n257790 , n257789 );
buf ( n257791 , n37613 );
not ( n257792 , n55146 );
nand ( n257793 , n250750 , n257792 );
not ( n257794 , n255724 );
not ( n257795 , n256131 );
or ( n257796 , n257794 , n257795 );
or ( n257797 , n249541 , n255724 );
nand ( n257798 , n257796 , n257797 );
and ( n257799 , n257798 , n249549 );
not ( n257800 , n257798 );
and ( n257801 , n257800 , n249546 );
nor ( n257802 , n257799 , n257801 );
nand ( n257803 , n257802 , n253901 );
or ( n257804 , n257793 , n257803 );
nand ( n257805 , n250751 , n257803 );
nand ( n257806 , n255116 , n205168 );
nand ( n257807 , n257804 , n257805 , n257806 );
buf ( n257808 , n257807 );
buf ( n257809 , n32832 );
not ( n257810 , n32648 );
not ( n257811 , n233501 );
or ( n257812 , n257810 , n257811 );
not ( n257813 , n253151 );
not ( n257814 , n223827 );
or ( n257815 , n257813 , n257814 );
not ( n257816 , n253151 );
nand ( n257817 , n257816 , n46074 );
nand ( n257818 , n257815 , n257817 );
and ( n257819 , n257818 , n244508 );
not ( n257820 , n257818 );
and ( n257821 , n257820 , n244509 );
nor ( n257822 , n257819 , n257821 );
not ( n257823 , n257822 );
not ( n257824 , n41575 );
not ( n257825 , n233026 );
or ( n257826 , n257824 , n257825 );
not ( n257827 , n41575 );
nand ( n257828 , n257827 , n233035 );
nand ( n257829 , n257826 , n257828 );
and ( n257830 , n257829 , n233091 );
not ( n257831 , n257829 );
and ( n257832 , n257831 , n233084 );
nor ( n257833 , n257830 , n257832 );
not ( n257834 , n257833 );
nand ( n257835 , n257823 , n257834 );
not ( n257836 , n251647 );
not ( n257837 , n46941 );
or ( n257838 , n257836 , n257837 );
not ( n257839 , n251647 );
nand ( n257840 , n257839 , n46950 );
nand ( n257841 , n257838 , n257840 );
and ( n257842 , n257841 , n224925 );
not ( n257843 , n257841 );
and ( n257844 , n257843 , n47157 );
nor ( n257845 , n257842 , n257844 );
not ( n257846 , n257845 );
and ( n257847 , n257835 , n257846 );
not ( n257848 , n257835 );
and ( n257849 , n257848 , n257845 );
nor ( n257850 , n257847 , n257849 );
buf ( n257851 , n253544 );
or ( n257852 , n257850 , n257851 );
nand ( n257853 , n257812 , n257852 );
buf ( n257854 , n257853 );
not ( n257855 , n234813 );
not ( n257856 , n234540 );
nand ( n257857 , n257855 , n257856 );
not ( n257858 , n244932 );
not ( n257859 , n34439 );
or ( n257860 , n257858 , n257859 );
not ( n257861 , n244932 );
nand ( n257862 , n257861 , n34448 );
nand ( n257863 , n257860 , n257862 );
and ( n257864 , n257863 , n33709 );
not ( n257865 , n257863 );
and ( n257866 , n257865 , n235042 );
nor ( n257867 , n257864 , n257866 );
nand ( n257868 , n257867 , n241373 );
or ( n257869 , n257857 , n257868 );
nor ( n257870 , n257867 , n31572 );
nand ( n257871 , n257857 , n257870 );
nand ( n257872 , n234024 , n206401 );
nand ( n257873 , n257869 , n257871 , n257872 );
buf ( n257874 , n257873 );
buf ( n257875 , n35842 );
buf ( n257876 , n25620 );
buf ( n257877 , n26459 );
buf ( n257878 , n32426 );
not ( n257879 , n242201 );
not ( n257880 , n236861 );
and ( n257881 , n257879 , n257880 );
and ( n257882 , n242201 , n236861 );
nor ( n257883 , n257881 , n257882 );
and ( n257884 , n257883 , n255160 );
not ( n257885 , n257883 );
and ( n257886 , n257885 , n255163 );
nor ( n257887 , n257884 , n257886 );
nand ( n257888 , n257887 , n254528 );
not ( n257889 , n253827 );
not ( n257890 , n257889 );
not ( n257891 , n46506 );
or ( n257892 , n257890 , n257891 );
not ( n257893 , n257889 );
nand ( n257894 , n257893 , n46514 );
nand ( n257895 , n257892 , n257894 );
and ( n257896 , n257895 , n224478 );
not ( n257897 , n257895 );
and ( n257898 , n257897 , n251333 );
nor ( n257899 , n257896 , n257898 );
not ( n257900 , n257899 );
not ( n257901 , n252414 );
not ( n257902 , n240893 );
not ( n257903 , n257902 );
not ( n257904 , n250626 );
nand ( n257905 , n257904 , n37586 );
not ( n257906 , n257905 );
or ( n257907 , n257903 , n257906 );
or ( n257908 , n257905 , n257902 );
nand ( n257909 , n257907 , n257908 );
not ( n257910 , n257909 );
nand ( n257911 , n252391 , n37542 );
not ( n257912 , n257911 );
not ( n257913 , n240874 );
and ( n257914 , n257912 , n257913 );
not ( n257915 , n37541 );
nand ( n257916 , n257915 , n252391 );
and ( n257917 , n257916 , n240874 );
nor ( n257918 , n257914 , n257917 );
not ( n257919 , n257918 );
or ( n257920 , n257910 , n257919 );
or ( n257921 , n257918 , n257909 );
nand ( n257922 , n257920 , n257921 );
nand ( n257923 , n37693 , n250658 );
and ( n257924 , n257923 , n240852 );
not ( n257925 , n257923 );
and ( n257926 , n257925 , n240853 );
nor ( n257927 , n257924 , n257926 );
xor ( n257928 , n257922 , n257927 );
not ( n257929 , n240929 );
nand ( n257930 , n252428 , n37361 );
not ( n257931 , n257930 );
or ( n257932 , n257929 , n257931 );
or ( n257933 , n257930 , n240929 );
nand ( n257934 , n257932 , n257933 );
not ( n257935 , n257934 );
not ( n257936 , n240908 );
not ( n257937 , n240834 );
nand ( n257938 , n257937 , n37475 );
not ( n257939 , n257938 );
and ( n257940 , n257936 , n257939 );
and ( n257941 , n240908 , n257938 );
nor ( n257942 , n257940 , n257941 );
not ( n257943 , n257942 );
or ( n257944 , n257935 , n257943 );
or ( n257945 , n257942 , n257934 );
nand ( n257946 , n257944 , n257945 );
and ( n257947 , n257928 , n257946 );
not ( n257948 , n257928 );
not ( n257949 , n257946 );
and ( n257950 , n257948 , n257949 );
nor ( n257951 , n257947 , n257950 );
buf ( n257952 , n257951 );
not ( n257953 , n257952 );
or ( n257954 , n257901 , n257953 );
not ( n257955 , n252414 );
not ( n257956 , n257951 );
nand ( n257957 , n257955 , n257956 );
nand ( n257958 , n257954 , n257957 );
not ( n257959 , n39598 );
not ( n257960 , n257959 );
and ( n257961 , n257958 , n257960 );
not ( n257962 , n257958 );
not ( n257963 , n39595 );
not ( n257964 , n257963 );
and ( n257965 , n257962 , n257964 );
nor ( n257966 , n257961 , n257965 );
not ( n257967 , n257966 );
nand ( n257968 , n257900 , n257967 );
or ( n257969 , n257888 , n257968 );
not ( n257970 , n257900 );
not ( n257971 , n257887 );
or ( n257972 , n257970 , n257971 );
nand ( n257973 , n257966 , n38638 );
not ( n257974 , n257973 );
nand ( n257975 , n257972 , n257974 );
nand ( n257976 , n31577 , n33879 );
nand ( n257977 , n257969 , n257975 , n257976 );
buf ( n257978 , n257977 );
not ( n257979 , n41245 );
not ( n257980 , n233501 );
or ( n257981 , n257979 , n257980 );
not ( n257982 , n248284 );
not ( n257983 , n247163 );
not ( n257984 , n257983 );
not ( n257985 , n253474 );
or ( n257986 , n257984 , n257985 );
nand ( n257987 , n248276 , n247163 );
nand ( n257988 , n257986 , n257987 );
not ( n257989 , n257988 );
or ( n257990 , n257982 , n257989 );
or ( n257991 , n257988 , n248284 );
nand ( n257992 , n257990 , n257991 );
not ( n257993 , n250790 );
not ( n257994 , n257993 );
not ( n257995 , n251154 );
or ( n257996 , n257994 , n257995 );
not ( n257997 , n257993 );
nand ( n257998 , n257997 , n251253 );
nand ( n257999 , n257996 , n257998 );
and ( n258000 , n257999 , n251314 );
not ( n258001 , n257999 );
and ( n258002 , n258001 , n251299 );
nor ( n258003 , n258000 , n258002 );
not ( n258004 , n258003 );
nand ( n258005 , n257992 , n258004 );
not ( n258006 , n36403 );
not ( n258007 , n253855 );
or ( n258008 , n258006 , n258007 );
not ( n258009 , n36403 );
nand ( n258010 , n258009 , n253863 );
nand ( n258011 , n258008 , n258010 );
not ( n258012 , n239858 );
not ( n258013 , n258012 );
and ( n258014 , n258011 , n258013 );
not ( n258015 , n258011 );
and ( n258016 , n258015 , n258012 );
nor ( n258017 , n258014 , n258016 );
not ( n258018 , n258017 );
and ( n258019 , n258005 , n258018 );
not ( n258020 , n258005 );
and ( n258021 , n258020 , n258017 );
nor ( n258022 , n258019 , n258021 );
or ( n258023 , n258022 , n257851 );
nand ( n258024 , n257981 , n258023 );
buf ( n258025 , n258024 );
not ( n258026 , n33543 );
not ( n258027 , n245702 );
or ( n258028 , n258026 , n258027 );
nand ( n258029 , n249095 , n249115 );
buf ( n258030 , n236732 );
not ( n258031 , n258030 );
not ( n258032 , n43218 );
not ( n258033 , n258032 );
not ( n258034 , n258033 );
or ( n258035 , n258031 , n258034 );
or ( n258036 , n43219 , n258030 );
nand ( n258037 , n258035 , n258036 );
buf ( n258038 , n45023 );
not ( n258039 , n258038 );
and ( n258040 , n258037 , n258039 );
not ( n258041 , n258037 );
and ( n258042 , n258041 , n45027 );
nor ( n258043 , n258040 , n258042 );
not ( n258044 , n258043 );
and ( n258045 , n258029 , n258044 );
not ( n258046 , n258029 );
and ( n258047 , n258046 , n258043 );
nor ( n258048 , n258045 , n258047 );
or ( n258049 , n258048 , n253544 );
nand ( n258050 , n258028 , n258049 );
buf ( n258051 , n258050 );
not ( n258052 , n239319 );
not ( n258053 , n252922 );
or ( n258054 , n258052 , n258053 );
not ( n258055 , n252917 );
or ( n258056 , n258055 , n239319 );
nand ( n258057 , n258054 , n258056 );
buf ( n258058 , n42149 );
and ( n258059 , n258057 , n258058 );
not ( n258060 , n258057 );
buf ( n258061 , n42156 );
and ( n258062 , n258060 , n258061 );
nor ( n258063 , n258059 , n258062 );
not ( n258064 , n258063 );
nand ( n258065 , n258064 , n249009 );
buf ( n258066 , n228965 );
not ( n258067 , n258066 );
not ( n258068 , n258067 );
not ( n258069 , n256761 );
or ( n258070 , n258068 , n258069 );
nand ( n258071 , n256762 , n258066 );
nand ( n258072 , n258070 , n258071 );
and ( n258073 , n258072 , n256765 );
not ( n258074 , n258072 );
and ( n258075 , n258074 , n253673 );
nor ( n258076 , n258073 , n258075 );
buf ( n258077 , n256862 );
not ( n258078 , n258077 );
not ( n258079 , n52941 );
not ( n258080 , n246882 );
or ( n258081 , n258079 , n258080 );
nand ( n258082 , n246891 , n230701 );
nand ( n258083 , n258081 , n258082 );
not ( n258084 , n258083 );
or ( n258085 , n258078 , n258084 );
or ( n258086 , n258077 , n258083 );
nand ( n258087 , n258085 , n258086 );
not ( n258088 , n258087 );
nand ( n258089 , n258076 , n258088 );
or ( n258090 , n258065 , n258089 );
not ( n258091 , n258088 );
not ( n258092 , n258064 );
or ( n258093 , n258091 , n258092 );
nor ( n258094 , n258076 , n33253 );
nand ( n258095 , n258093 , n258094 );
nand ( n258096 , n31577 , n42598 );
nand ( n258097 , n258090 , n258095 , n258096 );
buf ( n258098 , n258097 );
not ( n258099 , n31489 );
not ( n258100 , n51381 );
or ( n258101 , n258099 , n258100 );
not ( n258102 , n38760 );
not ( n258103 , n258102 );
not ( n258104 , n251298 );
or ( n258105 , n258103 , n258104 );
not ( n258106 , n258102 );
nand ( n258107 , n258106 , n251313 );
nand ( n258108 , n258105 , n258107 );
and ( n258109 , n258108 , n256008 );
not ( n258110 , n258108 );
and ( n258111 , n258110 , n256012 );
nor ( n258112 , n258109 , n258111 );
not ( n258113 , n258112 );
not ( n258114 , n242108 );
not ( n258115 , n204544 );
or ( n258116 , n258114 , n258115 );
not ( n258117 , n242108 );
nand ( n258118 , n258117 , n204553 );
nand ( n258119 , n258116 , n258118 );
and ( n258120 , n258119 , n27878 );
not ( n258121 , n258119 );
and ( n258122 , n258121 , n27870 );
nor ( n258123 , n258120 , n258122 );
nand ( n258124 , n258113 , n258123 );
and ( n258125 , n258124 , n240510 );
not ( n258126 , n258124 );
not ( n258127 , n240510 );
and ( n258128 , n258126 , n258127 );
nor ( n258129 , n258125 , n258128 );
or ( n258130 , n258129 , n256376 );
nand ( n258131 , n258101 , n258130 );
buf ( n258132 , n258131 );
not ( n258133 , RI19ac12b0_2321);
or ( n258134 , n25328 , n258133 );
or ( n258135 , n25336 , n248823 );
nand ( n258136 , n258134 , n258135 );
buf ( n258137 , n258136 );
not ( n258138 , n28354 );
not ( n258139 , n257764 );
or ( n258140 , n258138 , n258139 );
not ( n258141 , n226551 );
not ( n258142 , n239220 );
or ( n258143 , n258141 , n258142 );
not ( n258144 , n226551 );
nand ( n258145 , n258144 , n239228 );
nand ( n258146 , n258143 , n258145 );
and ( n258147 , n258146 , n250580 );
not ( n258148 , n258146 );
and ( n258149 , n258148 , n250577 );
nor ( n258150 , n258147 , n258149 );
not ( n258151 , n258150 );
not ( n258152 , n244336 );
not ( n258153 , n258152 );
not ( n258154 , n258153 );
not ( n258155 , n233853 );
not ( n258156 , n244273 );
or ( n258157 , n258155 , n258156 );
nand ( n258158 , n244282 , n233854 );
nand ( n258159 , n258157 , n258158 );
not ( n258160 , n258159 );
or ( n258161 , n258154 , n258160 );
or ( n258162 , n258159 , n258153 );
nand ( n258163 , n258161 , n258162 );
nand ( n258164 , n258151 , n258163 );
not ( n258165 , n237256 );
not ( n258166 , n253080 );
or ( n258167 , n258165 , n258166 );
or ( n258168 , n257658 , n237256 );
nand ( n258169 , n258167 , n258168 );
and ( n258170 , n258169 , n249207 );
not ( n258171 , n258169 );
and ( n258172 , n258171 , n249208 );
nor ( n258173 , n258170 , n258172 );
not ( n258174 , n258173 );
and ( n258175 , n258164 , n258174 );
not ( n258176 , n258164 );
and ( n258177 , n258176 , n258173 );
nor ( n258178 , n258175 , n258177 );
buf ( n258179 , n236795 );
or ( n258180 , n258178 , n258179 );
nand ( n258181 , n258140 , n258180 );
buf ( n258182 , n258181 );
not ( n258183 , RI1754be18_19);
or ( n258184 , n255977 , n258183 );
not ( n258185 , n226822 );
nand ( n258186 , n258185 , n29281 );
nand ( n258187 , n258184 , n258186 );
buf ( n258188 , n258187 );
not ( n258189 , RI19a98630_2623);
or ( n258190 , n25328 , n258189 );
not ( n258191 , RI19a8e478_2695);
or ( n258192 , n25335 , n258191 );
nand ( n258193 , n258190 , n258192 );
buf ( n258194 , n258193 );
buf ( n258195 , n245455 );
not ( n258196 , n258195 );
not ( n258197 , n241962 );
or ( n258198 , n258196 , n258197 );
or ( n258199 , n241962 , n258195 );
nand ( n258200 , n258198 , n258199 );
not ( n258201 , n258200 );
not ( n258202 , n250501 );
and ( n258203 , n258201 , n258202 );
and ( n258204 , n258200 , n250501 );
nor ( n258205 , n258203 , n258204 );
not ( n258206 , n258179 );
nand ( n258207 , n258205 , n258206 );
not ( n258208 , n256883 );
nand ( n258209 , n258208 , n256910 );
or ( n258210 , n258207 , n258209 );
nor ( n258211 , n258205 , n226004 );
nand ( n258212 , n258211 , n258209 );
buf ( n258213 , n35431 );
nand ( n258214 , n258213 , n32734 );
nand ( n258215 , n258210 , n258212 , n258214 );
buf ( n258216 , n258215 );
not ( n258217 , n255440 );
not ( n258218 , n33246 );
or ( n258219 , n258217 , n258218 );
not ( n258220 , n255440 );
nand ( n258221 , n258220 , n253530 );
nand ( n258222 , n258219 , n258221 );
and ( n258223 , n258222 , n253536 );
not ( n258224 , n258222 );
and ( n258225 , n258224 , n253533 );
nor ( n258226 , n258223 , n258225 );
buf ( n258227 , n248037 );
not ( n258228 , n258227 );
not ( n258229 , n238792 );
or ( n258230 , n258228 , n258229 );
or ( n258231 , n238792 , n258227 );
nand ( n258232 , n258230 , n258231 );
buf ( n258233 , n246077 );
and ( n258234 , n258232 , n258233 );
not ( n258235 , n258232 );
and ( n258236 , n258235 , n238895 );
nor ( n258237 , n258234 , n258236 );
nor ( n258238 , n251709 , n258226 , n258237 );
not ( n258239 , n258238 );
nor ( n258240 , n251633 , n235050 );
nand ( n258241 , n258240 , n258226 );
not ( n258242 , n258226 );
nor ( n258243 , n258242 , n234818 );
nand ( n258244 , n258243 , n258237 );
nand ( n258245 , n256673 , n236140 );
nand ( n258246 , n258239 , n258241 , n258244 , n258245 );
buf ( n258247 , n258246 );
not ( n258248 , n248248 );
not ( n258249 , n240312 );
or ( n258250 , n258248 , n258249 );
not ( n258251 , n248248 );
nand ( n258252 , n258251 , n240316 );
nand ( n258253 , n258250 , n258252 );
xor ( n258254 , n258253 , n240508 );
not ( n258255 , n246065 );
not ( n258256 , n243783 );
not ( n258257 , n236762 );
not ( n258258 , n258257 );
or ( n258259 , n258256 , n258258 );
nand ( n258260 , n236762 , n243782 );
nand ( n258261 , n258259 , n258260 );
not ( n258262 , n258261 );
or ( n258263 , n258255 , n258262 );
or ( n258264 , n258261 , n246065 );
nand ( n258265 , n258263 , n258264 );
not ( n258266 , n258265 );
nand ( n258267 , n258254 , n258266 );
or ( n258268 , n253394 , n258267 );
not ( n258269 , n258266 );
not ( n258270 , n253392 );
or ( n258271 , n258269 , n258270 );
nor ( n258272 , n258254 , n235050 );
nand ( n258273 , n258271 , n258272 );
nand ( n258274 , n31577 , n207930 );
nand ( n258275 , n258268 , n258273 , n258274 );
buf ( n258276 , n258275 );
not ( n258277 , n258254 );
nand ( n258278 , n258277 , n253400 );
or ( n258279 , n253398 , n258278 );
buf ( n258280 , n43517 );
nor ( n258281 , n253379 , n258280 );
nand ( n258282 , n258281 , n258278 );
nand ( n258283 , n255116 , n25437 );
nand ( n258284 , n258279 , n258282 , n258283 );
buf ( n258285 , n258284 );
not ( n258286 , n34513 );
not ( n258287 , n245702 );
or ( n258288 , n258286 , n258287 );
not ( n258289 , n50354 );
not ( n258290 , n53811 );
or ( n258291 , n258289 , n258290 );
not ( n258292 , n50354 );
nand ( n258293 , n258292 , n53820 );
nand ( n258294 , n258291 , n258293 );
and ( n258295 , n258294 , n231776 );
not ( n258296 , n258294 );
and ( n258297 , n258296 , n253730 );
nor ( n258298 , n258295 , n258297 );
not ( n258299 , n45180 );
not ( n258300 , n244054 );
or ( n258301 , n258299 , n258300 );
not ( n258302 , n45180 );
nand ( n258303 , n258302 , n253557 );
nand ( n258304 , n258301 , n258303 );
and ( n258305 , n258304 , n245517 );
not ( n258306 , n258304 );
and ( n258307 , n258306 , n253560 );
nor ( n258308 , n258305 , n258307 );
nand ( n258309 , n258298 , n258308 );
not ( n258310 , n46888 );
not ( n258311 , n250019 );
or ( n258312 , n258310 , n258311 );
not ( n258313 , n46888 );
nand ( n258314 , n258313 , n250028 );
nand ( n258315 , n258312 , n258314 );
buf ( n258316 , n252823 );
and ( n258317 , n258315 , n258316 );
not ( n258318 , n258315 );
buf ( n258319 , n252831 );
and ( n258320 , n258318 , n258319 );
nor ( n258321 , n258317 , n258320 );
not ( n258322 , n258321 );
and ( n258323 , n258309 , n258322 );
not ( n258324 , n258309 );
and ( n258325 , n258324 , n258321 );
nor ( n258326 , n258323 , n258325 );
buf ( n258327 , n37724 );
buf ( n258328 , n258327 );
or ( n258329 , n258326 , n258328 );
nand ( n258330 , n258288 , n258329 );
buf ( n258331 , n258330 );
not ( n258332 , n246374 );
not ( n258333 , n44539 );
or ( n258334 , n258332 , n258333 );
or ( n258335 , n44539 , n246374 );
nand ( n258336 , n258334 , n258335 );
and ( n258337 , n258336 , n222525 );
not ( n258338 , n258336 );
and ( n258339 , n258338 , n44761 );
nor ( n258340 , n258337 , n258339 );
nand ( n258341 , n258340 , n233973 );
not ( n258342 , n248921 );
not ( n258343 , n250098 );
or ( n258344 , n258342 , n258343 );
not ( n258345 , n248921 );
nand ( n258346 , n258345 , n250099 );
nand ( n258347 , n258344 , n258346 );
and ( n258348 , n258347 , n250108 );
not ( n258349 , n258347 );
and ( n258350 , n258349 , n250105 );
nor ( n258351 , n258348 , n258350 );
not ( n258352 , n247733 );
not ( n258353 , n238164 );
not ( n258354 , n45727 );
or ( n258355 , n258353 , n258354 );
not ( n258356 , n238164 );
nand ( n258357 , n258356 , n247727 );
nand ( n258358 , n258355 , n258357 );
not ( n258359 , n258358 );
or ( n258360 , n258352 , n258359 );
or ( n258361 , n258358 , n247733 );
nand ( n258362 , n258360 , n258361 );
not ( n258363 , n258362 );
nand ( n258364 , n258351 , n258363 );
or ( n258365 , n258341 , n258364 );
not ( n258366 , n258363 );
not ( n258367 , n258340 );
or ( n258368 , n258366 , n258367 );
not ( n258369 , n222532 );
nor ( n258370 , n258351 , n258369 );
nand ( n258371 , n258368 , n258370 );
nand ( n258372 , n31577 , n30122 );
nand ( n258373 , n258365 , n258371 , n258372 );
buf ( n258374 , n258373 );
not ( n258375 , n255774 );
not ( n258376 , n246548 );
or ( n258377 , n258375 , n258376 );
not ( n258378 , n255774 );
nand ( n258379 , n258378 , n246553 );
nand ( n258380 , n258377 , n258379 );
and ( n258381 , n258380 , n246654 );
not ( n258382 , n258380 );
and ( n258383 , n258382 , n246661 );
nor ( n258384 , n258381 , n258383 );
nand ( n258385 , n258384 , n253565 );
not ( n258386 , n27862 );
not ( n258387 , n228364 );
or ( n258388 , n258386 , n258387 );
not ( n258389 , n27862 );
nand ( n258390 , n258389 , n50539 );
nand ( n258391 , n258388 , n258390 );
and ( n258392 , n258391 , n55726 );
not ( n258393 , n258391 );
and ( n258394 , n258393 , n55727 );
nor ( n258395 , n258392 , n258394 );
not ( n258396 , n258395 );
not ( n258397 , n237833 );
not ( n258398 , n254916 );
or ( n258399 , n258397 , n258398 );
not ( n258400 , n237833 );
nand ( n258401 , n258400 , n251684 );
nand ( n258402 , n258399 , n258401 );
and ( n258403 , n258402 , n251692 );
not ( n258404 , n258402 );
and ( n258405 , n258404 , n251693 );
nor ( n258406 , n258403 , n258405 );
not ( n258407 , n258406 );
nand ( n258408 , n258396 , n258407 );
or ( n258409 , n258385 , n258408 );
not ( n258410 , n258407 );
not ( n258411 , n258384 );
or ( n258412 , n258410 , n258411 );
nor ( n258413 , n258396 , n37725 );
nand ( n258414 , n258412 , n258413 );
nand ( n258415 , n31577 , n205344 );
nand ( n258416 , n258409 , n258414 , n258415 );
buf ( n258417 , n258416 );
nand ( n258418 , n245801 , n245932 );
nor ( n258419 , n226001 , n256413 );
not ( n258420 , n258419 );
or ( n258421 , n258418 , n258420 );
nand ( n258422 , n48244 , n258418 );
nand ( n258423 , n234453 , n33423 );
nand ( n258424 , n258421 , n258422 , n258423 );
buf ( n258425 , n258424 );
not ( n258426 , n248069 );
not ( n258427 , n258426 );
not ( n258428 , n248083 );
or ( n258429 , n258427 , n258428 );
nand ( n258430 , n258429 , n226010 );
not ( n258431 , n248524 );
not ( n258432 , n243659 );
or ( n258433 , n258431 , n258432 );
or ( n258434 , n243659 , n248524 );
nand ( n258435 , n258433 , n258434 );
and ( n258436 , n258435 , n251846 );
not ( n258437 , n258435 );
and ( n258438 , n258437 , n251856 );
nor ( n258439 , n258436 , n258438 );
or ( n258440 , n258430 , n258439 );
nor ( n258441 , n248069 , n249030 );
nand ( n258442 , n258441 , n248083 , n258439 );
nand ( n258443 , n239240 , n38457 );
nand ( n258444 , n258440 , n258442 , n258443 );
buf ( n258445 , n258444 );
not ( n258446 , n239157 );
not ( n258447 , n244386 );
or ( n258448 , n258446 , n258447 );
or ( n258449 , n244386 , n239157 );
nand ( n258450 , n258448 , n258449 );
not ( n258451 , n258450 );
not ( n258452 , n240153 );
and ( n258453 , n258451 , n258452 );
and ( n258454 , n258450 , n255353 );
nor ( n258455 , n258453 , n258454 );
nor ( n258456 , n258455 , n240080 );
not ( n258457 , n246059 );
not ( n258458 , n45026 );
or ( n258459 , n258457 , n258458 );
not ( n258460 , n246059 );
nand ( n258461 , n258460 , n45023 );
nand ( n258462 , n258459 , n258461 );
and ( n258463 , n258462 , n223016 );
not ( n258464 , n258462 );
and ( n258465 , n258464 , n45261 );
nor ( n258466 , n258463 , n258465 );
not ( n258467 , n249371 );
nand ( n258468 , n258467 , n248663 );
not ( n258469 , n258468 );
not ( n258470 , n249372 );
not ( n258471 , n258470 );
and ( n258472 , n258469 , n258471 );
and ( n258473 , n258468 , n258470 );
nor ( n258474 , n258472 , n258473 );
not ( n258475 , n250151 );
nand ( n258476 , n258475 , n248640 );
not ( n258477 , n258476 );
not ( n258478 , n243171 );
and ( n258479 , n258477 , n258478 );
and ( n258480 , n258476 , n243171 );
nor ( n258481 , n258479 , n258480 );
not ( n258482 , n258481 );
not ( n258483 , n258482 );
not ( n258484 , n250934 );
not ( n258485 , n258484 );
or ( n258486 , n258483 , n258485 );
nand ( n258487 , n250934 , n258481 );
nand ( n258488 , n258486 , n258487 );
xor ( n258489 , n258474 , n258488 );
nand ( n258490 , n248581 , n251835 );
and ( n258491 , n258490 , n243017 );
not ( n258492 , n258490 );
not ( n258493 , n243017 );
and ( n258494 , n258492 , n258493 );
nor ( n258495 , n258491 , n258494 );
not ( n258496 , n258495 );
nand ( n258497 , n248596 , n250214 );
and ( n258498 , n258497 , n243052 );
not ( n258499 , n258497 );
and ( n258500 , n258499 , n243053 );
nor ( n258501 , n258498 , n258500 );
not ( n258502 , n258501 );
not ( n258503 , n258502 );
or ( n258504 , n258496 , n258503 );
not ( n258505 , n258490 );
not ( n258506 , n258493 );
and ( n258507 , n258505 , n258506 );
and ( n258508 , n258490 , n258493 );
nor ( n258509 , n258507 , n258508 );
nand ( n258510 , n258501 , n258509 );
nand ( n258511 , n258504 , n258510 );
xor ( n258512 , n258489 , n258511 );
not ( n258513 , n243566 );
not ( n258514 , n254728 );
and ( n258515 , n258513 , n258514 );
not ( n258516 , n258513 );
not ( n258517 , n255100 );
and ( n258518 , n258516 , n258517 );
nor ( n258519 , n258515 , n258518 );
and ( n258520 , n258512 , n258519 );
not ( n258521 , n258512 );
not ( n258522 , n258519 );
and ( n258523 , n258521 , n258522 );
nor ( n258524 , n258520 , n258523 );
nor ( n258525 , n258466 , n258524 );
nand ( n258526 , n258456 , n258525 );
not ( n258527 , n258524 );
not ( n258528 , n258527 );
not ( n258529 , n258455 );
not ( n258530 , n258529 );
or ( n258531 , n258528 , n258530 );
not ( n258532 , n258466 );
nor ( n258533 , n258532 , n252200 );
nand ( n258534 , n258531 , n258533 );
nand ( n258535 , n244987 , n29983 );
nand ( n258536 , n258526 , n258534 , n258535 );
buf ( n258537 , n258536 );
not ( n258538 , n237604 );
not ( n258539 , n258538 );
not ( n258540 , n233987 );
or ( n258541 , n258539 , n258540 );
or ( n258542 , n233987 , n258538 );
nand ( n258543 , n258541 , n258542 );
and ( n258544 , n258543 , n253206 );
not ( n258545 , n258543 );
and ( n258546 , n258545 , n233990 );
nor ( n258547 , n258544 , n258546 );
not ( n258548 , n258547 );
nor ( n258549 , n258548 , n244399 );
buf ( n258550 , n237985 );
not ( n258551 , n258550 );
not ( n258552 , n257110 );
not ( n258553 , n258552 );
or ( n258554 , n258551 , n258553 );
or ( n258555 , n226319 , n258550 );
nand ( n258556 , n258554 , n258555 );
not ( n258557 , n257116 );
and ( n258558 , n258556 , n258557 );
not ( n258559 , n258556 );
not ( n258560 , n257113 );
and ( n258561 , n258559 , n258560 );
nor ( n258562 , n258558 , n258561 );
not ( n258563 , n230428 );
not ( n258564 , n230443 );
nand ( n258565 , n258564 , n40261 );
not ( n258566 , n258565 );
not ( n258567 , n235828 );
and ( n258568 , n258566 , n258567 );
and ( n258569 , n258565 , n235828 );
nor ( n258570 , n258568 , n258569 );
not ( n258571 , n258570 );
nand ( n258572 , n52649 , n52663 );
and ( n258573 , n258572 , n40246 );
not ( n258574 , n258572 );
and ( n258575 , n258574 , n235819 );
nor ( n258576 , n258573 , n258575 );
not ( n258577 , n258576 );
or ( n258578 , n258571 , n258577 );
or ( n258579 , n258570 , n258576 );
nand ( n258580 , n258578 , n258579 );
nand ( n258581 , n40315 , n230387 );
not ( n258582 , n258581 );
not ( n258583 , n235841 );
and ( n258584 , n258582 , n258583 );
and ( n258585 , n258581 , n235841 );
nor ( n258586 , n258584 , n258585 );
and ( n258587 , n258580 , n258586 );
not ( n258588 , n258580 );
not ( n258589 , n258586 );
and ( n258590 , n258588 , n258589 );
nor ( n258591 , n258587 , n258590 );
nand ( n258592 , n40349 , n52709 );
not ( n258593 , n258592 );
not ( n258594 , n235863 );
and ( n258595 , n258593 , n258594 );
and ( n258596 , n258592 , n235863 );
nor ( n258597 , n258595 , n258596 );
not ( n258598 , n258597 );
nand ( n258599 , n52742 , n230488 );
not ( n258600 , n258599 );
not ( n258601 , n258600 );
not ( n258602 , n40416 );
or ( n258603 , n258601 , n258602 );
nand ( n258604 , n235855 , n258599 );
nand ( n258605 , n258603 , n258604 );
not ( n258606 , n258605 );
or ( n258607 , n258598 , n258606 );
or ( n258608 , n258605 , n258597 );
nand ( n258609 , n258607 , n258608 );
xor ( n258610 , n258591 , n258609 );
not ( n258611 , n258610 );
not ( n258612 , n258611 );
not ( n258613 , n258612 );
or ( n258614 , n258563 , n258613 );
not ( n258615 , n230428 );
nand ( n258616 , n258615 , n258611 );
nand ( n258617 , n258614 , n258616 );
buf ( n258618 , n242520 );
and ( n258619 , n258617 , n258618 );
not ( n258620 , n258617 );
not ( n258621 , n242527 );
not ( n258622 , n258621 );
and ( n258623 , n258620 , n258622 );
nor ( n258624 , n258619 , n258623 );
nor ( n258625 , n258562 , n258624 );
nand ( n258626 , n258549 , n258625 );
not ( n258627 , n258562 );
not ( n258628 , n258627 );
not ( n258629 , n258547 );
or ( n258630 , n258628 , n258629 );
not ( n258631 , n258624 );
nor ( n258632 , n258631 , n226003 );
nand ( n258633 , n258630 , n258632 );
nand ( n258634 , n245943 , n211219 );
nand ( n258635 , n258626 , n258633 , n258634 );
buf ( n258636 , n258635 );
not ( n258637 , n222383 );
not ( n258638 , n237810 );
or ( n258639 , n258637 , n258638 );
not ( n258640 , n222383 );
nand ( n258641 , n258640 , n237817 );
nand ( n258642 , n258639 , n258641 );
xor ( n258643 , n258642 , n237868 );
not ( n258644 , n258643 );
not ( n258645 , n254539 );
nand ( n258646 , n258644 , n258645 );
or ( n258647 , n258646 , n254529 );
nor ( n258648 , n254527 , n219702 );
nand ( n258649 , n258648 , n258646 );
nand ( n258650 , n244987 , n215143 );
nand ( n258651 , n258647 , n258649 , n258650 );
buf ( n258652 , n258651 );
not ( n258653 , RI19abba90_2370);
or ( n258654 , n25335 , n258653 );
not ( n258655 , n229127 );
nand ( n258656 , n258655 , RI1754b350_42);
nor ( n258657 , n249124 , n51364 );
and ( n258658 , n51363 , n258657 );
nor ( n258659 , RI1754a630_70 , RI1754a5b8_71);
nand ( n258660 , n258658 , n258659 );
nand ( n258661 , n258654 , n258656 , n258660 );
buf ( n258662 , n258661 );
not ( n258663 , n257646 );
not ( n258664 , n258663 );
not ( n258665 , n252232 );
not ( n258666 , n246385 );
or ( n258667 , n258665 , n258666 );
not ( n258668 , n252232 );
nand ( n258669 , n258668 , n255822 );
nand ( n258670 , n258667 , n258669 );
and ( n258671 , n258670 , n246441 );
not ( n258672 , n258670 );
and ( n258673 , n258672 , n246449 );
nor ( n258674 , n258671 , n258673 );
not ( n258675 , n258674 );
not ( n258676 , n255497 );
not ( n258677 , n246787 );
not ( n258678 , n249927 );
or ( n258679 , n258677 , n258678 );
not ( n258680 , n246787 );
nand ( n258681 , n258680 , n255493 );
nand ( n258682 , n258679 , n258681 );
not ( n258683 , n258682 );
or ( n258684 , n258676 , n258683 );
or ( n258685 , n258682 , n255497 );
nand ( n258686 , n258684 , n258685 );
not ( n258687 , n258686 );
nand ( n258688 , n258675 , n258687 );
not ( n258689 , n258688 );
and ( n258690 , n258664 , n258689 );
and ( n258691 , n237714 , n37254 );
nor ( n258692 , n258690 , n258691 );
not ( n258693 , n257622 );
nand ( n258694 , n258693 , n258674 );
nand ( n258695 , n258674 , n245241 );
not ( n258696 , n258695 );
nand ( n258697 , n258696 , n258686 );
nand ( n258698 , n258692 , n258694 , n258697 );
buf ( n258699 , n258698 );
not ( n258700 , n238557 );
not ( n258701 , n241131 );
or ( n258702 , n258700 , n258701 );
or ( n258703 , n241131 , n238557 );
nand ( n258704 , n258702 , n258703 );
and ( n258705 , n258704 , n241180 );
not ( n258706 , n258704 );
and ( n258707 , n258706 , n241181 );
nor ( n258708 , n258705 , n258707 );
nor ( n258709 , n258708 , n249531 );
not ( n258710 , n258709 );
buf ( n258711 , n37698 );
not ( n258712 , n258711 );
not ( n258713 , n257724 );
or ( n258714 , n258712 , n258713 );
buf ( n258715 , n252443 );
or ( n258716 , n258715 , n258711 );
nand ( n258717 , n258714 , n258716 );
and ( n258718 , n258717 , n257729 );
not ( n258719 , n258717 );
not ( n258720 , n257729 );
and ( n258721 , n258719 , n258720 );
nor ( n258722 , n258718 , n258721 );
buf ( n258723 , n258722 );
not ( n258724 , n220863 );
not ( n258725 , n246671 );
or ( n258726 , n258724 , n258725 );
not ( n258727 , n220863 );
nand ( n258728 , n258727 , n244453 );
nand ( n258729 , n258726 , n258728 );
and ( n258730 , n258729 , n249789 );
not ( n258731 , n258729 );
and ( n258732 , n258731 , n249792 );
nor ( n258733 , n258730 , n258732 );
not ( n258734 , n258733 );
nand ( n258735 , n258723 , n258734 );
or ( n258736 , n258710 , n258735 );
not ( n258737 , n258734 );
not ( n258738 , n258708 );
not ( n258739 , n258738 );
or ( n258740 , n258737 , n258739 );
nor ( n258741 , n258723 , n40465 );
nand ( n258742 , n258740 , n258741 );
buf ( n258743 , n35431 );
nand ( n258744 , n258743 , n32226 );
nand ( n258745 , n258736 , n258742 , n258744 );
buf ( n258746 , n258745 );
buf ( n258747 , n33346 );
buf ( n258748 , n35978 );
buf ( n258749 , n205117 );
not ( n258750 , n38646 );
not ( n258751 , n252711 );
or ( n258752 , n258750 , n258751 );
nand ( n258753 , n253117 , n250694 );
not ( n258754 , n250725 );
and ( n258755 , n258753 , n258754 );
not ( n258756 , n258753 );
and ( n258757 , n258756 , n250725 );
nor ( n258758 , n258755 , n258757 );
buf ( n258759 , n253358 );
or ( n258760 , n258758 , n258759 );
nand ( n258761 , n258752 , n258760 );
buf ( n258762 , n258761 );
not ( n258763 , n254967 );
not ( n258764 , n258763 );
not ( n258765 , n236781 );
or ( n258766 , n258764 , n258765 );
or ( n258767 , n236781 , n258763 );
nand ( n258768 , n258766 , n258767 );
and ( n258769 , n258768 , n234889 );
not ( n258770 , n258768 );
and ( n258771 , n258770 , n236789 );
nor ( n258772 , n258769 , n258771 );
nand ( n258773 , n258772 , n205649 );
not ( n258774 , n258340 );
nand ( n258775 , n258774 , n258363 );
or ( n258776 , n258773 , n258775 );
not ( n258777 , n258774 );
not ( n258778 , n258772 );
or ( n258779 , n258777 , n258778 );
nor ( n258780 , n258363 , n52445 );
nand ( n258781 , n258779 , n258780 );
nand ( n258782 , n35431 , n49423 );
nand ( n258783 , n258776 , n258781 , n258782 );
buf ( n258784 , n258783 );
not ( n258785 , RI19ac0338_2330);
or ( n258786 , n25328 , n258785 );
not ( n258787 , RI19ab73c8_2400);
or ( n258788 , n226822 , n258787 );
nand ( n258789 , n258786 , n258788 );
buf ( n258790 , n258789 );
not ( n258791 , n38273 );
not ( n258792 , n234453 );
or ( n258793 , n258791 , n258792 );
buf ( n258794 , n52360 );
not ( n258795 , n258794 );
not ( n258796 , n256547 );
or ( n258797 , n258795 , n258796 );
or ( n258798 , n256547 , n258794 );
nand ( n258799 , n258797 , n258798 );
and ( n258800 , n258799 , n248067 );
not ( n258801 , n258799 );
and ( n258802 , n258801 , n248062 );
nor ( n258803 , n258800 , n258802 );
not ( n258804 , n244553 );
not ( n258805 , n239705 );
or ( n258806 , n258804 , n258805 );
not ( n258807 , n244553 );
nand ( n258808 , n258807 , n239715 );
nand ( n258809 , n258806 , n258808 );
not ( n258810 , n255625 );
and ( n258811 , n258809 , n258810 );
not ( n258812 , n258809 );
and ( n258813 , n258812 , n255625 );
nor ( n258814 , n258811 , n258813 );
nand ( n258815 , n258803 , n258814 );
buf ( n258816 , n244876 );
not ( n258817 , n258816 );
not ( n258818 , n231421 );
or ( n258819 , n258817 , n258818 );
or ( n258820 , n231421 , n258816 );
nand ( n258821 , n258819 , n258820 );
and ( n258822 , n258821 , n53665 );
not ( n258823 , n258821 );
and ( n258824 , n258823 , n53669 );
nor ( n258825 , n258822 , n258824 );
and ( n258826 , n258815 , n258825 );
not ( n258827 , n258815 );
not ( n258828 , n258825 );
and ( n258829 , n258827 , n258828 );
nor ( n258830 , n258826 , n258829 );
or ( n258831 , n258830 , n235052 );
nand ( n258832 , n258793 , n258831 );
buf ( n258833 , n258832 );
buf ( n258834 , n29850 );
or ( n258835 , n25328 , n235058 );
or ( n258836 , n25335 , n252206 );
nand ( n258837 , n258835 , n258836 );
buf ( n258838 , n258837 );
buf ( n258839 , n221492 );
buf ( n258840 , n25755 );
not ( n258841 , n28749 );
not ( n258842 , n37728 );
or ( n258843 , n258841 , n258842 );
not ( n258844 , n238288 );
not ( n258845 , n231480 );
not ( n258846 , n258845 );
and ( n258847 , n258844 , n258846 );
and ( n258848 , n238288 , n258845 );
nor ( n258849 , n258847 , n258848 );
and ( n258850 , n258849 , n238401 );
not ( n258851 , n258849 );
and ( n258852 , n258851 , n238409 );
nor ( n258853 , n258850 , n258852 );
not ( n258854 , n35494 );
not ( n258855 , n258854 );
not ( n258856 , n236881 );
or ( n258857 , n258855 , n258856 );
or ( n258858 , n236883 , n258854 );
nand ( n258859 , n258857 , n258858 );
not ( n258860 , n236993 );
and ( n258861 , n258859 , n258860 );
not ( n258862 , n258859 );
and ( n258863 , n258862 , n236993 );
nor ( n258864 , n258861 , n258863 );
nand ( n258865 , n258853 , n258864 );
not ( n258866 , n55863 );
not ( n258867 , n49181 );
or ( n258868 , n258866 , n258867 );
not ( n258869 , n55863 );
nand ( n258870 , n258869 , n49190 );
nand ( n258871 , n258868 , n258870 );
and ( n258872 , n258871 , n238183 );
not ( n258873 , n258871 );
and ( n258874 , n258873 , n238186 );
nor ( n258875 , n258872 , n258874 );
not ( n258876 , n258875 );
and ( n258877 , n258865 , n258876 );
not ( n258878 , n258865 );
and ( n258879 , n258878 , n258875 );
nor ( n258880 , n258877 , n258879 );
or ( n258881 , n258880 , n257851 );
nand ( n258882 , n258843 , n258881 );
buf ( n258883 , n258882 );
buf ( n258884 , n33209 );
not ( n258885 , n251160 );
nand ( n258886 , n258885 , n251173 );
not ( n258887 , n238866 );
not ( n258888 , n247500 );
or ( n258889 , n258887 , n258888 );
not ( n258890 , n238866 );
nand ( n258891 , n258890 , n247499 );
nand ( n258892 , n258889 , n258891 );
and ( n258893 , n258892 , n247553 );
not ( n258894 , n258892 );
and ( n258895 , n258894 , n247563 );
nor ( n258896 , n258893 , n258895 );
not ( n258897 , n258896 );
nor ( n258898 , n258897 , n252358 );
not ( n258899 , n258898 );
or ( n258900 , n258886 , n258899 );
nor ( n258901 , n258896 , n233971 );
nand ( n258902 , n258886 , n258901 );
nand ( n258903 , n231444 , n25941 );
nand ( n258904 , n258900 , n258902 , n258903 );
buf ( n258905 , n258904 );
not ( n258906 , RI19a95930_2643);
or ( n258907 , n25328 , n258906 );
not ( n258908 , RI19a8b700_2715);
or ( n258909 , n25335 , n258908 );
nand ( n258910 , n258907 , n258909 );
buf ( n258911 , n258910 );
not ( n258912 , RI19aa5560_2527);
or ( n258913 , n25328 , n258912 );
not ( n258914 , RI19a9bfd8_2598);
or ( n258915 , n226822 , n258914 );
nand ( n258916 , n258913 , n258915 );
buf ( n258917 , n258916 );
not ( n258918 , n226955 );
nand ( n258919 , n255828 , n258918 );
not ( n258920 , n45863 );
not ( n258921 , n258920 );
not ( n258922 , n36729 );
or ( n258923 , n258921 , n258922 );
not ( n258924 , n258920 );
nand ( n258925 , n258924 , n249482 );
nand ( n258926 , n258923 , n258925 );
and ( n258927 , n258926 , n249495 );
not ( n258928 , n258926 );
and ( n258929 , n258928 , n249491 );
nor ( n258930 , n258927 , n258929 );
not ( n258931 , n48355 );
not ( n258932 , n254947 );
or ( n258933 , n258931 , n258932 );
not ( n258934 , n48355 );
nand ( n258935 , n258934 , n254946 );
nand ( n258936 , n258933 , n258935 );
not ( n258937 , n254974 );
and ( n258938 , n258936 , n258937 );
not ( n258939 , n258936 );
and ( n258940 , n258939 , n254974 );
nor ( n258941 , n258938 , n258940 );
not ( n258942 , n258941 );
nand ( n258943 , n258930 , n258942 );
or ( n258944 , n258919 , n258943 );
not ( n258945 , n258942 );
not ( n258946 , n255828 );
or ( n258947 , n258945 , n258946 );
nor ( n258948 , n258930 , n53680 );
nand ( n258949 , n258947 , n258948 );
nand ( n258950 , n39767 , n32258 );
nand ( n258951 , n258944 , n258949 , n258950 );
buf ( n258952 , n258951 );
not ( n258953 , n234174 );
not ( n258954 , n251619 );
or ( n258955 , n258953 , n258954 );
not ( n258956 , n234174 );
nand ( n258957 , n258956 , n251627 );
nand ( n258958 , n258955 , n258957 );
and ( n258959 , n258958 , n251573 );
not ( n258960 , n258958 );
buf ( n258961 , n239994 );
and ( n258962 , n258960 , n258961 );
nor ( n258963 , n258959 , n258962 );
nor ( n258964 , n258963 , n253904 );
not ( n258965 , n258964 );
not ( n258966 , n44529 );
not ( n258967 , n241360 );
or ( n258968 , n258966 , n258967 );
not ( n258969 , n44529 );
nand ( n258970 , n258969 , n241369 );
nand ( n258971 , n258968 , n258970 );
buf ( n258972 , n237817 );
and ( n258973 , n258971 , n258972 );
not ( n258974 , n258971 );
buf ( n258975 , n237810 );
and ( n258976 , n258974 , n258975 );
nor ( n258977 , n258973 , n258976 );
not ( n258978 , n239679 );
not ( n258979 , n238975 );
or ( n258980 , n258978 , n258979 );
not ( n258981 , n239679 );
nand ( n258982 , n258981 , n238985 );
nand ( n258983 , n258980 , n258982 );
and ( n258984 , n258983 , n239108 );
not ( n258985 , n258983 );
and ( n258986 , n258985 , n239100 );
nor ( n258987 , n258984 , n258986 );
nand ( n258988 , n258977 , n258987 );
or ( n258989 , n258965 , n258988 );
not ( n258990 , n258963 );
not ( n258991 , n258990 );
not ( n258992 , n258977 );
or ( n258993 , n258991 , n258992 );
nor ( n258994 , n258987 , n55104 );
nand ( n258995 , n258993 , n258994 );
nand ( n258996 , n31577 , n32628 );
nand ( n258997 , n258989 , n258995 , n258996 );
buf ( n258998 , n258997 );
not ( n258999 , n252395 );
not ( n259000 , n258999 );
not ( n259001 , n257952 );
or ( n259002 , n259000 , n259001 );
or ( n259003 , n257952 , n258999 );
nand ( n259004 , n259002 , n259003 );
and ( n259005 , n259004 , n257964 );
not ( n259006 , n259004 );
and ( n259007 , n259006 , n257963 );
nor ( n259008 , n259005 , n259007 );
not ( n259009 , n39763 );
nand ( n259010 , n259008 , n259009 );
not ( n259011 , n35401 );
not ( n259012 , n223951 );
or ( n259013 , n259011 , n259012 );
or ( n259014 , n255071 , n35401 );
nand ( n259015 , n259013 , n259014 );
and ( n259016 , n259015 , n46420 );
not ( n259017 , n259015 );
not ( n259018 , n257541 );
and ( n259019 , n259017 , n259018 );
nor ( n259020 , n259016 , n259019 );
not ( n259021 , n259020 );
not ( n259022 , n246819 );
not ( n259023 , n249927 );
or ( n259024 , n259022 , n259023 );
not ( n259025 , n246819 );
nand ( n259026 , n259025 , n255493 );
nand ( n259027 , n259024 , n259026 );
and ( n259028 , n259027 , n255497 );
not ( n259029 , n259027 );
and ( n259030 , n259029 , n255500 );
nor ( n259031 , n259028 , n259030 );
nand ( n259032 , n259021 , n259031 );
or ( n259033 , n259010 , n259032 );
nor ( n259034 , n259008 , n247212 );
nand ( n259035 , n259034 , n259032 );
nand ( n259036 , n238114 , n207340 );
nand ( n259037 , n259033 , n259035 , n259036 );
buf ( n259038 , n259037 );
buf ( n259039 , n32398 );
buf ( n259040 , n55653 );
not ( n259041 , RI19ac96e0_2259);
or ( n259042 , n25328 , n259041 );
or ( n259043 , n226822 , n249038 );
nand ( n259044 , n259042 , n259043 );
buf ( n259045 , n259044 );
not ( n259046 , n30266 );
not ( n259047 , n245701 );
or ( n259048 , n259046 , n259047 );
not ( n259049 , n54459 );
not ( n259050 , n251162 );
or ( n259051 , n259049 , n259050 );
not ( n259052 , n54459 );
nand ( n259053 , n259052 , n245473 );
nand ( n259054 , n259051 , n259053 );
and ( n259055 , n259054 , n251168 );
not ( n259056 , n259054 );
and ( n259057 , n259056 , n251171 );
nor ( n259058 , n259055 , n259057 );
not ( n259059 , n259058 );
not ( n259060 , n50530 );
not ( n259061 , n35804 );
or ( n259062 , n259060 , n259061 );
not ( n259063 , n50530 );
nand ( n259064 , n259063 , n35811 );
nand ( n259065 , n259062 , n259064 );
and ( n259066 , n259065 , n253336 );
not ( n259067 , n259065 );
and ( n259068 , n259067 , n257757 );
nor ( n259069 , n259066 , n259068 );
nand ( n259070 , n259059 , n259069 );
not ( n259071 , n235709 );
not ( n259072 , n259071 );
not ( n259073 , n238461 );
or ( n259074 , n259072 , n259073 );
nand ( n259075 , n238470 , n235709 );
nand ( n259076 , n259074 , n259075 );
not ( n259077 , n259076 );
buf ( n259078 , n32472 );
not ( n259079 , n259078 );
and ( n259080 , n259077 , n259079 );
and ( n259081 , n259076 , n259078 );
nor ( n259082 , n259080 , n259081 );
not ( n259083 , n259082 );
and ( n259084 , n259070 , n259083 );
not ( n259085 , n259070 );
and ( n259086 , n259085 , n259082 );
nor ( n259087 , n259084 , n259086 );
or ( n259088 , n259087 , n254882 );
nand ( n259089 , n259048 , n259088 );
buf ( n259090 , n259089 );
buf ( n259091 , n235536 );
not ( n259092 , n259091 );
not ( n259093 , n248135 );
or ( n259094 , n259092 , n259093 );
or ( n259095 , n248135 , n259091 );
nand ( n259096 , n259094 , n259095 );
and ( n259097 , n259096 , n248149 );
not ( n259098 , n259096 );
and ( n259099 , n259098 , n248146 );
nor ( n259100 , n259097 , n259099 );
not ( n259101 , n259100 );
nand ( n259102 , n259101 , n235051 );
buf ( n259103 , n234279 );
not ( n259104 , n259103 );
buf ( n259105 , n43722 );
not ( n259106 , n259105 );
or ( n259107 , n259104 , n259106 );
or ( n259108 , n259105 , n259103 );
nand ( n259109 , n259107 , n259108 );
and ( n259110 , n259109 , n43956 );
not ( n259111 , n259109 );
and ( n259112 , n259111 , n43964 );
nor ( n259113 , n259110 , n259112 );
not ( n259114 , n239373 );
not ( n259115 , n259114 );
not ( n259116 , n258055 );
or ( n259117 , n259115 , n259116 );
or ( n259118 , n258055 , n259114 );
nand ( n259119 , n259117 , n259118 );
and ( n259120 , n259119 , n258061 );
not ( n259121 , n259119 );
and ( n259122 , n259121 , n258058 );
nor ( n259123 , n259120 , n259122 );
not ( n259124 , n259123 );
nand ( n259125 , n259113 , n259124 );
or ( n259126 , n259102 , n259125 );
not ( n259127 , n259113 );
not ( n259128 , n259101 );
or ( n259129 , n259127 , n259128 );
nor ( n259130 , n259124 , n33253 );
nand ( n259131 , n259129 , n259130 );
nand ( n259132 , n237361 , n209207 );
nand ( n259133 , n259126 , n259131 , n259132 );
buf ( n259134 , n259133 );
or ( n259135 , n233507 , n255659 );
not ( n259136 , RI19ac6620_2282);
or ( n259137 , n25335 , n259136 );
nand ( n259138 , n259135 , n259137 );
buf ( n259139 , n259138 );
not ( n259140 , RI19aac6d0_2480);
or ( n259141 , n233507 , n259140 );
not ( n259142 , RI19aa2068_2552);
or ( n259143 , n25335 , n259142 );
nand ( n259144 , n259141 , n259143 );
buf ( n259145 , n259144 );
not ( n259146 , n258495 );
not ( n259147 , n250229 );
or ( n259148 , n259146 , n259147 );
not ( n259149 , n258495 );
not ( n259150 , n250229 );
nand ( n259151 , n259149 , n259150 );
nand ( n259152 , n259148 , n259151 );
buf ( n259153 , n228042 );
and ( n259154 , n259152 , n259153 );
not ( n259155 , n259152 );
and ( n259156 , n259155 , n250942 );
nor ( n259157 , n259154 , n259156 );
not ( n259158 , n259157 );
nand ( n259159 , n259158 , n256197 );
buf ( n259160 , n254337 );
not ( n259161 , n259160 );
not ( n259162 , n238279 );
not ( n259163 , n259162 );
not ( n259164 , n236166 );
or ( n259165 , n259163 , n259164 );
or ( n259166 , n254275 , n259162 );
nand ( n259167 , n259165 , n259166 );
not ( n259168 , n259167 );
not ( n259169 , n259168 );
or ( n259170 , n259161 , n259169 );
not ( n259171 , n254344 );
not ( n259172 , n259171 );
nand ( n259173 , n259172 , n259167 );
nand ( n259174 , n259170 , n259173 );
nand ( n259175 , n259174 , n239934 );
or ( n259176 , n259159 , n259175 );
not ( n259177 , n259174 );
not ( n259178 , n259158 );
or ( n259179 , n259177 , n259178 );
nor ( n259180 , n256197 , n46425 );
nand ( n259181 , n259179 , n259180 );
nand ( n259182 , n253486 , n35756 );
nand ( n259183 , n259176 , n259181 , n259182 );
buf ( n259184 , n259183 );
not ( n259185 , n253904 );
not ( n259186 , n239687 );
not ( n259187 , n238975 );
or ( n259188 , n259186 , n259187 );
not ( n259189 , n239687 );
nand ( n259190 , n259189 , n238985 );
nand ( n259191 , n259188 , n259190 );
and ( n259192 , n259191 , n239100 );
not ( n259193 , n259191 );
and ( n259194 , n259193 , n239108 );
nor ( n259195 , n259192 , n259194 );
nand ( n259196 , n259185 , n259195 );
not ( n259197 , n243649 );
not ( n259198 , n259197 );
not ( n259199 , n255100 );
or ( n259200 , n259198 , n259199 );
or ( n259201 , n258514 , n259197 );
nand ( n259202 , n259200 , n259201 );
not ( n259203 , n258511 );
and ( n259204 , n258488 , n258474 );
not ( n259205 , n258488 );
not ( n259206 , n258474 );
and ( n259207 , n259205 , n259206 );
nor ( n259208 , n259204 , n259207 );
not ( n259209 , n259208 );
or ( n259210 , n259203 , n259209 );
not ( n259211 , n258511 );
not ( n259212 , n259208 );
nand ( n259213 , n259211 , n259212 );
nand ( n259214 , n259210 , n259213 );
buf ( n259215 , n259214 );
and ( n259216 , n259202 , n259215 );
not ( n259217 , n259202 );
buf ( n259218 , n258512 );
and ( n259219 , n259217 , n259218 );
nor ( n259220 , n259216 , n259219 );
not ( n259221 , n259220 );
not ( n259222 , n237072 );
not ( n259223 , n253072 );
or ( n259224 , n259222 , n259223 );
nand ( n259225 , n253073 , n237076 );
nand ( n259226 , n259224 , n259225 );
and ( n259227 , n259226 , n257659 );
not ( n259228 , n259226 );
and ( n259229 , n259228 , n253081 );
nor ( n259230 , n259227 , n259229 );
nand ( n259231 , n259221 , n259230 );
or ( n259232 , n259196 , n259231 );
not ( n259233 , n259221 );
not ( n259234 , n259195 );
or ( n259235 , n259233 , n259234 );
nor ( n259236 , n259230 , n37725 );
nand ( n259237 , n259235 , n259236 );
nand ( n259238 , n236798 , n204612 );
nand ( n259239 , n259232 , n259237 , n259238 );
buf ( n259240 , n259239 );
not ( n259241 , RI19aab0c8_2488);
or ( n259242 , n233507 , n259241 );
not ( n259243 , RI19aa10f0_2560);
or ( n259244 , n25335 , n259243 );
nand ( n259245 , n259242 , n259244 );
buf ( n259246 , n259245 );
buf ( n259247 , n31379 );
buf ( n259248 , n38871 );
buf ( n259249 , n40002 );
buf ( n259250 , n40162 );
not ( n259251 , n237217 );
not ( n259252 , n249204 );
or ( n259253 , n259251 , n259252 );
or ( n259254 , n249204 , n237217 );
nand ( n259255 , n259253 , n259254 );
xor ( n259256 , n259255 , n249207 );
not ( n259257 , n239020 );
not ( n259258 , n52221 );
or ( n259259 , n259257 , n259258 );
not ( n259260 , n239020 );
nand ( n259261 , n259260 , n52229 );
nand ( n259262 , n259259 , n259261 );
not ( n259263 , n246385 );
not ( n259264 , n259263 );
and ( n259265 , n259262 , n259264 );
not ( n259266 , n259262 );
and ( n259267 , n259266 , n246389 );
nor ( n259268 , n259265 , n259267 );
not ( n259269 , n259268 );
nand ( n259270 , n259256 , n259269 );
not ( n259271 , n39588 );
not ( n259272 , n34956 );
or ( n259273 , n259271 , n259272 );
not ( n259274 , n39588 );
nand ( n259275 , n259274 , n34968 );
nand ( n259276 , n259273 , n259275 );
and ( n259277 , n259276 , n35418 );
not ( n259278 , n259276 );
and ( n259279 , n259278 , n35410 );
nor ( n259280 , n259277 , n259279 );
not ( n259281 , n259280 );
nand ( n259282 , n259281 , n234111 );
or ( n259283 , n259270 , n259282 );
nor ( n259284 , n259281 , n50944 );
nand ( n259285 , n259270 , n259284 );
nand ( n259286 , n31577 , n42610 );
nand ( n259287 , n259283 , n259285 , n259286 );
buf ( n259288 , n259287 );
buf ( n259289 , n29196 );
buf ( n259290 , n222721 );
not ( n259291 , n259290 );
not ( n259292 , n244009 );
or ( n259293 , n259291 , n259292 );
or ( n259294 , n244009 , n259290 );
nand ( n259295 , n259293 , n259294 );
and ( n259296 , n259295 , n244056 );
not ( n259297 , n259295 );
and ( n259298 , n259297 , n257630 );
nor ( n259299 , n259296 , n259298 );
not ( n259300 , n259299 );
not ( n259301 , n234069 );
not ( n259302 , n38232 );
or ( n259303 , n259301 , n259302 );
or ( n259304 , n38232 , n234069 );
nand ( n259305 , n259303 , n259304 );
not ( n259306 , n259305 );
not ( n259307 , n38634 );
and ( n259308 , n259306 , n259307 );
and ( n259309 , n259305 , n38634 );
nor ( n259310 , n259308 , n259309 );
nand ( n259311 , n259300 , n259310 );
nor ( n259312 , n237647 , n220412 );
not ( n259313 , n259312 );
not ( n259314 , n220413 );
nand ( n259315 , n259314 , n237647 );
nand ( n259316 , n259313 , n259315 );
and ( n259317 , n259316 , n237704 );
not ( n259318 , n259316 );
and ( n259319 , n259318 , n237701 );
nor ( n259320 , n259317 , n259319 );
nor ( n259321 , n259320 , n244216 );
not ( n259322 , n259321 );
or ( n259323 , n259311 , n259322 );
not ( n259324 , n259320 );
nor ( n259325 , n259324 , n39763 );
nand ( n259326 , n259325 , n259311 );
nand ( n259327 , n31576 , n204952 );
nand ( n259328 , n259323 , n259326 , n259327 );
buf ( n259329 , n259328 );
buf ( n259330 , n33751 );
not ( n259331 , n45987 );
not ( n259332 , n249489 );
not ( n259333 , n259332 );
or ( n259334 , n259331 , n259333 );
or ( n259335 , n249494 , n45987 );
nand ( n259336 , n259334 , n259335 );
and ( n259337 , n259336 , n248000 );
not ( n259338 , n259336 );
buf ( n259339 , n247991 );
and ( n259340 , n259338 , n259339 );
nor ( n259341 , n259337 , n259340 );
not ( n259342 , n259341 );
not ( n259343 , n235203 );
not ( n259344 , n53098 );
not ( n259345 , n259344 );
not ( n259346 , n252348 );
or ( n259347 , n259345 , n259346 );
nand ( n259348 , n42436 , n53098 );
nand ( n259349 , n259347 , n259348 );
not ( n259350 , n259349 );
or ( n259351 , n259343 , n259350 );
or ( n259352 , n259349 , n235203 );
nand ( n259353 , n259351 , n259352 );
not ( n259354 , n259353 );
nand ( n259355 , n241376 , n259342 , n259354 );
not ( n259356 , n241372 );
not ( n259357 , n259356 );
not ( n259358 , n259342 );
or ( n259359 , n259357 , n259358 );
not ( n259360 , n259353 );
nor ( n259361 , n259360 , n39763 );
nand ( n259362 , n259359 , n259361 );
nand ( n259363 , n233501 , n205330 );
nand ( n259364 , n259355 , n259362 , n259363 );
buf ( n259365 , n259364 );
buf ( n259366 , n250315 );
not ( n259367 , n259366 );
not ( n259368 , n237148 );
or ( n259369 , n259367 , n259368 );
not ( n259370 , n237148 );
not ( n259371 , n259370 );
or ( n259372 , n259371 , n259366 );
nand ( n259373 , n259369 , n259372 );
and ( n259374 , n259373 , n237342 );
not ( n259375 , n259373 );
and ( n259376 , n259375 , n250412 );
nor ( n259377 , n259374 , n259376 );
nand ( n259378 , n259377 , n222531 );
not ( n259379 , n48157 );
not ( n259380 , n226557 );
or ( n259381 , n259379 , n259380 );
not ( n259382 , n48157 );
nand ( n259383 , n259382 , n48804 );
nand ( n259384 , n259381 , n259383 );
not ( n259385 , n253807 );
and ( n259386 , n259384 , n259385 );
not ( n259387 , n259384 );
buf ( n259388 , n253807 );
and ( n259389 , n259387 , n259388 );
nor ( n259390 , n259386 , n259389 );
or ( n259391 , n259378 , n259390 );
nor ( n259392 , n259377 , n251190 );
not ( n259393 , n244532 );
not ( n259394 , n252790 );
not ( n259395 , n259394 );
not ( n259396 , n50940 );
or ( n259397 , n259395 , n259396 );
nand ( n259398 , n50930 , n252790 );
nand ( n259399 , n259397 , n259398 );
not ( n259400 , n259399 );
or ( n259401 , n259393 , n259400 );
or ( n259402 , n259399 , n244532 );
nand ( n259403 , n259401 , n259402 );
not ( n259404 , n259390 );
nor ( n259405 , n259403 , n259404 );
nand ( n259406 , n259392 , n259405 );
not ( n259407 , n244789 );
not ( n259408 , n259407 );
not ( n259409 , n30783 );
and ( n259410 , n259408 , n259409 );
nor ( n259411 , n259390 , n249030 );
and ( n259412 , n259411 , n259403 );
nor ( n259413 , n259410 , n259412 );
nand ( n259414 , n259391 , n259406 , n259413 );
buf ( n259415 , n259414 );
buf ( n259416 , n31698 );
not ( n259417 , n32522 );
not ( n259418 , n254441 );
or ( n259419 , n259417 , n259418 );
nand ( n259420 , n256140 , n256155 );
and ( n259421 , n259420 , n257246 );
not ( n259422 , n259420 );
and ( n259423 , n259422 , n257245 );
nor ( n259424 , n259421 , n259423 );
buf ( n259425 , n35816 );
or ( n259426 , n259424 , n259425 );
nand ( n259427 , n259419 , n259426 );
buf ( n259428 , n259427 );
buf ( n259429 , n42337 );
not ( n259430 , RI19a89e28_2725);
or ( n259431 , n25335 , n259430 );
not ( n259432 , RI1754a630_70);
and ( n259433 , n51375 , n259432 );
nor ( n259434 , n259433 , RI1754c250_10);
not ( n259435 , n259434 );
nand ( n259436 , n259435 , n51363 );
nand ( n259437 , n259431 , n259436 );
buf ( n259438 , n259437 );
nand ( n259439 , n256651 , n205649 );
nor ( n259440 , n256664 , n255701 );
or ( n259441 , n259439 , n259440 );
nor ( n259442 , n256651 , n236795 );
nand ( n259443 , n259442 , n259440 );
nand ( n259444 , n251465 , n28561 );
nand ( n259445 , n259441 , n259443 , n259444 );
buf ( n259446 , n259445 );
or ( n259447 , n25328 , n246097 );
not ( n259448 , RI19a964e8_2638);
or ( n259449 , n25335 , n259448 );
nand ( n259450 , n259447 , n259449 );
buf ( n259451 , n259450 );
not ( n259452 , n255250 );
nand ( n259453 , n259452 , n43969 );
buf ( n259454 , n246601 );
nor ( n259455 , n255464 , n259454 );
not ( n259456 , n259455 );
nand ( n259457 , n255464 , n259454 );
nand ( n259458 , n259456 , n259457 );
buf ( n259459 , n253074 );
not ( n259460 , n259459 );
and ( n259461 , n259458 , n259460 );
not ( n259462 , n259458 );
buf ( n259463 , n253073 );
not ( n259464 , n259463 );
and ( n259465 , n259462 , n259464 );
nor ( n259466 , n259461 , n259465 );
nand ( n259467 , n259466 , n255262 );
or ( n259468 , n259453 , n259467 );
not ( n259469 , n259466 );
not ( n259470 , n259452 );
or ( n259471 , n259469 , n259470 );
nor ( n259472 , n255262 , n55108 );
nand ( n259473 , n259471 , n259472 );
nand ( n259474 , n244987 , n32740 );
nand ( n259475 , n259468 , n259473 , n259474 );
buf ( n259476 , n259475 );
buf ( n259477 , n241438 );
not ( n259478 , n259477 );
not ( n259479 , n225301 );
or ( n259480 , n259478 , n259479 );
or ( n259481 , n225301 , n259477 );
nand ( n259482 , n259480 , n259481 );
and ( n259483 , n259482 , n225536 );
not ( n259484 , n259482 );
and ( n259485 , n259484 , n256892 );
nor ( n259486 , n259483 , n259485 );
nand ( n259487 , n259486 , n223839 );
not ( n259488 , n237623 );
not ( n259489 , n41216 );
or ( n259490 , n259488 , n259489 );
not ( n259491 , n237623 );
nand ( n259492 , n259491 , n233987 );
nand ( n259493 , n259490 , n259492 );
and ( n259494 , n259493 , n233990 );
not ( n259495 , n259493 );
and ( n259496 , n259495 , n253206 );
nor ( n259497 , n259494 , n259496 );
not ( n259498 , n259497 );
not ( n259499 , n251658 );
not ( n259500 , n46941 );
or ( n259501 , n259499 , n259500 );
not ( n259502 , n251658 );
nand ( n259503 , n259502 , n46950 );
nand ( n259504 , n259501 , n259503 );
and ( n259505 , n259504 , n47157 );
not ( n259506 , n259504 );
and ( n259507 , n259506 , n224925 );
nor ( n259508 , n259505 , n259507 );
not ( n259509 , n259508 );
nand ( n259510 , n259498 , n259509 );
or ( n259511 , n259487 , n259510 );
not ( n259512 , n259498 );
not ( n259513 , n259486 );
or ( n259514 , n259512 , n259513 );
nand ( n259515 , n259508 , n247444 );
not ( n259516 , n259515 );
nand ( n259517 , n259514 , n259516 );
nand ( n259518 , n247585 , n28691 );
nand ( n259519 , n259511 , n259517 , n259518 );
buf ( n259520 , n259519 );
not ( n259521 , n237802 );
not ( n259522 , n245392 );
or ( n259523 , n259521 , n259522 );
nand ( n259524 , n245402 , n237799 );
nand ( n259525 , n259523 , n259524 );
not ( n259526 , n259525 );
buf ( n259527 , n254916 );
not ( n259528 , n259527 );
and ( n259529 , n259526 , n259528 );
not ( n259530 , n254916 );
not ( n259531 , n259530 );
and ( n259532 , n259525 , n259531 );
nor ( n259533 , n259529 , n259532 );
nor ( n259534 , n259533 , n39763 );
not ( n259535 , n43768 );
not ( n259536 , n252552 );
or ( n259537 , n259535 , n259536 );
not ( n259538 , n43768 );
nand ( n259539 , n259538 , n252561 );
nand ( n259540 , n259537 , n259539 );
and ( n259541 , n259540 , n255673 );
not ( n259542 , n259540 );
not ( n259543 , n255673 );
and ( n259544 , n259542 , n259543 );
nor ( n259545 , n259541 , n259544 );
not ( n259546 , n259545 );
not ( n259547 , n53032 );
not ( n259548 , n42149 );
or ( n259549 , n259547 , n259548 );
not ( n259550 , n53032 );
nand ( n259551 , n259550 , n42156 );
nand ( n259552 , n259549 , n259551 );
not ( n259553 , n252348 );
and ( n259554 , n259552 , n259553 );
not ( n259555 , n259552 );
and ( n259556 , n259555 , n220201 );
nor ( n259557 , n259554 , n259556 );
not ( n259558 , n259557 );
nand ( n259559 , n259534 , n259546 , n259558 );
not ( n259560 , n259533 );
not ( n259561 , n259560 );
not ( n259562 , n259546 );
or ( n259563 , n259561 , n259562 );
nor ( n259564 , n259558 , n250431 );
nand ( n259565 , n259563 , n259564 );
nand ( n259566 , n31577 , n35563 );
nand ( n259567 , n259559 , n259565 , n259566 );
buf ( n259568 , n259567 );
not ( n259569 , n241935 );
not ( n259570 , n256152 );
or ( n259571 , n259569 , n259570 );
not ( n259572 , n241935 );
nand ( n259573 , n259572 , n237590 );
nand ( n259574 , n259571 , n259573 );
not ( n259575 , n253385 );
and ( n259576 , n259574 , n259575 );
not ( n259577 , n259574 );
buf ( n259578 , n234682 );
and ( n259579 , n259577 , n259578 );
nor ( n259580 , n259576 , n259579 );
nand ( n259581 , n259580 , n234111 );
not ( n259582 , n249679 );
not ( n259583 , n255830 );
or ( n259584 , n259582 , n259583 );
not ( n259585 , n249679 );
not ( n259586 , n248339 );
not ( n259587 , n248380 );
and ( n259588 , n259586 , n259587 );
and ( n259589 , n248339 , n248380 );
nor ( n259590 , n259588 , n259589 );
nand ( n259591 , n259585 , n259590 );
nand ( n259592 , n259584 , n259591 );
and ( n259593 , n259592 , n255885 );
not ( n259594 , n259592 );
buf ( n259595 , n255879 );
and ( n259596 , n259594 , n259595 );
nor ( n259597 , n259593 , n259596 );
not ( n259598 , n255408 );
buf ( n259599 , n246541 );
not ( n259600 , n259599 );
and ( n259601 , n259598 , n259600 );
and ( n259602 , n236502 , n259599 );
nor ( n259603 , n259601 , n259602 );
and ( n259604 , n259603 , n255455 );
not ( n259605 , n259603 );
and ( n259606 , n259605 , n255465 );
nor ( n259607 , n259604 , n259606 );
not ( n259608 , n259607 );
nand ( n259609 , n259597 , n259608 );
or ( n259610 , n259581 , n259609 );
not ( n259611 , n259597 );
not ( n259612 , n259580 );
or ( n259613 , n259611 , n259612 );
nor ( n259614 , n259608 , n40465 );
nand ( n259615 , n259613 , n259614 );
nand ( n259616 , n234024 , n205690 );
nand ( n259617 , n259610 , n259615 , n259616 );
buf ( n259618 , n259617 );
not ( n259619 , n40465 );
nand ( n259620 , n259341 , n259619 );
not ( n259621 , n241185 );
nand ( n259622 , n259621 , n259354 );
or ( n259623 , n259620 , n259622 );
not ( n259624 , n259360 );
not ( n259625 , n259341 );
or ( n259626 , n259624 , n259625 );
nor ( n259627 , n259621 , n235050 );
nand ( n259628 , n259626 , n259627 );
nand ( n259629 , n234024 , n205333 );
nand ( n259630 , n259623 , n259628 , n259629 );
buf ( n259631 , n259630 );
not ( n259632 , n31039 );
not ( n259633 , n258213 );
or ( n259634 , n259632 , n259633 );
nand ( n259635 , n251360 , n251352 );
not ( n259636 , n237402 );
not ( n259637 , n247813 );
or ( n259638 , n259636 , n259637 );
not ( n259639 , n237402 );
nand ( n259640 , n259639 , n247822 );
nand ( n259641 , n259638 , n259640 );
and ( n259642 , n259641 , n247872 );
not ( n259643 , n259641 );
and ( n259644 , n259643 , n247873 );
nor ( n259645 , n259642 , n259644 );
not ( n259646 , n259645 );
and ( n259647 , n259635 , n259646 );
not ( n259648 , n259635 );
and ( n259649 , n259648 , n259645 );
nor ( n259650 , n259647 , n259649 );
buf ( n259651 , n55152 );
or ( n259652 , n259650 , n259651 );
nand ( n259653 , n259634 , n259652 );
buf ( n259654 , n259653 );
not ( n259655 , n224463 );
not ( n259656 , n253196 );
or ( n259657 , n259655 , n259656 );
not ( n259658 , n224463 );
nand ( n259659 , n259658 , n253188 );
nand ( n259660 , n259657 , n259659 );
and ( n259661 , n259660 , n253948 );
not ( n259662 , n259660 );
and ( n259663 , n259662 , n253949 );
nor ( n259664 , n259661 , n259663 );
not ( n259665 , n259664 );
not ( n259666 , n247491 );
not ( n259667 , n243510 );
or ( n259668 , n259666 , n259667 );
not ( n259669 , n247491 );
nand ( n259670 , n259669 , n243503 );
nand ( n259671 , n259668 , n259670 );
and ( n259672 , n259671 , n248481 );
not ( n259673 , n259671 );
and ( n259674 , n259673 , n248478 );
nor ( n259675 , n259672 , n259674 );
not ( n259676 , n259675 );
nand ( n259677 , n259665 , n259676 );
or ( n259678 , n259378 , n259677 );
nand ( n259679 , n259392 , n259677 );
nand ( n259680 , n245943 , n33500 );
nand ( n259681 , n259678 , n259679 , n259680 );
buf ( n259682 , n259681 );
not ( n259683 , n251896 );
buf ( n259684 , n239214 );
not ( n259685 , n259684 );
not ( n259686 , n240141 );
or ( n259687 , n259685 , n259686 );
or ( n259688 , n240148 , n259684 );
nand ( n259689 , n259687 , n259688 );
and ( n259690 , n259689 , n255353 );
not ( n259691 , n259689 );
and ( n259692 , n259691 , n255356 );
nor ( n259693 , n259690 , n259692 );
buf ( n259694 , n254564 );
not ( n259695 , n259694 );
not ( n259696 , n249462 );
or ( n259697 , n259695 , n259696 );
not ( n259698 , n259694 );
nand ( n259699 , n259698 , n249469 );
nand ( n259700 , n259697 , n259699 );
buf ( n259701 , n233660 );
and ( n259702 , n259700 , n259701 );
not ( n259703 , n259700 );
buf ( n259704 , n55889 );
and ( n259705 , n259703 , n259704 );
nor ( n259706 , n259702 , n259705 );
nor ( n259707 , n259693 , n259706 );
or ( n259708 , n259683 , n259707 );
nand ( n259709 , n251883 , n259707 );
nand ( n259710 , n249622 , n34185 );
nand ( n259711 , n259708 , n259709 , n259710 );
buf ( n259712 , n259711 );
buf ( n259713 , n25367 );
not ( n259714 , RI19ab65b8_2406);
or ( n259715 , n25328 , n259714 );
not ( n259716 , RI19aacbf8_2477);
or ( n259717 , n25335 , n259716 );
nand ( n259718 , n259715 , n259717 );
buf ( n259719 , n259718 );
buf ( n259720 , n204289 );
not ( n259721 , n28198 );
not ( n259722 , n255116 );
or ( n259723 , n259721 , n259722 );
not ( n259724 , n42035 );
not ( n259725 , n234243 );
or ( n259726 , n259724 , n259725 );
not ( n259727 , n42035 );
nand ( n259728 , n259727 , n234252 );
nand ( n259729 , n259726 , n259728 );
and ( n259730 , n259729 , n234306 );
not ( n259731 , n259729 );
and ( n259732 , n259731 , n234299 );
nor ( n259733 , n259730 , n259732 );
and ( n259734 , n243403 , n243410 );
not ( n259735 , n243403 );
and ( n259736 , n259735 , n243413 );
nor ( n259737 , n259734 , n259736 );
not ( n259738 , n259737 );
not ( n259739 , n259738 );
not ( n259740 , n49674 );
and ( n259741 , n259739 , n259740 );
and ( n259742 , n246693 , n49674 );
nor ( n259743 , n259741 , n259742 );
buf ( n259744 , n245862 );
and ( n259745 , n259743 , n259744 );
not ( n259746 , n259743 );
buf ( n259747 , n245872 );
and ( n259748 , n259746 , n259747 );
nor ( n259749 , n259745 , n259748 );
nand ( n259750 , n259733 , n259749 );
and ( n259751 , n247613 , n48232 );
not ( n259752 , n247613 );
and ( n259753 , n259752 , n48233 );
or ( n259754 , n259751 , n259753 );
not ( n259755 , n253464 );
not ( n259756 , n259755 );
xnor ( n259757 , n259754 , n259756 );
and ( n259758 , n259750 , n259757 );
not ( n259759 , n259750 );
not ( n259760 , n259757 );
and ( n259761 , n259759 , n259760 );
nor ( n259762 , n259758 , n259761 );
or ( n259763 , n259762 , n49959 );
nand ( n259764 , n259723 , n259763 );
buf ( n259765 , n259764 );
not ( n259766 , RI19ab8d90_2389);
or ( n259767 , n226819 , n259766 );
not ( n259768 , RI19aaf088_2461);
or ( n259769 , n25335 , n259768 );
nand ( n259770 , n259767 , n259769 );
buf ( n259771 , n259770 );
not ( n259772 , n250566 );
not ( n259773 , n227174 );
or ( n259774 , n259772 , n259773 );
not ( n259775 , n250566 );
nand ( n259776 , n259775 , n49420 );
nand ( n259777 , n259774 , n259776 );
and ( n259778 , n259777 , n49618 );
not ( n259779 , n259777 );
and ( n259780 , n259779 , n49627 );
nor ( n259781 , n259778 , n259780 );
not ( n259782 , n259781 );
not ( n259783 , n234818 );
nand ( n259784 , n259782 , n259783 );
not ( n259785 , n238199 );
nand ( n259786 , n238188 , n259785 );
or ( n259787 , n259784 , n259786 );
not ( n259788 , n259785 );
not ( n259789 , n259782 );
or ( n259790 , n259788 , n259789 );
nor ( n259791 , n238188 , n221279 );
nand ( n259792 , n259790 , n259791 );
nand ( n259793 , n35431 , n26374 );
nand ( n259794 , n259787 , n259792 , n259793 );
buf ( n259795 , n259794 );
nand ( n259796 , n246770 , n249772 );
or ( n259797 , n246698 , n259796 );
not ( n259798 , n246770 );
not ( n259799 , n246696 );
or ( n259800 , n259798 , n259799 );
not ( n259801 , n205649 );
nor ( n259802 , n249772 , n259801 );
nand ( n259803 , n259800 , n259802 );
nand ( n259804 , n239240 , n33108 );
nand ( n259805 , n259797 , n259803 , n259804 );
buf ( n259806 , n259805 );
buf ( n259807 , n241752 );
not ( n259808 , n259807 );
not ( n259809 , n248892 );
or ( n259810 , n259808 , n259809 );
or ( n259811 , n248892 , n259807 );
nand ( n259812 , n259810 , n259811 );
and ( n259813 , n259812 , n248904 );
not ( n259814 , n259812 );
and ( n259815 , n259814 , n248907 );
nor ( n259816 , n259813 , n259815 );
not ( n259817 , n39690 );
not ( n259818 , n35409 );
or ( n259819 , n259817 , n259818 );
not ( n259820 , n39690 );
nand ( n259821 , n259820 , n35417 );
nand ( n259822 , n259819 , n259821 );
and ( n259823 , n259822 , n249601 );
not ( n259824 , n259822 );
and ( n259825 , n259824 , n249611 );
nor ( n259826 , n259823 , n259825 );
nand ( n259827 , n259816 , n259826 );
or ( n259828 , n259515 , n259827 );
not ( n259829 , n259816 );
not ( n259830 , n259508 );
or ( n259831 , n259829 , n259830 );
nor ( n259832 , n259826 , n226003 );
nand ( n259833 , n259831 , n259832 );
nand ( n259834 , n50615 , n25984 );
nand ( n259835 , n259828 , n259833 , n259834 );
buf ( n259836 , n259835 );
not ( n259837 , n243190 );
not ( n259838 , n253293 );
or ( n259839 , n259837 , n259838 );
or ( n259840 , n248677 , n243190 );
nand ( n259841 , n259839 , n259840 );
and ( n259842 , n259841 , n253287 );
not ( n259843 , n259841 );
and ( n259844 , n259843 , n253288 );
nor ( n259845 , n259842 , n259844 );
not ( n259846 , n259845 );
not ( n259847 , n235732 );
nand ( n259848 , n259846 , n259847 );
not ( n259849 , n40336 );
not ( n259850 , n235878 );
or ( n259851 , n259849 , n259850 );
not ( n259852 , n40336 );
nand ( n259853 , n259852 , n235887 );
nand ( n259854 , n259851 , n259853 );
buf ( n259855 , n243363 );
and ( n259856 , n259854 , n259855 );
not ( n259857 , n259854 );
buf ( n259858 , n243372 );
and ( n259859 , n259857 , n259858 );
nor ( n259860 , n259856 , n259859 );
not ( n259861 , n37237 );
not ( n259862 , n259861 );
not ( n259863 , n240799 );
or ( n259864 , n259862 , n259863 );
not ( n259865 , n259861 );
nand ( n259866 , n259865 , n240810 );
nand ( n259867 , n259864 , n259866 );
and ( n259868 , n259867 , n252444 );
not ( n259869 , n259867 );
and ( n259870 , n259869 , n252447 );
nor ( n259871 , n259868 , n259870 );
nand ( n259872 , n259860 , n259871 );
or ( n259873 , n259848 , n259872 );
not ( n259874 , n259871 );
not ( n259875 , n259846 );
or ( n259876 , n259874 , n259875 );
nor ( n259877 , n259860 , n50944 );
nand ( n259878 , n259876 , n259877 );
nand ( n259879 , n31576 , n27804 );
nand ( n259880 , n259873 , n259878 , n259879 );
buf ( n259881 , n259880 );
buf ( n259882 , n243357 );
and ( n259883 , n259882 , n250805 );
not ( n259884 , n259882 );
and ( n259885 , n259884 , n250811 );
nor ( n259886 , n259883 , n259885 );
not ( n259887 , n259886 );
not ( n259888 , n257379 );
and ( n259889 , n259887 , n259888 );
and ( n259890 , n259886 , n257379 );
nor ( n259891 , n259889 , n259890 );
not ( n259892 , n239912 );
not ( n259893 , n247569 );
or ( n259894 , n259892 , n259893 );
not ( n259895 , n239912 );
nand ( n259896 , n259895 , n230199 );
nand ( n259897 , n259894 , n259896 );
and ( n259898 , n259897 , n242696 );
not ( n259899 , n259897 );
and ( n259900 , n259899 , n247575 );
nor ( n259901 , n259898 , n259900 );
not ( n259902 , n259901 );
nand ( n259903 , n259891 , n259902 );
not ( n259904 , n241953 );
not ( n259905 , n237590 );
not ( n259906 , n259905 );
or ( n259907 , n259904 , n259906 );
not ( n259908 , n241953 );
nand ( n259909 , n259908 , n237590 );
nand ( n259910 , n259907 , n259909 );
and ( n259911 , n259910 , n259575 );
not ( n259912 , n259910 );
and ( n259913 , n259912 , n259578 );
nor ( n259914 , n259911 , n259913 );
nand ( n259915 , n259903 , n259914 , n252259 );
nor ( n259916 , n259901 , n40465 );
not ( n259917 , n259914 );
nand ( n259918 , n259916 , n259917 , n259891 );
nand ( n259919 , n31577 , n40038 );
nand ( n259920 , n259915 , n259918 , n259919 );
buf ( n259921 , n259920 );
nor ( n259922 , n244594 , n235050 );
not ( n259923 , n248512 );
not ( n259924 , n243659 );
or ( n259925 , n259923 , n259924 );
or ( n259926 , n243659 , n248512 );
nand ( n259927 , n259925 , n259926 );
and ( n259928 , n259927 , n251846 );
not ( n259929 , n259927 );
and ( n259930 , n259929 , n251856 );
nor ( n259931 , n259928 , n259930 );
not ( n259932 , n234492 );
not ( n259933 , n49043 );
or ( n259934 , n259932 , n259933 );
not ( n259935 , n234492 );
nand ( n259936 , n259935 , n234121 );
nand ( n259937 , n259934 , n259936 );
and ( n259938 , n259937 , n234186 );
not ( n259939 , n259937 );
and ( n259940 , n259939 , n234185 );
nor ( n259941 , n259938 , n259940 );
nand ( n259942 , n259922 , n259931 , n259941 );
not ( n259943 , n259931 );
nand ( n259944 , n259941 , n244593 );
nand ( n259945 , n259943 , n259944 , n239934 );
nand ( n259946 , n224937 , n36291 );
nand ( n259947 , n259942 , n259945 , n259946 );
buf ( n259948 , n259947 );
not ( n259949 , n238007 );
not ( n259950 , n226319 );
or ( n259951 , n259949 , n259950 );
nand ( n259952 , n257110 , n238006 );
nand ( n259953 , n259951 , n259952 );
and ( n259954 , n259953 , n257116 );
not ( n259955 , n259953 );
and ( n259956 , n259955 , n258557 );
nor ( n259957 , n259954 , n259956 );
not ( n259958 , n259957 );
nor ( n259959 , n259958 , n235050 );
not ( n259960 , n259959 );
not ( n259961 , n39546 );
not ( n259962 , n34956 );
or ( n259963 , n259961 , n259962 );
not ( n259964 , n39546 );
nand ( n259965 , n259964 , n34968 );
nand ( n259966 , n259963 , n259965 );
and ( n259967 , n259966 , n35410 );
not ( n259968 , n259966 );
and ( n259969 , n259968 , n35418 );
nor ( n259970 , n259967 , n259969 );
not ( n259971 , n43335 );
not ( n259972 , n238894 );
or ( n259973 , n259971 , n259972 );
not ( n259974 , n43335 );
nand ( n259975 , n259974 , n246077 );
nand ( n259976 , n259973 , n259975 );
and ( n259977 , n259976 , n246082 );
not ( n259978 , n259976 );
and ( n259979 , n259978 , n244453 );
nor ( n259980 , n259977 , n259979 );
not ( n259981 , n259980 );
nand ( n259982 , n259970 , n259981 );
or ( n259983 , n259960 , n259982 );
not ( n259984 , n259970 );
not ( n259985 , n259957 );
or ( n259986 , n259984 , n259985 );
nor ( n259987 , n259981 , n27889 );
nand ( n259988 , n259986 , n259987 );
nand ( n259989 , n252711 , n39303 );
nand ( n259990 , n259983 , n259988 , n259989 );
buf ( n259991 , n259990 );
not ( n259992 , n235772 );
not ( n259993 , n245738 );
or ( n259994 , n259992 , n259993 );
nand ( n259995 , n245743 , n235775 );
nand ( n259996 , n259994 , n259995 );
and ( n259997 , n259996 , n245794 );
not ( n259998 , n259996 );
and ( n259999 , n259998 , n245799 );
nor ( n260000 , n259997 , n259999 );
nand ( n260001 , n260000 , n54200 );
buf ( n260002 , n36899 );
not ( n260003 , n260002 );
not ( n260004 , n240810 );
or ( n260005 , n260003 , n260004 );
or ( n260006 , n240810 , n260002 );
nand ( n260007 , n260005 , n260006 );
not ( n260008 , n260007 );
not ( n260009 , n252444 );
and ( n260010 , n260008 , n260009 );
not ( n260011 , n258715 );
and ( n260012 , n260007 , n260011 );
nor ( n260013 , n260010 , n260012 );
not ( n260014 , n246957 );
not ( n260015 , n256191 );
or ( n260016 , n260014 , n260015 );
not ( n260017 , n246957 );
nand ( n260018 , n260017 , n256190 );
nand ( n260019 , n260016 , n260018 );
and ( n260020 , n260019 , n249849 );
not ( n260021 , n260019 );
buf ( n260022 , n242155 );
and ( n260023 , n260021 , n260022 );
nor ( n260024 , n260020 , n260023 );
nand ( n260025 , n260013 , n260024 );
or ( n260026 , n260001 , n260025 );
not ( n260027 , n260013 );
not ( n260028 , n260000 );
or ( n260029 , n260027 , n260028 );
nor ( n260030 , n260024 , n226955 );
nand ( n260031 , n260029 , n260030 );
nand ( n260032 , n35431 , n38518 );
nand ( n260033 , n260026 , n260031 , n260032 );
buf ( n260034 , n260033 );
not ( n260035 , n44107 );
not ( n260036 , n255320 );
or ( n260037 , n260035 , n260036 );
or ( n260038 , n255320 , n44107 );
nand ( n260039 , n260037 , n260038 );
and ( n260040 , n260039 , n234098 );
not ( n260041 , n260039 );
and ( n260042 , n260041 , n234107 );
nor ( n260043 , n260040 , n260042 );
nand ( n260044 , n260043 , n245241 );
not ( n260045 , n238102 );
not ( n260046 , n47667 );
not ( n260047 , n238033 );
or ( n260048 , n260046 , n260047 );
not ( n260049 , n47667 );
nand ( n260050 , n260049 , n238040 );
nand ( n260051 , n260048 , n260050 );
not ( n260052 , n260051 );
or ( n260053 , n260045 , n260052 );
or ( n260054 , n260051 , n238102 );
nand ( n260055 , n260053 , n260054 );
not ( n260056 , n243401 );
not ( n260057 , n39052 );
or ( n260058 , n260056 , n260057 );
not ( n260059 , n243401 );
nand ( n260060 , n260059 , n39059 );
nand ( n260061 , n260058 , n260060 );
and ( n260062 , n260061 , n39435 );
not ( n260063 , n260061 );
and ( n260064 , n260063 , n39445 );
nor ( n260065 , n260062 , n260064 );
nand ( n260066 , n260055 , n260065 );
or ( n260067 , n260044 , n260066 );
not ( n260068 , n260055 );
not ( n260069 , n260043 );
or ( n260070 , n260068 , n260069 );
nor ( n260071 , n260065 , n234818 );
nand ( n260072 , n260070 , n260071 );
nand ( n260073 , n247585 , n218775 );
nand ( n260074 , n260067 , n260072 , n260073 );
buf ( n260075 , n260074 );
not ( n260076 , n239484 );
not ( n260077 , n260076 );
not ( n260078 , n249640 );
nand ( n260079 , n239455 , n239479 );
and ( n260080 , n260079 , n248305 );
not ( n260081 , n260079 );
and ( n260082 , n260081 , n248306 );
nor ( n260083 , n260080 , n260082 );
not ( n260084 , n260083 );
not ( n260085 , n260084 );
or ( n260086 , n260078 , n260085 );
nand ( n260087 , n260083 , n249639 );
nand ( n260088 , n260086 , n260087 );
and ( n260089 , n260088 , n251519 );
not ( n260090 , n260088 );
and ( n260091 , n260090 , n251520 );
nor ( n260092 , n260089 , n260091 );
buf ( n260093 , n248350 );
not ( n260094 , n260093 );
not ( n260095 , n239558 );
nand ( n260096 , n260095 , n244098 );
not ( n260097 , n260096 );
or ( n260098 , n260094 , n260097 );
or ( n260099 , n260096 , n260093 );
nand ( n260100 , n260098 , n260099 );
not ( n260101 , n260100 );
nand ( n260102 , n239520 , n246300 );
not ( n260103 , n249650 );
and ( n260104 , n260102 , n260103 );
not ( n260105 , n260102 );
and ( n260106 , n260105 , n249650 );
nor ( n260107 , n260104 , n260106 );
not ( n260108 , n260107 );
and ( n260109 , n260101 , n260108 );
and ( n260110 , n260100 , n260107 );
nor ( n260111 , n260109 , n260110 );
xor ( n260112 , n260092 , n260111 );
not ( n260113 , n260112 );
or ( n260114 , n260077 , n260113 );
not ( n260115 , n260076 );
not ( n260116 , n260111 );
not ( n260117 , n260092 );
or ( n260118 , n260116 , n260117 );
not ( n260119 , n260092 );
not ( n260120 , n260111 );
nand ( n260121 , n260119 , n260120 );
nand ( n260122 , n260118 , n260121 );
nand ( n260123 , n260115 , n260122 );
nand ( n260124 , n260114 , n260123 );
buf ( n260125 , n36368 );
and ( n260126 , n260124 , n260125 );
not ( n260127 , n260124 );
and ( n260128 , n260127 , n36372 );
nor ( n260129 , n260126 , n260128 );
nand ( n260130 , n246681 , n260129 );
not ( n260131 , n251961 );
not ( n260132 , n251689 );
not ( n260133 , n260132 );
or ( n260134 , n260131 , n260133 );
nand ( n260135 , n251689 , n251960 );
nand ( n260136 , n260134 , n260135 );
and ( n260137 , n260136 , n257307 );
not ( n260138 , n260136 );
and ( n260139 , n260138 , n257308 );
nor ( n260140 , n260137 , n260139 );
not ( n260141 , n260140 );
or ( n260142 , n260130 , n260141 );
nand ( n260143 , n260129 , n246675 );
nand ( n260144 , n260143 , n260141 , n249009 );
nand ( n260145 , n239240 , n31440 );
nand ( n260146 , n260142 , n260144 , n260145 );
buf ( n260147 , n260146 );
not ( n260148 , n40685 );
not ( n260149 , n251450 );
or ( n260150 , n260148 , n260149 );
nand ( n260151 , n251443 , n40686 );
nand ( n260152 , n260150 , n260151 );
not ( n260153 , n260152 );
not ( n260154 , n253106 );
and ( n260155 , n260153 , n260154 );
and ( n260156 , n260152 , n253106 );
nor ( n260157 , n260155 , n260156 );
nand ( n260158 , n260157 , n259619 );
not ( n260159 , n243454 );
nand ( n260160 , n255129 , n260159 );
or ( n260161 , n260158 , n260160 );
not ( n260162 , n255129 );
not ( n260163 , n260157 );
or ( n260164 , n260162 , n260163 );
nor ( n260165 , n260159 , n234440 );
nand ( n260166 , n260164 , n260165 );
nand ( n260167 , n31577 , n34869 );
nand ( n260168 , n260161 , n260166 , n260167 );
buf ( n260169 , n260168 );
not ( n260170 , n49629 );
nand ( n260171 , n260170 , n49953 );
nand ( n260172 , n244464 , n244809 );
or ( n260173 , n260171 , n260172 );
nand ( n260174 , n244465 , n260171 );
nand ( n260175 , n39767 , n28860 );
nand ( n260176 , n260173 , n260174 , n260175 );
buf ( n260177 , n260176 );
not ( n260178 , RI19abd6b0_2355);
or ( n260179 , n25328 , n260178 );
not ( n260180 , RI19ab3840_2427);
or ( n260181 , n25335 , n260180 );
nand ( n260182 , n260179 , n260181 );
buf ( n260183 , n260182 );
not ( n260184 , RI1754b1e8_45);
or ( n260185 , n249126 , n260184 );
nand ( n260186 , n249131 , n28363 );
nand ( n260187 , n260185 , n260186 );
buf ( n260188 , n260187 );
not ( n260189 , n249701 );
not ( n260190 , n255884 );
or ( n260191 , n260189 , n260190 );
not ( n260192 , n249701 );
nand ( n260193 , n260192 , n255879 );
nand ( n260194 , n260191 , n260193 );
buf ( n260195 , n46506 );
and ( n260196 , n260194 , n260195 );
not ( n260197 , n260194 );
buf ( n260198 , n46514 );
and ( n260199 , n260197 , n260198 );
nor ( n260200 , n260196 , n260199 );
nor ( n260201 , n259466 , n260200 );
or ( n260202 , n255251 , n260201 );
nor ( n260203 , n255250 , n236795 );
nand ( n260204 , n260203 , n260201 );
nand ( n260205 , n239240 , n26112 );
nand ( n260206 , n260202 , n260204 , n260205 );
buf ( n260207 , n260206 );
buf ( n260208 , n254544 );
not ( n260209 , n260208 );
not ( n260210 , n249462 );
or ( n260211 , n260209 , n260210 );
or ( n260212 , n249462 , n260208 );
nand ( n260213 , n260211 , n260212 );
not ( n260214 , n260213 );
not ( n260215 , n259704 );
and ( n260216 , n260214 , n260215 );
and ( n260217 , n260213 , n259704 );
nor ( n260218 , n260216 , n260217 );
nand ( n260219 , n260218 , n43969 );
buf ( n260220 , n248945 );
not ( n260221 , n260220 );
not ( n260222 , n250099 );
or ( n260223 , n260221 , n260222 );
or ( n260224 , n250102 , n260220 );
nand ( n260225 , n260223 , n260224 );
and ( n260226 , n260225 , n250108 );
not ( n260227 , n260225 );
and ( n260228 , n260227 , n250105 );
nor ( n260229 , n260226 , n260228 );
not ( n260230 , n260229 );
nand ( n260231 , n260230 , n246084 );
or ( n260232 , n260219 , n260231 );
not ( n260233 , n260218 );
not ( n260234 , n260230 );
or ( n260235 , n260233 , n260234 );
nor ( n260236 , n246084 , n31571 );
nand ( n260237 , n260235 , n260236 );
nand ( n260238 , n234453 , n36152 );
nand ( n260239 , n260232 , n260237 , n260238 );
buf ( n260240 , n260239 );
not ( n260241 , RI19a98d38_2620);
or ( n260242 , n25328 , n260241 );
not ( n260243 , RI19a8ed60_2691);
or ( n260244 , n25336 , n260243 );
nand ( n260245 , n260242 , n260244 );
buf ( n260246 , n260245 );
not ( n260247 , n54125 );
not ( n260248 , n242307 );
not ( n260249 , n260248 );
or ( n260250 , n260247 , n260249 );
or ( n260251 , n260248 , n54125 );
nand ( n260252 , n260250 , n260251 );
and ( n260253 , n260252 , n242374 );
not ( n260254 , n260252 );
and ( n260255 , n260254 , n242381 );
nor ( n260256 , n260253 , n260255 );
nand ( n260257 , n260256 , n241704 );
not ( n260258 , n259749 );
nand ( n260259 , n259733 , n260258 );
or ( n260260 , n260257 , n260259 );
not ( n260261 , n260258 );
not ( n260262 , n260256 );
or ( n260263 , n260261 , n260262 );
nor ( n260264 , n259733 , n35427 );
nand ( n260265 , n260263 , n260264 );
nand ( n260266 , n241976 , n25718 );
nand ( n260267 , n260260 , n260265 , n260266 );
buf ( n260268 , n260267 );
not ( n260269 , n236385 );
not ( n260270 , n51901 );
and ( n260271 , n260269 , n260270 );
and ( n260272 , n245201 , n51901 );
nor ( n260273 , n260271 , n260272 );
and ( n260274 , n260273 , n245211 );
not ( n260275 , n260273 );
and ( n260276 , n260275 , n236392 );
nor ( n260277 , n260274 , n260276 );
nand ( n260278 , n241667 , n260277 );
nand ( n260279 , n241679 , n248981 );
or ( n260280 , n260278 , n260279 );
not ( n260281 , n241679 );
not ( n260282 , n241667 );
or ( n260283 , n260281 , n260282 );
nor ( n260284 , n260277 , n250431 );
nand ( n260285 , n260283 , n260284 );
nand ( n260286 , n252711 , n38449 );
nand ( n260287 , n260280 , n260285 , n260286 );
buf ( n260288 , n260287 );
not ( n260289 , RI19ab92b8_2387);
or ( n260290 , n25328 , n260289 );
or ( n260291 , n25335 , n251916 );
nand ( n260292 , n260290 , n260291 );
buf ( n260293 , n260292 );
not ( n260294 , n255551 );
not ( n260295 , n238628 );
or ( n260296 , n260294 , n260295 );
or ( n260297 , n238628 , n255551 );
nand ( n260298 , n260296 , n260297 );
and ( n260299 , n260298 , n257185 );
not ( n260300 , n260298 );
and ( n260301 , n260300 , n257188 );
nor ( n260302 , n260299 , n260301 );
not ( n260303 , n260302 );
nor ( n260304 , n260303 , n226955 );
nand ( n260305 , n260304 , n254225 );
nor ( n260306 , n260302 , n38637 );
not ( n260307 , n259160 );
not ( n260308 , n238256 );
not ( n260309 , n236166 );
not ( n260310 , n260309 );
or ( n260311 , n260308 , n260310 );
nand ( n260312 , n236166 , n238259 );
nand ( n260313 , n260311 , n260312 );
not ( n260314 , n260313 );
not ( n260315 , n260314 );
or ( n260316 , n260307 , n260315 );
nand ( n260317 , n259172 , n260313 );
nand ( n260318 , n260316 , n260317 );
nor ( n260319 , n254225 , n260318 );
nand ( n260320 , n260306 , n260319 );
not ( n260321 , n254228 );
nand ( n260322 , n260321 , n260318 );
nand ( n260323 , n39766 , n39215 );
nand ( n260324 , n260305 , n260320 , n260322 , n260323 );
buf ( n260325 , n260324 );
nand ( n260326 , n247198 , n257792 );
nor ( n260327 , n251481 , n247021 );
or ( n260328 , n260326 , n260327 );
nand ( n260329 , n247215 , n260327 );
nand ( n260330 , n245414 , n43693 );
nand ( n260331 , n260328 , n260329 , n260330 );
buf ( n260332 , n260331 );
nand ( n260333 , n258624 , n253397 );
not ( n260334 , n52838 );
not ( n260335 , n246882 );
or ( n260336 , n260334 , n260335 );
not ( n260337 , n52838 );
nand ( n260338 , n260337 , n246891 );
nand ( n260339 , n260336 , n260338 );
buf ( n260340 , n256870 );
and ( n260341 , n260339 , n260340 );
not ( n260342 , n260339 );
and ( n260343 , n260342 , n258077 );
nor ( n260344 , n260341 , n260343 );
not ( n260345 , n260344 );
not ( n260346 , n48724 );
not ( n260347 , n239220 );
or ( n260348 , n260346 , n260347 );
not ( n260349 , n48724 );
nand ( n260350 , n260349 , n239228 );
nand ( n260351 , n260348 , n260350 );
xnor ( n260352 , n260351 , n250580 );
nand ( n260353 , n260345 , n260352 );
or ( n260354 , n260333 , n260353 );
not ( n260355 , n260345 );
not ( n260356 , n258624 );
or ( n260357 , n260355 , n260356 );
nor ( n260358 , n260352 , n221279 );
nand ( n260359 , n260357 , n260358 );
nand ( n260360 , n31577 , n29386 );
nand ( n260361 , n260354 , n260359 , n260360 );
buf ( n260362 , n260361 );
not ( n260363 , n53495 );
not ( n260364 , n250496 );
or ( n260365 , n260363 , n260364 );
not ( n260366 , n53495 );
nand ( n260367 , n260366 , n255291 );
nand ( n260368 , n260365 , n260367 );
not ( n260369 , n244199 );
not ( n260370 , n260369 );
and ( n260371 , n260368 , n260370 );
not ( n260372 , n260368 );
and ( n260373 , n260372 , n255295 );
nor ( n260374 , n260371 , n260373 );
not ( n260375 , n50944 );
nand ( n260376 , n260374 , n260375 );
not ( n260377 , n238091 );
not ( n260378 , n260377 );
not ( n260379 , n247669 );
not ( n260380 , n247684 );
or ( n260381 , n260379 , n260380 );
nand ( n260382 , n247685 , n247670 );
nand ( n260383 , n260381 , n260382 );
not ( n260384 , n260383 );
not ( n260385 , n260384 );
or ( n260386 , n260378 , n260385 );
not ( n260387 , n260377 );
nand ( n260388 , n260387 , n260383 );
nand ( n260389 , n260386 , n260388 );
and ( n260390 , n260389 , n247645 );
not ( n260391 , n260389 );
and ( n260392 , n260391 , n247646 );
nor ( n260393 , n260390 , n260392 );
not ( n260394 , n260393 );
not ( n260395 , n37715 );
not ( n260396 , n245572 );
not ( n260397 , n37290 );
or ( n260398 , n260396 , n260397 );
nand ( n260399 , n37289 , n245573 );
nand ( n260400 , n260398 , n260399 );
not ( n260401 , n260400 );
or ( n260402 , n260395 , n260401 );
or ( n260403 , n260400 , n37715 );
nand ( n260404 , n260402 , n260403 );
not ( n260405 , n260404 );
nand ( n260406 , n260394 , n260405 );
or ( n260407 , n260376 , n260406 );
not ( n260408 , n260405 );
not ( n260409 , n260374 );
or ( n260410 , n260408 , n260409 );
nor ( n260411 , n260394 , n47173 );
nand ( n260412 , n260410 , n260411 );
nand ( n260413 , n255116 , n204691 );
nand ( n260414 , n260407 , n260412 , n260413 );
buf ( n260415 , n260414 );
not ( n260416 , n260055 );
nor ( n260417 , n246028 , n243793 );
not ( n260418 , n260417 );
not ( n260419 , n243792 );
nand ( n260420 , n260419 , n246028 );
nand ( n260421 , n260418 , n260420 );
buf ( n260422 , n246705 );
and ( n260423 , n260421 , n260422 );
not ( n260424 , n260421 );
and ( n260425 , n260424 , n246065 );
nor ( n260426 , n260423 , n260425 );
nand ( n260427 , n260416 , n260426 );
or ( n260428 , n260427 , n260044 );
nor ( n260429 , n260043 , n252070 );
nand ( n260430 , n260429 , n260427 );
nand ( n260431 , n246460 , n38419 );
nand ( n260432 , n260428 , n260430 , n260431 );
buf ( n260433 , n260432 );
nand ( n260434 , n254509 , n254487 );
buf ( n260435 , n246352 );
not ( n260436 , n260435 );
not ( n260437 , n44539 );
or ( n260438 , n260436 , n260437 );
or ( n260439 , n44539 , n260435 );
nand ( n260440 , n260438 , n260439 );
not ( n260441 , n260440 );
buf ( n260442 , n256742 );
not ( n260443 , n260442 );
and ( n260444 , n260441 , n260443 );
and ( n260445 , n260440 , n44761 );
nor ( n260446 , n260444 , n260445 );
not ( n260447 , n260446 );
nor ( n260448 , n260447 , n237358 );
not ( n260449 , n260448 );
or ( n260450 , n260434 , n260449 );
nor ( n260451 , n260446 , n43968 );
nand ( n260452 , n260451 , n260434 );
nand ( n260453 , n231444 , n35259 );
nand ( n260454 , n260450 , n260452 , n260453 );
buf ( n260455 , n260454 );
not ( n260456 , RI19ab4dd0_2417);
or ( n260457 , n25328 , n260456 );
or ( n260458 , n25336 , n259241 );
nand ( n260459 , n260457 , n260458 );
buf ( n260460 , n260459 );
not ( n260461 , n259031 );
not ( n260462 , n225829 );
not ( n260463 , n260462 );
not ( n260464 , n226557 );
or ( n260465 , n260463 , n260464 );
not ( n260466 , n260462 );
nand ( n260467 , n260466 , n48804 );
nand ( n260468 , n260465 , n260467 );
and ( n260469 , n260468 , n259388 );
not ( n260470 , n260468 );
not ( n260471 , n259388 );
and ( n260472 , n260470 , n260471 );
nor ( n260473 , n260469 , n260472 );
not ( n260474 , n260473 );
nand ( n260475 , n260461 , n260474 );
or ( n260476 , n259010 , n260475 );
not ( n260477 , n260461 );
not ( n260478 , n259008 );
or ( n260479 , n260477 , n260478 );
nor ( n260480 , n260474 , n43517 );
nand ( n260481 , n260479 , n260480 );
nand ( n260482 , n244987 , n38889 );
nand ( n260483 , n260476 , n260481 , n260482 );
buf ( n260484 , n260483 );
not ( n260485 , n253041 );
not ( n260486 , n260485 );
not ( n260487 , n244704 );
or ( n260488 , n260486 , n260487 );
not ( n260489 , n260485 );
nand ( n260490 , n260489 , n244711 );
nand ( n260491 , n260488 , n260490 );
not ( n260492 , n260491 );
not ( n260493 , n244778 );
and ( n260494 , n260492 , n260493 );
and ( n260495 , n260491 , n244778 );
nor ( n260496 , n260494 , n260495 );
nand ( n260497 , n260496 , n254227 );
not ( n260498 , n53242 );
not ( n260499 , n256765 );
or ( n260500 , n260498 , n260499 );
not ( n260501 , n53242 );
nand ( n260502 , n260501 , n253673 );
nand ( n260503 , n260500 , n260502 );
and ( n260504 , n260503 , n253679 );
not ( n260505 , n260503 );
and ( n260506 , n260505 , n253676 );
nor ( n260507 , n260504 , n260506 );
not ( n260508 , n251800 );
not ( n260509 , n258512 );
or ( n260510 , n260508 , n260509 );
not ( n260511 , n251800 );
nand ( n260512 , n260511 , n259214 );
nand ( n260513 , n260510 , n260512 );
not ( n260514 , n257147 );
not ( n260515 , n50192 );
nand ( n260516 , n260515 , n235936 );
and ( n260517 , n260516 , n50203 );
not ( n260518 , n260516 );
and ( n260519 , n260518 , n50202 );
nor ( n260520 , n260517 , n260519 );
not ( n260521 , n260520 );
and ( n260522 , n260514 , n260521 );
and ( n260523 , n257147 , n260520 );
nor ( n260524 , n260522 , n260523 );
not ( n260525 , n260524 );
not ( n260526 , n227838 );
nand ( n260527 , n50154 , n236006 );
not ( n260528 , n260527 );
not ( n260529 , n50146 );
and ( n260530 , n260528 , n260529 );
and ( n260531 , n260527 , n50146 );
nor ( n260532 , n260530 , n260531 );
not ( n260533 , n260532 );
or ( n260534 , n260526 , n260533 );
or ( n260535 , n260532 , n227838 );
nand ( n260536 , n260534 , n260535 );
nand ( n260537 , n236028 , n236044 );
buf ( n260538 , n227862 );
xnor ( n260539 , n260537 , n260538 );
and ( n260540 , n260536 , n260539 );
not ( n260541 , n260536 );
not ( n260542 , n260539 );
and ( n260543 , n260541 , n260542 );
nor ( n260544 , n260540 , n260543 );
not ( n260545 , n260544 );
or ( n260546 , n260525 , n260545 );
not ( n260547 , n260544 );
not ( n260548 , n260524 );
nand ( n260549 , n260547 , n260548 );
nand ( n260550 , n260546 , n260549 );
buf ( n260551 , n260550 );
and ( n260552 , n260513 , n260551 );
not ( n260553 , n260513 );
and ( n260554 , n260547 , n260548 );
not ( n260555 , n260547 );
and ( n260556 , n260555 , n260524 );
nor ( n260557 , n260554 , n260556 );
buf ( n260558 , n260557 );
and ( n260559 , n260553 , n260558 );
nor ( n260560 , n260552 , n260559 );
not ( n260561 , n260560 );
nand ( n260562 , n260507 , n260561 );
or ( n260563 , n260497 , n260562 );
not ( n260564 , n260507 );
not ( n260565 , n260496 );
or ( n260566 , n260564 , n260565 );
not ( n260567 , n241373 );
nor ( n260568 , n260561 , n260567 );
nand ( n260569 , n260566 , n260568 );
nand ( n260570 , n35431 , n205267 );
nand ( n260571 , n260563 , n260569 , n260570 );
buf ( n260572 , n260571 );
not ( n260573 , n245306 );
not ( n260574 , n252235 );
or ( n260575 , n260573 , n260574 );
not ( n260576 , n245306 );
nand ( n260577 , n260576 , n252236 );
nand ( n260578 , n260575 , n260577 );
and ( n260579 , n260578 , n252239 );
not ( n260580 , n260578 );
and ( n260581 , n260580 , n252242 );
nor ( n260582 , n260579 , n260581 );
not ( n260583 , n260582 );
nand ( n260584 , n260583 , n253902 );
not ( n260585 , n252308 );
not ( n260586 , n243959 );
or ( n260587 , n260585 , n260586 );
not ( n260588 , n252308 );
nand ( n260589 , n260588 , n243953 );
nand ( n260590 , n260587 , n260589 );
and ( n260591 , n260590 , n250275 );
not ( n260592 , n260590 );
and ( n260593 , n260592 , n250272 );
nor ( n260594 , n260591 , n260593 );
not ( n260595 , n259756 );
not ( n260596 , n225920 );
not ( n260597 , n48227 );
or ( n260598 , n260596 , n260597 );
or ( n260599 , n48227 , n225920 );
nand ( n260600 , n260598 , n260599 );
not ( n260601 , n247601 );
nor ( n260602 , n260600 , n260601 );
not ( n260603 , n260602 );
nand ( n260604 , n260600 , n260601 );
nand ( n260605 , n260603 , n260604 );
not ( n260606 , n260605 );
and ( n260607 , n260595 , n260606 );
and ( n260608 , n253578 , n260605 );
nor ( n260609 , n260607 , n260608 );
nand ( n260610 , n260594 , n260609 );
or ( n260611 , n260584 , n260610 );
not ( n260612 , n260594 );
not ( n260613 , n260583 );
or ( n260614 , n260612 , n260613 );
nor ( n260615 , n260609 , n237384 );
nand ( n260616 , n260614 , n260615 );
nand ( n260617 , n234453 , n30474 );
nand ( n260618 , n260611 , n260616 , n260617 );
buf ( n260619 , n260618 );
not ( n260620 , n235149 );
not ( n260621 , n248455 );
or ( n260622 , n260620 , n260621 );
or ( n260623 , n248455 , n235149 );
nand ( n260624 , n260622 , n260623 );
not ( n260625 , n248386 );
and ( n260626 , n260624 , n260625 );
not ( n260627 , n260624 );
and ( n260628 , n260627 , n248386 );
nor ( n260629 , n260626 , n260628 );
not ( n260630 , n260629 );
nor ( n260631 , n260630 , n52445 );
not ( n260632 , n260631 );
buf ( n260633 , n250991 );
and ( n260634 , n260633 , n245114 );
not ( n260635 , n260633 );
not ( n260636 , n245072 );
not ( n260637 , n245105 );
and ( n260638 , n260636 , n260637 );
and ( n260639 , n245072 , n245105 );
nor ( n260640 , n260638 , n260639 );
and ( n260641 , n260635 , n260640 );
or ( n260642 , n260634 , n260641 );
not ( n260643 , n260642 );
not ( n260644 , n245171 );
not ( n260645 , n260644 );
and ( n260646 , n260643 , n260645 );
not ( n260647 , n245171 );
and ( n260648 , n260642 , n260647 );
nor ( n260649 , n260646 , n260648 );
not ( n260650 , n247912 );
not ( n260651 , n239858 );
or ( n260652 , n260650 , n260651 );
nand ( n260653 , n239854 , n247913 );
nand ( n260654 , n260652 , n260653 );
and ( n260655 , n260654 , n239931 );
not ( n260656 , n260654 );
and ( n260657 , n260656 , n239924 );
nor ( n260658 , n260655 , n260657 );
nand ( n260659 , n260649 , n260658 );
or ( n260660 , n260632 , n260659 );
not ( n260661 , n260658 );
not ( n260662 , n260629 );
or ( n260663 , n260661 , n260662 );
nor ( n260664 , n260649 , n235732 );
nand ( n260665 , n260663 , n260664 );
nand ( n260666 , n244789 , n30985 );
nand ( n260667 , n260660 , n260665 , n260666 );
buf ( n260668 , n260667 );
nand ( n260669 , n249971 , n223839 );
not ( n260670 , n241647 );
not ( n260671 , n243363 );
or ( n260672 , n260670 , n260671 );
not ( n260673 , n241647 );
nand ( n260674 , n260673 , n243372 );
nand ( n260675 , n260672 , n260674 );
and ( n260676 , n260675 , n256069 );
not ( n260677 , n260675 );
and ( n260678 , n260677 , n246694 );
nor ( n260679 , n260676 , n260678 );
not ( n260680 , n247119 );
not ( n260681 , n240124 );
not ( n260682 , n255992 );
or ( n260683 , n260681 , n260682 );
or ( n260684 , n256695 , n240124 );
nand ( n260685 , n260683 , n260684 );
not ( n260686 , n260685 );
or ( n260687 , n260680 , n260686 );
or ( n260688 , n255998 , n260685 );
nand ( n260689 , n260687 , n260688 );
not ( n260690 , n260689 );
nand ( n260691 , n260679 , n260690 );
or ( n260692 , n260669 , n260691 );
not ( n260693 , n260690 );
not ( n260694 , n249971 );
or ( n260695 , n260693 , n260694 );
nor ( n260696 , n260679 , n255014 );
nand ( n260697 , n260695 , n260696 );
nand ( n260698 , n234024 , n42272 );
nand ( n260699 , n260692 , n260697 , n260698 );
buf ( n260700 , n260699 );
not ( n260701 , n35141 );
not ( n260702 , n37728 );
or ( n260703 , n260701 , n260702 );
nand ( n260704 , n254406 , n254410 );
not ( n260705 , n241170 );
not ( n260706 , n235728 );
or ( n260707 , n260705 , n260706 );
not ( n260708 , n241170 );
nand ( n260709 , n260708 , n235718 );
nand ( n260710 , n260707 , n260709 );
buf ( n260711 , n236502 );
not ( n260712 , n260711 );
and ( n260713 , n260710 , n260712 );
not ( n260714 , n260710 );
and ( n260715 , n260714 , n260711 );
nor ( n260716 , n260713 , n260715 );
not ( n260717 , n260716 );
and ( n260718 , n260704 , n260717 );
not ( n260719 , n260704 );
and ( n260720 , n260719 , n260716 );
nor ( n260721 , n260718 , n260720 );
or ( n260722 , n260721 , n254882 );
nand ( n260723 , n260703 , n260722 );
buf ( n260724 , n260723 );
not ( n260725 , n30526 );
not ( n260726 , n50615 );
or ( n260727 , n260725 , n260726 );
not ( n260728 , n49355 );
not ( n260729 , n247119 );
or ( n260730 , n260728 , n260729 );
not ( n260731 , n49355 );
nand ( n260732 , n260731 , n247126 );
nand ( n260733 , n260730 , n260732 );
and ( n260734 , n260733 , n247250 );
not ( n260735 , n260733 );
and ( n260736 , n260735 , n247196 );
nor ( n260737 , n260734 , n260736 );
buf ( n260738 , n44080 );
not ( n260739 , n260738 );
not ( n260740 , n255320 );
or ( n260741 , n260739 , n260740 );
or ( n260742 , n255320 , n260738 );
nand ( n260743 , n260741 , n260742 );
not ( n260744 , n260743 );
not ( n260745 , n234098 );
and ( n260746 , n260744 , n260745 );
and ( n260747 , n260743 , n234098 );
nor ( n260748 , n260746 , n260747 );
nand ( n260749 , n260737 , n260748 );
not ( n260750 , n260749 );
not ( n260751 , n227548 );
xor ( n260752 , n242491 , n260751 );
not ( n260753 , n253377 );
xor ( n260754 , n260752 , n260753 );
not ( n260755 , n260754 );
not ( n260756 , n260755 );
and ( n260757 , n260750 , n260756 );
and ( n260758 , n260749 , n260755 );
nor ( n260759 , n260757 , n260758 );
buf ( n260760 , n52445 );
or ( n260761 , n260759 , n260760 );
nand ( n260762 , n260727 , n260761 );
buf ( n260763 , n260762 );
not ( n260764 , n205649 );
not ( n260765 , n234087 );
not ( n260766 , n38222 );
or ( n260767 , n260765 , n260766 );
not ( n260768 , n234087 );
nand ( n260769 , n260768 , n38232 );
nand ( n260770 , n260767 , n260769 );
and ( n260771 , n260770 , n38634 );
not ( n260772 , n260770 );
and ( n260773 , n260772 , n38625 );
nor ( n260774 , n260771 , n260773 );
nor ( n260775 , n260764 , n260774 );
nor ( n260776 , n257822 , n257834 );
nand ( n260777 , n260775 , n260776 );
not ( n260778 , n257833 );
not ( n260779 , n260774 );
not ( n260780 , n260779 );
or ( n260781 , n260778 , n260780 );
nor ( n260782 , n257823 , n234021 );
nand ( n260783 , n260781 , n260782 );
nand ( n260784 , n241378 , n32615 );
nand ( n260785 , n260777 , n260783 , n260784 );
buf ( n260786 , n260785 );
not ( n260787 , RI19aa0b50_2563);
or ( n260788 , n25328 , n260787 );
not ( n260789 , RI19a97028_2633);
or ( n260790 , n25336 , n260789 );
nand ( n260791 , n260788 , n260790 );
buf ( n260792 , n260791 );
not ( n260793 , n252815 );
not ( n260794 , n50940 );
or ( n260795 , n260793 , n260794 );
not ( n260796 , n252815 );
nand ( n260797 , n260796 , n50930 );
nand ( n260798 , n260795 , n260797 );
and ( n260799 , n260798 , n244532 );
not ( n260800 , n260798 );
and ( n260801 , n260800 , n244529 );
nor ( n260802 , n260799 , n260801 );
nor ( n260803 , n260802 , n52445 );
not ( n260804 , n234502 );
not ( n260805 , n234121 );
or ( n260806 , n260804 , n260805 );
not ( n260807 , n49043 );
or ( n260808 , n260807 , n234502 );
nand ( n260809 , n260806 , n260808 );
not ( n260810 , n260809 );
not ( n260811 , n234186 );
and ( n260812 , n260810 , n260811 );
and ( n260813 , n260809 , n248154 );
nor ( n260814 , n260812 , n260813 );
not ( n260815 , n260814 );
not ( n260816 , n226084 );
not ( n260817 , n260816 );
not ( n260818 , n254947 );
or ( n260819 , n260817 , n260818 );
not ( n260820 , n260816 );
nand ( n260821 , n260820 , n254946 );
nand ( n260822 , n260819 , n260821 );
not ( n260823 , n254974 );
and ( n260824 , n260822 , n260823 );
not ( n260825 , n260822 );
and ( n260826 , n260825 , n254974 );
nor ( n260827 , n260824 , n260826 );
nor ( n260828 , n260815 , n260827 );
nand ( n260829 , n260803 , n260828 );
not ( n260830 , n260827 );
not ( n260831 , n260830 );
not ( n260832 , n260802 );
not ( n260833 , n260832 );
or ( n260834 , n260831 , n260833 );
nor ( n260835 , n260814 , n50944 );
nand ( n260836 , n260834 , n260835 );
nand ( n260837 , n35431 , n38126 );
nand ( n260838 , n260829 , n260836 , n260837 );
buf ( n260839 , n260838 );
not ( n260840 , n34276 );
not ( n260841 , n244789 );
or ( n260842 , n260840 , n260841 );
not ( n260843 , n54152 );
not ( n260844 , n242380 );
or ( n260845 , n260843 , n260844 );
not ( n260846 , n54152 );
nand ( n260847 , n260846 , n242373 );
nand ( n260848 , n260845 , n260847 );
and ( n260849 , n260848 , n243660 );
not ( n260850 , n260848 );
and ( n260851 , n260850 , n243659 );
nor ( n260852 , n260849 , n260851 );
not ( n260853 , n260852 );
nand ( n260854 , n238411 , n260853 );
not ( n260855 , n260854 );
not ( n260856 , n238478 );
not ( n260857 , n260856 );
and ( n260858 , n260855 , n260857 );
and ( n260859 , n260854 , n260856 );
nor ( n260860 , n260858 , n260859 );
buf ( n260861 , n260567 );
or ( n260862 , n260860 , n260861 );
nand ( n260863 , n260842 , n260862 );
buf ( n260864 , n260863 );
not ( n260865 , n253056 );
not ( n260866 , n244704 );
or ( n260867 , n260865 , n260866 );
not ( n260868 , n253056 );
nand ( n260869 , n260868 , n244711 );
nand ( n260870 , n260867 , n260869 );
not ( n260871 , n260870 );
not ( n260872 , n244778 );
and ( n260873 , n260871 , n260872 );
and ( n260874 , n260870 , n244778 );
nor ( n260875 , n260873 , n260874 );
nand ( n260876 , n260875 , n256811 );
or ( n260877 , n260876 , n237735 );
not ( n260878 , n260875 );
not ( n260879 , n249531 );
nand ( n260880 , n260878 , n260879 );
not ( n260881 , n260880 );
not ( n260882 , n237657 );
not ( n260883 , n233997 );
or ( n260884 , n260882 , n260883 );
not ( n260885 , n237657 );
nand ( n260886 , n260885 , n44176 );
nand ( n260887 , n260884 , n260886 );
and ( n260888 , n260887 , n44325 );
not ( n260889 , n260887 );
and ( n260890 , n260889 , n44316 );
nor ( n260891 , n260888 , n260890 );
not ( n260892 , n260891 );
nand ( n260893 , n260892 , n237735 );
not ( n260894 , n260893 );
and ( n260895 , n260881 , n260894 );
and ( n260896 , n245221 , n205036 );
nor ( n260897 , n260895 , n260896 );
nand ( n260898 , n237736 , n260891 );
nand ( n260899 , n260877 , n260897 , n260898 );
buf ( n260900 , n260899 );
not ( n260901 , RI19ac7f70_2270);
or ( n260902 , n226819 , n260901 );
or ( n260903 , n25336 , n256302 );
nand ( n260904 , n260902 , n260903 );
buf ( n260905 , n260904 );
or ( n260906 , n25328 , n245696 );
not ( n260907 , RI19a82790_2777);
or ( n260908 , n226822 , n260907 );
nand ( n260909 , n260906 , n260908 );
buf ( n260910 , n260909 );
not ( n260911 , n253103 );
nand ( n260912 , n260911 , n235051 );
not ( n260913 , n260912 );
nand ( n260914 , n253118 , n250694 );
not ( n260915 , n260914 );
and ( n260916 , n260913 , n260915 );
and ( n260917 , n245702 , n40867 );
nor ( n260918 , n260916 , n260917 );
not ( n260919 , n253104 );
nand ( n260920 , n260919 , n250727 );
nand ( n260921 , n250695 , n253117 );
nand ( n260922 , n260918 , n260920 , n260921 );
buf ( n260923 , n260922 );
not ( n260924 , RI19ab1ba8_2441);
or ( n260925 , n25328 , n260924 );
not ( n260926 , RI19aa7c48_2511);
or ( n260927 , n25335 , n260926 );
nand ( n260928 , n260925 , n260927 );
buf ( n260929 , n260928 );
not ( n260930 , n253904 );
nand ( n260931 , n55780 , n260930 );
or ( n260932 , n260931 , n256408 );
and ( n260933 , n234441 , n55780 );
and ( n260934 , n30625 , n35431 );
nor ( n260935 , n260933 , n260934 );
nand ( n260936 , n234446 , n55781 , n256408 );
nand ( n260937 , n260932 , n260935 , n260936 );
buf ( n260938 , n260937 );
nor ( n260939 , n233959 , n233192 );
not ( n260940 , n260939 );
nand ( n260941 , n233192 , n233959 );
nand ( n260942 , n260940 , n260941 );
and ( n260943 , n260942 , n238629 );
not ( n260944 , n260942 );
and ( n260945 , n260944 , n238621 );
nor ( n260946 , n260943 , n260945 );
nand ( n260947 , n260946 , n241459 );
not ( n260948 , n55289 );
not ( n260949 , n260948 );
not ( n260950 , n53080 );
or ( n260951 , n260949 , n260950 );
not ( n260952 , n260948 );
nand ( n260953 , n260952 , n255385 );
nand ( n260954 , n260951 , n260953 );
and ( n260955 , n260954 , n230906 );
not ( n260956 , n260954 );
buf ( n260957 , n249298 );
and ( n260958 , n260956 , n260957 );
nor ( n260959 , n260955 , n260958 );
not ( n260960 , n248601 );
not ( n260961 , n251845 );
or ( n260962 , n260960 , n260961 );
not ( n260963 , n248601 );
nand ( n260964 , n260963 , n251855 );
nand ( n260965 , n260962 , n260964 );
buf ( n260966 , n236055 );
not ( n260967 , n260966 );
and ( n260968 , n260965 , n260967 );
not ( n260969 , n260965 );
and ( n260970 , n260969 , n260966 );
nor ( n260971 , n260968 , n260970 );
not ( n260972 , n260971 );
nand ( n260973 , n260959 , n260972 );
or ( n260974 , n260947 , n260973 );
nor ( n260975 , n260946 , n38637 );
nand ( n260976 , n260975 , n260973 );
nand ( n260977 , n31576 , n204496 );
nand ( n260978 , n260974 , n260976 , n260977 );
buf ( n260979 , n260978 );
not ( n260980 , n204650 );
not ( n260981 , n245701 );
or ( n260982 , n260980 , n260981 );
not ( n260983 , n246302 );
not ( n260984 , n260983 );
not ( n260985 , n244116 );
not ( n260986 , n260985 );
or ( n260987 , n260984 , n260986 );
not ( n260988 , n260983 );
nand ( n260989 , n260988 , n244116 );
nand ( n260990 , n260987 , n260989 );
and ( n260991 , n260990 , n239654 );
not ( n260992 , n260990 );
and ( n260993 , n260992 , n244127 );
nor ( n260994 , n260991 , n260993 );
not ( n260995 , n260994 );
not ( n260996 , n52430 );
not ( n260997 , n248056 );
or ( n260998 , n260996 , n260997 );
not ( n260999 , n52430 );
nand ( n261000 , n260999 , n248055 );
nand ( n261001 , n260998 , n261000 );
xor ( n261002 , n261001 , n248063 );
nand ( n261003 , n260995 , n261002 );
and ( n261004 , n261003 , n256969 );
not ( n261005 , n261003 );
not ( n261006 , n256969 );
and ( n261007 , n261005 , n261006 );
nor ( n261008 , n261004 , n261007 );
not ( n261009 , n205649 );
or ( n261010 , n261008 , n261009 );
nand ( n261011 , n260982 , n261010 );
buf ( n261012 , n261011 );
not ( n261013 , RI19aa27e8_2549);
or ( n261014 , n25328 , n261013 );
not ( n261015 , RI19a98f90_2619);
or ( n261016 , n25336 , n261015 );
nand ( n261017 , n261014 , n261016 );
buf ( n261018 , n261017 );
not ( n261019 , RI19abeda8_2342);
or ( n261020 , n25328 , n261019 );
not ( n261021 , RI19ab5820_2412);
or ( n261022 , n226822 , n261021 );
nand ( n261023 , n261020 , n261022 );
buf ( n261024 , n261023 );
not ( n261025 , n44909 );
not ( n261026 , n31577 );
or ( n261027 , n261025 , n261026 );
not ( n261028 , n245510 );
not ( n261029 , n241893 );
or ( n261030 , n261028 , n261029 );
or ( n261031 , n55067 , n245510 );
nand ( n261032 , n261030 , n261031 );
not ( n261033 , n261032 );
not ( n261034 , n241963 );
or ( n261035 , n261033 , n261034 );
not ( n261036 , n241962 );
not ( n261037 , n261036 );
or ( n261038 , n261037 , n261032 );
nand ( n261039 , n261035 , n261038 );
not ( n261040 , n258512 );
not ( n261041 , n243598 );
not ( n261042 , n254728 );
or ( n261043 , n261041 , n261042 );
or ( n261044 , n254728 , n243598 );
nand ( n261045 , n261043 , n261044 );
not ( n261046 , n261045 );
and ( n261047 , n261040 , n261046 );
and ( n261048 , n259218 , n261045 );
nor ( n261049 , n261047 , n261048 );
nand ( n261050 , n261039 , n261049 );
not ( n261051 , n261050 );
not ( n261052 , n234233 );
not ( n261053 , n41929 );
or ( n261054 , n261052 , n261053 );
not ( n261055 , n234233 );
nand ( n261056 , n261055 , n41933 );
nand ( n261057 , n261054 , n261056 );
buf ( n261058 , n43725 );
and ( n261059 , n261057 , n261058 );
not ( n261060 , n261057 );
and ( n261061 , n261060 , n259105 );
nor ( n261062 , n261059 , n261061 );
not ( n261063 , n261062 );
not ( n261064 , n261063 );
and ( n261065 , n261051 , n261064 );
and ( n261066 , n261050 , n261063 );
nor ( n261067 , n261065 , n261066 );
or ( n261068 , n261067 , n55108 );
nand ( n261069 , n261027 , n261068 );
buf ( n261070 , n261069 );
not ( n261071 , n236708 );
not ( n261072 , n43219 );
or ( n261073 , n261071 , n261072 );
or ( n261074 , n43219 , n236708 );
nand ( n261075 , n261073 , n261074 );
not ( n261076 , n45023 );
buf ( n261077 , n261076 );
and ( n261078 , n261075 , n261077 );
not ( n261079 , n261075 );
and ( n261080 , n261079 , n45027 );
nor ( n261081 , n261078 , n261080 );
nor ( n261082 , n261081 , n55332 );
nand ( n261083 , n55513 , n50945 );
or ( n261084 , n261082 , n261083 );
nand ( n261085 , n233496 , n261082 );
nand ( n261086 , n239240 , n39833 );
nand ( n261087 , n261084 , n261085 , n261086 );
buf ( n261088 , n261087 );
not ( n261089 , n37042 );
not ( n261090 , n55760 );
or ( n261091 , n261089 , n261090 );
not ( n261092 , n52878 );
not ( n261093 , n246882 );
or ( n261094 , n261092 , n261093 );
not ( n261095 , n52878 );
nand ( n261096 , n261095 , n246891 );
nand ( n261097 , n261094 , n261096 );
and ( n261098 , n261097 , n260340 );
not ( n261099 , n261097 );
and ( n261100 , n261099 , n258077 );
nor ( n261101 , n261098 , n261100 );
not ( n261102 , n237907 );
not ( n261103 , n261102 );
not ( n261104 , n246767 );
or ( n261105 , n261103 , n261104 );
not ( n261106 , n261102 );
nand ( n261107 , n261106 , n246759 );
nand ( n261108 , n261105 , n261107 );
and ( n261109 , n261108 , n254010 );
not ( n261110 , n261108 );
and ( n261111 , n261110 , n254006 );
nor ( n261112 , n261109 , n261111 );
nand ( n261113 , n261101 , n261112 );
and ( n261114 , n261113 , n259113 );
not ( n261115 , n261113 );
not ( n261116 , n259113 );
and ( n261117 , n261115 , n261116 );
nor ( n261118 , n261114 , n261117 );
or ( n261119 , n261118 , n46425 );
nand ( n261120 , n261091 , n261119 );
buf ( n261121 , n261120 );
not ( n261122 , n254286 );
not ( n261123 , n261122 );
not ( n261124 , n251029 );
or ( n261125 , n261123 , n261124 );
not ( n261126 , n261122 );
not ( n261127 , n251028 );
nand ( n261128 , n261126 , n261127 );
nand ( n261129 , n261125 , n261128 );
buf ( n261130 , n47310 );
and ( n261131 , n261129 , n261130 );
not ( n261132 , n261129 );
buf ( n261133 , n47319 );
and ( n261134 , n261132 , n261133 );
nor ( n261135 , n261131 , n261134 );
not ( n261136 , n249419 );
not ( n261137 , n261136 );
not ( n261138 , n38633 );
or ( n261139 , n261137 , n261138 );
not ( n261140 , n261136 );
nand ( n261141 , n261140 , n38625 );
nand ( n261142 , n261139 , n261141 );
and ( n261143 , n261142 , n49182 );
not ( n261144 , n261142 );
and ( n261145 , n261144 , n49191 );
nor ( n261146 , n261143 , n261145 );
not ( n261147 , n261146 );
nand ( n261148 , n261135 , n261147 );
not ( n261149 , n239286 );
not ( n261150 , n248755 );
or ( n261151 , n261149 , n261150 );
not ( n261152 , n239286 );
nand ( n261153 , n261152 , n248762 );
nand ( n261154 , n261151 , n261153 );
and ( n261155 , n261154 , n252924 );
not ( n261156 , n261154 );
and ( n261157 , n261156 , n252923 );
nor ( n261158 , n261155 , n261157 );
not ( n261159 , n261158 );
nor ( n261160 , n261159 , n236795 );
not ( n261161 , n261160 );
or ( n261162 , n261148 , n261161 );
nor ( n261163 , n261158 , n259801 );
nand ( n261164 , n261148 , n261163 );
nand ( n261165 , n31577 , n34358 );
nand ( n261166 , n261162 , n261164 , n261165 );
buf ( n261167 , n261166 );
buf ( n261168 , n33641 );
buf ( n261169 , n204452 );
not ( n261170 , n258576 );
not ( n261171 , n40460 );
or ( n261172 , n261170 , n261171 );
not ( n261173 , n258576 );
nand ( n261174 , n261173 , n251345 );
nand ( n261175 , n261172 , n261174 );
buf ( n261176 , n241657 );
not ( n261177 , n261176 );
and ( n261178 , n261175 , n261177 );
not ( n261179 , n261175 );
and ( n261180 , n261179 , n253378 );
nor ( n261181 , n261178 , n261180 );
nand ( n261182 , n261181 , n254227 );
buf ( n261183 , n256837 );
not ( n261184 , n261183 );
not ( n261185 , n30968 );
not ( n261186 , n261185 );
or ( n261187 , n261184 , n261186 );
or ( n261188 , n208725 , n261183 );
nand ( n261189 , n261187 , n261188 );
and ( n261190 , n261189 , n31552 );
not ( n261191 , n261189 );
and ( n261192 , n261191 , n31561 );
nor ( n261193 , n261190 , n261192 );
not ( n261194 , n53609 );
not ( n261195 , n261194 );
not ( n261196 , n250496 );
or ( n261197 , n261195 , n261196 );
nand ( n261198 , n255291 , n53609 );
nand ( n261199 , n261197 , n261198 );
and ( n261200 , n261199 , n244190 );
not ( n261201 , n261199 );
and ( n261202 , n261201 , n260370 );
nor ( n261203 , n261200 , n261202 );
nor ( n261204 , n261193 , n261203 );
or ( n261205 , n261182 , n261204 );
nor ( n261206 , n261193 , n31571 );
nor ( n261207 , n261203 , n261181 );
nand ( n261208 , n261206 , n261207 );
nand ( n261209 , n247585 , n37630 );
nand ( n261210 , n261205 , n261208 , n261209 );
buf ( n261211 , n261210 );
not ( n261212 , n30093 );
not ( n261213 , n254441 );
or ( n261214 , n261212 , n261213 );
nand ( n261215 , n257436 , n257420 );
and ( n261216 , n261215 , n255602 );
not ( n261217 , n261215 );
and ( n261218 , n261217 , n255601 );
nor ( n261219 , n261216 , n261218 );
or ( n261220 , n261219 , n251498 );
nand ( n261221 , n261214 , n261220 );
buf ( n261222 , n261221 );
or ( n261223 , n25328 , n248825 );
not ( n261224 , RI19aa48b8_2533);
or ( n261225 , n226822 , n261224 );
nand ( n261226 , n261223 , n261225 );
buf ( n261227 , n261226 );
not ( n261228 , n253817 );
nand ( n261229 , n261228 , n55147 );
not ( n261230 , n233768 );
not ( n261231 , n238182 );
or ( n261232 , n261230 , n261231 );
not ( n261233 , n233768 );
nand ( n261234 , n261233 , n251217 );
nand ( n261235 , n261232 , n261234 );
and ( n261236 , n261235 , n251220 );
not ( n261237 , n261235 );
and ( n261238 , n261237 , n251224 );
nor ( n261239 , n261236 , n261238 );
nand ( n261240 , n253878 , n261239 );
or ( n261241 , n261229 , n261240 );
not ( n261242 , n253878 );
not ( n261243 , n261228 );
or ( n261244 , n261242 , n261243 );
not ( n261245 , n205649 );
nor ( n261246 , n261245 , n261239 );
nand ( n261247 , n261244 , n261246 );
nand ( n261248 , n253486 , n25556 );
nand ( n261249 , n261241 , n261247 , n261248 );
buf ( n261250 , n261249 );
not ( n261251 , RI19acd358_2230);
or ( n261252 , n25328 , n261251 );
not ( n261253 , RI19ac46b8_2296);
or ( n261254 , n25335 , n261253 );
nand ( n261255 , n261252 , n261254 );
buf ( n261256 , n261255 );
not ( n261257 , n242184 );
not ( n261258 , n27876 );
or ( n261259 , n261257 , n261258 );
not ( n261260 , n242184 );
nand ( n261261 , n261260 , n27869 );
nand ( n261262 , n261259 , n261261 );
and ( n261263 , n261262 , n248763 );
not ( n261264 , n261262 );
and ( n261265 , n261264 , n248756 );
nor ( n261266 , n261263 , n261265 );
not ( n261267 , n251029 );
not ( n261268 , n236157 );
not ( n261269 , n256950 );
not ( n261270 , n261269 );
or ( n261271 , n261268 , n261270 );
not ( n261272 , n236157 );
nand ( n261273 , n261272 , n251082 );
nand ( n261274 , n261271 , n261273 );
not ( n261275 , n261274 );
and ( n261276 , n261267 , n261275 );
and ( n261277 , n251029 , n261274 );
nor ( n261278 , n261276 , n261277 );
nor ( n261279 , n261266 , n261278 );
or ( n261280 , n261279 , n259848 );
nor ( n261281 , n259846 , n235050 );
nand ( n261282 , n261279 , n261281 );
nand ( n261283 , n247744 , n33199 );
nand ( n261284 , n261280 , n261282 , n261283 );
buf ( n261285 , n261284 );
not ( n261286 , n245040 );
not ( n261287 , n231768 );
or ( n261288 , n261286 , n261287 );
not ( n261289 , n253729 );
or ( n261290 , n261289 , n245040 );
nand ( n261291 , n261288 , n261290 );
not ( n261292 , n40918 );
and ( n261293 , n261291 , n261292 );
not ( n261294 , n261291 );
not ( n261295 , n261292 );
and ( n261296 , n261294 , n261295 );
nor ( n261297 , n261293 , n261296 );
not ( n261298 , n261297 );
nand ( n261299 , n261298 , n244515 );
not ( n261300 , n261299 );
not ( n261301 , n40095 );
not ( n261302 , n235807 );
or ( n261303 , n261301 , n261302 );
not ( n261304 , n40095 );
nand ( n261305 , n261304 , n235815 );
nand ( n261306 , n261303 , n261305 );
and ( n261307 , n261306 , n235888 );
not ( n261308 , n261306 );
and ( n261309 , n261308 , n235879 );
nor ( n261310 , n261307 , n261309 );
not ( n261311 , n261310 );
not ( n261312 , n237139 );
not ( n261313 , n253072 );
or ( n261314 , n261312 , n261313 );
nand ( n261315 , n253073 , n237033 );
nand ( n261316 , n261314 , n261315 );
and ( n261317 , n261316 , n249195 );
not ( n261318 , n261316 );
and ( n261319 , n261318 , n253081 );
nor ( n261320 , n261317 , n261319 );
nand ( n261321 , n261311 , n261320 );
not ( n261322 , n261321 );
and ( n261323 , n261300 , n261322 );
and ( n261324 , n234823 , n26490 );
nor ( n261325 , n261323 , n261324 );
nand ( n261326 , n261297 , n258918 );
not ( n261327 , n261326 );
not ( n261328 , n261320 );
nand ( n261329 , n261327 , n261328 );
nor ( n261330 , n261320 , n235050 );
nand ( n261331 , n261330 , n261310 );
nand ( n261332 , n261325 , n261329 , n261331 );
buf ( n261333 , n261332 );
not ( n261334 , RI19ab2b98_2434);
or ( n261335 , n25328 , n261334 );
not ( n261336 , RI19aa8bc0_2505);
or ( n261337 , n226822 , n261336 );
nand ( n261338 , n261335 , n261337 );
buf ( n261339 , n261338 );
buf ( n261340 , n26358 );
buf ( n261341 , n33171 );
buf ( n261342 , n25578 );
buf ( n261343 , n29590 );
not ( n261344 , n250930 );
buf ( n261345 , n250886 );
not ( n261346 , n261345 );
not ( n261347 , n245950 );
or ( n261348 , n261346 , n261347 );
or ( n261349 , n245950 , n261345 );
nand ( n261350 , n261348 , n261349 );
not ( n261351 , n226319 );
and ( n261352 , n261350 , n261351 );
not ( n261353 , n261350 );
and ( n261354 , n261353 , n226319 );
nor ( n261355 , n261352 , n261354 );
nand ( n261356 , n261355 , n252259 );
not ( n261357 , n261356 );
or ( n261358 , n261344 , n261357 );
not ( n261359 , n239765 );
not ( n261360 , n261359 );
not ( n261361 , n239107 );
or ( n261362 , n261360 , n261361 );
not ( n261363 , n261359 );
nand ( n261364 , n261363 , n239099 );
nand ( n261365 , n261362 , n261364 );
and ( n261366 , n261365 , n242079 );
not ( n261367 , n261365 );
and ( n261368 , n261367 , n242080 );
nor ( n261369 , n261366 , n261368 );
nand ( n261370 , n261358 , n261369 );
nor ( n261371 , n261355 , n261369 );
and ( n261372 , n250970 , n261371 );
and ( n261373 , n234453 , n36315 );
nor ( n261374 , n261372 , n261373 );
nand ( n261375 , n261370 , n261374 );
buf ( n261376 , n261375 );
nor ( n261377 , n256000 , n43968 );
not ( n261378 , n45876 );
buf ( n261379 , n51440 );
not ( n261380 , n261379 );
not ( n261381 , n261380 );
not ( n261382 , n239653 );
or ( n261383 , n261381 , n261382 );
nand ( n261384 , n244125 , n261379 );
nand ( n261385 , n261383 , n261384 );
not ( n261386 , n261385 );
or ( n261387 , n261378 , n261386 );
or ( n261388 , n261385 , n244978 );
nand ( n261389 , n261387 , n261388 );
nand ( n261390 , n261377 , n256014 , n261389 );
not ( n261391 , n256029 );
not ( n261392 , n261389 );
or ( n261393 , n261391 , n261392 );
nor ( n261394 , n256014 , n221279 );
nand ( n261395 , n261393 , n261394 );
nand ( n261396 , n48251 , n205187 );
nand ( n261397 , n261390 , n261395 , n261396 );
buf ( n261398 , n261397 );
nand ( n261399 , n257435 , n54200 );
nand ( n261400 , n255601 , n255614 );
or ( n261401 , n261399 , n261400 );
not ( n261402 , n255601 );
not ( n261403 , n257435 );
or ( n261404 , n261402 , n261403 );
nor ( n261405 , n255614 , n27889 );
nand ( n261406 , n261404 , n261405 );
nand ( n261407 , n31577 , n40718 );
nand ( n261408 , n261401 , n261406 , n261407 );
buf ( n261409 , n261408 );
xor ( n261410 , n250631 , n240996 );
xnor ( n261411 , n261410 , n245618 );
not ( n261412 , n261411 );
nand ( n261413 , n261412 , n252858 );
not ( n261414 , n229478 );
not ( n261415 , n256862 );
or ( n261416 , n261414 , n261415 );
not ( n261417 , n229478 );
nand ( n261418 , n261417 , n256870 );
nand ( n261419 , n261416 , n261418 );
and ( n261420 , n261419 , n256878 );
not ( n261421 , n261419 );
and ( n261422 , n261421 , n256879 );
nor ( n261423 , n261420 , n261422 );
not ( n261424 , n261423 );
not ( n261425 , n45642 );
not ( n261426 , n248210 );
or ( n261427 , n261425 , n261426 );
not ( n261428 , n45642 );
nand ( n261429 , n261428 , n248219 );
nand ( n261430 , n261427 , n261429 );
buf ( n261431 , n230374 );
and ( n261432 , n261430 , n261431 );
not ( n261433 , n261430 );
buf ( n261434 , n230367 );
and ( n261435 , n261433 , n261434 );
nor ( n261436 , n261432 , n261435 );
not ( n261437 , n261436 );
nand ( n261438 , n261424 , n261437 );
or ( n261439 , n261413 , n261438 );
not ( n261440 , n261437 );
not ( n261441 , n261412 );
or ( n261442 , n261440 , n261441 );
nor ( n261443 , n261424 , n33254 );
nand ( n261444 , n261442 , n261443 );
nand ( n261445 , n246217 , n35150 );
nand ( n261446 , n261439 , n261444 , n261445 );
buf ( n261447 , n261446 );
not ( n261448 , RI19a9ff20_2569);
or ( n261449 , n25328 , n261448 );
not ( n261450 , RI19a96038_2640);
or ( n261451 , n25335 , n261450 );
nand ( n261452 , n261449 , n261451 );
buf ( n261453 , n261452 );
not ( n261454 , n248927 );
not ( n261455 , n250099 );
or ( n261456 , n261454 , n261455 );
or ( n261457 , n250102 , n248927 );
nand ( n261458 , n261456 , n261457 );
and ( n261459 , n261458 , n250108 );
not ( n261460 , n261458 );
and ( n261461 , n261460 , n250105 );
nor ( n261462 , n261459 , n261461 );
nor ( n261463 , n261462 , n55104 );
not ( n261464 , n242585 );
not ( n261465 , n236488 );
and ( n261466 , n261464 , n261465 );
and ( n261467 , n32473 , n236488 );
nor ( n261468 , n261466 , n261467 );
and ( n261469 , n261468 , n33247 );
not ( n261470 , n261468 );
buf ( n261471 , n253530 );
and ( n261472 , n261470 , n261471 );
nor ( n261473 , n261469 , n261472 );
not ( n261474 , n45727 );
not ( n261475 , n49115 );
not ( n261476 , n223266 );
or ( n261477 , n261475 , n261476 );
not ( n261478 , n49115 );
nand ( n261479 , n45506 , n261478 );
nand ( n261480 , n261477 , n261479 );
not ( n261481 , n261480 );
or ( n261482 , n261474 , n261481 );
not ( n261483 , n45727 );
not ( n261484 , n261483 );
or ( n261485 , n261480 , n261484 );
nand ( n261486 , n261482 , n261485 );
nor ( n261487 , n261473 , n261486 );
nand ( n261488 , n261463 , n261487 );
nand ( n261489 , n261473 , n205649 );
not ( n261490 , n261489 );
not ( n261491 , n261462 );
not ( n261492 , n261486 );
nand ( n261493 , n261491 , n261492 );
nand ( n261494 , n261490 , n261493 );
nand ( n261495 , n241378 , n204741 );
nand ( n261496 , n261488 , n261494 , n261495 );
buf ( n261497 , n261496 );
not ( n261498 , n254309 );
not ( n261499 , n251029 );
or ( n261500 , n261498 , n261499 );
not ( n261501 , n254309 );
nand ( n261502 , n261501 , n261127 );
nand ( n261503 , n261500 , n261502 );
and ( n261504 , n261503 , n261130 );
not ( n261505 , n261503 );
and ( n261506 , n261505 , n261133 );
nor ( n261507 , n261504 , n261506 );
not ( n261508 , n261507 );
buf ( n261509 , n51240 );
not ( n261510 , n261509 );
not ( n261511 , n255813 );
or ( n261512 , n261510 , n261511 );
or ( n261513 , n255813 , n261509 );
nand ( n261514 , n261512 , n261513 );
and ( n261515 , n261514 , n256768 );
not ( n261516 , n261514 );
and ( n261517 , n261516 , n253669 );
nor ( n261518 , n261515 , n261517 );
not ( n261519 , n261518 );
nand ( n261520 , n261508 , n261519 );
not ( n261521 , n241113 );
not ( n261522 , n235580 );
or ( n261523 , n261521 , n261522 );
not ( n261524 , n241113 );
nand ( n261525 , n261524 , n235590 );
nand ( n261526 , n261523 , n261525 );
and ( n261527 , n261526 , n235720 );
not ( n261528 , n261526 );
and ( n261529 , n261528 , n243244 );
nor ( n261530 , n261527 , n261529 );
nand ( n261531 , n261530 , n259619 );
or ( n261532 , n261520 , n261531 );
nor ( n261533 , n261530 , n244399 );
nand ( n261534 , n261533 , n261520 );
nand ( n261535 , n31576 , n205298 );
nand ( n261536 , n261532 , n261534 , n261535 );
buf ( n261537 , n261536 );
not ( n261538 , n252511 );
not ( n261539 , n249358 );
not ( n261540 , n249332 );
or ( n261541 , n261539 , n261540 );
nand ( n261542 , n261541 , n249361 );
not ( n261543 , n261542 );
or ( n261544 , n261538 , n261543 );
or ( n261545 , n261542 , n252511 );
nand ( n261546 , n261544 , n261545 );
buf ( n261547 , n260122 );
and ( n261548 , n261546 , n261547 );
not ( n261549 , n261546 );
buf ( n261550 , n260112 );
and ( n261551 , n261549 , n261550 );
nor ( n261552 , n261548 , n261551 );
not ( n261553 , n261552 );
nand ( n261554 , n261553 , n226010 );
not ( n261555 , n234057 );
not ( n261556 , n261555 );
not ( n261557 , n38222 );
or ( n261558 , n261556 , n261557 );
not ( n261559 , n261555 );
nand ( n261560 , n261559 , n38232 );
nand ( n261561 , n261558 , n261560 );
and ( n261562 , n261561 , n38634 );
not ( n261563 , n261561 );
and ( n261564 , n261563 , n38625 );
nor ( n261565 , n261562 , n261564 );
not ( n261566 , n261565 );
not ( n261567 , n243909 );
not ( n261568 , n246064 );
or ( n261569 , n261567 , n261568 );
not ( n261570 , n243909 );
nand ( n261571 , n261570 , n246705 );
nand ( n261572 , n261569 , n261571 );
and ( n261573 , n261572 , n246760 );
not ( n261574 , n261572 );
and ( n261575 , n261574 , n246768 );
nor ( n261576 , n261573 , n261575 );
not ( n261577 , n261576 );
nand ( n261578 , n261566 , n261577 );
or ( n261579 , n261554 , n261578 );
not ( n261580 , n261566 );
not ( n261581 , n261553 );
or ( n261582 , n261580 , n261581 );
nor ( n261583 , n261577 , n235895 );
nand ( n261584 , n261582 , n261583 );
buf ( n261585 , n35431 );
nand ( n261586 , n261585 , n36927 );
nand ( n261587 , n261579 , n261584 , n261586 );
buf ( n261588 , n261587 );
not ( n261589 , n29377 );
not ( n261590 , n37728 );
or ( n261591 , n261589 , n261590 );
not ( n261592 , n51274 );
nand ( n261593 , n261592 , n229112 );
not ( n261594 , n239879 );
not ( n261595 , n261594 );
not ( n261596 , n256438 );
or ( n261597 , n261595 , n261596 );
or ( n261598 , n247572 , n261594 );
nand ( n261599 , n261597 , n261598 );
and ( n261600 , n261599 , n247575 );
not ( n261601 , n261599 );
and ( n261602 , n261601 , n242696 );
nor ( n261603 , n261600 , n261602 );
and ( n261604 , n261593 , n261603 );
not ( n261605 , n261593 );
not ( n261606 , n261603 );
and ( n261607 , n261605 , n261606 );
nor ( n261608 , n261604 , n261607 );
or ( n261609 , n261608 , n49959 );
nand ( n261610 , n261591 , n261609 );
buf ( n261611 , n261610 );
or ( n261612 , n25328 , n260180 );
not ( n261613 , RI19aa9d90_2497);
or ( n261614 , n25336 , n261613 );
nand ( n261615 , n261612 , n261614 );
buf ( n261616 , n261615 );
buf ( n261617 , n204468 );
buf ( n261618 , n36960 );
buf ( n261619 , n42750 );
buf ( n261620 , n36452 );
buf ( n261621 , n34071 );
buf ( n261622 , n30681 );
not ( n261623 , n256437 );
not ( n261624 , n246412 );
not ( n261625 , n256742 );
or ( n261626 , n261624 , n261625 );
not ( n261627 , n246412 );
nand ( n261628 , n261627 , n256738 );
nand ( n261629 , n261626 , n261628 );
buf ( n261630 , n50776 );
and ( n261631 , n261629 , n261630 );
not ( n261632 , n261629 );
and ( n261633 , n261632 , n228527 );
nor ( n261634 , n261631 , n261633 );
nand ( n261635 , n256462 , n261634 );
or ( n261636 , n261623 , n261635 );
nor ( n261637 , n256435 , n236795 );
nand ( n261638 , n261637 , n261635 );
nand ( n261639 , n238638 , n36452 );
nand ( n261640 , n261636 , n261638 , n261639 );
buf ( n261641 , n261640 );
buf ( n261642 , n30920 );
or ( n261643 , n233507 , n258914 );
not ( n261644 , RI19a91e98_2669);
or ( n261645 , n226822 , n261644 );
nand ( n261646 , n261643 , n261645 );
buf ( n261647 , n261646 );
buf ( n261648 , n31421 );
buf ( n261649 , n28076 );
not ( n261650 , n204655 );
not ( n261651 , n245702 );
or ( n261652 , n261650 , n261651 );
not ( n261653 , n238431 );
not ( n261654 , n228918 );
or ( n261655 , n261653 , n261654 );
not ( n261656 , n238431 );
nand ( n261657 , n261656 , n51167 );
nand ( n261658 , n261655 , n261657 );
and ( n261659 , n261658 , n51269 );
not ( n261660 , n261658 );
and ( n261661 , n261660 , n51272 );
nor ( n261662 , n261659 , n261661 );
nand ( n261663 , n249497 , n261662 );
buf ( n261664 , n245284 );
not ( n261665 , n261664 );
not ( n261666 , n252236 );
or ( n261667 , n261665 , n261666 );
or ( n261668 , n252236 , n261664 );
nand ( n261669 , n261667 , n261668 );
and ( n261670 , n261669 , n252242 );
not ( n261671 , n261669 );
and ( n261672 , n261671 , n252239 );
nor ( n261673 , n261670 , n261672 );
not ( n261674 , n261673 );
and ( n261675 , n261663 , n261674 );
not ( n261676 , n261663 );
and ( n261677 , n261676 , n261673 );
nor ( n261678 , n261675 , n261677 );
or ( n261679 , n261678 , n254470 );
nand ( n261680 , n261652 , n261679 );
buf ( n261681 , n261680 );
not ( n261682 , n31808 );
not ( n261683 , n244789 );
or ( n261684 , n261682 , n261683 );
not ( n261685 , n248418 );
not ( n261686 , n221715 );
or ( n261687 , n261685 , n261686 );
not ( n261688 , n248418 );
nand ( n261689 , n261688 , n43962 );
nand ( n261690 , n261687 , n261689 );
and ( n261691 , n261690 , n255612 );
not ( n261692 , n261690 );
and ( n261693 , n261692 , n255609 );
nor ( n261694 , n261691 , n261693 );
not ( n261695 , n261694 );
not ( n261696 , n234913 );
not ( n261697 , n254117 );
not ( n261698 , n261697 );
or ( n261699 , n261696 , n261698 );
not ( n261700 , n234913 );
nand ( n261701 , n261700 , n254117 );
nand ( n261702 , n261699 , n261701 );
and ( n261703 , n261702 , n254122 );
not ( n261704 , n261702 );
and ( n261705 , n261704 , n254125 );
nor ( n261706 , n261703 , n261705 );
nand ( n261707 , n261695 , n261706 );
not ( n261708 , n46411 );
not ( n261709 , n248557 );
or ( n261710 , n261708 , n261709 );
not ( n261711 , n46411 );
nand ( n261712 , n261711 , n248565 );
nand ( n261713 , n261710 , n261712 );
and ( n261714 , n261713 , n248679 );
not ( n261715 , n261713 );
and ( n261716 , n261715 , n248678 );
nor ( n261717 , n261714 , n261716 );
not ( n261718 , n261717 );
and ( n261719 , n261707 , n261718 );
not ( n261720 , n261707 );
and ( n261721 , n261720 , n261717 );
nor ( n261722 , n261719 , n261721 );
or ( n261723 , n261722 , n255135 );
nand ( n261724 , n261684 , n261723 );
buf ( n261725 , n261724 );
not ( n261726 , n35065 );
not ( n261727 , n255116 );
or ( n261728 , n261726 , n261727 );
nand ( n261729 , n241887 , n241968 );
not ( n261730 , n47147 );
not ( n261731 , n252823 );
or ( n261732 , n261730 , n261731 );
not ( n261733 , n47147 );
nand ( n261734 , n261733 , n252831 );
nand ( n261735 , n261732 , n261734 );
and ( n261736 , n261735 , n252834 );
not ( n261737 , n261735 );
and ( n261738 , n261737 , n252837 );
nor ( n261739 , n261736 , n261738 );
and ( n261740 , n261729 , n261739 );
not ( n261741 , n261729 );
not ( n261742 , n261739 );
and ( n261743 , n261741 , n261742 );
nor ( n261744 , n261740 , n261743 );
or ( n261745 , n261744 , n251498 );
nand ( n261746 , n261728 , n261745 );
buf ( n261747 , n261746 );
not ( n261748 , RI19a9cc08_2592);
or ( n261749 , n25328 , n261748 );
not ( n261750 , RI19aced20_2219);
or ( n261751 , n25335 , n261750 );
nand ( n261752 , n261749 , n261751 );
buf ( n261753 , n261752 );
not ( n261754 , n39696 );
not ( n261755 , n245221 );
or ( n261756 , n261754 , n261755 );
not ( n261757 , n221138 );
not ( n261758 , n261757 );
not ( n261759 , n238894 );
or ( n261760 , n261758 , n261759 );
not ( n261761 , n261757 );
nand ( n261762 , n261761 , n246077 );
nand ( n261763 , n261760 , n261762 );
and ( n261764 , n261763 , n246082 );
not ( n261765 , n261763 );
and ( n261766 , n261765 , n244453 );
nor ( n261767 , n261764 , n261766 );
not ( n261768 , n239524 );
not ( n261769 , n260112 );
or ( n261770 , n261768 , n261769 );
not ( n261771 , n239524 );
nand ( n261772 , n261771 , n260122 );
nand ( n261773 , n261770 , n261772 );
and ( n261774 , n261773 , n237746 );
not ( n261775 , n261773 );
not ( n261776 , n260125 );
and ( n261777 , n261775 , n261776 );
nor ( n261778 , n261774 , n261777 );
nand ( n261779 , n261767 , n261778 );
and ( n261780 , n261779 , n256771 );
not ( n261781 , n261779 );
and ( n261782 , n261781 , n256770 );
nor ( n261783 , n261780 , n261782 );
or ( n261784 , n261783 , n35816 );
nand ( n261785 , n261756 , n261784 );
buf ( n261786 , n261785 );
not ( n261787 , n31573 );
not ( n261788 , n246133 );
not ( n261789 , n261788 );
not ( n261790 , n245602 );
or ( n261791 , n261789 , n261790 );
nand ( n261792 , n245611 , n246133 );
nand ( n261793 , n261791 , n261792 );
not ( n261794 , n261793 );
not ( n261795 , n245615 );
and ( n261796 , n261794 , n261795 );
and ( n261797 , n261793 , n253746 );
nor ( n261798 , n261796 , n261797 );
not ( n261799 , n241422 );
not ( n261800 , n47531 );
or ( n261801 , n261799 , n261800 );
not ( n261802 , n241422 );
nand ( n261803 , n261802 , n225301 );
nand ( n261804 , n261801 , n261803 );
and ( n261805 , n261804 , n225525 );
not ( n261806 , n261804 );
and ( n261807 , n261806 , n225536 );
nor ( n261808 , n261805 , n261807 );
nand ( n261809 , n261798 , n261808 );
or ( n261810 , n261787 , n261809 );
not ( n261811 , n261808 );
not ( n261812 , n29968 );
or ( n261813 , n261811 , n261812 );
nor ( n261814 , n261798 , n47173 );
nand ( n261815 , n261813 , n261814 );
nand ( n261816 , n31577 , n25367 );
nand ( n261817 , n261810 , n261815 , n261816 );
buf ( n261818 , n261817 );
not ( n261819 , RI19a998f0_2615);
or ( n261820 , n25328 , n261819 );
not ( n261821 , RI19a8f8a0_2686);
or ( n261822 , n25335 , n261821 );
nand ( n261823 , n261820 , n261822 );
buf ( n261824 , n261823 );
not ( n261825 , n234792 );
not ( n261826 , n242645 );
not ( n261827 , n242670 );
and ( n261828 , n261826 , n261827 );
and ( n261829 , n242645 , n242670 );
nor ( n261830 , n261828 , n261829 );
not ( n261831 , n261830 );
or ( n261832 , n261825 , n261831 );
not ( n261833 , n234792 );
not ( n261834 , n261830 );
nand ( n261835 , n261833 , n261834 );
nand ( n261836 , n261832 , n261835 );
and ( n261837 , n261836 , n242680 );
not ( n261838 , n261836 );
and ( n261839 , n261838 , n242683 );
nor ( n261840 , n261837 , n261839 );
not ( n261841 , n51307 );
not ( n261842 , n43005 );
or ( n261843 , n261841 , n261842 );
not ( n261844 , n51307 );
nand ( n261845 , n261844 , n43010 );
nand ( n261846 , n261843 , n261845 );
and ( n261847 , n261846 , n227796 );
not ( n261848 , n261846 );
and ( n261849 , n261848 , n50028 );
nor ( n261850 , n261847 , n261849 );
nand ( n261851 , n261840 , n261850 );
not ( n261852 , n238669 );
not ( n261853 , n261852 );
not ( n261854 , n247991 );
or ( n261855 , n261853 , n261854 );
not ( n261856 , n261852 );
nand ( n261857 , n261856 , n247999 );
nand ( n261858 , n261855 , n261857 );
buf ( n261859 , n247499 );
and ( n261860 , n261858 , n261859 );
not ( n261861 , n261858 );
not ( n261862 , n261859 );
and ( n261863 , n261861 , n261862 );
nor ( n261864 , n261860 , n261863 );
not ( n261865 , n261864 );
nor ( n261866 , n261865 , n234110 );
not ( n261867 , n261866 );
or ( n261868 , n261851 , n261867 );
not ( n261869 , n261864 );
not ( n261870 , n261840 );
or ( n261871 , n261869 , n261870 );
nor ( n261872 , n261850 , n40465 );
nand ( n261873 , n261871 , n261872 );
nand ( n261874 , n35431 , n30632 );
nand ( n261875 , n261868 , n261873 , n261874 );
buf ( n261876 , n261875 );
not ( n261877 , n230043 );
not ( n261878 , n248056 );
or ( n261879 , n261877 , n261878 );
not ( n261880 , n230043 );
nand ( n261881 , n261880 , n256547 );
nand ( n261882 , n261879 , n261881 );
and ( n261883 , n261882 , n248062 );
not ( n261884 , n261882 );
and ( n261885 , n261884 , n248067 );
nor ( n261886 , n261883 , n261885 );
nor ( n261887 , n261886 , n54208 );
not ( n261888 , n226524 );
not ( n261889 , n239220 );
or ( n261890 , n261888 , n261889 );
not ( n261891 , n226524 );
nand ( n261892 , n261891 , n239228 );
nand ( n261893 , n261890 , n261892 );
and ( n261894 , n261893 , n250577 );
not ( n261895 , n261893 );
and ( n261896 , n261895 , n250580 );
nor ( n261897 , n261894 , n261896 );
nand ( n261898 , n261887 , n261897 , n247762 );
not ( n261899 , n261886 );
not ( n261900 , n261899 );
not ( n261901 , n261897 );
or ( n261902 , n261900 , n261901 );
nor ( n261903 , n247762 , n242391 );
nand ( n261904 , n261902 , n261903 );
nand ( n261905 , n31577 , n25896 );
nand ( n261906 , n261898 , n261904 , n261905 );
buf ( n261907 , n261906 );
not ( n261908 , n257100 );
not ( n261909 , n249229 );
not ( n261910 , n244889 );
or ( n261911 , n261909 , n261910 );
not ( n261912 , n249229 );
nand ( n261913 , n261912 , n244899 );
nand ( n261914 , n261911 , n261913 );
and ( n261915 , n261914 , n244955 );
not ( n261916 , n261914 );
and ( n261917 , n261916 , n244940 );
nor ( n261918 , n261915 , n261917 );
not ( n261919 , n261918 );
not ( n261920 , n261919 );
or ( n261921 , n261908 , n261920 );
not ( n261922 , n254908 );
nor ( n261923 , n261922 , n251190 );
nand ( n261924 , n261921 , n261923 );
nand ( n261925 , n257095 , n261919 , n261922 );
nand ( n261926 , n31577 , n33337 );
nand ( n261927 , n261924 , n261925 , n261926 );
buf ( n261928 , n261927 );
not ( n261929 , n44285 );
not ( n261930 , n234106 );
or ( n261931 , n261929 , n261930 );
or ( n261932 , n234106 , n44285 );
nand ( n261933 , n261931 , n261932 );
and ( n261934 , n261933 , n249463 );
not ( n261935 , n261933 );
and ( n261936 , n261935 , n249470 );
nor ( n261937 , n261934 , n261936 );
not ( n261938 , n242238 );
not ( n261939 , n249298 );
or ( n261940 , n261938 , n261939 );
not ( n261941 , n242238 );
nand ( n261942 , n261941 , n53140 );
nand ( n261943 , n261940 , n261942 );
and ( n261944 , n261943 , n249366 );
not ( n261945 , n261943 );
and ( n261946 , n261945 , n249363 );
nor ( n261947 , n261944 , n261946 );
not ( n261948 , n261947 );
nand ( n261949 , n261937 , n261948 );
nor ( n261950 , n239233 , n49959 );
not ( n261951 , n261950 );
or ( n261952 , n261949 , n261951 );
nand ( n261953 , n238901 , n261949 );
nand ( n261954 , n247585 , n35082 );
nand ( n261955 , n261952 , n261953 , n261954 );
buf ( n261956 , n261955 );
not ( n261957 , RI19abd4d0_2356);
or ( n261958 , n233507 , n261957 );
or ( n261959 , n226822 , n246221 );
nand ( n261960 , n261958 , n261959 );
buf ( n261961 , n261960 );
buf ( n261962 , n249710 );
not ( n261963 , n261962 );
not ( n261964 , n255879 );
or ( n261965 , n261963 , n261964 );
or ( n261966 , n255879 , n261962 );
nand ( n261967 , n261965 , n261966 );
not ( n261968 , n261967 );
not ( n261969 , n260195 );
and ( n261970 , n261968 , n261969 );
and ( n261971 , n261967 , n260195 );
nor ( n261972 , n261970 , n261971 );
not ( n261973 , n261972 );
nand ( n261974 , n261973 , n237385 );
not ( n261975 , n261974 );
not ( n261976 , n240861 );
not ( n261977 , n37714 );
or ( n261978 , n261976 , n261977 );
not ( n261979 , n240861 );
nand ( n261980 , n261979 , n37708 );
nand ( n261981 , n261978 , n261980 );
and ( n261982 , n261981 , n244805 );
not ( n261983 , n261981 );
and ( n261984 , n261983 , n244802 );
nor ( n261985 , n261982 , n261984 );
not ( n261986 , n239775 );
not ( n261987 , n244543 );
not ( n261988 , n239705 );
or ( n261989 , n261987 , n261988 );
nand ( n261990 , n239715 , n244544 );
nand ( n261991 , n261989 , n261990 );
not ( n261992 , n261991 );
or ( n261993 , n261986 , n261992 );
or ( n261994 , n261991 , n258810 );
nand ( n261995 , n261993 , n261994 );
not ( n261996 , n261995 );
nand ( n261997 , n261985 , n261996 );
not ( n261998 , n261997 );
and ( n261999 , n261975 , n261998 );
buf ( n262000 , n35431 );
and ( n262001 , n262000 , n35713 );
nor ( n262002 , n261999 , n262001 );
nand ( n262003 , n261972 , n223839 );
not ( n262004 , n262003 );
not ( n262005 , n261985 );
nand ( n262006 , n262004 , n262005 );
nor ( n262007 , n261985 , n47173 );
nand ( n262008 , n262007 , n261995 );
nand ( n262009 , n262002 , n262006 , n262008 );
buf ( n262010 , n262009 );
not ( n262011 , n241868 );
not ( n262012 , n262011 );
not ( n262013 , n248892 );
or ( n262014 , n262012 , n262013 );
nand ( n262015 , n248901 , n241868 );
nand ( n262016 , n262014 , n262015 );
xnor ( n262017 , n262016 , n248907 );
not ( n262018 , n262017 );
not ( n262019 , n47166 );
or ( n262020 , n262018 , n262019 );
not ( n262021 , n234082 );
not ( n262022 , n38222 );
or ( n262023 , n262021 , n262022 );
not ( n262024 , n234082 );
nand ( n262025 , n262024 , n38232 );
nand ( n262026 , n262023 , n262025 );
and ( n262027 , n262026 , n38634 );
not ( n262028 , n262026 );
and ( n262029 , n262028 , n38627 );
nor ( n262030 , n262027 , n262029 );
nor ( n262031 , n262030 , n257769 );
nand ( n262032 , n262020 , n262031 );
nand ( n262033 , n262017 , n239934 );
not ( n262034 , n262033 );
nand ( n262035 , n262034 , n262030 , n47166 );
nand ( n262036 , n46083 , n28213 );
nand ( n262037 , n262032 , n262035 , n262036 );
buf ( n262038 , n262037 );
buf ( n262039 , RI19a24320_2787);
not ( n262040 , n262039 );
not ( n262041 , n257347 );
or ( n262042 , n262040 , n262041 );
buf ( n262043 , RI19a24578_2786);
nand ( n262044 , n257351 , n262043 );
nand ( n262045 , n262042 , n262044 );
buf ( n262046 , n262045 );
not ( n262047 , n257236 );
nand ( n262048 , n262047 , n256158 );
or ( n262049 , n257226 , n262048 );
not ( n262050 , n262047 );
not ( n262051 , n256124 );
or ( n262052 , n262050 , n262051 );
nor ( n262053 , n256158 , n37724 );
nand ( n262054 , n262052 , n262053 );
nand ( n262055 , n237361 , n29135 );
nand ( n262056 , n262049 , n262054 , n262055 );
buf ( n262057 , n262056 );
not ( n262058 , n249871 );
not ( n262059 , n254855 );
not ( n262060 , n55345 );
or ( n262061 , n262059 , n262060 );
not ( n262062 , n254855 );
nand ( n262063 , n262062 , n33708 );
nand ( n262064 , n262061 , n262063 );
and ( n262065 , n262064 , n233265 );
not ( n262066 , n262064 );
and ( n262067 , n262066 , n55511 );
nor ( n262068 , n262065 , n262067 );
not ( n262069 , n262068 );
not ( n262070 , n252436 );
not ( n262071 , n257952 );
or ( n262072 , n262070 , n262071 );
not ( n262073 , n252436 );
nand ( n262074 , n262073 , n257956 );
nand ( n262075 , n262072 , n262074 );
and ( n262076 , n262075 , n257960 );
not ( n262077 , n262075 );
and ( n262078 , n262077 , n257964 );
nor ( n262079 , n262076 , n262078 );
not ( n262080 , n262079 );
nand ( n262081 , n262069 , n262080 );
or ( n262082 , n262058 , n262081 );
not ( n262083 , n262069 );
not ( n262084 , n249794 );
or ( n262085 , n262083 , n262084 );
nor ( n262086 , n262080 , n252258 );
nand ( n262087 , n262085 , n262086 );
nand ( n262088 , n39766 , n35455 );
nand ( n262089 , n262082 , n262087 , n262088 );
buf ( n262090 , n262089 );
buf ( n262091 , n35692 );
nor ( n262092 , n258547 , n256413 );
not ( n262093 , n262092 );
nand ( n262094 , n258631 , n260345 );
or ( n262095 , n262093 , n262094 );
not ( n262096 , n258631 );
not ( n262097 , n258548 );
or ( n262098 , n262096 , n262097 );
nor ( n262099 , n260345 , n35427 );
nand ( n262100 , n262098 , n262099 );
nand ( n262101 , n244987 , n230239 );
nand ( n262102 , n262095 , n262100 , n262101 );
buf ( n262103 , n262102 );
not ( n262104 , n35174 );
not ( n262105 , n258213 );
or ( n262106 , n262104 , n262105 );
xor ( n262107 , n51639 , n256877 );
xor ( n262108 , n262107 , n256870 );
not ( n262109 , n262108 );
not ( n262110 , n251674 );
not ( n262111 , n46941 );
or ( n262112 , n262110 , n262111 );
not ( n262113 , n251674 );
nand ( n262114 , n262113 , n46950 );
nand ( n262115 , n262112 , n262114 );
and ( n262116 , n262115 , n224925 );
not ( n262117 , n262115 );
and ( n262118 , n262117 , n47157 );
nor ( n262119 , n262116 , n262118 );
nand ( n262120 , n262109 , n262119 );
and ( n262121 , n262120 , n247272 );
not ( n262122 , n262120 );
and ( n262123 , n262122 , n247271 );
nor ( n262124 , n262121 , n262123 );
or ( n262125 , n262124 , n259651 );
nand ( n262126 , n262106 , n262125 );
buf ( n262127 , n262126 );
buf ( n262128 , n28769 );
buf ( n262129 , n25817 );
buf ( n262130 , n27985 );
not ( n262131 , RI19ac6878_2281);
or ( n262132 , n25328 , n262131 );
or ( n262133 , n25336 , n242603 );
nand ( n262134 , n262132 , n262133 );
buf ( n262135 , n262134 );
buf ( n262136 , n38419 );
not ( n262137 , RI19ac8e70_2263);
or ( n262138 , n226819 , n262137 );
not ( n262139 , RI19abfd98_2333);
or ( n262140 , n25335 , n262139 );
nand ( n262141 , n262138 , n262140 );
buf ( n262142 , n262141 );
not ( n262143 , RI19a9f908_2572);
or ( n262144 , n25328 , n262143 );
or ( n262145 , n25335 , n234040 );
nand ( n262146 , n262144 , n262145 );
buf ( n262147 , n262146 );
not ( n262148 , n242656 );
not ( n262149 , n244954 );
or ( n262150 , n262148 , n262149 );
or ( n262151 , n244954 , n242656 );
nand ( n262152 , n262150 , n262151 );
and ( n262153 , n262152 , n254867 );
not ( n262154 , n262152 );
and ( n262155 , n262154 , n254874 );
nor ( n262156 , n262153 , n262155 );
nand ( n262157 , n262156 , n244809 );
not ( n262158 , n253813 );
buf ( n262159 , n253420 );
not ( n262160 , n262159 );
not ( n262161 , n253807 );
or ( n262162 , n262160 , n262161 );
or ( n262163 , n253807 , n262159 );
nand ( n262164 , n262162 , n262163 );
not ( n262165 , n262164 );
or ( n262166 , n262158 , n262165 );
buf ( n262167 , n240312 );
or ( n262168 , n262164 , n262167 );
nand ( n262169 , n262166 , n262168 );
not ( n262170 , n222615 );
not ( n262171 , n262170 );
not ( n262172 , n244459 );
or ( n262173 , n262171 , n262172 );
or ( n262174 , n244459 , n262170 );
nand ( n262175 , n262173 , n262174 );
and ( n262176 , n262175 , n257630 );
not ( n262177 , n262175 );
and ( n262178 , n262177 , n244056 );
nor ( n262179 , n262176 , n262178 );
not ( n262180 , n262179 );
nand ( n262181 , n262169 , n262180 );
or ( n262182 , n262157 , n262181 );
not ( n262183 , n262169 );
not ( n262184 , n262156 );
or ( n262185 , n262183 , n262184 );
nor ( n262186 , n262180 , n37724 );
nand ( n262187 , n262185 , n262186 );
nand ( n262188 , n238638 , n41837 );
nand ( n262189 , n262182 , n262187 , n262188 );
buf ( n262190 , n262189 );
not ( n262191 , n237973 );
not ( n262192 , n248170 );
not ( n262193 , n240001 );
or ( n262194 , n262192 , n262193 );
not ( n262195 , n248170 );
nand ( n262196 , n262195 , n239994 );
nand ( n262197 , n262194 , n262196 );
and ( n262198 , n262197 , n240053 );
not ( n262199 , n262197 );
and ( n262200 , n262199 , n240057 );
nor ( n262201 , n262198 , n262200 );
not ( n262202 , n262201 );
nand ( n262203 , n262191 , n262202 );
not ( n262204 , n238112 );
or ( n262205 , n262203 , n262204 );
nor ( n262206 , n237953 , n249030 );
nand ( n262207 , n262203 , n262206 );
nand ( n262208 , n247744 , n33517 );
nand ( n262209 , n262205 , n262207 , n262208 );
buf ( n262210 , n262209 );
buf ( n262211 , n257934 );
not ( n262212 , n262211 );
not ( n262213 , n250681 );
or ( n262214 , n262212 , n262213 );
or ( n262215 , n250681 , n262211 );
nand ( n262216 , n262214 , n262215 );
buf ( n262217 , n34968 );
and ( n262218 , n262216 , n262217 );
not ( n262219 , n262216 );
buf ( n262220 , n34956 );
and ( n262221 , n262219 , n262220 );
nor ( n262222 , n262218 , n262221 );
nand ( n262223 , n262222 , n254528 );
not ( n262224 , n255391 );
nand ( n262225 , n262224 , n255402 );
or ( n262226 , n262223 , n262225 );
not ( n262227 , n262224 );
not ( n262228 , n262222 );
or ( n262229 , n262227 , n262228 );
nor ( n262230 , n255402 , n259801 );
nand ( n262231 , n262229 , n262230 );
nand ( n262232 , n241976 , n40989 );
nand ( n262233 , n262226 , n262231 , n262232 );
buf ( n262234 , n262233 );
nor ( n262235 , n258384 , n258406 );
not ( n262236 , n260083 );
not ( n262237 , n249689 );
or ( n262238 , n262236 , n262237 );
not ( n262239 , n260083 );
nand ( n262240 , n262239 , n251526 );
nand ( n262241 , n262238 , n262240 );
and ( n262242 , n262241 , n249750 );
not ( n262243 , n262241 );
and ( n262244 , n262243 , n251532 );
nor ( n262245 , n262242 , n262244 );
not ( n262246 , n262245 );
nor ( n262247 , n262246 , n257769 );
nand ( n262248 , n262235 , n262247 );
not ( n262249 , n262245 );
not ( n262250 , n258384 );
not ( n262251 , n262250 );
or ( n262252 , n262249 , n262251 );
nor ( n262253 , n258407 , n244216 );
nand ( n262254 , n262252 , n262253 );
nand ( n262255 , n238114 , n31866 );
nand ( n262256 , n262248 , n262254 , n262255 );
buf ( n262257 , n262256 );
nor ( n262258 , n241458 , n47173 );
not ( n262259 , n262258 );
not ( n262260 , n238884 );
not ( n262261 , n261859 );
or ( n262262 , n262260 , n262261 );
or ( n262263 , n261859 , n238884 );
nand ( n262264 , n262262 , n262263 );
and ( n262265 , n262264 , n247563 );
not ( n262266 , n262264 );
and ( n262267 , n262266 , n247553 );
nor ( n262268 , n262265 , n262267 );
nand ( n262269 , n262268 , n241680 );
or ( n262270 , n262259 , n262269 );
not ( n262271 , n262268 );
not ( n262272 , n241458 );
not ( n262273 , n262272 );
or ( n262274 , n262271 , n262273 );
not ( n262275 , n260279 );
nand ( n262276 , n262274 , n262275 );
nand ( n262277 , n39767 , n40398 );
nand ( n262278 , n262270 , n262276 , n262277 );
buf ( n262279 , n262278 );
not ( n262280 , n232299 );
not ( n262281 , n247803 );
not ( n262282 , n232514 );
or ( n262283 , n262281 , n262282 );
nand ( n262284 , n232520 , n247804 );
nand ( n262285 , n262283 , n262284 );
not ( n262286 , n262285 );
and ( n262287 , n262280 , n262286 );
and ( n262288 , n232299 , n262285 );
nor ( n262289 , n262287 , n262288 );
not ( n262290 , n262289 );
not ( n262291 , n256371 );
or ( n262292 , n262290 , n262291 );
xor ( n262293 , n250645 , n240996 );
xor ( n262294 , n262293 , n245618 );
nor ( n262295 , n262294 , n234440 );
nand ( n262296 , n262292 , n262295 );
not ( n262297 , n262289 );
nor ( n262298 , n262297 , n33254 );
nand ( n262299 , n262298 , n262294 , n256371 );
nand ( n262300 , n245414 , n26069 );
nand ( n262301 , n262296 , n262299 , n262300 );
buf ( n262302 , n262301 );
not ( n262303 , n52761 );
not ( n262304 , n228346 );
not ( n262305 , n31560 );
or ( n262306 , n262304 , n262305 );
not ( n262307 , n228346 );
nand ( n262308 , n262307 , n209312 );
nand ( n262309 , n262306 , n262308 );
and ( n262310 , n262309 , n35813 );
not ( n262311 , n262309 );
and ( n262312 , n262311 , n35805 );
nor ( n262313 , n262310 , n262312 );
not ( n262314 , n262313 );
nand ( n262315 , n262303 , n262314 );
or ( n262316 , n230208 , n262315 );
not ( n262317 , n262303 );
not ( n262318 , n230205 );
or ( n262319 , n262317 , n262318 );
nor ( n262320 , n262314 , n39763 );
nand ( n262321 , n262319 , n262320 );
nand ( n262322 , n35431 , n37602 );
nand ( n262323 , n262316 , n262321 , n262322 );
buf ( n262324 , n262323 );
not ( n262325 , n26431 );
not ( n262326 , n237361 );
or ( n262327 , n262325 , n262326 );
nand ( n262328 , n261985 , n261995 );
not ( n262329 , n53998 );
not ( n262330 , n262329 );
not ( n262331 , n238400 );
or ( n262332 , n262330 , n262331 );
not ( n262333 , n262329 );
nand ( n262334 , n262333 , n238408 );
nand ( n262335 , n262332 , n262334 );
and ( n262336 , n262335 , n251451 );
not ( n262337 , n262335 );
and ( n262338 , n262337 , n251444 );
nor ( n262339 , n262336 , n262338 );
not ( n262340 , n262339 );
and ( n262341 , n262328 , n262340 );
not ( n262342 , n262328 );
and ( n262343 , n262342 , n262339 );
nor ( n262344 , n262341 , n262343 );
or ( n262345 , n262344 , n260760 );
nand ( n262346 , n262327 , n262345 );
buf ( n262347 , n262346 );
buf ( n262348 , n258597 );
not ( n262349 , n262348 );
not ( n262350 , n251345 );
or ( n262351 , n262349 , n262350 );
or ( n262352 , n251345 , n262348 );
nand ( n262353 , n262351 , n262352 );
not ( n262354 , n262353 );
not ( n262355 , n261176 );
and ( n262356 , n262354 , n262355 );
and ( n262357 , n262353 , n253378 );
nor ( n262358 , n262356 , n262357 );
nand ( n262359 , n262358 , n246697 );
buf ( n262360 , n256851 );
not ( n262361 , n262360 );
not ( n262362 , n261185 );
or ( n262363 , n262361 , n262362 );
or ( n262364 , n261185 , n262360 );
nand ( n262365 , n262363 , n262364 );
and ( n262366 , n262365 , n31561 );
not ( n262367 , n262365 );
and ( n262368 , n262367 , n31552 );
nor ( n262369 , n262366 , n262368 );
not ( n262370 , n262369 );
not ( n262371 , n244264 );
not ( n262372 , n28929 );
or ( n262373 , n262371 , n262372 );
not ( n262374 , n244264 );
nand ( n262375 , n262374 , n28936 );
nand ( n262376 , n262373 , n262375 );
and ( n262377 , n262376 , n29965 );
not ( n262378 , n262376 );
not ( n262379 , n29965 );
and ( n262380 , n262378 , n262379 );
nor ( n262381 , n262377 , n262380 );
not ( n262382 , n262381 );
nand ( n262383 , n262370 , n262382 );
or ( n262384 , n262359 , n262383 );
not ( n262385 , n262370 );
not ( n262386 , n262358 );
or ( n262387 , n262385 , n262386 );
nor ( n262388 , n262382 , n233971 );
nand ( n262389 , n262387 , n262388 );
nand ( n262390 , n247423 , n39609 );
nand ( n262391 , n262384 , n262389 , n262390 );
buf ( n262392 , n262391 );
not ( n262393 , RI1754b5a8_37);
or ( n262394 , n249128 , n262393 );
nand ( n262395 , n249131 , n26347 );
nand ( n262396 , n262394 , n262395 );
buf ( n262397 , n262396 );
not ( n262398 , RI19a23858_2792);
or ( n262399 , n226819 , n262398 );
not ( n262400 , RI19a85e68_2753);
or ( n262401 , n25335 , n262400 );
nand ( n262402 , n262399 , n262401 );
buf ( n262403 , n262402 );
not ( n262404 , n28412 );
not ( n262405 , n245943 );
or ( n262406 , n262404 , n262405 );
not ( n262407 , n36123 );
not ( n262408 , n249757 );
or ( n262409 , n262407 , n262408 );
not ( n262410 , n36123 );
nand ( n262411 , n262410 , n249749 );
nand ( n262412 , n262409 , n262411 );
and ( n262413 , n262412 , n254644 );
not ( n262414 , n262412 );
and ( n262415 , n262414 , n254647 );
nor ( n262416 , n262413 , n262415 );
not ( n262417 , n262416 );
not ( n262418 , n252032 );
not ( n262419 , n49617 );
or ( n262420 , n262418 , n262419 );
not ( n262421 , n252032 );
nand ( n262422 , n262421 , n49626 );
nand ( n262423 , n262420 , n262422 );
and ( n262424 , n262423 , n253272 );
not ( n262425 , n262423 );
and ( n262426 , n262425 , n253265 );
nor ( n262427 , n262424 , n262426 );
nand ( n262428 , n262417 , n262427 );
not ( n262429 , n56029 );
not ( n262430 , n238182 );
not ( n262431 , n262430 );
or ( n262432 , n262429 , n262431 );
or ( n262433 , n262430 , n56029 );
nand ( n262434 , n262432 , n262433 );
and ( n262435 , n262434 , n251220 );
not ( n262436 , n262434 );
and ( n262437 , n262436 , n251224 );
nor ( n262438 , n262435 , n262437 );
not ( n262439 , n262438 );
and ( n262440 , n262428 , n262439 );
not ( n262441 , n262428 );
and ( n262442 , n262441 , n262438 );
nor ( n262443 , n262440 , n262442 );
or ( n262444 , n262443 , n246091 );
nand ( n262445 , n262406 , n262444 );
buf ( n262446 , n262445 );
not ( n262447 , n204775 );
not ( n262448 , n233501 );
or ( n262449 , n262447 , n262448 );
nand ( n262450 , n258532 , n258524 );
not ( n262451 , n52972 );
not ( n262452 , n246882 );
or ( n262453 , n262451 , n262452 );
nand ( n262454 , n246891 , n52973 );
nand ( n262455 , n262453 , n262454 );
not ( n262456 , n262455 );
not ( n262457 , n258077 );
and ( n262458 , n262456 , n262457 );
and ( n262459 , n262455 , n258077 );
nor ( n262460 , n262458 , n262459 );
not ( n262461 , n262460 );
and ( n262462 , n262450 , n262461 );
not ( n262463 , n262450 );
and ( n262464 , n262463 , n262460 );
nor ( n262465 , n262462 , n262464 );
or ( n262466 , n262465 , n257851 );
nand ( n262467 , n262449 , n262466 );
buf ( n262468 , n262467 );
not ( n262469 , n36171 );
not ( n262470 , n234453 );
or ( n262471 , n262469 , n262470 );
not ( n262472 , n247359 );
not ( n262473 , n262472 );
not ( n262474 , n240508 );
or ( n262475 , n262473 , n262474 );
not ( n262476 , n262472 );
nand ( n262477 , n262476 , n240503 );
nand ( n262478 , n262475 , n262477 );
and ( n262479 , n262478 , n246173 );
not ( n262480 , n262478 );
and ( n262481 , n262480 , n246168 );
nor ( n262482 , n262479 , n262481 );
not ( n262483 , n262482 );
buf ( n262484 , n234840 );
not ( n262485 , n262484 );
not ( n262486 , n47773 );
or ( n262487 , n262485 , n262486 );
or ( n262488 , n47773 , n262484 );
nand ( n262489 , n262487 , n262488 );
not ( n262490 , n262489 );
not ( n262491 , n234437 );
and ( n262492 , n262490 , n262491 );
not ( n262493 , n234420 );
not ( n262494 , n262493 );
and ( n262495 , n262489 , n262494 );
nor ( n262496 , n262492 , n262495 );
nand ( n262497 , n262483 , n262496 );
and ( n262498 , n262497 , n244820 );
not ( n262499 , n262497 );
not ( n262500 , n244820 );
and ( n262501 , n262499 , n262500 );
nor ( n262502 , n262498 , n262501 );
or ( n262503 , n262502 , n254882 );
nand ( n262504 , n262471 , n262503 );
buf ( n262505 , n262504 );
not ( n262506 , n46294 );
not ( n262507 , n248557 );
or ( n262508 , n262506 , n262507 );
not ( n262509 , n46294 );
nand ( n262510 , n262509 , n248565 );
nand ( n262511 , n262508 , n262510 );
and ( n262512 , n262511 , n248679 );
not ( n262513 , n262511 );
and ( n262514 , n262513 , n248678 );
nor ( n262515 , n262512 , n262514 );
nand ( n262516 , n242595 , n262515 );
not ( n262517 , n253622 );
not ( n262518 , n262517 );
not ( n262519 , n246660 );
or ( n262520 , n262518 , n262519 );
not ( n262521 , n262517 );
nand ( n262522 , n262521 , n246653 );
nand ( n262523 , n262520 , n262522 );
and ( n262524 , n262523 , n259371 );
not ( n262525 , n262523 );
buf ( n262526 , n237135 );
and ( n262527 , n262525 , n262526 );
nor ( n262528 , n262524 , n262527 );
not ( n262529 , n262528 );
nand ( n262530 , n262529 , n241704 );
or ( n262531 , n262516 , n262530 );
not ( n262532 , n262529 );
not ( n262533 , n242595 );
or ( n262534 , n262532 , n262533 );
nor ( n262535 , n262515 , n55146 );
nand ( n262536 , n262534 , n262535 );
nand ( n262537 , n238114 , n25535 );
nand ( n262538 , n262531 , n262536 , n262537 );
buf ( n262539 , n262538 );
or ( n262540 , n25328 , n256679 );
not ( n262541 , RI19a91100_2675);
or ( n262542 , n226822 , n262541 );
nand ( n262543 , n262540 , n262542 );
buf ( n262544 , n262543 );
not ( n262545 , RI19accc50_2233);
or ( n262546 , n25328 , n262545 );
not ( n262547 , RI19ac40a0_2299);
or ( n262548 , n226822 , n262547 );
nand ( n262549 , n262546 , n262548 );
buf ( n262550 , n262549 );
or ( n262551 , n25328 , n255713 );
not ( n262552 , RI19a9d400_2589);
or ( n262553 , n25335 , n262552 );
nand ( n262554 , n262551 , n262553 );
buf ( n262555 , n262554 );
not ( n262556 , RI19a9f188_2576);
or ( n262557 , n25328 , n262556 );
or ( n262558 , n25335 , n257605 );
nand ( n262559 , n262557 , n262558 );
buf ( n262560 , n262559 );
nor ( n262561 , n256479 , n254226 );
not ( n262562 , n39867 );
not ( n262563 , n235807 );
or ( n262564 , n262562 , n262563 );
not ( n262565 , n39867 );
nand ( n262566 , n262565 , n235815 );
nand ( n262567 , n262564 , n262566 );
and ( n262568 , n262567 , n235888 );
not ( n262569 , n262567 );
and ( n262570 , n262569 , n235879 );
nor ( n262571 , n262568 , n262570 );
nor ( n262572 , n256492 , n262571 );
nand ( n262573 , n262561 , n262572 );
not ( n262574 , n262571 );
not ( n262575 , n262574 );
nand ( n262576 , n256511 , n256480 );
nand ( n262577 , n262575 , n262576 , n43969 );
nand ( n262578 , n231444 , n207296 );
nand ( n262579 , n262573 , n262577 , n262578 );
buf ( n262580 , n262579 );
not ( n262581 , RI19ab9498_2386);
or ( n262582 , n25328 , n262581 );
not ( n262583 , RI19aaf790_2457);
or ( n262584 , n25336 , n262583 );
nand ( n262585 , n262582 , n262584 );
buf ( n262586 , n262585 );
not ( n262587 , RI19ab8f70_2388);
or ( n262588 , n226819 , n262587 );
not ( n262589 , RI19aaf268_2460);
or ( n262590 , n25336 , n262589 );
nand ( n262591 , n262588 , n262590 );
buf ( n262592 , n262591 );
not ( n262593 , n237927 );
not ( n262594 , n246767 );
or ( n262595 , n262593 , n262594 );
or ( n262596 , n246767 , n237927 );
nand ( n262597 , n262595 , n262596 );
and ( n262598 , n262597 , n254006 );
not ( n262599 , n262597 );
and ( n262600 , n262599 , n254010 );
nor ( n262601 , n262598 , n262600 );
nand ( n262602 , n262601 , n222532 );
not ( n262603 , n252517 );
not ( n262604 , n262603 );
not ( n262605 , n249362 );
or ( n262606 , n262604 , n262605 );
not ( n262607 , n262603 );
not ( n262608 , n249362 );
nand ( n262609 , n262607 , n262608 );
nand ( n262610 , n262606 , n262609 );
and ( n262611 , n262610 , n261547 );
not ( n262612 , n262610 );
and ( n262613 , n262612 , n261550 );
nor ( n262614 , n262611 , n262613 );
not ( n262615 , n262614 );
not ( n262616 , n48441 );
not ( n262617 , n254973 );
or ( n262618 , n262616 , n262617 );
not ( n262619 , n48441 );
and ( n262620 , n254959 , n234832 );
not ( n262621 , n254959 );
and ( n262622 , n262621 , n234831 );
nor ( n262623 , n262620 , n262622 );
not ( n262624 , n254972 );
and ( n262625 , n262623 , n262624 );
not ( n262626 , n262623 );
and ( n262627 , n262626 , n254972 );
nor ( n262628 , n262625 , n262627 );
not ( n262629 , n262628 );
nand ( n262630 , n262619 , n262629 );
nand ( n262631 , n262618 , n262630 );
not ( n262632 , n48019 );
not ( n262633 , n262632 );
xor ( n262634 , n262631 , n262633 );
nand ( n262635 , n262615 , n262634 );
or ( n262636 , n262602 , n262635 );
not ( n262637 , n262615 );
not ( n262638 , n262601 );
or ( n262639 , n262637 , n262638 );
nor ( n262640 , n262634 , n37725 );
nand ( n262641 , n262639 , n262640 );
nand ( n262642 , n241378 , n28952 );
nand ( n262643 , n262636 , n262641 , n262642 );
buf ( n262644 , n262643 );
not ( n262645 , n209367 );
not ( n262646 , n245701 );
or ( n262647 , n262645 , n262646 );
nand ( n262648 , n257052 , n257062 );
not ( n262649 , n39521 );
not ( n262650 , n34956 );
or ( n262651 , n262649 , n262650 );
not ( n262652 , n39521 );
nand ( n262653 , n262652 , n34968 );
nand ( n262654 , n262651 , n262653 );
and ( n262655 , n262654 , n35410 );
not ( n262656 , n262654 );
and ( n262657 , n262656 , n35418 );
nor ( n262658 , n262655 , n262657 );
not ( n262659 , n262658 );
and ( n262660 , n262648 , n262659 );
not ( n262661 , n262648 );
and ( n262662 , n262661 , n262658 );
nor ( n262663 , n262660 , n262662 );
or ( n262664 , n262663 , n254882 );
nand ( n262665 , n262647 , n262664 );
buf ( n262666 , n262665 );
not ( n262667 , RI19ac4b68_2294);
or ( n262668 , n25328 , n262667 );
not ( n262669 , RI19abc4e0_2365);
or ( n262670 , n25335 , n262669 );
nand ( n262671 , n262668 , n262670 );
buf ( n262672 , n262671 );
or ( n262673 , n25328 , n255022 );
not ( n262674 , RI19a95750_2644);
or ( n262675 , n226822 , n262674 );
nand ( n262676 , n262673 , n262675 );
buf ( n262677 , n262676 );
or ( n262678 , n25328 , n262400 );
not ( n262679 , RI19aca9a0_2251);
or ( n262680 , n226822 , n262679 );
nand ( n262681 , n262678 , n262680 );
buf ( n262682 , n262681 );
buf ( n262683 , n249813 );
xnor ( n262684 , n262683 , n51747 );
and ( n262685 , n262684 , n51753 );
not ( n262686 , n262684 );
and ( n262687 , n262686 , n229518 );
nor ( n262688 , n262685 , n262687 );
not ( n262689 , n262688 );
nand ( n262690 , n262689 , n260879 );
not ( n262691 , n249906 );
not ( n262692 , n262691 );
not ( n262693 , n227707 );
or ( n262694 , n262692 , n262693 );
or ( n262695 , n227707 , n262691 );
nand ( n262696 , n262694 , n262695 );
and ( n262697 , n262696 , n242978 );
not ( n262698 , n262696 );
and ( n262699 , n262698 , n242970 );
nor ( n262700 , n262697 , n262699 );
not ( n262701 , n232818 );
not ( n262702 , n237444 );
or ( n262703 , n262701 , n262702 );
or ( n262704 , n237444 , n232818 );
nand ( n262705 , n262703 , n262704 );
not ( n262706 , n262705 );
not ( n262707 , n262706 );
not ( n262708 , n237590 );
or ( n262709 , n262707 , n262708 );
nand ( n262710 , n256153 , n262705 );
nand ( n262711 , n262709 , n262710 );
not ( n262712 , n262711 );
nand ( n262713 , n262700 , n262712 );
or ( n262714 , n262690 , n262713 );
not ( n262715 , n262712 );
not ( n262716 , n262688 );
not ( n262717 , n262716 );
or ( n262718 , n262715 , n262717 );
not ( n262719 , n205649 );
nor ( n262720 , n262700 , n262719 );
nand ( n262721 , n262718 , n262720 );
nand ( n262722 , n247423 , n40109 );
nand ( n262723 , n262714 , n262721 , n262722 );
buf ( n262724 , n262723 );
not ( n262725 , n29972 );
not ( n262726 , n241068 );
or ( n262727 , n262725 , n262726 );
not ( n262728 , n244029 );
not ( n262729 , n262728 );
not ( n262730 , n54917 );
or ( n262731 , n262729 , n262730 );
not ( n262732 , n262728 );
nand ( n262733 , n262732 , n54926 );
nand ( n262734 , n262731 , n262733 );
xor ( n262735 , n262734 , n55068 );
buf ( n262736 , n239643 );
not ( n262737 , n262736 );
not ( n262738 , n36368 );
not ( n262739 , n262738 );
or ( n262740 , n262737 , n262739 );
or ( n262741 , n262738 , n262736 );
nand ( n262742 , n262740 , n262741 );
and ( n262743 , n262742 , n249482 );
not ( n262744 , n262742 );
and ( n262745 , n262744 , n36730 );
nor ( n262746 , n262743 , n262745 );
nand ( n262747 , n262735 , n262746 );
not ( n262748 , n244910 );
not ( n262749 , n34448 );
or ( n262750 , n262748 , n262749 );
or ( n262751 , n34448 , n244910 );
nand ( n262752 , n262750 , n262751 );
not ( n262753 , n262752 );
not ( n262754 , n33709 );
and ( n262755 , n262753 , n262754 );
and ( n262756 , n262752 , n33709 );
nor ( n262757 , n262755 , n262756 );
not ( n262758 , n262757 );
and ( n262759 , n262747 , n262758 );
not ( n262760 , n262747 );
and ( n262761 , n262760 , n262757 );
nor ( n262762 , n262759 , n262761 );
or ( n262763 , n262762 , n237358 );
nand ( n262764 , n262727 , n262763 );
buf ( n262765 , n262764 );
not ( n262766 , n252537 );
not ( n262767 , n262766 );
not ( n262768 , n261542 );
or ( n262769 , n262767 , n262768 );
or ( n262770 , n249362 , n262766 );
nand ( n262771 , n262769 , n262770 );
and ( n262772 , n262771 , n261547 );
not ( n262773 , n262771 );
and ( n262774 , n262773 , n261550 );
nor ( n262775 , n262772 , n262774 );
nand ( n262776 , n262775 , n259619 );
not ( n262777 , n234200 );
not ( n262778 , n41929 );
or ( n262779 , n262777 , n262778 );
not ( n262780 , n234200 );
nand ( n262781 , n262780 , n41933 );
nand ( n262782 , n262779 , n262781 );
not ( n262783 , n259105 );
and ( n262784 , n262782 , n262783 );
not ( n262785 , n262782 );
not ( n262786 , n262783 );
and ( n262787 , n262785 , n262786 );
nor ( n262788 , n262784 , n262787 );
not ( n262789 , n255814 );
not ( n262790 , n51106 );
not ( n262791 , n257184 );
or ( n262792 , n262790 , n262791 );
not ( n262793 , n51106 );
nand ( n262794 , n262793 , n255762 );
nand ( n262795 , n262792 , n262794 );
not ( n262796 , n262795 );
or ( n262797 , n262789 , n262796 );
or ( n262798 , n255814 , n262795 );
nand ( n262799 , n262797 , n262798 );
not ( n262800 , n262799 );
nand ( n262801 , n262788 , n262800 );
or ( n262802 , n262776 , n262801 );
not ( n262803 , n262800 );
not ( n262804 , n262775 );
or ( n262805 , n262803 , n262804 );
nor ( n262806 , n262788 , n242391 );
nand ( n262807 , n262805 , n262806 );
nand ( n262808 , n261585 , n25784 );
nand ( n262809 , n262802 , n262807 , n262808 );
buf ( n262810 , n262809 );
not ( n262811 , n27839 );
not ( n262812 , n37728 );
or ( n262813 , n262811 , n262812 );
not ( n262814 , n250576 );
not ( n262815 , n253787 );
and ( n262816 , n262814 , n262815 );
and ( n262817 , n250576 , n253787 );
nor ( n262818 , n262816 , n262817 );
and ( n262819 , n262818 , n252037 );
not ( n262820 , n262818 );
and ( n262821 , n262820 , n252052 );
nor ( n262822 , n262819 , n262821 );
not ( n262823 , n257927 );
not ( n262824 , n250681 );
or ( n262825 , n262823 , n262824 );
not ( n262826 , n257927 );
nand ( n262827 , n262826 , n250691 );
nand ( n262828 , n262825 , n262827 );
and ( n262829 , n262828 , n262220 );
not ( n262830 , n262828 );
and ( n262831 , n262830 , n262217 );
nor ( n262832 , n262829 , n262831 );
nand ( n262833 , n262822 , n262832 );
not ( n262834 , n241947 );
not ( n262835 , n262834 );
not ( n262836 , n256152 );
or ( n262837 , n262835 , n262836 );
not ( n262838 , n262834 );
nand ( n262839 , n262838 , n237590 );
nand ( n262840 , n262837 , n262839 );
and ( n262841 , n262840 , n259578 );
not ( n262842 , n262840 );
and ( n262843 , n262842 , n259575 );
nor ( n262844 , n262841 , n262843 );
not ( n262845 , n262844 );
and ( n262846 , n262833 , n262845 );
not ( n262847 , n262833 );
and ( n262848 , n262847 , n262844 );
nor ( n262849 , n262846 , n262848 );
or ( n262850 , n262849 , n251462 );
nand ( n262851 , n262813 , n262850 );
buf ( n262852 , n262851 );
nand ( n262853 , n254103 , n254095 );
not ( n262854 , n249564 );
not ( n262855 , n257541 );
or ( n262856 , n262854 , n262855 );
not ( n262857 , n249564 );
nand ( n262858 , n262857 , n243006 );
nand ( n262859 , n262856 , n262858 );
and ( n262860 , n262859 , n243199 );
not ( n262861 , n262859 );
and ( n262862 , n262861 , n243198 );
nor ( n262863 , n262860 , n262862 );
nand ( n262864 , n262863 , n237385 );
or ( n262865 , n262853 , n262864 );
nor ( n262866 , n262863 , n50944 );
nand ( n262867 , n262866 , n262853 );
nand ( n262868 , n238114 , n32415 );
nand ( n262869 , n262865 , n262867 , n262868 );
buf ( n262870 , n262869 );
not ( n262871 , n234731 );
not ( n262872 , n242675 );
or ( n262873 , n262871 , n262872 );
or ( n262874 , n242675 , n234731 );
nand ( n262875 , n262873 , n262874 );
and ( n262876 , n262875 , n242683 );
not ( n262877 , n262875 );
and ( n262878 , n262877 , n242680 );
nor ( n262879 , n262876 , n262878 );
nand ( n262880 , n262879 , n241704 );
not ( n262881 , n233091 );
not ( n262882 , n41423 );
not ( n262883 , n233026 );
or ( n262884 , n262882 , n262883 );
or ( n262885 , n233026 , n41423 );
nand ( n262886 , n262884 , n262885 );
not ( n262887 , n262886 );
or ( n262888 , n262881 , n262887 );
or ( n262889 , n262886 , n233091 );
nand ( n262890 , n262888 , n262889 );
not ( n262891 , n42318 );
not ( n262892 , n234305 );
or ( n262893 , n262891 , n262892 );
not ( n262894 , n42318 );
nand ( n262895 , n262894 , n234298 );
nand ( n262896 , n262893 , n262895 );
and ( n262897 , n262896 , n257164 );
not ( n262898 , n262896 );
and ( n262899 , n262898 , n256928 );
nor ( n262900 , n262897 , n262899 );
nor ( n262901 , n262890 , n262900 );
or ( n262902 , n262880 , n262901 );
nor ( n262903 , n262879 , n250909 );
nand ( n262904 , n262903 , n262901 );
nand ( n262905 , n247585 , n31719 );
nand ( n262906 , n262902 , n262904 , n262905 );
buf ( n262907 , n262906 );
not ( n262908 , n236046 );
not ( n262909 , n260550 );
or ( n262910 , n262908 , n262909 );
not ( n262911 , n236046 );
nand ( n262912 , n262911 , n260557 );
nand ( n262913 , n262910 , n262912 );
buf ( n262914 , n256950 );
not ( n262915 , n262914 );
and ( n262916 , n262913 , n262915 );
not ( n262917 , n262913 );
and ( n262918 , n262917 , n262914 );
nor ( n262919 , n262916 , n262918 );
nor ( n262920 , n262919 , n43968 );
not ( n262921 , n237763 );
not ( n262922 , n245392 );
or ( n262923 , n262921 , n262922 );
not ( n262924 , n237763 );
nand ( n262925 , n262924 , n245402 );
nand ( n262926 , n262923 , n262925 );
not ( n262927 , n262926 );
not ( n262928 , n259527 );
and ( n262929 , n262927 , n262928 );
and ( n262930 , n262926 , n259531 );
nor ( n262931 , n262929 , n262930 );
nand ( n262932 , n262920 , n262931 , n261565 );
not ( n262933 , n262919 );
not ( n262934 , n262933 );
not ( n262935 , n262931 );
or ( n262936 , n262934 , n262935 );
nor ( n262937 , n261565 , n256481 );
nand ( n262938 , n262936 , n262937 );
nand ( n262939 , n237361 , n35238 );
nand ( n262940 , n262932 , n262938 , n262939 );
buf ( n262941 , n262940 );
not ( n262942 , n26236 );
not ( n262943 , n245943 );
or ( n262944 , n262942 , n262943 );
not ( n262945 , n245100 );
not ( n262946 , n231768 );
or ( n262947 , n262945 , n262946 );
not ( n262948 , n245100 );
nand ( n262949 , n262948 , n231775 );
nand ( n262950 , n262947 , n262949 );
buf ( n262951 , n40918 );
and ( n262952 , n262950 , n262951 );
not ( n262953 , n262950 );
and ( n262954 , n262953 , n261292 );
nor ( n262955 , n262952 , n262954 );
nand ( n262956 , n254635 , n262955 );
and ( n262957 , n262956 , n254649 );
not ( n262958 , n262956 );
and ( n262959 , n262958 , n254650 );
nor ( n262960 , n262957 , n262959 );
not ( n262961 , n258327 );
not ( n262962 , n262961 );
or ( n262963 , n262960 , n262962 );
nand ( n262964 , n262944 , n262963 );
buf ( n262965 , n262964 );
or ( n262966 , n25328 , n241384 );
not ( n262967 , RI19ac3920_2302);
or ( n262968 , n25336 , n262967 );
nand ( n262969 , n262966 , n262968 );
buf ( n262970 , n262969 );
not ( n262971 , n30993 );
not ( n262972 , n237361 );
or ( n262973 , n262971 , n262972 );
nand ( n262974 , n243246 , n243267 );
not ( n262975 , n236182 );
not ( n262976 , n241255 );
or ( n262977 , n262975 , n262976 );
or ( n262978 , n241255 , n236182 );
nand ( n262979 , n262977 , n262978 );
and ( n262980 , n262979 , n241370 );
not ( n262981 , n262979 );
and ( n262982 , n262981 , n241361 );
nor ( n262983 , n262980 , n262982 );
and ( n262984 , n262974 , n262983 );
not ( n262985 , n262974 );
not ( n262986 , n262983 );
and ( n262987 , n262985 , n262986 );
nor ( n262988 , n262984 , n262987 );
or ( n262989 , n262988 , n255967 );
nand ( n262990 , n262973 , n262989 );
buf ( n262991 , n262990 );
not ( n262992 , n244663 );
not ( n262993 , n241723 );
or ( n262994 , n262992 , n262993 );
or ( n262995 , n231211 , n244663 );
nand ( n262996 , n262994 , n262995 );
and ( n262997 , n262996 , n241878 );
not ( n262998 , n262996 );
and ( n262999 , n262998 , n241885 );
nor ( n263000 , n262997 , n262999 );
nand ( n263001 , n263000 , n241459 );
not ( n263002 , n250084 );
not ( n263003 , n236063 );
or ( n263004 , n263002 , n263003 );
not ( n263005 , n236056 );
or ( n263006 , n263005 , n250084 );
nand ( n263007 , n263004 , n263006 );
and ( n263008 , n263007 , n236172 );
not ( n263009 , n263007 );
and ( n263010 , n263009 , n236171 );
nor ( n263011 , n263008 , n263010 );
not ( n263012 , n253243 );
not ( n263013 , n240684 );
or ( n263014 , n263012 , n263013 );
not ( n263015 , n253243 );
nand ( n263016 , n263015 , n240676 );
nand ( n263017 , n263014 , n263016 );
and ( n263018 , n263017 , n240801 );
not ( n263019 , n263017 );
and ( n263020 , n263019 , n240811 );
nor ( n263021 , n263018 , n263020 );
nand ( n263022 , n263011 , n263021 );
or ( n263023 , n263001 , n263022 );
not ( n263024 , n263021 );
not ( n263025 , n263000 );
or ( n263026 , n263024 , n263025 );
nor ( n263027 , n263011 , n55104 );
nand ( n263028 , n263026 , n263027 );
nand ( n263029 , n239240 , n33929 );
nand ( n263030 , n263023 , n263028 , n263029 );
buf ( n263031 , n263030 );
not ( n263032 , n246745 );
not ( n263033 , n45261 );
or ( n263034 , n263032 , n263033 );
not ( n263035 , n246745 );
nand ( n263036 , n263035 , n45253 );
nand ( n263037 , n263034 , n263036 );
and ( n263038 , n263037 , n255245 );
not ( n263039 , n263037 );
and ( n263040 , n263039 , n255248 );
nor ( n263041 , n263038 , n263040 );
not ( n263042 , n263041 );
nor ( n263043 , n263042 , n226003 );
not ( n263044 , n263043 );
not ( n263045 , n236994 );
not ( n263046 , n35654 );
not ( n263047 , n236881 );
or ( n263048 , n263046 , n263047 );
or ( n263049 , n236881 , n35654 );
nand ( n263050 , n263048 , n263049 );
not ( n263051 , n263050 );
or ( n263052 , n263045 , n263051 );
not ( n263053 , n263050 );
nand ( n263054 , n263053 , n236993 );
nand ( n263055 , n263052 , n263054 );
not ( n263056 , n249584 );
not ( n263057 , n243006 );
not ( n263058 , n263057 );
or ( n263059 , n263056 , n263058 );
not ( n263060 , n249584 );
nand ( n263061 , n263060 , n243006 );
nand ( n263062 , n263059 , n263061 );
and ( n263063 , n263062 , n243198 );
not ( n263064 , n263062 );
and ( n263065 , n263064 , n243199 );
nor ( n263066 , n263063 , n263065 );
not ( n263067 , n263066 );
nor ( n263068 , n263055 , n263067 );
or ( n263069 , n263044 , n263068 );
nor ( n263070 , n263041 , n40465 );
nand ( n263071 , n263070 , n263068 );
nand ( n263072 , n31577 , n31962 );
nand ( n263073 , n263069 , n263071 , n263072 );
buf ( n263074 , n263073 );
buf ( n263075 , n35713 );
not ( n263076 , n31370 );
not ( n263077 , n245943 );
or ( n263078 , n263076 , n263077 );
not ( n263079 , n257729 );
not ( n263080 , n37661 );
not ( n263081 , n252444 );
or ( n263082 , n263080 , n263081 );
not ( n263083 , n37661 );
nand ( n263084 , n263083 , n257724 );
nand ( n263085 , n263082 , n263084 );
not ( n263086 , n263085 );
or ( n263087 , n263079 , n263086 );
or ( n263088 , n263085 , n257729 );
nand ( n263089 , n263087 , n263088 );
nand ( n263090 , n259901 , n263089 );
not ( n263091 , n259891 );
and ( n263092 , n263090 , n263091 );
not ( n263093 , n263090 );
and ( n263094 , n263093 , n259891 );
nor ( n263095 , n263092 , n263094 );
or ( n263096 , n263095 , n260760 );
nand ( n263097 , n263078 , n263096 );
buf ( n263098 , n263097 );
and ( n263099 , n51187 , n256762 );
not ( n263100 , n51187 );
and ( n263101 , n263100 , n256761 );
or ( n263102 , n263099 , n263101 );
and ( n263103 , n263102 , n256765 );
not ( n263104 , n263102 );
and ( n263105 , n263104 , n253673 );
nor ( n263106 , n263103 , n263105 );
nor ( n263107 , n263106 , n256481 );
not ( n263108 , n263107 );
buf ( n263109 , n243619 );
not ( n263110 , n263109 );
not ( n263111 , n255100 );
or ( n263112 , n263110 , n263111 );
or ( n263113 , n258514 , n263109 );
nand ( n263114 , n263112 , n263113 );
not ( n263115 , n263114 );
not ( n263116 , n258512 );
and ( n263117 , n263115 , n263116 );
and ( n263118 , n263114 , n259218 );
nor ( n263119 , n263117 , n263118 );
not ( n263120 , n247109 );
not ( n263121 , n253578 );
or ( n263122 , n263120 , n263121 );
not ( n263123 , n247109 );
not ( n263124 , n253464 );
nand ( n263125 , n263123 , n263124 );
nand ( n263126 , n263122 , n263125 );
and ( n263127 , n263126 , n253478 );
not ( n263128 , n263126 );
and ( n263129 , n263128 , n253475 );
nor ( n263130 , n263127 , n263129 );
not ( n263131 , n263130 );
nand ( n263132 , n263119 , n263131 );
or ( n263133 , n263108 , n263132 );
not ( n263134 , n263131 );
not ( n263135 , n263106 );
not ( n263136 , n263135 );
or ( n263137 , n263134 , n263136 );
nor ( n263138 , n263119 , n234110 );
nand ( n263139 , n263137 , n263138 );
nand ( n263140 , n35431 , n32811 );
nand ( n263141 , n263133 , n263139 , n263140 );
buf ( n263142 , n263141 );
buf ( n263143 , n28552 );
not ( n263144 , n250913 );
not ( n263145 , n250858 );
not ( n263146 , n263145 );
or ( n263147 , n263144 , n263146 );
not ( n263148 , n245586 );
not ( n263149 , n232899 );
or ( n263150 , n263148 , n263149 );
not ( n263151 , n245586 );
nand ( n263152 , n263151 , n37289 );
nand ( n263153 , n263150 , n263152 );
and ( n263154 , n263153 , n37709 );
not ( n263155 , n263153 );
and ( n263156 , n263155 , n37715 );
nor ( n263157 , n263154 , n263156 );
not ( n263158 , n263157 );
nor ( n263159 , n263158 , n254740 );
nand ( n263160 , n263147 , n263159 );
nor ( n263161 , n250858 , n263157 );
nand ( n263162 , n250910 , n263161 );
nand ( n263163 , n256673 , n208179 );
nand ( n263164 , n263160 , n263162 , n263163 );
buf ( n263165 , n263164 );
buf ( n263166 , n240098 );
not ( n263167 , n263166 );
not ( n263168 , n255992 );
or ( n263169 , n263167 , n263168 );
or ( n263170 , n256695 , n263166 );
nand ( n263171 , n263169 , n263170 );
not ( n263172 , n263171 );
not ( n263173 , n247119 );
or ( n263174 , n263172 , n263173 );
or ( n263175 , n255998 , n263171 );
nand ( n263176 , n263174 , n263175 );
not ( n263177 , n263176 );
nand ( n263178 , n260856 , n263177 );
or ( n263179 , n238633 , n263178 );
not ( n263180 , n238632 );
not ( n263181 , n260856 );
or ( n263182 , n263180 , n263181 );
and ( n263183 , n263176 , n250111 );
nand ( n263184 , n263182 , n263183 );
nand ( n263185 , n246460 , n35195 );
nand ( n263186 , n263179 , n263184 , n263185 );
buf ( n263187 , n263186 );
not ( n263188 , RI19abd2f0_2357);
or ( n263189 , n25328 , n263188 );
not ( n263190 , RI19ab34f8_2429);
or ( n263191 , n25336 , n263190 );
nand ( n263192 , n263189 , n263191 );
buf ( n263193 , n263192 );
not ( n263194 , RI19ab6cc0_2403);
or ( n263195 , n233507 , n263194 );
not ( n263196 , RI19a83690_2770);
or ( n263197 , n226822 , n263196 );
nand ( n263198 , n263195 , n263197 );
buf ( n263199 , n263198 );
not ( n263200 , n29346 );
not ( n263201 , n263200 );
not ( n263202 , n256711 );
or ( n263203 , n263201 , n263202 );
not ( n263204 , n263200 );
nand ( n263205 , n263204 , n253009 );
nand ( n263206 , n263203 , n263205 );
buf ( n263207 , n248143 );
and ( n263208 , n263206 , n263207 );
not ( n263209 , n263206 );
and ( n263210 , n263209 , n253015 );
nor ( n263211 , n263208 , n263210 );
nand ( n263212 , n263211 , n222531 );
not ( n263213 , n233601 );
not ( n263214 , n49181 );
or ( n263215 , n263213 , n263214 );
not ( n263216 , n233601 );
nand ( n263217 , n263216 , n49190 );
nand ( n263218 , n263215 , n263217 );
and ( n263219 , n263218 , n238183 );
not ( n263220 , n263218 );
and ( n263221 , n263220 , n238186 );
nor ( n263222 , n263219 , n263221 );
not ( n263223 , n240768 );
not ( n263224 , n247348 );
or ( n263225 , n263223 , n263224 );
not ( n263226 , n240768 );
and ( n263227 , n247327 , n247343 );
not ( n263228 , n247327 );
and ( n263229 , n263228 , n247344 );
nor ( n263230 , n263227 , n263229 );
nand ( n263231 , n263226 , n263230 );
nand ( n263232 , n263225 , n263231 );
and ( n263233 , n263232 , n257952 );
not ( n263234 , n263232 );
not ( n263235 , n257952 );
and ( n263236 , n263234 , n263235 );
nor ( n263237 , n263233 , n263236 );
not ( n263238 , n263237 );
nand ( n263239 , n263222 , n263238 );
or ( n263240 , n263212 , n263239 );
not ( n263241 , n263238 );
not ( n263242 , n263211 );
or ( n263243 , n263241 , n263242 );
nor ( n263244 , n263222 , n244399 );
nand ( n263245 , n263243 , n263244 );
nand ( n263246 , n35431 , n31248 );
nand ( n263247 , n263240 , n263245 , n263246 );
buf ( n263248 , n263247 );
nor ( n263249 , n254793 , n39763 );
not ( n263250 , n263249 );
not ( n263251 , n257155 );
nand ( n263252 , n263251 , n257168 );
or ( n263253 , n263250 , n263252 );
nand ( n263254 , n254758 , n263252 );
nand ( n263255 , n234453 , n31991 );
nand ( n263256 , n263253 , n263254 , n263255 );
buf ( n263257 , n263256 );
not ( n263258 , RI19ac6e18_2278);
or ( n263259 , n25328 , n263258 );
not ( n263260 , RI19abdf98_2350);
or ( n263261 , n25335 , n263260 );
nand ( n263262 , n263259 , n263261 );
buf ( n263263 , n263262 );
buf ( n263264 , RI17539218_590);
and ( n263265 , n27883 , n263264 );
buf ( n263266 , n263265 );
nand ( n263267 , n231459 , n54018 );
not ( n263268 , n49703 );
not ( n263269 , n263268 );
not ( n263270 , n259738 );
or ( n263271 , n263269 , n263270 );
or ( n263272 , n246693 , n263268 );
nand ( n263273 , n263271 , n263272 );
and ( n263274 , n263273 , n259744 );
not ( n263275 , n263273 );
and ( n263276 , n263275 , n259747 );
nor ( n263277 , n263274 , n263276 );
not ( n263278 , n263277 );
nand ( n263279 , n263278 , n249288 );
or ( n263280 , n263267 , n263279 );
not ( n263281 , n263278 );
not ( n263282 , n231459 );
or ( n263283 , n263281 , n263282 );
nor ( n263284 , n54018 , n39763 );
nand ( n263285 , n263283 , n263284 );
buf ( n263286 , RI173f7b58_1548);
nand ( n263287 , n31577 , n263286 );
nand ( n263288 , n263280 , n263285 , n263287 );
buf ( n263289 , n263288 );
buf ( n263290 , n226233 );
not ( n263291 , n263290 );
not ( n263292 , n262629 );
or ( n263293 , n263291 , n263292 );
not ( n263294 , n254973 );
or ( n263295 , n263294 , n263290 );
nand ( n263296 , n263293 , n263295 );
buf ( n263297 , n48015 );
and ( n263298 , n263296 , n263297 );
not ( n263299 , n263296 );
and ( n263300 , n263299 , n262633 );
nor ( n263301 , n263298 , n263300 );
nand ( n263302 , n263301 , n241459 );
not ( n263303 , n252402 );
not ( n263304 , n257952 );
or ( n263305 , n263303 , n263304 );
not ( n263306 , n252402 );
nand ( n263307 , n263306 , n257956 );
nand ( n263308 , n263305 , n263307 );
and ( n263309 , n263308 , n257960 );
not ( n263310 , n263308 );
and ( n263311 , n263310 , n257964 );
nor ( n263312 , n263309 , n263311 );
not ( n263313 , n263312 );
not ( n263314 , n248668 );
not ( n263315 , n251845 );
or ( n263316 , n263314 , n263315 );
not ( n263317 , n248668 );
nand ( n263318 , n263317 , n251855 );
nand ( n263319 , n263316 , n263318 );
and ( n263320 , n263319 , n260967 );
not ( n263321 , n263319 );
and ( n263322 , n263321 , n260966 );
nor ( n263323 , n263320 , n263322 );
nand ( n263324 , n263313 , n263323 );
or ( n263325 , n263302 , n263324 );
not ( n263326 , n263313 );
not ( n263327 , n263301 );
or ( n263328 , n263326 , n263327 );
nor ( n263329 , n263323 , n247212 );
nand ( n263330 , n263328 , n263329 );
nand ( n263331 , n246460 , n34971 );
nand ( n263332 , n263325 , n263330 , n263331 );
buf ( n263333 , n263332 );
and ( n263334 , n250998 , n260640 );
not ( n263335 , n250998 );
not ( n263336 , n260640 );
and ( n263337 , n263335 , n263336 );
or ( n263338 , n263334 , n263337 );
not ( n263339 , n245174 );
and ( n263340 , n263338 , n263339 );
not ( n263341 , n263338 );
and ( n263342 , n263341 , n260647 );
nor ( n263343 , n263340 , n263342 );
not ( n263344 , n255073 );
not ( n263345 , n34947 );
not ( n263346 , n255080 );
or ( n263347 , n263345 , n263346 );
or ( n263348 , n255080 , n34947 );
nand ( n263349 , n263347 , n263348 );
not ( n263350 , n263349 );
and ( n263351 , n263344 , n263350 );
not ( n263352 , n255088 );
and ( n263353 , n263352 , n263349 );
nor ( n263354 , n263351 , n263353 );
nor ( n263355 , n263354 , n236795 );
not ( n263356 , n241839 );
not ( n263357 , n248892 );
or ( n263358 , n263356 , n263357 );
not ( n263359 , n241839 );
nand ( n263360 , n263359 , n248901 );
nand ( n263361 , n263358 , n263360 );
and ( n263362 , n263361 , n248904 );
not ( n263363 , n263361 );
and ( n263364 , n263363 , n248907 );
nor ( n263365 , n263362 , n263364 );
nand ( n263366 , n263355 , n263365 );
or ( n263367 , n263343 , n263366 );
not ( n263368 , n263343 );
not ( n263369 , n263354 );
nand ( n263370 , n263365 , n263369 );
nand ( n263371 , n263370 , n255152 );
or ( n263372 , n263368 , n263371 );
nand ( n263373 , n31577 , n25578 );
nand ( n263374 , n263367 , n263372 , n263373 );
buf ( n263375 , n263374 );
not ( n263376 , n235835 );
not ( n263377 , n245797 );
or ( n263378 , n263376 , n263377 );
not ( n263379 , n245791 );
or ( n263380 , n263379 , n235835 );
nand ( n263381 , n263378 , n263380 );
buf ( n263382 , n250805 );
and ( n263383 , n263381 , n263382 );
not ( n263384 , n263381 );
and ( n263385 , n263384 , n250813 );
nor ( n263386 , n263383 , n263385 );
nor ( n263387 , n263386 , n252358 );
nor ( n263388 , n235024 , n234893 );
nand ( n263389 , n263387 , n263388 );
not ( n263390 , n263386 );
nor ( n263391 , n263390 , n251361 );
nand ( n263392 , n263391 , n234893 );
nand ( n263393 , n234893 , n256957 );
not ( n263394 , n263393 );
nand ( n263395 , n263394 , n235024 );
nand ( n263396 , n39766 , n28658 );
nand ( n263397 , n263389 , n263392 , n263395 , n263396 );
buf ( n263398 , n263397 );
nand ( n263399 , n254769 , n256751 );
nand ( n263400 , n257155 , n254789 );
or ( n263401 , n263399 , n263400 );
not ( n263402 , n254789 );
not ( n263403 , n254769 );
or ( n263404 , n263402 , n263403 );
nor ( n263405 , n257155 , n53680 );
nand ( n263406 , n263404 , n263405 );
nand ( n263407 , n244840 , n41338 );
nand ( n263408 , n263401 , n263406 , n263407 );
buf ( n263409 , n263408 );
not ( n263410 , n37547 );
not ( n263411 , n258715 );
or ( n263412 , n263410 , n263411 );
or ( n263413 , n258715 , n37547 );
nand ( n263414 , n263412 , n263413 );
and ( n263415 , n263414 , n257729 );
not ( n263416 , n263414 );
and ( n263417 , n263416 , n258720 );
nor ( n263418 , n263415 , n263417 );
not ( n263419 , n263418 );
nand ( n263420 , n263419 , n233973 );
not ( n263421 , n238336 );
not ( n263422 , n254337 );
or ( n263423 , n263421 , n263422 );
not ( n263424 , n238336 );
nand ( n263425 , n263424 , n254344 );
nand ( n263426 , n263423 , n263425 );
and ( n263427 , n263426 , n256646 );
not ( n263428 , n263426 );
and ( n263429 , n263428 , n256649 );
nor ( n263430 , n263427 , n263429 );
not ( n263431 , n263430 );
not ( n263432 , n222011 );
not ( n263433 , n234097 );
or ( n263434 , n263432 , n263433 );
not ( n263435 , n222011 );
nand ( n263436 , n263435 , n234106 );
nand ( n263437 , n263434 , n263436 );
and ( n263438 , n263437 , n249470 );
not ( n263439 , n263437 );
and ( n263440 , n263439 , n249463 );
nor ( n263441 , n263438 , n263440 );
not ( n263442 , n263441 );
nand ( n263443 , n263431 , n263442 );
or ( n263444 , n263420 , n263443 );
not ( n263445 , n263419 );
not ( n263446 , n263431 );
or ( n263447 , n263445 , n263446 );
nor ( n263448 , n263442 , n52445 );
nand ( n263449 , n263447 , n263448 );
nand ( n263450 , n238638 , n42576 );
nand ( n263451 , n263444 , n263449 , n263450 );
buf ( n263452 , n263451 );
not ( n263453 , n249613 );
not ( n263454 , n263453 );
not ( n263455 , n257118 );
or ( n263456 , n263454 , n263455 );
nor ( n263457 , n257130 , n240080 );
nand ( n263458 , n263456 , n263457 );
nand ( n263459 , n249620 , n257118 , n257130 );
nand ( n263460 , n252711 , n30974 );
nand ( n263461 , n263458 , n263459 , n263460 );
buf ( n263462 , n263461 );
not ( n263463 , RI19ac30b0_2306);
or ( n263464 , n233507 , n263463 );
not ( n263465 , RI19aba8c0_2377);
or ( n263466 , n25335 , n263465 );
nand ( n263467 , n263464 , n263466 );
buf ( n263468 , n263467 );
not ( n263469 , n258570 );
not ( n263470 , n263469 );
not ( n263471 , n40460 );
or ( n263472 , n263470 , n263471 );
not ( n263473 , n263469 );
nand ( n263474 , n263473 , n251345 );
nand ( n263475 , n263472 , n263474 );
and ( n263476 , n263475 , n253377 );
not ( n263477 , n263475 );
and ( n263478 , n263477 , n253378 );
nor ( n263479 , n263476 , n263478 );
nand ( n263480 , n263479 , n247275 );
not ( n263481 , n243978 );
not ( n263482 , n252317 );
or ( n263483 , n263481 , n263482 );
or ( n263484 , n252317 , n243978 );
nand ( n263485 , n263483 , n263484 );
and ( n263486 , n263485 , n252327 );
not ( n263487 , n263485 );
and ( n263488 , n263487 , n252324 );
nor ( n263489 , n263486 , n263488 );
not ( n263490 , n239673 );
not ( n263491 , n238975 );
or ( n263492 , n263490 , n263491 );
not ( n263493 , n239673 );
nand ( n263494 , n263493 , n238985 );
nand ( n263495 , n263492 , n263494 );
and ( n263496 , n263495 , n239100 );
not ( n263497 , n263495 );
and ( n263498 , n263497 , n239108 );
nor ( n263499 , n263496 , n263498 );
not ( n263500 , n263499 );
nand ( n263501 , n263489 , n263500 );
or ( n263502 , n263480 , n263501 );
not ( n263503 , n263479 );
not ( n263504 , n263489 );
or ( n263505 , n263503 , n263504 );
nor ( n263506 , n263500 , n31572 );
nand ( n263507 , n263505 , n263506 );
nand ( n263508 , n46083 , n42665 );
nand ( n263509 , n263502 , n263507 , n263508 );
buf ( n263510 , n263509 );
not ( n263511 , n52088 );
not ( n263512 , n263511 );
not ( n263513 , n236267 );
or ( n263514 , n263512 , n263513 );
nand ( n263515 , n245210 , n52088 );
nand ( n263516 , n263514 , n263515 );
not ( n263517 , n263516 );
not ( n263518 , n251181 );
and ( n263519 , n263517 , n263518 );
and ( n263520 , n263516 , n251181 );
nor ( n263521 , n263519 , n263520 );
not ( n263522 , n255998 );
not ( n263523 , n240094 );
not ( n263524 , n247644 );
or ( n263525 , n263523 , n263524 );
not ( n263526 , n240094 );
nand ( n263527 , n263526 , n255992 );
nand ( n263528 , n263525 , n263527 );
not ( n263529 , n263528 );
and ( n263530 , n263522 , n263529 );
and ( n263531 , n255998 , n263528 );
nor ( n263532 , n263530 , n263531 );
nand ( n263533 , n263521 , n263532 );
not ( n263534 , n248488 );
or ( n263535 , n263533 , n263534 );
not ( n263536 , n248483 );
not ( n263537 , n263521 );
or ( n263538 , n263536 , n263537 );
nor ( n263539 , n263532 , n31572 );
nand ( n263540 , n263538 , n263539 );
nand ( n263541 , n241378 , n30845 );
nand ( n263542 , n263535 , n263540 , n263541 );
buf ( n263543 , n263542 );
not ( n263544 , RI19aa0790_2565);
or ( n263545 , n25328 , n263544 );
not ( n263546 , RI19a96bf0_2635);
or ( n263547 , n25335 , n263546 );
nand ( n263548 , n263545 , n263547 );
buf ( n263549 , n263548 );
not ( n263550 , n248843 );
not ( n263551 , n237340 );
or ( n263552 , n263550 , n263551 );
not ( n263553 , n248843 );
nand ( n263554 , n263553 , n237350 );
nand ( n263555 , n263552 , n263554 );
xnor ( n263556 , n263555 , n256279 );
not ( n263557 , n263556 );
not ( n263558 , n237559 );
not ( n263559 , n247871 );
or ( n263560 , n263558 , n263559 );
not ( n263561 , n237559 );
not ( n263562 , n247870 );
nand ( n263563 , n263561 , n263562 );
nand ( n263564 , n263560 , n263563 );
not ( n263565 , n263564 );
not ( n263566 , n249285 );
and ( n263567 , n263565 , n263566 );
not ( n263568 , n249274 );
and ( n263569 , n263564 , n263568 );
nor ( n263570 , n263567 , n263569 );
nand ( n263571 , n263557 , n263570 );
nor ( n263572 , n252677 , n235050 );
not ( n263573 , n263572 );
or ( n263574 , n263571 , n263573 );
nand ( n263575 , n263571 , n252680 );
nand ( n263576 , n245414 , n220493 );
nand ( n263577 , n263574 , n263575 , n263576 );
buf ( n263578 , n263577 );
not ( n263579 , n243251 );
not ( n263580 , n41209 );
not ( n263581 , n54263 );
or ( n263582 , n263580 , n263581 );
nand ( n263583 , n54273 , n41205 );
nand ( n263584 , n263582 , n263583 );
and ( n263585 , n263584 , n255321 );
not ( n263586 , n263584 );
and ( n263587 , n263586 , n255324 );
nor ( n263588 , n263585 , n263587 );
not ( n263589 , n263588 );
nand ( n263590 , n262986 , n263589 );
or ( n263591 , n263579 , n263590 );
not ( n263592 , n243246 );
not ( n263593 , n263592 );
not ( n263594 , n262986 );
or ( n263595 , n263593 , n263594 );
nor ( n263596 , n263589 , n49959 );
nand ( n263597 , n263595 , n263596 );
buf ( n263598 , n35431 );
nand ( n263599 , n263598 , n35094 );
nand ( n263600 , n263591 , n263597 , n263599 );
buf ( n263601 , n263600 );
not ( n263602 , n207164 );
not ( n263603 , n234453 );
or ( n263604 , n263602 , n263603 );
not ( n263605 , n46649 );
not ( n263606 , n253196 );
or ( n263607 , n263605 , n263606 );
not ( n263608 , n46649 );
nand ( n263609 , n263608 , n253188 );
nand ( n263610 , n263607 , n263609 );
and ( n263611 , n263610 , n253949 );
not ( n263612 , n263610 );
not ( n263613 , n255303 );
and ( n263614 , n263612 , n263613 );
nor ( n263615 , n263611 , n263614 );
not ( n263616 , n242559 );
not ( n263617 , n227548 );
or ( n263618 , n263616 , n263617 );
not ( n263619 , n242559 );
nand ( n263620 , n263619 , n49786 );
nand ( n263621 , n263618 , n263620 );
and ( n263622 , n263621 , n49947 );
not ( n263623 , n263621 );
and ( n263624 , n263623 , n49950 );
nor ( n263625 , n263622 , n263624 );
nand ( n263626 , n263615 , n263625 );
and ( n263627 , n263626 , n257022 );
not ( n263628 , n263626 );
and ( n263629 , n263628 , n257021 );
nor ( n263630 , n263627 , n263629 );
or ( n263631 , n263630 , n256376 );
nand ( n263632 , n263604 , n263631 );
buf ( n263633 , n263632 );
not ( n263634 , n37952 );
not ( n263635 , n263634 );
not ( n263636 , n50027 );
or ( n263637 , n263635 , n263636 );
not ( n263638 , n263634 );
nand ( n263639 , n263638 , n227795 );
nand ( n263640 , n263637 , n263639 );
and ( n263641 , n263640 , n234522 );
not ( n263642 , n263640 );
and ( n263643 , n263642 , n234514 );
nor ( n263644 , n263641 , n263643 );
not ( n263645 , n263644 );
not ( n263646 , n246872 );
not ( n263647 , n242852 );
or ( n263648 , n263646 , n263647 );
or ( n263649 , n242852 , n246872 );
nand ( n263650 , n263648 , n263649 );
not ( n263651 , n263650 );
not ( n263652 , n208725 );
and ( n263653 , n263651 , n263652 );
and ( n263654 , n263650 , n261185 );
nor ( n263655 , n263653 , n263654 );
nand ( n263656 , n263645 , n260411 , n263655 );
nand ( n263657 , n263655 , n260393 );
nand ( n263658 , n263644 , n263657 , n205649 );
nand ( n263659 , n239240 , n32929 );
nand ( n263660 , n263656 , n263658 , n263659 );
buf ( n263661 , n263660 );
not ( n263662 , n240245 );
not ( n263663 , n252051 );
or ( n263664 , n263662 , n263663 );
not ( n263665 , n240245 );
nand ( n263666 , n263665 , n252036 );
nand ( n263667 , n263664 , n263666 );
and ( n263668 , n263667 , n254223 );
not ( n263669 , n263667 );
and ( n263670 , n263669 , n256227 );
nor ( n263671 , n263668 , n263670 );
nor ( n263672 , n263671 , n221279 );
not ( n263673 , n246619 );
not ( n263674 , n255455 );
or ( n263675 , n263673 , n263674 );
not ( n263676 , n246619 );
nand ( n263677 , n263676 , n255464 );
nand ( n263678 , n263675 , n263677 );
and ( n263679 , n263678 , n259459 );
not ( n263680 , n263678 );
and ( n263681 , n263680 , n259463 );
nor ( n263682 , n263679 , n263681 );
not ( n263683 , n263682 );
nand ( n263684 , n263672 , n263683 );
not ( n263685 , n230851 );
not ( n263686 , n235072 );
not ( n263687 , n263686 );
or ( n263688 , n263685 , n263687 );
not ( n263689 , n230851 );
nand ( n263690 , n263689 , n235072 );
nand ( n263691 , n263688 , n263690 );
and ( n263692 , n263691 , n235203 );
not ( n263693 , n263691 );
and ( n263694 , n263693 , n235211 );
nor ( n263695 , n263692 , n263694 );
nand ( n263696 , n263695 , n250111 );
not ( n263697 , n263696 );
not ( n263698 , n263671 );
and ( n263699 , n263697 , n263698 );
and ( n263700 , n236798 , n207855 );
nor ( n263701 , n263699 , n263700 );
nor ( n263702 , n263695 , n31571 );
nand ( n263703 , n263702 , n263671 , n263682 );
nand ( n263704 , n263684 , n263701 , n263703 );
buf ( n263705 , n263704 );
not ( n263706 , n241401 );
not ( n263707 , n225301 );
or ( n263708 , n263706 , n263707 );
or ( n263709 , n225301 , n241401 );
nand ( n263710 , n263708 , n263709 );
not ( n263711 , n263710 );
not ( n263712 , n256892 );
and ( n263713 , n263711 , n263712 );
and ( n263714 , n263710 , n256892 );
nor ( n263715 , n263713 , n263714 );
nand ( n263716 , n263715 , n245241 );
not ( n263717 , n263089 );
nand ( n263718 , n259914 , n263717 );
or ( n263719 , n263716 , n263718 );
not ( n263720 , n259914 );
not ( n263721 , n263715 );
or ( n263722 , n263720 , n263721 );
nor ( n263723 , n263717 , n233972 );
nand ( n263724 , n263722 , n263723 );
nand ( n263725 , n238638 , n40883 );
nand ( n263726 , n263719 , n263724 , n263725 );
buf ( n263727 , n263726 );
buf ( n263728 , n218281 );
buf ( n263729 , n35259 );
not ( n263730 , n36672 );
not ( n263731 , n253855 );
or ( n263732 , n263730 , n263731 );
not ( n263733 , n36672 );
nand ( n263734 , n263733 , n253863 );
nand ( n263735 , n263732 , n263734 );
and ( n263736 , n263735 , n258013 );
not ( n263737 , n263735 );
and ( n263738 , n263737 , n258012 );
nor ( n263739 , n263736 , n263738 );
nor ( n263740 , n263739 , n52445 );
not ( n263741 , n263740 );
not ( n263742 , n250350 );
not ( n263743 , n237135 );
or ( n263744 , n263742 , n263743 );
not ( n263745 , n250350 );
nand ( n263746 , n263745 , n237148 );
nand ( n263747 , n263744 , n263746 );
and ( n263748 , n263747 , n250412 );
not ( n263749 , n263747 );
and ( n263750 , n263749 , n250408 );
nor ( n263751 , n263748 , n263750 );
not ( n263752 , n263751 );
not ( n263753 , n244131 );
nand ( n263754 , n263752 , n263753 );
or ( n263755 , n263741 , n263754 );
not ( n263756 , n263752 );
not ( n263757 , n263739 );
not ( n263758 , n263757 );
or ( n263759 , n263756 , n263758 );
nor ( n263760 , n263753 , n260567 );
nand ( n263761 , n263759 , n263760 );
nand ( n263762 , n246217 , n204484 );
nand ( n263763 , n263755 , n263761 , n263762 );
buf ( n263764 , n263763 );
not ( n263765 , n243882 );
not ( n263766 , n263765 );
not ( n263767 , n246064 );
or ( n263768 , n263766 , n263767 );
not ( n263769 , n263765 );
nand ( n263770 , n263769 , n246705 );
nand ( n263771 , n263768 , n263770 );
and ( n263772 , n263771 , n246768 );
not ( n263773 , n263771 );
and ( n263774 , n263773 , n246760 );
nor ( n263775 , n263772 , n263774 );
nor ( n263776 , n263775 , n243204 );
not ( n263777 , n253642 );
not ( n263778 , n246660 );
or ( n263779 , n263777 , n263778 );
not ( n263780 , n253642 );
nand ( n263781 , n263780 , n246653 );
nand ( n263782 , n263779 , n263781 );
and ( n263783 , n263782 , n259371 );
not ( n263784 , n263782 );
not ( n263785 , n237135 );
not ( n263786 , n263785 );
and ( n263787 , n263784 , n263786 );
nor ( n263788 , n263783 , n263787 );
not ( n263789 , n244315 );
not ( n263790 , n29962 );
or ( n263791 , n263789 , n263790 );
not ( n263792 , n244315 );
nand ( n263793 , n263792 , n256362 );
nand ( n263794 , n263791 , n263793 );
and ( n263795 , n263794 , n256366 );
not ( n263796 , n263794 );
buf ( n263797 , n235590 );
and ( n263798 , n263796 , n263797 );
nor ( n263799 , n263795 , n263798 );
not ( n263800 , n263799 );
nor ( n263801 , n263788 , n263800 );
nand ( n263802 , n263776 , n263801 );
not ( n263803 , n263775 );
not ( n263804 , n263803 );
not ( n263805 , n263799 );
or ( n263806 , n263804 , n263805 );
not ( n263807 , n263788 );
nor ( n263808 , n263807 , n27889 );
nand ( n263809 , n263806 , n263808 );
nand ( n263810 , n236798 , n205078 );
nand ( n263811 , n263802 , n263809 , n263810 );
buf ( n263812 , n263811 );
or ( n263813 , n25328 , n258653 );
not ( n263814 , RI19a83f78_2766);
or ( n263815 , n25336 , n263814 );
nand ( n263816 , n263813 , n263815 );
buf ( n263817 , n263816 );
not ( n263818 , n29375 );
buf ( n263819 , n35431 );
not ( n263820 , n263819 );
or ( n263821 , n263818 , n263820 );
not ( n263822 , n49856 );
not ( n263823 , n245862 );
or ( n263824 , n263822 , n263823 );
not ( n263825 , n49856 );
nand ( n263826 , n263825 , n245872 );
nand ( n263827 , n263824 , n263826 );
and ( n263828 , n263827 , n245920 );
not ( n263829 , n263827 );
and ( n263830 , n263829 , n245930 );
nor ( n263831 , n263828 , n263830 );
nand ( n263832 , n263831 , n254127 );
and ( n263833 , n263832 , n252329 );
not ( n263834 , n263832 );
not ( n263835 , n252329 );
and ( n263836 , n263834 , n263835 );
nor ( n263837 , n263833 , n263836 );
or ( n263838 , n263837 , n255135 );
nand ( n263839 , n263821 , n263838 );
buf ( n263840 , n263839 );
buf ( n263841 , n33119 );
not ( n263842 , n251056 );
not ( n263843 , n50474 );
or ( n263844 , n263842 , n263843 );
not ( n263845 , n251056 );
nand ( n263846 , n263845 , n50482 );
nand ( n263847 , n263844 , n263846 );
buf ( n263848 , n260640 );
and ( n263849 , n263847 , n263848 );
not ( n263850 , n263847 );
not ( n263851 , n263848 );
and ( n263852 , n263850 , n263851 );
nor ( n263853 , n263849 , n263852 );
not ( n263854 , n244181 );
not ( n263855 , n234810 );
or ( n263856 , n263854 , n263855 );
not ( n263857 , n244181 );
nand ( n263858 , n263857 , n234803 );
nand ( n263859 , n263856 , n263858 );
and ( n263860 , n263859 , n250398 );
not ( n263861 , n263859 );
and ( n263862 , n263861 , n250395 );
nor ( n263863 , n263860 , n263862 );
nand ( n263864 , n263853 , n263863 );
or ( n263865 , n263864 , n239787 );
nand ( n263866 , n263863 , n239780 );
not ( n263867 , n263853 );
nand ( n263868 , n263866 , n263867 , n205649 );
nand ( n263869 , n241976 , n25609 );
nand ( n263870 , n263865 , n263868 , n263869 );
buf ( n263871 , n263870 );
not ( n263872 , RI19aacdd8_2476);
or ( n263873 , n25328 , n263872 );
not ( n263874 , RI19aa2c20_2547);
or ( n263875 , n226822 , n263874 );
nand ( n263876 , n263873 , n263875 );
buf ( n263877 , n263876 );
not ( n263878 , n226585 );
not ( n263879 , n44315 );
or ( n263880 , n263878 , n263879 );
not ( n263881 , n226585 );
nand ( n263882 , n263881 , n44324 );
nand ( n263883 , n263880 , n263882 );
xnor ( n263884 , n263883 , n256460 );
not ( n263885 , n263884 );
nand ( n263886 , n263885 , n245267 );
or ( n263887 , n263886 , n245242 );
nor ( n263888 , n245240 , n247698 );
nand ( n263889 , n263886 , n263888 );
nand ( n263890 , n234024 , n39908 );
nand ( n263891 , n263887 , n263889 , n263890 );
buf ( n263892 , n263891 );
not ( n263893 , n50890 );
not ( n263894 , n251970 );
or ( n263895 , n263893 , n263894 );
not ( n263896 , n50890 );
not ( n263897 , n251970 );
nand ( n263898 , n263896 , n263897 );
nand ( n263899 , n263895 , n263898 );
not ( n263900 , n250896 );
and ( n263901 , n263899 , n263900 );
not ( n263902 , n263899 );
and ( n263903 , n263902 , n250900 );
nor ( n263904 , n263901 , n263903 );
not ( n263905 , n263904 );
not ( n263906 , n257846 );
or ( n263907 , n263905 , n263906 );
nand ( n263908 , n263907 , n260775 );
not ( n263909 , n263904 );
nor ( n263910 , n263909 , n256481 );
nand ( n263911 , n263910 , n260774 , n257846 );
nand ( n263912 , n238114 , n33119 );
nand ( n263913 , n263908 , n263911 , n263912 );
buf ( n263914 , n263913 );
buf ( n263915 , n37394 );
buf ( n263916 , n35577 );
not ( n263917 , n249723 );
not ( n263918 , n255884 );
or ( n263919 , n263917 , n263918 );
not ( n263920 , n249723 );
nand ( n263921 , n263920 , n255879 );
nand ( n263922 , n263919 , n263921 );
and ( n263923 , n263922 , n260195 );
not ( n263924 , n263922 );
and ( n263925 , n263924 , n260198 );
nor ( n263926 , n263923 , n263925 );
not ( n263927 , n234206 );
not ( n263928 , n263927 );
not ( n263929 , n41929 );
or ( n263930 , n263928 , n263929 );
not ( n263931 , n263927 );
nand ( n263932 , n263931 , n41933 );
nand ( n263933 , n263930 , n263932 );
xor ( n263934 , n263933 , n261058 );
not ( n263935 , n263934 );
nand ( n263936 , n263926 , n263935 );
not ( n263937 , n228024 );
not ( n263938 , n248967 );
or ( n263939 , n263937 , n263938 );
not ( n263940 , n228024 );
nand ( n263941 , n263940 , n249394 );
nand ( n263942 , n263939 , n263941 );
and ( n263943 , n263942 , n248975 );
not ( n263944 , n263942 );
and ( n263945 , n263944 , n248972 );
nor ( n263946 , n263943 , n263945 );
not ( n263947 , n263946 );
nor ( n263948 , n263947 , n33254 );
not ( n263949 , n263948 );
or ( n263950 , n263936 , n263949 );
nor ( n263951 , n263946 , n235732 );
nand ( n263952 , n263936 , n263951 );
nand ( n263953 , n241068 , n208497 );
nand ( n263954 , n263950 , n263952 , n263953 );
buf ( n263955 , n263954 );
not ( n263956 , n251404 );
not ( n263957 , n252132 );
or ( n263958 , n263956 , n263957 );
not ( n263959 , n251404 );
nand ( n263960 , n263959 , n252139 );
nand ( n263961 , n263958 , n263960 );
not ( n263962 , n263961 );
not ( n263963 , n252194 );
and ( n263964 , n263962 , n263963 );
not ( n263965 , n252192 );
not ( n263966 , n263965 );
and ( n263967 , n263961 , n263966 );
nor ( n263968 , n263964 , n263967 );
nand ( n263969 , n263968 , n246177 );
nand ( n263970 , n256554 , n257310 );
or ( n263971 , n263969 , n263970 );
nor ( n263972 , n263968 , n247698 );
nand ( n263973 , n263972 , n263970 );
nand ( n263974 , n255116 , n32132 );
nand ( n263975 , n263971 , n263973 , n263974 );
buf ( n263976 , n263975 );
not ( n263977 , n249395 );
not ( n263978 , n250157 );
not ( n263979 , n249388 );
or ( n263980 , n263978 , n263979 );
or ( n263981 , n249388 , n250157 );
nand ( n263982 , n263980 , n263981 );
not ( n263983 , n263982 );
or ( n263984 , n263977 , n263983 );
or ( n263985 , n263982 , n249395 );
nand ( n263986 , n263984 , n263985 );
nor ( n263987 , n245405 , n263986 );
not ( n263988 , n263987 );
not ( n263989 , n263888 );
or ( n263990 , n263988 , n263989 );
not ( n263991 , n35431 );
not ( n263992 , n263991 );
not ( n263993 , n37997 );
and ( n263994 , n263992 , n263993 );
nand ( n263995 , n245239 , n245406 );
not ( n263996 , n263986 );
nor ( n263997 , n263996 , n37725 );
and ( n263998 , n263995 , n263997 );
nor ( n263999 , n263994 , n263998 );
nand ( n264000 , n263990 , n263999 );
buf ( n264001 , n264000 );
not ( n264002 , n238356 );
not ( n264003 , n254337 );
or ( n264004 , n264002 , n264003 );
not ( n264005 , n238356 );
nand ( n264006 , n264005 , n254344 );
nand ( n264007 , n264004 , n264006 );
and ( n264008 , n264007 , n256646 );
not ( n264009 , n264007 );
and ( n264010 , n264009 , n256649 );
nor ( n264011 , n264008 , n264010 );
not ( n264012 , n264011 );
not ( n264013 , n256152 );
not ( n264014 , n232726 );
not ( n264015 , n237443 );
or ( n264016 , n264014 , n264015 );
not ( n264017 , n232726 );
nand ( n264018 , n237444 , n264017 );
nand ( n264019 , n264016 , n264018 );
not ( n264020 , n264019 );
and ( n264021 , n264013 , n264020 );
and ( n264022 , n237591 , n264019 );
nor ( n264023 , n264021 , n264022 );
nand ( n264024 , n264012 , n264023 );
not ( n264025 , n51421 );
not ( n264026 , n239653 );
or ( n264027 , n264025 , n264026 );
not ( n264028 , n51421 );
nand ( n264029 , n264028 , n244125 );
nand ( n264030 , n264027 , n264029 );
and ( n264031 , n264030 , n45873 );
not ( n264032 , n264030 );
and ( n264033 , n264032 , n45876 );
nor ( n264034 , n264031 , n264033 );
not ( n264035 , n264034 );
nor ( n264036 , n264035 , n226955 );
not ( n264037 , n264036 );
or ( n264038 , n264024 , n264037 );
nand ( n264039 , n264034 , n264023 );
nand ( n264040 , n264039 , n264011 , n260879 );
nand ( n264041 , n247585 , n44132 );
nand ( n264042 , n264038 , n264040 , n264041 );
buf ( n264043 , n264042 );
not ( n264044 , n251009 );
not ( n264045 , n260640 );
or ( n264046 , n264044 , n264045 );
not ( n264047 , n251009 );
nand ( n264048 , n264047 , n263336 );
nand ( n264049 , n264046 , n264048 );
and ( n264050 , n264049 , n263339 );
not ( n264051 , n264049 );
and ( n264052 , n264051 , n260644 );
nor ( n264053 , n264050 , n264052 );
not ( n264054 , n264053 );
nor ( n264055 , n264054 , n46425 );
not ( n264056 , n264055 );
not ( n264057 , n240306 );
not ( n264058 , n264057 );
not ( n264059 , n252051 );
or ( n264060 , n264058 , n264059 );
not ( n264061 , n264057 );
nand ( n264062 , n264061 , n252036 );
nand ( n264063 , n264060 , n264062 );
and ( n264064 , n264063 , n256227 );
not ( n264065 , n264063 );
and ( n264066 , n264065 , n254223 );
nor ( n264067 , n264064 , n264066 );
not ( n264068 , n264067 );
not ( n264069 , n248178 );
not ( n264070 , n240001 );
or ( n264071 , n264069 , n264070 );
not ( n264072 , n248178 );
nand ( n264073 , n264072 , n239994 );
nand ( n264074 , n264071 , n264073 );
not ( n264075 , n240053 );
and ( n264076 , n264074 , n264075 );
not ( n264077 , n264074 );
and ( n264078 , n264077 , n240053 );
nor ( n264079 , n264076 , n264078 );
not ( n264080 , n264079 );
nand ( n264081 , n264068 , n264080 );
or ( n264082 , n264056 , n264081 );
not ( n264083 , n264053 );
not ( n264084 , n264068 );
or ( n264085 , n264083 , n264084 );
nor ( n264086 , n264080 , n40465 );
nand ( n264087 , n264085 , n264086 );
nand ( n264088 , n237361 , n33586 );
nand ( n264089 , n264082 , n264087 , n264088 );
buf ( n264090 , n264089 );
nand ( n264091 , n252066 , n33255 );
not ( n264092 , n45246 );
not ( n264093 , n244054 );
or ( n264094 , n264092 , n264093 );
not ( n264095 , n45246 );
nand ( n264096 , n264095 , n253557 );
nand ( n264097 , n264094 , n264096 );
not ( n264098 , n257706 );
and ( n264099 , n264097 , n264098 );
not ( n264100 , n264097 );
not ( n264101 , n257703 );
and ( n264102 , n264100 , n264101 );
nor ( n264103 , n264099 , n264102 );
not ( n264104 , n251400 );
not ( n264105 , n252132 );
or ( n264106 , n264104 , n264105 );
not ( n264107 , n251400 );
nand ( n264108 , n264107 , n252139 );
nand ( n264109 , n264106 , n264108 );
and ( n264110 , n264109 , n252194 );
not ( n264111 , n264109 );
and ( n264112 , n264111 , n252186 );
nor ( n264113 , n264110 , n264112 );
nand ( n264114 , n264103 , n264113 );
or ( n264115 , n264091 , n264114 );
not ( n264116 , n252066 );
not ( n264117 , n264113 );
or ( n264118 , n264116 , n264117 );
nor ( n264119 , n264103 , n49051 );
nand ( n264120 , n264118 , n264119 );
nand ( n264121 , n236798 , n205079 );
nand ( n264122 , n264115 , n264120 , n264121 );
buf ( n264123 , n264122 );
nor ( n264124 , n235891 , n255647 );
nand ( n264125 , n55105 , n264124 );
not ( n264126 , n232864 );
not ( n264127 , n255647 );
nand ( n264128 , n264126 , n264127 );
nand ( n264129 , n264128 , n235891 , n256584 );
nand ( n264130 , n247585 , n33557 );
nand ( n264131 , n264125 , n264129 , n264130 );
buf ( n264132 , n264131 );
not ( n264133 , RI19ac0158_2331);
or ( n264134 , n25328 , n264133 );
not ( n264135 , RI19ab71e8_2401);
or ( n264136 , n25335 , n264135 );
nand ( n264137 , n264134 , n264136 );
buf ( n264138 , n264137 );
not ( n264139 , RI19abebc8_2343);
or ( n264140 , n25328 , n264139 );
not ( n264141 , RI19ab5640_2413);
or ( n264142 , n25335 , n264141 );
nand ( n264143 , n264140 , n264142 );
buf ( n264144 , n264143 );
not ( n264145 , n261002 );
nand ( n264146 , n261006 , n264145 );
or ( n264147 , n256958 , n264146 );
nor ( n264148 , n256956 , n235050 );
nand ( n264149 , n264148 , n264146 );
nand ( n264150 , n35431 , n220505 );
nand ( n264151 , n264147 , n264149 , n264150 );
buf ( n264152 , n264151 );
not ( n264153 , n28789 );
not ( n264154 , n244073 );
or ( n264155 , n264153 , n264154 );
not ( n264156 , n253849 );
not ( n264157 , n46506 );
or ( n264158 , n264156 , n264157 );
not ( n264159 , n253849 );
nand ( n264160 , n264159 , n46514 );
nand ( n264161 , n264158 , n264160 );
and ( n264162 , n264161 , n224478 );
not ( n264163 , n264161 );
and ( n264164 , n264163 , n251333 );
nor ( n264165 , n264162 , n264164 );
nand ( n264166 , n264165 , n261146 );
not ( n264167 , n261135 );
and ( n264168 , n264166 , n264167 );
not ( n264169 , n264166 );
and ( n264170 , n264169 , n261135 );
nor ( n264171 , n264168 , n264170 );
or ( n264172 , n264171 , n254515 );
nand ( n264173 , n264155 , n264172 );
buf ( n264174 , n264173 );
not ( n264175 , n31150 );
not ( n264176 , n237361 );
or ( n264177 , n264175 , n264176 );
not ( n264178 , n245423 );
not ( n264179 , n241962 );
or ( n264180 , n264178 , n264179 );
not ( n264181 , n245423 );
nand ( n264182 , n264181 , n250439 );
nand ( n264183 , n264180 , n264182 );
and ( n264184 , n264183 , n257572 );
not ( n264185 , n264183 );
and ( n264186 , n264185 , n250498 );
nor ( n264187 , n264184 , n264186 );
not ( n264188 , n245654 );
not ( n264189 , n241448 );
not ( n264190 , n264189 );
or ( n264191 , n264188 , n264190 );
not ( n264192 , n245654 );
nand ( n264193 , n264192 , n243687 );
nand ( n264194 , n264191 , n264193 );
and ( n264195 , n264194 , n234881 );
not ( n264196 , n264194 );
not ( n264197 , n234881 );
and ( n264198 , n264196 , n264197 );
nor ( n264199 , n264195 , n264198 );
nand ( n264200 , n264187 , n264199 );
not ( n264201 , n255798 );
not ( n264202 , n246548 );
or ( n264203 , n264201 , n264202 );
not ( n264204 , n255798 );
nand ( n264205 , n264204 , n246553 );
nand ( n264206 , n264203 , n264205 );
and ( n264207 , n264206 , n246661 );
not ( n264208 , n264206 );
and ( n264209 , n264208 , n246654 );
nor ( n264210 , n264207 , n264209 );
not ( n264211 , n264210 );
and ( n264212 , n264200 , n264211 );
not ( n264213 , n264200 );
and ( n264214 , n264213 , n264210 );
nor ( n264215 , n264212 , n264214 );
or ( n264216 , n264215 , n254882 );
nand ( n264217 , n264177 , n264216 );
buf ( n264218 , n264217 );
or ( n264219 , n25328 , n253221 );
not ( n264220 , RI19ac8510_2267);
or ( n264221 , n25335 , n264220 );
nand ( n264222 , n264219 , n264221 );
buf ( n264223 , n264222 );
buf ( n264224 , n29681 );
buf ( n264225 , n33278 );
buf ( n264226 , n32713 );
not ( n264227 , n32295 );
not ( n264228 , n234453 );
or ( n264229 , n264227 , n264228 );
not ( n264230 , n49454 );
not ( n264231 , n247187 );
or ( n264232 , n264230 , n264231 );
not ( n264233 , n49454 );
nand ( n264234 , n264233 , n247195 );
nand ( n264235 , n264232 , n264234 );
and ( n264236 , n264235 , n254400 );
not ( n264237 , n264235 );
and ( n264238 , n264237 , n254403 );
nor ( n264239 , n264236 , n264238 );
not ( n264240 , n264239 );
nand ( n264241 , n264240 , n252737 );
not ( n264242 , n48303 );
not ( n264243 , n254947 );
or ( n264244 , n264242 , n264243 );
not ( n264245 , n48303 );
nand ( n264246 , n264245 , n245677 );
nand ( n264247 , n264244 , n264246 );
and ( n264248 , n264247 , n254974 );
not ( n264249 , n264247 );
and ( n264250 , n264249 , n260823 );
nor ( n264251 , n264248 , n264250 );
not ( n264252 , n264251 );
and ( n264253 , n264241 , n264252 );
not ( n264254 , n264241 );
and ( n264255 , n264254 , n264251 );
nor ( n264256 , n264253 , n264255 );
not ( n264257 , n234111 );
or ( n264258 , n264256 , n264257 );
nand ( n264259 , n264229 , n264258 );
buf ( n264260 , n264259 );
or ( n264261 , n25328 , n257469 );
not ( n264262 , RI19ac1148_2322);
or ( n264263 , n25335 , n264262 );
nand ( n264264 , n264261 , n264263 );
buf ( n264265 , n264264 );
not ( n264266 , n245898 );
not ( n264267 , n52982 );
or ( n264268 , n264266 , n264267 );
not ( n264269 , n245898 );
nand ( n264270 , n264269 , n52989 );
nand ( n264271 , n264268 , n264270 );
and ( n264272 , n264271 , n52997 );
not ( n264273 , n264271 );
and ( n264274 , n264273 , n52996 );
nor ( n264275 , n264272 , n264274 );
nand ( n264276 , n264275 , n239934 );
nand ( n264277 , n260959 , n260971 );
or ( n264278 , n264276 , n264277 );
not ( n264279 , n260971 );
not ( n264280 , n264275 );
or ( n264281 , n264279 , n264280 );
nor ( n264282 , n260959 , n46425 );
nand ( n264283 , n264281 , n264282 );
nand ( n264284 , n55760 , n27985 );
nand ( n264285 , n264278 , n264283 , n264284 );
buf ( n264286 , n264285 );
not ( n264287 , RI19abd188_2358);
or ( n264288 , n25328 , n264287 );
not ( n264289 , RI19ab3318_2430);
or ( n264290 , n25335 , n264289 );
nand ( n264291 , n264288 , n264290 );
buf ( n264292 , n264291 );
not ( n264293 , n257802 );
nand ( n264294 , n264293 , n250826 );
or ( n264295 , n257793 , n264294 );
not ( n264296 , n264293 );
not ( n264297 , n250750 );
or ( n264298 , n264296 , n264297 );
nand ( n264299 , n264298 , n253905 );
nand ( n264300 , n251465 , n204432 );
nand ( n264301 , n264295 , n264299 , n264300 );
buf ( n264302 , n264301 );
not ( n264303 , n252123 );
not ( n264304 , n47319 );
or ( n264305 , n264303 , n264304 );
or ( n264306 , n47319 , n252123 );
nand ( n264307 , n264305 , n264306 );
and ( n264308 , n264307 , n225086 );
not ( n264309 , n264307 );
and ( n264310 , n264309 , n225083 );
nor ( n264311 , n264308 , n264310 );
not ( n264312 , n264311 );
nor ( n264313 , n264312 , n260567 );
not ( n264314 , n264313 );
not ( n264315 , n36253 );
not ( n264316 , n249757 );
or ( n264317 , n264315 , n264316 );
not ( n264318 , n36253 );
nand ( n264319 , n264318 , n249749 );
nand ( n264320 , n264317 , n264319 );
and ( n264321 , n264320 , n254644 );
not ( n264322 , n264320 );
and ( n264323 , n264322 , n254647 );
nor ( n264324 , n264321 , n264323 );
not ( n264325 , n264324 );
not ( n264326 , n46067 );
not ( n264327 , n51571 );
not ( n264328 , n45873 );
or ( n264329 , n264327 , n264328 );
or ( n264330 , n45873 , n51571 );
nand ( n264331 , n264329 , n264330 );
not ( n264332 , n264331 );
or ( n264333 , n264326 , n264332 );
or ( n264334 , n264331 , n241701 );
nand ( n264335 , n264333 , n264334 );
not ( n264336 , n264335 );
nand ( n264337 , n264325 , n264336 );
or ( n264338 , n264314 , n264337 );
not ( n264339 , n264325 );
not ( n264340 , n264311 );
or ( n264341 , n264339 , n264340 );
not ( n264342 , n250111 );
nor ( n264343 , n264342 , n264336 );
nand ( n264344 , n264341 , n264343 );
nand ( n264345 , n31577 , n218281 );
nand ( n264346 , n264338 , n264344 , n264345 );
buf ( n264347 , n264346 );
not ( n264348 , n263615 );
not ( n264349 , n264348 );
not ( n264350 , n257021 );
or ( n264351 , n264349 , n264350 );
nor ( n264352 , n257012 , n247276 );
nand ( n264353 , n264351 , n264352 );
nor ( n264354 , n263615 , n238900 );
nand ( n264355 , n264354 , n257021 , n257012 );
nand ( n264356 , n35431 , n40162 );
nand ( n264357 , n264353 , n264355 , n264356 );
buf ( n264358 , n264357 );
not ( n264359 , RI19aae110_2467);
or ( n264360 , n25328 , n264359 );
or ( n264361 , n25335 , n254046 );
nand ( n264362 , n264360 , n264361 );
buf ( n264363 , n264362 );
buf ( n264364 , n34365 );
buf ( n264365 , n37937 );
not ( n264366 , n238372 );
not ( n264367 , n254337 );
or ( n264368 , n264366 , n264367 );
not ( n264369 , n238372 );
nand ( n264370 , n264369 , n254344 );
nand ( n264371 , n264368 , n264370 );
and ( n264372 , n264371 , n256649 );
not ( n264373 , n264371 );
and ( n264374 , n264373 , n256646 );
nor ( n264375 , n264372 , n264374 );
buf ( n264376 , n245147 );
not ( n264377 , n264376 );
not ( n264378 , n40914 );
or ( n264379 , n264377 , n264378 );
or ( n264380 , n40918 , n264376 );
nand ( n264381 , n264379 , n264380 );
not ( n264382 , n264381 );
not ( n264383 , n218981 );
not ( n264384 , n264383 );
and ( n264385 , n264382 , n264384 );
and ( n264386 , n264381 , n41217 );
nor ( n264387 , n264385 , n264386 );
nand ( n264388 , n264375 , n264387 );
not ( n264389 , n257290 );
or ( n264390 , n264388 , n264389 );
not ( n264391 , n257285 );
not ( n264392 , n264375 );
or ( n264393 , n264391 , n264392 );
nor ( n264394 , n264387 , n254150 );
nand ( n264395 , n264393 , n264394 );
nand ( n264396 , n39767 , n26086 );
nand ( n264397 , n264390 , n264395 , n264396 );
buf ( n264398 , n264397 );
buf ( n264399 , n38543 );
not ( n264400 , RI19a846f8_2763);
or ( n264401 , n25328 , n264400 );
not ( n264402 , RI19ac9500_2260);
or ( n264403 , n226822 , n264402 );
nand ( n264404 , n264401 , n264403 );
buf ( n264405 , n264404 );
buf ( n264406 , n29515 );
not ( n264407 , n33254 );
not ( n264408 , n253927 );
nand ( n264409 , n264407 , n264408 );
not ( n264410 , n245881 );
not ( n264411 , n264410 );
not ( n264412 , n52982 );
or ( n264413 , n264411 , n264412 );
not ( n264414 , n264410 );
nand ( n264415 , n264414 , n52989 );
nand ( n264416 , n264413 , n264415 );
and ( n264417 , n264416 , n52996 );
not ( n264418 , n264416 );
and ( n264419 , n264418 , n52997 );
nor ( n264420 , n264417 , n264419 );
not ( n264421 , n252000 );
not ( n264422 , n49617 );
or ( n264423 , n264421 , n264422 );
not ( n264424 , n252000 );
nand ( n264425 , n264424 , n49626 );
nand ( n264426 , n264423 , n264425 );
and ( n264427 , n264426 , n253272 );
not ( n264428 , n264426 );
and ( n264429 , n264428 , n253265 );
nor ( n264430 , n264427 , n264429 );
nand ( n264431 , n264420 , n264430 );
or ( n264432 , n264409 , n264431 );
not ( n264433 , n253929 );
nand ( n264434 , n264433 , n264431 );
nand ( n264435 , n51381 , n205295 );
nand ( n264436 , n264432 , n264434 , n264435 );
buf ( n264437 , n264436 );
not ( n264438 , n29546 );
not ( n264439 , n41945 );
or ( n264440 , n264438 , n264439 );
not ( n264441 , n259206 );
not ( n264442 , n250229 );
or ( n264443 , n264441 , n264442 );
not ( n264444 , n259206 );
nand ( n264445 , n264444 , n259150 );
nand ( n264446 , n264443 , n264445 );
and ( n264447 , n264446 , n250942 );
not ( n264448 , n264446 );
and ( n264449 , n264448 , n259153 );
nor ( n264450 , n264447 , n264449 );
not ( n264451 , n264450 );
buf ( n264452 , n49985 );
not ( n264453 , n264452 );
not ( n264454 , n48883 );
or ( n264455 , n264453 , n264454 );
or ( n264456 , n48883 , n264452 );
nand ( n264457 , n264455 , n264456 );
not ( n264458 , n264457 );
not ( n264459 , n246479 );
and ( n264460 , n264458 , n264459 );
and ( n264461 , n264457 , n246479 );
nor ( n264462 , n264460 , n264461 );
nand ( n264463 , n264451 , n264462 );
and ( n264464 , n264463 , n247579 );
not ( n264465 , n264463 );
not ( n264466 , n247579 );
and ( n264467 , n264465 , n264466 );
nor ( n264468 , n264464 , n264467 );
not ( n264469 , n222532 );
or ( n264470 , n264468 , n264469 );
nand ( n264471 , n264440 , n264470 );
buf ( n264472 , n264471 );
not ( n264473 , n255231 );
not ( n264474 , n240656 );
not ( n264475 , n247393 );
or ( n264476 , n264474 , n264475 );
nand ( n264477 , n247399 , n240657 );
nand ( n264478 , n264476 , n264477 );
not ( n264479 , n264478 );
not ( n264480 , n247349 );
and ( n264481 , n264479 , n264480 );
and ( n264482 , n264478 , n247349 );
nor ( n264483 , n264481 , n264482 );
not ( n264484 , n264483 );
or ( n264485 , n264473 , n264484 );
not ( n264486 , n245888 );
not ( n264487 , n52982 );
or ( n264488 , n264486 , n264487 );
not ( n264489 , n245888 );
nand ( n264490 , n264489 , n52989 );
nand ( n264491 , n264488 , n264490 );
and ( n264492 , n264491 , n52997 );
not ( n264493 , n264491 );
and ( n264494 , n264493 , n52996 );
nor ( n264495 , n264492 , n264494 );
not ( n264496 , n264495 );
nor ( n264497 , n264496 , n258327 );
nand ( n264498 , n264485 , n264497 );
nand ( n264499 , n255206 , n264483 , n264496 );
nand ( n264500 , n50615 , n36335 );
nand ( n264501 , n264498 , n264499 , n264500 );
buf ( n264502 , n264501 );
not ( n264503 , n43945 );
not ( n264504 , n264503 );
not ( n264505 , n252552 );
or ( n264506 , n264504 , n264505 );
not ( n264507 , n264503 );
nand ( n264508 , n264507 , n252561 );
nand ( n264509 , n264506 , n264508 );
and ( n264510 , n264509 , n255676 );
not ( n264511 , n264509 );
and ( n264512 , n264511 , n255673 );
nor ( n264513 , n264510 , n264512 );
buf ( n264514 , n221994 );
not ( n264515 , n264514 );
not ( n264516 , n234106 );
or ( n264517 , n264515 , n264516 );
or ( n264518 , n234106 , n264514 );
nand ( n264519 , n264517 , n264518 );
and ( n264520 , n264519 , n249463 );
not ( n264521 , n264519 );
and ( n264522 , n264521 , n249470 );
nor ( n264523 , n264520 , n264522 );
not ( n264524 , n264523 );
nand ( n264525 , n264513 , n264524 );
not ( n264526 , n49768 );
not ( n264527 , n246693 );
or ( n264528 , n264526 , n264527 );
or ( n264529 , n246693 , n49768 );
nand ( n264530 , n264528 , n264529 );
and ( n264531 , n264530 , n259744 );
not ( n264532 , n264530 );
and ( n264533 , n264532 , n259747 );
nor ( n264534 , n264531 , n264533 );
nand ( n264535 , n264534 , n222532 );
or ( n264536 , n264525 , n264535 );
nor ( n264537 , n264534 , n37725 );
nand ( n264538 , n264525 , n264537 );
nand ( n264539 , n262000 , n33069 );
nand ( n264540 , n264536 , n264538 , n264539 );
buf ( n264541 , n264540 );
not ( n264542 , RI19ab6900_2405);
or ( n264543 , n25328 , n264542 );
or ( n264544 , n25335 , n263872 );
nand ( n264545 , n264543 , n264544 );
buf ( n264546 , n264545 );
not ( n264547 , n248190 );
not ( n264548 , n264547 );
not ( n264549 , n240001 );
or ( n264550 , n264548 , n264549 );
not ( n264551 , n264547 );
nand ( n264552 , n264551 , n239994 );
nand ( n264553 , n264550 , n264552 );
and ( n264554 , n264553 , n240057 );
not ( n264555 , n264553 );
and ( n264556 , n264555 , n240053 );
nor ( n264557 , n264554 , n264556 );
not ( n264558 , n264557 );
not ( n264559 , n256830 );
not ( n264560 , n264559 );
not ( n264561 , n208725 );
or ( n264562 , n264560 , n264561 );
not ( n264563 , n264559 );
nand ( n264564 , n264563 , n30968 );
nand ( n264565 , n264562 , n264564 );
and ( n264566 , n264565 , n31561 );
not ( n264567 , n264565 );
and ( n264568 , n264567 , n31552 );
nor ( n264569 , n264566 , n264568 );
nand ( n264570 , n264558 , n264569 );
or ( n264571 , n240815 , n264570 );
not ( n264572 , n264558 );
not ( n264573 , n240814 );
or ( n264574 , n264572 , n264573 );
nor ( n264575 , n264569 , n250431 );
nand ( n264576 , n264574 , n264575 );
nand ( n264577 , n35431 , n25902 );
nand ( n264578 , n264571 , n264576 , n264577 );
buf ( n264579 , n264578 );
not ( n264580 , n239237 );
nand ( n264581 , n264580 , n259157 );
nand ( n264582 , n256180 , n256197 );
or ( n264583 , n264581 , n264582 );
not ( n264584 , n256197 );
not ( n264585 , n259157 );
or ( n264586 , n264584 , n264585 );
nor ( n264587 , n256180 , n247698 );
nand ( n264588 , n264586 , n264587 );
nand ( n264589 , n251712 , n38055 );
nand ( n264590 , n264583 , n264588 , n264589 );
buf ( n264591 , n264590 );
not ( n264592 , n246921 );
not ( n264593 , n256190 );
or ( n264594 , n264592 , n264593 );
not ( n264595 , n246921 );
nand ( n264596 , n264595 , n256191 );
nand ( n264597 , n264594 , n264596 );
and ( n264598 , n264597 , n260022 );
not ( n264599 , n264597 );
buf ( n264600 , n242148 );
and ( n264601 , n264599 , n264600 );
nor ( n264602 , n264598 , n264601 );
not ( n264603 , n264602 );
nor ( n264604 , n264603 , n39763 );
not ( n264605 , n264604 );
not ( n264606 , n234712 );
not ( n264607 , n261830 );
or ( n264608 , n264606 , n264607 );
not ( n264609 , n234712 );
nand ( n264610 , n264609 , n261834 );
nand ( n264611 , n264608 , n264610 );
and ( n264612 , n264611 , n242683 );
not ( n264613 , n264611 );
and ( n264614 , n264613 , n242680 );
nor ( n264615 , n264612 , n264614 );
not ( n264616 , n264615 );
not ( n264617 , n48917 );
not ( n264618 , n264617 );
not ( n264619 , n254603 );
or ( n264620 , n264618 , n264619 );
not ( n264621 , n264617 );
nand ( n264622 , n264621 , n254594 );
nand ( n264623 , n264620 , n264622 );
and ( n264624 , n264623 , n254611 );
not ( n264625 , n264623 );
not ( n264626 , n251627 );
not ( n264627 , n264626 );
and ( n264628 , n264625 , n264627 );
nor ( n264629 , n264624 , n264628 );
nand ( n264630 , n264616 , n264629 );
or ( n264631 , n264605 , n264630 );
nand ( n264632 , n264602 , n264629 );
nand ( n264633 , n264632 , n264615 , n233973 );
nand ( n264634 , n48251 , n204737 );
nand ( n264635 , n264631 , n264633 , n264634 );
buf ( n264636 , n264635 );
not ( n264637 , RI19ab96f0_2385);
or ( n264638 , n25328 , n264637 );
not ( n264639 , RI19aafad8_2456);
or ( n264640 , n226822 , n264639 );
nand ( n264641 , n264638 , n264640 );
buf ( n264642 , n264641 );
not ( n264643 , n248045 );
not ( n264644 , n264643 );
not ( n264645 , n238792 );
or ( n264646 , n264644 , n264645 );
or ( n264647 , n238792 , n264643 );
nand ( n264648 , n264646 , n264647 );
and ( n264649 , n264648 , n238895 );
not ( n264650 , n264648 );
and ( n264651 , n264650 , n258233 );
nor ( n264652 , n264649 , n264651 );
nor ( n264653 , n264652 , n55146 );
not ( n264654 , n246393 );
not ( n264655 , n264654 );
not ( n264656 , n256742 );
or ( n264657 , n264655 , n264656 );
not ( n264658 , n264654 );
nand ( n264659 , n264658 , n256738 );
nand ( n264660 , n264657 , n264659 );
and ( n264661 , n264660 , n228527 );
not ( n264662 , n264660 );
and ( n264663 , n264662 , n261630 );
nor ( n264664 , n264661 , n264663 );
not ( n264665 , n248716 );
not ( n264666 , n264665 );
not ( n264667 , n55725 );
or ( n264668 , n264666 , n264667 );
not ( n264669 , n264665 );
nand ( n264670 , n264669 , n55724 );
nand ( n264671 , n264668 , n264670 );
buf ( n264672 , n241050 );
and ( n264673 , n264671 , n264672 );
not ( n264674 , n264671 );
not ( n264675 , n264672 );
and ( n264676 , n264674 , n264675 );
nor ( n264677 , n264673 , n264676 );
nand ( n264678 , n264653 , n264664 , n264677 );
not ( n264679 , n264652 );
not ( n264680 , n264679 );
not ( n264681 , n264677 );
or ( n264682 , n264680 , n264681 );
nor ( n264683 , n264664 , n235895 );
nand ( n264684 , n264682 , n264683 );
nand ( n264685 , n35431 , n44724 );
nand ( n264686 , n264678 , n264684 , n264685 );
buf ( n264687 , n264686 );
not ( n264688 , n37624 );
not ( n264689 , n51381 );
or ( n264690 , n264688 , n264689 );
not ( n264691 , n239066 );
not ( n264692 , n52221 );
or ( n264693 , n264691 , n264692 );
not ( n264694 , n239066 );
nand ( n264695 , n264694 , n52229 );
nand ( n264696 , n264693 , n264695 );
and ( n264697 , n264696 , n259264 );
not ( n264698 , n264696 );
buf ( n264699 , n246385 );
not ( n264700 , n264699 );
and ( n264701 , n264698 , n264700 );
nor ( n264702 , n264697 , n264701 );
not ( n264703 , n252887 );
not ( n264704 , n241050 );
not ( n264705 , n264704 );
not ( n264706 , n264705 );
or ( n264707 , n264703 , n264706 );
not ( n264708 , n252887 );
nand ( n264709 , n264708 , n264704 );
nand ( n264710 , n264707 , n264709 );
and ( n264711 , n264710 , n241060 );
not ( n264712 , n264710 );
and ( n264713 , n264712 , n241057 );
nor ( n264714 , n264711 , n264713 );
nand ( n264715 , n264702 , n264714 );
not ( n264716 , n206371 );
not ( n264717 , n254866 );
or ( n264718 , n264716 , n264717 );
not ( n264719 , n206371 );
nand ( n264720 , n264719 , n254873 );
nand ( n264721 , n264718 , n264720 );
and ( n264722 , n264721 , n256712 );
not ( n264723 , n264721 );
and ( n264724 , n264723 , n256716 );
nor ( n264725 , n264722 , n264724 );
not ( n264726 , n264725 );
and ( n264727 , n264715 , n264726 );
not ( n264728 , n264715 );
and ( n264729 , n264728 , n264725 );
nor ( n264730 , n264727 , n264729 );
or ( n264731 , n264730 , n258327 );
nand ( n264732 , n264690 , n264731 );
buf ( n264733 , n264732 );
not ( n264734 , RI19aa38c8_2541);
or ( n264735 , n25328 , n264734 );
not ( n264736 , RI19a9a160_2611);
or ( n264737 , n25335 , n264736 );
nand ( n264738 , n264735 , n264737 );
buf ( n264739 , n264738 );
not ( n264740 , n247946 );
not ( n264741 , n239922 );
or ( n264742 , n264740 , n264741 );
or ( n264743 , n239922 , n247946 );
nand ( n264744 , n264742 , n264743 );
not ( n264745 , n264744 );
not ( n264746 , n243511 );
and ( n264747 , n264745 , n264746 );
and ( n264748 , n264744 , n243511 );
nor ( n264749 , n264747 , n264748 );
nor ( n264750 , n264749 , n49051 );
not ( n264751 , n264750 );
nand ( n264752 , n260802 , n260830 );
or ( n264753 , n264751 , n264752 );
not ( n264754 , n260802 );
not ( n264755 , n264749 );
not ( n264756 , n264755 );
or ( n264757 , n264754 , n264756 );
nor ( n264758 , n260830 , n33254 );
nand ( n264759 , n264757 , n264758 );
nand ( n264760 , n237714 , n37851 );
nand ( n264761 , n264753 , n264759 , n264760 );
buf ( n264762 , n264761 );
not ( n264763 , n30790 );
not ( n264764 , n245702 );
or ( n264765 , n264763 , n264764 );
not ( n264766 , n260100 );
not ( n264767 , n251525 );
or ( n264768 , n264766 , n264767 );
not ( n264769 , n260100 );
nand ( n264770 , n264769 , n251526 );
nand ( n264771 , n264768 , n264770 );
not ( n264772 , n264771 );
not ( n264773 , n249757 );
or ( n264774 , n264772 , n264773 );
or ( n264775 , n251532 , n264771 );
nand ( n264776 , n264774 , n264775 );
nand ( n264777 , n264776 , n254065 );
and ( n264778 , n264777 , n254095 );
not ( n264779 , n264777 );
and ( n264780 , n264779 , n254098 );
nor ( n264781 , n264778 , n264780 );
or ( n264782 , n264781 , n260760 );
nand ( n264783 , n264765 , n264782 );
buf ( n264784 , n264783 );
not ( n264785 , n241924 );
not ( n264786 , n264785 );
not ( n264787 , n259905 );
or ( n264788 , n264786 , n264787 );
not ( n264789 , n264785 );
nand ( n264790 , n264789 , n237590 );
nand ( n264791 , n264788 , n264790 );
and ( n264792 , n264791 , n259578 );
not ( n264793 , n264791 );
and ( n264794 , n264793 , n259575 );
nor ( n264795 , n264792 , n264794 );
not ( n264796 , n261389 );
nand ( n264797 , n264795 , n264796 );
not ( n264798 , n256027 );
or ( n264799 , n264797 , n264798 );
not ( n264800 , n256026 );
not ( n264801 , n264800 );
not ( n264802 , n264795 );
or ( n264803 , n264801 , n264802 );
nor ( n264804 , n264796 , n35427 );
nand ( n264805 , n264803 , n264804 );
nand ( n264806 , n241976 , n25514 );
nand ( n264807 , n264799 , n264805 , n264806 );
buf ( n264808 , n264807 );
buf ( n264809 , n35877 );
buf ( n264810 , n35304 );
buf ( n264811 , n32162 );
buf ( n264812 , n41136 );
buf ( n264813 , n31857 );
buf ( n264814 , n25922 );
buf ( n264815 , n30266 );
buf ( n264816 , n39626 );
not ( n264817 , n226763 );
not ( n264818 , n254603 );
or ( n264819 , n264817 , n264818 );
not ( n264820 , n226763 );
nand ( n264821 , n264820 , n254594 );
nand ( n264822 , n264819 , n264821 );
and ( n264823 , n264822 , n264627 );
not ( n264824 , n264822 );
and ( n264825 , n264824 , n254608 );
nor ( n264826 , n264823 , n264825 );
not ( n264827 , n264826 );
nor ( n264828 , n264827 , n244399 );
not ( n264829 , n249309 );
not ( n264830 , n235202 );
or ( n264831 , n264829 , n264830 );
not ( n264832 , n249309 );
nand ( n264833 , n264832 , n235211 );
nand ( n264834 , n264831 , n264833 );
xor ( n264835 , n264834 , n250721 );
nand ( n264836 , n264828 , n264835 , n257584 );
not ( n264837 , n264826 );
not ( n264838 , n264835 );
or ( n264839 , n264837 , n264838 );
nor ( n264840 , n257584 , n33254 );
nand ( n264841 , n264839 , n264840 );
nand ( n264842 , n35431 , n31404 );
nand ( n264843 , n264836 , n264841 , n264842 );
buf ( n264844 , n264843 );
buf ( n264845 , n29658 );
buf ( n264846 , n39485 );
buf ( n264847 , n30625 );
buf ( n264848 , n33793 );
buf ( n264849 , n209798 );
not ( n264850 , n258814 );
not ( n264851 , n264850 );
not ( n264852 , n258828 );
or ( n264853 , n264851 , n264852 );
and ( n264854 , n48527 , n254973 );
not ( n264855 , n48527 );
and ( n264856 , n264855 , n263294 );
nor ( n264857 , n264854 , n264856 );
and ( n264858 , n264857 , n262633 );
not ( n264859 , n264857 );
and ( n264860 , n264859 , n263297 );
nor ( n264861 , n264858 , n264860 );
nor ( n264862 , n264861 , n252872 );
nand ( n264863 , n264853 , n264862 );
nor ( n264864 , n258814 , n243434 );
nand ( n264865 , n264864 , n264861 , n258828 );
nand ( n264866 , n255116 , n208623 );
nand ( n264867 , n264863 , n264865 , n264866 );
buf ( n264868 , n264867 );
buf ( n264869 , n34792 );
not ( n264870 , n28487 );
not ( n264871 , n255116 );
or ( n264872 , n264870 , n264871 );
not ( n264873 , n46181 );
not ( n264874 , n54195 );
or ( n264875 , n264873 , n264874 );
not ( n264876 , n46181 );
nand ( n264877 , n264876 , n231952 );
nand ( n264878 , n264875 , n264877 );
buf ( n264879 , n248557 );
and ( n264880 , n264878 , n264879 );
not ( n264881 , n264878 );
buf ( n264882 , n248565 );
and ( n264883 , n264881 , n264882 );
nor ( n264884 , n264880 , n264883 );
not ( n264885 , n240141 );
buf ( n264886 , n239138 );
not ( n264887 , n264886 );
and ( n264888 , n264885 , n264887 );
and ( n264889 , n244386 , n264886 );
nor ( n264890 , n264888 , n264889 );
and ( n264891 , n264890 , n255353 );
not ( n264892 , n264890 );
and ( n264893 , n264892 , n255356 );
nor ( n264894 , n264891 , n264893 );
nand ( n264895 , n264884 , n264894 );
not ( n264896 , n264895 );
not ( n264897 , n234999 );
not ( n264898 , n254117 );
or ( n264899 , n264897 , n264898 );
or ( n264900 , n254117 , n234999 );
nand ( n264901 , n264899 , n264900 );
and ( n264902 , n264901 , n254122 );
not ( n264903 , n264901 );
and ( n264904 , n264903 , n254125 );
nor ( n264905 , n264902 , n264904 );
not ( n264906 , n264905 );
and ( n264907 , n264896 , n264906 );
and ( n264908 , n264895 , n264905 );
nor ( n264909 , n264907 , n264908 );
or ( n264910 , n264909 , n244837 );
nand ( n264911 , n264872 , n264910 );
buf ( n264912 , n264911 );
not ( n264913 , n31597 );
not ( n264914 , n31577 );
or ( n264915 , n264913 , n264914 );
not ( n264916 , n242665 );
not ( n264917 , n244939 );
or ( n264918 , n264916 , n264917 );
not ( n264919 , n242665 );
nand ( n264920 , n264919 , n244954 );
nand ( n264921 , n264918 , n264920 );
and ( n264922 , n264921 , n254874 );
not ( n264923 , n264921 );
and ( n264924 , n264923 , n254867 );
nor ( n264925 , n264922 , n264924 );
not ( n264926 , n264925 );
not ( n264927 , n225083 );
not ( n264928 , n252107 );
not ( n264929 , n47310 );
or ( n264930 , n264928 , n264929 );
not ( n264931 , n252107 );
nand ( n264932 , n264931 , n47319 );
nand ( n264933 , n264930 , n264932 );
not ( n264934 , n264933 );
or ( n264935 , n264927 , n264934 );
or ( n264936 , n264933 , n225083 );
nand ( n264937 , n264935 , n264936 );
nand ( n264938 , n264926 , n264937 );
not ( n264939 , n252894 );
not ( n264940 , n241054 );
or ( n264941 , n264939 , n264940 );
or ( n264942 , n241054 , n252894 );
nand ( n264943 , n264941 , n264942 );
and ( n264944 , n264943 , n241057 );
not ( n264945 , n264943 );
and ( n264946 , n264945 , n241060 );
nor ( n264947 , n264944 , n264946 );
not ( n264948 , n264947 );
and ( n264949 , n264938 , n264948 );
not ( n264950 , n264938 );
and ( n264951 , n264950 , n264947 );
nor ( n264952 , n264949 , n264951 );
or ( n264953 , n264952 , n252859 );
nand ( n264954 , n264915 , n264953 );
buf ( n264955 , n264954 );
or ( n264956 , n25328 , n260789 );
not ( n264957 , RI19a8cd80_2705);
or ( n264958 , n226822 , n264957 );
nand ( n264959 , n264956 , n264958 );
buf ( n264960 , n264959 );
not ( n264961 , RI19aad648_2472);
or ( n264962 , n25328 , n264961 );
not ( n264963 , RI19aa3418_2543);
or ( n264964 , n25336 , n264963 );
nand ( n264965 , n264962 , n264964 );
buf ( n264966 , n264965 );
buf ( n264967 , n249260 );
not ( n264968 , n264967 );
not ( n264969 , n264968 );
not ( n264970 , n244889 );
or ( n264971 , n264969 , n264970 );
nand ( n264972 , n244899 , n264967 );
nand ( n264973 , n264971 , n264972 );
not ( n264974 , n264973 );
not ( n264975 , n244940 );
and ( n264976 , n264974 , n264975 );
and ( n264977 , n264973 , n244940 );
nor ( n264978 , n264976 , n264977 );
not ( n264979 , n264978 );
not ( n264980 , n253869 );
nand ( n264981 , n264979 , n264980 );
or ( n264982 , n253818 , n264981 );
nor ( n264983 , n253817 , n236795 );
nand ( n264984 , n264983 , n264981 );
nand ( n264985 , n55760 , n31771 );
nand ( n264986 , n264982 , n264984 , n264985 );
buf ( n264987 , n264986 );
not ( n264988 , n253577 );
not ( n264989 , n40251 );
not ( n264990 , n235878 );
or ( n264991 , n264989 , n264990 );
not ( n264992 , n40251 );
nand ( n264993 , n264992 , n235887 );
nand ( n264994 , n264991 , n264993 );
and ( n264995 , n264994 , n259858 );
not ( n264996 , n264994 );
and ( n264997 , n264996 , n259855 );
nor ( n264998 , n264995 , n264997 );
nand ( n264999 , n264988 , n264998 );
or ( n265000 , n264999 , n253566 );
nor ( n265001 , n253564 , n55152 );
nand ( n265002 , n264999 , n265001 );
nand ( n265003 , n246460 , n34022 );
nand ( n265004 , n265000 , n265002 , n265003 );
buf ( n265005 , n265004 );
not ( n265006 , n27683 );
not ( n265007 , n55760 );
or ( n265008 , n265006 , n265007 );
nand ( n265009 , n258254 , n258265 );
not ( n265010 , n265009 );
not ( n265011 , n253374 );
and ( n265012 , n265010 , n265011 );
and ( n265013 , n265009 , n253374 );
nor ( n265014 , n265012 , n265013 );
or ( n265015 , n265014 , n254515 );
nand ( n265016 , n265008 , n265015 );
buf ( n265017 , n265016 );
not ( n265018 , RI19ac2390_2312);
or ( n265019 , n226819 , n265018 );
not ( n265020 , RI19ab98d0_2384);
or ( n265021 , n25335 , n265020 );
nand ( n265022 , n265019 , n265021 );
buf ( n265023 , n265022 );
not ( n265024 , n49147 );
not ( n265025 , n243426 );
or ( n265026 , n265024 , n265025 );
or ( n265027 , n243426 , n49147 );
nand ( n265028 , n265026 , n265027 );
buf ( n265029 , n247727 );
and ( n265030 , n265028 , n265029 );
not ( n265031 , n265028 );
and ( n265032 , n265031 , n261484 );
nor ( n265033 , n265030 , n265032 );
nand ( n265034 , n265033 , n226010 );
not ( n265035 , n238247 );
not ( n265036 , n260309 );
or ( n265037 , n265035 , n265036 );
not ( n265038 , n238247 );
nand ( n265039 , n265038 , n236166 );
nand ( n265040 , n265037 , n265039 );
and ( n265041 , n265040 , n259172 );
not ( n265042 , n265040 );
and ( n265043 , n265042 , n259160 );
nor ( n265044 , n265041 , n265043 );
not ( n265045 , n247039 );
not ( n265046 , n253578 );
or ( n265047 , n265045 , n265046 );
not ( n265048 , n247039 );
nand ( n265049 , n265048 , n263124 );
nand ( n265050 , n265047 , n265049 );
and ( n265051 , n265050 , n253478 );
not ( n265052 , n265050 );
and ( n265053 , n265052 , n253475 );
nor ( n265054 , n265051 , n265053 );
nor ( n265055 , n265044 , n265054 );
or ( n265056 , n265034 , n265055 );
nor ( n265057 , n265033 , n49051 );
nand ( n265058 , n265057 , n265055 );
nand ( n265059 , n234448 , n34200 );
nand ( n265060 , n265056 , n265058 , n265059 );
buf ( n265061 , n265060 );
not ( n265062 , n205318 );
not ( n265063 , n37728 );
or ( n265064 , n265062 , n265063 );
not ( n265065 , n248992 );
not ( n265066 , n42105 );
not ( n265067 , n234243 );
or ( n265068 , n265066 , n265067 );
not ( n265069 , n42105 );
nand ( n265070 , n265069 , n234252 );
nand ( n265071 , n265068 , n265070 );
and ( n265072 , n265071 , n234299 );
not ( n265073 , n265071 );
and ( n265074 , n265073 , n234306 );
nor ( n265075 , n265072 , n265074 );
not ( n265076 , n265075 );
nand ( n265077 , n265065 , n265076 );
and ( n265078 , n265077 , n257664 );
not ( n265079 , n265077 );
and ( n265080 , n265079 , n257663 );
nor ( n265081 , n265078 , n265080 );
or ( n265082 , n265081 , n257851 );
nand ( n265083 , n265064 , n265082 );
buf ( n265084 , n265083 );
not ( n265085 , n242453 );
not ( n265086 , n241657 );
or ( n265087 , n265085 , n265086 );
not ( n265088 , n242453 );
nand ( n265089 , n265088 , n241656 );
nand ( n265090 , n265087 , n265089 );
and ( n265091 , n265090 , n241662 );
not ( n265092 , n265090 );
and ( n265093 , n265092 , n244826 );
nor ( n265094 , n265091 , n265093 );
nor ( n265095 , n265094 , n50944 );
not ( n265096 , n265095 );
not ( n265097 , n242297 );
not ( n265098 , n39595 );
or ( n265099 , n265097 , n265098 );
nand ( n265100 , n39598 , n242296 );
nand ( n265101 , n265099 , n265100 );
and ( n265102 , n265101 , n217515 );
not ( n265103 , n265101 );
and ( n265104 , n265103 , n234013 );
nor ( n265105 , n265102 , n265104 );
not ( n265106 , n261706 );
nand ( n265107 , n265105 , n265106 );
or ( n265108 , n265096 , n265107 );
not ( n265109 , n265105 );
not ( n265110 , n265094 );
not ( n265111 , n265110 );
or ( n265112 , n265109 , n265111 );
nor ( n265113 , n265106 , n252872 );
nand ( n265114 , n265112 , n265113 );
nand ( n265115 , n41945 , n31846 );
nand ( n265116 , n265108 , n265114 , n265115 );
buf ( n265117 , n265116 );
buf ( n265118 , n34696 );
buf ( n265119 , n34638 );
not ( n265120 , n240702 );
not ( n265121 , n265120 );
not ( n265122 , n247348 );
or ( n265123 , n265121 , n265122 );
not ( n265124 , n265120 );
nand ( n265125 , n265124 , n263230 );
nand ( n265126 , n265123 , n265125 );
and ( n265127 , n265126 , n263235 );
not ( n265128 , n265126 );
and ( n265129 , n265128 , n257952 );
nor ( n265130 , n265127 , n265129 );
nand ( n265131 , n235044 , n265130 );
or ( n265132 , n263393 , n265131 );
not ( n265133 , n235044 );
not ( n265134 , n234893 );
or ( n265135 , n265133 , n265134 );
nor ( n265136 , n265130 , n234021 );
nand ( n265137 , n265135 , n265136 );
nand ( n265138 , n37728 , n46571 );
nand ( n265139 , n265132 , n265137 , n265138 );
buf ( n265140 , n265139 );
not ( n265141 , RI19aaaa38_2491);
or ( n265142 , n25328 , n265141 );
or ( n265143 , n25336 , n260787 );
nand ( n265144 , n265142 , n265143 );
buf ( n265145 , n265144 );
nand ( n265146 , n252692 , n263556 );
nand ( n265147 , n252702 , n243233 );
or ( n265148 , n265146 , n265147 );
not ( n265149 , n252702 );
not ( n265150 , n252692 );
or ( n265151 , n265149 , n265150 );
nor ( n265152 , n263556 , n251361 );
nand ( n265153 , n265151 , n265152 );
nand ( n265154 , n237714 , n35048 );
nand ( n265155 , n265148 , n265153 , n265154 );
buf ( n265156 , n265155 );
not ( n265157 , n53802 );
not ( n265158 , n238288 );
or ( n265159 , n265157 , n265158 );
not ( n265160 , n53802 );
nand ( n265161 , n265160 , n238297 );
nand ( n265162 , n265159 , n265161 );
and ( n265163 , n265162 , n238401 );
not ( n265164 , n265162 );
and ( n265165 , n265164 , n238409 );
nor ( n265166 , n265163 , n265165 );
not ( n265167 , n265166 );
not ( n265168 , n43810 );
not ( n265169 , n252561 );
or ( n265170 , n265168 , n265169 );
or ( n265171 , n252561 , n43810 );
nand ( n265172 , n265170 , n265171 );
and ( n265173 , n265172 , n255673 );
not ( n265174 , n265172 );
and ( n265175 , n265174 , n255676 );
nor ( n265176 , n265173 , n265175 );
not ( n265177 , n265176 );
nand ( n265178 , n265167 , n265177 );
buf ( n265179 , n238421 );
not ( n265180 , n265179 );
not ( n265181 , n51167 );
or ( n265182 , n265180 , n265181 );
or ( n265183 , n51167 , n265179 );
nand ( n265184 , n265182 , n265183 );
and ( n265185 , n265184 , n51272 );
not ( n265186 , n265184 );
not ( n265187 , n51272 );
and ( n265188 , n265186 , n265187 );
nor ( n265189 , n265185 , n265188 );
not ( n265190 , n265189 );
nand ( n265191 , n265190 , n248981 );
or ( n265192 , n265178 , n265191 );
not ( n265193 , n245241 );
not ( n265194 , n265189 );
nor ( n265195 , n265193 , n265194 );
nand ( n265196 , n265195 , n265178 );
nand ( n265197 , n234823 , n30184 );
nand ( n265198 , n265192 , n265196 , n265197 );
buf ( n265199 , n265198 );
buf ( n265200 , n257909 );
not ( n265201 , n265200 );
not ( n265202 , n250681 );
or ( n265203 , n265201 , n265202 );
or ( n265204 , n250681 , n265200 );
nand ( n265205 , n265203 , n265204 );
not ( n265206 , n265205 );
not ( n265207 , n262220 );
and ( n265208 , n265206 , n265207 );
and ( n265209 , n265205 , n262220 );
nor ( n265210 , n265208 , n265209 );
not ( n265211 , n265210 );
nand ( n265212 , n265211 , n248981 );
not ( n265213 , n233476 );
not ( n265214 , n235008 );
or ( n265215 , n265213 , n265214 );
not ( n265216 , n233476 );
nand ( n265217 , n265216 , n235016 );
nand ( n265218 , n265215 , n265217 );
and ( n265219 , n265218 , n235022 );
not ( n265220 , n265218 );
and ( n265221 , n265220 , n235019 );
nor ( n265222 , n265219 , n265221 );
not ( n265223 , n236017 );
not ( n265224 , n265223 );
not ( n265225 , n260550 );
or ( n265226 , n265224 , n265225 );
or ( n265227 , n260550 , n265223 );
nand ( n265228 , n265226 , n265227 );
not ( n265229 , n265228 );
not ( n265230 , n261269 );
and ( n265231 , n265229 , n265230 );
and ( n265232 , n265228 , n262915 );
nor ( n265233 , n265231 , n265232 );
not ( n265234 , n265233 );
nor ( n265235 , n265222 , n265234 );
or ( n265236 , n265212 , n265235 );
nor ( n265237 , n265211 , n265222 );
nor ( n265238 , n265234 , n258280 );
nand ( n265239 , n265237 , n265238 );
nand ( n265240 , n35431 , n27775 );
nand ( n265241 , n265236 , n265239 , n265240 );
buf ( n265242 , n265241 );
nand ( n265243 , n244513 , n222531 );
not ( n265244 , n259941 );
nand ( n265245 , n265244 , n259931 );
or ( n265246 , n265243 , n265245 );
nor ( n265247 , n244513 , n235050 );
nand ( n265248 , n265247 , n265245 );
nand ( n265249 , n31577 , n31026 );
nand ( n265250 , n265246 , n265248 , n265249 );
buf ( n265251 , n265250 );
not ( n265252 , RI19a97dc0_2627);
or ( n265253 , n25328 , n265252 );
not ( n265254 , RI19a8dd70_2698);
or ( n265255 , n25335 , n265254 );
nand ( n265256 , n265253 , n265255 );
buf ( n265257 , n265256 );
not ( n265258 , RI19abcdc8_2360);
or ( n265259 , n25328 , n265258 );
not ( n265260 , RI19ab3138_2431);
or ( n265261 , n25335 , n265260 );
nand ( n265262 , n265259 , n265261 );
buf ( n265263 , n265262 );
not ( n265264 , n249648 );
not ( n265265 , n265264 );
not ( n265266 , n259590 );
or ( n265267 , n265265 , n265266 );
or ( n265268 , n248385 , n265264 );
nand ( n265269 , n265267 , n265268 );
and ( n265270 , n265269 , n255881 );
not ( n265271 , n265269 );
and ( n265272 , n265271 , n255885 );
nor ( n265273 , n265270 , n265272 );
not ( n265274 , n265273 );
nand ( n265275 , n265274 , n249288 );
buf ( n265276 , n234474 );
not ( n265277 , n265276 );
not ( n265278 , n234121 );
or ( n265279 , n265277 , n265278 );
or ( n265280 , n260807 , n265276 );
nand ( n265281 , n265279 , n265280 );
not ( n265282 , n265281 );
not ( n265283 , n234186 );
and ( n265284 , n265282 , n265283 );
and ( n265285 , n265281 , n248154 );
nor ( n265286 , n265284 , n265285 );
not ( n265287 , n265286 );
not ( n265288 , n258308 );
nand ( n265289 , n265287 , n265288 );
or ( n265290 , n265275 , n265289 );
not ( n265291 , n265287 );
not ( n265292 , n265274 );
or ( n265293 , n265291 , n265292 );
nor ( n265294 , n265288 , n222533 );
nand ( n265295 , n265293 , n265294 );
nand ( n265296 , n31577 , n36845 );
nand ( n265297 , n265290 , n265295 , n265296 );
buf ( n265298 , n265297 );
not ( n265299 , n247924 );
not ( n265300 , n239855 );
or ( n265301 , n265299 , n265300 );
not ( n265302 , n247924 );
nand ( n265303 , n265302 , n239854 );
nand ( n265304 , n265301 , n265303 );
and ( n265305 , n265304 , n239931 );
not ( n265306 , n265304 );
and ( n265307 , n265306 , n239924 );
nor ( n265308 , n265305 , n265307 );
not ( n265309 , n265308 );
not ( n265310 , n249996 );
not ( n265311 , n228527 );
or ( n265312 , n265310 , n265311 );
not ( n265313 , n249996 );
nand ( n265314 , n265313 , n50776 );
nand ( n265315 , n265312 , n265314 );
and ( n265316 , n265315 , n50941 );
not ( n265317 , n265315 );
and ( n265318 , n265317 , n50931 );
nor ( n265319 , n265316 , n265318 );
nand ( n265320 , n265309 , n265319 );
or ( n265321 , n261326 , n265320 );
not ( n265322 , n261299 );
nand ( n265323 , n265322 , n265320 );
nand ( n265324 , n251465 , n40508 );
nand ( n265325 , n265321 , n265323 , n265324 );
buf ( n265326 , n265325 );
not ( n265327 , n39199 );
not ( n265328 , n233501 );
or ( n265329 , n265327 , n265328 );
nand ( n265330 , n258242 , n258237 );
and ( n265331 , n265330 , n251695 );
not ( n265332 , n265330 );
not ( n265333 , n251695 );
and ( n265334 , n265332 , n265333 );
nor ( n265335 , n265331 , n265334 );
or ( n265336 , n265335 , n235732 );
nand ( n265337 , n265329 , n265336 );
buf ( n265338 , n265337 );
buf ( n265339 , n32386 );
buf ( n265340 , n55176 );
not ( n265341 , n265340 );
not ( n265342 , n239390 );
or ( n265343 , n265341 , n265342 );
or ( n265344 , n239390 , n265340 );
nand ( n265345 , n265343 , n265344 );
and ( n265346 , n265345 , n249018 );
not ( n265347 , n265345 );
and ( n265348 , n265347 , n249021 );
nor ( n265349 , n265346 , n265348 );
nand ( n265350 , n265349 , n241459 );
not ( n265351 , n223680 );
not ( n265352 , n249489 );
or ( n265353 , n265351 , n265352 );
not ( n265354 , n223680 );
nand ( n265355 , n265354 , n259332 );
nand ( n265356 , n265353 , n265355 );
and ( n265357 , n265356 , n248000 );
not ( n265358 , n265356 );
and ( n265359 , n265358 , n259339 );
nor ( n265360 , n265357 , n265359 );
not ( n265361 , n265360 );
nand ( n265362 , n265361 , n259299 );
or ( n265363 , n265350 , n265362 );
not ( n265364 , n265361 );
not ( n265365 , n265349 );
or ( n265366 , n265364 , n265365 );
nor ( n265367 , n259299 , n27889 );
nand ( n265368 , n265366 , n265367 );
nand ( n265369 , n238114 , n28387 );
nand ( n265370 , n265363 , n265368 , n265369 );
buf ( n265371 , n265370 );
not ( n265372 , n253629 );
not ( n265373 , n246660 );
or ( n265374 , n265372 , n265373 );
not ( n265375 , n253629 );
nand ( n265376 , n265375 , n246653 );
nand ( n265377 , n265374 , n265376 );
and ( n265378 , n265377 , n259371 );
not ( n265379 , n265377 );
and ( n265380 , n265379 , n262526 );
nor ( n265381 , n265378 , n265380 );
nand ( n265382 , n265381 , n223839 );
not ( n265383 , n250666 );
not ( n265384 , n240941 );
or ( n265385 , n265383 , n265384 );
not ( n265386 , n250666 );
nand ( n265387 , n265386 , n240948 );
nand ( n265388 , n265385 , n265387 );
and ( n265389 , n265388 , n240997 );
not ( n265390 , n265388 );
and ( n265391 , n265390 , n244374 );
nor ( n265392 , n265389 , n265391 );
not ( n265393 , n265392 );
not ( n265394 , n50758 );
not ( n265395 , n237867 );
or ( n265396 , n265394 , n265395 );
not ( n265397 , n50758 );
nand ( n265398 , n265397 , n255503 );
nand ( n265399 , n265396 , n265398 );
and ( n265400 , n265399 , n255515 );
not ( n265401 , n265399 );
buf ( n265402 , n256497 );
and ( n265403 , n265401 , n265402 );
nor ( n265404 , n265400 , n265403 );
nand ( n265405 , n265393 , n265404 );
or ( n265406 , n265382 , n265405 );
not ( n265407 , n265393 );
not ( n265408 , n265381 );
or ( n265409 , n265407 , n265408 );
nor ( n265410 , n265404 , n235050 );
nand ( n265411 , n265409 , n265410 );
nand ( n265412 , n246217 , n30043 );
nand ( n265413 , n265406 , n265411 , n265412 );
buf ( n265414 , n265413 );
not ( n265415 , RI19a99ad0_2614);
or ( n265416 , n25328 , n265415 );
not ( n265417 , RI19ace870_2221);
or ( n265418 , n226822 , n265417 );
nand ( n265419 , n265416 , n265418 );
buf ( n265420 , n265419 );
not ( n265421 , n28438 );
not ( n265422 , n51381 );
or ( n265423 , n265421 , n265422 );
not ( n265424 , n39334 );
not ( n265425 , n246826 );
or ( n265426 , n265424 , n265425 );
not ( n265427 , n39334 );
nand ( n265428 , n265427 , n246835 );
nand ( n265429 , n265426 , n265428 );
and ( n265430 , n265429 , n246883 );
not ( n265431 , n265429 );
and ( n265432 , n265431 , n246892 );
nor ( n265433 , n265430 , n265432 );
not ( n265434 , n265433 );
not ( n265435 , n244412 );
not ( n265436 , n247561 );
or ( n265437 , n265435 , n265436 );
or ( n265438 , n247561 , n244412 );
nand ( n265439 , n265437 , n265438 );
and ( n265440 , n265439 , n255006 );
not ( n265441 , n265439 );
not ( n265442 , n255006 );
and ( n265443 , n265441 , n265442 );
nor ( n265444 , n265440 , n265443 );
nand ( n265445 , n265434 , n265444 );
not ( n265446 , n265445 );
not ( n265447 , n33378 );
not ( n265448 , n244203 );
not ( n265449 , n265448 );
or ( n265450 , n265447 , n265449 );
or ( n265451 , n244207 , n33378 );
nand ( n265452 , n265450 , n265451 );
and ( n265453 , n265452 , n233968 );
not ( n265454 , n265452 );
and ( n265455 , n265454 , n233960 );
nor ( n265456 , n265453 , n265455 );
not ( n265457 , n265456 );
not ( n265458 , n265457 );
and ( n265459 , n265446 , n265458 );
and ( n265460 , n265445 , n265457 );
nor ( n265461 , n265459 , n265460 );
or ( n265462 , n265461 , n256376 );
nand ( n265463 , n265423 , n265462 );
buf ( n265464 , n265463 );
buf ( n265465 , n34084 );
buf ( n265466 , n205345 );
nor ( n265467 , n254177 , n234440 );
not ( n265468 , n254694 );
not ( n265469 , n265468 );
not ( n265470 , n249610 );
or ( n265471 , n265469 , n265470 );
or ( n265472 , n249610 , n265468 );
nand ( n265473 , n265471 , n265472 );
and ( n265474 , n265473 , n250234 );
not ( n265475 , n265473 );
not ( n265476 , n250234 );
and ( n265477 , n265475 , n265476 );
nor ( n265478 , n265474 , n265477 );
nor ( n265479 , n254162 , n265478 );
nand ( n265480 , n265467 , n265479 );
not ( n265481 , n265478 );
not ( n265482 , n265481 );
not ( n265483 , n254149 );
or ( n265484 , n265482 , n265483 );
nor ( n265485 , n254163 , n251361 );
nand ( n265486 , n265484 , n265485 );
nand ( n265487 , n31577 , n32107 );
nand ( n265488 , n265480 , n265486 , n265487 );
buf ( n265489 , n265488 );
not ( n265490 , n252627 );
not ( n265491 , n265490 );
not ( n265492 , n253264 );
or ( n265493 , n265491 , n265492 );
not ( n265494 , n265490 );
nand ( n265495 , n265494 , n253271 );
nand ( n265496 , n265493 , n265495 );
and ( n265497 , n265496 , n232899 );
not ( n265498 , n265496 );
and ( n265499 , n265498 , n232900 );
nor ( n265500 , n265497 , n265499 );
nand ( n265501 , n265500 , n245241 );
not ( n265502 , n246810 );
not ( n265503 , n249927 );
or ( n265504 , n265502 , n265503 );
not ( n265505 , n246810 );
nand ( n265506 , n265505 , n255493 );
nand ( n265507 , n265504 , n265506 );
xnor ( n265508 , n265507 , n255500 );
not ( n265509 , n48975 );
not ( n265510 , n254603 );
or ( n265511 , n265509 , n265510 );
not ( n265512 , n48975 );
nand ( n265513 , n265512 , n254594 );
nand ( n265514 , n265511 , n265513 );
and ( n265515 , n265514 , n264627 );
not ( n265516 , n265514 );
and ( n265517 , n265516 , n254611 );
nor ( n265518 , n265515 , n265517 );
not ( n265519 , n265518 );
nand ( n265520 , n265508 , n265519 );
or ( n265521 , n265501 , n265520 );
not ( n265522 , n265519 );
not ( n265523 , n265500 );
or ( n265524 , n265522 , n265523 );
nor ( n265525 , n265508 , n37725 );
nand ( n265526 , n265524 , n265525 );
nand ( n265527 , n35431 , n27808 );
nand ( n265528 , n265521 , n265526 , n265527 );
buf ( n265529 , n265528 );
not ( n265530 , n44924 );
not ( n265531 , n257764 );
or ( n265532 , n265530 , n265531 );
not ( n265533 , n247839 );
not ( n265534 , n265533 );
not ( n265535 , n54537 );
or ( n265536 , n265534 , n265535 );
not ( n265537 , n265533 );
nand ( n265538 , n265537 , n246188 );
nand ( n265539 , n265536 , n265538 );
and ( n265540 , n265539 , n246193 );
not ( n265541 , n265539 );
and ( n265542 , n265541 , n246196 );
nor ( n265543 , n265540 , n265542 );
not ( n265544 , n254943 );
nand ( n265545 , n265543 , n265544 );
not ( n265546 , n254978 );
and ( n265547 , n265545 , n265546 );
not ( n265548 , n265545 );
and ( n265549 , n265548 , n254978 );
nor ( n265550 , n265547 , n265549 );
or ( n265551 , n265550 , n49959 );
nand ( n265552 , n265532 , n265551 );
buf ( n265553 , n265552 );
not ( n265554 , n40451 );
not ( n265555 , n235878 );
or ( n265556 , n265554 , n265555 );
not ( n265557 , n40451 );
nand ( n265558 , n265557 , n235887 );
nand ( n265559 , n265556 , n265558 );
and ( n265560 , n265559 , n259858 );
not ( n265561 , n265559 );
and ( n265562 , n265561 , n259855 );
nor ( n265563 , n265560 , n265562 );
not ( n265564 , n265563 );
nand ( n265565 , n265564 , n262758 );
buf ( n265566 , n45678 );
not ( n265567 , n265566 );
not ( n265568 , n248210 );
or ( n265569 , n265567 , n265568 );
or ( n265570 , n248210 , n265566 );
nand ( n265571 , n265569 , n265570 );
and ( n265572 , n265571 , n261431 );
not ( n265573 , n265571 );
and ( n265574 , n265573 , n261434 );
nor ( n265575 , n265572 , n265574 );
not ( n265576 , n265575 );
nand ( n265577 , n265576 , n226010 );
or ( n265578 , n265565 , n265577 );
nor ( n265579 , n265576 , n234440 );
nand ( n265580 , n265565 , n265579 );
nand ( n265581 , n238114 , n28211 );
nand ( n265582 , n265578 , n265580 , n265581 );
buf ( n265583 , n265582 );
nand ( n265584 , n249096 , n222532 );
not ( n265585 , n238751 );
not ( n265586 , n247991 );
or ( n265587 , n265585 , n265586 );
not ( n265588 , n238751 );
nand ( n265589 , n265588 , n247999 );
nand ( n265590 , n265587 , n265589 );
and ( n265591 , n265590 , n261862 );
not ( n265592 , n265590 );
and ( n265593 , n265592 , n261859 );
nor ( n265594 , n265591 , n265593 );
nand ( n265595 , n258043 , n265594 );
or ( n265596 , n265584 , n265595 );
not ( n265597 , n258043 );
not ( n265598 , n249096 );
or ( n265599 , n265597 , n265598 );
nor ( n265600 , n265594 , n234440 );
nand ( n265601 , n265599 , n265600 );
nand ( n265602 , n261585 , n35336 );
nand ( n265603 , n265596 , n265601 , n265602 );
buf ( n265604 , n265603 );
nor ( n265605 , n261798 , n31563 );
nand ( n265606 , n27880 , n205649 );
or ( n265607 , n265605 , n265606 );
nand ( n265608 , n265605 , n205651 );
nand ( n265609 , n35431 , n204594 );
nand ( n265610 , n265607 , n265608 , n265609 );
buf ( n265611 , n265610 );
or ( n265612 , n226819 , n262547 );
not ( n265613 , RI19abb748_2371);
or ( n265614 , n226822 , n265613 );
nand ( n265615 , n265612 , n265614 );
buf ( n265616 , n265615 );
not ( n265617 , n26216 );
not ( n265618 , n244073 );
or ( n265619 , n265617 , n265618 );
not ( n265620 , n252802 );
not ( n265621 , n50930 );
or ( n265622 , n265620 , n265621 );
or ( n265623 , n50930 , n252802 );
nand ( n265624 , n265622 , n265623 );
and ( n265625 , n265624 , n244532 );
not ( n265626 , n265624 );
and ( n265627 , n265626 , n244529 );
nor ( n265628 , n265625 , n265627 );
not ( n265629 , n265628 );
not ( n265630 , n265629 );
not ( n265631 , n223310 );
not ( n265632 , n265631 );
not ( n265633 , n248210 );
or ( n265634 , n265632 , n265633 );
not ( n265635 , n265631 );
nand ( n265636 , n265635 , n248219 );
nand ( n265637 , n265634 , n265636 );
and ( n265638 , n265637 , n261431 );
not ( n265639 , n265637 );
and ( n265640 , n265639 , n261434 );
nor ( n265641 , n265638 , n265640 );
not ( n265642 , n31438 );
not ( n265643 , n247013 );
or ( n265644 , n265642 , n265643 );
or ( n265645 , n247013 , n31438 );
nand ( n265646 , n265644 , n265645 );
not ( n265647 , n265646 );
not ( n265648 , n250113 );
and ( n265649 , n265647 , n265648 );
and ( n265650 , n265646 , n250123 );
nor ( n265651 , n265649 , n265650 );
nand ( n265652 , n265641 , n265651 );
not ( n265653 , n265652 );
and ( n265654 , n265630 , n265653 );
and ( n265655 , n265629 , n265652 );
nor ( n265656 , n265654 , n265655 );
or ( n265657 , n265656 , n259651 );
nand ( n265658 , n265619 , n265657 );
buf ( n265659 , n265658 );
nor ( n265660 , n264311 , n253544 );
not ( n265661 , n242289 );
not ( n265662 , n257963 );
or ( n265663 , n265661 , n265662 );
or ( n265664 , n39598 , n242289 );
nand ( n265665 , n265663 , n265664 );
xnor ( n265666 , n265665 , n39755 );
nor ( n265667 , n265666 , n264324 );
nand ( n265668 , n265660 , n265667 );
not ( n265669 , n265666 );
not ( n265670 , n265669 );
not ( n265671 , n264312 );
or ( n265672 , n265670 , n265671 );
nor ( n265673 , n264325 , n235050 );
nand ( n265674 , n265672 , n265673 );
nand ( n265675 , n247744 , n35568 );
nand ( n265676 , n265668 , n265674 , n265675 );
buf ( n265677 , n265676 );
not ( n265678 , RI19ac6080_2284);
or ( n265679 , n25328 , n265678 );
or ( n265680 , n25335 , n260178 );
nand ( n265681 , n265679 , n265680 );
buf ( n265682 , n265681 );
not ( n265683 , n259597 );
nand ( n265684 , n265683 , n239934 );
not ( n265685 , n242223 );
not ( n265686 , n249298 );
or ( n265687 , n265685 , n265686 );
not ( n265688 , n242223 );
nand ( n265689 , n265688 , n53140 );
nand ( n265690 , n265687 , n265689 );
and ( n265691 , n265690 , n249366 );
not ( n265692 , n265690 );
and ( n265693 , n265692 , n249363 );
nor ( n265694 , n265691 , n265693 );
nand ( n265695 , n265694 , n259608 );
or ( n265696 , n265684 , n265695 );
not ( n265697 , n259608 );
not ( n265698 , n265683 );
or ( n265699 , n265697 , n265698 );
buf ( n265700 , n236795 );
nor ( n265701 , n265694 , n265700 );
nand ( n265702 , n265699 , n265701 );
nand ( n265703 , n31576 , n27931 );
nand ( n265704 , n265696 , n265702 , n265703 );
buf ( n265705 , n265704 );
not ( n265706 , n243634 );
not ( n265707 , n245701 );
or ( n265708 , n265706 , n265707 );
not ( n265709 , n246639 );
not ( n265710 , n265709 );
not ( n265711 , n255455 );
or ( n265712 , n265710 , n265711 );
not ( n265713 , n265709 );
nand ( n265714 , n265713 , n255464 );
nand ( n265715 , n265712 , n265714 );
and ( n265716 , n265715 , n259459 );
not ( n265717 , n265715 );
and ( n265718 , n265717 , n259463 );
nor ( n265719 , n265716 , n265718 );
not ( n265720 , n265719 );
not ( n265721 , n261039 );
nand ( n265722 , n265720 , n265721 );
not ( n265723 , n261049 );
and ( n265724 , n265722 , n265723 );
not ( n265725 , n265722 );
and ( n265726 , n265725 , n261049 );
nor ( n265727 , n265724 , n265726 );
or ( n265728 , n265727 , n244217 );
nand ( n265729 , n265708 , n265728 );
buf ( n265730 , n265729 );
buf ( n265731 , n234780 );
not ( n265732 , n265731 );
not ( n265733 , n261834 );
or ( n265734 , n265732 , n265733 );
or ( n265735 , n242675 , n265731 );
nand ( n265736 , n265734 , n265735 );
and ( n265737 , n265736 , n242683 );
not ( n265738 , n265736 );
and ( n265739 , n265738 , n242680 );
nor ( n265740 , n265737 , n265739 );
nand ( n265741 , n265740 , n222532 );
not ( n265742 , n248745 );
not ( n265743 , n55725 );
or ( n265744 , n265742 , n265743 );
not ( n265745 , n248745 );
not ( n265746 , n55725 );
nand ( n265747 , n265745 , n265746 );
nand ( n265748 , n265744 , n265747 );
and ( n265749 , n265748 , n264675 );
not ( n265750 , n265748 );
and ( n265751 , n265750 , n264672 );
nor ( n265752 , n265749 , n265751 );
nor ( n265753 , n265752 , n257395 );
or ( n265754 , n265741 , n265753 );
nor ( n265755 , n265740 , n31572 );
nand ( n265756 , n265755 , n265753 );
nand ( n265757 , n49054 , n41265 );
nand ( n265758 , n265754 , n265756 , n265757 );
buf ( n265759 , n265758 );
not ( n265760 , n246385 );
not ( n265761 , n239003 );
not ( n265762 , n52221 );
or ( n265763 , n265761 , n265762 );
nand ( n265764 , n52229 , n239004 );
nand ( n265765 , n265763 , n265764 );
not ( n265766 , n265765 );
or ( n265767 , n265760 , n265766 );
or ( n265768 , n265765 , n259264 );
nand ( n265769 , n265767 , n265768 );
not ( n265770 , n265769 );
nor ( n265771 , n265770 , n244399 );
not ( n265772 , n265771 );
not ( n265773 , n258482 );
not ( n265774 , n259150 );
not ( n265775 , n265774 );
or ( n265776 , n265773 , n265775 );
not ( n265777 , n258482 );
nand ( n265778 , n265777 , n259150 );
nand ( n265779 , n265776 , n265778 );
and ( n265780 , n265779 , n250942 );
not ( n265781 , n265779 );
and ( n265782 , n265781 , n259153 );
nor ( n265783 , n265780 , n265782 );
not ( n265784 , n254585 );
not ( n265785 , n249462 );
or ( n265786 , n265784 , n265785 );
not ( n265787 , n254585 );
nand ( n265788 , n265787 , n249469 );
nand ( n265789 , n265786 , n265788 );
and ( n265790 , n265789 , n259701 );
not ( n265791 , n265789 );
and ( n265792 , n265791 , n259704 );
nor ( n265793 , n265790 , n265792 );
not ( n265794 , n265793 );
nand ( n265795 , n265783 , n265794 );
or ( n265796 , n265772 , n265795 );
not ( n265797 , n265783 );
not ( n265798 , n265769 );
or ( n265799 , n265797 , n265798 );
nor ( n265800 , n265794 , n31572 );
nand ( n265801 , n265799 , n265800 );
nand ( n265802 , n31576 , n32946 );
nand ( n265803 , n265796 , n265801 , n265802 );
buf ( n265804 , n265803 );
not ( n265805 , n252580 );
not ( n265806 , n252564 );
not ( n265807 , n265806 );
or ( n265808 , n265805 , n265807 );
not ( n265809 , n241160 );
not ( n265810 , n235728 );
or ( n265811 , n265809 , n265810 );
not ( n265812 , n241160 );
nand ( n265813 , n265812 , n235718 );
nand ( n265814 , n265811 , n265813 );
and ( n265815 , n265814 , n260711 );
not ( n265816 , n265814 );
and ( n265817 , n265816 , n236504 );
nor ( n265818 , n265815 , n265817 );
not ( n265819 , n265818 );
nor ( n265820 , n265819 , n244399 );
nand ( n265821 , n265808 , n265820 );
nand ( n265822 , n265806 , n252577 , n265819 );
nand ( n265823 , n238114 , n42936 );
nand ( n265824 , n265821 , n265822 , n265823 );
buf ( n265825 , n265824 );
not ( n265826 , n241141 );
not ( n265827 , n235728 );
or ( n265828 , n265826 , n265827 );
not ( n265829 , n241141 );
nand ( n265830 , n265829 , n235718 );
nand ( n265831 , n265828 , n265830 );
and ( n265832 , n265831 , n260711 );
not ( n265833 , n265831 );
and ( n265834 , n265833 , n260712 );
nor ( n265835 , n265832 , n265834 );
nor ( n265836 , n265835 , n55152 );
buf ( n265837 , n54076 );
not ( n265838 , n265837 );
not ( n265839 , n242315 );
or ( n265840 , n265838 , n265839 );
or ( n265841 , n260248 , n265837 );
nand ( n265842 , n265840 , n265841 );
and ( n265843 , n265842 , n242381 );
not ( n265844 , n265842 );
and ( n265845 , n265844 , n242374 );
nor ( n265846 , n265843 , n265845 );
not ( n265847 , n265846 );
not ( n265848 , n248124 );
not ( n265849 , n265848 );
not ( n265850 , n256901 );
or ( n265851 , n265849 , n265850 );
not ( n265852 , n265848 );
nand ( n265853 , n265852 , n255593 );
nand ( n265854 , n265851 , n265853 );
and ( n265855 , n265854 , n255599 );
not ( n265856 , n265854 );
and ( n265857 , n265856 , n255596 );
nor ( n265858 , n265855 , n265857 );
not ( n265859 , n265858 );
nor ( n265860 , n265847 , n265859 );
nand ( n265861 , n265836 , n265860 );
not ( n265862 , n265858 );
not ( n265863 , n265835 );
not ( n265864 , n265863 );
or ( n265865 , n265862 , n265864 );
nor ( n265866 , n265846 , n235895 );
nand ( n265867 , n265865 , n265866 );
nand ( n265868 , n51381 , n30426 );
nand ( n265869 , n265861 , n265867 , n265868 );
buf ( n265870 , n265869 );
not ( n265871 , n204717 );
not ( n265872 , n245702 );
or ( n265873 , n265871 , n265872 );
not ( n265874 , n263021 );
nand ( n265875 , n265874 , n263011 );
not ( n265876 , n242251 );
not ( n265877 , n249298 );
or ( n265878 , n265876 , n265877 );
not ( n265879 , n242251 );
nand ( n265880 , n265879 , n53140 );
nand ( n265881 , n265878 , n265880 );
and ( n265882 , n265881 , n249366 );
not ( n265883 , n265881 );
and ( n265884 , n265883 , n249363 );
nor ( n265885 , n265882 , n265884 );
not ( n265886 , n265885 );
and ( n265887 , n265875 , n265886 );
not ( n265888 , n265875 );
and ( n265889 , n265888 , n265885 );
nor ( n265890 , n265887 , n265889 );
or ( n265891 , n265890 , n253544 );
nand ( n265892 , n265873 , n265891 );
buf ( n265893 , n265892 );
not ( n265894 , n236394 );
nand ( n265895 , n265894 , n236508 );
not ( n265896 , n252595 );
not ( n265897 , n253271 );
or ( n265898 , n265896 , n265897 );
or ( n265899 , n253271 , n252595 );
nand ( n265900 , n265898 , n265899 );
and ( n265901 , n265900 , n55135 );
not ( n265902 , n265900 );
and ( n265903 , n265902 , n253348 );
nor ( n265904 , n265901 , n265903 );
not ( n265905 , n265904 );
nand ( n265906 , n265895 , n265905 , n33255 );
nor ( n265907 , n236394 , n234021 );
nand ( n265908 , n265904 , n236508 , n265907 );
nand ( n265909 , n50615 , n31333 );
nand ( n265910 , n265906 , n265908 , n265909 );
buf ( n265911 , n265910 );
not ( n265912 , RI19ac5720_2288);
or ( n265913 , n25328 , n265912 );
or ( n265914 , n25336 , n265258 );
nand ( n265915 , n265913 , n265914 );
buf ( n265916 , n265915 );
nand ( n265917 , n261918 , n261922 );
or ( n265918 , n265917 , n254923 );
nand ( n265919 , n265917 , n257077 );
nand ( n265920 , n241378 , n208320 );
nand ( n265921 , n265918 , n265919 , n265920 );
buf ( n265922 , n265921 );
buf ( n265923 , n39464 );
buf ( n265924 , n40888 );
not ( n265925 , n204312 );
not ( n265926 , n41945 );
or ( n265927 , n265925 , n265926 );
not ( n265928 , n243284 );
buf ( n265929 , n249655 );
not ( n265930 , n265929 );
not ( n265931 , n259590 );
or ( n265932 , n265930 , n265931 );
or ( n265933 , n259590 , n265929 );
nand ( n265934 , n265932 , n265933 );
and ( n265935 , n265934 , n259595 );
not ( n265936 , n265934 );
and ( n265937 , n265936 , n255880 );
nor ( n265938 , n265935 , n265937 );
nand ( n265939 , n265928 , n265938 );
and ( n265940 , n265939 , n257771 );
not ( n265941 , n265939 );
and ( n265942 , n265941 , n243417 );
nor ( n265943 , n265940 , n265942 );
or ( n265944 , n265943 , n264469 );
nand ( n265945 , n265927 , n265944 );
buf ( n265946 , n265945 );
not ( n265947 , n28883 );
not ( n265948 , n51381 );
or ( n265949 , n265947 , n265948 );
nand ( n265950 , n265360 , n259299 );
not ( n265951 , n265950 );
not ( n265952 , n259310 );
not ( n265953 , n265952 );
and ( n265954 , n265951 , n265953 );
and ( n265955 , n265950 , n265952 );
nor ( n265956 , n265954 , n265955 );
or ( n265957 , n265956 , n251498 );
nand ( n265958 , n265949 , n265957 );
buf ( n265959 , n265958 );
not ( n265960 , n32790 );
not ( n265961 , n53257 );
or ( n265962 , n265960 , n265961 );
or ( n265963 , n53257 , n32790 );
nand ( n265964 , n265962 , n265963 );
and ( n265965 , n265964 , n53451 );
not ( n265966 , n265964 );
and ( n265967 , n265966 , n53454 );
nor ( n265968 , n265965 , n265967 );
nor ( n265969 , n265968 , n39763 );
not ( n265970 , n265969 );
not ( n265971 , n36720 );
not ( n265972 , n253863 );
or ( n265973 , n265971 , n265972 );
not ( n265974 , n36720 );
nand ( n265975 , n265974 , n253855 );
nand ( n265976 , n265973 , n265975 );
and ( n265977 , n265976 , n239854 );
not ( n265978 , n265976 );
and ( n265979 , n265978 , n258013 );
nor ( n265980 , n265977 , n265979 );
not ( n265981 , n251664 );
not ( n265982 , n265981 );
not ( n265983 , n46941 );
or ( n265984 , n265982 , n265983 );
not ( n265985 , n265981 );
nand ( n265986 , n265985 , n46950 );
nand ( n265987 , n265984 , n265986 );
and ( n265988 , n265987 , n47157 );
not ( n265989 , n265987 );
and ( n265990 , n265989 , n224925 );
nor ( n265991 , n265988 , n265990 );
not ( n265992 , n265991 );
nand ( n265993 , n265980 , n265992 );
or ( n265994 , n265970 , n265993 );
not ( n265995 , n265980 );
not ( n265996 , n265968 );
not ( n265997 , n265996 );
or ( n265998 , n265995 , n265997 );
nand ( n265999 , n265991 , n205649 );
not ( n266000 , n265999 );
nand ( n266001 , n265998 , n266000 );
nand ( n266002 , n237714 , n32378 );
nand ( n266003 , n265994 , n266001 , n266002 );
buf ( n266004 , n266003 );
buf ( n266005 , n32344 );
not ( n266006 , n252278 );
not ( n266007 , n243953 );
or ( n266008 , n266006 , n266007 );
or ( n266009 , n243953 , n252278 );
nand ( n266010 , n266008 , n266009 );
and ( n266011 , n266010 , n250272 );
not ( n266012 , n266010 );
and ( n266013 , n266012 , n250275 );
nor ( n266014 , n266011 , n266013 );
not ( n266015 , n266014 );
nor ( n266016 , n266015 , n235050 );
not ( n266017 , n266016 );
not ( n266018 , n255104 );
not ( n266019 , n228364 );
and ( n266020 , n204535 , n50594 );
not ( n266021 , n204535 );
and ( n266022 , n266021 , n50595 );
nor ( n266023 , n266020 , n266022 );
not ( n266024 , n266023 );
not ( n266025 , n266024 );
or ( n266026 , n266019 , n266025 );
nand ( n266027 , n266023 , n50539 );
nand ( n266028 , n266026 , n266027 );
not ( n266029 , n266028 );
nand ( n266030 , n266018 , n266029 );
or ( n266031 , n266017 , n266030 );
nor ( n266032 , n266014 , n258280 );
nand ( n266033 , n266032 , n266030 );
nand ( n266034 , n252711 , n204468 );
nand ( n266035 , n266031 , n266033 , n266034 );
buf ( n266036 , n266035 );
buf ( n266037 , n240635 );
not ( n266038 , n226164 );
not ( n266039 , n245680 );
or ( n266040 , n266038 , n266039 );
or ( n266041 , n245680 , n226164 );
nand ( n266042 , n266040 , n266041 );
and ( n266043 , n266042 , n258937 );
not ( n266044 , n266042 );
and ( n266045 , n266044 , n254974 );
nor ( n266046 , n266043 , n266045 );
not ( n266047 , n266046 );
nor ( n266048 , n266047 , n55108 );
not ( n266049 , n266048 );
not ( n266050 , n237383 );
nand ( n266051 , n266050 , n237706 );
or ( n266052 , n266049 , n266051 );
not ( n266053 , n266050 );
not ( n266054 , n266046 );
or ( n266055 , n266053 , n266054 );
nor ( n266056 , n237706 , n221279 );
nand ( n266057 , n266055 , n266056 );
nand ( n266058 , n246217 , n34776 );
nand ( n266059 , n266052 , n266057 , n266058 );
buf ( n266060 , n266059 );
not ( n266061 , n40156 );
not ( n266062 , n234453 );
or ( n266063 , n266061 , n266062 );
nand ( n266064 , n260344 , n260352 );
and ( n266065 , n266064 , n258627 );
not ( n266066 , n266064 );
and ( n266067 , n266066 , n258562 );
nor ( n266068 , n266065 , n266067 );
or ( n266069 , n266068 , n52445 );
nand ( n266070 , n266063 , n266069 );
buf ( n266071 , n266070 );
buf ( n266072 , RI175379b8_594);
and ( n266073 , n27883 , n266072 );
buf ( n266074 , n266073 );
not ( n266075 , n31110 );
not ( n266076 , n255116 );
or ( n266077 , n266075 , n266076 );
not ( n266078 , n226606 );
not ( n266079 , n44315 );
or ( n266080 , n266078 , n266079 );
not ( n266081 , n226606 );
nand ( n266082 , n266081 , n44324 );
nand ( n266083 , n266080 , n266082 );
not ( n266084 , n256460 );
and ( n266085 , n266083 , n266084 );
not ( n266086 , n266083 );
and ( n266087 , n266086 , n256460 );
nor ( n266088 , n266085 , n266087 );
not ( n266089 , n266088 );
not ( n266090 , n48222 );
not ( n266091 , n266090 );
not ( n266092 , n226557 );
or ( n266093 , n266091 , n266092 );
not ( n266094 , n266090 );
nand ( n266095 , n266094 , n48804 );
nand ( n266096 , n266093 , n266095 );
and ( n266097 , n266096 , n260471 );
not ( n266098 , n266096 );
not ( n266099 , n259385 );
and ( n266100 , n266098 , n266099 );
nor ( n266101 , n266097 , n266100 );
nand ( n266102 , n266089 , n266101 );
not ( n266103 , n250778 );
not ( n266104 , n251154 );
or ( n266105 , n266103 , n266104 );
not ( n266106 , n250778 );
nand ( n266107 , n266106 , n251253 );
nand ( n266108 , n266105 , n266107 );
and ( n266109 , n266108 , n251299 );
not ( n266110 , n266108 );
and ( n266111 , n266110 , n251314 );
nor ( n266112 , n266109 , n266111 );
not ( n266113 , n266112 );
and ( n266114 , n266102 , n266113 );
not ( n266115 , n266102 );
and ( n266116 , n266115 , n266112 );
nor ( n266117 , n266114 , n266116 );
or ( n266118 , n266117 , n251498 );
nand ( n266119 , n266077 , n266118 );
buf ( n266120 , n266119 );
nor ( n266121 , n264387 , n49959 );
not ( n266122 , n257262 );
nand ( n266123 , n266121 , n266122 , n257273 );
not ( n266124 , n264387 );
not ( n266125 , n266124 );
not ( n266126 , n266122 );
or ( n266127 , n266125 , n266126 );
nor ( n266128 , n257273 , n237384 );
nand ( n266129 , n266127 , n266128 );
nand ( n266130 , n31577 , n39485 );
nand ( n266131 , n266123 , n266129 , n266130 );
buf ( n266132 , n266131 );
nand ( n266133 , n251893 , n253565 );
not ( n266134 , n259706 );
nand ( n266135 , n266134 , n259693 );
or ( n266136 , n266133 , n266135 );
not ( n266137 , n259693 );
not ( n266138 , n251893 );
or ( n266139 , n266137 , n266138 );
nor ( n266140 , n266134 , n39763 );
nand ( n266141 , n266139 , n266140 );
nand ( n266142 , n31577 , n35557 );
nand ( n266143 , n266136 , n266141 , n266142 );
buf ( n266144 , n266143 );
buf ( n266145 , n33697 );
not ( n266146 , n266145 );
not ( n266147 , n233904 );
or ( n266148 , n266146 , n266147 );
not ( n266149 , n244203 );
or ( n266150 , n266149 , n266145 );
nand ( n266151 , n266148 , n266150 );
not ( n266152 , n266151 );
not ( n266153 , n233968 );
and ( n266154 , n266152 , n266153 );
and ( n266155 , n266151 , n233968 );
nor ( n266156 , n266154 , n266155 );
nand ( n266157 , n266156 , n40466 );
not ( n266158 , n263222 );
buf ( n266159 , n242951 );
not ( n266160 , n266159 );
not ( n266161 , n245929 );
or ( n266162 , n266160 , n266161 );
or ( n266163 , n245929 , n266159 );
nand ( n266164 , n266162 , n266163 );
not ( n266165 , n256191 );
and ( n266166 , n266164 , n266165 );
not ( n266167 , n266164 );
buf ( n266168 , n256190 );
not ( n266169 , n266168 );
and ( n266170 , n266167 , n266169 );
nor ( n266171 , n266166 , n266170 );
not ( n266172 , n266171 );
nand ( n266173 , n266158 , n266172 );
or ( n266174 , n266157 , n266173 );
nor ( n266175 , n266156 , n260567 );
nand ( n266176 , n266175 , n266173 );
nand ( n266177 , n247585 , n33346 );
nand ( n266178 , n266174 , n266176 , n266177 );
buf ( n266179 , n266178 );
buf ( n266180 , n253237 );
not ( n266181 , n266180 );
not ( n266182 , n240684 );
or ( n266183 , n266181 , n266182 );
or ( n266184 , n240684 , n266180 );
nand ( n266185 , n266183 , n266184 );
and ( n266186 , n266185 , n240801 );
not ( n266187 , n266185 );
and ( n266188 , n266187 , n240811 );
nor ( n266189 , n266186 , n266188 );
nand ( n266190 , n266189 , n246177 );
not ( n266191 , n251072 );
not ( n266192 , n50474 );
or ( n266193 , n266191 , n266192 );
not ( n266194 , n251072 );
nand ( n266195 , n266194 , n50482 );
nand ( n266196 , n266193 , n266195 );
and ( n266197 , n266196 , n263851 );
not ( n266198 , n266196 );
and ( n266199 , n266198 , n263848 );
nor ( n266200 , n266197 , n266199 );
not ( n266201 , n266200 );
nand ( n266202 , n259083 , n266201 );
or ( n266203 , n266190 , n266202 );
not ( n266204 , n266189 );
not ( n266205 , n259083 );
or ( n266206 , n266204 , n266205 );
nor ( n266207 , n266201 , n244216 );
nand ( n266208 , n266206 , n266207 );
nand ( n266209 , n247744 , n30133 );
nand ( n266210 , n266203 , n266208 , n266209 );
buf ( n266211 , n266210 );
not ( n266212 , RI19abcbe8_2361);
or ( n266213 , n25328 , n266212 );
not ( n266214 , RI19ab2f58_2432);
or ( n266215 , n25335 , n266214 );
nand ( n266216 , n266213 , n266215 );
buf ( n266217 , n266216 );
not ( n266218 , n33537 );
not ( n266219 , n241068 );
or ( n266220 , n266218 , n266219 );
not ( n266221 , n234467 );
not ( n266222 , n234125 );
or ( n266223 , n266221 , n266222 );
not ( n266224 , n234467 );
nand ( n266225 , n266224 , n234124 );
nand ( n266226 , n266223 , n266225 );
and ( n266227 , n266226 , n234184 );
not ( n266228 , n266226 );
and ( n266229 , n266228 , n234186 );
nor ( n266230 , n266227 , n266229 );
not ( n266231 , n266230 );
nand ( n266232 , n260473 , n266231 );
and ( n266233 , n266232 , n259021 );
not ( n266234 , n266232 );
and ( n266235 , n266234 , n259020 );
nor ( n266236 , n266233 , n266235 );
or ( n266237 , n266236 , n261009 );
nand ( n266238 , n266220 , n266237 );
buf ( n266239 , n266238 );
not ( n266240 , RI19aceac8_2220);
or ( n266241 , n25328 , n266240 );
not ( n266242 , RI19ac5e28_2285);
or ( n266243 , n25336 , n266242 );
nand ( n266244 , n266241 , n266243 );
buf ( n266245 , n266244 );
not ( n266246 , n235976 );
not ( n266247 , n260550 );
or ( n266248 , n266246 , n266247 );
not ( n266249 , n235976 );
nand ( n266250 , n266249 , n260557 );
nand ( n266251 , n266248 , n266250 );
and ( n266252 , n266251 , n262915 );
not ( n266253 , n266251 );
not ( n266254 , n261269 );
and ( n266255 , n266253 , n266254 );
nor ( n266256 , n266252 , n266255 );
nand ( n266257 , n255467 , n266256 );
not ( n266258 , n262230 );
or ( n266259 , n266257 , n266258 );
not ( n266260 , n255401 );
not ( n266261 , n255467 );
or ( n266262 , n266260 , n266261 );
nor ( n266263 , n266256 , n235895 );
nand ( n266264 , n266262 , n266263 );
nand ( n266265 , n244987 , n32252 );
nand ( n266266 , n266259 , n266264 , n266265 );
buf ( n266267 , n266266 );
not ( n266268 , n241962 );
not ( n266269 , n245490 );
not ( n266270 , n241892 );
or ( n266271 , n266269 , n266270 );
not ( n266272 , n245490 );
nand ( n266273 , n241893 , n266272 );
nand ( n266274 , n266271 , n266273 );
not ( n266275 , n266274 );
and ( n266276 , n266268 , n266275 );
and ( n266277 , n241962 , n266274 );
nor ( n266278 , n266276 , n266277 );
not ( n266279 , n266278 );
not ( n266280 , n266279 );
and ( n266281 , n246503 , n236503 );
not ( n266282 , n246503 );
and ( n266283 , n266282 , n255408 );
nor ( n266284 , n266281 , n266283 );
and ( n266285 , n266284 , n255455 );
not ( n266286 , n266284 );
and ( n266287 , n266286 , n255465 );
nor ( n266288 , n266285 , n266287 );
not ( n266289 , n266288 );
not ( n266290 , n266289 );
or ( n266291 , n266280 , n266290 );
not ( n266292 , n260000 );
nor ( n266293 , n266292 , n49959 );
nand ( n266294 , n266291 , n266293 );
nor ( n266295 , n266278 , n234445 );
not ( n266296 , n266288 );
nand ( n266297 , n266295 , n266292 , n266296 );
nand ( n266298 , n50615 , n32356 );
nand ( n266299 , n266294 , n266297 , n266298 );
buf ( n266300 , n266299 );
not ( n266301 , n244160 );
not ( n266302 , n234810 );
or ( n266303 , n266301 , n266302 );
not ( n266304 , n244160 );
nand ( n266305 , n266304 , n234803 );
nand ( n266306 , n266303 , n266305 );
and ( n266307 , n266306 , n250395 );
not ( n266308 , n266306 );
and ( n266309 , n266308 , n250398 );
nor ( n266310 , n266307 , n266309 );
nor ( n266311 , n266310 , n219702 );
not ( n266312 , n266311 );
not ( n266313 , n239089 );
not ( n266314 , n52221 );
or ( n266315 , n266313 , n266314 );
not ( n266316 , n239089 );
nand ( n266317 , n266316 , n52229 );
nand ( n266318 , n266315 , n266317 );
and ( n266319 , n266318 , n259264 );
not ( n266320 , n266318 );
and ( n266321 , n266320 , n264700 );
nor ( n266322 , n266319 , n266321 );
not ( n266323 , n266322 );
not ( n266324 , n48651 );
not ( n266325 , n234420 );
or ( n266326 , n266324 , n266325 );
not ( n266327 , n48651 );
nand ( n266328 , n266327 , n239119 );
nand ( n266329 , n266326 , n266328 );
and ( n266330 , n266329 , n239221 );
not ( n266331 , n266329 );
and ( n266332 , n266331 , n239229 );
nor ( n266333 , n266330 , n266332 );
nand ( n266334 , n266323 , n266333 );
or ( n266335 , n266312 , n266334 );
not ( n266336 , n266323 );
not ( n266337 , n266310 );
not ( n266338 , n266337 );
or ( n266339 , n266336 , n266338 );
nor ( n266340 , n266333 , n258327 );
nand ( n266341 , n266339 , n266340 );
nand ( n266342 , n256673 , n26295 );
nand ( n266343 , n266335 , n266341 , n266342 );
buf ( n266344 , n266343 );
not ( n266345 , n204644 );
not ( n266346 , n251465 );
or ( n266347 , n266345 , n266346 );
not ( n266348 , n252692 );
nand ( n266349 , n266348 , n263556 );
not ( n266350 , n263570 );
and ( n266351 , n266349 , n266350 );
not ( n266352 , n266349 );
and ( n266353 , n266352 , n263570 );
nor ( n266354 , n266351 , n266353 );
or ( n266355 , n266354 , n256214 );
nand ( n266356 , n266347 , n266355 );
buf ( n266357 , n266356 );
not ( n266358 , RI19ab5118_2416);
or ( n266359 , n233507 , n266358 );
not ( n266360 , RI19aab410_2487);
or ( n266361 , n25335 , n266360 );
nand ( n266362 , n266359 , n266361 );
buf ( n266363 , n266362 );
not ( n266364 , RI19a86318_2751);
or ( n266365 , n25328 , n266364 );
or ( n266366 , n25336 , n254185 );
nand ( n266367 , n266365 , n266366 );
buf ( n266368 , n266367 );
not ( n266369 , n43603 );
not ( n266370 , n242270 );
or ( n266371 , n266369 , n266370 );
not ( n266372 , n43603 );
nand ( n266373 , n266372 , n252503 );
nand ( n266374 , n266371 , n266373 );
and ( n266375 , n266374 , n252553 );
not ( n266376 , n266374 );
and ( n266377 , n266376 , n252562 );
nor ( n266378 , n266375 , n266377 );
not ( n266379 , n266378 );
not ( n266380 , n39152 );
not ( n266381 , n246826 );
or ( n266382 , n266380 , n266381 );
not ( n266383 , n39152 );
nand ( n266384 , n266383 , n246835 );
nand ( n266385 , n266382 , n266384 );
and ( n266386 , n266385 , n246883 );
not ( n266387 , n266385 );
and ( n266388 , n266387 , n246892 );
nor ( n266389 , n266386 , n266388 );
not ( n266390 , n39724 );
not ( n266391 , n266390 );
not ( n266392 , n35409 );
or ( n266393 , n266391 , n266392 );
not ( n266394 , n266390 );
nand ( n266395 , n266394 , n35417 );
nand ( n266396 , n266393 , n266395 );
and ( n266397 , n266396 , n249601 );
not ( n266398 , n266396 );
and ( n266399 , n266398 , n249611 );
nor ( n266400 , n266397 , n266399 );
not ( n266401 , n266400 );
nand ( n266402 , n266389 , n266401 );
nand ( n266403 , n266379 , n266402 , n253393 );
nor ( n266404 , n266400 , n37724 );
nand ( n266405 , n266378 , n266404 , n266389 );
nand ( n266406 , n35431 , n205559 );
nand ( n266407 , n266403 , n266405 , n266406 );
buf ( n266408 , n266407 );
buf ( n266409 , n30317 );
buf ( n266410 , n205267 );
buf ( n266411 , n204606 );
or ( n266412 , n25328 , n262583 );
not ( n266413 , RI19aa53f8_2528);
or ( n266414 , n25335 , n266413 );
nand ( n266415 , n266412 , n266414 );
buf ( n266416 , n266415 );
not ( n266417 , n252424 );
not ( n266418 , n257952 );
or ( n266419 , n266417 , n266418 );
not ( n266420 , n252424 );
nand ( n266421 , n266420 , n257956 );
nand ( n266422 , n266419 , n266421 );
and ( n266423 , n266422 , n257964 );
not ( n266424 , n266422 );
and ( n266425 , n266424 , n257960 );
nor ( n266426 , n266423 , n266425 );
nand ( n266427 , n264615 , n266426 );
nor ( n266428 , n226557 , n225956 );
not ( n266429 , n266428 );
not ( n266430 , n225957 );
nand ( n266431 , n266430 , n226557 );
nand ( n266432 , n266429 , n266431 );
and ( n266433 , n266432 , n266099 );
not ( n266434 , n266432 );
and ( n266435 , n266434 , n260471 );
nor ( n266436 , n266433 , n266435 );
nor ( n266437 , n266436 , n31572 );
not ( n266438 , n266437 );
or ( n266439 , n266427 , n266438 );
not ( n266440 , n266436 );
nor ( n266441 , n266440 , n256413 );
nand ( n266442 , n266441 , n266427 );
nand ( n266443 , n238638 , n32964 );
nand ( n266444 , n266439 , n266442 , n266443 );
buf ( n266445 , n266444 );
not ( n266446 , RI19aa71f8_2515);
or ( n266447 , n226819 , n266446 );
not ( n266448 , RI19a9dbf8_2586);
or ( n266449 , n226822 , n266448 );
nand ( n266450 , n266447 , n266449 );
buf ( n266451 , n266450 );
buf ( n266452 , n33089 );
buf ( n266453 , n205127 );
buf ( n266454 , n34857 );
buf ( n266455 , n39953 );
buf ( n266456 , n33359 );
not ( n266457 , n248102 );
not ( n266458 , n266457 );
not ( n266459 , n256901 );
or ( n266460 , n266458 , n266459 );
or ( n266461 , n256901 , n266457 );
nand ( n266462 , n266460 , n266461 );
not ( n266463 , n266462 );
not ( n266464 , n255596 );
and ( n266465 , n266463 , n266464 );
and ( n266466 , n266462 , n255596 );
nor ( n266467 , n266465 , n266466 );
nand ( n266468 , n266467 , n254528 );
not ( n266469 , n246123 );
not ( n266470 , n245602 );
or ( n266471 , n266469 , n266470 );
not ( n266472 , n246123 );
nand ( n266473 , n266472 , n245611 );
nand ( n266474 , n266471 , n266473 );
and ( n266475 , n266474 , n253746 );
not ( n266476 , n266474 );
and ( n266477 , n266476 , n245618 );
nor ( n266478 , n266475 , n266477 );
not ( n266479 , n266478 );
not ( n266480 , n264187 );
nand ( n266481 , n266479 , n266480 );
or ( n266482 , n266468 , n266481 );
not ( n266483 , n266479 );
not ( n266484 , n266467 );
or ( n266485 , n266483 , n266484 );
nor ( n266486 , n266480 , n33254 );
nand ( n266487 , n266485 , n266486 );
nand ( n266488 , n39766 , n205042 );
nand ( n266489 , n266482 , n266487 , n266488 );
buf ( n266490 , n266489 );
not ( n266491 , n34542 );
not ( n266492 , n255116 );
or ( n266493 , n266491 , n266492 );
not ( n266494 , n46836 );
not ( n266495 , n266494 );
not ( n266496 , n250019 );
or ( n266497 , n266495 , n266496 );
not ( n266498 , n266494 );
nand ( n266499 , n266498 , n250028 );
nand ( n266500 , n266497 , n266499 );
and ( n266501 , n266500 , n258316 );
not ( n266502 , n266500 );
and ( n266503 , n266502 , n258319 );
nor ( n266504 , n266501 , n266503 );
not ( n266505 , n237868 );
not ( n266506 , n44750 );
not ( n266507 , n237810 );
or ( n266508 , n266506 , n266507 );
nand ( n266509 , n237817 , n222512 );
nand ( n266510 , n266508 , n266509 );
not ( n266511 , n266510 );
or ( n266512 , n266505 , n266511 );
or ( n266513 , n266510 , n237868 );
nand ( n266514 , n266512 , n266513 );
nand ( n266515 , n266504 , n266514 );
not ( n266516 , n237666 );
not ( n266517 , n266516 );
not ( n266518 , n233997 );
or ( n266519 , n266517 , n266518 );
not ( n266520 , n266516 );
nand ( n266521 , n266520 , n44176 );
nand ( n266522 , n266519 , n266521 );
and ( n266523 , n266522 , n44316 );
not ( n266524 , n266522 );
and ( n266525 , n266524 , n44325 );
nor ( n266526 , n266523 , n266525 );
not ( n266527 , n266526 );
and ( n266528 , n266515 , n266527 );
not ( n266529 , n266515 );
and ( n266530 , n266529 , n266526 );
nor ( n266531 , n266528 , n266530 );
or ( n266532 , n266531 , n255135 );
nand ( n266533 , n266493 , n266532 );
buf ( n266534 , n266533 );
buf ( n266535 , n216717 );
buf ( n266536 , n26168 );
buf ( n266537 , n26329 );
buf ( n266538 , n30343 );
not ( n266539 , n244329 );
not ( n266540 , n29962 );
or ( n266541 , n266539 , n266540 );
not ( n266542 , n244329 );
nand ( n266543 , n266542 , n256362 );
nand ( n266544 , n266541 , n266543 );
and ( n266545 , n266544 , n256366 );
not ( n266546 , n266544 );
and ( n266547 , n266546 , n263797 );
nor ( n266548 , n266545 , n266547 );
not ( n266549 , n266548 );
buf ( n266550 , n53130 );
not ( n266551 , n266550 );
not ( n266552 , n235072 );
or ( n266553 , n266551 , n266552 );
or ( n266554 , n42436 , n266550 );
nand ( n266555 , n266553 , n266554 );
not ( n266556 , n266555 );
not ( n266557 , n235203 );
and ( n266558 , n266556 , n266557 );
and ( n266559 , n266555 , n235203 );
nor ( n266560 , n266558 , n266559 );
nand ( n266561 , n266549 , n266560 );
not ( n266562 , n248853 );
not ( n266563 , n237340 );
or ( n266564 , n266562 , n266563 );
not ( n266565 , n248853 );
nand ( n266566 , n266565 , n237350 );
nand ( n266567 , n266564 , n266566 );
and ( n266568 , n266567 , n252567 );
not ( n266569 , n266567 );
and ( n266570 , n266569 , n256279 );
nor ( n266571 , n266568 , n266570 );
not ( n266572 , n266571 );
nor ( n266573 , n266572 , n243434 );
not ( n266574 , n266573 );
or ( n266575 , n266561 , n266574 );
nor ( n266576 , n266571 , n43517 );
nand ( n266577 , n266561 , n266576 );
nand ( n266578 , n239240 , n30075 );
nand ( n266579 , n266575 , n266577 , n266578 );
buf ( n266580 , n266579 );
or ( n266581 , n25328 , n265020 );
not ( n266582 , RI19aafcb8_2455);
or ( n266583 , n25335 , n266582 );
nand ( n266584 , n266581 , n266583 );
buf ( n266585 , n266584 );
not ( n266586 , n28587 );
not ( n266587 , n254441 );
or ( n266588 , n266586 , n266587 );
nand ( n266589 , n243698 , n251090 );
not ( n266590 , n226933 );
not ( n266591 , n223266 );
or ( n266592 , n266590 , n266591 );
not ( n266593 , n226933 );
nand ( n266594 , n266593 , n45506 );
nand ( n266595 , n266592 , n266594 );
and ( n266596 , n266595 , n45728 );
not ( n266597 , n266595 );
and ( n266598 , n266597 , n265029 );
nor ( n266599 , n266596 , n266598 );
not ( n266600 , n266599 );
and ( n266601 , n266589 , n266600 );
not ( n266602 , n266589 );
and ( n266603 , n266602 , n266599 );
nor ( n266604 , n266601 , n266603 );
or ( n266605 , n266604 , n254470 );
nand ( n266606 , n266588 , n266605 );
buf ( n266607 , n266606 );
nor ( n266608 , n258088 , n256481 );
not ( n266609 , n246752 );
not ( n266610 , n45261 );
or ( n266611 , n266609 , n266610 );
not ( n266612 , n246752 );
nand ( n266613 , n266612 , n45253 );
nand ( n266614 , n266611 , n266613 );
and ( n266615 , n266614 , n255245 );
not ( n266616 , n266614 );
and ( n266617 , n266616 , n255248 );
nor ( n266618 , n266615 , n266617 );
not ( n266619 , n266618 );
nand ( n266620 , n266608 , n258076 , n266619 );
not ( n266621 , n258087 );
not ( n266622 , n258076 );
or ( n266623 , n266621 , n266622 );
nor ( n266624 , n266619 , n239237 );
nand ( n266625 , n266623 , n266624 );
nand ( n266626 , n31577 , n34525 );
nand ( n266627 , n266620 , n266625 , n266626 );
buf ( n266628 , n266627 );
buf ( n266629 , n29450 );
buf ( n266630 , n240166 );
not ( n266631 , n25319 );
nand ( n266632 , n266631 , n25326 );
not ( n266633 , n25324 );
or ( n266634 , n266632 , n266633 );
not ( n266635 , RI19ad04a8_2209);
or ( n266636 , n266635 , RI1754c610_2);
nand ( n266637 , n266634 , n266636 );
buf ( n266638 , n266637 );
not ( n266639 , n247861 );
not ( n266640 , n54537 );
or ( n266641 , n266639 , n266640 );
not ( n266642 , n247861 );
nand ( n266643 , n266642 , n246188 );
nand ( n266644 , n266641 , n266643 );
and ( n266645 , n266644 , n244889 );
not ( n266646 , n266644 );
and ( n266647 , n266646 , n246193 );
nor ( n266648 , n266645 , n266647 );
nand ( n266649 , n266648 , n262313 );
nand ( n266650 , n266649 , n53001 , n205649 );
nor ( n266651 , n262314 , n55146 );
not ( n266652 , n53001 );
nand ( n266653 , n266651 , n266652 , n266648 );
nand ( n266654 , n234453 , n34151 );
nand ( n266655 , n266650 , n266653 , n266654 );
buf ( n266656 , n266655 );
or ( n266657 , n25328 , n256570 );
not ( n266658 , RI19a9c5f0_2595);
or ( n266659 , n25335 , n266658 );
nand ( n266660 , n266657 , n266659 );
buf ( n266661 , n266660 );
not ( n266662 , n253435 );
not ( n266663 , n253807 );
or ( n266664 , n266662 , n266663 );
or ( n266665 , n253807 , n253435 );
nand ( n266666 , n266664 , n266665 );
not ( n266667 , n266666 );
not ( n266668 , n262167 );
or ( n266669 , n266667 , n266668 );
or ( n266670 , n253813 , n266666 );
nand ( n266671 , n266669 , n266670 );
not ( n266672 , n266671 );
nand ( n266673 , n261518 , n266672 );
or ( n266674 , n261531 , n266673 );
not ( n266675 , n261530 );
not ( n266676 , n261518 );
or ( n266677 , n266675 , n266676 );
nor ( n266678 , n266672 , n237384 );
nand ( n266679 , n266677 , n266678 );
nand ( n266680 , n256673 , n34849 );
nand ( n266681 , n266674 , n266679 , n266680 );
buf ( n266682 , n266681 );
not ( n266683 , n253843 );
not ( n266684 , n46514 );
or ( n266685 , n266683 , n266684 );
or ( n266686 , n46514 , n253843 );
nand ( n266687 , n266685 , n266686 );
and ( n266688 , n266687 , n251333 );
not ( n266689 , n266687 );
and ( n266690 , n266689 , n224478 );
nor ( n266691 , n266688 , n266690 );
nand ( n266692 , n266691 , n205649 );
not ( n266693 , n248727 );
not ( n266694 , n55724 );
not ( n266695 , n266694 );
or ( n266696 , n266693 , n266695 );
not ( n266697 , n248727 );
nand ( n266698 , n266697 , n55724 );
nand ( n266699 , n266696 , n266698 );
and ( n266700 , n266699 , n264675 );
not ( n266701 , n266699 );
buf ( n266702 , n264705 );
and ( n266703 , n266701 , n266702 );
nor ( n266704 , n266700 , n266703 );
not ( n266705 , n266514 );
nand ( n266706 , n266704 , n266705 );
or ( n266707 , n266692 , n266706 );
not ( n266708 , n266704 );
not ( n266709 , n266691 );
or ( n266710 , n266708 , n266709 );
nor ( n266711 , n266705 , n250909 );
nand ( n266712 , n266710 , n266711 );
nand ( n266713 , n254798 , n36796 );
nand ( n266714 , n266707 , n266712 , n266713 );
buf ( n266715 , n266714 );
not ( n266716 , RI19ab0ff0_2446);
or ( n266717 , n25328 , n266716 );
not ( n266718 , RI19aa6d48_2517);
or ( n266719 , n25336 , n266718 );
nand ( n266720 , n266717 , n266719 );
buf ( n266721 , n266720 );
not ( n266722 , n245357 );
not ( n266723 , n235366 );
or ( n266724 , n266722 , n266723 );
or ( n266725 , n235366 , n245357 );
nand ( n266726 , n266724 , n266725 );
and ( n266727 , n266726 , n235372 );
not ( n266728 , n266726 );
and ( n266729 , n266728 , n235369 );
nor ( n266730 , n266727 , n266729 );
not ( n266731 , n266730 );
nand ( n266732 , n266731 , n241704 );
not ( n266733 , n253692 );
not ( n266734 , n236096 );
not ( n266735 , n261269 );
or ( n266736 , n266734 , n266735 );
not ( n266737 , n236096 );
nand ( n266738 , n266737 , n256950 );
nand ( n266739 , n266736 , n266738 );
not ( n266740 , n261127 );
xnor ( n266741 , n266739 , n266740 );
not ( n266742 , n266741 );
nand ( n266743 , n266733 , n266742 );
or ( n266744 , n266732 , n266743 );
not ( n266745 , n266733 );
not ( n266746 , n266731 );
or ( n266747 , n266745 , n266746 );
nor ( n266748 , n266742 , n226004 );
nand ( n266749 , n266747 , n266748 );
nand ( n266750 , n231444 , n31698 );
nand ( n266751 , n266744 , n266749 , n266750 );
buf ( n266752 , n266751 );
nand ( n266753 , n258063 , n244809 );
and ( n266754 , n46141 , n231952 );
not ( n266755 , n46141 );
and ( n266756 , n266755 , n54195 );
or ( n266757 , n266754 , n266756 );
and ( n266758 , n266757 , n264879 );
not ( n266759 , n266757 );
and ( n266760 , n266759 , n264882 );
nor ( n266761 , n266758 , n266760 );
nand ( n266762 , n266761 , n266618 );
or ( n266763 , n266753 , n266762 );
nor ( n266764 , n258063 , n49959 );
nand ( n266765 , n266764 , n266762 );
nand ( n266766 , n51381 , n33063 );
nand ( n266767 , n266763 , n266765 , n266766 );
buf ( n266768 , n266767 );
not ( n266769 , RI19aa2248_2551);
or ( n266770 , n226819 , n266769 );
not ( n266771 , RI19a98ae0_2621);
or ( n266772 , n25335 , n266771 );
nand ( n266773 , n266770 , n266772 );
buf ( n266774 , n266773 );
not ( n266775 , n30153 );
not ( n266776 , n39766 );
or ( n266777 , n266775 , n266776 );
not ( n266778 , n49406 );
not ( n266779 , n247119 );
or ( n266780 , n266778 , n266779 );
not ( n266781 , n49406 );
nand ( n266782 , n266781 , n247126 );
nand ( n266783 , n266780 , n266782 );
and ( n266784 , n266783 , n247188 );
not ( n266785 , n266783 );
and ( n266786 , n266785 , n247196 );
nor ( n266787 , n266784 , n266786 );
nand ( n266788 , n251182 , n266787 );
and ( n266789 , n266788 , n258885 );
not ( n266790 , n266788 );
and ( n266791 , n266790 , n251160 );
nor ( n266792 , n266789 , n266791 );
or ( n266793 , n266792 , n49959 );
nand ( n266794 , n266777 , n266793 );
buf ( n266795 , n266794 );
not ( n266796 , n261778 );
not ( n266797 , n266796 );
not ( n266798 , n256770 );
or ( n266799 , n266797 , n266798 );
nor ( n266800 , n256781 , n235895 );
nand ( n266801 , n266799 , n266800 );
nor ( n266802 , n261778 , n258280 );
nand ( n266803 , n266802 , n256770 , n256781 );
nand ( n266804 , n31576 , n30730 );
nand ( n266805 , n266801 , n266803 , n266804 );
buf ( n266806 , n266805 );
not ( n266807 , RI19a9c398_2596);
or ( n266808 , n25328 , n266807 );
not ( n266809 , RI19a922d0_2667);
or ( n266810 , n226822 , n266809 );
nand ( n266811 , n266808 , n266810 );
buf ( n266812 , n266811 );
not ( n266813 , n257643 );
nand ( n266814 , n266813 , n258687 );
or ( n266815 , n257622 , n266814 );
not ( n266816 , n266813 );
not ( n266817 , n257621 );
or ( n266818 , n266816 , n266817 );
nor ( n266819 , n258687 , n244216 );
nand ( n266820 , n266818 , n266819 );
nand ( n266821 , n249622 , n210076 );
nand ( n266822 , n266815 , n266820 , n266821 );
buf ( n266823 , n266822 );
not ( n266824 , n204321 );
not ( n266825 , n234823 );
or ( n266826 , n266824 , n266825 );
nand ( n266827 , n263312 , n263323 );
not ( n266828 , n266827 );
not ( n266829 , n252957 );
not ( n266830 , n233271 );
or ( n266831 , n266829 , n266830 );
not ( n266832 , n252957 );
nand ( n266833 , n266832 , n233264 );
nand ( n266834 , n266831 , n266833 );
not ( n266835 , n256901 );
and ( n266836 , n266834 , n266835 );
not ( n266837 , n266834 );
not ( n266838 , n266835 );
and ( n266839 , n266837 , n266838 );
nor ( n266840 , n266836 , n266839 );
not ( n266841 , n266840 );
not ( n266842 , n266841 );
and ( n266843 , n266828 , n266842 );
and ( n266844 , n266827 , n266841 );
nor ( n266845 , n266843 , n266844 );
or ( n266846 , n266845 , n238223 );
nand ( n266847 , n266826 , n266846 );
buf ( n266848 , n266847 );
not ( n266849 , n245089 );
not ( n266850 , n231768 );
or ( n266851 , n266849 , n266850 );
not ( n266852 , n245089 );
nand ( n266853 , n266852 , n231775 );
nand ( n266854 , n266851 , n266853 );
and ( n266855 , n266854 , n261292 );
not ( n266856 , n266854 );
and ( n266857 , n266856 , n262951 );
nor ( n266858 , n266855 , n266857 );
not ( n266859 , n266858 );
nand ( n266860 , n266859 , n265222 );
not ( n266861 , n265238 );
or ( n266862 , n266860 , n266861 );
nor ( n266863 , n265233 , n252358 );
nand ( n266864 , n266860 , n266863 );
nand ( n266865 , n31577 , n30553 );
nand ( n266866 , n266862 , n266864 , n266865 );
buf ( n266867 , n266866 );
not ( n266868 , n249508 );
nand ( n266869 , n261674 , n266868 );
or ( n266870 , n266869 , n249473 );
nor ( n266871 , n249472 , n244837 );
nand ( n266872 , n266869 , n266871 );
nand ( n266873 , n35431 , n35907 );
nand ( n266874 , n266870 , n266872 , n266873 );
buf ( n266875 , n266874 );
not ( n266876 , RI19abca80_2362);
or ( n266877 , n25328 , n266876 );
not ( n266878 , RI19ab2d78_2433);
or ( n266879 , n226822 , n266878 );
nand ( n266880 , n266877 , n266879 );
buf ( n266881 , n266880 );
nand ( n266882 , n259100 , n260375 );
not ( n266883 , n261101 );
nand ( n266884 , n259124 , n266883 );
or ( n266885 , n266882 , n266884 );
not ( n266886 , n259124 );
not ( n266887 , n259100 );
or ( n266888 , n266886 , n266887 );
nor ( n266889 , n266883 , n234818 );
nand ( n266890 , n266888 , n266889 );
nand ( n266891 , n255116 , n29426 );
nand ( n266892 , n266885 , n266890 , n266891 );
buf ( n266893 , n266892 );
nand ( n266894 , n226569 , n49048 );
not ( n266895 , n251807 );
not ( n266896 , n258512 );
or ( n266897 , n266895 , n266896 );
not ( n266898 , n251807 );
nand ( n266899 , n266898 , n259214 );
nand ( n266900 , n266897 , n266899 );
and ( n266901 , n266900 , n260558 );
not ( n266902 , n266900 );
and ( n266903 , n266902 , n260551 );
nor ( n266904 , n266901 , n266903 );
nor ( n266905 , n266904 , n244399 );
not ( n266906 , n266905 );
or ( n266907 , n266894 , n266906 );
not ( n266908 , n266904 );
not ( n266909 , n266908 );
not ( n266910 , n226569 );
or ( n266911 , n266909 , n266910 );
nor ( n266912 , n49048 , n236795 );
nand ( n266913 , n266911 , n266912 );
nand ( n266914 , n247585 , n26444 );
nand ( n266915 , n266907 , n266913 , n266914 );
buf ( n266916 , n266915 );
not ( n266917 , n204755 );
not ( n266918 , n228364 );
or ( n266919 , n266917 , n266918 );
not ( n266920 , n204755 );
nand ( n266921 , n266920 , n50539 );
nand ( n266922 , n266919 , n266921 );
and ( n266923 , n266922 , n55727 );
not ( n266924 , n266922 );
and ( n266925 , n266924 , n55730 );
nor ( n266926 , n266923 , n266925 );
nand ( n266927 , n266926 , n262658 );
or ( n266928 , n257072 , n266927 );
not ( n266929 , n262658 );
not ( n266930 , n257051 );
or ( n266931 , n266929 , n266930 );
nor ( n266932 , n266926 , n265700 );
nand ( n266933 , n266931 , n266932 );
nand ( n266934 , n238638 , n205127 );
nand ( n266935 , n266928 , n266933 , n266934 );
buf ( n266936 , n266935 );
not ( n266937 , RI19acfb30_2213);
or ( n266938 , n25328 , n266937 );
or ( n266939 , n25336 , n43524 );
nand ( n266940 , n266938 , n266939 );
buf ( n266941 , n266940 );
not ( n266942 , RI19a82970_2776);
or ( n266943 , n25328 , n266942 );
not ( n266944 , RI19ac7b38_2272);
or ( n266945 , n25335 , n266944 );
nand ( n266946 , n266943 , n266945 );
buf ( n266947 , n266946 );
not ( n266948 , n254317 );
not ( n266949 , n251029 );
or ( n266950 , n266948 , n266949 );
not ( n266951 , n254317 );
nand ( n266952 , n266951 , n261127 );
nand ( n266953 , n266950 , n266952 );
and ( n266954 , n266953 , n261130 );
not ( n266955 , n266953 );
and ( n266956 , n266955 , n261133 );
nor ( n266957 , n266954 , n266956 );
nor ( n266958 , n266957 , n262245 );
or ( n266959 , n258385 , n266958 );
nor ( n266960 , n258384 , n266957 );
nor ( n266961 , n262245 , n40465 );
nand ( n266962 , n266960 , n266961 );
nand ( n266963 , n241976 , n25494 );
nand ( n266964 , n266959 , n266962 , n266963 );
buf ( n266965 , n266964 );
not ( n266966 , n248537 );
not ( n266967 , n243659 );
or ( n266968 , n266966 , n266967 );
or ( n266969 , n243659 , n248537 );
nand ( n266970 , n266968 , n266969 );
and ( n266971 , n266970 , n251856 );
not ( n266972 , n266970 );
and ( n266973 , n266972 , n251846 );
nor ( n266974 , n266971 , n266973 );
not ( n266975 , n266974 );
not ( n266976 , n263926 );
nand ( n266977 , n263948 , n266975 , n266976 );
not ( n266978 , n263946 );
not ( n266979 , n266976 );
or ( n266980 , n266978 , n266979 );
nor ( n266981 , n266975 , n238635 );
nand ( n266982 , n266980 , n266981 );
nand ( n266983 , n238114 , n31625 );
nand ( n266984 , n266977 , n266982 , n266983 );
buf ( n266985 , n266984 );
not ( n266986 , RI19a23a38_2791);
or ( n266987 , n25328 , n266986 );
not ( n266988 , RI19a860c0_2752);
or ( n266989 , n25335 , n266988 );
nand ( n266990 , n266987 , n266989 );
buf ( n266991 , n266990 );
buf ( n266992 , n234361 );
not ( n266993 , n266992 );
not ( n266994 , n238106 );
or ( n266995 , n266993 , n266994 );
or ( n266996 , n238106 , n266992 );
nand ( n266997 , n266995 , n266996 );
not ( n266998 , n244390 );
and ( n266999 , n266997 , n266998 );
not ( n267000 , n266997 );
not ( n267001 , n244387 );
and ( n267002 , n267000 , n267001 );
nor ( n267003 , n266999 , n267002 );
not ( n267004 , n265054 );
nor ( n267005 , n267003 , n267004 );
nand ( n267006 , n265057 , n267005 );
not ( n267007 , n265054 );
not ( n267008 , n265033 );
not ( n267009 , n267008 );
or ( n267010 , n267007 , n267009 );
not ( n267011 , n267003 );
nor ( n267012 , n267011 , n258280 );
nand ( n267013 , n267010 , n267012 );
nand ( n267014 , n35431 , n32113 );
nand ( n267015 , n267006 , n267013 , n267014 );
buf ( n267016 , n267015 );
not ( n267017 , n224748 );
not ( n267018 , n267017 );
not ( n267019 , n252823 );
or ( n267020 , n267018 , n267019 );
not ( n267021 , n267017 );
nand ( n267022 , n267021 , n252831 );
nand ( n267023 , n267020 , n267022 );
xnor ( n267024 , n267023 , n252834 );
not ( n267025 , n267024 );
not ( n267026 , n234959 );
not ( n267027 , n236993 );
or ( n267028 , n267026 , n267027 );
or ( n267029 , n236993 , n234959 );
nand ( n267030 , n267028 , n267029 );
and ( n267031 , n267030 , n254125 );
not ( n267032 , n267030 );
and ( n267033 , n267032 , n254122 );
nor ( n267034 , n267031 , n267033 );
nand ( n267035 , n267025 , n267034 );
buf ( n267036 , n245134 );
or ( n267037 , n267036 , n40918 );
nand ( n267038 , n40914 , n267036 );
nand ( n267039 , n267037 , n267038 );
not ( n267040 , n267039 );
not ( n267041 , n264383 );
and ( n267042 , n267040 , n267041 );
and ( n267043 , n267039 , n41217 );
nor ( n267044 , n267042 , n267043 );
not ( n267045 , n267044 );
nor ( n267046 , n267045 , n31572 );
not ( n267047 , n267046 );
or ( n267048 , n267035 , n267047 );
nor ( n267049 , n267044 , n243434 );
nand ( n267050 , n267035 , n267049 );
nand ( n267051 , n234453 , n37434 );
nand ( n267052 , n267048 , n267050 , n267051 );
buf ( n267053 , n267052 );
not ( n267054 , n37377 );
not ( n267055 , n31577 );
or ( n267056 , n267054 , n267055 );
or ( n267057 , n248026 , n238792 );
nand ( n267058 , n238792 , n248026 );
nand ( n267059 , n267057 , n267058 );
not ( n267060 , n267059 );
not ( n267061 , n238895 );
and ( n267062 , n267060 , n267061 );
and ( n267063 , n267059 , n238895 );
nor ( n267064 , n267062 , n267063 );
not ( n267065 , n238073 );
not ( n267066 , n256094 );
or ( n267067 , n267065 , n267066 );
not ( n267068 , n238073 );
nand ( n267069 , n267068 , n260383 );
nand ( n267070 , n267067 , n267069 );
and ( n267071 , n267070 , n247646 );
not ( n267072 , n267070 );
and ( n267073 , n267072 , n247645 );
nor ( n267074 , n267071 , n267073 );
not ( n267075 , n267074 );
nand ( n267076 , n267064 , n267075 );
and ( n267077 , n267076 , n265980 );
not ( n267078 , n267076 );
not ( n267079 , n265980 );
and ( n267080 , n267078 , n267079 );
nor ( n267081 , n267077 , n267080 );
or ( n267082 , n267081 , n238223 );
nand ( n267083 , n267056 , n267082 );
buf ( n267084 , n267083 );
buf ( n267085 , n32560 );
not ( n267086 , n246040 );
not ( n267087 , n267086 );
not ( n267088 , n261076 );
or ( n267089 , n267087 , n267088 );
not ( n267090 , n267086 );
nand ( n267091 , n267090 , n45023 );
nand ( n267092 , n267089 , n267091 );
and ( n267093 , n267092 , n223016 );
not ( n267094 , n267092 );
and ( n267095 , n267094 , n45262 );
nor ( n267096 , n267093 , n267095 );
nand ( n267097 , n267096 , n251859 );
nor ( n267098 , n261739 , n241968 );
or ( n267099 , n267097 , n267098 );
nor ( n267100 , n267096 , n49959 );
nand ( n267101 , n267100 , n267098 );
nand ( n267102 , n256673 , n38062 );
nand ( n267103 , n267099 , n267101 , n267102 );
buf ( n267104 , n267103 );
or ( n267105 , n25328 , n266448 );
not ( n267106 , RI19a93950_2657);
or ( n267107 , n25336 , n267106 );
nand ( n267108 , n267105 , n267107 );
buf ( n267109 , n267108 );
buf ( n267110 , n37090 );
buf ( n267111 , n31962 );
not ( n267112 , n243687 );
not ( n267113 , n245641 );
not ( n267114 , n267113 );
and ( n267115 , n267112 , n267114 );
and ( n267116 , n243687 , n267113 );
nor ( n267117 , n267115 , n267116 );
and ( n267118 , n267117 , n234881 );
not ( n267119 , n267117 );
and ( n267120 , n267119 , n264197 );
nor ( n267121 , n267118 , n267120 );
nand ( n267122 , n267121 , n223839 );
not ( n267123 , n50737 );
not ( n267124 , n255503 );
or ( n267125 , n267123 , n267124 );
or ( n267126 , n255508 , n50737 );
nand ( n267127 , n267125 , n267126 );
and ( n267128 , n267127 , n265402 );
not ( n267129 , n267127 );
and ( n267130 , n267129 , n255515 );
nor ( n267131 , n267128 , n267130 );
not ( n267132 , n267131 );
not ( n267133 , n263848 );
buf ( n267134 , n251063 );
not ( n267135 , n267134 );
not ( n267136 , n267135 );
not ( n267137 , n50474 );
or ( n267138 , n267136 , n267137 );
nand ( n267139 , n50482 , n267134 );
nand ( n267140 , n267138 , n267139 );
not ( n267141 , n267140 );
or ( n267142 , n267133 , n267141 );
or ( n267143 , n267140 , n263848 );
nand ( n267144 , n267142 , n267143 );
not ( n267145 , n267144 );
nand ( n267146 , n267132 , n267145 );
or ( n267147 , n267122 , n267146 );
not ( n267148 , n267132 );
not ( n267149 , n267121 );
or ( n267150 , n267148 , n267149 );
nor ( n267151 , n267145 , n251190 );
nand ( n267152 , n267150 , n267151 );
nand ( n267153 , n241068 , n28852 );
nand ( n267154 , n267147 , n267152 , n267153 );
buf ( n267155 , n267154 );
not ( n267156 , n255574 );
not ( n267157 , n238628 );
or ( n267158 , n267156 , n267157 );
not ( n267159 , n255574 );
nand ( n267160 , n267159 , n238620 );
nand ( n267161 , n267158 , n267160 );
and ( n267162 , n267161 , n257185 );
not ( n267163 , n267161 );
and ( n267164 , n267163 , n257188 );
nor ( n267165 , n267162 , n267164 );
not ( n267166 , n267165 );
nor ( n267167 , n267166 , n260567 );
not ( n267168 , n244299 );
not ( n267169 , n267168 );
not ( n267170 , n29962 );
or ( n267171 , n267169 , n267170 );
nand ( n267172 , n256362 , n244299 );
nand ( n267173 , n267171 , n267172 );
not ( n267174 , n267173 );
not ( n267175 , n256366 );
and ( n267176 , n267174 , n267175 );
and ( n267177 , n267173 , n256366 );
nor ( n267178 , n267176 , n267177 );
not ( n267179 , n267178 );
nand ( n267180 , n267167 , n261411 , n267179 );
nor ( n267181 , n261411 , n37725 );
nand ( n267182 , n267179 , n267165 );
nand ( n267183 , n267181 , n267182 );
nand ( n267184 , n49054 , n29328 );
nand ( n267185 , n267180 , n267183 , n267184 );
buf ( n267186 , n267185 );
buf ( n267187 , n53184 );
not ( n267188 , n267187 );
not ( n267189 , n253673 );
or ( n267190 , n267188 , n267189 );
or ( n267191 , n256768 , n267187 );
nand ( n267192 , n267190 , n267191 );
not ( n267193 , n267192 );
not ( n267194 , n253676 );
and ( n267195 , n267193 , n267194 );
and ( n267196 , n267192 , n253676 );
nor ( n267197 , n267195 , n267196 );
not ( n267198 , n267197 );
nand ( n267199 , n267198 , n226010 );
not ( n267200 , n267199 );
not ( n267201 , n258163 );
nand ( n267202 , n258151 , n267201 );
not ( n267203 , n267202 );
and ( n267204 , n267200 , n267203 );
and ( n267205 , n51381 , n204565 );
nor ( n267206 , n267204 , n267205 );
nand ( n267207 , n267197 , n245241 );
not ( n267208 , n267207 );
nand ( n267209 , n267208 , n258150 );
nand ( n267210 , n258150 , n237385 );
not ( n267211 , n267210 );
nand ( n267212 , n267211 , n258163 );
nand ( n267213 , n267206 , n267209 , n267212 );
buf ( n267214 , n267213 );
not ( n267215 , RI19aa46d8_2534);
or ( n267216 , n25328 , n267215 );
or ( n267217 , n25335 , n250287 );
nand ( n267218 , n267216 , n267217 );
buf ( n267219 , n267218 );
not ( n267220 , n262169 );
not ( n267221 , n233165 );
not ( n267222 , n233967 );
or ( n267223 , n267221 , n267222 );
not ( n267224 , n233165 );
nand ( n267225 , n267224 , n233959 );
nand ( n267226 , n267223 , n267225 );
and ( n267227 , n267226 , n238621 );
not ( n267228 , n267226 );
and ( n267229 , n267228 , n238629 );
nor ( n267230 , n267227 , n267229 );
nand ( n267231 , n267220 , n267230 );
or ( n267232 , n262157 , n267231 );
nor ( n267233 , n262156 , n55152 );
nand ( n267234 , n267233 , n267231 );
nand ( n267235 , n245943 , n43234 );
nand ( n267236 , n267232 , n267234 , n267235 );
buf ( n267237 , n267236 );
buf ( n267238 , n251264 );
not ( n267239 , n267238 );
not ( n267240 , n249006 );
or ( n267241 , n267239 , n267240 );
or ( n267242 , n242574 , n267238 );
nand ( n267243 , n267241 , n267242 );
and ( n267244 , n267243 , n249929 );
not ( n267245 , n267243 );
not ( n267246 , n255493 );
not ( n267247 , n267246 );
and ( n267248 , n267245 , n267247 );
nor ( n267249 , n267244 , n267248 );
not ( n267250 , n267249 );
not ( n267251 , n267250 );
not ( n267252 , n258708 );
or ( n267253 , n267251 , n267252 );
nor ( n267254 , n258734 , n265700 );
nand ( n267255 , n267253 , n267254 );
nor ( n267256 , n267249 , n252258 );
nand ( n267257 , n258708 , n267256 , n258734 );
nand ( n267258 , n245701 , n36901 );
nand ( n267259 , n267255 , n267257 , n267258 );
buf ( n267260 , n267259 );
or ( n267261 , n233507 , n256087 );
not ( n267262 , RI19a89270_2730);
or ( n267263 , n25336 , n267262 );
nand ( n267264 , n267261 , n267263 );
buf ( n267265 , n267264 );
buf ( n267266 , n36221 );
not ( n267267 , n28365 );
not ( n267268 , n245702 );
or ( n267269 , n267267 , n267268 );
nand ( n267270 , n256241 , n256251 );
not ( n267271 , n242132 );
not ( n267272 , n204553 );
or ( n267273 , n267271 , n267272 );
or ( n267274 , n204553 , n242132 );
nand ( n267275 , n267273 , n267274 );
not ( n267276 , n267275 );
not ( n267277 , n27878 );
and ( n267278 , n267276 , n267277 );
and ( n267279 , n267275 , n27878 );
nor ( n267280 , n267278 , n267279 );
not ( n267281 , n267280 );
and ( n267282 , n267270 , n267281 );
not ( n267283 , n267270 );
and ( n267284 , n267283 , n267280 );
nor ( n267285 , n267282 , n267284 );
or ( n267286 , n267285 , n245938 );
nand ( n267287 , n267269 , n267286 );
buf ( n267288 , n267287 );
not ( n267289 , RI19a96740_2637);
or ( n267290 , n25328 , n267289 );
not ( n267291 , RI19a8c6f0_2708);
or ( n267292 , n25336 , n267291 );
nand ( n267293 , n267290 , n267292 );
buf ( n267294 , n267293 );
nor ( n267295 , n249551 , n257130 );
nand ( n267296 , n249530 , n205649 );
or ( n267297 , n267295 , n267296 );
nand ( n267298 , n249532 , n267295 );
nand ( n267299 , n237361 , n35071 );
nand ( n267300 , n267297 , n267298 , n267299 );
buf ( n267301 , n267300 );
not ( n267302 , n26418 );
not ( n267303 , n256877 );
or ( n267304 , n267302 , n267303 );
not ( n267305 , n256876 );
or ( n267306 , n267305 , n26418 );
nand ( n267307 , n267304 , n267306 );
and ( n267308 , n267307 , n50604 );
not ( n267309 , n267307 );
and ( n267310 , n267309 , n50540 );
nor ( n267311 , n267308 , n267310 );
nor ( n267312 , n267311 , n240080 );
not ( n267313 , n242806 );
not ( n267314 , n242977 );
or ( n267315 , n267313 , n267314 );
nand ( n267316 , n242969 , n242807 );
nand ( n267317 , n267315 , n267316 );
and ( n267318 , n267317 , n254063 );
not ( n267319 , n267317 );
and ( n267320 , n267319 , n254060 );
nor ( n267321 , n267318 , n267320 );
nor ( n267322 , n263803 , n267321 );
nand ( n267323 , n267312 , n267322 );
not ( n267324 , n267321 );
not ( n267325 , n267324 );
not ( n267326 , n267311 );
not ( n267327 , n267326 );
or ( n267328 , n267325 , n267327 );
nand ( n267329 , n267328 , n263776 );
nand ( n267330 , n252711 , n55476 );
nand ( n267331 , n267323 , n267329 , n267330 );
buf ( n267332 , n267331 );
not ( n267333 , n248584 );
not ( n267334 , n251855 );
or ( n267335 , n267333 , n267334 );
or ( n267336 , n251855 , n248584 );
nand ( n267337 , n267335 , n267336 );
and ( n267338 , n267337 , n260967 );
not ( n267339 , n267337 );
buf ( n267340 , n236056 );
not ( n267341 , n267340 );
and ( n267342 , n267339 , n267341 );
nor ( n267343 , n267338 , n267342 );
nand ( n267344 , n267343 , n253397 );
nand ( n267345 , n232090 , n52233 );
or ( n267346 , n267344 , n267345 );
nor ( n267347 , n267343 , n258179 );
nand ( n267348 , n267345 , n267347 );
nand ( n267349 , n244484 , n29571 );
nand ( n267350 , n267346 , n267348 , n267349 );
buf ( n267351 , n267350 );
not ( n267352 , n240623 );
not ( n267353 , n247393 );
or ( n267354 , n267352 , n267353 );
not ( n267355 , n240623 );
nand ( n267356 , n267355 , n247399 );
nand ( n267357 , n267354 , n267356 );
buf ( n267358 , n263230 );
and ( n267359 , n267357 , n267358 );
not ( n267360 , n267357 );
and ( n267361 , n267360 , n247349 );
nor ( n267362 , n267359 , n267361 );
nand ( n267363 , n267362 , n262369 );
or ( n267364 , n262359 , n267363 );
nor ( n267365 , n262358 , n31572 );
nand ( n267366 , n267365 , n267363 );
nand ( n267367 , n241976 , n28159 );
nand ( n267368 , n267364 , n267366 , n267367 );
buf ( n267369 , n267368 );
buf ( n267370 , n247365 );
not ( n267371 , n267370 );
not ( n267372 , n240508 );
or ( n267373 , n267371 , n267372 );
or ( n267374 , n240504 , n267370 );
nand ( n267375 , n267373 , n267374 );
and ( n267376 , n267375 , n246168 );
not ( n267377 , n267375 );
and ( n267378 , n267377 , n246173 );
nor ( n267379 , n267376 , n267378 );
not ( n267380 , n242366 );
not ( n267381 , n234013 );
or ( n267382 , n267380 , n267381 );
not ( n267383 , n242366 );
nand ( n267384 , n267383 , n39749 );
nand ( n267385 , n267382 , n267384 );
xnor ( n267386 , n267385 , n258517 );
nand ( n267387 , n267379 , n267386 );
not ( n267388 , n34315 );
not ( n267389 , n244190 );
or ( n267390 , n267388 , n267389 );
not ( n267391 , n34315 );
nand ( n267392 , n267391 , n244199 );
nand ( n267393 , n267390 , n267392 );
and ( n267394 , n267393 , n244204 );
not ( n267395 , n267393 );
and ( n267396 , n267395 , n244208 );
nor ( n267397 , n267394 , n267396 );
not ( n267398 , n267397 );
nor ( n267399 , n267398 , n35427 );
not ( n267400 , n267399 );
or ( n267401 , n267387 , n267400 );
nor ( n267402 , n267397 , n234021 );
nand ( n267403 , n267387 , n267402 );
nand ( n267404 , n245414 , n35133 );
nand ( n267405 , n267401 , n267403 , n267404 );
buf ( n267406 , n267405 );
not ( n267407 , n39454 );
not ( n267408 , n234453 );
or ( n267409 , n267407 , n267408 );
nand ( n267410 , n255261 , n255273 );
not ( n267411 , n260200 );
and ( n267412 , n267410 , n267411 );
not ( n267413 , n267410 );
and ( n267414 , n267413 , n260200 );
nor ( n267415 , n267412 , n267414 );
or ( n267416 , n267415 , n244837 );
nand ( n267417 , n267409 , n267416 );
buf ( n267418 , n267417 );
not ( n267419 , n44477 );
not ( n267420 , n241360 );
or ( n267421 , n267419 , n267420 );
not ( n267422 , n44477 );
nand ( n267423 , n267422 , n241369 );
nand ( n267424 , n267421 , n267423 );
and ( n267425 , n267424 , n258975 );
not ( n267426 , n267424 );
and ( n267427 , n267426 , n258972 );
nor ( n267428 , n267425 , n267427 );
nand ( n267429 , n267428 , n256718 );
or ( n267430 , n267429 , n256726 );
nor ( n267431 , n256703 , n258280 );
nand ( n267432 , n267429 , n267431 );
nand ( n267433 , n256673 , n204949 );
nand ( n267434 , n267430 , n267432 , n267433 );
buf ( n267435 , n267434 );
not ( n267436 , n32148 );
not ( n267437 , n258213 );
or ( n267438 , n267436 , n267437 );
not ( n267439 , n46796 );
not ( n267440 , n250019 );
or ( n267441 , n267439 , n267440 );
not ( n267442 , n46796 );
nand ( n267443 , n267442 , n250028 );
nand ( n267444 , n267441 , n267443 );
and ( n267445 , n267444 , n258316 );
not ( n267446 , n267444 );
and ( n267447 , n267446 , n258319 );
nor ( n267448 , n267445 , n267447 );
not ( n267449 , n267448 );
nand ( n267450 , n267449 , n264054 );
and ( n267451 , n267450 , n264067 );
not ( n267452 , n267450 );
and ( n267453 , n267452 , n264068 );
nor ( n267454 , n267451 , n267453 );
or ( n267455 , n267454 , n255707 );
nand ( n267456 , n267438 , n267455 );
buf ( n267457 , n267456 );
not ( n267458 , n267428 );
not ( n267459 , n243748 );
not ( n267460 , n258257 );
or ( n267461 , n267459 , n267460 );
not ( n267462 , n243748 );
nand ( n267463 , n267462 , n236762 );
nand ( n267464 , n267461 , n267463 );
and ( n267465 , n267464 , n260422 );
not ( n267466 , n267464 );
and ( n267467 , n267466 , n246065 );
nor ( n267468 , n267465 , n267467 );
not ( n267469 , n267468 );
nand ( n267470 , n267458 , n267469 );
or ( n267471 , n256692 , n267470 );
not ( n267472 , n267469 );
not ( n267473 , n256691 );
or ( n267474 , n267472 , n267473 );
nor ( n267475 , n267458 , n246680 );
nand ( n267476 , n267474 , n267475 );
nand ( n267477 , n31577 , n28394 );
nand ( n267478 , n267471 , n267476 , n267477 );
buf ( n267479 , n267478 );
not ( n267480 , n254327 );
not ( n267481 , n261127 );
or ( n267482 , n267480 , n267481 );
or ( n267483 , n261127 , n254327 );
nand ( n267484 , n267482 , n267483 );
and ( n267485 , n267484 , n261133 );
not ( n267486 , n267484 );
and ( n267487 , n267486 , n261130 );
nor ( n267488 , n267485 , n267487 );
nand ( n267489 , n267488 , n253397 );
buf ( n267490 , n264652 );
nand ( n267491 , n264677 , n267490 );
or ( n267492 , n267489 , n267491 );
not ( n267493 , n264652 );
not ( n267494 , n267488 );
or ( n267495 , n267493 , n267494 );
nor ( n267496 , n264677 , n238900 );
nand ( n267497 , n267495 , n267496 );
nand ( n267498 , n49054 , n30462 );
nand ( n267499 , n267492 , n267497 , n267498 );
buf ( n267500 , n267499 );
not ( n267501 , n255429 );
not ( n267502 , n267501 );
not ( n267503 , n33246 );
or ( n267504 , n267502 , n267503 );
not ( n267505 , n267501 );
nand ( n267506 , n267505 , n253530 );
nand ( n267507 , n267504 , n267506 );
and ( n267508 , n267507 , n253536 );
not ( n267509 , n267507 );
and ( n267510 , n267509 , n253533 );
nor ( n267511 , n267508 , n267510 );
not ( n267512 , n245669 );
not ( n267513 , n264189 );
or ( n267514 , n267512 , n267513 );
not ( n267515 , n245669 );
nand ( n267516 , n267515 , n241448 );
nand ( n267517 , n267514 , n267516 );
and ( n267518 , n267517 , n241454 );
not ( n267519 , n267517 );
and ( n267520 , n267519 , n241453 );
nor ( n267521 , n267518 , n267520 );
nor ( n267522 , n267511 , n267521 );
not ( n267523 , n267522 );
and ( n267524 , n249743 , n255879 );
not ( n267525 , n249743 );
and ( n267526 , n267525 , n255884 );
or ( n267527 , n267524 , n267526 );
not ( n267528 , n267527 );
not ( n267529 , n260195 );
and ( n267530 , n267528 , n267529 );
and ( n267531 , n267527 , n260195 );
nor ( n267532 , n267530 , n267531 );
nor ( n267533 , n267532 , n238900 );
not ( n267534 , n267533 );
or ( n267535 , n267523 , n267534 );
not ( n267536 , n267511 );
nor ( n267537 , n267536 , n265700 );
nand ( n267538 , n267537 , n267521 );
nand ( n267539 , n267535 , n267538 );
not ( n267540 , n267539 );
nand ( n267541 , n267532 , n226010 );
not ( n267542 , n267541 );
nand ( n267543 , n267542 , n267511 );
nand ( n267544 , n46083 , n29351 );
nand ( n267545 , n267540 , n267543 , n267544 );
buf ( n267546 , n267545 );
not ( n267547 , n242765 );
not ( n267548 , n242977 );
or ( n267549 , n267547 , n267548 );
not ( n267550 , n242765 );
nand ( n267551 , n267550 , n242969 );
nand ( n267552 , n267549 , n267551 );
and ( n267553 , n267552 , n254063 );
not ( n267554 , n267552 );
and ( n267555 , n267554 , n254060 );
nor ( n267556 , n267553 , n267555 );
nand ( n267557 , n267556 , n241373 );
not ( n267558 , n267557 );
not ( n267559 , n254346 );
and ( n267560 , n267558 , n267559 );
nand ( n267561 , n254269 , n226010 );
nor ( n267562 , n267561 , n267556 );
and ( n267563 , n267562 , n254346 );
nor ( n267564 , n267560 , n267563 );
not ( n267565 , n254271 );
not ( n267566 , n267556 );
not ( n267567 , n267566 );
and ( n267568 , n267565 , n267567 );
and ( n267569 , n41945 , n34365 );
nor ( n267570 , n267568 , n267569 );
nand ( n267571 , n267564 , n267570 );
buf ( n267572 , n267571 );
not ( n267573 , n238452 );
not ( n267574 , n51167 );
or ( n267575 , n267573 , n267574 );
or ( n267576 , n51167 , n238452 );
nand ( n267577 , n267575 , n267576 );
and ( n267578 , n267577 , n51272 );
not ( n267579 , n267577 );
and ( n267580 , n267579 , n265187 );
nor ( n267581 , n267578 , n267580 );
nand ( n267582 , n267581 , n226010 );
not ( n267583 , n246581 );
not ( n267584 , n255455 );
or ( n267585 , n267583 , n267584 );
not ( n267586 , n246581 );
nand ( n267587 , n267586 , n255464 );
nand ( n267588 , n267585 , n267587 );
and ( n267589 , n267588 , n259460 );
not ( n267590 , n267588 );
and ( n267591 , n267590 , n259464 );
nor ( n267592 , n267589 , n267591 );
nor ( n267593 , n267592 , n253285 );
or ( n267594 , n267582 , n267593 );
nor ( n267595 , n267581 , n37725 );
nand ( n267596 , n267595 , n267593 );
nand ( n267597 , n55760 , n28168 );
nand ( n267598 , n267594 , n267596 , n267597 );
buf ( n267599 , n267598 );
not ( n267600 , RI19abc8a0_2363);
or ( n267601 , n25328 , n267600 );
or ( n267602 , n25335 , n261334 );
nand ( n267603 , n267601 , n267602 );
buf ( n267604 , n267603 );
not ( n267605 , n266467 );
nand ( n267606 , n267605 , n223839 );
not ( n267607 , n267606 );
nand ( n267608 , n266480 , n264199 );
not ( n267609 , n267608 );
and ( n267610 , n267607 , n267609 );
and ( n267611 , n51381 , n32059 );
nor ( n267612 , n267610 , n267611 );
not ( n267613 , n266468 );
not ( n267614 , n264199 );
nand ( n267615 , n267613 , n267614 );
nor ( n267616 , n264199 , n251361 );
nand ( n267617 , n267616 , n264187 );
nand ( n267618 , n267612 , n267615 , n267617 );
buf ( n267619 , n267618 );
or ( n267620 , n233507 , n254048 );
not ( n267621 , RI19a905c0_2680);
or ( n267622 , n226822 , n267621 );
nand ( n267623 , n267620 , n267622 );
buf ( n267624 , n267623 );
not ( n267625 , n41173 );
not ( n267626 , n37728 );
or ( n267627 , n267625 , n267626 );
not ( n267628 , n235374 );
nand ( n267629 , n267628 , n235730 );
not ( n267630 , n237615 );
not ( n267631 , n41216 );
or ( n267632 , n267630 , n267631 );
not ( n267633 , n237615 );
nand ( n267634 , n267633 , n233987 );
nand ( n267635 , n267632 , n267634 );
and ( n267636 , n267635 , n233990 );
not ( n267637 , n267635 );
and ( n267638 , n267637 , n253206 );
nor ( n267639 , n267636 , n267638 );
and ( n267640 , n267629 , n267639 );
not ( n267641 , n267629 );
not ( n267642 , n267639 );
and ( n267643 , n267641 , n267642 );
nor ( n267644 , n267640 , n267643 );
or ( n267645 , n267644 , n251462 );
nand ( n267646 , n267627 , n267645 );
buf ( n267647 , n267646 );
not ( n267648 , RI19ad0700_2208);
not ( n267649 , RI19ad21b8_2198);
and ( n267650 , n267648 , n267649 );
nor ( n267651 , n267650 , RI1754c610_2);
buf ( n267652 , n267651 );
not ( n267653 , n48628 );
not ( n267654 , n234420 );
or ( n267655 , n267653 , n267654 );
not ( n267656 , n48628 );
nand ( n267657 , n267656 , n239119 );
nand ( n267658 , n267655 , n267657 );
and ( n267659 , n267658 , n239221 );
not ( n267660 , n267658 );
and ( n267661 , n267660 , n239229 );
nor ( n267662 , n267659 , n267661 );
nor ( n267663 , n267662 , n43968 );
not ( n267664 , n260539 );
not ( n267665 , n50274 );
or ( n267666 , n267664 , n267665 );
not ( n267667 , n260539 );
nand ( n267668 , n267667 , n228042 );
nand ( n267669 , n267666 , n267668 );
and ( n267670 , n267669 , n50475 );
not ( n267671 , n267669 );
and ( n267672 , n267671 , n50483 );
nor ( n267673 , n267670 , n267672 );
not ( n267674 , n267673 );
not ( n267675 , n34773 );
not ( n267676 , n244373 );
or ( n267677 , n267675 , n267676 );
not ( n267678 , n34773 );
nand ( n267679 , n267678 , n240996 );
nand ( n267680 , n267677 , n267679 );
buf ( n267681 , n255071 );
not ( n267682 , n267681 );
and ( n267683 , n267680 , n267682 );
not ( n267684 , n267680 );
and ( n267685 , n267684 , n267681 );
nor ( n267686 , n267683 , n267685 );
nor ( n267687 , n267674 , n267686 );
nand ( n267688 , n267663 , n267687 );
not ( n267689 , n267686 );
not ( n267690 , n267689 );
not ( n267691 , n267662 );
not ( n267692 , n267691 );
or ( n267693 , n267690 , n267692 );
nor ( n267694 , n267673 , n233972 );
nand ( n267695 , n267693 , n267694 );
nand ( n267696 , n237714 , n33868 );
nand ( n267697 , n267688 , n267695 , n267696 );
buf ( n267698 , n267697 );
nor ( n267699 , n264835 , n251862 );
not ( n267700 , n257574 );
nor ( n267701 , n267700 , n257585 );
nand ( n267702 , n267699 , n267701 );
not ( n267703 , n257584 );
not ( n267704 , n264835 );
not ( n267705 , n267704 );
or ( n267706 , n267703 , n267705 );
nor ( n267707 , n257574 , n247212 );
nand ( n267708 , n267706 , n267707 );
nand ( n267709 , n41945 , n204993 );
nand ( n267710 , n267702 , n267708 , n267709 );
buf ( n267711 , n267710 );
not ( n267712 , n54907 );
not ( n267713 , n237936 );
or ( n267714 , n267712 , n267713 );
not ( n267715 , n54907 );
nand ( n267716 , n267715 , n237944 );
nand ( n267717 , n267714 , n267716 );
and ( n267718 , n267717 , n237948 );
not ( n267719 , n267717 );
and ( n267720 , n267719 , n237947 );
nor ( n267721 , n267718 , n267720 );
nand ( n267722 , n267721 , n259847 );
nor ( n267723 , n263230 , n240790 );
not ( n267724 , n267723 );
nand ( n267725 , n263230 , n240790 );
nand ( n267726 , n267724 , n267725 );
and ( n267727 , n267726 , n263235 );
not ( n267728 , n267726 );
not ( n267729 , n263235 );
and ( n267730 , n267728 , n267729 );
nor ( n267731 , n267727 , n267730 );
not ( n267732 , n255516 );
nand ( n267733 , n267731 , n267732 );
or ( n267734 , n267722 , n267733 );
not ( n267735 , n267731 );
not ( n267736 , n267721 );
or ( n267737 , n267735 , n267736 );
nor ( n267738 , n267732 , n39763 );
nand ( n267739 , n267737 , n267738 );
nand ( n267740 , n39767 , n31640 );
nand ( n267741 , n267734 , n267739 , n267740 );
buf ( n267742 , n267741 );
not ( n267743 , RI19ab03c0_2452);
or ( n267744 , n25328 , n267743 );
not ( n267745 , RI19aa6190_2522);
or ( n267746 , n25335 , n267745 );
nand ( n267747 , n267744 , n267746 );
buf ( n267748 , n267747 );
not ( n267749 , n238020 );
not ( n267750 , n258552 );
or ( n267751 , n267749 , n267750 );
or ( n267752 , n258552 , n238020 );
nand ( n267753 , n267751 , n267752 );
and ( n267754 , n267753 , n258557 );
not ( n267755 , n267753 );
and ( n267756 , n267755 , n258560 );
nor ( n267757 , n267754 , n267756 );
nand ( n267758 , n267757 , n253393 );
not ( n267759 , n46331 );
not ( n267760 , n248557 );
or ( n267761 , n267759 , n267760 );
not ( n267762 , n46331 );
nand ( n267763 , n267762 , n248565 );
nand ( n267764 , n267761 , n267763 );
and ( n267765 , n267764 , n248679 );
not ( n267766 , n267764 );
and ( n267767 , n267766 , n248678 );
nor ( n267768 , n267765 , n267767 );
not ( n267769 , n267768 );
not ( n267770 , n232077 );
not ( n267771 , n51336 );
or ( n267772 , n267770 , n267771 );
or ( n267773 , n51343 , n232077 );
nand ( n267774 , n267772 , n267773 );
not ( n267775 , n267774 );
not ( n267776 , n38222 );
or ( n267777 , n267775 , n267776 );
or ( n267778 , n51349 , n267774 );
nand ( n267779 , n267777 , n267778 );
not ( n267780 , n267779 );
nand ( n267781 , n267769 , n267780 );
or ( n267782 , n267758 , n267781 );
not ( n267783 , n267769 );
not ( n267784 , n267757 );
or ( n267785 , n267783 , n267784 );
nor ( n267786 , n267780 , n31572 );
nand ( n267787 , n267785 , n267786 );
nand ( n267788 , n49054 , n32970 );
nand ( n267789 , n267782 , n267787 , n267788 );
buf ( n267790 , n267789 );
not ( n267791 , n34501 );
not ( n267792 , n50615 );
or ( n267793 , n267791 , n267792 );
nand ( n267794 , n255180 , n255183 );
not ( n267795 , n239630 );
not ( n267796 , n36368 );
or ( n267797 , n267795 , n267796 );
nand ( n267798 , n36372 , n239631 );
nand ( n267799 , n267797 , n267798 );
not ( n267800 , n267799 );
not ( n267801 , n36730 );
and ( n267802 , n267800 , n267801 );
and ( n267803 , n267799 , n36730 );
nor ( n267804 , n267802 , n267803 );
not ( n267805 , n267804 );
and ( n267806 , n267794 , n267805 );
not ( n267807 , n267794 );
and ( n267808 , n267807 , n267804 );
nor ( n267809 , n267806 , n267808 );
or ( n267810 , n267809 , n245938 );
nand ( n267811 , n267793 , n267810 );
buf ( n267812 , n267811 );
not ( n267813 , n263365 );
nand ( n267814 , n267813 , n263368 );
and ( n267815 , n248706 , n266694 );
not ( n267816 , n248706 );
and ( n267817 , n267816 , n265746 );
or ( n267818 , n267815 , n267817 );
not ( n267819 , n266702 );
and ( n267820 , n267818 , n267819 );
not ( n267821 , n267818 );
and ( n267822 , n267821 , n264672 );
nor ( n267823 , n267820 , n267822 );
nor ( n267824 , n267823 , n40465 );
not ( n267825 , n267824 );
or ( n267826 , n267814 , n267825 );
not ( n267827 , n267823 );
nor ( n267828 , n267827 , n254150 );
nand ( n267829 , n267814 , n267828 );
nand ( n267830 , n241976 , n36646 );
nand ( n267831 , n267826 , n267829 , n267830 );
buf ( n267832 , n267831 );
nand ( n267833 , n234340 , n56075 );
or ( n267834 , n260931 , n267833 );
not ( n267835 , n56075 );
not ( n267836 , n55780 );
or ( n267837 , n267835 , n267836 );
nor ( n267838 , n234340 , n55152 );
nand ( n267839 , n267837 , n267838 );
nand ( n267840 , n31576 , n25662 );
nand ( n267841 , n267834 , n267839 , n267840 );
buf ( n267842 , n267841 );
not ( n267843 , RI19aabb90_2484);
or ( n267844 , n25328 , n267843 );
not ( n267845 , RI19aa19d8_2555);
or ( n267846 , n25335 , n267845 );
nand ( n267847 , n267844 , n267846 );
buf ( n267848 , n267847 );
not ( n267849 , n261463 );
not ( n267850 , n44517 );
not ( n267851 , n267850 );
not ( n267852 , n241360 );
or ( n267853 , n267851 , n267852 );
not ( n267854 , n267850 );
nand ( n267855 , n267854 , n241369 );
nand ( n267856 , n267853 , n267855 );
and ( n267857 , n267856 , n258972 );
not ( n267858 , n267856 );
and ( n267859 , n267858 , n258975 );
nor ( n267860 , n267857 , n267859 );
not ( n267861 , n267860 );
not ( n267862 , n249735 );
not ( n267863 , n255884 );
or ( n267864 , n267862 , n267863 );
not ( n267865 , n249735 );
nand ( n267866 , n267865 , n255879 );
nand ( n267867 , n267864 , n267866 );
and ( n267868 , n267867 , n260195 );
not ( n267869 , n267867 );
and ( n267870 , n267869 , n260198 );
nor ( n267871 , n267868 , n267870 );
nor ( n267872 , n267861 , n267871 );
or ( n267873 , n267849 , n267872 );
nor ( n267874 , n261491 , n247698 );
nand ( n267875 , n267874 , n267872 );
nand ( n267876 , n241976 , n29893 );
nand ( n267877 , n267873 , n267875 , n267876 );
buf ( n267878 , n267877 );
not ( n267879 , n45956 );
not ( n267880 , n247931 );
or ( n267881 , n267879 , n267880 );
nand ( n267882 , n247934 , n45957 );
nand ( n267883 , n267881 , n267882 );
xnor ( n267884 , n267883 , n248000 );
not ( n267885 , n267884 );
not ( n267886 , n258605 );
not ( n267887 , n40460 );
or ( n267888 , n267886 , n267887 );
not ( n267889 , n258605 );
nand ( n267890 , n267889 , n251345 );
nand ( n267891 , n267888 , n267890 );
and ( n267892 , n267891 , n253378 );
not ( n267893 , n267891 );
and ( n267894 , n267893 , n261177 );
nor ( n267895 , n267892 , n267894 );
nand ( n267896 , n267885 , n267895 );
nor ( n267897 , n245685 , n249531 );
not ( n267898 , n267897 );
or ( n267899 , n267896 , n267898 );
nand ( n267900 , n267896 , n245527 );
nand ( n267901 , n241378 , n42917 );
nand ( n267902 , n267899 , n267900 , n267901 );
buf ( n267903 , n267902 );
nand ( n267904 , n261330 , n265308 , n265319 );
nand ( n267905 , n265308 , n261328 );
not ( n267906 , n265319 );
nand ( n267907 , n267905 , n267906 , n223839 );
nand ( n267908 , n49054 , n35577 );
nand ( n267909 , n267904 , n267907 , n267908 );
buf ( n267910 , n267909 );
not ( n267911 , n54192 );
not ( n267912 , n240962 );
not ( n267913 , n267912 );
not ( n267914 , n249858 );
or ( n267915 , n267913 , n267914 );
not ( n267916 , n267912 );
nand ( n267917 , n267916 , n257082 );
nand ( n267918 , n267915 , n267917 );
not ( n267919 , n267918 );
or ( n267920 , n267911 , n267919 );
or ( n267921 , n231957 , n267918 );
nand ( n267922 , n267920 , n267921 );
not ( n267923 , n267922 );
nor ( n267924 , n267923 , n40465 );
not ( n267925 , n251433 );
not ( n267926 , n252132 );
or ( n267927 , n267925 , n267926 );
not ( n267928 , n251433 );
nand ( n267929 , n267928 , n252139 );
nand ( n267930 , n267927 , n267929 );
and ( n267931 , n267930 , n252186 );
not ( n267932 , n267930 );
and ( n267933 , n267932 , n263966 );
nor ( n267934 , n267931 , n267933 );
or ( n267935 , n242535 , n227556 );
nand ( n267936 , n227556 , n242535 );
nand ( n267937 , n267935 , n267936 );
and ( n267938 , n267937 , n49950 );
not ( n267939 , n267937 );
and ( n267940 , n267939 , n227707 );
nor ( n267941 , n267938 , n267940 );
not ( n267942 , n267941 );
nor ( n267943 , n267934 , n267942 );
nand ( n267944 , n267924 , n267943 );
nand ( n267945 , n267922 , n267941 );
nand ( n267946 , n267945 , n267934 , n241459 );
nand ( n267947 , n252711 , n35126 );
nand ( n267948 , n267944 , n267946 , n267947 );
buf ( n267949 , n267948 );
buf ( n267950 , n53577 );
not ( n267951 , n267950 );
not ( n267952 , n250496 );
or ( n267953 , n267951 , n267952 );
or ( n267954 , n250498 , n267950 );
nand ( n267955 , n267953 , n267954 );
and ( n267956 , n267955 , n255295 );
not ( n267957 , n267955 );
and ( n267958 , n267957 , n260370 );
nor ( n267959 , n267956 , n267958 );
nand ( n267960 , n267959 , n205649 );
not ( n267961 , n230926 );
not ( n267962 , n253669 );
or ( n267963 , n267961 , n267962 );
not ( n267964 , n230926 );
nand ( n267965 , n267964 , n253673 );
nand ( n267966 , n267963 , n267965 );
and ( n267967 , n267966 , n253679 );
not ( n267968 , n267966 );
and ( n267969 , n267968 , n253676 );
nor ( n267970 , n267967 , n267969 );
not ( n267971 , n267970 );
not ( n267972 , n248738 );
not ( n267973 , n55725 );
or ( n267974 , n267972 , n267973 );
not ( n267975 , n248738 );
nand ( n267976 , n267975 , n55726 );
nand ( n267977 , n267974 , n267976 );
and ( n267978 , n267977 , n267819 );
not ( n267979 , n267977 );
and ( n267980 , n267979 , n264672 );
nor ( n267981 , n267978 , n267980 );
nand ( n267982 , n267971 , n267981 );
or ( n267983 , n267960 , n267982 );
not ( n267984 , n267981 );
not ( n267985 , n267959 );
or ( n267986 , n267984 , n267985 );
nand ( n267987 , n267970 , n244809 );
not ( n267988 , n267987 );
nand ( n267989 , n267986 , n267988 );
nand ( n267990 , n244789 , n32875 );
nand ( n267991 , n267983 , n267989 , n267990 );
buf ( n267992 , n267991 );
nor ( n267993 , n258772 , n235050 );
not ( n267994 , n236610 );
not ( n267995 , n248062 );
or ( n267996 , n267994 , n267995 );
not ( n267997 , n236610 );
not ( n267998 , n248062 );
nand ( n267999 , n267997 , n267998 );
nand ( n268000 , n267996 , n267999 );
and ( n268001 , n268000 , n258033 );
not ( n268002 , n268000 );
not ( n268003 , n258033 );
and ( n268004 , n268002 , n268003 );
nor ( n268005 , n268001 , n268004 );
not ( n268006 , n268005 );
nor ( n268007 , n258340 , n268006 );
nand ( n268008 , n267993 , n268007 );
not ( n268009 , n268005 );
not ( n268010 , n258772 );
not ( n268011 , n268010 );
or ( n268012 , n268009 , n268011 );
nor ( n268013 , n258774 , n254740 );
nand ( n268014 , n268012 , n268013 );
nand ( n268015 , n39767 , n30249 );
nand ( n268016 , n268008 , n268014 , n268015 );
buf ( n268017 , n268016 );
buf ( n268018 , n32811 );
buf ( n268019 , n219510 );
buf ( n268020 , n42917 );
buf ( n268021 , n29725 );
not ( n268022 , n36344 );
not ( n268023 , n245943 );
or ( n268024 , n268022 , n268023 );
not ( n268025 , n256241 );
nand ( n268026 , n268025 , n267280 );
and ( n268027 , n268026 , n256582 );
not ( n268028 , n268026 );
and ( n268029 , n268028 , n256581 );
nor ( n268030 , n268027 , n268029 );
or ( n268031 , n268030 , n262962 );
nand ( n268032 , n268024 , n268031 );
buf ( n268033 , n268032 );
buf ( n268034 , n204922 );
buf ( n268035 , n46027 );
not ( n268036 , n268035 );
not ( n268037 , n247934 );
or ( n268038 , n268036 , n268037 );
or ( n268039 , n259332 , n268035 );
nand ( n268040 , n268038 , n268039 );
and ( n268041 , n268040 , n248000 );
not ( n268042 , n268040 );
and ( n268043 , n268042 , n259339 );
nor ( n268044 , n268041 , n268043 );
nand ( n268045 , n268044 , n222531 );
nor ( n268046 , n235730 , n267639 );
or ( n268047 , n268045 , n268046 );
nor ( n268048 , n268044 , n265700 );
nand ( n268049 , n268048 , n268046 );
nand ( n268050 , n234453 , n33411 );
nand ( n268051 , n268047 , n268049 , n268050 );
buf ( n268052 , n268051 );
not ( n268053 , n256781 );
not ( n268054 , n261767 );
nand ( n268055 , n268053 , n268054 );
or ( n268056 , n256752 , n268055 );
not ( n268057 , n268053 );
not ( n268058 , n256750 );
or ( n268059 , n268057 , n268058 );
nor ( n268060 , n268054 , n39763 );
nand ( n268061 , n268059 , n268060 );
nand ( n268062 , n250916 , n26075 );
nand ( n268063 , n268056 , n268061 , n268062 );
buf ( n268064 , n268063 );
not ( n268065 , n250198 );
not ( n268066 , n249388 );
or ( n268067 , n268065 , n268066 );
or ( n268068 , n243197 , n250198 );
nand ( n268069 , n268067 , n268068 );
and ( n268070 , n268069 , n249395 );
not ( n268071 , n268069 );
and ( n268072 , n268071 , n249398 );
nor ( n268073 , n268070 , n268072 );
not ( n268074 , n52212 );
not ( n268075 , n268074 );
not ( n268076 , n236267 );
or ( n268077 , n268075 , n268076 );
nand ( n268078 , n245210 , n52212 );
nand ( n268079 , n268077 , n268078 );
not ( n268080 , n268079 );
not ( n268081 , n251181 );
and ( n268082 , n268080 , n268081 );
not ( n268083 , n44539 );
and ( n268084 , n268079 , n268083 );
nor ( n268085 , n268082 , n268084 );
not ( n268086 , n268085 );
nand ( n268087 , n268073 , n268086 );
not ( n268088 , n244748 );
not ( n268089 , n268088 );
not ( n268090 , n241877 );
or ( n268091 , n268089 , n268090 );
nand ( n268092 , n241884 , n244748 );
nand ( n268093 , n268091 , n268092 );
not ( n268094 , n268093 );
not ( n268095 , n254235 );
and ( n268096 , n268094 , n268095 );
and ( n268097 , n268093 , n254235 );
nor ( n268098 , n268096 , n268097 );
not ( n268099 , n268098 );
nor ( n268100 , n268099 , n39763 );
not ( n268101 , n268100 );
or ( n268102 , n268087 , n268101 );
nor ( n268103 , n268098 , n254226 );
nand ( n268104 , n268087 , n268103 );
nand ( n268105 , n49054 , n205875 );
nand ( n268106 , n268102 , n268104 , n268105 );
buf ( n268107 , n268106 );
nor ( n268108 , n244983 , n221279 );
not ( n268109 , n253336 );
not ( n268110 , n50492 );
not ( n268111 , n268110 );
not ( n268112 , n35804 );
or ( n268113 , n268111 , n268112 );
nand ( n268114 , n35811 , n50492 );
nand ( n268115 , n268113 , n268114 );
not ( n268116 , n268115 );
or ( n268117 , n268109 , n268116 );
or ( n268118 , n268115 , n253336 );
nand ( n268119 , n268117 , n268118 );
not ( n268120 , n268119 );
nor ( n268121 , n268120 , n244980 );
nand ( n268122 , n268108 , n268121 );
not ( n268123 , n268119 );
not ( n268124 , n244957 );
or ( n268125 , n268123 , n268124 );
nor ( n268126 , n244984 , n252070 );
nand ( n268127 , n268125 , n268126 );
nand ( n268128 , n256673 , n27897 );
nand ( n268129 , n268122 , n268127 , n268128 );
buf ( n268130 , n268129 );
buf ( n268131 , n40127 );
not ( n268132 , RI19ab3de0_2424);
or ( n268133 , n226819 , n268132 );
or ( n268134 , n25336 , n246095 );
nand ( n268135 , n268133 , n268134 );
buf ( n268136 , n268135 );
not ( n268137 , n207116 );
not ( n268138 , n252711 );
or ( n268139 , n268137 , n268138 );
not ( n268140 , n262788 );
not ( n268141 , n30456 );
not ( n268142 , n268141 );
not ( n268143 , n246963 );
or ( n268144 , n268142 , n268143 );
not ( n268145 , n268141 );
nand ( n268146 , n268145 , n246968 );
nand ( n268147 , n268144 , n268146 );
and ( n268148 , n268147 , n247019 );
not ( n268149 , n268147 );
and ( n268150 , n268149 , n247014 );
nor ( n268151 , n268148 , n268150 );
nand ( n268152 , n268140 , n268151 );
buf ( n268153 , n54689 );
not ( n268154 , n268153 );
not ( n268155 , n245517 );
or ( n268156 , n268154 , n268155 );
or ( n268157 , n257706 , n268153 );
nand ( n268158 , n268156 , n268157 );
not ( n268159 , n251162 );
and ( n268160 , n268158 , n268159 );
not ( n268161 , n268158 );
and ( n268162 , n268161 , n251162 );
nor ( n268163 , n268160 , n268162 );
and ( n268164 , n268152 , n268163 );
not ( n268165 , n268152 );
not ( n268166 , n268163 );
and ( n268167 , n268165 , n268166 );
nor ( n268168 , n268164 , n268167 );
or ( n268169 , n268168 , n258759 );
nand ( n268170 , n268139 , n268169 );
buf ( n268171 , n268170 );
not ( n268172 , n245046 );
not ( n268173 , n268172 );
not ( n268174 , n231768 );
or ( n268175 , n268173 , n268174 );
not ( n268176 , n268172 );
nand ( n268177 , n268176 , n231775 );
nand ( n268178 , n268175 , n268177 );
and ( n268179 , n268178 , n262951 );
not ( n268180 , n268178 );
and ( n268181 , n268180 , n261292 );
nor ( n268182 , n268179 , n268181 );
not ( n268183 , n268182 );
nor ( n268184 , n268183 , n40465 );
not ( n268185 , n40294 );
not ( n268186 , n268185 );
not ( n268187 , n235878 );
or ( n268188 , n268186 , n268187 );
not ( n268189 , n268185 );
nand ( n268190 , n268189 , n235887 );
nand ( n268191 , n268188 , n268190 );
and ( n268192 , n268191 , n259858 );
not ( n268193 , n268191 );
and ( n268194 , n268193 , n259855 );
nor ( n268195 , n268192 , n268194 );
nand ( n268196 , n268184 , n268195 );
not ( n268197 , n46934 );
not ( n268198 , n250019 );
or ( n268199 , n268197 , n268198 );
not ( n268200 , n46934 );
nand ( n268201 , n268200 , n250028 );
nand ( n268202 , n268199 , n268201 );
and ( n268203 , n268202 , n258316 );
not ( n268204 , n268202 );
and ( n268205 , n268204 , n258319 );
nor ( n268206 , n268203 , n268205 );
not ( n268207 , n268206 );
nor ( n268208 , n268207 , n47173 );
nand ( n268209 , n268208 , n268182 );
nor ( n268210 , n268206 , n244399 );
not ( n268211 , n268195 );
nand ( n268212 , n268210 , n268211 , n268183 );
nand ( n268213 , n237714 , n206190 );
nand ( n268214 , n268196 , n268209 , n268212 , n268213 );
buf ( n268215 , n268214 );
buf ( n268216 , n33833 );
buf ( n268217 , n32074 );
not ( n268218 , n260520 );
not ( n268219 , n50274 );
or ( n268220 , n268218 , n268219 );
not ( n268221 , n260520 );
nand ( n268222 , n268221 , n228042 );
nand ( n268223 , n268220 , n268222 );
not ( n268224 , n268223 );
not ( n268225 , n50475 );
and ( n268226 , n268224 , n268225 );
and ( n268227 , n268223 , n50475 );
nor ( n268228 , n268226 , n268227 );
nand ( n268229 , n268228 , n239934 );
not ( n268230 , n45809 );
not ( n268231 , n268230 );
not ( n268232 , n36729 );
or ( n268233 , n268231 , n268232 );
not ( n268234 , n268230 );
nand ( n268235 , n268234 , n249482 );
nand ( n268236 , n268233 , n268235 );
and ( n268237 , n268236 , n249494 );
not ( n268238 , n268236 );
and ( n268239 , n268238 , n249495 );
nor ( n268240 , n268237 , n268239 );
not ( n268241 , n268240 );
not ( n268242 , n229078 );
not ( n268243 , n43005 );
or ( n268244 , n268242 , n268243 );
not ( n268245 , n229078 );
nand ( n268246 , n268245 , n43010 );
nand ( n268247 , n268244 , n268246 );
and ( n268248 , n268247 , n50028 );
not ( n268249 , n268247 );
and ( n268250 , n268249 , n227796 );
nor ( n268251 , n268248 , n268250 );
nand ( n268252 , n268241 , n268251 );
or ( n268253 , n268229 , n268252 );
not ( n268254 , n268251 );
not ( n268255 , n268228 );
or ( n268256 , n268254 , n268255 );
nor ( n268257 , n268241 , n55146 );
nand ( n268258 , n268256 , n268257 );
nand ( n268259 , n252711 , n26171 );
nand ( n268260 , n268253 , n268258 , n268259 );
buf ( n268261 , n268260 );
not ( n268262 , n234613 );
not ( n268263 , n249274 );
or ( n268264 , n268262 , n268263 );
or ( n268265 , n249274 , n234613 );
nand ( n268266 , n268264 , n268265 );
and ( n268267 , n268266 , n249528 );
not ( n268268 , n268266 );
not ( n268269 , n249528 );
and ( n268270 , n268268 , n268269 );
nor ( n268271 , n268267 , n268270 );
nand ( n268272 , n268271 , n257527 );
not ( n268273 , n54527 );
not ( n268274 , n268273 );
not ( n268275 , n251162 );
or ( n268276 , n268274 , n268275 );
not ( n268277 , n268273 );
nand ( n268278 , n268277 , n245473 );
nand ( n268279 , n268276 , n268278 );
and ( n268280 , n268279 , n251168 );
not ( n268281 , n268279 );
and ( n268282 , n268281 , n251171 );
nor ( n268283 , n268280 , n268282 );
nand ( n268284 , n260755 , n268283 );
or ( n268285 , n268272 , n268284 );
not ( n268286 , n268271 );
nand ( n268287 , n268286 , n246697 );
not ( n268288 , n268287 );
nand ( n268289 , n268288 , n268284 );
nand ( n268290 , n31577 , n35692 );
nand ( n268291 , n268285 , n268289 , n268290 );
buf ( n268292 , n268291 );
or ( n268293 , n25328 , n242879 );
or ( n268294 , n226822 , n235062 );
nand ( n268295 , n268293 , n268294 );
buf ( n268296 , n268295 );
not ( n268297 , n239814 );
not ( n268298 , n46708 );
or ( n268299 , n268297 , n268298 );
not ( n268300 , n239814 );
nand ( n268301 , n268300 , n46716 );
nand ( n268302 , n268299 , n268301 );
and ( n268303 , n268302 , n256438 );
not ( n268304 , n268302 );
and ( n268305 , n268304 , n52439 );
nor ( n268306 , n268303 , n268305 );
not ( n268307 , n51499 );
not ( n268308 , n268307 );
not ( n268309 , n239653 );
or ( n268310 , n268308 , n268309 );
not ( n268311 , n268307 );
nand ( n268312 , n268311 , n244125 );
nand ( n268313 , n268310 , n268312 );
and ( n268314 , n268313 , n244978 );
not ( n268315 , n268313 );
and ( n268316 , n268315 , n45877 );
nor ( n268317 , n268314 , n268316 );
not ( n268318 , n268317 );
nor ( n268319 , n268306 , n268318 );
not ( n268320 , n246510 );
nor ( n268321 , n268320 , n255408 );
not ( n268322 , n268321 );
not ( n268323 , n246510 );
nand ( n268324 , n268323 , n236502 );
nand ( n268325 , n268322 , n268324 );
and ( n268326 , n268325 , n255465 );
not ( n268327 , n268325 );
and ( n268328 , n268327 , n255457 );
nor ( n268329 , n268326 , n268328 );
nand ( n268330 , n268329 , n234111 );
or ( n268331 , n268319 , n268330 );
nor ( n268332 , n268329 , n40465 );
nand ( n268333 , n268332 , n268319 );
nand ( n268334 , n251717 , n38340 );
nand ( n268335 , n268331 , n268333 , n268334 );
buf ( n268336 , n268335 );
not ( n268337 , RI19abff78_2332);
or ( n268338 , n25328 , n268337 );
not ( n268339 , RI19ab7008_2402);
or ( n268340 , n25335 , n268339 );
nand ( n268341 , n268338 , n268340 );
buf ( n268342 , n268341 );
or ( n268343 , n233507 , n257479 );
not ( n268344 , RI19ab0000_2454);
or ( n268345 , n25335 , n268344 );
nand ( n268346 , n268343 , n268345 );
buf ( n268347 , n268346 );
not ( n268348 , n28889 );
not ( n268349 , n255116 );
or ( n268350 , n268348 , n268349 );
not ( n268351 , n251016 );
not ( n268352 , n268351 );
not ( n268353 , n245110 );
or ( n268354 , n268352 , n268353 );
not ( n268355 , n268351 );
nand ( n268356 , n268355 , n245114 );
nand ( n268357 , n268354 , n268356 );
and ( n268358 , n268357 , n245171 );
not ( n268359 , n268357 );
and ( n268360 , n268359 , n245174 );
nor ( n268361 , n268358 , n268360 );
nand ( n268362 , n252492 , n268361 );
not ( n268363 , n268362 );
not ( n268364 , n265806 );
and ( n268365 , n268363 , n268364 );
and ( n268366 , n268362 , n265806 );
nor ( n268367 , n268365 , n268366 );
or ( n268368 , n268367 , n35816 );
nand ( n268369 , n268350 , n268368 );
buf ( n268370 , n268369 );
not ( n268371 , n235572 );
not ( n268372 , n248143 );
or ( n268373 , n268371 , n268372 );
not ( n268374 , n235572 );
nand ( n268375 , n268374 , n248135 );
nand ( n268376 , n268373 , n268375 );
and ( n268377 , n268376 , n248149 );
not ( n268378 , n268376 );
and ( n268379 , n268378 , n248146 );
nor ( n268380 , n268377 , n268379 );
nand ( n268381 , n268380 , n38638 );
and ( n268382 , n263042 , n263055 );
or ( n268383 , n268381 , n268382 );
not ( n268384 , n268380 );
nand ( n268385 , n263070 , n268384 , n263055 );
nand ( n268386 , n234453 , n29066 );
nand ( n268387 , n268383 , n268385 , n268386 );
buf ( n268388 , n268387 );
buf ( n268389 , n205053 );
buf ( n268390 , n37187 );
not ( n268391 , n255870 );
not ( n268392 , n51549 );
or ( n268393 , n268391 , n268392 );
or ( n268394 , n51549 , n255870 );
nand ( n268395 , n268393 , n268394 );
and ( n268396 , n268395 , n51598 );
not ( n268397 , n268395 );
and ( n268398 , n268397 , n51607 );
nor ( n268399 , n268396 , n268398 );
nand ( n268400 , n268399 , n254013 );
not ( n268401 , n228680 );
not ( n268402 , n256497 );
or ( n268403 , n268401 , n268402 );
or ( n268404 , n256497 , n228680 );
nand ( n268405 , n268403 , n268404 );
and ( n268406 , n268405 , n251975 );
not ( n268407 , n268405 );
and ( n268408 , n268407 , n256500 );
nor ( n268409 , n268406 , n268408 );
not ( n268410 , n250702 );
buf ( n268411 , n241245 );
not ( n268412 , n268411 );
and ( n268413 , n268410 , n268412 );
and ( n268414 , n250705 , n268411 );
nor ( n268415 , n268413 , n268414 );
xor ( n268416 , n268415 , n250712 );
nor ( n268417 , n268409 , n268416 );
or ( n268418 , n268400 , n268417 );
nor ( n268419 , n268399 , n221279 );
nand ( n268420 , n268419 , n268417 );
nand ( n268421 , n39766 , n32151 );
nand ( n268422 , n268418 , n268420 , n268421 );
buf ( n268423 , n268422 );
or ( n268424 , n25328 , n239795 );
or ( n268425 , n226822 , n266942 );
nand ( n268426 , n268424 , n268425 );
buf ( n268427 , n268426 );
buf ( n268428 , n36359 );
not ( n268429 , n268428 );
not ( n268430 , n249749 );
or ( n268431 , n268429 , n268430 );
or ( n268432 , n249749 , n268428 );
nand ( n268433 , n268431 , n268432 );
and ( n268434 , n268433 , n254644 );
not ( n268435 , n268433 );
and ( n268436 , n268435 , n254647 );
nor ( n268437 , n268434 , n268436 );
nand ( n268438 , n268437 , n255152 );
not ( n268439 , n264714 );
nand ( n268440 , n264702 , n268439 );
or ( n268441 , n268438 , n268440 );
not ( n268442 , n268439 );
not ( n268443 , n268437 );
or ( n268444 , n268442 , n268443 );
nor ( n268445 , n264702 , n234021 );
nand ( n268446 , n268444 , n268445 );
nand ( n268447 , n256673 , n28843 );
nand ( n268448 , n268441 , n268446 , n268447 );
buf ( n268449 , n268448 );
nor ( n268450 , n259486 , n31571 );
not ( n268451 , n268450 );
not ( n268452 , n259826 );
nand ( n268453 , n259498 , n268452 );
or ( n268454 , n268451 , n268453 );
not ( n268455 , n268452 );
not ( n268456 , n259486 );
not ( n268457 , n268456 );
or ( n268458 , n268455 , n268457 );
nor ( n268459 , n259498 , n247276 );
nand ( n268460 , n268458 , n268459 );
nand ( n268461 , n245414 , n204697 );
nand ( n268462 , n268454 , n268460 , n268461 );
buf ( n268463 , n268462 );
not ( n268464 , n247830 );
not ( n268465 , n54537 );
or ( n268466 , n268464 , n268465 );
not ( n268467 , n247830 );
nand ( n268468 , n268467 , n246188 );
nand ( n268469 , n268466 , n268468 );
and ( n268470 , n268469 , n246196 );
not ( n268471 , n268469 );
and ( n268472 , n268471 , n246193 );
nor ( n268473 , n268470 , n268472 );
nand ( n268474 , n268473 , n237385 );
not ( n268475 , n244590 );
and ( n268476 , n236376 , n244583 );
not ( n268477 , n236376 );
and ( n268478 , n268477 , n244574 );
nor ( n268479 , n268476 , n268478 );
not ( n268480 , n268479 );
or ( n268481 , n268475 , n268480 );
not ( n268482 , n268479 );
nand ( n268483 , n268482 , n244586 );
nand ( n268484 , n268481 , n268483 );
not ( n268485 , n268484 );
or ( n268486 , n268474 , n268485 );
nor ( n268487 , n268473 , n39763 );
not ( n268488 , n242585 );
buf ( n268489 , n236467 );
not ( n268490 , n268489 );
and ( n268491 , n268488 , n268490 );
and ( n268492 , n242585 , n268489 );
nor ( n268493 , n268491 , n268492 );
and ( n268494 , n268493 , n33247 );
not ( n268495 , n268493 );
and ( n268496 , n268495 , n261471 );
nor ( n268497 , n268494 , n268496 );
nor ( n268498 , n268497 , n268484 );
nand ( n268499 , n268487 , n268498 );
nand ( n268500 , n268484 , n256957 );
not ( n268501 , n268500 );
not ( n268502 , n268497 );
not ( n268503 , n268502 );
and ( n268504 , n268501 , n268503 );
and ( n268505 , n258743 , n25983 );
nor ( n268506 , n268504 , n268505 );
nand ( n268507 , n268486 , n268499 , n268506 );
buf ( n268508 , n268507 );
not ( n268509 , n259325 );
not ( n268510 , n265349 );
nand ( n268511 , n268510 , n265361 );
or ( n268512 , n268509 , n268511 );
not ( n268513 , n259320 );
not ( n268514 , n268510 );
or ( n268515 , n268513 , n268514 );
nor ( n268516 , n265361 , n254226 );
nand ( n268517 , n268515 , n268516 );
nand ( n268518 , n50615 , n39227 );
nand ( n268519 , n268512 , n268517 , n268518 );
buf ( n268520 , n268519 );
not ( n268521 , n235121 );
not ( n268522 , n248446 );
or ( n268523 , n268521 , n268522 );
not ( n268524 , n235121 );
nand ( n268525 , n268524 , n248455 );
nand ( n268526 , n268523 , n268525 );
and ( n268527 , n268526 , n255830 );
not ( n268528 , n268526 );
and ( n268529 , n268528 , n248386 );
nor ( n268530 , n268527 , n268529 );
nor ( n268531 , n244969 , n268530 );
nand ( n268532 , n268531 , n268126 );
not ( n268533 , n244980 );
not ( n268534 , n244969 );
not ( n268535 , n268534 );
or ( n268536 , n268533 , n268535 );
not ( n268537 , n268530 );
nor ( n268538 , n268537 , n250909 );
nand ( n268539 , n268536 , n268538 );
nand ( n268540 , n255116 , n29022 );
nand ( n268541 , n268532 , n268539 , n268540 );
buf ( n268542 , n268541 );
not ( n268543 , n27752 );
not ( n268544 , n233501 );
or ( n268545 , n268543 , n268544 );
nand ( n268546 , n53679 , n231432 );
not ( n268547 , n235949 );
not ( n268548 , n260557 );
or ( n268549 , n268547 , n268548 );
not ( n268550 , n235949 );
nand ( n268551 , n268550 , n260550 );
nand ( n268552 , n268549 , n268551 );
and ( n268553 , n268552 , n262915 );
not ( n268554 , n268552 );
and ( n268555 , n268554 , n266254 );
nor ( n268556 , n268553 , n268555 );
not ( n268557 , n268556 );
and ( n268558 , n268546 , n268557 );
not ( n268559 , n268546 );
and ( n268560 , n268559 , n268556 );
nor ( n268561 , n268558 , n268560 );
or ( n268562 , n268561 , n235732 );
nand ( n268563 , n268545 , n268562 );
buf ( n268564 , n268563 );
not ( n268565 , n259756 );
not ( n268566 , n247594 );
not ( n268567 , n260600 );
or ( n268568 , n268566 , n268567 );
or ( n268569 , n260600 , n247594 );
nand ( n268570 , n268568 , n268569 );
not ( n268571 , n268570 );
and ( n268572 , n268565 , n268571 );
and ( n268573 , n259756 , n268570 );
nor ( n268574 , n268572 , n268573 );
not ( n268575 , n268574 );
nand ( n268576 , n267448 , n268575 );
not ( n268577 , n268576 );
not ( n268578 , n264055 );
or ( n268579 , n268577 , n268578 );
nor ( n268580 , n268574 , n43517 );
nand ( n268581 , n268580 , n267448 );
not ( n268582 , n268581 );
not ( n268583 , n264053 );
and ( n268584 , n268582 , n268583 );
and ( n268585 , n244789 , n38444 );
nor ( n268586 , n268584 , n268585 );
nand ( n268587 , n268579 , n268586 );
buf ( n268588 , n268587 );
buf ( n268589 , n236687 );
not ( n268590 , n268589 );
not ( n268591 , n43219 );
or ( n268592 , n268590 , n268591 );
or ( n268593 , n43219 , n268589 );
nand ( n268594 , n268592 , n268593 );
and ( n268595 , n268594 , n45027 );
not ( n268596 , n268594 );
and ( n268597 , n268596 , n258039 );
nor ( n268598 , n268595 , n268597 );
nand ( n268599 , n268598 , n230207 );
not ( n268600 , n251753 );
nand ( n268601 , n251743 , n268600 );
or ( n268602 , n268599 , n268601 );
not ( n268603 , n268600 );
not ( n268604 , n268598 );
or ( n268605 , n268603 , n268604 );
nor ( n268606 , n251743 , n252872 );
nand ( n268607 , n268605 , n268606 );
nand ( n268608 , n241378 , n40845 );
nand ( n268609 , n268602 , n268607 , n268608 );
buf ( n268610 , n268609 );
not ( n268611 , n239965 );
not ( n268612 , n255926 );
or ( n268613 , n268611 , n268612 );
not ( n268614 , n239965 );
not ( n268615 , n56039 );
nand ( n268616 , n268614 , n268615 );
nand ( n268617 , n268613 , n268616 );
and ( n268618 , n268617 , n251730 );
not ( n268619 , n268617 );
buf ( n268620 , n40203 );
and ( n268621 , n268619 , n268620 );
nor ( n268622 , n268618 , n268621 );
nor ( n268623 , n268622 , n49959 );
not ( n268624 , n233043 );
not ( n268625 , n53080 );
or ( n268626 , n268624 , n268625 );
not ( n268627 , n233043 );
nand ( n268628 , n268627 , n53077 );
nand ( n268629 , n268626 , n268628 );
and ( n268630 , n268629 , n260957 );
not ( n268631 , n268629 );
and ( n268632 , n268631 , n230903 );
nor ( n268633 , n268630 , n268632 );
not ( n268634 , n54217 );
not ( n268635 , n252185 );
or ( n268636 , n268634 , n268635 );
not ( n268637 , n54217 );
nand ( n268638 , n268637 , n252192 );
nand ( n268639 , n268636 , n268638 );
buf ( n268640 , n51342 );
and ( n268641 , n268639 , n268640 );
not ( n268642 , n268639 );
not ( n268643 , n268640 );
and ( n268644 , n268642 , n268643 );
nor ( n268645 , n268641 , n268644 );
not ( n268646 , n268645 );
nor ( n268647 , n268633 , n268646 );
nand ( n268648 , n268623 , n268647 );
not ( n268649 , n268645 );
not ( n268650 , n268622 );
not ( n268651 , n268650 );
or ( n268652 , n268649 , n268651 );
not ( n268653 , n268633 );
nor ( n268654 , n268653 , n252258 );
nand ( n268655 , n268652 , n268654 );
nand ( n268656 , n31576 , n32223 );
nand ( n268657 , n268648 , n268655 , n268656 );
buf ( n268658 , n268657 );
not ( n268659 , n234217 );
not ( n268660 , n41929 );
or ( n268661 , n268659 , n268660 );
not ( n268662 , n234217 );
nand ( n268663 , n268662 , n41933 );
nand ( n268664 , n268661 , n268663 );
and ( n268665 , n268664 , n262783 );
not ( n268666 , n268664 );
and ( n268667 , n268666 , n262786 );
nor ( n268668 , n268665 , n268667 );
nor ( n268669 , n268668 , n235050 );
not ( n268670 , n239823 );
not ( n268671 , n46708 );
or ( n268672 , n268670 , n268671 );
not ( n268673 , n239823 );
nand ( n268674 , n268673 , n46716 );
nand ( n268675 , n268672 , n268674 );
and ( n268676 , n268675 , n230201 );
not ( n268677 , n268675 );
not ( n268678 , n256438 );
and ( n268679 , n268677 , n268678 );
nor ( n268680 , n268676 , n268679 );
not ( n268681 , n268680 );
not ( n268682 , n42912 );
not ( n268683 , n268682 );
not ( n268684 , n243222 );
or ( n268685 , n268683 , n268684 );
or ( n268686 , n237700 , n268682 );
nand ( n268687 , n268685 , n268686 );
and ( n268688 , n268687 , n243230 );
not ( n268689 , n268687 );
and ( n268690 , n268689 , n243226 );
nor ( n268691 , n268688 , n268690 );
nor ( n268692 , n268681 , n268691 );
nand ( n268693 , n268669 , n268692 );
not ( n268694 , n268691 );
not ( n268695 , n268694 );
not ( n268696 , n268668 );
not ( n268697 , n268696 );
or ( n268698 , n268695 , n268697 );
nor ( n268699 , n268680 , n244216 );
nand ( n268700 , n268698 , n268699 );
nand ( n268701 , n252711 , n32751 );
nand ( n268702 , n268693 , n268700 , n268701 );
buf ( n268703 , n268702 );
not ( n268704 , RI1754c160_12);
or ( n268705 , n51369 , n268704 );
nand ( n268706 , n258185 , n37338 );
nand ( n268707 , n268705 , n268706 );
buf ( n268708 , n268707 );
or ( n268709 , n25328 , n262669 );
not ( n268710 , RI19ab2670_2436);
or ( n268711 , n25335 , n268710 );
nand ( n268712 , n268709 , n268711 );
buf ( n268713 , n268712 );
not ( n268714 , n266175 );
not ( n268715 , n263211 );
nand ( n268716 , n268715 , n263238 );
or ( n268717 , n268714 , n268716 );
not ( n268718 , n268715 );
not ( n268719 , n266156 );
not ( n268720 , n268719 );
or ( n268721 , n268718 , n268720 );
nor ( n268722 , n263238 , n242391 );
nand ( n268723 , n268721 , n268722 );
nand ( n268724 , n234453 , n27786 );
nand ( n268725 , n268717 , n268723 , n268724 );
buf ( n268726 , n268725 );
not ( n268727 , n208980 );
not ( n268728 , n268727 );
not ( n268729 , n247018 );
or ( n268730 , n268728 , n268729 );
nand ( n268731 , n247013 , n208980 );
nand ( n268732 , n268730 , n268731 );
not ( n268733 , n268732 );
not ( n268734 , n250113 );
and ( n268735 , n268733 , n268734 );
and ( n268736 , n268732 , n257128 );
nor ( n268737 , n268735 , n268736 );
nor ( n268738 , n265858 , n268737 );
nand ( n268739 , n265835 , n226010 );
or ( n268740 , n268738 , n268739 );
nand ( n268741 , n265836 , n268738 );
nand ( n268742 , n50615 , n204299 );
nand ( n268743 , n268740 , n268741 , n268742 );
buf ( n268744 , n268743 );
not ( n268745 , n43655 );
not ( n268746 , n242270 );
or ( n268747 , n268745 , n268746 );
not ( n268748 , n43655 );
nand ( n268749 , n268748 , n252503 );
nand ( n268750 , n268747 , n268749 );
and ( n268751 , n268750 , n252562 );
not ( n268752 , n268750 );
and ( n268753 , n268752 , n252553 );
nor ( n268754 , n268751 , n268753 );
nand ( n268755 , n268754 , n43969 );
not ( n268756 , n247792 );
not ( n268757 , n232514 );
or ( n268758 , n268756 , n268757 );
not ( n268759 , n247792 );
nand ( n268760 , n268759 , n232520 );
nand ( n268761 , n268758 , n268760 );
and ( n268762 , n268761 , n232299 );
not ( n268763 , n268761 );
and ( n268764 , n268763 , n247269 );
nor ( n268765 , n268762 , n268764 );
not ( n268766 , n43400 );
not ( n268767 , n238894 );
or ( n268768 , n268766 , n268767 );
not ( n268769 , n43400 );
nand ( n268770 , n268769 , n246077 );
nand ( n268771 , n268768 , n268770 );
and ( n268772 , n268771 , n244453 );
not ( n268773 , n268771 );
and ( n268774 , n268773 , n246082 );
nor ( n268775 , n268772 , n268774 );
nand ( n268776 , n268765 , n268775 );
or ( n268777 , n268755 , n268776 );
not ( n268778 , n268775 );
not ( n268779 , n268754 );
or ( n268780 , n268778 , n268779 );
nor ( n268781 , n268765 , n226955 );
nand ( n268782 , n268780 , n268781 );
nand ( n268783 , n234024 , n31351 );
nand ( n268784 , n268777 , n268782 , n268783 );
buf ( n268785 , n268784 );
not ( n268786 , n38438 );
not ( n268787 , n244789 );
or ( n268788 , n268786 , n268787 );
not ( n268789 , n241041 );
not ( n268790 , n219396 );
or ( n268791 , n268789 , n268790 );
not ( n268792 , n241041 );
nand ( n268793 , n268792 , n41632 );
nand ( n268794 , n268791 , n268793 );
and ( n268795 , n268794 , n41935 );
not ( n268796 , n268794 );
and ( n268797 , n268796 , n41929 );
nor ( n268798 , n268795 , n268797 );
not ( n268799 , n268798 );
not ( n268800 , n235826 );
not ( n268801 , n250754 );
or ( n268802 , n268800 , n268801 );
nand ( n268803 , n245797 , n235825 );
nand ( n268804 , n268802 , n268803 );
not ( n268805 , n263382 );
and ( n268806 , n268804 , n268805 );
not ( n268807 , n268804 );
and ( n268808 , n268807 , n250808 );
nor ( n268809 , n268806 , n268808 );
not ( n268810 , n268809 );
nand ( n268811 , n268799 , n268810 );
not ( n268812 , n255814 );
not ( n268813 , n51061 );
not ( n268814 , n257184 );
or ( n268815 , n268813 , n268814 );
nand ( n268816 , n255762 , n51060 );
nand ( n268817 , n268815 , n268816 );
not ( n268818 , n268817 );
or ( n268819 , n268812 , n268818 );
or ( n268820 , n255814 , n268817 );
nand ( n268821 , n268819 , n268820 );
and ( n268822 , n268811 , n268821 );
not ( n268823 , n268811 );
not ( n268824 , n268821 );
and ( n268825 , n268823 , n268824 );
nor ( n268826 , n268822 , n268825 );
or ( n268827 , n268826 , n258328 );
nand ( n268828 , n268788 , n268827 );
buf ( n268829 , n268828 );
not ( n268830 , RI19ab6ae0_2404);
or ( n268831 , n25328 , n268830 );
not ( n268832 , RI19aad120_2475);
or ( n268833 , n226822 , n268832 );
nand ( n268834 , n268831 , n268833 );
buf ( n268835 , n268834 );
not ( n268836 , RI19a96998_2636);
or ( n268837 , n25328 , n268836 );
not ( n268838 , RI19ace3c0_2223);
or ( n268839 , n226822 , n268838 );
nand ( n268840 , n268837 , n268839 );
buf ( n268841 , n268840 );
not ( n268842 , n35371 );
not ( n268843 , n234453 );
or ( n268844 , n268842 , n268843 );
not ( n268845 , n267681 );
not ( n268846 , n34883 );
not ( n268847 , n268846 );
not ( n268848 , n240996 );
or ( n268849 , n268847 , n268848 );
or ( n268850 , n268846 , n255080 );
nand ( n268851 , n268849 , n268850 );
not ( n268852 , n268851 );
or ( n268853 , n268845 , n268852 );
or ( n268854 , n268851 , n267681 );
nand ( n268855 , n268853 , n268854 );
nand ( n268856 , n251785 , n268855 );
and ( n268857 , n268856 , n251773 );
not ( n268858 , n268856 );
and ( n268859 , n268858 , n251774 );
nor ( n268860 , n268857 , n268859 );
or ( n268861 , n268860 , n35816 );
nand ( n268862 , n268844 , n268861 );
buf ( n268863 , n268862 );
nand ( n268864 , n264450 , n264462 );
or ( n268865 , n247445 , n268864 );
not ( n268866 , n247443 );
not ( n268867 , n264450 );
or ( n268868 , n268866 , n268867 );
nor ( n268869 , n264462 , n235050 );
nand ( n268870 , n268868 , n268869 );
nand ( n268871 , n48251 , n32266 );
nand ( n268872 , n268865 , n268870 , n268871 );
buf ( n268873 , n268872 );
not ( n268874 , n240494 );
not ( n268875 , n268874 );
not ( n268876 , n252644 );
or ( n268877 , n268875 , n268876 );
not ( n268878 , n268874 );
nand ( n268879 , n268878 , n252649 );
nand ( n268880 , n268877 , n268879 );
and ( n268881 , n268880 , n252652 );
not ( n268882 , n268880 );
and ( n268883 , n268882 , n252656 );
nor ( n268884 , n268881 , n268883 );
not ( n268885 , n239984 );
not ( n268886 , n255926 );
or ( n268887 , n268885 , n268886 );
not ( n268888 , n239984 );
nand ( n268889 , n268888 , n268615 );
nand ( n268890 , n268887 , n268889 );
and ( n268891 , n268890 , n251721 );
not ( n268892 , n268890 );
and ( n268893 , n268892 , n268620 );
nor ( n268894 , n268891 , n268893 );
nand ( n268895 , n268884 , n268894 );
not ( n268896 , n255808 );
not ( n268897 , n228789 );
not ( n268898 , n257184 );
or ( n268899 , n268897 , n268898 );
not ( n268900 , n228789 );
nand ( n268901 , n268900 , n255762 );
nand ( n268902 , n268899 , n268901 );
not ( n268903 , n268902 );
or ( n268904 , n268896 , n268903 );
or ( n268905 , n255810 , n268902 );
nand ( n268906 , n268904 , n268905 );
nand ( n268907 , n268906 , n205649 );
or ( n268908 , n268895 , n268907 );
not ( n268909 , n268906 );
not ( n268910 , n268894 );
or ( n268911 , n268909 , n268910 );
nor ( n268912 , n268884 , n260567 );
nand ( n268913 , n268911 , n268912 );
nand ( n268914 , n41945 , n33428 );
nand ( n268915 , n268908 , n268913 , n268914 );
buf ( n268916 , n268915 );
nand ( n268917 , n267662 , n249009 );
not ( n268918 , n206683 );
not ( n268919 , n254866 );
or ( n268920 , n268918 , n268919 );
not ( n268921 , n206683 );
nand ( n268922 , n268921 , n254873 );
nand ( n268923 , n268920 , n268922 );
and ( n268924 , n268923 , n256716 );
not ( n268925 , n268923 );
and ( n268926 , n268925 , n256712 );
nor ( n268927 , n268924 , n268926 );
nand ( n268928 , n268927 , n267689 );
or ( n268929 , n268917 , n268928 );
not ( n268930 , n267662 );
not ( n268931 , n268927 );
or ( n268932 , n268930 , n268931 );
nor ( n268933 , n267689 , n37724 );
nand ( n268934 , n268932 , n268933 );
nand ( n268935 , n237714 , n25526 );
nand ( n268936 , n268929 , n268934 , n268935 );
buf ( n268937 , n268936 );
not ( n268938 , RI19ac74a8_2275);
or ( n268939 , n25328 , n268938 );
not ( n268940 , RI19abe6a0_2346);
or ( n268941 , n25335 , n268940 );
nand ( n268942 , n268939 , n268941 );
buf ( n268943 , n268942 );
buf ( n268944 , n27752 );
buf ( n268945 , n26034 );
buf ( n268946 , n46571 );
buf ( n268947 , n38149 );
not ( n268948 , RI19aa7540_2514);
or ( n268949 , n25328 , n268948 );
not ( n268950 , RI19acfd88_2212);
or ( n268951 , n226822 , n268950 );
nand ( n268952 , n268949 , n268951 );
buf ( n268953 , n268952 );
or ( n268954 , n25328 , n266878 );
not ( n268955 , RI19aa8da0_2504);
or ( n268956 , n25335 , n268955 );
nand ( n268957 , n268954 , n268956 );
buf ( n268958 , n268957 );
not ( n268959 , RI1754a900_64);
or ( n268960 , n249125 , n268959 );
not ( n268961 , RI19ab3a20_2426);
or ( n268962 , n25335 , n268961 );
nand ( n268963 , n268960 , n268962 );
buf ( n268964 , n268963 );
buf ( n268965 , n32763 );
buf ( n268966 , n38073 );
buf ( n268967 , n35271 );
buf ( n268968 , RI19a24c80_2783);
not ( n268969 , n268968 );
not ( n268970 , n257347 );
or ( n268971 , n268969 , n268970 );
nand ( n268972 , n257351 , n257345 );
nand ( n268973 , n268971 , n268972 );
buf ( n268974 , n268973 );
buf ( n268975 , n40845 );
nand ( n268976 , n254405 , n259783 );
not ( n268977 , n46372 );
not ( n268978 , n248557 );
or ( n268979 , n268977 , n268978 );
not ( n268980 , n46372 );
nand ( n268981 , n268980 , n248565 );
nand ( n268982 , n268979 , n268981 );
and ( n268983 , n268982 , n248678 );
not ( n268984 , n268982 );
and ( n268985 , n268984 , n248679 );
nor ( n268986 , n268983 , n268985 );
not ( n268987 , n268986 );
nand ( n268988 , n260716 , n268987 );
or ( n268989 , n268976 , n268988 );
not ( n268990 , n260716 );
not ( n268991 , n254405 );
or ( n268992 , n268990 , n268991 );
nor ( n268993 , n268987 , n247276 );
nand ( n268994 , n268992 , n268993 );
nand ( n268995 , n39766 , n29003 );
nand ( n268996 , n268989 , n268994 , n268995 );
buf ( n268997 , n268996 );
or ( n268998 , n226819 , n261450 );
not ( n268999 , RI19a8bfe8_2711);
or ( n269000 , n226822 , n268999 );
nand ( n269001 , n268998 , n269000 );
buf ( n269002 , n269001 );
nor ( n269003 , n254452 , n236795 );
not ( n269004 , n244650 );
nand ( n269005 , n269003 , n269004 , n254464 );
not ( n269006 , n254452 );
nand ( n269007 , n254464 , n269006 );
nand ( n269008 , n269007 , n244650 , n259783 );
nand ( n269009 , n49054 , n26019 );
nand ( n269010 , n269005 , n269008 , n269009 );
buf ( n269011 , n269010 );
not ( n269012 , n255862 );
not ( n269013 , n269012 );
not ( n269014 , n51549 );
or ( n269015 , n269013 , n269014 );
or ( n269016 , n51549 , n269012 );
nand ( n269017 , n269015 , n269016 );
and ( n269018 , n269017 , n51598 );
not ( n269019 , n269017 );
and ( n269020 , n269019 , n51607 );
nor ( n269021 , n269018 , n269020 );
not ( n269022 , n269021 );
not ( n269023 , n255418 );
not ( n269024 , n33246 );
or ( n269025 , n269023 , n269024 );
not ( n269026 , n255418 );
nand ( n269027 , n269026 , n253530 );
nand ( n269028 , n269025 , n269027 );
and ( n269029 , n269028 , n253533 );
not ( n269030 , n269028 );
and ( n269031 , n269030 , n253536 );
nor ( n269032 , n269029 , n269031 );
nand ( n269033 , n267049 , n269022 , n269032 );
not ( n269034 , n267045 );
not ( n269035 , n269022 );
or ( n269036 , n269034 , n269035 );
nor ( n269037 , n269032 , n251361 );
nand ( n269038 , n269036 , n269037 );
nand ( n269039 , n247423 , n205380 );
nand ( n269040 , n269033 , n269038 , n269039 );
buf ( n269041 , n269040 );
buf ( n269042 , n34211 );
buf ( n269043 , n36145 );
not ( n269044 , n242063 );
not ( n269045 , n246385 );
or ( n269046 , n269044 , n269045 );
not ( n269047 , n242063 );
nand ( n269048 , n269047 , n255822 );
nand ( n269049 , n269046 , n269048 );
and ( n269050 , n269049 , n246449 );
not ( n269051 , n269049 );
and ( n269052 , n269051 , n246441 );
nor ( n269053 , n269050 , n269052 );
or ( n269054 , n255153 , n255180 , n269053 );
not ( n269055 , n255151 );
not ( n269056 , n269053 );
not ( n269057 , n269056 );
or ( n269058 , n269055 , n269057 );
nor ( n269059 , n255181 , n53680 );
nand ( n269060 , n269058 , n269059 );
nand ( n269061 , n247744 , n36836 );
nand ( n269062 , n269054 , n269060 , n269061 );
buf ( n269063 , n269062 );
buf ( n269064 , n28027 );
buf ( n269065 , n217071 );
not ( n269066 , n260352 );
nand ( n269067 , n269066 , n258562 );
not ( n269068 , n258549 );
or ( n269069 , n269067 , n269068 );
nand ( n269070 , n262092 , n269067 );
nand ( n269071 , n234453 , n38538 );
nand ( n269072 , n269069 , n269070 , n269071 );
buf ( n269073 , n269072 );
or ( n269074 , n25328 , n260926 );
not ( n269075 , RI19a9e288_2583);
or ( n269076 , n25336 , n269075 );
nand ( n269077 , n269074 , n269076 );
buf ( n269078 , n269077 );
not ( n269079 , n250462 );
not ( n269080 , n234682 );
or ( n269081 , n269079 , n269080 );
not ( n269082 , n250462 );
nand ( n269083 , n269082 , n234691 );
nand ( n269084 , n269081 , n269083 );
and ( n269085 , n269084 , n234804 );
not ( n269086 , n269084 );
and ( n269087 , n269086 , n234811 );
nor ( n269088 , n269085 , n269087 );
not ( n269089 , n269088 );
nand ( n269090 , n269089 , n257190 );
not ( n269091 , n247969 );
not ( n269092 , n239922 );
or ( n269093 , n269091 , n269092 );
not ( n269094 , n247969 );
nand ( n269095 , n269094 , n239930 );
nand ( n269096 , n269093 , n269095 );
and ( n269097 , n269096 , n243511 );
not ( n269098 , n269096 );
and ( n269099 , n269098 , n243504 );
nor ( n269100 , n269097 , n269099 );
not ( n269101 , n269100 );
nand ( n269102 , n269101 , n241459 );
or ( n269103 , n269090 , n269102 );
not ( n269104 , n269101 );
not ( n269105 , n269089 );
or ( n269106 , n269104 , n269105 );
nor ( n269107 , n257190 , n54208 );
nand ( n269108 , n269106 , n269107 );
nand ( n269109 , n256292 , n28054 );
nand ( n269110 , n269103 , n269108 , n269109 );
buf ( n269111 , n269110 );
buf ( n269112 , n29905 );
not ( n269113 , n240932 );
not ( n269114 , n37714 );
or ( n269115 , n269113 , n269114 );
not ( n269116 , n240932 );
nand ( n269117 , n269116 , n37708 );
nand ( n269118 , n269115 , n269117 );
and ( n269119 , n269118 , n246233 );
not ( n269120 , n269118 );
and ( n269121 , n269120 , n244802 );
nor ( n269122 , n269119 , n269121 );
nor ( n269123 , n269122 , n252258 );
not ( n269124 , n269123 );
not ( n269125 , n230869 );
not ( n269126 , n42436 );
or ( n269127 , n269125 , n269126 );
or ( n269128 , n42436 , n230869 );
nand ( n269129 , n269127 , n269128 );
not ( n269130 , n269129 );
not ( n269131 , n235203 );
and ( n269132 , n269130 , n269131 );
and ( n269133 , n269129 , n235203 );
nor ( n269134 , n269132 , n269133 );
not ( n269135 , n39740 );
not ( n269136 , n35409 );
or ( n269137 , n269135 , n269136 );
not ( n269138 , n39740 );
nand ( n269139 , n269138 , n35417 );
nand ( n269140 , n269137 , n269139 );
and ( n269141 , n269140 , n249611 );
not ( n269142 , n269140 );
and ( n269143 , n269142 , n249601 );
nor ( n269144 , n269141 , n269143 );
nor ( n269145 , n269134 , n269144 );
or ( n269146 , n269124 , n269145 );
nor ( n269147 , n269144 , n247698 );
not ( n269148 , n269134 );
nand ( n269149 , n269147 , n269122 , n269148 );
nand ( n269150 , n39767 , n29188 );
nand ( n269151 , n269146 , n269149 , n269150 );
buf ( n269152 , n269151 );
buf ( n269153 , n29328 );
not ( n269154 , n250414 );
nand ( n269155 , n269154 , n250425 );
not ( n269156 , n254295 );
not ( n269157 , n251029 );
or ( n269158 , n269156 , n269157 );
not ( n269159 , n254295 );
nand ( n269160 , n269159 , n261127 );
nand ( n269161 , n269158 , n269160 );
and ( n269162 , n269161 , n261130 );
not ( n269163 , n269161 );
and ( n269164 , n269163 , n261133 );
nor ( n269165 , n269162 , n269164 );
nand ( n269166 , n269165 , n50945 );
or ( n269167 , n269155 , n269166 );
nor ( n269168 , n269165 , n252070 );
nand ( n269169 , n269155 , n269168 );
nand ( n269170 , n244789 , n205372 );
nand ( n269171 , n269167 , n269169 , n269170 );
buf ( n269172 , n269171 );
not ( n269173 , RI19a9b8d0_2601);
or ( n269174 , n25328 , n269173 );
not ( n269175 , RI19a915b0_2673);
or ( n269176 , n226822 , n269175 );
nand ( n269177 , n269174 , n269176 );
buf ( n269178 , n269177 );
buf ( n269179 , n218775 );
buf ( n269180 , n28738 );
nand ( n269181 , n268824 , n268809 );
not ( n269182 , n253287 );
not ( n269183 , n243079 );
not ( n269184 , n253293 );
or ( n269185 , n269183 , n269184 );
or ( n269186 , n253293 , n243079 );
nand ( n269187 , n269185 , n269186 );
not ( n269188 , n269187 );
or ( n269189 , n269182 , n269188 );
or ( n269190 , n253287 , n269187 );
nand ( n269191 , n269189 , n269190 );
not ( n269192 , n269191 );
nand ( n269193 , n269192 , n256811 );
or ( n269194 , n269181 , n269193 );
nor ( n269195 , n269192 , n55146 );
nand ( n269196 , n269181 , n269195 );
nand ( n269197 , n237361 , n32142 );
nand ( n269198 , n269194 , n269196 , n269197 );
buf ( n269199 , n269198 );
not ( n269200 , n37717 );
not ( n269201 , n36734 );
nand ( n269202 , n269200 , n269201 );
not ( n269203 , n237135 );
not ( n269204 , n253660 );
not ( n269205 , n246660 );
or ( n269206 , n269204 , n269205 );
not ( n269207 , n253660 );
nand ( n269208 , n269207 , n246653 );
nand ( n269209 , n269206 , n269208 );
not ( n269210 , n269209 );
or ( n269211 , n269203 , n269210 );
or ( n269212 , n269209 , n263786 );
nand ( n269213 , n269211 , n269212 );
not ( n269214 , n269213 );
nand ( n269215 , n269214 , n253902 );
or ( n269216 , n269202 , n269215 );
nor ( n269217 , n269214 , n37725 );
nand ( n269218 , n269217 , n269202 );
nand ( n269219 , n35431 , n204339 );
nand ( n269220 , n269216 , n269218 , n269219 );
buf ( n269221 , n269220 );
not ( n269222 , RI19ab1ef0_2440);
or ( n269223 , n25328 , n269222 );
not ( n269224 , RI19aa7e28_2510);
or ( n269225 , n226822 , n269224 );
nand ( n269226 , n269223 , n269225 );
buf ( n269227 , n269226 );
not ( n269228 , RI1754bf08_17);
or ( n269229 , n51369 , n269228 );
nand ( n269230 , n249131 , n25629 );
nand ( n269231 , n269229 , n269230 );
buf ( n269232 , n269231 );
not ( n269233 , n251602 );
not ( n269234 , n55889 );
or ( n269235 , n269233 , n269234 );
not ( n269236 , n251602 );
nand ( n269237 , n269236 , n233660 );
nand ( n269238 , n269235 , n269237 );
not ( n269239 , n56040 );
and ( n269240 , n269238 , n269239 );
not ( n269241 , n269238 );
and ( n269242 , n269241 , n251771 );
nor ( n269243 , n269240 , n269242 );
nand ( n269244 , n269243 , n33255 );
nand ( n269245 , n264035 , n264023 );
or ( n269246 , n269244 , n269245 );
not ( n269247 , n264035 );
not ( n269248 , n269243 );
or ( n269249 , n269247 , n269248 );
nor ( n269250 , n264023 , n246680 );
nand ( n269251 , n269249 , n269250 );
nand ( n269252 , n31577 , n34554 );
nand ( n269253 , n269246 , n269251 , n269252 );
buf ( n269254 , n269253 );
not ( n269255 , RI19a86750_2749);
or ( n269256 , n25328 , n269255 );
not ( n269257 , RI19acb120_2247);
or ( n269258 , n25335 , n269257 );
nand ( n269259 , n269256 , n269258 );
buf ( n269260 , n269259 );
nor ( n269261 , n266504 , n31571 );
nor ( n269262 , n266527 , n266704 );
nand ( n269263 , n269261 , n269262 );
not ( n269264 , n266504 );
not ( n269265 , n269264 );
not ( n269266 , n266526 );
or ( n269267 , n269265 , n269266 );
not ( n269268 , n266704 );
nor ( n269269 , n269268 , n236795 );
nand ( n269270 , n269267 , n269269 );
nand ( n269271 , n252711 , n33057 );
nand ( n269272 , n269263 , n269270 , n269271 );
buf ( n269273 , n269272 );
not ( n269274 , RI19aaa150_2495);
or ( n269275 , n25328 , n269274 );
not ( n269276 , RI19aa05b0_2566);
or ( n269277 , n25336 , n269276 );
nand ( n269278 , n269275 , n269277 );
buf ( n269279 , n269278 );
buf ( n269280 , n29600 );
buf ( n269281 , n32955 );
not ( n269282 , n30051 );
not ( n269283 , n251465 );
or ( n269284 , n269282 , n269283 );
nand ( n269285 , n265392 , n265404 );
not ( n269286 , n269285 );
not ( n269287 , n53950 );
not ( n269288 , n238400 );
or ( n269289 , n269287 , n269288 );
not ( n269290 , n53950 );
nand ( n269291 , n269290 , n238408 );
nand ( n269292 , n269289 , n269291 );
and ( n269293 , n269292 , n251444 );
not ( n269294 , n269292 );
and ( n269295 , n269294 , n251451 );
nor ( n269296 , n269293 , n269295 );
not ( n269297 , n269296 );
and ( n269298 , n269286 , n269297 );
and ( n269299 , n269285 , n269296 );
nor ( n269300 , n269298 , n269299 );
or ( n269301 , n269300 , n256214 );
nand ( n269302 , n269284 , n269301 );
buf ( n269303 , n269302 );
buf ( n269304 , n247339 );
not ( n269305 , n269304 );
not ( n269306 , n251372 );
or ( n269307 , n269305 , n269306 );
or ( n269308 , n246166 , n269304 );
nand ( n269309 , n269307 , n269308 );
and ( n269310 , n269309 , n250692 );
not ( n269311 , n269309 );
and ( n269312 , n269311 , n250682 );
nor ( n269313 , n269310 , n269312 );
not ( n269314 , n269313 );
nand ( n269315 , n269314 , n254013 );
nand ( n269316 , n242277 , n242390 );
or ( n269317 , n269315 , n269316 );
nor ( n269318 , n269314 , n234021 );
nand ( n269319 , n269318 , n269316 );
nand ( n269320 , n256673 , n25947 );
nand ( n269321 , n269317 , n269319 , n269320 );
buf ( n269322 , n269321 );
nand ( n269323 , n257632 , n257643 );
or ( n269324 , n258695 , n269323 );
not ( n269325 , n258674 );
not ( n269326 , n257632 );
or ( n269327 , n269325 , n269326 );
nor ( n269328 , n257643 , n55146 );
nand ( n269329 , n269327 , n269328 );
nand ( n269330 , n237361 , n36145 );
nand ( n269331 , n269324 , n269329 , n269330 );
buf ( n269332 , n269331 );
nand ( n269333 , n262068 , n260879 );
nand ( n269334 , n249867 , n262080 );
or ( n269335 , n269333 , n269334 );
not ( n269336 , n262080 );
not ( n269337 , n262068 );
or ( n269338 , n269336 , n269337 );
nor ( n269339 , n249867 , n33254 );
nand ( n269340 , n269338 , n269339 );
nand ( n269341 , n233501 , n27949 );
nand ( n269342 , n269335 , n269340 , n269341 );
buf ( n269343 , n269342 );
not ( n269344 , n268287 );
not ( n269345 , n260737 );
nand ( n269346 , n269345 , n260748 );
not ( n269347 , n269346 );
and ( n269348 , n269344 , n269347 );
and ( n269349 , n31577 , n28659 );
nor ( n269350 , n269348 , n269349 );
not ( n269351 , n268272 );
not ( n269352 , n260748 );
nand ( n269353 , n269351 , n269352 );
not ( n269354 , n269345 );
nor ( n269355 , n260748 , n244837 );
nand ( n269356 , n269354 , n269355 );
nand ( n269357 , n269350 , n269353 , n269356 );
buf ( n269358 , n269357 );
not ( n269359 , n251883 );
not ( n269360 , n251906 );
nand ( n269361 , n269360 , n259706 );
or ( n269362 , n269359 , n269361 );
not ( n269363 , n259706 );
not ( n269364 , n251895 );
or ( n269365 , n269363 , n269364 );
nor ( n269366 , n269360 , n254740 );
nand ( n269367 , n269365 , n269366 );
nand ( n269368 , n35431 , n33630 );
nand ( n269369 , n269362 , n269367 , n269368 );
buf ( n269370 , n269369 );
not ( n269371 , n223924 );
not ( n269372 , n269371 );
not ( n269373 , n54195 );
or ( n269374 , n269372 , n269373 );
not ( n269375 , n269371 );
nand ( n269376 , n269375 , n231952 );
nand ( n269377 , n269374 , n269376 );
and ( n269378 , n269377 , n264879 );
not ( n269379 , n269377 );
and ( n269380 , n269379 , n264882 );
nor ( n269381 , n269378 , n269380 );
not ( n269382 , n269381 );
nand ( n269383 , n269382 , n267201 );
or ( n269384 , n267207 , n269383 );
not ( n269385 , n269382 );
not ( n269386 , n267197 );
or ( n269387 , n269385 , n269386 );
nor ( n269388 , n267201 , n221279 );
nand ( n269389 , n269387 , n269388 );
nand ( n269390 , n247585 , n34896 );
nand ( n269391 , n269384 , n269389 , n269390 );
buf ( n269392 , n269391 );
not ( n269393 , n260426 );
not ( n269394 , n241229 );
not ( n269395 , n250702 );
or ( n269396 , n269394 , n269395 );
or ( n269397 , n250702 , n241229 );
nand ( n269398 , n269396 , n269397 );
not ( n269399 , n269398 );
not ( n269400 , n245333 );
or ( n269401 , n269399 , n269400 );
not ( n269402 , n245338 );
or ( n269403 , n269402 , n269398 );
nand ( n269404 , n269401 , n269403 );
not ( n269405 , n269404 );
nand ( n269406 , n260071 , n269393 , n269405 );
not ( n269407 , n260065 );
nand ( n269408 , n269407 , n269405 );
not ( n269409 , n251361 );
nand ( n269410 , n269408 , n260426 , n269409 );
nand ( n269411 , n244484 , n32272 );
nand ( n269412 , n269406 , n269410 , n269411 );
buf ( n269413 , n269412 );
buf ( n269414 , n27997 );
buf ( n269415 , n221738 );
buf ( n269416 , n37164 );
not ( n269417 , n234626 );
not ( n269418 , n249522 );
not ( n269419 , n269418 );
or ( n269420 , n269417 , n269419 );
nand ( n269421 , n249522 , n234629 );
nand ( n269422 , n269420 , n269421 );
and ( n269423 , n269422 , n249528 );
not ( n269424 , n269422 );
and ( n269425 , n269424 , n249525 );
nor ( n269426 , n269423 , n269425 );
not ( n269427 , n246046 );
not ( n269428 , n45026 );
or ( n269429 , n269427 , n269428 );
not ( n269430 , n246046 );
nand ( n269431 , n269430 , n45023 );
nand ( n269432 , n269429 , n269431 );
and ( n269433 , n269432 , n223016 );
not ( n269434 , n269432 );
and ( n269435 , n269434 , n45262 );
nor ( n269436 , n269433 , n269435 );
nand ( n269437 , n269426 , n269436 );
not ( n269438 , n52567 );
not ( n269439 , n240052 );
not ( n269440 , n269439 );
not ( n269441 , n269440 );
or ( n269442 , n269438 , n269441 );
or ( n269443 , n240056 , n52567 );
nand ( n269444 , n269442 , n269443 );
not ( n269445 , n269444 );
not ( n269446 , n258610 );
not ( n269447 , n269446 );
not ( n269448 , n269447 );
and ( n269449 , n269445 , n269448 );
and ( n269450 , n269444 , n269447 );
nor ( n269451 , n269449 , n269450 );
nand ( n269452 , n269451 , n248981 );
or ( n269453 , n269437 , n269452 );
nor ( n269454 , n269451 , n55152 );
nand ( n269455 , n269454 , n269437 );
nand ( n269456 , n237714 , n31156 );
nand ( n269457 , n269453 , n269455 , n269456 );
buf ( n269458 , n269457 );
not ( n269459 , n266101 );
nand ( n269460 , n266112 , n269459 );
not ( n269461 , n243475 );
not ( n269462 , n269461 );
not ( n269463 , n236631 );
or ( n269464 , n269462 , n269463 );
not ( n269465 , n269461 );
nand ( n269466 , n269465 , n236637 );
nand ( n269467 , n269464 , n269466 );
and ( n269468 , n269467 , n236763 );
not ( n269469 , n269467 );
and ( n269470 , n269469 , n242699 );
or ( n269471 , n269468 , n269470 );
nor ( n269472 , n269471 , n226003 );
not ( n269473 , n269472 );
or ( n269474 , n269460 , n269473 );
not ( n269475 , n269471 );
nor ( n269476 , n269475 , n226004 );
nand ( n269477 , n269476 , n269460 );
nand ( n269478 , n244789 , n34174 );
nand ( n269479 , n269474 , n269477 , n269478 );
buf ( n269480 , n269479 );
not ( n269481 , RI19abcfa8_2359);
or ( n269482 , n25328 , n269481 );
or ( n269483 , n25335 , n256562 );
nand ( n269484 , n269482 , n269483 );
buf ( n269485 , n269484 );
not ( n269486 , RI19ab8778_2392);
or ( n269487 , n25328 , n269486 );
not ( n269488 , RI19a838e8_2769);
or ( n269489 , n25336 , n269488 );
nand ( n269490 , n269487 , n269489 );
buf ( n269491 , n269490 );
not ( n269492 , n240719 );
not ( n269493 , n247348 );
or ( n269494 , n269492 , n269493 );
not ( n269495 , n240719 );
nand ( n269496 , n269495 , n263230 );
nand ( n269497 , n269494 , n269496 );
and ( n269498 , n269497 , n263235 );
not ( n269499 , n269497 );
and ( n269500 , n269499 , n267729 );
nor ( n269501 , n269498 , n269500 );
nor ( n269502 , n269501 , n233972 );
not ( n269503 , n235319 );
not ( n269504 , n246448 );
or ( n269505 , n269503 , n269504 );
not ( n269506 , n235319 );
nand ( n269507 , n269506 , n246439 );
nand ( n269508 , n269505 , n269507 );
and ( n269509 , n269508 , n250021 );
not ( n269510 , n269508 );
and ( n269511 , n269510 , n250030 );
nor ( n269512 , n269509 , n269511 );
not ( n269513 , n251043 );
not ( n269514 , n50474 );
or ( n269515 , n269513 , n269514 );
not ( n269516 , n251043 );
nand ( n269517 , n269516 , n50482 );
nand ( n269518 , n269515 , n269517 );
and ( n269519 , n269518 , n263851 );
not ( n269520 , n269518 );
and ( n269521 , n269520 , n263848 );
nor ( n269522 , n269519 , n269521 );
not ( n269523 , n269522 );
nand ( n269524 , n269502 , n269512 , n269523 );
not ( n269525 , n269501 );
not ( n269526 , n269525 );
not ( n269527 , n269512 );
or ( n269528 , n269526 , n269527 );
nor ( n269529 , n269523 , n252872 );
nand ( n269530 , n269528 , n269529 );
nand ( n269531 , n256292 , n28476 );
nand ( n269532 , n269524 , n269530 , n269531 );
buf ( n269533 , n269532 );
not ( n269534 , RI19a9e030_2584);
or ( n269535 , n25328 , n269534 );
or ( n269536 , n25335 , n256574 );
nand ( n269537 , n269535 , n269536 );
buf ( n269538 , n269537 );
not ( n269539 , n205010 );
not ( n269540 , n244606 );
or ( n269541 , n269539 , n269540 );
or ( n269542 , n255976 , n51364 );
nand ( n269543 , n269542 , n249125 );
not ( n269544 , n269543 );
not ( n269545 , RI1754ac48_57);
or ( n269546 , n269544 , n269545 );
nand ( n269547 , n269541 , n269546 );
buf ( n269548 , n269547 );
not ( n269549 , n246401 );
not ( n269550 , n256739 );
or ( n269551 , n269549 , n269550 );
or ( n269552 , n256742 , n246401 );
nand ( n269553 , n269551 , n269552 );
not ( n269554 , n269553 );
not ( n269555 , n256748 );
and ( n269556 , n269554 , n269555 );
and ( n269557 , n269553 , n256748 );
nor ( n269558 , n269556 , n269557 );
nor ( n269559 , n269558 , n258369 );
not ( n269560 , n262832 );
nor ( n269561 , n262822 , n269560 );
nand ( n269562 , n269559 , n269561 );
nor ( n269563 , n262832 , n234021 );
not ( n269564 , n269558 );
not ( n269565 , n262822 );
nand ( n269566 , n269564 , n269565 );
nand ( n269567 , n269563 , n269566 );
nand ( n269568 , n231444 , n231153 );
nand ( n269569 , n269562 , n269567 , n269568 );
buf ( n269570 , n269569 );
nand ( n269571 , n253480 , n245241 );
not ( n269572 , n254552 );
not ( n269573 , n269572 );
not ( n269574 , n249462 );
or ( n269575 , n269573 , n269574 );
not ( n269576 , n269572 );
nand ( n269577 , n269576 , n249469 );
nand ( n269578 , n269575 , n269577 );
and ( n269579 , n269578 , n259704 );
not ( n269580 , n269578 );
and ( n269581 , n269580 , n259701 );
nor ( n269582 , n269579 , n269581 );
nand ( n269583 , n253352 , n269582 );
or ( n269584 , n269571 , n269583 );
not ( n269585 , n253352 );
not ( n269586 , n253480 );
or ( n269587 , n269585 , n269586 );
nor ( n269588 , n269582 , n40465 );
nand ( n269589 , n269587 , n269588 );
nand ( n269590 , n31577 , n27943 );
nand ( n269591 , n269584 , n269589 , n269590 );
buf ( n269592 , n269591 );
not ( n269593 , n250702 );
not ( n269594 , n241237 );
not ( n269595 , n269594 );
and ( n269596 , n269593 , n269595 );
and ( n269597 , n250705 , n269594 );
nor ( n269598 , n269596 , n269597 );
and ( n269599 , n269598 , n250708 );
not ( n269600 , n269598 );
and ( n269601 , n269600 , n269402 );
nor ( n269602 , n269599 , n269601 );
not ( n269603 , n269602 );
nor ( n269604 , n269603 , n54208 );
not ( n269605 , n31916 );
not ( n269606 , n250738 );
or ( n269607 , n269605 , n269606 );
not ( n269608 , n31916 );
nand ( n269609 , n269608 , n51269 );
nand ( n269610 , n269607 , n269609 );
and ( n269611 , n269610 , n250746 );
not ( n269612 , n269610 );
buf ( n269613 , n53257 );
and ( n269614 , n269612 , n269613 );
nor ( n269615 , n269611 , n269614 );
nand ( n269616 , n269604 , n269615 , n269522 );
not ( n269617 , n269602 );
not ( n269618 , n269522 );
or ( n269619 , n269617 , n269618 );
nor ( n269620 , n269615 , n234021 );
nand ( n269621 , n269619 , n269620 );
nand ( n269622 , n236798 , n33257 );
nand ( n269623 , n269616 , n269621 , n269622 );
buf ( n269624 , n269623 );
nand ( n269625 , n261552 , n235051 );
nand ( n269626 , n261577 , n262919 );
or ( n269627 , n269625 , n269626 );
not ( n269628 , n261577 );
not ( n269629 , n261552 );
or ( n269630 , n269628 , n269629 );
nand ( n269631 , n269630 , n262920 );
nand ( n269632 , n246217 , n32230 );
nand ( n269633 , n269627 , n269631 , n269632 );
buf ( n269634 , n269633 );
not ( n269635 , RI19ab9c18_2382);
or ( n269636 , n25328 , n269635 );
or ( n269637 , n25335 , n256568 );
nand ( n269638 , n269636 , n269637 );
buf ( n269639 , n269638 );
not ( n269640 , n228151 );
not ( n269641 , n53811 );
or ( n269642 , n269640 , n269641 );
not ( n269643 , n228151 );
nand ( n269644 , n269643 , n53820 );
nand ( n269645 , n269642 , n269644 );
and ( n269646 , n269645 , n231769 );
not ( n269647 , n269645 );
and ( n269648 , n269647 , n231776 );
nor ( n269649 , n269646 , n269648 );
nand ( n269650 , n269649 , n260930 );
nand ( n269651 , n267923 , n267941 );
or ( n269652 , n269650 , n269651 );
not ( n269653 , n267923 );
not ( n269654 , n269649 );
or ( n269655 , n269653 , n269654 );
nor ( n269656 , n267941 , n55104 );
nand ( n269657 , n269655 , n269656 );
nand ( n269658 , n31577 , n205409 );
nand ( n269659 , n269652 , n269657 , n269658 );
buf ( n269660 , n269659 );
not ( n269661 , RI19acb4e0_2245);
or ( n269662 , n25328 , n269661 );
or ( n269663 , n25335 , n265018 );
nand ( n269664 , n269662 , n269663 );
buf ( n269665 , n269664 );
not ( n269666 , n43968 );
buf ( n269667 , n30778 );
not ( n269668 , n269667 );
not ( n269669 , n246968 );
or ( n269670 , n269668 , n269669 );
or ( n269671 , n246968 , n269667 );
nand ( n269672 , n269670 , n269671 );
and ( n269673 , n269672 , n247019 );
not ( n269674 , n269672 );
and ( n269675 , n269674 , n247014 );
nor ( n269676 , n269673 , n269675 );
nand ( n269677 , n269666 , n269676 );
nand ( n269678 , n265719 , n261063 );
or ( n269679 , n269677 , n269678 );
not ( n269680 , n269676 );
not ( n269681 , n261063 );
or ( n269682 , n269680 , n269681 );
nor ( n269683 , n265719 , n235050 );
nand ( n269684 , n269682 , n269683 );
nand ( n269685 , n239240 , n35947 );
nand ( n269686 , n269679 , n269684 , n269685 );
buf ( n269687 , n269686 );
not ( n269688 , RI1754bf80_16);
or ( n269689 , n51369 , n269688 );
nand ( n269690 , n258185 , n30642 );
nand ( n269691 , n269689 , n269690 );
buf ( n269692 , n269691 );
not ( n269693 , n258205 );
nand ( n269694 , n269693 , n252873 );
nor ( n269695 , n242315 , n231821 );
not ( n269696 , n269695 );
nand ( n269697 , n260248 , n231821 );
nand ( n269698 , n269696 , n269697 );
and ( n269699 , n269698 , n242381 );
not ( n269700 , n269698 );
and ( n269701 , n269700 , n242374 );
nor ( n269702 , n269699 , n269701 );
not ( n269703 , n256894 );
nand ( n269704 , n269702 , n269703 );
or ( n269705 , n269694 , n269704 );
not ( n269706 , n269702 );
not ( n269707 , n269693 );
or ( n269708 , n269706 , n269707 );
nor ( n269709 , n269703 , n40465 );
nand ( n269710 , n269708 , n269709 );
nand ( n269711 , n234453 , n39448 );
nand ( n269712 , n269705 , n269710 , n269711 );
buf ( n269713 , n269712 );
buf ( n269714 , n35662 );
buf ( n269715 , n25998 );
not ( n269716 , n29225 );
not ( n269717 , n245943 );
or ( n269718 , n269716 , n269717 );
not ( n269719 , n36029 );
not ( n269720 , n249757 );
or ( n269721 , n269719 , n269720 );
not ( n269722 , n36029 );
nand ( n269723 , n269722 , n249749 );
nand ( n269724 , n269721 , n269723 );
and ( n269725 , n269724 , n254644 );
not ( n269726 , n269724 );
and ( n269727 , n269726 , n254647 );
nor ( n269728 , n269725 , n269727 );
not ( n269729 , n269728 );
not ( n269730 , n249158 );
not ( n269731 , n244776 );
or ( n269732 , n269730 , n269731 );
not ( n269733 , n249158 );
nand ( n269734 , n269733 , n244768 );
nand ( n269735 , n269732 , n269734 );
and ( n269736 , n269735 , n252934 );
not ( n269737 , n269735 );
and ( n269738 , n269737 , n249059 );
nor ( n269739 , n269736 , n269738 );
nand ( n269740 , n269729 , n269739 );
buf ( n269741 , n252906 );
not ( n269742 , n269741 );
not ( n269743 , n264704 );
or ( n269744 , n269742 , n269743 );
or ( n269745 , n264704 , n269741 );
nand ( n269746 , n269744 , n269745 );
and ( n269747 , n269746 , n241057 );
not ( n269748 , n269746 );
and ( n269749 , n269748 , n241060 );
nor ( n269750 , n269747 , n269749 );
not ( n269751 , n269750 );
and ( n269752 , n269740 , n269751 );
not ( n269753 , n269740 );
and ( n269754 , n269753 , n269750 );
nor ( n269755 , n269752 , n269754 );
or ( n269756 , n269755 , n246091 );
nand ( n269757 , n269718 , n269756 );
buf ( n269758 , n269757 );
not ( n269759 , n253767 );
not ( n269760 , n250576 );
or ( n269761 , n269759 , n269760 );
or ( n269762 , n250576 , n253767 );
nand ( n269763 , n269761 , n269762 );
and ( n269764 , n269763 , n252037 );
not ( n269765 , n269763 );
and ( n269766 , n269765 , n252052 );
nor ( n269767 , n269764 , n269766 );
nand ( n269768 , n269767 , n254013 );
not ( n269769 , n257992 );
not ( n269770 , n232790 );
not ( n269771 , n256042 );
or ( n269772 , n269770 , n269771 );
not ( n269773 , n232790 );
nand ( n269774 , n269773 , n237447 );
nand ( n269775 , n269772 , n269774 );
and ( n269776 , n269775 , n237594 );
not ( n269777 , n269775 );
and ( n269778 , n269777 , n237590 );
nor ( n269779 , n269776 , n269778 );
not ( n269780 , n269779 );
nand ( n269781 , n269769 , n269780 );
or ( n269782 , n269768 , n269781 );
not ( n269783 , n269780 );
not ( n269784 , n269767 );
or ( n269785 , n269783 , n269784 );
nor ( n269786 , n269769 , n234440 );
nand ( n269787 , n269785 , n269786 );
nand ( n269788 , n254798 , n38184 );
nand ( n269789 , n269782 , n269787 , n269788 );
buf ( n269790 , n269789 );
buf ( n269791 , n247542 );
not ( n269792 , n269791 );
not ( n269793 , n243810 );
or ( n269794 , n269792 , n269793 );
or ( n269795 , n243810 , n269791 );
nand ( n269796 , n269794 , n269795 );
and ( n269797 , n269796 , n243960 );
not ( n269798 , n269796 );
and ( n269799 , n269798 , n243954 );
nor ( n269800 , n269797 , n269799 );
not ( n269801 , n269800 );
not ( n269802 , n267521 );
nand ( n269803 , n269801 , n269802 );
or ( n269804 , n267541 , n269803 );
not ( n269805 , n269801 );
not ( n269806 , n267532 );
or ( n269807 , n269805 , n269806 );
nor ( n269808 , n269802 , n249531 );
nand ( n269809 , n269807 , n269808 );
nand ( n269810 , n237714 , n25778 );
nand ( n269811 , n269804 , n269809 , n269810 );
buf ( n269812 , n269811 );
not ( n269813 , n31005 );
not ( n269814 , n31577 );
or ( n269815 , n269813 , n269814 );
not ( n269816 , n239231 );
nand ( n269817 , n261947 , n269816 );
not ( n269818 , n261937 );
and ( n269819 , n269817 , n269818 );
not ( n269820 , n269817 );
and ( n269821 , n269820 , n261937 );
nor ( n269822 , n269819 , n269821 );
or ( n269823 , n269822 , n254515 );
nand ( n269824 , n269815 , n269823 );
buf ( n269825 , n269824 );
nand ( n269826 , n258226 , n205649 );
nand ( n269827 , n265333 , n251706 );
or ( n269828 , n269826 , n269827 );
not ( n269829 , n265333 );
not ( n269830 , n258226 );
or ( n269831 , n269829 , n269830 );
nor ( n269832 , n251706 , n219702 );
nand ( n269833 , n269831 , n269832 );
nand ( n269834 , n245701 , n26269 );
nand ( n269835 , n269828 , n269833 , n269834 );
buf ( n269836 , n269835 );
not ( n269837 , RI19a84ba8_2761);
or ( n269838 , n226819 , n269837 );
not ( n269839 , RI19ac9938_2258);
or ( n269840 , n226822 , n269839 );
nand ( n269841 , n269838 , n269840 );
buf ( n269842 , n269841 );
buf ( n269843 , n34022 );
not ( n269844 , n257505 );
not ( n269845 , n243203 );
nand ( n269846 , n269844 , n269845 );
or ( n269847 , n269846 , n257495 );
not ( n269848 , n257493 );
nor ( n269849 , n269848 , n39763 );
nand ( n269850 , n269849 , n269846 );
nand ( n269851 , n241378 , n205795 );
nand ( n269852 , n269847 , n269850 , n269851 );
buf ( n269853 , n269852 );
buf ( n269854 , n205380 );
not ( n269855 , RI19a976b8_2630);
or ( n269856 , n25328 , n269855 );
not ( n269857 , RI19a8d668_2701);
or ( n269858 , n25335 , n269857 );
nand ( n269859 , n269856 , n269858 );
buf ( n269860 , n269859 );
buf ( n269861 , n41698 );
buf ( n269862 , n42665 );
not ( n269863 , n257026 );
not ( n269864 , n263625 );
nand ( n269865 , n263615 , n269864 );
not ( n269866 , n269865 );
and ( n269867 , n269863 , n269866 );
and ( n269868 , n234453 , n210118 );
nor ( n269869 , n269867 , n269868 );
not ( n269870 , n257001 );
nand ( n269871 , n269870 , n264348 );
nand ( n269872 , n264354 , n263625 );
nand ( n269873 , n269869 , n269871 , n269872 );
buf ( n269874 , n269873 );
nand ( n269875 , n259845 , n257527 );
nand ( n269876 , n261266 , n259871 );
or ( n269877 , n269875 , n269876 );
not ( n269878 , n259845 );
not ( n269879 , n261266 );
or ( n269880 , n269878 , n269879 );
nor ( n269881 , n259871 , n226004 );
nand ( n269882 , n269880 , n269881 );
nand ( n269883 , n241068 , n25693 );
nand ( n269884 , n269877 , n269882 , n269883 );
buf ( n269885 , n269884 );
not ( n269886 , n32935 );
not ( n269887 , n51381 );
or ( n269888 , n269886 , n269887 );
nand ( n269889 , n259497 , n259509 );
not ( n269890 , n259816 );
and ( n269891 , n269889 , n269890 );
not ( n269892 , n269889 );
and ( n269893 , n269892 , n259816 );
nor ( n269894 , n269891 , n269893 );
or ( n269895 , n269894 , n238223 );
nand ( n269896 , n269888 , n269895 );
buf ( n269897 , n269896 );
nor ( n269898 , n265110 , n244399 );
nor ( n269899 , n261694 , n261706 );
nand ( n269900 , n269898 , n269899 );
not ( n269901 , n265106 );
not ( n269902 , n265094 );
or ( n269903 , n269901 , n269902 );
nor ( n269904 , n261695 , n40465 );
nand ( n269905 , n269903 , n269904 );
nand ( n269906 , n31577 , n46879 );
nand ( n269907 , n269900 , n269905 , n269906 );
buf ( n269908 , n269907 );
not ( n269909 , n44406 );
not ( n269910 , n269909 );
not ( n269911 , n241360 );
or ( n269912 , n269910 , n269911 );
nand ( n269913 , n241369 , n44406 );
nand ( n269914 , n269912 , n269913 );
not ( n269915 , n269914 );
not ( n269916 , n258972 );
and ( n269917 , n269915 , n269916 );
and ( n269918 , n269914 , n258972 );
nor ( n269919 , n269917 , n269918 );
not ( n269920 , n269919 );
nand ( n269921 , n269920 , n241459 );
not ( n269922 , n35214 );
not ( n269923 , n255072 );
or ( n269924 , n269922 , n269923 );
not ( n269925 , n35214 );
nand ( n269926 , n269925 , n255071 );
nand ( n269927 , n269924 , n269926 );
not ( n269928 , n46420 );
and ( n269929 , n269927 , n269928 );
not ( n269930 , n269927 );
not ( n269931 , n259018 );
and ( n269932 , n269930 , n269931 );
nor ( n269933 , n269929 , n269932 );
not ( n269934 , n269933 );
nand ( n269935 , n253210 , n269934 );
or ( n269936 , n269921 , n269935 );
not ( n269937 , n269934 );
not ( n269938 , n269920 );
or ( n269939 , n269937 , n269938 );
nor ( n269940 , n253210 , n244216 );
nand ( n269941 , n269939 , n269940 );
nand ( n269942 , n263819 , n40547 );
nand ( n269943 , n269936 , n269941 , n269942 );
buf ( n269944 , n269943 );
and ( n269945 , n27883 , n204514 );
buf ( n269946 , n269945 );
or ( n269947 , n25328 , n251918 );
not ( n269948 , RI19a9bb28_2600);
or ( n269949 , n226822 , n269948 );
nand ( n269950 , n269947 , n269949 );
buf ( n269951 , n269950 );
buf ( n269952 , n204399 );
not ( n269953 , n239955 );
not ( n269954 , n56040 );
or ( n269955 , n269953 , n269954 );
not ( n269956 , n239955 );
not ( n269957 , n268615 );
nand ( n269958 , n269956 , n269957 );
nand ( n269959 , n269955 , n269958 );
and ( n269960 , n269959 , n268620 );
not ( n269961 , n269959 );
and ( n269962 , n269961 , n251730 );
nor ( n269963 , n269960 , n269962 );
not ( n269964 , n269963 );
nor ( n269965 , n269964 , n50944 );
not ( n269966 , n258033 );
buf ( n269967 , n236666 );
not ( n269968 , n269967 );
and ( n269969 , n269966 , n269968 );
and ( n269970 , n258033 , n269967 );
nor ( n269971 , n269969 , n269970 );
and ( n269972 , n269971 , n45026 );
not ( n269973 , n269971 );
and ( n269974 , n269973 , n258038 );
nor ( n269975 , n269972 , n269974 );
not ( n269976 , n268640 );
not ( n269977 , n54246 );
not ( n269978 , n252185 );
or ( n269979 , n269977 , n269978 );
or ( n269980 , n252185 , n54246 );
nand ( n269981 , n269979 , n269980 );
not ( n269982 , n269981 );
or ( n269983 , n269976 , n269982 );
or ( n269984 , n269981 , n268640 );
nand ( n269985 , n269983 , n269984 );
nor ( n269986 , n269975 , n269985 );
nand ( n269987 , n269965 , n269986 );
not ( n269988 , n269975 );
nor ( n269989 , n269988 , n235050 );
not ( n269990 , n269985 );
nand ( n269991 , n269963 , n269990 );
nand ( n269992 , n269989 , n269991 );
nand ( n269993 , n256673 , n30547 );
nand ( n269994 , n269987 , n269992 , n269993 );
buf ( n269995 , n269994 );
buf ( n269996 , n28374 );
not ( n269997 , RI19ac2f48_2307);
or ( n269998 , n233507 , n269997 );
not ( n269999 , RI19aba578_2378);
or ( n270000 , n25335 , n269999 );
nand ( n270001 , n269998 , n270000 );
buf ( n270002 , n270001 );
not ( n270003 , n208049 );
not ( n270004 , n254441 );
or ( n270005 , n270003 , n270004 );
nand ( n270006 , n262614 , n262634 );
not ( n270007 , n52747 );
not ( n270008 , n270007 );
not ( n270009 , n258612 );
or ( n270010 , n270008 , n270009 );
not ( n270011 , n270007 );
nand ( n270012 , n270011 , n258611 );
nand ( n270013 , n270010 , n270012 );
and ( n270014 , n270013 , n258622 );
not ( n270015 , n270013 );
and ( n270016 , n270015 , n258618 );
nor ( n270017 , n270014 , n270016 );
not ( n270018 , n270017 );
and ( n270019 , n270006 , n270018 );
not ( n270020 , n270006 );
and ( n270021 , n270020 , n270017 );
nor ( n270022 , n270019 , n270021 );
or ( n270023 , n270022 , n259425 );
nand ( n270024 , n270005 , n270023 );
buf ( n270025 , n270024 );
not ( n270026 , n258589 );
not ( n270027 , n40460 );
or ( n270028 , n270026 , n270027 );
not ( n270029 , n258589 );
nand ( n270030 , n270029 , n251345 );
nand ( n270031 , n270028 , n270030 );
and ( n270032 , n270031 , n253377 );
not ( n270033 , n270031 );
and ( n270034 , n270033 , n253378 );
nor ( n270035 , n270032 , n270034 );
not ( n270036 , n270035 );
nand ( n270037 , n270036 , n250063 );
buf ( n270038 , n251945 );
nor ( n270039 , n246011 , n270038 );
not ( n270040 , n270039 );
nand ( n270041 , n257298 , n270038 );
nand ( n270042 , n270040 , n270041 );
and ( n270043 , n270042 , n257308 );
not ( n270044 , n270042 );
and ( n270045 , n270044 , n246017 );
nor ( n270046 , n270043 , n270045 );
not ( n270047 , n270046 );
nand ( n270048 , n270047 , n253393 );
or ( n270049 , n270037 , n270048 );
nor ( n270050 , n270047 , n53680 );
nand ( n270051 , n270050 , n270037 );
nand ( n270052 , n239240 , n31091 );
nand ( n270053 , n270049 , n270051 , n270052 );
buf ( n270054 , n270053 );
not ( n270055 , RI1754bc38_23);
or ( n270056 , n255977 , n270055 );
nand ( n270057 , n244606 , n205196 );
nand ( n270058 , n270056 , n270057 );
buf ( n270059 , n270058 );
not ( n270060 , n204830 );
not ( n270061 , n252711 );
or ( n270062 , n270060 , n270061 );
not ( n270063 , n236833 );
not ( n270064 , n257360 );
or ( n270065 , n270063 , n270064 );
not ( n270066 , n236833 );
nand ( n270067 , n270066 , n242201 );
nand ( n270068 , n270065 , n270067 );
and ( n270069 , n270068 , n255160 );
not ( n270070 , n270068 );
and ( n270071 , n270070 , n255163 );
nor ( n270072 , n270069 , n270071 );
not ( n270073 , n248012 );
nor ( n270074 , n238792 , n270073 );
not ( n270075 , n270074 );
not ( n270076 , n248012 );
nand ( n270077 , n270076 , n238792 );
nand ( n270078 , n270075 , n270077 );
not ( n270079 , n270078 );
not ( n270080 , n238895 );
and ( n270081 , n270079 , n270080 );
and ( n270082 , n270078 , n238895 );
nor ( n270083 , n270081 , n270082 );
not ( n270084 , n270083 );
nand ( n270085 , n270072 , n270084 );
not ( n270086 , n261203 );
and ( n270087 , n270085 , n270086 );
not ( n270088 , n270085 );
and ( n270089 , n270088 , n261203 );
nor ( n270090 , n270087 , n270089 );
or ( n270091 , n270090 , n258759 );
nand ( n270092 , n270062 , n270091 );
buf ( n270093 , n270092 );
or ( n270094 , n226819 , n266771 );
not ( n270095 , RI19a8e8b0_2693);
or ( n270096 , n25336 , n270095 );
nand ( n270097 , n270094 , n270096 );
buf ( n270098 , n270097 );
not ( n270099 , n263011 );
nand ( n270100 , n265885 , n270099 );
not ( n270101 , n248397 );
not ( n270102 , n43962 );
or ( n270103 , n270101 , n270102 );
not ( n270104 , n248397 );
nand ( n270105 , n270104 , n221715 );
nand ( n270106 , n270103 , n270105 );
and ( n270107 , n270106 , n255612 );
not ( n270108 , n270106 );
and ( n270109 , n270108 , n255609 );
nor ( n270110 , n270107 , n270109 );
nor ( n270111 , n270110 , n251190 );
not ( n270112 , n270111 );
or ( n270113 , n270100 , n270112 );
not ( n270114 , n270110 );
nor ( n270115 , n270114 , n55152 );
nand ( n270116 , n270115 , n270100 );
nand ( n270117 , n254798 , n28702 );
nand ( n270118 , n270113 , n270116 , n270117 );
buf ( n270119 , n270118 );
nor ( n270120 , n266046 , n55146 );
buf ( n270121 , n49578 );
not ( n270122 , n270121 );
not ( n270123 , n247187 );
or ( n270124 , n270122 , n270123 );
or ( n270125 , n247187 , n270121 );
nand ( n270126 , n270124 , n270125 );
not ( n270127 , n270126 );
not ( n270128 , n254403 );
and ( n270129 , n270127 , n270128 );
and ( n270130 , n270126 , n254403 );
nor ( n270131 , n270129 , n270130 );
not ( n270132 , n270131 );
nand ( n270133 , n270120 , n270132 , n266050 );
not ( n270134 , n266047 );
not ( n270135 , n270132 );
or ( n270136 , n270134 , n270135 );
nor ( n270137 , n266050 , n233972 );
nand ( n270138 , n270136 , n270137 );
nand ( n270139 , n50615 , n33286 );
nand ( n270140 , n270133 , n270138 , n270139 );
buf ( n270141 , n270140 );
not ( n270142 , n243348 );
not ( n270143 , n250807 );
or ( n270144 , n270142 , n270143 );
not ( n270145 , n243348 );
nand ( n270146 , n270145 , n250811 );
nand ( n270147 , n270144 , n270146 );
and ( n270148 , n270147 , n257382 );
not ( n270149 , n270147 );
buf ( n270150 , n39052 );
and ( n270151 , n270149 , n270150 );
nor ( n270152 , n270148 , n270151 );
not ( n270153 , n270152 );
nor ( n270154 , n270153 , n235050 );
not ( n270155 , n270154 );
not ( n270156 , n246156 );
not ( n270157 , n245611 );
or ( n270158 , n270156 , n270157 );
or ( n270159 , n245611 , n246156 );
nand ( n270160 , n270158 , n270159 );
not ( n270161 , n270160 );
not ( n270162 , n245615 );
and ( n270163 , n270161 , n270162 );
and ( n270164 , n270160 , n253746 );
nor ( n270165 , n270163 , n270164 );
not ( n270166 , n247003 );
not ( n270167 , n242148 );
or ( n270168 , n270166 , n270167 );
not ( n270169 , n247003 );
nand ( n270170 , n270169 , n242155 );
nand ( n270171 , n270168 , n270170 );
and ( n270172 , n270171 , n242206 );
not ( n270173 , n270171 );
and ( n270174 , n270173 , n242202 );
nor ( n270175 , n270172 , n270174 );
nor ( n270176 , n270165 , n270175 );
not ( n270177 , n270176 );
not ( n270178 , n270177 );
or ( n270179 , n270155 , n270178 );
not ( n270180 , n256292 );
not ( n270181 , n270180 );
not ( n270182 , n32208 );
and ( n270183 , n270181 , n270182 );
nor ( n270184 , n270152 , n252258 );
and ( n270185 , n270176 , n270184 );
nor ( n270186 , n270183 , n270185 );
nand ( n270187 , n270179 , n270186 );
buf ( n270188 , n270187 );
not ( n270189 , n29361 );
not ( n270190 , n233501 );
or ( n270191 , n270189 , n270190 );
nand ( n270192 , n267536 , n267521 );
not ( n270193 , n254575 );
not ( n270194 , n249462 );
or ( n270195 , n270193 , n270194 );
not ( n270196 , n254575 );
nand ( n270197 , n270196 , n249469 );
nand ( n270198 , n270195 , n270197 );
and ( n270199 , n270198 , n259704 );
not ( n270200 , n270198 );
and ( n270201 , n270200 , n259701 );
nor ( n270202 , n270199 , n270201 );
not ( n270203 , n270202 );
and ( n270204 , n270192 , n270203 );
not ( n270205 , n270192 );
and ( n270206 , n270205 , n270202 );
nor ( n270207 , n270204 , n270206 );
or ( n270208 , n270207 , n254470 );
nand ( n270209 , n270191 , n270208 );
buf ( n270210 , n270209 );
not ( n270211 , RI19acabf8_2250);
or ( n270212 , n226819 , n270211 );
not ( n270213 , RI19ac1670_2319);
or ( n270214 , n25335 , n270213 );
nand ( n270215 , n270212 , n270214 );
buf ( n270216 , n270215 );
not ( n270217 , n25512 );
not ( n270218 , n244789 );
or ( n270219 , n270217 , n270218 );
not ( n270220 , n256014 );
nand ( n270221 , n256026 , n270220 );
not ( n270222 , n264795 );
and ( n270223 , n270221 , n270222 );
not ( n270224 , n270221 );
and ( n270225 , n270224 , n264795 );
nor ( n270226 , n270223 , n270225 );
or ( n270227 , n270226 , n260861 );
nand ( n270228 , n270219 , n270227 );
buf ( n270229 , n270228 );
buf ( n270230 , n204356 );
buf ( n270231 , n45207 );
buf ( n270232 , n33466 );
xor ( n270233 , n53364 , n250370 );
xnor ( n270234 , n270233 , n250359 );
nand ( n270235 , n270234 , n259619 );
not ( n270236 , n223603 );
not ( n270237 , n36729 );
or ( n270238 , n270236 , n270237 );
not ( n270239 , n223603 );
nand ( n270240 , n270239 , n249482 );
nand ( n270241 , n270238 , n270240 );
and ( n270242 , n270241 , n249491 );
not ( n270243 , n270241 );
and ( n270244 , n270243 , n249495 );
nor ( n270245 , n270242 , n270244 );
not ( n270246 , n54254 );
not ( n270247 , n270246 );
not ( n270248 , n252185 );
or ( n270249 , n270247 , n270248 );
nand ( n270250 , n252192 , n54254 );
nand ( n270251 , n270249 , n270250 );
not ( n270252 , n270251 );
not ( n270253 , n268640 );
and ( n270254 , n270252 , n270253 );
and ( n270255 , n270251 , n268640 );
nor ( n270256 , n270254 , n270255 );
nor ( n270257 , n270245 , n270256 );
or ( n270258 , n270235 , n270257 );
nor ( n270259 , n270234 , n55152 );
nand ( n270260 , n270259 , n270257 );
nand ( n270261 , n39766 , n26095 );
nand ( n270262 , n270258 , n270260 , n270261 );
buf ( n270263 , n270262 );
not ( n270264 , n242201 );
not ( n270265 , n236840 );
and ( n270266 , n270264 , n270265 );
and ( n270267 , n242205 , n236840 );
nor ( n270268 , n270266 , n270267 );
not ( n270269 , n255163 );
and ( n270270 , n270268 , n270269 );
not ( n270271 , n270268 );
and ( n270272 , n270271 , n255163 );
nor ( n270273 , n270270 , n270272 );
not ( n270274 , n270273 );
nor ( n270275 , n268485 , n40465 );
not ( n270276 , n241024 );
not ( n270277 , n219396 );
or ( n270278 , n270276 , n270277 );
not ( n270279 , n241024 );
nand ( n270280 , n270279 , n41632 );
nand ( n270281 , n270278 , n270280 );
and ( n270282 , n270281 , n41935 );
not ( n270283 , n270281 );
and ( n270284 , n270283 , n41930 );
nor ( n270285 , n270282 , n270284 );
nand ( n270286 , n270274 , n270275 , n270285 );
nand ( n270287 , n268484 , n270285 );
nand ( n270288 , n270287 , n270273 , n222532 );
nand ( n270289 , n238638 , n204703 );
nand ( n270290 , n270286 , n270288 , n270289 );
buf ( n270291 , n270290 );
buf ( n270292 , n204594 );
buf ( n270293 , n41686 );
not ( n270294 , n41128 );
not ( n270295 , n245943 );
or ( n270296 , n270294 , n270295 );
not ( n270297 , n249597 );
not ( n270298 , n46420 );
or ( n270299 , n270297 , n270298 );
not ( n270300 , n249597 );
nand ( n270301 , n270300 , n243006 );
nand ( n270302 , n270299 , n270301 );
and ( n270303 , n270302 , n243199 );
not ( n270304 , n270302 );
and ( n270305 , n270304 , n243198 );
nor ( n270306 , n270303 , n270305 );
not ( n270307 , n270306 );
nand ( n270308 , n270307 , n250847 );
and ( n270309 , n270308 , n263145 );
not ( n270310 , n270308 );
and ( n270311 , n270310 , n250858 );
nor ( n270312 , n270309 , n270311 );
or ( n270313 , n270312 , n244217 );
nand ( n270314 , n270296 , n270313 );
buf ( n270315 , n270314 );
nand ( n270316 , n244060 , n243438 );
nand ( n270317 , n266600 , n243963 );
or ( n270318 , n270316 , n270317 );
nand ( n270319 , n270317 , n250981 );
nand ( n270320 , n49054 , n217113 );
nand ( n270321 , n270318 , n270319 , n270320 );
buf ( n270322 , n270321 );
not ( n270323 , n269352 );
not ( n270324 , n260754 );
or ( n270325 , n270323 , n270324 );
nor ( n270326 , n268283 , n31572 );
nand ( n270327 , n270325 , n270326 );
nand ( n270328 , n260754 , n268283 , n269355 );
nand ( n270329 , n244484 , n46583 );
nand ( n270330 , n270327 , n270328 , n270329 );
buf ( n270331 , n270330 );
not ( n270332 , RI19a991e8_2618);
or ( n270333 , n233507 , n270332 );
not ( n270334 , RI19a8f210_2689);
or ( n270335 , n25335 , n270334 );
nand ( n270336 , n270333 , n270335 );
buf ( n270337 , n270336 );
not ( n270338 , n53756 );
not ( n270339 , n238297 );
or ( n270340 , n270338 , n270339 );
or ( n270341 , n238297 , n53756 );
nand ( n270342 , n270340 , n270341 );
and ( n270343 , n270342 , n238409 );
not ( n270344 , n270342 );
and ( n270345 , n270344 , n238401 );
nor ( n270346 , n270343 , n270345 );
not ( n270347 , n270346 );
nor ( n270348 , n270347 , n250909 );
not ( n270349 , n270348 );
nand ( n270350 , n53147 , n53674 );
or ( n270351 , n270349 , n270350 );
not ( n270352 , n53147 );
not ( n270353 , n270346 );
or ( n270354 , n270352 , n270353 );
nor ( n270355 , n53674 , n226955 );
nand ( n270356 , n270354 , n270355 );
nand ( n270357 , n35431 , n205345 );
nand ( n270358 , n270351 , n270356 , n270357 );
buf ( n270359 , n270358 );
buf ( n270360 , n30845 );
buf ( n270361 , n32675 );
not ( n270362 , RI19a99f80_2612);
or ( n270363 , n233507 , n270362 );
not ( n270364 , RI19a8fd50_2684);
or ( n270365 , n25336 , n270364 );
nand ( n270366 , n270363 , n270365 );
buf ( n270367 , n270366 );
nand ( n270368 , n268680 , n268691 );
not ( n270369 , n237292 );
not ( n270370 , n249204 );
or ( n270371 , n270369 , n270370 );
or ( n270372 , n257658 , n237292 );
nand ( n270373 , n270371 , n270372 );
and ( n270374 , n270373 , n249207 );
not ( n270375 , n270373 );
and ( n270376 , n270375 , n249208 );
nor ( n270377 , n270374 , n270376 );
nand ( n270378 , n270377 , n241459 );
or ( n270379 , n270368 , n270378 );
nor ( n270380 , n270377 , n234021 );
nand ( n270381 , n270380 , n270368 );
nand ( n270382 , n31577 , n35759 );
nand ( n270383 , n270379 , n270381 , n270382 );
buf ( n270384 , n270383 );
nor ( n270385 , n50485 , n234021 );
buf ( n270386 , n226794 );
not ( n270387 , n270386 );
not ( n270388 , n254594 );
or ( n270389 , n270387 , n270388 );
or ( n270390 , n256460 , n270386 );
nand ( n270391 , n270389 , n270390 );
not ( n270392 , n270391 );
not ( n270393 , n254611 );
and ( n270394 , n270392 , n270393 );
and ( n270395 , n270391 , n254608 );
nor ( n270396 , n270394 , n270395 );
nand ( n270397 , n270385 , n270396 , n50607 );
not ( n270398 , n50607 );
not ( n270399 , n50485 );
not ( n270400 , n270399 );
or ( n270401 , n270398 , n270400 );
nor ( n270402 , n270396 , n234021 );
nand ( n270403 , n270401 , n270402 );
nand ( n270404 , n241068 , n29744 );
nand ( n270405 , n270397 , n270403 , n270404 );
buf ( n270406 , n270405 );
not ( n270407 , n25744 );
not ( n270408 , n51381 );
or ( n270409 , n270407 , n270408 );
not ( n270410 , n244392 );
nand ( n270411 , n249023 , n270410 );
not ( n270412 , n244349 );
and ( n270413 , n270411 , n270412 );
not ( n270414 , n270411 );
and ( n270415 , n270414 , n244349 );
nor ( n270416 , n270413 , n270415 );
or ( n270417 , n270416 , n258327 );
nand ( n270418 , n270409 , n270417 );
buf ( n270419 , n270418 );
not ( n270420 , n261850 );
nor ( n270421 , n270420 , n261840 );
not ( n270422 , n238083 );
not ( n270423 , n260383 );
or ( n270424 , n270422 , n270423 );
or ( n270425 , n260383 , n238083 );
nand ( n270426 , n270424 , n270425 );
and ( n270427 , n270426 , n247645 );
not ( n270428 , n270426 );
and ( n270429 , n270428 , n247646 );
nor ( n270430 , n270427 , n270429 );
nand ( n270431 , n270430 , n254528 );
or ( n270432 , n270421 , n270431 );
nor ( n270433 , n270430 , n238635 );
nand ( n270434 , n270433 , n270421 );
nand ( n270435 , n39767 , n25631 );
nand ( n270436 , n270432 , n270434 , n270435 );
buf ( n270437 , n270436 );
nor ( n270438 , n263757 , n226003 );
nor ( n270439 , n263751 , n244210 );
nand ( n270440 , n270438 , n270439 );
not ( n270441 , n244211 );
not ( n270442 , n263739 );
or ( n270443 , n270441 , n270442 );
nor ( n270444 , n263752 , n54208 );
nand ( n270445 , n270443 , n270444 );
nand ( n270446 , n256673 , n27973 );
nand ( n270447 , n270440 , n270445 , n270446 );
buf ( n270448 , n270447 );
nand ( n270449 , n245213 , n55147 );
not ( n270450 , n270449 );
not ( n270451 , n249353 );
not ( n270452 , n235211 );
or ( n270453 , n270451 , n270452 );
or ( n270454 , n235211 , n249353 );
nand ( n270455 , n270453 , n270454 );
and ( n270456 , n270455 , n250721 );
not ( n270457 , n270455 );
and ( n270458 , n270457 , n254375 );
nor ( n270459 , n270456 , n270458 );
nand ( n270460 , n270459 , n257792 );
not ( n270461 , n270460 );
or ( n270462 , n270450 , n270461 );
nand ( n270463 , n270462 , n245192 );
nor ( n270464 , n270459 , n236795 );
nor ( n270465 , n245213 , n245192 );
and ( n270466 , n270464 , n270465 );
and ( n270467 , n39766 , n42505 );
nor ( n270468 , n270466 , n270467 );
nand ( n270469 , n270463 , n270468 );
buf ( n270470 , n270469 );
not ( n270471 , n34637 );
not ( n270472 , n245943 );
or ( n270473 , n270471 , n270472 );
not ( n270474 , n269032 );
nand ( n270475 , n270474 , n267024 );
not ( n270476 , n267034 );
and ( n270477 , n270475 , n270476 );
not ( n270478 , n270475 );
and ( n270479 , n270478 , n267034 );
nor ( n270480 , n270477 , n270479 );
or ( n270481 , n270480 , n258327 );
nand ( n270482 , n270473 , n270481 );
buf ( n270483 , n270482 );
nand ( n270484 , n263430 , n263442 );
not ( n270485 , n244560 );
not ( n270486 , n239705 );
or ( n270487 , n270485 , n270486 );
not ( n270488 , n244560 );
nand ( n270489 , n270488 , n239715 );
nand ( n270490 , n270487 , n270489 );
and ( n270491 , n270490 , n239775 );
not ( n270492 , n270490 );
and ( n270493 , n270492 , n239776 );
nor ( n270494 , n270491 , n270493 );
not ( n270495 , n270494 );
nor ( n270496 , n270495 , n234021 );
not ( n270497 , n270496 );
or ( n270498 , n270484 , n270497 );
nor ( n270499 , n270494 , n252358 );
nand ( n270500 , n270484 , n270499 );
nand ( n270501 , n246460 , n34496 );
nand ( n270502 , n270498 , n270500 , n270501 );
buf ( n270503 , n270502 );
and ( n270504 , n27883 , n204521 );
buf ( n270505 , n270504 );
not ( n270506 , RI19ac4910_2295);
or ( n270507 , n25328 , n270506 );
not ( n270508 , RI19abc378_2366);
or ( n270509 , n25335 , n270508 );
nand ( n270510 , n270507 , n270509 );
buf ( n270511 , n270510 );
or ( n270512 , n25328 , n252208 );
or ( n270513 , n25335 , n255711 );
nand ( n270514 , n270512 , n270513 );
buf ( n270515 , n270514 );
not ( n270516 , n39694 );
not ( n270517 , n257764 );
or ( n270518 , n270516 , n270517 );
not ( n270519 , n255497 );
not ( n270520 , n246780 );
not ( n270521 , n270520 );
not ( n270522 , n249927 );
or ( n270523 , n270521 , n270522 );
nand ( n270524 , n255493 , n246780 );
nand ( n270525 , n270523 , n270524 );
not ( n270526 , n270525 );
or ( n270527 , n270519 , n270526 );
or ( n270528 , n270525 , n255497 );
nand ( n270529 , n270527 , n270528 );
nand ( n270530 , n263934 , n270529 );
and ( n270531 , n270530 , n266976 );
not ( n270532 , n270530 );
and ( n270533 , n270532 , n263926 );
nor ( n270534 , n270531 , n270533 );
or ( n270535 , n270534 , n258179 );
nand ( n270536 , n270518 , n270535 );
buf ( n270537 , n270536 );
not ( n270538 , n253063 );
not ( n270539 , n270538 );
not ( n270540 , n244704 );
or ( n270541 , n270539 , n270540 );
not ( n270542 , n270538 );
nand ( n270543 , n270542 , n244711 );
nand ( n270544 , n270541 , n270543 );
and ( n270545 , n270544 , n244778 );
not ( n270546 , n270544 );
and ( n270547 , n270546 , n244769 );
nor ( n270548 , n270545 , n270547 );
nand ( n270549 , n254275 , n238269 );
not ( n270550 , n270549 );
nor ( n270551 , n254275 , n238269 );
nor ( n270552 , n270550 , n270551 );
not ( n270553 , n270552 );
not ( n270554 , n259160 );
and ( n270555 , n270553 , n270554 );
and ( n270556 , n270552 , n259160 );
nor ( n270557 , n270555 , n270556 );
not ( n270558 , n270557 );
nor ( n270559 , n270548 , n270558 );
or ( n270560 , n257888 , n270559 );
nor ( n270561 , n257887 , n38637 );
nand ( n270562 , n270561 , n270559 );
nand ( n270563 , n41945 , n35010 );
nand ( n270564 , n270560 , n270562 , n270563 );
buf ( n270565 , n270564 );
not ( n270566 , n205026 );
not ( n270567 , n245702 );
or ( n270568 , n270566 , n270567 );
not ( n270569 , n237914 );
not ( n270570 , n246767 );
or ( n270571 , n270569 , n270570 );
not ( n270572 , n237914 );
nand ( n270573 , n270572 , n246759 );
nand ( n270574 , n270571 , n270573 );
and ( n270575 , n270574 , n254010 );
not ( n270576 , n270574 );
and ( n270577 , n270576 , n254006 );
nor ( n270578 , n270575 , n270577 );
not ( n270579 , n270578 );
not ( n270580 , n229805 );
not ( n270581 , n236267 );
or ( n270582 , n270580 , n270581 );
not ( n270583 , n229805 );
nand ( n270584 , n270583 , n245210 );
nand ( n270585 , n270582 , n270584 );
not ( n270586 , n251181 );
and ( n270587 , n270585 , n270586 );
not ( n270588 , n270585 );
and ( n270589 , n270588 , n222301 );
nor ( n270590 , n270587 , n270589 );
not ( n270591 , n270590 );
nand ( n270592 , n270579 , n270591 );
not ( n270593 , n48667 );
not ( n270594 , n234420 );
or ( n270595 , n270593 , n270594 );
not ( n270596 , n48667 );
nand ( n270597 , n270596 , n239119 );
nand ( n270598 , n270595 , n270597 );
and ( n270599 , n270598 , n239229 );
not ( n270600 , n270598 );
and ( n270601 , n270600 , n239221 );
nor ( n270602 , n270599 , n270601 );
and ( n270603 , n270592 , n270602 );
not ( n270604 , n270592 );
not ( n270605 , n270602 );
and ( n270606 , n270604 , n270605 );
nor ( n270607 , n270603 , n270606 );
or ( n270608 , n270607 , n245938 );
nand ( n270609 , n270568 , n270608 );
buf ( n270610 , n270609 );
not ( n270611 , RI19ac21b0_2313);
or ( n270612 , n25328 , n270611 );
or ( n270613 , n25336 , n264637 );
nand ( n270614 , n270612 , n270613 );
buf ( n270615 , n270614 );
buf ( n270616 , n35341 );
buf ( n270617 , n31466 );
buf ( n270618 , n34804 );
buf ( n270619 , n29867 );
nor ( n270620 , n269702 , n234021 );
not ( n270621 , n270620 );
nand ( n270622 , n256883 , n269703 );
or ( n270623 , n270621 , n270622 );
not ( n270624 , n269703 );
not ( n270625 , n269702 );
not ( n270626 , n270625 );
or ( n270627 , n270624 , n270626 );
nor ( n270628 , n256883 , n31572 );
nand ( n270629 , n270627 , n270628 );
nand ( n270630 , n238638 , n29994 );
nand ( n270631 , n270623 , n270629 , n270630 );
buf ( n270632 , n270631 );
not ( n270633 , RI19a93518_2659);
or ( n270634 , n226819 , n270633 );
or ( n270635 , n25335 , n257406 );
nand ( n270636 , n270634 , n270635 );
buf ( n270637 , n270636 );
buf ( n270638 , n29157 );
buf ( n270639 , n36927 );
buf ( n270640 , n28900 );
nand ( n270641 , n255679 , n256665 );
or ( n270642 , n259439 , n270641 );
not ( n270643 , n256665 );
not ( n270644 , n256651 );
or ( n270645 , n270643 , n270644 );
nor ( n270646 , n255679 , n33253 );
nand ( n270647 , n270645 , n270646 );
nand ( n270648 , n31576 , n39336 );
nand ( n270649 , n270642 , n270647 , n270648 );
buf ( n270650 , n270649 );
not ( n270651 , n36825 );
not ( n270652 , n245943 );
or ( n270653 , n270651 , n270652 );
not ( n270654 , n53297 );
not ( n270655 , n250359 );
or ( n270656 , n270654 , n270655 );
not ( n270657 , n53297 );
nand ( n270658 , n270657 , n250366 );
nand ( n270659 , n270656 , n270658 );
and ( n270660 , n270659 , n250374 );
not ( n270661 , n270659 );
and ( n270662 , n270661 , n250371 );
nor ( n270663 , n270660 , n270662 );
not ( n270664 , n270663 );
nand ( n270665 , n270664 , n263418 );
and ( n270666 , n270665 , n263430 );
not ( n270667 , n270665 );
and ( n270668 , n270667 , n263431 );
nor ( n270669 , n270666 , n270668 );
or ( n270670 , n270669 , n258327 );
nand ( n270671 , n270653 , n270670 );
buf ( n270672 , n270671 );
buf ( n270673 , n30526 );
not ( n270674 , n246860 );
not ( n270675 , n242852 );
or ( n270676 , n270674 , n270675 );
or ( n270677 , n242860 , n246860 );
nand ( n270678 , n270676 , n270677 );
and ( n270679 , n270678 , n208725 );
not ( n270680 , n270678 );
and ( n270681 , n270680 , n242866 );
nor ( n270682 , n270679 , n270681 );
not ( n270683 , n270682 );
not ( n270684 , n241152 );
not ( n270685 , n235728 );
or ( n270686 , n270684 , n270685 );
not ( n270687 , n241152 );
nand ( n270688 , n270687 , n235718 );
nand ( n270689 , n270686 , n270688 );
and ( n270690 , n270689 , n260711 );
not ( n270691 , n270689 );
and ( n270692 , n270691 , n236504 );
nor ( n270693 , n270690 , n270692 );
not ( n270694 , n270693 );
or ( n270695 , n270683 , n270694 );
not ( n270696 , n227538 );
not ( n270697 , n259737 );
or ( n270698 , n270696 , n270697 );
or ( n270699 , n243415 , n227538 );
nand ( n270700 , n270698 , n270699 );
not ( n270701 , n270700 );
not ( n270702 , n259744 );
and ( n270703 , n270701 , n270702 );
and ( n270704 , n270700 , n259744 );
nor ( n270705 , n270703 , n270704 );
nor ( n270706 , n270705 , n37724 );
nand ( n270707 , n270695 , n270706 );
not ( n270708 , n270705 );
not ( n270709 , n270708 );
not ( n270710 , n270682 );
nor ( n270711 , n270710 , n241065 );
nand ( n270712 , n270709 , n270693 , n270711 );
nand ( n270713 , n238114 , n31293 );
nand ( n270714 , n270707 , n270712 , n270713 );
buf ( n270715 , n270714 );
not ( n270716 , RI19aba050_2380);
or ( n270717 , n25328 , n270716 );
or ( n270718 , n25335 , n267743 );
nand ( n270719 , n270717 , n270718 );
buf ( n270720 , n270719 );
nand ( n270721 , n242685 , n222532 );
not ( n270722 , n245555 );
not ( n270723 , n270722 );
not ( n270724 , n232899 );
or ( n270725 , n270723 , n270724 );
not ( n270726 , n270722 );
nand ( n270727 , n270726 , n55135 );
nand ( n270728 , n270725 , n270727 );
and ( n270729 , n270728 , n37709 );
not ( n270730 , n270728 );
and ( n270731 , n270730 , n37715 );
nor ( n270732 , n270729 , n270731 );
not ( n270733 , n270732 );
nand ( n270734 , n270733 , n242703 );
or ( n270735 , n270721 , n270734 );
not ( n270736 , n242703 );
not ( n270737 , n242685 );
or ( n270738 , n270736 , n270737 );
nor ( n270739 , n270733 , n265700 );
nand ( n270740 , n270738 , n270739 );
nand ( n270741 , n250916 , n25817 );
nand ( n270742 , n270735 , n270740 , n270741 );
buf ( n270743 , n270742 );
or ( n270744 , n233507 , n268838 );
or ( n270745 , n226822 , n265912 );
nand ( n270746 , n270744 , n270745 );
buf ( n270747 , n270746 );
not ( n270748 , n205001 );
not ( n270749 , n262000 );
or ( n270750 , n270748 , n270749 );
not ( n270751 , n251936 );
not ( n270752 , n257298 );
or ( n270753 , n270751 , n270752 );
or ( n270754 , n251689 , n251936 );
nand ( n270755 , n270753 , n270754 );
not ( n270756 , n270755 );
not ( n270757 , n246017 );
and ( n270758 , n270756 , n270757 );
and ( n270759 , n270755 , n246017 );
nor ( n270760 , n270758 , n270759 );
not ( n270761 , n247781 );
not ( n270762 , n232514 );
or ( n270763 , n270761 , n270762 );
not ( n270764 , n247781 );
nand ( n270765 , n270764 , n232520 );
nand ( n270766 , n270763 , n270765 );
and ( n270767 , n270766 , n247269 );
not ( n270768 , n270766 );
and ( n270769 , n270768 , n232299 );
nor ( n270770 , n270767 , n270769 );
nand ( n270771 , n270760 , n270770 );
not ( n270772 , n270771 );
not ( n270773 , n238445 );
not ( n270774 , n228918 );
or ( n270775 , n270773 , n270774 );
not ( n270776 , n238445 );
nand ( n270777 , n270776 , n51167 );
nand ( n270778 , n270775 , n270777 );
and ( n270779 , n270778 , n51269 );
not ( n270780 , n270778 );
and ( n270781 , n270780 , n51272 );
nor ( n270782 , n270779 , n270781 );
not ( n270783 , n270782 );
not ( n270784 , n270783 );
and ( n270785 , n270772 , n270784 );
and ( n270786 , n270771 , n270783 );
nor ( n270787 , n270785 , n270786 );
or ( n270788 , n270787 , n31572 );
nand ( n270789 , n270750 , n270788 );
buf ( n270790 , n270789 );
or ( n270791 , n25328 , n269488 );
not ( n270792 , RI19ac89c0_2265);
or ( n270793 , n25335 , n270792 );
nand ( n270794 , n270791 , n270793 );
buf ( n270795 , n270794 );
not ( n270796 , n248429 );
not ( n270797 , n43962 );
or ( n270798 , n270796 , n270797 );
not ( n270799 , n248429 );
nand ( n270800 , n270799 , n221715 );
nand ( n270801 , n270798 , n270800 );
and ( n270802 , n270801 , n255612 );
not ( n270803 , n270801 );
and ( n270804 , n270803 , n255609 );
nor ( n270805 , n270802 , n270804 );
not ( n270806 , n270805 );
nor ( n270807 , n270806 , n49959 );
not ( n270808 , n270807 );
not ( n270809 , n50943 );
nand ( n270810 , n51274 , n270809 );
or ( n270811 , n270808 , n270810 );
not ( n270812 , n270809 );
not ( n270813 , n270805 );
or ( n270814 , n270812 , n270813 );
nor ( n270815 , n51274 , n31572 );
nand ( n270816 , n270814 , n270815 );
nand ( n270817 , n245701 , n33449 );
nand ( n270818 , n270811 , n270816 , n270817 );
buf ( n270819 , n270818 );
not ( n270820 , n244918 );
not ( n270821 , n34439 );
or ( n270822 , n270820 , n270821 );
not ( n270823 , n244918 );
nand ( n270824 , n270823 , n34448 );
nand ( n270825 , n270822 , n270824 );
and ( n270826 , n270825 , n33709 );
not ( n270827 , n270825 );
and ( n270828 , n270827 , n235042 );
nor ( n270829 , n270826 , n270828 );
not ( n270830 , n270829 );
not ( n270831 , n255962 );
or ( n270832 , n270830 , n270831 );
nand ( n270833 , n270832 , n248684 );
not ( n270834 , n270829 );
nor ( n270835 , n270834 , n254226 );
nand ( n270836 , n270835 , n255962 , n248683 );
nand ( n270837 , n253486 , n35891 );
nand ( n270838 , n270833 , n270836 , n270837 );
buf ( n270839 , n270838 );
nand ( n270840 , n254389 , n250111 );
nand ( n270841 , n268986 , n254377 );
or ( n270842 , n270840 , n270841 );
not ( n270843 , n268986 );
not ( n270844 , n254389 );
or ( n270845 , n270843 , n270844 );
nor ( n270846 , n254377 , n46425 );
nand ( n270847 , n270845 , n270846 );
nand ( n270848 , n31577 , n29319 );
nand ( n270849 , n270842 , n270847 , n270848 );
buf ( n270850 , n270849 );
not ( n270851 , n239444 );
not ( n270852 , n260112 );
or ( n270853 , n270851 , n270852 );
not ( n270854 , n239444 );
nand ( n270855 , n270854 , n260122 );
nand ( n270856 , n270853 , n270855 );
not ( n270857 , n270856 );
not ( n270858 , n260125 );
and ( n270859 , n270857 , n270858 );
and ( n270860 , n270856 , n260125 );
nor ( n270861 , n270859 , n270860 );
nor ( n270862 , n270861 , n252358 );
nand ( n270863 , n270862 , n265770 , n265783 );
not ( n270864 , n270861 );
not ( n270865 , n270864 );
not ( n270866 , n265770 );
or ( n270867 , n270865 , n270866 );
nor ( n270868 , n265783 , n234440 );
nand ( n270869 , n270867 , n270868 );
nand ( n270870 , n255116 , n28714 );
nand ( n270871 , n270863 , n270869 , n270870 );
buf ( n270872 , n270871 );
buf ( n270873 , n32203 );
not ( n270874 , RI19a9c848_2594);
or ( n270875 , n25328 , n270874 );
not ( n270876 , RI19a92708_2665);
or ( n270877 , n25335 , n270876 );
nand ( n270878 , n270875 , n270877 );
buf ( n270879 , n270878 );
buf ( n270880 , n40045 );
nor ( n270881 , n264602 , n266426 );
nand ( n270882 , n266437 , n270881 );
not ( n270883 , n266426 );
not ( n270884 , n270883 );
not ( n270885 , n266440 );
or ( n270886 , n270884 , n270885 );
nand ( n270887 , n270886 , n264604 );
nand ( n270888 , n49054 , n29875 );
nand ( n270889 , n270882 , n270887 , n270888 );
buf ( n270890 , n270889 );
not ( n270891 , n251610 );
not ( n270892 , n55889 );
or ( n270893 , n270891 , n270892 );
not ( n270894 , n251610 );
nand ( n270895 , n270894 , n233660 );
nand ( n270896 , n270893 , n270895 );
and ( n270897 , n270896 , n233805 );
not ( n270898 , n270896 );
and ( n270899 , n270898 , n269239 );
nor ( n270900 , n270897 , n270899 );
not ( n270901 , n268765 );
nand ( n270902 , n270900 , n270901 );
not ( n270903 , n38214 );
not ( n270904 , n50027 );
or ( n270905 , n270903 , n270904 );
not ( n270906 , n38214 );
nand ( n270907 , n270906 , n227795 );
nand ( n270908 , n270905 , n270907 );
and ( n270909 , n270908 , n234522 );
not ( n270910 , n270908 );
and ( n270911 , n270910 , n234514 );
nor ( n270912 , n270909 , n270911 );
nor ( n270913 , n270912 , n55152 );
not ( n270914 , n270913 );
or ( n270915 , n270902 , n270914 );
not ( n270916 , n270912 );
nor ( n270917 , n270916 , n251462 );
nand ( n270918 , n270917 , n270902 );
nand ( n270919 , n241068 , n40027 );
nand ( n270920 , n270915 , n270918 , n270919 );
buf ( n270921 , n270920 );
not ( n270922 , RI19a23c18_2790);
or ( n270923 , n25328 , n270922 );
or ( n270924 , n25335 , n266364 );
nand ( n270925 , n270923 , n270924 );
buf ( n270926 , n270925 );
not ( n270927 , RI19a9e468_2582);
or ( n270928 , n25328 , n270927 );
not ( n270929 , RI19a94238_2653);
or ( n270930 , n226822 , n270929 );
nand ( n270931 , n270928 , n270930 );
buf ( n270932 , n270931 );
not ( n270933 , RI19ab52f8_2415);
or ( n270934 , n233507 , n270933 );
not ( n270935 , RI19aab5f0_2486);
or ( n270936 , n25335 , n270935 );
nand ( n270937 , n270934 , n270936 );
buf ( n270938 , n270937 );
nor ( n270939 , n270829 , n243204 );
nand ( n270940 , n270939 , n248694 , n248683 );
nand ( n270941 , n248683 , n270834 );
nand ( n270942 , n270941 , n255949 , n40466 );
nand ( n270943 , n237714 , n208577 );
nand ( n270944 , n270940 , n270942 , n270943 );
buf ( n270945 , n270944 );
not ( n270946 , RI19a94490_2652);
or ( n270947 , n25328 , n270946 );
not ( n270948 , RI19a8a530_2722);
or ( n270949 , n25335 , n270948 );
nand ( n270950 , n270947 , n270949 );
buf ( n270951 , n270950 );
buf ( n270952 , RI19a240c8_2788);
not ( n270953 , n270952 );
not ( n270954 , n257347 );
or ( n270955 , n270953 , n270954 );
nand ( n270956 , n257351 , n262039 );
nand ( n270957 , n270955 , n270956 );
buf ( n270958 , n270957 );
buf ( n270959 , n36796 );
buf ( n270960 , n26282 );
buf ( n270961 , n39476 );
buf ( n270962 , n30993 );
not ( n270963 , n205649 );
nor ( n270964 , n261662 , n270963 );
nand ( n270965 , n270964 , n249497 );
not ( n270966 , n249473 );
not ( n270967 , n261662 );
and ( n270968 , n270966 , n270967 );
and ( n270969 , n50615 , n35057 );
nor ( n270970 , n270968 , n270969 );
nand ( n270971 , n266871 , n249498 , n261662 );
nand ( n270972 , n270965 , n270970 , n270971 );
buf ( n270973 , n270972 );
not ( n270974 , n264513 );
not ( n270975 , n244443 );
not ( n270976 , n247551 );
or ( n270977 , n270975 , n270976 );
not ( n270978 , n244443 );
nand ( n270979 , n270978 , n247561 );
nand ( n270980 , n270977 , n270979 );
not ( n270981 , n255006 );
and ( n270982 , n270980 , n270981 );
not ( n270983 , n270980 );
and ( n270984 , n270983 , n255006 );
nor ( n270985 , n270982 , n270984 );
not ( n270986 , n270985 );
nand ( n270987 , n270974 , n270986 );
or ( n270988 , n264535 , n270987 );
not ( n270989 , n264534 );
not ( n270990 , n270974 );
or ( n270991 , n270989 , n270990 );
nor ( n270992 , n270986 , n264469 );
nand ( n270993 , n270991 , n270992 );
nand ( n270994 , n35431 , n36779 );
nand ( n270995 , n270988 , n270993 , n270994 );
buf ( n270996 , n270995 );
or ( n270997 , n25328 , n255972 );
or ( n270998 , n25335 , n256677 );
nand ( n270999 , n270997 , n270998 );
buf ( n271000 , n270999 );
buf ( n271001 , n253654 );
not ( n271002 , n271001 );
not ( n271003 , n246653 );
or ( n271004 , n271002 , n271003 );
or ( n271005 , n246653 , n271001 );
nand ( n271006 , n271004 , n271005 );
not ( n271007 , n271006 );
not ( n271008 , n262526 );
and ( n271009 , n271007 , n271008 );
and ( n271010 , n271006 , n262526 );
nor ( n271011 , n271009 , n271010 );
nand ( n271012 , n271011 , n246177 );
not ( n271013 , n252177 );
not ( n271014 , n220460 );
or ( n271015 , n271013 , n271014 );
not ( n271016 , n252177 );
nand ( n271017 , n271016 , n220467 );
nand ( n271018 , n271015 , n271017 );
and ( n271019 , n271018 , n43006 );
not ( n271020 , n271018 );
and ( n271021 , n271020 , n43011 );
nor ( n271022 , n271019 , n271021 );
not ( n271023 , n271022 );
nand ( n271024 , n271023 , n246451 );
or ( n271025 , n271012 , n271024 );
not ( n271026 , n246451 );
not ( n271027 , n271011 );
or ( n271028 , n271026 , n271027 );
nor ( n271029 , n271023 , n35427 );
nand ( n271030 , n271028 , n271029 );
nand ( n271031 , n256673 , n31180 );
nand ( n271032 , n271025 , n271030 , n271031 );
buf ( n271033 , n271032 );
not ( n271034 , RI1754c070_14);
or ( n271035 , n51369 , n271034 );
nand ( n271036 , n258185 , n33078 );
nand ( n271037 , n271035 , n271036 );
buf ( n271038 , n271037 );
not ( n271039 , RI19a86c00_2747);
or ( n271040 , n25328 , n271039 );
or ( n271041 , n25335 , n269661 );
nand ( n271042 , n271040 , n271041 );
buf ( n271043 , n271042 );
not ( n271044 , n49823 );
not ( n271045 , n245872 );
or ( n271046 , n271044 , n271045 );
or ( n271047 , n245872 , n49823 );
nand ( n271048 , n271046 , n271047 );
and ( n271049 , n271048 , n245930 );
not ( n271050 , n271048 );
and ( n271051 , n271050 , n245920 );
nor ( n271052 , n271049 , n271051 );
not ( n271053 , n271052 );
nor ( n271054 , n271053 , n250431 );
not ( n271055 , n271054 );
not ( n271056 , n241914 );
not ( n271057 , n259905 );
or ( n271058 , n271056 , n271057 );
not ( n271059 , n241914 );
nand ( n271060 , n271059 , n237590 );
nand ( n271061 , n271058 , n271060 );
and ( n271062 , n271061 , n259578 );
not ( n271063 , n271061 );
and ( n271064 , n271063 , n259575 );
nor ( n271065 , n271062 , n271064 );
not ( n271066 , n235270 );
not ( n271067 , n271066 );
not ( n271068 , n246448 );
or ( n271069 , n271067 , n271068 );
not ( n271070 , n271066 );
nand ( n271071 , n271070 , n246439 );
nand ( n271072 , n271069 , n271071 );
and ( n271073 , n271072 , n250021 );
not ( n271074 , n271072 );
and ( n271075 , n271074 , n250030 );
nor ( n271076 , n271073 , n271075 );
nand ( n271077 , n271065 , n271076 );
or ( n271078 , n271055 , n271077 );
not ( n271079 , n271052 );
not ( n271080 , n271065 );
or ( n271081 , n271079 , n271080 );
nor ( n271082 , n271076 , n52445 );
nand ( n271083 , n271081 , n271082 );
nand ( n271084 , n35431 , n29984 );
nand ( n271085 , n271078 , n271083 , n271084 );
buf ( n271086 , n271085 );
not ( n271087 , RI19aa1f00_2553);
or ( n271088 , n25328 , n271087 );
or ( n271089 , n226822 , n258189 );
nand ( n271090 , n271088 , n271089 );
buf ( n271091 , n271090 );
not ( n271092 , n29052 );
not ( n271093 , n251465 );
or ( n271094 , n271092 , n271093 );
not ( n271095 , n264569 );
nand ( n271096 , n271095 , n241062 );
and ( n271097 , n271096 , n240998 );
not ( n271098 , n271096 );
not ( n271099 , n240998 );
and ( n271100 , n271098 , n271099 );
nor ( n271101 , n271097 , n271100 );
or ( n271102 , n271101 , n237358 );
nand ( n271103 , n271094 , n271102 );
buf ( n271104 , n271103 );
not ( n271105 , n251513 );
not ( n271106 , n46870 );
not ( n271107 , n250019 );
or ( n271108 , n271106 , n271107 );
not ( n271109 , n46870 );
nand ( n271110 , n271109 , n250028 );
nand ( n271111 , n271108 , n271110 );
xnor ( n271112 , n271111 , n252831 );
not ( n271113 , n271112 );
nand ( n271114 , n271113 , n251536 );
or ( n271115 , n271105 , n271114 );
nor ( n271116 , n251552 , n255896 );
nand ( n271117 , n271116 , n271114 );
nand ( n271118 , n251717 , n34203 );
nand ( n271119 , n271115 , n271117 , n271118 );
buf ( n271120 , n271119 );
not ( n271121 , n40529 );
not ( n271122 , n39766 );
or ( n271123 , n271121 , n271122 );
not ( n271124 , n254173 );
not ( n271125 , n235501 );
not ( n271126 , n248135 );
or ( n271127 , n271125 , n271126 );
not ( n271128 , n235501 );
nand ( n271129 , n271128 , n248143 );
nand ( n271130 , n271127 , n271129 );
and ( n271131 , n271130 , n248146 );
not ( n271132 , n271130 );
and ( n271133 , n271132 , n248149 );
nor ( n271134 , n271131 , n271133 );
nand ( n271135 , n271124 , n271134 );
and ( n271136 , n271135 , n265481 );
not ( n271137 , n271135 );
and ( n271138 , n271137 , n265478 );
nor ( n271139 , n271136 , n271138 );
or ( n271140 , n271139 , n237358 );
nand ( n271141 , n271123 , n271140 );
buf ( n271142 , n271141 );
or ( n271143 , n25328 , n267845 );
not ( n271144 , RI19a98018_2626);
or ( n271145 , n226822 , n271144 );
nand ( n271146 , n271143 , n271145 );
buf ( n271147 , n271146 );
not ( n271148 , n41035 );
not ( n271149 , n54273 );
or ( n271150 , n271148 , n271149 );
or ( n271151 , n54273 , n41035 );
nand ( n271152 , n271150 , n271151 );
and ( n271153 , n271152 , n255324 );
not ( n271154 , n271152 );
and ( n271155 , n271154 , n255321 );
nor ( n271156 , n271153 , n271155 );
nand ( n271157 , n271156 , n257792 );
not ( n271158 , n249343 );
not ( n271159 , n235202 );
or ( n271160 , n271158 , n271159 );
not ( n271161 , n249343 );
nand ( n271162 , n271161 , n235211 );
nand ( n271163 , n271160 , n271162 );
and ( n271164 , n271163 , n254375 );
not ( n271165 , n271163 );
and ( n271166 , n271165 , n250721 );
nor ( n271167 , n271164 , n271166 );
not ( n271168 , n248627 );
not ( n271169 , n251845 );
or ( n271170 , n271168 , n271169 );
not ( n271171 , n248627 );
nand ( n271172 , n271171 , n251855 );
nand ( n271173 , n271170 , n271172 );
and ( n271174 , n271173 , n260966 );
not ( n271175 , n271173 );
and ( n271176 , n271175 , n267340 );
nor ( n271177 , n271174 , n271176 );
not ( n271178 , n271177 );
nand ( n271179 , n271167 , n271178 );
or ( n271180 , n271157 , n271179 );
not ( n271181 , n271167 );
not ( n271182 , n271156 );
or ( n271183 , n271181 , n271182 );
nor ( n271184 , n271178 , n251862 );
nand ( n271185 , n271183 , n271184 );
nand ( n271186 , n251712 , n25520 );
nand ( n271187 , n271180 , n271185 , n271186 );
buf ( n271188 , n271187 );
not ( n271189 , RI19abad70_2375);
or ( n271190 , n25328 , n271189 );
or ( n271191 , n25336 , n266716 );
nand ( n271192 , n271190 , n271191 );
buf ( n271193 , n271192 );
not ( n271194 , n246276 );
not ( n271195 , n239607 );
or ( n271196 , n271194 , n271195 );
or ( n271197 , n239610 , n246276 );
nand ( n271198 , n271196 , n271197 );
and ( n271199 , n271198 , n244127 );
not ( n271200 , n271198 );
and ( n271201 , n271200 , n239654 );
nor ( n271202 , n271199 , n271201 );
not ( n271203 , n271202 );
nand ( n271204 , n271203 , n262340 );
or ( n271205 , n262003 , n271204 );
not ( n271206 , n261974 );
nand ( n271207 , n271206 , n271204 );
nand ( n271208 , n245702 , n209468 );
nand ( n271209 , n271205 , n271207 , n271208 );
buf ( n271210 , n271209 );
not ( n271211 , n31421 );
not ( n271212 , n39766 );
or ( n271213 , n271211 , n271212 );
not ( n271214 , n249240 );
not ( n271215 , n244889 );
or ( n271216 , n271214 , n271215 );
not ( n271217 , n249240 );
nand ( n271218 , n271217 , n244899 );
nand ( n271219 , n271216 , n271218 );
and ( n271220 , n271219 , n244940 );
not ( n271221 , n271219 );
and ( n271222 , n271221 , n244955 );
nor ( n271223 , n271220 , n271222 );
not ( n271224 , n271223 );
nand ( n271225 , n271224 , n259958 );
not ( n271226 , n259970 );
and ( n271227 , n271225 , n271226 );
not ( n271228 , n271225 );
and ( n271229 , n271228 , n259970 );
nor ( n271230 , n271227 , n271229 );
or ( n271231 , n271230 , n253358 );
nand ( n271232 , n271213 , n271231 );
buf ( n271233 , n271232 );
not ( n271234 , n236261 );
not ( n271235 , n241255 );
or ( n271236 , n271234 , n271235 );
or ( n271237 , n241255 , n236261 );
nand ( n271238 , n271236 , n271237 );
and ( n271239 , n271238 , n241370 );
not ( n271240 , n271238 );
and ( n271241 , n271240 , n241361 );
nor ( n271242 , n271239 , n271241 );
not ( n271243 , n268251 );
nand ( n271244 , n271242 , n271243 );
or ( n271245 , n271244 , n268229 );
nor ( n271246 , n268228 , n237384 );
nand ( n271247 , n271244 , n271246 );
nand ( n271248 , n254798 , n36488 );
nand ( n271249 , n271245 , n271247 , n271248 );
buf ( n271250 , n271249 );
not ( n271251 , RI1754b3c8_41);
or ( n271252 , n249128 , n271251 );
nand ( n271253 , n249131 , n32166 );
nand ( n271254 , n271252 , n271253 );
buf ( n271255 , n271254 );
not ( n271256 , n30388 );
not ( n271257 , n233501 );
or ( n271258 , n271256 , n271257 );
not ( n271259 , n250815 );
nand ( n271260 , n253900 , n271259 );
and ( n271261 , n271260 , n264293 );
not ( n271262 , n271260 );
and ( n271263 , n271262 , n257802 );
nor ( n271264 , n271261 , n271263 );
or ( n271265 , n271264 , n258280 );
nand ( n271266 , n271258 , n271265 );
buf ( n271267 , n271266 );
buf ( n271268 , n40508 );
nand ( n271269 , n268530 , n268120 );
not ( n271270 , n268108 );
or ( n271271 , n271269 , n271270 );
nand ( n271272 , n244958 , n271269 );
nand ( n271273 , n39767 , n204463 );
nand ( n271274 , n271271 , n271272 , n271273 );
buf ( n271275 , n271274 );
not ( n271276 , n30125 );
not ( n271277 , n31577 );
or ( n271278 , n271276 , n271277 );
nand ( n271279 , n269100 , n257214 );
and ( n271280 , n271279 , n269088 );
not ( n271281 , n271279 );
and ( n271282 , n271281 , n269089 );
nor ( n271283 , n271280 , n271282 );
or ( n271284 , n271283 , n258328 );
nand ( n271285 , n271278 , n271284 );
buf ( n271286 , n271285 );
buf ( n271287 , n28587 );
not ( n271288 , n255073 );
not ( n271289 , n34622 );
not ( n271290 , n244373 );
or ( n271291 , n271289 , n271290 );
not ( n271292 , n34622 );
nand ( n271293 , n271292 , n255080 );
nand ( n271294 , n271291 , n271293 );
not ( n271295 , n271294 );
or ( n271296 , n271288 , n271295 );
or ( n271297 , n271294 , n255089 );
nand ( n271298 , n271296 , n271297 );
nor ( n271299 , n238217 , n271298 );
or ( n271300 , n259784 , n271299 );
nor ( n271301 , n271298 , n38637 );
nand ( n271302 , n259781 , n271301 , n238218 );
nand ( n271303 , n251465 , n26438 );
nand ( n271304 , n271300 , n271302 , n271303 );
buf ( n271305 , n271304 );
not ( n271306 , n263588 );
nand ( n271307 , n271306 , n262983 );
or ( n271308 , n271307 , n243234 );
nand ( n271309 , n271307 , n243270 );
nand ( n271310 , n31577 , n38085 );
nand ( n271311 , n271308 , n271309 , n271310 );
buf ( n271312 , n271311 );
not ( n271313 , RI19ac7d90_2271);
or ( n271314 , n25328 , n271313 );
or ( n271315 , n25336 , n261019 );
nand ( n271316 , n271314 , n271315 );
buf ( n271317 , n271316 );
or ( n271318 , n25328 , n264963 );
not ( n271319 , RI19a99d28_2613);
or ( n271320 , n25335 , n271319 );
nand ( n271321 , n271318 , n271320 );
buf ( n271322 , n271321 );
not ( n271323 , n34484 );
not ( n271324 , n245702 );
or ( n271325 , n271323 , n271324 );
not ( n271326 , n217329 );
not ( n271327 , n34956 );
or ( n271328 , n271326 , n271327 );
not ( n271329 , n217329 );
nand ( n271330 , n271329 , n34968 );
nand ( n271331 , n271328 , n271330 );
xor ( n271332 , n271331 , n35410 );
not ( n271333 , n250272 );
not ( n271334 , n252293 );
not ( n271335 , n243959 );
or ( n271336 , n271334 , n271335 );
nand ( n271337 , n243953 , n252290 );
nand ( n271338 , n271336 , n271337 );
not ( n271339 , n271338 );
or ( n271340 , n271333 , n271339 );
or ( n271341 , n271338 , n250272 );
nand ( n271342 , n271340 , n271341 );
nand ( n271343 , n271332 , n271342 );
not ( n271344 , n234981 );
not ( n271345 , n236993 );
or ( n271346 , n271344 , n271345 );
or ( n271347 , n236993 , n234981 );
nand ( n271348 , n271346 , n271347 );
and ( n271349 , n271348 , n254125 );
not ( n271350 , n271348 );
and ( n271351 , n271350 , n254122 );
nor ( n271352 , n271349 , n271351 );
not ( n271353 , n271352 );
and ( n271354 , n271343 , n271353 );
not ( n271355 , n271343 );
and ( n271356 , n271355 , n271352 );
nor ( n271357 , n271354 , n271356 );
or ( n271358 , n271357 , n260760 );
nand ( n271359 , n271325 , n271358 );
buf ( n271360 , n271359 );
not ( n271361 , n264483 );
nand ( n271362 , n271361 , n264496 );
not ( n271363 , n255230 );
or ( n271364 , n271362 , n271363 );
nand ( n271365 , n271362 , n255234 );
nand ( n271366 , n239240 , n31069 );
nand ( n271367 , n271364 , n271365 , n271366 );
buf ( n271368 , n271367 );
not ( n271369 , n44305 );
not ( n271370 , n234097 );
or ( n271371 , n271369 , n271370 );
not ( n271372 , n44305 );
nand ( n271373 , n271372 , n234106 );
nand ( n271374 , n271371 , n271373 );
and ( n271375 , n271374 , n249470 );
not ( n271376 , n271374 );
and ( n271377 , n271376 , n249463 );
nor ( n271378 , n271375 , n271377 );
not ( n271379 , n271378 );
not ( n271380 , n262601 );
not ( n271381 , n271380 );
or ( n271382 , n271379 , n271381 );
nor ( n271383 , n262615 , n40465 );
nand ( n271384 , n271382 , n271383 );
not ( n271385 , n271378 );
nor ( n271386 , n271385 , n256413 );
nand ( n271387 , n271386 , n271380 , n262615 );
nand ( n271388 , n245414 , n30409 );
nand ( n271389 , n271384 , n271387 , n271388 );
buf ( n271390 , n271389 );
nand ( n271391 , n260302 , n248981 );
not ( n271392 , n260318 );
not ( n271393 , n254240 );
nand ( n271394 , n271392 , n271393 );
or ( n271395 , n271391 , n271394 );
and ( n271396 , n260302 , n271393 );
nand ( n271397 , n260318 , n254227 );
nor ( n271398 , n271396 , n271397 );
not ( n271399 , n35997 );
not ( n271400 , n234024 );
nor ( n271401 , n271399 , n271400 );
nor ( n271402 , n271398 , n271401 );
nand ( n271403 , n271395 , n271402 );
buf ( n271404 , n271403 );
nand ( n271405 , n269021 , n235051 );
nand ( n271406 , n269032 , n267024 );
or ( n271407 , n271405 , n271406 );
not ( n271408 , n269032 );
not ( n271409 , n269021 );
or ( n271410 , n271408 , n271409 );
nor ( n271411 , n267024 , n234440 );
nand ( n271412 , n271410 , n271411 );
nand ( n271413 , n263819 , n31669 );
nand ( n271414 , n271407 , n271412 , n271413 );
buf ( n271415 , n271414 );
not ( n271416 , n247213 );
not ( n271417 , n251492 );
nand ( n271418 , n251481 , n271417 );
or ( n271419 , n271416 , n271418 );
not ( n271420 , n271417 );
not ( n271421 , n247216 );
or ( n271422 , n271420 , n271421 );
nor ( n271423 , n251481 , n35427 );
nand ( n271424 , n271422 , n271423 );
nand ( n271425 , n238638 , n207190 );
nand ( n271426 , n271419 , n271424 , n271425 );
buf ( n271427 , n271426 );
not ( n271428 , n253398 );
not ( n271429 , n253394 );
or ( n271430 , n271428 , n271429 );
nand ( n271431 , n271430 , n258265 );
nor ( n271432 , n253392 , n258265 );
and ( n271433 , n258281 , n271432 );
and ( n271434 , n245943 , n206940 );
nor ( n271435 , n271433 , n271434 );
nand ( n271436 , n271431 , n271435 );
buf ( n271437 , n271436 );
nand ( n271438 , n261950 , n269818 , n239111 );
not ( n271439 , n238899 );
not ( n271440 , n269818 );
or ( n271441 , n271439 , n271440 );
not ( n271442 , n205649 );
nor ( n271443 , n271442 , n239111 );
nand ( n271444 , n271441 , n271443 );
nand ( n271445 , n241378 , n38073 );
nand ( n271446 , n271438 , n271444 , n271445 );
buf ( n271447 , n271446 );
not ( n271448 , n234673 );
not ( n271449 , n271448 );
not ( n271450 , n249284 );
or ( n271451 , n271449 , n271450 );
nand ( n271452 , n249522 , n234673 );
nand ( n271453 , n271451 , n271452 );
and ( n271454 , n271453 , n249528 );
not ( n271455 , n271453 );
and ( n271456 , n271455 , n249525 );
nor ( n271457 , n271454 , n271456 );
not ( n271458 , n271457 );
nand ( n271459 , n271458 , n43969 );
buf ( n271460 , n250869 );
not ( n271461 , n271460 );
not ( n271462 , n245950 );
or ( n271463 , n271461 , n271462 );
or ( n271464 , n245950 , n271460 );
nand ( n271465 , n271463 , n271464 );
and ( n271466 , n271465 , n261351 );
not ( n271467 , n271465 );
and ( n271468 , n271467 , n226319 );
nor ( n271469 , n271466 , n271468 );
buf ( n271470 , n242163 );
not ( n271471 , n271470 );
not ( n271472 , n27876 );
or ( n271473 , n271471 , n271472 );
not ( n271474 , n271470 );
nand ( n271475 , n271474 , n27869 );
nand ( n271476 , n271473 , n271475 );
and ( n271477 , n271476 , n248756 );
not ( n271478 , n271476 );
and ( n271479 , n271478 , n248763 );
nor ( n271480 , n271477 , n271479 );
nor ( n271481 , n271469 , n271480 );
or ( n271482 , n271459 , n271481 );
nor ( n271483 , n271458 , n219702 );
nand ( n271484 , n271483 , n271481 );
nand ( n271485 , n247585 , n29630 );
nand ( n271486 , n271482 , n271484 , n271485 );
buf ( n271487 , n271486 );
not ( n271488 , n238183 );
not ( n271489 , n55881 );
not ( n271490 , n271489 );
not ( n271491 , n49181 );
or ( n271492 , n271490 , n271491 );
nand ( n271493 , n49190 , n55881 );
nand ( n271494 , n271492 , n271493 );
not ( n271495 , n271494 );
or ( n271496 , n271488 , n271495 );
or ( n271497 , n271494 , n238183 );
nand ( n271498 , n271496 , n271497 );
not ( n271499 , n271498 );
not ( n271500 , n271499 );
not ( n271501 , n269451 );
not ( n271502 , n271501 );
or ( n271503 , n271500 , n271502 );
not ( n271504 , n248356 );
not ( n271505 , n271504 );
not ( n271506 , n246321 );
or ( n271507 , n271505 , n271506 );
not ( n271508 , n271504 );
nand ( n271509 , n271508 , n246326 );
nand ( n271510 , n271507 , n271509 );
and ( n271511 , n271510 , n246331 );
not ( n271512 , n271510 );
and ( n271513 , n271512 , n254483 );
nor ( n271514 , n271511 , n271513 );
nor ( n271515 , n271514 , n240080 );
nand ( n271516 , n271503 , n271515 );
not ( n271517 , n271514 );
nor ( n271518 , n271517 , n271498 );
nand ( n271519 , n269454 , n271518 );
nand ( n271520 , n251712 , n204794 );
nand ( n271521 , n271516 , n271519 , n271520 );
buf ( n271522 , n271521 );
nand ( n271523 , n253719 , n260375 );
not ( n271524 , n256284 );
nand ( n271525 , n271524 , n253749 );
or ( n271526 , n271523 , n271525 );
not ( n271527 , n271524 );
not ( n271528 , n253719 );
or ( n271529 , n271527 , n271528 );
nor ( n271530 , n253749 , n254740 );
nand ( n271531 , n271529 , n271530 );
nand ( n271532 , n251465 , n35251 );
nand ( n271533 , n271526 , n271531 , n271532 );
buf ( n271534 , n271533 );
not ( n271535 , RI19a887a8_2735);
or ( n271536 , n25328 , n271535 );
not ( n271537 , RI19a86fc0_2745);
or ( n271538 , n25336 , n271537 );
nand ( n271539 , n271536 , n271538 );
buf ( n271540 , n271539 );
buf ( n271541 , n30397 );
not ( n271542 , n55255 );
not ( n271543 , n239390 );
or ( n271544 , n271542 , n271543 );
or ( n271545 , n239390 , n55255 );
nand ( n271546 , n271544 , n271545 );
and ( n271547 , n271546 , n249021 );
not ( n271548 , n271546 );
and ( n271549 , n271548 , n249018 );
nor ( n271550 , n271547 , n271549 );
nand ( n271551 , n271550 , n267934 );
not ( n271552 , n269649 );
nand ( n271553 , n271552 , n222531 );
or ( n271554 , n271551 , n271553 );
nor ( n271555 , n271552 , n249531 );
nand ( n271556 , n271551 , n271555 );
nand ( n271557 , n234453 , n30330 );
nand ( n271558 , n271554 , n271556 , n271557 );
buf ( n271559 , n271558 );
buf ( n271560 , n33269 );
not ( n271561 , n271156 );
nor ( n271562 , n271561 , n238635 );
not ( n271563 , n246950 );
not ( n271564 , n256191 );
or ( n271565 , n271563 , n271564 );
not ( n271566 , n246950 );
nand ( n271567 , n271566 , n256190 );
nand ( n271568 , n271565 , n271567 );
and ( n271569 , n271568 , n249849 );
not ( n271570 , n271568 );
and ( n271571 , n271570 , n260022 );
nor ( n271572 , n271569 , n271571 );
not ( n271573 , n271572 );
nand ( n271574 , n271562 , n271573 );
nor ( n271575 , n271156 , n249531 );
nor ( n271576 , n271573 , n271177 );
nand ( n271577 , n271575 , n271576 );
nor ( n271578 , n271572 , n246680 );
nand ( n271579 , n271578 , n271177 );
nand ( n271580 , n31577 , n33875 );
nand ( n271581 , n271574 , n271577 , n271579 , n271580 );
buf ( n271582 , n271581 );
nand ( n271583 , n248977 , n254013 );
nand ( n271584 , n248992 , n265076 );
or ( n271585 , n271583 , n271584 );
not ( n271586 , n248992 );
not ( n271587 , n248977 );
or ( n271588 , n271586 , n271587 );
nor ( n271589 , n265076 , n244216 );
nand ( n271590 , n271588 , n271589 );
nand ( n271591 , n263598 , n28769 );
nand ( n271592 , n271585 , n271590 , n271591 );
buf ( n271593 , n271592 );
not ( n271594 , n261886 );
not ( n271595 , n247877 );
or ( n271596 , n271594 , n271595 );
nor ( n271597 , n261897 , n49051 );
nand ( n271598 , n271596 , n271597 );
nor ( n271599 , n261899 , n33254 );
nand ( n271600 , n247877 , n271599 , n261897 );
nand ( n271601 , n239240 , n204478 );
nand ( n271602 , n271598 , n271600 , n271601 );
buf ( n271603 , n271602 );
not ( n271604 , RI19a93ba8_2656);
or ( n271605 , n233507 , n271604 );
not ( n271606 , RI19a89888_2727);
or ( n271607 , n25336 , n271606 );
nand ( n271608 , n271605 , n271607 );
buf ( n271609 , n271608 );
not ( n271610 , n231996 );
not ( n271611 , n252192 );
or ( n271612 , n271610 , n271611 );
not ( n271613 , n263965 );
or ( n271614 , n271613 , n231996 );
nand ( n271615 , n271612 , n271614 );
and ( n271616 , n271615 , n268643 );
not ( n271617 , n271615 );
and ( n271618 , n271617 , n268640 );
nor ( n271619 , n271616 , n271618 );
not ( n271620 , n271619 );
not ( n271621 , n247415 );
not ( n271622 , n271621 );
or ( n271623 , n271620 , n271622 );
nor ( n271624 , n247297 , n251862 );
nand ( n271625 , n271623 , n271624 );
nor ( n271626 , n247415 , n37725 );
nand ( n271627 , n271626 , n247297 , n271619 );
nand ( n271628 , n255116 , n32188 );
nand ( n271629 , n271625 , n271627 , n271628 );
buf ( n271630 , n271629 );
or ( n271631 , n25328 , n264402 );
or ( n271632 , n25336 , n258785 );
nand ( n271633 , n271631 , n271632 );
buf ( n271634 , n271633 );
or ( n271635 , n226819 , n246223 );
or ( n271636 , n25335 , n261448 );
nand ( n271637 , n271635 , n271636 );
buf ( n271638 , n271637 );
buf ( n271639 , n39914 );
not ( n271640 , n255614 );
nand ( n271641 , n271640 , n257421 );
or ( n271642 , n271641 , n255628 );
not ( n271643 , n255627 );
not ( n271644 , n271640 );
or ( n271645 , n271643 , n271644 );
nor ( n271646 , n257421 , n234110 );
nand ( n271647 , n271645 , n271646 );
nand ( n271648 , n241976 , n29157 );
nand ( n271649 , n271642 , n271647 , n271648 );
buf ( n271650 , n271649 );
buf ( n271651 , n36335 );
not ( n271652 , n38103 );
not ( n271653 , n245943 );
or ( n271654 , n271652 , n271653 );
not ( n271655 , n257708 );
nand ( n271656 , n271655 , n257696 );
not ( n271657 , n234155 );
not ( n271658 , n251619 );
or ( n271659 , n271657 , n271658 );
not ( n271660 , n234155 );
nand ( n271661 , n271660 , n251627 );
nand ( n271662 , n271659 , n271661 );
and ( n271663 , n271662 , n251573 );
not ( n271664 , n271662 );
and ( n271665 , n271664 , n258961 );
nor ( n271666 , n271663 , n271665 );
not ( n271667 , n271666 );
and ( n271668 , n271656 , n271667 );
not ( n271669 , n271656 );
and ( n271670 , n271669 , n271666 );
nor ( n271671 , n271668 , n271670 );
or ( n271672 , n271671 , n244217 );
nand ( n271673 , n271654 , n271672 );
buf ( n271674 , n271673 );
buf ( n271675 , n31991 );
buf ( n271676 , n26188 );
buf ( n271677 , n33929 );
buf ( n271678 , n37063 );
not ( n271679 , n252530 );
not ( n271680 , n249362 );
or ( n271681 , n271679 , n271680 );
not ( n271682 , n252530 );
not ( n271683 , n261542 );
nand ( n271684 , n271682 , n271683 );
nand ( n271685 , n271681 , n271684 );
and ( n271686 , n271685 , n261550 );
not ( n271687 , n271685 );
and ( n271688 , n271687 , n261547 );
nor ( n271689 , n271686 , n271688 );
not ( n271690 , n271689 );
nand ( n271691 , n247699 , n271690 );
nor ( n271692 , n247738 , n243434 );
nor ( n271693 , n271690 , n247735 );
nand ( n271694 , n271692 , n271693 );
nor ( n271695 , n271689 , n219702 );
nand ( n271696 , n271695 , n247735 );
nand ( n271697 , n253486 , n25620 );
nand ( n271698 , n271691 , n271694 , n271696 , n271697 );
buf ( n271699 , n271698 );
or ( n271700 , n25328 , n264262 );
not ( n271701 , RI19ab8430_2393);
or ( n271702 , n226822 , n271701 );
nand ( n271703 , n271700 , n271702 );
buf ( n271704 , n271703 );
not ( n271705 , RI19aa9430_2501);
or ( n271706 , n25328 , n271705 );
not ( n271707 , RI19a9f728_2573);
or ( n271708 , n25335 , n271707 );
nand ( n271709 , n271706 , n271708 );
buf ( n271710 , n271709 );
or ( n271711 , n233507 , n268339 );
not ( n271712 , RI19aad300_2474);
or ( n271713 , n25336 , n271712 );
nand ( n271714 , n271711 , n271713 );
buf ( n271715 , n271714 );
buf ( n271716 , n31457 );
not ( n271717 , n37054 );
not ( n271718 , n245702 );
or ( n271719 , n271717 , n271718 );
buf ( n271720 , n52642 );
not ( n271721 , n271720 );
not ( n271722 , n258610 );
not ( n271723 , n271722 );
or ( n271724 , n271721 , n271723 );
or ( n271725 , n269446 , n271720 );
nand ( n271726 , n271724 , n271725 );
not ( n271727 , n271726 );
not ( n271728 , n242527 );
and ( n271729 , n271727 , n271728 );
and ( n271730 , n271726 , n258622 );
nor ( n271731 , n271729 , n271730 );
not ( n271732 , n53454 );
not ( n271733 , n32537 );
not ( n271734 , n53248 );
or ( n271735 , n271733 , n271734 );
not ( n271736 , n32537 );
nand ( n271737 , n271736 , n53257 );
nand ( n271738 , n271735 , n271737 );
not ( n271739 , n271738 );
or ( n271740 , n271732 , n271739 );
or ( n271741 , n271738 , n53694 );
nand ( n271742 , n271740 , n271741 );
nand ( n271743 , n271731 , n271742 );
not ( n271744 , n257942 );
not ( n271745 , n271744 );
not ( n271746 , n250681 );
or ( n271747 , n271745 , n271746 );
not ( n271748 , n271744 );
nand ( n271749 , n271748 , n250691 );
nand ( n271750 , n271747 , n271749 );
and ( n271751 , n271750 , n262220 );
not ( n271752 , n271750 );
and ( n271753 , n271752 , n262217 );
nor ( n271754 , n271751 , n271753 );
not ( n271755 , n271754 );
and ( n271756 , n271743 , n271755 );
not ( n271757 , n271743 );
and ( n271758 , n271757 , n271754 );
nor ( n271759 , n271756 , n271758 );
or ( n271760 , n271759 , n254470 );
nand ( n271761 , n271719 , n271760 );
buf ( n271762 , n271761 );
not ( n271763 , n262633 );
buf ( n271764 , n48548 );
not ( n271765 , n271764 );
not ( n271766 , n262628 );
or ( n271767 , n271765 , n271766 );
or ( n271768 , n254973 , n271764 );
nand ( n271769 , n271767 , n271768 );
not ( n271770 , n271769 );
or ( n271771 , n271763 , n271770 );
or ( n271772 , n271769 , n262633 );
nand ( n271773 , n271771 , n271772 );
not ( n271774 , n271773 );
not ( n271775 , n271774 );
not ( n271776 , n270377 );
not ( n271777 , n271776 );
or ( n271778 , n271775 , n271777 );
nand ( n271779 , n271778 , n268669 );
nor ( n271780 , n268696 , n271773 );
nand ( n271781 , n270380 , n271780 );
nand ( n271782 , n247744 , n37503 );
nand ( n271783 , n271779 , n271781 , n271782 );
buf ( n271784 , n271783 );
buf ( n271785 , n36845 );
buf ( n271786 , n241300 );
not ( n271787 , n271786 );
not ( n271788 , n250708 );
or ( n271789 , n271787 , n271788 );
or ( n271790 , n245338 , n271786 );
nand ( n271791 , n271789 , n271790 );
not ( n271792 , n271791 );
not ( n271793 , n245393 );
and ( n271794 , n271792 , n271793 );
and ( n271795 , n271791 , n253363 );
nor ( n271796 , n271794 , n271795 );
nand ( n271797 , n271796 , n235051 );
not ( n271798 , n236755 );
not ( n271799 , n43219 );
or ( n271800 , n271798 , n271799 );
or ( n271801 , n43219 , n236755 );
nand ( n271802 , n271800 , n271801 );
and ( n271803 , n271802 , n261077 );
not ( n271804 , n271802 );
and ( n271805 , n271804 , n45027 );
nor ( n271806 , n271803 , n271805 );
not ( n271807 , n271806 );
not ( n271808 , n253442 );
not ( n271809 , n271808 );
not ( n271810 , n253807 );
or ( n271811 , n271809 , n271810 );
or ( n271812 , n253807 , n271808 );
nand ( n271813 , n271811 , n271812 );
not ( n271814 , n271813 );
not ( n271815 , n253813 );
or ( n271816 , n271814 , n271815 );
or ( n271817 , n262167 , n271813 );
nand ( n271818 , n271816 , n271817 );
not ( n271819 , n271818 );
nand ( n271820 , n271807 , n271819 );
or ( n271821 , n271797 , n271820 );
not ( n271822 , n271807 );
not ( n271823 , n271796 );
or ( n271824 , n271822 , n271823 );
nor ( n271825 , n271819 , n238635 );
nand ( n271826 , n271824 , n271825 );
nand ( n271827 , n31577 , n26257 );
nand ( n271828 , n271821 , n271826 , n271827 );
buf ( n271829 , n271828 );
buf ( n271830 , n206160 );
buf ( n271831 , n41350 );
not ( n271832 , n270710 );
not ( n271833 , n270705 );
or ( n271834 , n271832 , n271833 );
not ( n271835 , n236583 );
not ( n271836 , n43504 );
or ( n271837 , n271835 , n271836 );
or ( n271838 , n43504 , n236583 );
nand ( n271839 , n271837 , n271838 );
and ( n271840 , n271839 , n43219 );
not ( n271841 , n271839 );
and ( n271842 , n271841 , n268003 );
nor ( n271843 , n271840 , n271842 );
not ( n271844 , n271843 );
nor ( n271845 , n271844 , n250431 );
nand ( n271846 , n271834 , n271845 );
nor ( n271847 , n270682 , n235732 );
nand ( n271848 , n270705 , n271847 , n271844 );
nand ( n271849 , n31577 , n28088 );
nand ( n271850 , n271846 , n271848 , n271849 );
buf ( n271851 , n271850 );
not ( n271852 , RI19aac838_2479);
or ( n271853 , n25328 , n271852 );
or ( n271854 , n25335 , n266769 );
nand ( n271855 , n271853 , n271854 );
buf ( n271856 , n271855 );
not ( n271857 , n257371 );
nand ( n271858 , n271857 , n257384 );
or ( n271859 , n265741 , n271858 );
not ( n271860 , n271857 );
not ( n271861 , n265740 );
or ( n271862 , n271860 , n271861 );
nor ( n271863 , n257384 , n235050 );
nand ( n271864 , n271862 , n271863 );
nand ( n271865 , n245414 , n34673 );
nand ( n271866 , n271859 , n271864 , n271865 );
buf ( n271867 , n271866 );
not ( n271868 , RI19abaf50_2374);
or ( n271869 , n226819 , n271868 );
not ( n271870 , RI19ab11d0_2445);
or ( n271871 , n25335 , n271870 );
nand ( n271872 , n271869 , n271871 );
buf ( n271873 , n271872 );
not ( n271874 , RI19aba398_2379);
or ( n271875 , n226819 , n271874 );
not ( n271876 , RI19ab0528_2451);
or ( n271877 , n25336 , n271876 );
nand ( n271878 , n271875 , n271877 );
buf ( n271879 , n271878 );
not ( n271880 , n252987 );
not ( n271881 , n233264 );
or ( n271882 , n271880 , n271881 );
or ( n271883 , n233264 , n252987 );
nand ( n271884 , n271882 , n271883 );
and ( n271885 , n271884 , n266835 );
not ( n271886 , n271884 );
and ( n271887 , n271886 , n266838 );
nor ( n271888 , n271885 , n271887 );
nor ( n271889 , n271888 , n39763 );
not ( n271890 , n271889 );
not ( n271891 , n243484 );
not ( n271892 , n236631 );
or ( n271893 , n271891 , n271892 );
not ( n271894 , n243484 );
nand ( n271895 , n271894 , n236637 );
nand ( n271896 , n271893 , n271895 );
and ( n271897 , n271896 , n242699 );
not ( n271898 , n271896 );
and ( n271899 , n271898 , n236763 );
nor ( n271900 , n271897 , n271899 );
not ( n271901 , n271900 );
nand ( n271902 , n270165 , n271901 );
or ( n271903 , n271890 , n271902 );
not ( n271904 , n271901 );
not ( n271905 , n271888 );
not ( n271906 , n271905 );
or ( n271907 , n271904 , n271906 );
nor ( n271908 , n270165 , n234021 );
nand ( n271909 , n271907 , n271908 );
nand ( n271910 , n31577 , n28136 );
nand ( n271911 , n271903 , n271909 , n271910 );
buf ( n271912 , n271911 );
not ( n271913 , n248406 );
not ( n271914 , n221715 );
or ( n271915 , n271913 , n271914 );
not ( n271916 , n248406 );
nand ( n271917 , n271916 , n43962 );
nand ( n271918 , n271915 , n271917 );
and ( n271919 , n271918 , n255609 );
not ( n271920 , n271918 );
and ( n271921 , n271920 , n255612 );
nor ( n271922 , n271919 , n271921 );
not ( n271923 , n271922 );
nand ( n271924 , n252224 , n271923 );
or ( n271925 , n271924 , n252260 );
nand ( n271926 , n271924 , n256386 );
nand ( n271927 , n251712 , n37423 );
nand ( n271928 , n271925 , n271926 , n271927 );
buf ( n271929 , n271928 );
not ( n271930 , n249851 );
not ( n271931 , n249870 );
or ( n271932 , n271930 , n271931 );
nor ( n271933 , n262069 , n253904 );
nand ( n271934 , n271932 , n271933 );
not ( n271935 , n249851 );
nor ( n271936 , n262068 , n271935 );
nand ( n271937 , n249795 , n271936 );
nand ( n271938 , n244987 , n25843 );
nand ( n271939 , n271934 , n271937 , n271938 );
buf ( n271940 , n271939 );
not ( n271941 , RI19acba08_2242);
or ( n271942 , n25328 , n271941 );
not ( n271943 , RI19ac2a98_2309);
or ( n271944 , n25335 , n271943 );
nand ( n271945 , n271942 , n271944 );
buf ( n271946 , n271945 );
nand ( n271947 , n261462 , n223839 );
nand ( n271948 , n267861 , n261492 );
or ( n271949 , n271947 , n271948 );
not ( n271950 , n267861 );
not ( n271951 , n261462 );
or ( n271952 , n271950 , n271951 );
nor ( n271953 , n261492 , n246680 );
nand ( n271954 , n271952 , n271953 );
nand ( n271955 , n31577 , n32883 );
nand ( n271956 , n271949 , n271954 , n271955 );
buf ( n271957 , n271956 );
not ( n271958 , n259214 );
buf ( n271959 , n251832 );
not ( n271960 , n271959 );
and ( n271961 , n271958 , n271960 );
and ( n271962 , n259214 , n271959 );
nor ( n271963 , n271961 , n271962 );
and ( n271964 , n271963 , n260558 );
not ( n271965 , n271963 );
and ( n271966 , n271965 , n260551 );
nor ( n271967 , n271964 , n271966 );
nand ( n271968 , n271967 , n249009 );
not ( n271969 , n243381 );
not ( n271970 , n271969 );
not ( n271971 , n39052 );
or ( n271972 , n271970 , n271971 );
not ( n271973 , n271969 );
nand ( n271974 , n271973 , n39059 );
nand ( n271975 , n271972 , n271974 );
and ( n271976 , n271975 , n39445 );
not ( n271977 , n271975 );
and ( n271978 , n271977 , n39435 );
nor ( n271979 , n271976 , n271978 );
not ( n271980 , n271979 );
not ( n271981 , n257541 );
not ( n271982 , n35299 );
not ( n271983 , n255072 );
or ( n271984 , n271982 , n271983 );
not ( n271985 , n35299 );
nand ( n271986 , n271985 , n255071 );
nand ( n271987 , n271984 , n271986 );
not ( n271988 , n271987 );
or ( n271989 , n271981 , n271988 );
or ( n271990 , n271987 , n269931 );
nand ( n271991 , n271989 , n271990 );
not ( n271992 , n271991 );
nand ( n271993 , n271980 , n271992 );
or ( n271994 , n271968 , n271993 );
not ( n271995 , n271992 );
not ( n271996 , n271967 );
or ( n271997 , n271995 , n271996 );
nor ( n271998 , n271980 , n252070 );
nand ( n271999 , n271997 , n271998 );
nand ( n272000 , n247423 , n205367 );
nand ( n272001 , n271994 , n271999 , n272000 );
buf ( n272002 , n272001 );
not ( n272003 , RI19aa81e8_2508);
or ( n272004 , n25328 , n272003 );
not ( n272005 , RI19a9eaf8_2579);
or ( n272006 , n25335 , n272005 );
nand ( n272007 , n272004 , n272006 );
buf ( n272008 , n272007 );
not ( n272009 , n258648 );
not ( n272010 , n242927 );
not ( n272011 , n272010 );
not ( n272012 , n245929 );
or ( n272013 , n272011 , n272012 );
not ( n272014 , n272010 );
nand ( n272015 , n272014 , n245918 );
nand ( n272016 , n272013 , n272015 );
and ( n272017 , n272016 , n266165 );
not ( n272018 , n272016 );
and ( n272019 , n272018 , n266169 );
nor ( n272020 , n272017 , n272019 );
not ( n272021 , n272020 );
nand ( n272022 , n254613 , n272021 );
or ( n272023 , n272009 , n272022 );
not ( n272024 , n254613 );
not ( n272025 , n254527 );
not ( n272026 , n272025 );
or ( n272027 , n272024 , n272026 );
nor ( n272028 , n272021 , n250909 );
nand ( n272029 , n272027 , n272028 );
nand ( n272030 , n234453 , n32398 );
nand ( n272031 , n272023 , n272029 , n272030 );
buf ( n272032 , n272031 );
not ( n272033 , n36557 );
not ( n272034 , n253863 );
or ( n272035 , n272033 , n272034 );
or ( n272036 , n253863 , n36557 );
nand ( n272037 , n272035 , n272036 );
and ( n272038 , n272037 , n258013 );
not ( n272039 , n272037 );
and ( n272040 , n272039 , n239854 );
nor ( n272041 , n272038 , n272040 );
nand ( n272042 , n272041 , n239934 );
not ( n272043 , n265543 );
not ( n272044 , n254988 );
nand ( n272045 , n272043 , n272044 );
or ( n272046 , n272042 , n272045 );
not ( n272047 , n272044 );
not ( n272048 , n272041 );
or ( n272049 , n272047 , n272048 );
nor ( n272050 , n272043 , n249531 );
nand ( n272051 , n272049 , n272050 );
nand ( n272052 , n249622 , n33131 );
nand ( n272053 , n272046 , n272051 , n272052 );
buf ( n272054 , n272053 );
not ( n272055 , n34573 );
not ( n272056 , n31577 );
or ( n272057 , n272055 , n272056 );
nand ( n272058 , n259403 , n259390 );
and ( n272059 , n272058 , n259676 );
not ( n272060 , n272058 );
and ( n272061 , n272060 , n259675 );
nor ( n272062 , n272059 , n272061 );
or ( n272063 , n272062 , n251498 );
nand ( n272064 , n272057 , n272063 );
buf ( n272065 , n272064 );
not ( n272066 , n37613 );
not ( n272067 , n244789 );
or ( n272068 , n272066 , n272067 );
nand ( n272069 , n271689 , n247735 );
not ( n272070 , n244440 );
not ( n272071 , n247561 );
or ( n272072 , n272070 , n272071 );
or ( n272073 , n247561 , n244440 );
nand ( n272074 , n272072 , n272073 );
and ( n272075 , n272074 , n255006 );
not ( n272076 , n272074 );
and ( n272077 , n272076 , n270981 );
nor ( n272078 , n272075 , n272077 );
not ( n272079 , n272078 );
and ( n272080 , n272069 , n272079 );
not ( n272081 , n272069 );
and ( n272082 , n272081 , n272078 );
nor ( n272083 , n272080 , n272082 );
or ( n272084 , n272083 , n260861 );
nand ( n272085 , n272068 , n272084 );
buf ( n272086 , n272085 );
nand ( n272087 , n253328 , n269582 );
or ( n272088 , n253482 , n272087 );
not ( n272089 , n269582 );
not ( n272090 , n253481 );
or ( n272091 , n272089 , n272090 );
nor ( n272092 , n253328 , n243204 );
nand ( n272093 , n272091 , n272092 );
nand ( n272094 , n31577 , n33828 );
nand ( n272095 , n272088 , n272093 , n272094 );
buf ( n272096 , n272095 );
or ( n272097 , n25328 , n272005 );
or ( n272098 , n25335 , n254416 );
nand ( n272099 , n272097 , n272098 );
buf ( n272100 , n272099 );
not ( n272101 , n266571 );
not ( n272102 , n266560 );
not ( n272103 , n272102 );
or ( n272104 , n272101 , n272103 );
not ( n272105 , n35163 );
not ( n272106 , n223951 );
or ( n272107 , n272105 , n272106 );
or ( n272108 , n255071 , n35163 );
nand ( n272109 , n272107 , n272108 );
not ( n272110 , n272109 );
not ( n272111 , n46420 );
and ( n272112 , n272110 , n272111 );
and ( n272113 , n272109 , n257541 );
nor ( n272114 , n272112 , n272113 );
nor ( n272115 , n272114 , n251361 );
nand ( n272116 , n272104 , n272115 );
nand ( n272117 , n266573 , n272102 , n272114 );
nand ( n272118 , n237714 , n33269 );
nand ( n272119 , n272116 , n272117 , n272118 );
buf ( n272120 , n272119 );
nand ( n272121 , n250714 , n258754 );
or ( n272122 , n253104 , n272121 );
nor ( n272123 , n253103 , n54208 );
nand ( n272124 , n272123 , n272121 );
nand ( n272125 , n234823 , n30900 );
nand ( n272126 , n272122 , n272124 , n272125 );
buf ( n272127 , n272126 );
or ( n272128 , n25328 , n261336 );
or ( n272129 , n25335 , n262556 );
nand ( n272130 , n272128 , n272129 );
buf ( n272131 , n272130 );
not ( n272132 , n54423 );
not ( n272133 , n251162 );
or ( n272134 , n272132 , n272133 );
not ( n272135 , n54423 );
nand ( n272136 , n272135 , n245473 );
nand ( n272137 , n272134 , n272136 );
and ( n272138 , n272137 , n251171 );
not ( n272139 , n272137 );
and ( n272140 , n272139 , n251168 );
nor ( n272141 , n272138 , n272140 );
not ( n272142 , n29478 );
not ( n272143 , n256711 );
or ( n272144 , n272142 , n272143 );
not ( n272145 , n29478 );
nand ( n272146 , n272145 , n253009 );
nand ( n272147 , n272144 , n272146 );
and ( n272148 , n272147 , n263207 );
not ( n272149 , n272147 );
and ( n272150 , n272149 , n253015 );
nor ( n272151 , n272148 , n272150 );
not ( n272152 , n272151 );
nand ( n272153 , n272141 , n272152 );
not ( n272154 , n242547 );
not ( n272155 , n227556 );
or ( n272156 , n272154 , n272155 );
or ( n272157 , n49786 , n242547 );
nand ( n272158 , n272156 , n272157 );
and ( n272159 , n272158 , n49950 );
not ( n272160 , n272158 );
and ( n272161 , n272160 , n49947 );
nor ( n272162 , n272159 , n272161 );
not ( n272163 , n272162 );
nor ( n272164 , n272163 , n251361 );
not ( n272165 , n272164 );
or ( n272166 , n272153 , n272165 );
nor ( n272167 , n272162 , n49051 );
nand ( n272168 , n272153 , n272167 );
nand ( n272169 , n253486 , n28357 );
nand ( n272170 , n272166 , n272168 , n272169 );
buf ( n272171 , n272170 );
not ( n272172 , RI19abb298_2373);
or ( n272173 , n25328 , n272172 );
not ( n272174 , RI19ab1518_2444);
or ( n272175 , n25335 , n272174 );
nand ( n272176 , n272173 , n272175 );
buf ( n272177 , n272176 );
nand ( n272178 , n48563 , n253397 );
nand ( n272179 , n266904 , n242083 );
or ( n272180 , n272178 , n272179 );
not ( n272181 , n242083 );
not ( n272182 , n48563 );
or ( n272183 , n272181 , n272182 );
nand ( n272184 , n272183 , n266905 );
nand ( n272185 , n244840 , n37770 );
nand ( n272186 , n272180 , n272184 , n272185 );
buf ( n272187 , n272186 );
not ( n272188 , n228311 );
not ( n272189 , n31560 );
or ( n272190 , n272188 , n272189 );
not ( n272191 , n228311 );
nand ( n272192 , n272191 , n209312 );
nand ( n272193 , n272190 , n272192 );
and ( n272194 , n272193 , n35813 );
not ( n272195 , n272193 );
and ( n272196 , n272195 , n35804 );
nor ( n272197 , n272194 , n272196 );
nor ( n272198 , n268240 , n272197 );
not ( n272199 , n272198 );
not ( n272200 , n271246 );
or ( n272201 , n272199 , n272200 );
not ( n272202 , n272197 );
nor ( n272203 , n272202 , n246680 );
nand ( n272204 , n272203 , n268240 );
nand ( n272205 , n272201 , n272204 );
not ( n272206 , n272205 );
not ( n272207 , n268229 );
nand ( n272208 , n272207 , n272197 );
nand ( n272209 , n250916 , n36593 );
nand ( n272210 , n272206 , n272208 , n272209 );
buf ( n272211 , n272210 );
or ( n272212 , n25328 , n253912 );
not ( n272213 , RI19abddb8_2351);
or ( n272214 , n226822 , n272213 );
nand ( n272215 , n272212 , n272214 );
buf ( n272216 , n272215 );
not ( n272217 , RI19ac3d58_2300);
or ( n272218 , n233507 , n272217 );
not ( n272219 , RI19abb5e0_2372);
or ( n272220 , n226822 , n272219 );
nand ( n272221 , n272218 , n272220 );
buf ( n272222 , n272221 );
not ( n272223 , n258722 );
not ( n272224 , n204985 );
not ( n272225 , n228364 );
or ( n272226 , n272224 , n272225 );
not ( n272227 , n204985 );
nand ( n272228 , n272227 , n50539 );
nand ( n272229 , n272226 , n272228 );
not ( n272230 , n272229 );
not ( n272231 , n55727 );
and ( n272232 , n272230 , n272231 );
and ( n272233 , n272229 , n55727 );
nor ( n272234 , n272232 , n272233 );
nand ( n272235 , n272223 , n272234 );
not ( n272236 , n35427 );
nand ( n272237 , n272236 , n267249 );
or ( n272238 , n272235 , n272237 );
nand ( n272239 , n272235 , n267256 );
nand ( n272240 , n39767 , n41730 );
nand ( n272241 , n272238 , n272239 , n272240 );
buf ( n272242 , n272241 );
not ( n272243 , n271065 );
nand ( n272244 , n272243 , n259847 );
not ( n272245 , n253413 );
not ( n272246 , n259385 );
or ( n272247 , n272245 , n272246 );
not ( n272248 , n253413 );
nand ( n272249 , n272248 , n253807 );
nand ( n272250 , n272247 , n272249 );
and ( n272251 , n272250 , n253813 );
not ( n272252 , n272250 );
not ( n272253 , n262167 );
and ( n272254 , n272252 , n272253 );
nor ( n272255 , n272251 , n272254 );
nand ( n272256 , n271076 , n272255 );
or ( n272257 , n272244 , n272256 );
not ( n272258 , n271076 );
not ( n272259 , n272243 );
or ( n272260 , n272258 , n272259 );
nor ( n272261 , n272255 , n55108 );
nand ( n272262 , n272260 , n272261 );
nand ( n272263 , n238638 , n204787 );
nand ( n272264 , n272257 , n272262 , n272263 );
buf ( n272265 , n272264 );
not ( n272266 , n204662 );
not ( n272267 , n244606 );
or ( n272268 , n272266 , n272267 );
not ( n272269 , RI1754af18_51);
or ( n272270 , n269544 , n272269 );
nand ( n272271 , n272268 , n272270 );
buf ( n272272 , n272271 );
nand ( n272273 , n269122 , n269144 );
not ( n272274 , n245770 );
not ( n272275 , n52756 );
or ( n272276 , n272274 , n272275 );
not ( n272277 , n245770 );
nand ( n272278 , n272277 , n245264 );
nand ( n272279 , n272276 , n272278 );
and ( n272280 , n272279 , n251156 );
not ( n272281 , n272279 );
and ( n272282 , n272281 , n252733 );
nor ( n272283 , n272280 , n272282 );
not ( n272284 , n272283 );
nand ( n272285 , n272273 , n272284 , n253393 );
not ( n272286 , n269144 );
nor ( n272287 , n272286 , n258179 );
nand ( n272288 , n272287 , n272283 , n269122 );
nand ( n272289 , n246460 , n27681 );
nand ( n272290 , n272285 , n272288 , n272289 );
buf ( n272291 , n272290 );
not ( n272292 , n248470 );
nand ( n272293 , n248484 , n263521 , n272292 );
not ( n272294 , n248487 );
not ( n272295 , n272292 );
or ( n272296 , n272294 , n272295 );
nor ( n272297 , n263521 , n55152 );
nand ( n272298 , n272296 , n272297 );
nand ( n272299 , n238638 , n35919 );
nand ( n272300 , n272293 , n272298 , n272299 );
buf ( n272301 , n272300 );
not ( n272302 , RI19a90368_2681);
or ( n272303 , n25328 , n272302 );
or ( n272304 , n25335 , n257473 );
nand ( n272305 , n272303 , n272304 );
buf ( n272306 , n272305 );
nand ( n272307 , n207728 , n261808 );
or ( n272308 , n265606 , n272307 );
not ( n272309 , n27880 );
not ( n272310 , n207728 );
or ( n272311 , n272309 , n272310 );
nor ( n272312 , n261808 , n52445 );
nand ( n272313 , n272311 , n272312 );
nand ( n272314 , n253486 , n39790 );
nand ( n272315 , n272308 , n272313 , n272314 );
buf ( n272316 , n272315 );
buf ( n272317 , n39965 );
buf ( n272318 , n207855 );
nand ( n272319 , n240813 , n243438 );
nand ( n272320 , n264558 , n240998 );
or ( n272321 , n272319 , n272320 );
not ( n272322 , n240998 );
not ( n272323 , n240813 );
or ( n272324 , n272322 , n272323 );
nor ( n272325 , n264558 , n40465 );
nand ( n272326 , n272324 , n272325 );
nand ( n272327 , n234024 , n204490 );
nand ( n272328 , n272321 , n272326 , n272327 );
buf ( n272329 , n272328 );
not ( n272330 , n261530 );
nand ( n272331 , n272330 , n254528 );
not ( n272332 , n250234 );
not ( n272333 , n254707 );
not ( n272334 , n249600 );
or ( n272335 , n272333 , n272334 );
or ( n272336 , n249600 , n254707 );
nand ( n272337 , n272335 , n272336 );
not ( n272338 , n272337 );
and ( n272339 , n272332 , n272338 );
and ( n272340 , n250234 , n272337 );
nor ( n272341 , n272339 , n272340 );
nand ( n272342 , n266672 , n272341 );
or ( n272343 , n272331 , n272342 );
not ( n272344 , n266672 );
not ( n272345 , n272330 );
or ( n272346 , n272344 , n272345 );
nor ( n272347 , n272341 , n50944 );
nand ( n272348 , n272346 , n272347 );
nand ( n272349 , n239240 , n34240 );
nand ( n272350 , n272343 , n272348 , n272349 );
buf ( n272351 , n272350 );
not ( n272352 , RI19abe9e8_2344);
or ( n272353 , n25328 , n272352 );
or ( n272354 , n226822 , n270933 );
nand ( n272355 , n272353 , n272354 );
buf ( n272356 , n272355 );
not ( n272357 , n46679 );
not ( n272358 , n253188 );
or ( n272359 , n272357 , n272358 );
or ( n272360 , n253188 , n46679 );
nand ( n272361 , n272359 , n272360 );
and ( n272362 , n272361 , n253949 );
not ( n272363 , n272361 );
and ( n272364 , n272363 , n263613 );
nor ( n272365 , n272362 , n272364 );
nand ( n272366 , n272365 , n269409 );
not ( n272367 , n244235 );
not ( n272368 , n28929 );
or ( n272369 , n272367 , n272368 );
not ( n272370 , n244235 );
nand ( n272371 , n272370 , n28936 );
nand ( n272372 , n272369 , n272371 );
and ( n272373 , n272372 , n262379 );
not ( n272374 , n272372 );
and ( n272375 , n272374 , n29965 );
nor ( n272376 , n272373 , n272375 );
not ( n272377 , n272376 );
not ( n272378 , n269739 );
nand ( n272379 , n272377 , n272378 );
or ( n272380 , n272366 , n272379 );
not ( n272381 , n272377 );
not ( n272382 , n272365 );
or ( n272383 , n272381 , n272382 );
nor ( n272384 , n272378 , n37725 );
nand ( n272385 , n272383 , n272384 );
nand ( n272386 , n35431 , n25935 );
nand ( n272387 , n272380 , n272385 , n272386 );
buf ( n272388 , n272387 );
not ( n272389 , RI1754b080_48);
or ( n272390 , n249126 , n272389 );
nand ( n272391 , n249131 , n31595 );
nand ( n272392 , n272390 , n272391 );
buf ( n272393 , n272392 );
not ( n272394 , n35056 );
not ( n272395 , n50615 );
or ( n272396 , n272394 , n272395 );
not ( n272397 , n263521 );
nand ( n272398 , n272397 , n263532 );
and ( n272399 , n272398 , n248461 );
not ( n272400 , n272398 );
not ( n272401 , n248461 );
and ( n272402 , n272400 , n272401 );
nor ( n272403 , n272399 , n272402 );
or ( n272404 , n272403 , n245938 );
nand ( n272405 , n272396 , n272404 );
buf ( n272406 , n272405 );
nand ( n272407 , n249063 , n252873 );
not ( n272408 , n249115 );
not ( n272409 , n265594 );
nand ( n272410 , n272408 , n272409 );
or ( n272411 , n272407 , n272410 );
not ( n272412 , n272409 );
not ( n272413 , n249063 );
or ( n272414 , n272412 , n272413 );
nor ( n272415 , n272408 , n50944 );
nand ( n272416 , n272414 , n272415 );
nand ( n272417 , n237361 , n38892 );
nand ( n272418 , n272411 , n272416 , n272417 );
buf ( n272419 , n272418 );
nand ( n272420 , n270175 , n270153 );
not ( n272421 , n272420 );
not ( n272422 , n271889 );
or ( n272423 , n272421 , n272422 );
and ( n272424 , n271888 , n270184 , n270175 );
not ( n272425 , n41725 );
nor ( n272426 , n272425 , n263991 );
nor ( n272427 , n272424 , n272426 );
nand ( n272428 , n272423 , n272427 );
buf ( n272429 , n272428 );
not ( n272430 , n233692 );
not ( n272431 , n262430 );
or ( n272432 , n272430 , n272431 );
or ( n272433 , n262430 , n233692 );
nand ( n272434 , n272432 , n272433 );
and ( n272435 , n272434 , n251220 );
not ( n272436 , n272434 );
and ( n272437 , n272436 , n251224 );
nor ( n272438 , n272435 , n272437 );
not ( n272439 , n223546 );
not ( n272440 , n36729 );
or ( n272441 , n272439 , n272440 );
not ( n272442 , n223546 );
nand ( n272443 , n272442 , n249482 );
nand ( n272444 , n272441 , n272443 );
and ( n272445 , n272444 , n249491 );
not ( n272446 , n272444 );
and ( n272447 , n272446 , n249495 );
nor ( n272448 , n272445 , n272447 );
not ( n272449 , n272448 );
nand ( n272450 , n262720 , n272438 , n272449 );
not ( n272451 , n262700 );
not ( n272452 , n272451 );
not ( n272453 , n272438 );
or ( n272454 , n272452 , n272453 );
nor ( n272455 , n272449 , n236795 );
nand ( n272456 , n272454 , n272455 );
nand ( n272457 , n31577 , n208380 );
nand ( n272458 , n272450 , n272456 , n272457 );
buf ( n272459 , n272458 );
not ( n272460 , n38149 );
not ( n272461 , n31577 );
or ( n272462 , n272460 , n272461 );
not ( n272463 , n268894 );
nand ( n272464 , n272463 , n268884 );
not ( n272465 , n246846 );
not ( n272466 , n272465 );
not ( n272467 , n255496 );
or ( n272468 , n272466 , n272467 );
or ( n272469 , n255496 , n272465 );
nand ( n272470 , n272468 , n272469 );
and ( n272471 , n272470 , n242866 );
not ( n272472 , n272470 );
and ( n272473 , n272472 , n208725 );
nor ( n272474 , n272471 , n272473 );
and ( n272475 , n272464 , n272474 );
not ( n272476 , n272464 );
not ( n272477 , n272474 );
and ( n272478 , n272476 , n272477 );
nor ( n272479 , n272475 , n272478 );
or ( n272480 , n272479 , n254515 );
nand ( n272481 , n272462 , n272480 );
buf ( n272482 , n272481 );
or ( n272483 , n25328 , n264220 );
not ( n272484 , RI19abf4b0_2338);
or ( n272485 , n25335 , n272484 );
nand ( n272486 , n272483 , n272485 );
buf ( n272487 , n272486 );
or ( n272488 , n233507 , n272219 );
not ( n272489 , RI19ab16f8_2443);
or ( n272490 , n25335 , n272489 );
nand ( n272491 , n272488 , n272490 );
buf ( n272492 , n272491 );
nand ( n272493 , n231217 , n268556 );
nor ( n272494 , n270346 , n33254 );
not ( n272495 , n272494 );
or ( n272496 , n272493 , n272495 );
nand ( n272497 , n270348 , n272493 );
nand ( n272498 , n244987 , n25482 );
nand ( n272499 , n272496 , n272497 , n272498 );
buf ( n272500 , n272499 );
not ( n272501 , n31327 );
not ( n272502 , n237361 );
or ( n272503 , n272501 , n272502 );
nand ( n272504 , n268183 , n268195 );
not ( n272505 , n246064 );
not ( n272506 , n243942 );
and ( n272507 , n272505 , n272506 );
and ( n272508 , n246064 , n243942 );
nor ( n272509 , n272507 , n272508 );
not ( n272510 , n272509 );
not ( n272511 , n272510 );
not ( n272512 , n246768 );
or ( n272513 , n272511 , n272512 );
nand ( n272514 , n246760 , n272509 );
nand ( n272515 , n272513 , n272514 );
and ( n272516 , n272504 , n272515 );
not ( n272517 , n272504 );
not ( n272518 , n272515 );
and ( n272519 , n272517 , n272518 );
nor ( n272520 , n272516 , n272519 );
or ( n272521 , n272520 , n255967 );
nand ( n272522 , n272503 , n272521 );
buf ( n272523 , n272522 );
not ( n272524 , n32580 );
not ( n272525 , n262000 );
or ( n272526 , n272524 , n272525 );
not ( n272527 , n269615 );
nand ( n272528 , n272527 , n269501 );
not ( n272529 , n269512 );
and ( n272530 , n272528 , n272529 );
not ( n272531 , n272528 );
and ( n272532 , n272531 , n269512 );
nor ( n272533 , n272530 , n272532 );
or ( n272534 , n272533 , n258179 );
nand ( n272535 , n272526 , n272534 );
buf ( n272536 , n272535 );
not ( n272537 , RI1754a720_68);
not ( n272538 , n25326 );
or ( n272539 , n272537 , n272538 );
nand ( n272540 , n272539 , n266632 );
buf ( n272541 , n272540 );
not ( n272542 , n237047 );
not ( n272543 , n253073 );
or ( n272544 , n272542 , n272543 );
or ( n272545 , n253073 , n237047 );
nand ( n272546 , n272544 , n272545 );
and ( n272547 , n272546 , n257658 );
not ( n272548 , n272546 );
and ( n272549 , n272548 , n257659 );
nor ( n272550 , n272547 , n272549 );
nand ( n272551 , n272550 , n223839 );
buf ( n272552 , n246362 );
not ( n272553 , n272552 );
not ( n272554 , n44539 );
or ( n272555 , n272553 , n272554 );
or ( n272556 , n44539 , n272552 );
nand ( n272557 , n272555 , n272556 );
and ( n272558 , n272557 , n260442 );
not ( n272559 , n272557 );
and ( n272560 , n272559 , n222525 );
nor ( n272561 , n272558 , n272560 );
nand ( n272562 , n262900 , n272561 );
or ( n272563 , n272551 , n272562 );
not ( n272564 , n272561 );
not ( n272565 , n272550 );
or ( n272566 , n272564 , n272565 );
nor ( n272567 , n262900 , n247698 );
nand ( n272568 , n272566 , n272567 );
nand ( n272569 , n236798 , n29941 );
nand ( n272570 , n272563 , n272568 , n272569 );
buf ( n272571 , n272570 );
not ( n272572 , n41916 );
not ( n272573 , n233090 );
or ( n272574 , n272572 , n272573 );
nand ( n272575 , n55322 , n41917 );
nand ( n272576 , n272574 , n272575 );
not ( n272577 , n272576 );
not ( n272578 , n242272 );
and ( n272579 , n272577 , n272578 );
and ( n272580 , n272576 , n242272 );
nor ( n272581 , n272579 , n272580 );
not ( n272582 , n272581 );
not ( n272583 , n244686 );
not ( n272584 , n241715 );
or ( n272585 , n272583 , n272584 );
not ( n272586 , n244686 );
nand ( n272587 , n272586 , n241723 );
nand ( n272588 , n272585 , n272587 );
and ( n272589 , n272588 , n241885 );
not ( n272590 , n272588 );
and ( n272591 , n272590 , n241878 );
nor ( n272592 , n272589 , n272591 );
nand ( n272593 , n272582 , n272592 );
not ( n272594 , n234017 );
nor ( n272595 , n272594 , n252070 );
not ( n272596 , n272595 );
or ( n272597 , n272593 , n272596 );
nand ( n272598 , n272593 , n234022 );
nand ( n272599 , n31577 , n32832 );
nand ( n272600 , n272597 , n272598 , n272599 );
buf ( n272601 , n272600 );
buf ( n272602 , n38126 );
buf ( n272603 , RI17539830_589);
and ( n272604 , n27883 , n272603 );
buf ( n272605 , n272604 );
not ( n272606 , n272378 );
not ( n272607 , n272365 );
not ( n272608 , n272607 );
or ( n272609 , n272606 , n272608 );
nor ( n272610 , n269729 , n40465 );
nand ( n272611 , n272609 , n272610 );
nor ( n272612 , n272365 , n55152 );
nor ( n272613 , n269728 , n269739 );
nand ( n272614 , n272612 , n272613 );
nand ( n272615 , n261585 , n31981 );
nand ( n272616 , n272611 , n272614 , n272615 );
buf ( n272617 , n272616 );
not ( n272618 , n237394 );
not ( n272619 , n247822 );
or ( n272620 , n272618 , n272619 );
or ( n272621 , n247822 , n237394 );
nand ( n272622 , n272620 , n272621 );
and ( n272623 , n272622 , n247872 );
not ( n272624 , n272622 );
and ( n272625 , n272624 , n247873 );
nor ( n272626 , n272623 , n272625 );
nand ( n272627 , n272626 , n239934 );
not ( n272628 , n264861 );
not ( n272629 , n258803 );
nand ( n272630 , n272628 , n272629 );
or ( n272631 , n272627 , n272630 );
not ( n272632 , n272628 );
not ( n272633 , n272626 );
or ( n272634 , n272632 , n272633 );
nor ( n272635 , n272629 , n234021 );
nand ( n272636 , n272634 , n272635 );
nand ( n272637 , n247744 , n26233 );
nand ( n272638 , n272631 , n272636 , n272637 );
buf ( n272639 , n272638 );
not ( n272640 , n271597 );
nand ( n272641 , n247773 , n247762 );
or ( n272642 , n272640 , n272641 );
not ( n272643 , n261897 );
nand ( n272644 , n272643 , n247762 );
not ( n272645 , n247773 );
nand ( n272646 , n272644 , n272645 , n50945 );
nand ( n272647 , n256673 , n31951 );
nand ( n272648 , n272642 , n272646 , n272647 );
buf ( n272649 , n272648 );
or ( n272650 , n25328 , n269999 );
not ( n272651 , RI19ab0870_2450);
or ( n272652 , n25336 , n272651 );
nand ( n272653 , n272650 , n272652 );
buf ( n272654 , n272653 );
nand ( n272655 , n260679 , n260689 );
nor ( n272656 , n249948 , n253904 );
not ( n272657 , n272656 );
or ( n272658 , n272655 , n272657 );
nand ( n272659 , n272655 , n249975 );
nand ( n272660 , n252711 , n204809 );
nand ( n272661 , n272658 , n272659 , n272660 );
buf ( n272662 , n272661 );
not ( n272663 , RI19aa4318_2536);
or ( n272664 , n25328 , n272663 );
not ( n272665 , RI19acf8d8_2214);
or ( n272666 , n226822 , n272665 );
nand ( n272667 , n272664 , n272666 );
buf ( n272668 , n272667 );
not ( n272669 , n224215 );
not ( n272670 , n51597 );
or ( n272671 , n272669 , n272670 );
or ( n272672 , n51597 , n224215 );
nand ( n272673 , n272671 , n272672 );
and ( n272674 , n272673 , n253197 );
not ( n272675 , n272673 );
and ( n272676 , n272675 , n253189 );
nor ( n272677 , n272674 , n272676 );
not ( n272678 , n272677 );
nand ( n272679 , n272678 , n257792 );
not ( n272680 , n272679 );
not ( n272681 , n41678 );
not ( n272682 , n233090 );
or ( n272683 , n272681 , n272682 );
not ( n272684 , n41678 );
nand ( n272685 , n272684 , n55322 );
nand ( n272686 , n272683 , n272685 );
buf ( n272687 , n252503 );
and ( n272688 , n272686 , n272687 );
not ( n272689 , n272686 );
and ( n272690 , n272689 , n242272 );
nor ( n272691 , n272688 , n272690 );
not ( n272692 , n272691 );
not ( n272693 , n253001 );
not ( n272694 , n233271 );
or ( n272695 , n272693 , n272694 );
not ( n272696 , n253001 );
nand ( n272697 , n272696 , n233264 );
nand ( n272698 , n272695 , n272697 );
and ( n272699 , n272698 , n266835 );
not ( n272700 , n272698 );
and ( n272701 , n272700 , n266838 );
nor ( n272702 , n272699 , n272701 );
nand ( n272703 , n272692 , n272702 );
not ( n272704 , n272703 );
and ( n272705 , n272680 , n272704 );
not ( n272706 , n39763 );
not ( n272707 , n272702 );
nand ( n272708 , n272706 , n272707 );
nor ( n272709 , n272708 , n272692 );
nor ( n272710 , n272705 , n272709 );
buf ( n272711 , n250111 );
nand ( n272712 , n272677 , n272711 );
not ( n272713 , n272712 );
nand ( n272714 , n272713 , n272707 );
nand ( n272715 , n37728 , n25443 );
nand ( n272716 , n272710 , n272714 , n272715 );
buf ( n272717 , n272716 );
not ( n272718 , n26349 );
not ( n272719 , n46083 );
or ( n272720 , n272718 , n272719 );
not ( n272721 , n261473 );
nand ( n272722 , n272721 , n261486 );
not ( n272723 , n267871 );
and ( n272724 , n272722 , n272723 );
not ( n272725 , n272722 );
and ( n272726 , n272725 , n267871 );
nor ( n272727 , n272724 , n272726 );
or ( n272728 , n272727 , n255707 );
nand ( n272729 , n272720 , n272728 );
buf ( n272730 , n272729 );
not ( n272731 , RI19a87218_2744);
or ( n272732 , n25328 , n272731 );
not ( n272733 , RI19acb828_2243);
or ( n272734 , n25336 , n272733 );
nand ( n272735 , n272732 , n272734 );
buf ( n272736 , n272735 );
or ( n272737 , n25328 , n266214 );
or ( n272738 , n25336 , n255020 );
nand ( n272739 , n272737 , n272738 );
buf ( n272740 , n272739 );
nor ( n272741 , n247565 , n46425 );
nand ( n272742 , n272741 , n247583 , n264450 );
not ( n272743 , n247566 );
not ( n272744 , n247583 );
or ( n272745 , n272743 , n272744 );
nor ( n272746 , n264450 , n265700 );
nand ( n272747 , n272745 , n272746 );
nand ( n272748 , n234453 , n41506 );
nand ( n272749 , n272742 , n272747 , n272748 );
buf ( n272750 , n272749 );
not ( n272751 , RI19a94b98_2649);
or ( n272752 , n226819 , n272751 );
not ( n272753 , RI19a8acb0_2719);
or ( n272754 , n25335 , n272753 );
nand ( n272755 , n272752 , n272754 );
buf ( n272756 , n272755 );
not ( n272757 , n244141 );
not ( n272758 , n234810 );
or ( n272759 , n272757 , n272758 );
not ( n272760 , n244141 );
nand ( n272761 , n272760 , n234803 );
nand ( n272762 , n272759 , n272761 );
and ( n272763 , n272762 , n250395 );
not ( n272764 , n272762 );
and ( n272765 , n272764 , n250398 );
nor ( n272766 , n272763 , n272765 );
not ( n272767 , n272766 );
not ( n272768 , n272767 );
not ( n272769 , n266841 );
or ( n272770 , n272768 , n272769 );
not ( n272771 , n55147 );
not ( n272772 , n263301 );
nor ( n272773 , n272771 , n272772 );
nand ( n272774 , n272770 , n272773 );
nor ( n272775 , n272766 , n254150 );
nand ( n272776 , n272775 , n266841 , n272772 );
nand ( n272777 , n39766 , n205165 );
nand ( n272778 , n272774 , n272776 , n272777 );
buf ( n272779 , n272778 );
nand ( n272780 , n264067 , n264080 );
nor ( n272781 , n268575 , n222533 );
not ( n272782 , n272781 );
or ( n272783 , n272780 , n272782 );
nand ( n272784 , n272780 , n268580 );
nand ( n272785 , n247585 , n29484 );
nand ( n272786 , n272783 , n272784 , n272785 );
buf ( n272787 , n272786 );
nor ( n272788 , n255408 , n246535 );
not ( n272789 , n272788 );
nand ( n272790 , n246535 , n236502 );
nand ( n272791 , n272789 , n272790 );
and ( n272792 , n272791 , n255465 );
not ( n272793 , n272791 );
and ( n272794 , n272793 , n255457 );
nor ( n272795 , n272792 , n272794 );
not ( n272796 , n272795 );
nand ( n272797 , n272796 , n259009 );
not ( n272798 , n241033 );
not ( n272799 , n272798 );
not ( n272800 , n219396 );
or ( n272801 , n272799 , n272800 );
not ( n272802 , n272798 );
nand ( n272803 , n272802 , n41632 );
nand ( n272804 , n272801 , n272803 );
and ( n272805 , n272804 , n41935 );
not ( n272806 , n272804 );
and ( n272807 , n272806 , n41930 );
nor ( n272808 , n272805 , n272807 );
not ( n272809 , n272808 );
not ( n272810 , n249284 );
not ( n272811 , n237526 );
not ( n272812 , n272811 );
not ( n272813 , n247871 );
or ( n272814 , n272812 , n272813 );
nand ( n272815 , n249276 , n237526 );
nand ( n272816 , n272814 , n272815 );
not ( n272817 , n272816 );
or ( n272818 , n272810 , n272817 );
or ( n272819 , n272816 , n263568 );
nand ( n272820 , n272818 , n272819 );
not ( n272821 , n272820 );
nand ( n272822 , n272809 , n272821 );
or ( n272823 , n272797 , n272822 );
nor ( n272824 , n272796 , n247698 );
nand ( n272825 , n272824 , n272822 );
nand ( n272826 , n247423 , n37937 );
nand ( n272827 , n272823 , n272825 , n272826 );
buf ( n272828 , n272827 );
buf ( n272829 , n36234 );
not ( n272830 , n252912 );
not ( n272831 , n241050 );
or ( n272832 , n272830 , n272831 );
not ( n272833 , n252912 );
nand ( n272834 , n272833 , n241054 );
nand ( n272835 , n272832 , n272834 );
and ( n272836 , n272835 , n241060 );
not ( n272837 , n272835 );
and ( n272838 , n272837 , n241057 );
nor ( n272839 , n272836 , n272838 );
not ( n272840 , n272839 );
not ( n272841 , n235607 );
not ( n272842 , n272841 );
not ( n272843 , n238461 );
or ( n272844 , n272842 , n272843 );
not ( n272845 , n272841 );
nand ( n272846 , n272845 , n238470 );
nand ( n272847 , n272844 , n272846 );
and ( n272848 , n272847 , n238473 );
not ( n272849 , n272847 );
and ( n272850 , n272849 , n238476 );
nor ( n272851 , n272848 , n272850 );
not ( n272852 , n272851 );
or ( n272853 , n272840 , n272852 );
not ( n272854 , n264894 );
nor ( n272855 , n272854 , n250909 );
nand ( n272856 , n272853 , n272855 );
not ( n272857 , n272839 );
nor ( n272858 , n272857 , n235732 );
nand ( n272859 , n272851 , n272858 , n272854 );
nand ( n272860 , n39767 , n49741 );
nand ( n272861 , n272856 , n272859 , n272860 );
buf ( n272862 , n272861 );
buf ( n272863 , n34554 );
buf ( n272864 , n236140 );
buf ( n272865 , n31753 );
not ( n272866 , n263831 );
nand ( n272867 , n263835 , n272866 );
or ( n272868 , n272867 , n252353 );
nand ( n272869 , n272867 , n254110 );
nand ( n272870 , n257764 , n29383 );
nand ( n272871 , n272868 , n272869 , n272870 );
buf ( n272872 , n272871 );
or ( n272873 , n233507 , n265613 );
not ( n272874 , RI19ab1860_2442);
or ( n272875 , n226822 , n272874 );
nand ( n272876 , n272873 , n272875 );
buf ( n272877 , n272876 );
or ( n272878 , n25328 , n255477 );
or ( n272879 , n25335 , n272751 );
nand ( n272880 , n272878 , n272879 );
buf ( n272881 , n272880 );
buf ( n272882 , n249834 );
not ( n272883 , n272882 );
not ( n272884 , n52995 );
not ( n272885 , n272884 );
or ( n272886 , n272883 , n272885 );
or ( n272887 , n272884 , n272882 );
nand ( n272888 , n272886 , n272887 );
and ( n272889 , n272888 , n51753 );
not ( n272890 , n272888 );
and ( n272891 , n272890 , n229518 );
nor ( n272892 , n272889 , n272891 );
nand ( n272893 , n272892 , n245176 );
or ( n272894 , n270460 , n272893 );
nand ( n272895 , n270464 , n272893 );
nand ( n272896 , n35431 , n36960 );
nand ( n272897 , n272894 , n272895 , n272896 );
buf ( n272898 , n272897 );
not ( n272899 , n235327 );
not ( n272900 , n246439 );
or ( n272901 , n272899 , n272900 );
or ( n272902 , n246439 , n235327 );
nand ( n272903 , n272901 , n272902 );
not ( n272904 , n272903 );
not ( n272905 , n254811 );
and ( n272906 , n272904 , n272905 );
and ( n272907 , n272903 , n250021 );
nor ( n272908 , n272906 , n272907 );
nor ( n272909 , n272908 , n254150 );
nor ( n272910 , n262416 , n262427 );
nand ( n272911 , n272909 , n272910 );
not ( n272912 , n262427 );
not ( n272913 , n272912 );
not ( n272914 , n272908 );
not ( n272915 , n272914 );
or ( n272916 , n272913 , n272915 );
nor ( n272917 , n262417 , n270963 );
nand ( n272918 , n272916 , n272917 );
nand ( n272919 , n31576 , n33979 );
nand ( n272920 , n272911 , n272918 , n272919 );
buf ( n272921 , n272920 );
buf ( n272922 , n29841 );
nand ( n272923 , n250282 , n248151 , n248222 );
not ( n272924 , n250277 );
not ( n272925 , n272924 );
not ( n272926 , n248151 );
or ( n272927 , n272925 , n272926 );
nor ( n272928 , n248222 , n40465 );
nand ( n272929 , n272927 , n272928 );
nand ( n272930 , n254441 , n204876 );
nand ( n272931 , n272923 , n272929 , n272930 );
buf ( n272932 , n272931 );
nand ( n272933 , n245682 , n226010 );
nand ( n272934 , n245620 , n267884 );
or ( n272935 , n272933 , n272934 );
not ( n272936 , n245682 );
not ( n272937 , n245620 );
or ( n272938 , n272936 , n272937 );
nor ( n272939 , n267884 , n247698 );
nand ( n272940 , n272938 , n272939 );
nand ( n272941 , n234024 , n28899 );
nand ( n272942 , n272935 , n272940 , n272941 );
buf ( n272943 , n272942 );
buf ( n272944 , n234411 );
not ( n272945 , n272944 );
not ( n272946 , n238106 );
or ( n272947 , n272945 , n272946 );
or ( n272948 , n238106 , n272944 );
nand ( n272949 , n272947 , n272948 );
and ( n272950 , n272949 , n244387 );
not ( n272951 , n272949 );
and ( n272952 , n272951 , n244390 );
nor ( n272953 , n272950 , n272952 );
nand ( n272954 , n272953 , n241704 );
not ( n272955 , n237770 );
not ( n272956 , n272955 );
not ( n272957 , n245392 );
or ( n272958 , n272956 , n272957 );
not ( n272959 , n272955 );
nand ( n272960 , n272959 , n245402 );
nand ( n272961 , n272958 , n272960 );
not ( n272962 , n272961 );
not ( n272963 , n259527 );
and ( n272964 , n272962 , n272963 );
and ( n272965 , n272961 , n259527 );
nor ( n272966 , n272964 , n272965 );
not ( n272967 , n52502 );
not ( n272968 , n272967 );
not ( n272969 , n269439 );
or ( n272970 , n272968 , n272969 );
nand ( n272971 , n240052 , n52502 );
nand ( n272972 , n272970 , n272971 );
not ( n272973 , n271722 );
and ( n272974 , n272972 , n272973 );
not ( n272975 , n272972 );
and ( n272976 , n272975 , n258611 );
or ( n272977 , n272974 , n272976 );
not ( n272978 , n272977 );
nand ( n272979 , n272966 , n272978 );
or ( n272980 , n272954 , n272979 );
not ( n272981 , n272966 );
not ( n272982 , n272953 );
or ( n272983 , n272981 , n272982 );
nor ( n272984 , n272978 , n55146 );
nand ( n272985 , n272983 , n272984 );
nand ( n272986 , n41945 , n28108 );
nand ( n272987 , n272980 , n272985 , n272986 );
buf ( n272988 , n272987 );
not ( n272989 , n256986 );
nand ( n272990 , n260994 , n261002 );
or ( n272991 , n272989 , n272990 );
not ( n272992 , n256980 );
not ( n272993 , n272992 );
not ( n272994 , n260994 );
or ( n272995 , n272993 , n272994 );
nor ( n272996 , n261002 , n49051 );
nand ( n272997 , n272995 , n272996 );
nand ( n272998 , n35431 , n35047 );
nand ( n272999 , n272991 , n272997 , n272998 );
buf ( n273000 , n272999 );
not ( n273001 , n32438 );
not ( n273002 , n245221 );
or ( n273003 , n273001 , n273002 );
not ( n273004 , n245068 );
not ( n273005 , n231768 );
or ( n273006 , n273004 , n273005 );
not ( n273007 , n245068 );
nand ( n273008 , n273007 , n231775 );
nand ( n273009 , n273006 , n273008 );
and ( n273010 , n273009 , n261292 );
not ( n273011 , n273009 );
and ( n273012 , n273011 , n262951 );
nor ( n273013 , n273010 , n273012 );
not ( n273014 , n273013 );
nand ( n273015 , n273014 , n262201 );
and ( n273016 , n273015 , n237973 );
not ( n273017 , n273015 );
and ( n273018 , n273017 , n262191 );
nor ( n273019 , n273016 , n273018 );
or ( n273020 , n273019 , n259651 );
nand ( n273021 , n273003 , n273020 );
buf ( n273022 , n273021 );
not ( n273023 , RI19ac8c18_2264);
or ( n273024 , n25328 , n273023 );
not ( n273025 , RI19abfc30_2334);
or ( n273026 , n25335 , n273025 );
nand ( n273027 , n273024 , n273026 );
buf ( n273028 , n273027 );
buf ( n273029 , n240881 );
not ( n273030 , n273029 );
not ( n273031 , n37708 );
or ( n273032 , n273030 , n273031 );
or ( n273033 , n37708 , n273029 );
nand ( n273034 , n273032 , n273033 );
and ( n273035 , n273034 , n244802 );
not ( n273036 , n273034 );
and ( n273037 , n273036 , n244805 );
nor ( n273038 , n273035 , n273037 );
not ( n273039 , n273038 );
nor ( n273040 , n273039 , n251862 );
not ( n273041 , n273040 );
not ( n273042 , n246569 );
not ( n273043 , n255455 );
or ( n273044 , n273042 , n273043 );
not ( n273045 , n246569 );
nand ( n273046 , n273045 , n255464 );
nand ( n273047 , n273044 , n273046 );
and ( n273048 , n273047 , n259459 );
not ( n273049 , n273047 );
and ( n273050 , n273049 , n259463 );
nor ( n273051 , n273048 , n273050 );
not ( n273052 , n273051 );
nor ( n273053 , n273052 , n264947 );
or ( n273054 , n273041 , n273053 );
nor ( n273055 , n273038 , n239237 );
nand ( n273056 , n273055 , n273053 );
nand ( n273057 , n246460 , n32551 );
nand ( n273058 , n273054 , n273056 , n273057 );
buf ( n273059 , n273058 );
not ( n273060 , n40379 );
not ( n273061 , n235878 );
or ( n273062 , n273060 , n273061 );
not ( n273063 , n40379 );
nand ( n273064 , n273063 , n235887 );
nand ( n273065 , n273062 , n273064 );
and ( n273066 , n273065 , n259855 );
not ( n273067 , n273065 );
and ( n273068 , n273067 , n259858 );
nor ( n273069 , n273066 , n273068 );
nand ( n273070 , n273069 , n261865 );
or ( n273071 , n270431 , n273070 );
not ( n273072 , n273069 );
not ( n273073 , n270430 );
or ( n273074 , n273072 , n273073 );
nand ( n273075 , n273074 , n261866 );
nand ( n273076 , n39767 , n40127 );
nand ( n273077 , n273071 , n273075 , n273076 );
buf ( n273078 , n273077 );
or ( n273079 , n25328 , n270508 );
not ( n273080 , RI19ab2328_2438);
or ( n273081 , n25335 , n273080 );
nand ( n273082 , n273079 , n273081 );
buf ( n273083 , n273082 );
not ( n273084 , RI19abbc70_2369);
or ( n273085 , n233507 , n273084 );
or ( n273086 , n226822 , n260924 );
nand ( n273087 , n273085 , n273086 );
buf ( n273088 , n273087 );
not ( n273089 , RI19ab4038_2423);
or ( n273090 , n25328 , n273089 );
or ( n273091 , n25335 , n269274 );
nand ( n273092 , n273090 , n273091 );
buf ( n273093 , n273092 );
not ( n273094 , RI19abc198_2367);
or ( n273095 , n25328 , n273094 );
not ( n273096 , RI19ab2148_2439);
or ( n273097 , n25335 , n273096 );
nand ( n273098 , n273095 , n273097 );
buf ( n273099 , n273098 );
not ( n273100 , RI19abbe50_2368);
or ( n273101 , n25328 , n273100 );
or ( n273102 , n25336 , n269222 );
nand ( n273103 , n273101 , n273102 );
buf ( n273104 , n273103 );
not ( n273105 , n29973 );
not ( n273106 , n234453 );
or ( n273107 , n273105 , n273106 );
not ( n273108 , n262030 );
nand ( n273109 , n273108 , n46424 );
not ( n273110 , n46719 );
and ( n273111 , n273109 , n273110 );
not ( n273112 , n273109 );
and ( n273113 , n273112 , n46719 );
nor ( n273114 , n273111 , n273113 );
or ( n273115 , n273114 , n52445 );
nand ( n273116 , n273107 , n273115 );
buf ( n273117 , n273116 );
buf ( n273118 , n234368 );
not ( n273119 , n273118 );
not ( n273120 , n238101 );
or ( n273121 , n273119 , n273120 );
or ( n273122 , n238101 , n273118 );
nand ( n273123 , n273121 , n273122 );
and ( n273124 , n273123 , n267001 );
not ( n273125 , n273123 );
and ( n273126 , n273125 , n266998 );
nor ( n273127 , n273124 , n273126 );
nor ( n273128 , n257455 , n273127 );
or ( n273129 , n254014 , n273128 );
nand ( n273130 , n257444 , n273128 );
nand ( n273131 , n247744 , n30512 );
nand ( n273132 , n273129 , n273130 , n273131 );
buf ( n273133 , n273132 );
not ( n273134 , n272953 );
nand ( n273135 , n273134 , n259009 );
not ( n273136 , n244433 );
not ( n273137 , n247551 );
or ( n273138 , n273136 , n273137 );
not ( n273139 , n244433 );
nand ( n273140 , n273139 , n247561 );
nand ( n273141 , n273138 , n273140 );
and ( n273142 , n273141 , n265442 );
not ( n273143 , n273141 );
and ( n273144 , n273143 , n255006 );
nor ( n273145 , n273142 , n273144 );
nand ( n273146 , n272966 , n273145 );
or ( n273147 , n273135 , n273146 );
not ( n273148 , n273145 );
not ( n273149 , n273134 );
or ( n273150 , n273148 , n273149 );
nor ( n273151 , n272966 , n260567 );
nand ( n273152 , n273150 , n273151 );
nand ( n273153 , n31577 , n209045 );
nand ( n273154 , n273147 , n273152 , n273153 );
buf ( n273155 , n273154 );
nand ( n273156 , n269213 , n244515 );
not ( n273157 , n227981 );
not ( n273158 , n248967 );
or ( n273159 , n273157 , n273158 );
not ( n273160 , n227981 );
nand ( n273161 , n273160 , n249394 );
nand ( n273162 , n273159 , n273161 );
and ( n273163 , n273162 , n248975 );
not ( n273164 , n273162 );
and ( n273165 , n273164 , n248972 );
nor ( n273166 , n273163 , n273165 );
nand ( n273167 , n273166 , n35815 );
or ( n273168 , n273156 , n273167 );
not ( n273169 , n273166 );
not ( n273170 , n269213 );
or ( n273171 , n273169 , n273170 );
nand ( n273172 , n273171 , n35817 );
nand ( n273173 , n31577 , n204399 );
nand ( n273174 , n273168 , n273172 , n273173 );
buf ( n273175 , n273174 );
buf ( n273176 , n36805 );
not ( n273177 , n204907 );
not ( n273178 , n245702 );
or ( n273179 , n273177 , n273178 );
not ( n273180 , n54377 );
not ( n273181 , n245473 );
not ( n273182 , n273181 );
or ( n273183 , n273180 , n273182 );
not ( n273184 , n54377 );
nand ( n273185 , n273184 , n245473 );
nand ( n273186 , n273183 , n273185 );
and ( n273187 , n273186 , n251171 );
not ( n273188 , n273186 );
and ( n273189 , n273188 , n251168 );
nor ( n273190 , n273187 , n273189 );
not ( n273191 , n273190 );
not ( n273192 , n266333 );
nand ( n273193 , n273191 , n273192 );
xor ( n273194 , n238833 , n247500 );
and ( n273195 , n273194 , n247553 );
not ( n273196 , n273194 );
and ( n273197 , n273196 , n247563 );
nor ( n273198 , n273195 , n273197 );
not ( n273199 , n273198 );
and ( n273200 , n273193 , n273199 );
not ( n273201 , n273193 );
and ( n273202 , n273201 , n273198 );
nor ( n273203 , n273200 , n273202 );
or ( n273204 , n273203 , n254470 );
nand ( n273205 , n273179 , n273204 );
buf ( n273206 , n273205 );
not ( n273207 , n234136 );
not ( n273208 , n251619 );
or ( n273209 , n273207 , n273208 );
not ( n273210 , n234136 );
nand ( n273211 , n273210 , n251627 );
nand ( n273212 , n273209 , n273211 );
and ( n273213 , n273212 , n251573 );
not ( n273214 , n273212 );
and ( n273215 , n273214 , n258961 );
nor ( n273216 , n273213 , n273215 );
not ( n273217 , n273216 );
nand ( n273218 , n271806 , n273217 );
or ( n273219 , n271797 , n273218 );
not ( n273220 , n271796 );
nand ( n273221 , n273220 , n40466 );
not ( n273222 , n273221 );
nand ( n273223 , n273222 , n273218 );
nand ( n273224 , n238638 , n36440 );
nand ( n273225 , n273219 , n273223 , n273224 );
buf ( n273226 , n273225 );
buf ( n273227 , n26269 );
not ( n273228 , n234263 );
not ( n273229 , n273228 );
not ( n273230 , n43722 );
or ( n273231 , n273229 , n273230 );
not ( n273232 , n273228 );
nand ( n273233 , n273232 , n43725 );
nand ( n273234 , n273231 , n273233 );
and ( n273235 , n273234 , n43964 );
not ( n273236 , n273234 );
and ( n273237 , n273236 , n43956 );
nor ( n273238 , n273235 , n273237 );
nor ( n273239 , n273238 , n234440 );
not ( n273240 , n235789 );
not ( n273241 , n273240 );
not ( n273242 , n245738 );
or ( n273243 , n273241 , n273242 );
nand ( n273244 , n245743 , n235789 );
nand ( n273245 , n273243 , n273244 );
and ( n273246 , n273245 , n245798 );
not ( n273247 , n273245 );
and ( n273248 , n273247 , n245799 );
nor ( n273249 , n273246 , n273248 );
not ( n273250 , n47467 );
not ( n273251 , n250899 );
or ( n273252 , n273250 , n273251 );
not ( n273253 , n47467 );
nand ( n273254 , n273253 , n250896 );
nand ( n273255 , n273252 , n273254 );
and ( n273256 , n273255 , n250903 );
not ( n273257 , n273255 );
and ( n273258 , n273257 , n250906 );
nor ( n273259 , n273256 , n273258 );
nor ( n273260 , n273249 , n273259 );
nand ( n273261 , n273239 , n273260 );
not ( n273262 , n273259 );
not ( n273263 , n273262 );
not ( n273264 , n273238 );
not ( n273265 , n273264 );
or ( n273266 , n273263 , n273265 );
not ( n273267 , n273249 );
nor ( n273268 , n273267 , n250909 );
nand ( n273269 , n273266 , n273268 );
nand ( n273270 , n37728 , n28971 );
nand ( n273271 , n273261 , n273269 , n273270 );
buf ( n273272 , n273271 );
nand ( n273273 , n238109 , n237952 );
nand ( n273274 , n273273 , n273014 , n254227 );
nand ( n273275 , n262206 , n273013 , n238109 );
nand ( n273276 , n37728 , n30801 );
nand ( n273277 , n273274 , n273275 , n273276 );
buf ( n273278 , n273277 );
or ( n273279 , n233507 , n266360 );
or ( n273280 , n226822 , n244616 );
nand ( n273281 , n273279 , n273280 );
buf ( n273282 , n273281 );
not ( n273283 , n233951 );
not ( n273284 , n244346 );
or ( n273285 , n273283 , n273284 );
or ( n273286 , n244346 , n233951 );
nand ( n273287 , n273285 , n273286 );
and ( n273288 , n273287 , n244472 );
not ( n273289 , n273287 );
and ( n273290 , n273289 , n244475 );
nor ( n273291 , n273288 , n273290 );
not ( n273292 , n273291 );
nand ( n273293 , n273292 , n247275 );
not ( n273294 , n223356 );
not ( n273295 , n248210 );
or ( n273296 , n273294 , n273295 );
not ( n273297 , n223356 );
nand ( n273298 , n273297 , n248219 );
nand ( n273299 , n273296 , n273298 );
and ( n273300 , n273299 , n261434 );
not ( n273301 , n273299 );
and ( n273302 , n273301 , n261431 );
nor ( n273303 , n273300 , n273302 );
not ( n273304 , n273303 );
not ( n273305 , n243660 );
not ( n273306 , n54176 );
not ( n273307 , n273306 );
not ( n273308 , n242380 );
or ( n273309 , n273307 , n273308 );
nand ( n273310 , n242373 , n54176 );
nand ( n273311 , n273309 , n273310 );
not ( n273312 , n273311 );
or ( n273313 , n273305 , n273312 );
or ( n273314 , n273311 , n243660 );
nand ( n273315 , n273313 , n273314 );
not ( n273316 , n273315 );
nand ( n273317 , n273304 , n273316 );
or ( n273318 , n273293 , n273317 );
not ( n273319 , n273304 );
not ( n273320 , n273292 );
or ( n273321 , n273319 , n273320 );
nor ( n273322 , n273316 , n55146 );
nand ( n273323 , n273321 , n273322 );
nand ( n273324 , n261585 , n29782 );
nand ( n273325 , n273318 , n273323 , n273324 );
buf ( n273326 , n273325 );
nand ( n273327 , n270557 , n270548 );
or ( n273328 , n257973 , n273327 );
not ( n273329 , n257966 );
not ( n273330 , n270548 );
or ( n273331 , n273329 , n273330 );
nor ( n273332 , n270557 , n219702 );
nand ( n273333 , n273331 , n273332 );
nand ( n273334 , n246217 , n204368 );
nand ( n273335 , n273328 , n273333 , n273334 );
buf ( n273336 , n273335 );
buf ( n273337 , n222908 );
not ( n273338 , n273337 );
not ( n273339 , n253557 );
or ( n273340 , n273338 , n273339 );
or ( n273341 , n253557 , n273337 );
nand ( n273342 , n273340 , n273341 );
and ( n273343 , n273342 , n264101 );
not ( n273344 , n273342 );
and ( n273345 , n273344 , n264098 );
nor ( n273346 , n273343 , n273345 );
nor ( n273347 , n273346 , n243434 );
not ( n273348 , n253050 );
not ( n273349 , n244704 );
or ( n273350 , n273348 , n273349 );
not ( n273351 , n253050 );
nand ( n273352 , n273351 , n244711 );
nand ( n273353 , n273350 , n273352 );
and ( n273354 , n273353 , n244769 );
not ( n273355 , n273353 );
and ( n273356 , n273355 , n244778 );
nor ( n273357 , n273354 , n273356 );
nand ( n273358 , n273347 , n273357 );
not ( n273359 , n273346 );
nor ( n273360 , n273359 , n260567 );
not ( n273361 , n255596 );
buf ( n273362 , n248099 );
not ( n273363 , n273362 );
not ( n273364 , n255589 );
or ( n273365 , n273363 , n273364 );
or ( n273366 , n256901 , n273362 );
nand ( n273367 , n273365 , n273366 );
not ( n273368 , n273367 );
or ( n273369 , n273361 , n273368 );
or ( n273370 , n273367 , n255596 );
nand ( n273371 , n273369 , n273370 );
nor ( n273372 , n273357 , n273371 );
nand ( n273373 , n273360 , n273372 );
not ( n273374 , n273357 );
nor ( n273375 , n273374 , n234021 );
nand ( n273376 , n273375 , n273371 );
nand ( n273377 , n239240 , n29121 );
nand ( n273378 , n273358 , n273373 , n273376 , n273377 );
buf ( n273379 , n273378 );
buf ( n273380 , n46105 );
not ( n273381 , n273380 );
not ( n273382 , n231952 );
or ( n273383 , n273381 , n273382 );
or ( n273384 , n231952 , n273380 );
nand ( n273385 , n273383 , n273384 );
and ( n273386 , n273385 , n264882 );
not ( n273387 , n273385 );
and ( n273388 , n273387 , n264879 );
nor ( n273389 , n273386 , n273388 );
not ( n273390 , n273389 );
nand ( n273391 , n273390 , n253902 );
not ( n273392 , n40957 );
not ( n273393 , n54263 );
or ( n273394 , n273392 , n273393 );
nand ( n273395 , n54273 , n40956 );
nand ( n273396 , n273394 , n273395 );
and ( n273397 , n273396 , n255321 );
not ( n273398 , n273396 );
and ( n273399 , n273398 , n255324 );
nor ( n273400 , n273397 , n273399 );
not ( n273401 , n273400 );
not ( n273402 , n258987 );
nand ( n273403 , n273401 , n273402 );
or ( n273404 , n273391 , n273403 );
not ( n273405 , n273402 );
not ( n273406 , n273390 );
or ( n273407 , n273405 , n273406 );
nor ( n273408 , n273401 , n250909 );
nand ( n273409 , n273407 , n273408 );
nand ( n273410 , n241976 , n33114 );
nand ( n273411 , n273404 , n273409 , n273410 );
buf ( n273412 , n273411 );
buf ( n273413 , n28244 );
buf ( n273414 , n34293 );
nand ( n273415 , n251379 , n226010 );
not ( n273416 , n229020 );
not ( n273417 , n255808 );
or ( n273418 , n273416 , n273417 );
not ( n273419 , n229020 );
nand ( n273420 , n273419 , n256762 );
nand ( n273421 , n273418 , n273420 );
and ( n273422 , n273421 , n256765 );
not ( n273423 , n273421 );
and ( n273424 , n273423 , n256768 );
nor ( n273425 , n273422 , n273424 );
not ( n273426 , n236982 );
not ( n273427 , n239298 );
or ( n273428 , n273426 , n273427 );
not ( n273429 , n236982 );
nand ( n273430 , n273429 , n239297 );
nand ( n273431 , n273428 , n273430 );
and ( n273432 , n273431 , n239399 );
not ( n273433 , n273431 );
and ( n273434 , n273433 , n239391 );
nor ( n273435 , n273432 , n273434 );
not ( n273436 , n273435 );
nand ( n273437 , n273425 , n273436 );
or ( n273438 , n273415 , n273437 );
nand ( n273439 , n251380 , n273437 );
nand ( n273440 , n236798 , n28103 );
nand ( n273441 , n273438 , n273439 , n273440 );
buf ( n273442 , n273441 );
buf ( n273443 , n28333 );
not ( n273444 , n32203 );
not ( n273445 , n255116 );
or ( n273446 , n273444 , n273445 );
not ( n273447 , n253287 );
not ( n273448 , n243153 );
not ( n273449 , n248677 );
not ( n273450 , n273449 );
or ( n273451 , n273448 , n273450 );
not ( n273452 , n243153 );
nand ( n273453 , n273452 , n253293 );
nand ( n273454 , n273451 , n273453 );
not ( n273455 , n273454 );
or ( n273456 , n273447 , n273455 );
or ( n273457 , n253287 , n273454 );
nand ( n273458 , n273456 , n273457 );
nand ( n273459 , n44766 , n273458 );
and ( n273460 , n273459 , n254999 );
not ( n273461 , n273459 );
and ( n273462 , n273461 , n44327 );
nor ( n273463 , n273460 , n273462 );
or ( n273464 , n273463 , n35816 );
nand ( n273465 , n273446 , n273464 );
buf ( n273466 , n273465 );
not ( n273467 , n230765 );
nand ( n273468 , n266648 , n262314 );
or ( n273469 , n273467 , n273468 );
not ( n273470 , n262314 );
not ( n273471 , n230205 );
not ( n273472 , n273471 );
or ( n273473 , n273470 , n273472 );
nor ( n273474 , n266648 , n265700 );
nand ( n273475 , n273473 , n273474 );
nand ( n273476 , n41944 , n31099 );
nand ( n273477 , n273469 , n273475 , n273476 );
buf ( n273478 , n273477 );
nand ( n273479 , n262688 , n256957 );
not ( n273480 , n272438 );
nand ( n273481 , n272449 , n273480 );
or ( n273482 , n273479 , n273481 );
nor ( n273483 , n262688 , n253358 );
nand ( n273484 , n273483 , n273481 );
nand ( n273485 , n35431 , n39902 );
nand ( n273486 , n273482 , n273484 , n273485 );
buf ( n273487 , n273486 );
not ( n273488 , RI19acf428_2216);
or ( n273489 , n233507 , n273488 );
not ( n273490 , RI19ac69e0_2280);
or ( n273491 , n226822 , n273490 );
nand ( n273492 , n273489 , n273491 );
buf ( n273493 , n273492 );
not ( n273494 , RI19acc020_2239);
or ( n273495 , n25328 , n273494 );
or ( n273496 , n226822 , n263463 );
nand ( n273497 , n273495 , n273496 );
buf ( n273498 , n273497 );
not ( n273499 , RI19ac5540_2289);
or ( n273500 , n233507 , n273499 );
or ( n273501 , n226822 , n266212 );
nand ( n273502 , n273500 , n273501 );
buf ( n273503 , n273502 );
nor ( n273504 , n263644 , n263655 );
or ( n273505 , n260376 , n273504 );
nor ( n273506 , n260374 , n239237 );
nand ( n273507 , n273506 , n273504 );
nand ( n273508 , n31576 , n25990 );
nand ( n273509 , n273505 , n273507 , n273508 );
buf ( n273510 , n273509 );
not ( n273511 , n268855 );
nand ( n273512 , n251785 , n273511 );
not ( n273513 , n242959 );
not ( n273514 , n273513 );
not ( n273515 , n245929 );
or ( n273516 , n273514 , n273515 );
not ( n273517 , n273513 );
nand ( n273518 , n273517 , n245918 );
nand ( n273519 , n273516 , n273518 );
and ( n273520 , n273519 , n256191 );
not ( n273521 , n273519 );
and ( n273522 , n273521 , n266168 );
nor ( n273523 , n273520 , n273522 );
nor ( n273524 , n273523 , n235050 );
not ( n273525 , n273524 );
or ( n273526 , n273512 , n273525 );
not ( n273527 , n273523 );
nand ( n273528 , n273527 , n273511 );
nand ( n273529 , n273528 , n251786 , n241459 );
nand ( n273530 , n46083 , n36599 );
nand ( n273531 , n273526 , n273529 , n273530 );
buf ( n273532 , n273531 );
nand ( n273533 , n270590 , n226010 );
not ( n273534 , n230478 );
not ( n273535 , n258610 );
or ( n273536 , n273534 , n273535 );
not ( n273537 , n230478 );
nand ( n273538 , n273537 , n271722 );
nand ( n273539 , n273536 , n273538 );
and ( n273540 , n273539 , n258622 );
not ( n273541 , n273539 );
and ( n273542 , n273541 , n258618 );
nor ( n273543 , n273540 , n273542 );
nand ( n273544 , n273543 , n270605 );
or ( n273545 , n273533 , n273544 );
not ( n273546 , n270605 );
not ( n273547 , n270590 );
or ( n273548 , n273546 , n273547 );
nor ( n273549 , n273543 , n226003 );
nand ( n273550 , n273548 , n273549 );
nand ( n273551 , n234448 , n32043 );
nand ( n273552 , n273545 , n273550 , n273551 );
buf ( n273553 , n273552 );
not ( n273554 , n205403 );
not ( n273555 , n55760 );
or ( n273556 , n273554 , n273555 );
buf ( n273557 , n243971 );
not ( n273558 , n273557 );
not ( n273559 , n252317 );
or ( n273560 , n273558 , n273559 );
or ( n273561 , n252317 , n273557 );
nand ( n273562 , n273560 , n273561 );
and ( n273563 , n273562 , n252324 );
not ( n273564 , n273562 );
and ( n273565 , n273564 , n252327 );
nor ( n273566 , n273563 , n273565 );
nand ( n273567 , n273238 , n273566 );
and ( n273568 , n273567 , n273259 );
not ( n273569 , n273567 );
and ( n273570 , n273569 , n273262 );
nor ( n273571 , n273568 , n273570 );
or ( n273572 , n273571 , n39763 );
nand ( n273573 , n273556 , n273572 );
buf ( n273574 , n273573 );
not ( n273575 , n259069 );
nand ( n273576 , n273575 , n259082 );
or ( n273577 , n266190 , n273576 );
nor ( n273578 , n266189 , n236795 );
nand ( n273579 , n273578 , n273576 );
nand ( n273580 , n246217 , n204606 );
nand ( n273581 , n273577 , n273579 , n273580 );
buf ( n273582 , n273581 );
not ( n273583 , RI19aa3058_2545);
or ( n273584 , n226819 , n273583 );
not ( n273585 , RI19a99698_2616);
or ( n273586 , n25335 , n273585 );
nand ( n273587 , n273584 , n273586 );
buf ( n273588 , n273587 );
not ( n273589 , n252976 );
not ( n273590 , n233271 );
or ( n273591 , n273589 , n273590 );
not ( n273592 , n252976 );
nand ( n273593 , n273592 , n233264 );
nand ( n273594 , n273591 , n273593 );
and ( n273595 , n273594 , n266838 );
not ( n273596 , n273594 );
and ( n273597 , n273596 , n266835 );
nor ( n273598 , n273595 , n273597 );
not ( n273599 , n273598 );
nand ( n273600 , n273599 , n257746 );
or ( n273601 , n257760 , n273600 );
nand ( n273602 , n257746 , n257759 );
nand ( n273603 , n273602 , n273598 , n235051 );
nand ( n273604 , n31576 , n25408 );
nand ( n273605 , n273601 , n273603 , n273604 );
buf ( n273606 , n273605 );
or ( n273607 , n233507 , n263465 );
not ( n273608 , RI19ab0a50_2449);
or ( n273609 , n25335 , n273608 );
nand ( n273610 , n273607 , n273609 );
buf ( n273611 , n273610 );
buf ( n273612 , n25907 );
not ( n273613 , n235008 );
not ( n273614 , n228280 );
not ( n273615 , n35804 );
or ( n273616 , n273614 , n273615 );
nand ( n273617 , n35811 , n228281 );
nand ( n273618 , n273616 , n273617 );
not ( n273619 , n273618 );
or ( n273620 , n273613 , n273619 );
or ( n273621 , n273618 , n253336 );
nand ( n273622 , n273620 , n273621 );
nor ( n273623 , n273622 , n40465 );
not ( n273624 , n248876 );
not ( n273625 , n237340 );
or ( n273626 , n273624 , n273625 );
not ( n273627 , n248876 );
nand ( n273628 , n273627 , n237350 );
nand ( n273629 , n273626 , n273628 );
and ( n273630 , n273629 , n256279 );
not ( n273631 , n273629 );
and ( n273632 , n273631 , n256280 );
nor ( n273633 , n273630 , n273632 );
not ( n273634 , n273633 );
nor ( n273635 , n273634 , n235732 );
nor ( n273636 , n273623 , n273635 );
not ( n273637 , n244857 );
not ( n273638 , n53657 );
or ( n273639 , n273637 , n273638 );
not ( n273640 , n244857 );
nand ( n273641 , n273640 , n231421 );
nand ( n273642 , n273639 , n273641 );
and ( n273643 , n273642 , n53665 );
not ( n273644 , n273642 );
and ( n273645 , n273644 , n34439 );
nor ( n273646 , n273643 , n273645 );
not ( n273647 , n273646 );
or ( n273648 , n273636 , n273647 );
nor ( n273649 , n273633 , n243434 );
and ( n273650 , n273649 , n273622 , n273647 );
not ( n273651 , n37976 );
nor ( n273652 , n273651 , n263991 );
nor ( n273653 , n273650 , n273652 );
nand ( n273654 , n273648 , n273653 );
buf ( n273655 , n273654 );
buf ( n273656 , n29366 );
not ( n273657 , n226596 );
not ( n273658 , n44324 );
or ( n273659 , n273657 , n273658 );
or ( n273660 , n44324 , n226596 );
nand ( n273661 , n273659 , n273660 );
not ( n273662 , n273661 );
not ( n273663 , n266084 );
and ( n273664 , n273662 , n273663 );
and ( n273665 , n273661 , n266084 );
nor ( n273666 , n273664 , n273665 );
nand ( n273667 , n273666 , n205649 );
not ( n273668 , n239621 );
not ( n273669 , n237746 );
or ( n273670 , n273668 , n273669 );
not ( n273671 , n239621 );
nand ( n273672 , n273671 , n262738 );
nand ( n273673 , n273670 , n273672 );
and ( n273674 , n273673 , n249482 );
not ( n273675 , n273673 );
and ( n273676 , n273675 , n36730 );
nor ( n273677 , n273674 , n273676 );
not ( n273678 , n273677 );
nand ( n273679 , n273678 , n258876 );
or ( n273680 , n273667 , n273679 );
nor ( n273681 , n273666 , n234110 );
nand ( n273682 , n273681 , n273679 );
nand ( n273683 , n234453 , n34846 );
nand ( n273684 , n273680 , n273682 , n273683 );
buf ( n273685 , n273684 );
not ( n273686 , RI19a9bd80_2599);
or ( n273687 , n25328 , n273686 );
not ( n273688 , RI19a919e8_2671);
or ( n273689 , n25335 , n273688 );
nand ( n273690 , n273687 , n273689 );
buf ( n273691 , n273690 );
not ( n273692 , RI19aa6640_2520);
or ( n273693 , n25328 , n273692 );
not ( n273694 , RI19a9ce60_2591);
or ( n273695 , n226822 , n273694 );
nand ( n273696 , n273693 , n273695 );
buf ( n273697 , n273696 );
not ( n273698 , n270245 );
not ( n273699 , n239379 );
not ( n273700 , n252917 );
or ( n273701 , n273699 , n273700 );
not ( n273702 , n239379 );
nand ( n273703 , n273702 , n252922 );
nand ( n273704 , n273701 , n273703 );
and ( n273705 , n273704 , n258058 );
not ( n273706 , n273704 );
and ( n273707 , n273706 , n258061 );
nor ( n273708 , n273705 , n273707 );
nor ( n273709 , n273708 , n258280 );
nand ( n273710 , n273698 , n273709 , n270256 );
not ( n273711 , n273708 );
nand ( n273712 , n273711 , n270256 );
nand ( n273713 , n273712 , n270245 , n237385 );
nand ( n273714 , n31577 , n26065 );
nand ( n273715 , n273710 , n273713 , n273714 );
buf ( n273716 , n273715 );
nand ( n273717 , n272581 , n272592 );
or ( n273718 , n233974 , n273717 );
not ( n273719 , n233970 );
not ( n273720 , n272581 );
or ( n273721 , n273719 , n273720 );
nor ( n273722 , n272592 , n234021 );
nand ( n273723 , n273721 , n273722 );
nand ( n273724 , n245701 , n28499 );
nand ( n273725 , n273718 , n273723 , n273724 );
buf ( n273726 , n273725 );
not ( n273727 , RI19a8d230_2703);
or ( n273728 , n233507 , n273727 );
not ( n273729 , RI19acd5b0_2229);
or ( n273730 , n25335 , n273729 );
nand ( n273731 , n273728 , n273730 );
buf ( n273732 , n273731 );
or ( n273733 , n25328 , n254436 );
or ( n273734 , n25335 , n254422 );
nand ( n273735 , n273733 , n273734 );
buf ( n273736 , n273735 );
or ( n273737 , n233507 , n262674 );
not ( n273738 , RI19a8b4a8_2716);
or ( n273739 , n25335 , n273738 );
nand ( n273740 , n273737 , n273739 );
buf ( n273741 , n273740 );
or ( n273742 , n233507 , n266242 );
or ( n273743 , n25336 , n261957 );
nand ( n273744 , n273742 , n273743 );
buf ( n273745 , n273744 );
not ( n273746 , n244228 );
not ( n273747 , n28929 );
or ( n273748 , n273746 , n273747 );
not ( n273749 , n244228 );
nand ( n273750 , n273749 , n28936 );
nand ( n273751 , n273748 , n273750 );
and ( n273752 , n273751 , n29962 );
not ( n273753 , n273751 );
and ( n273754 , n273753 , n29965 );
nor ( n273755 , n273752 , n273754 );
nand ( n273756 , n262461 , n273755 );
nand ( n273757 , n258455 , n250111 );
or ( n273758 , n273756 , n273757 );
nand ( n273759 , n258456 , n273756 );
nand ( n273760 , n238114 , n28244 );
nand ( n273761 , n273758 , n273759 , n273760 );
buf ( n273762 , n273761 );
nand ( n273763 , n256581 , n267281 );
or ( n273764 , n273763 , n256585 );
nor ( n273765 , n256229 , n240080 );
nand ( n273766 , n273763 , n273765 );
nand ( n273767 , n251717 , n31057 );
nand ( n273768 , n273764 , n273766 , n273767 );
buf ( n273769 , n273768 );
nand ( n273770 , n42442 , n259009 );
not ( n273771 , n250234 );
buf ( n273772 , n254713 );
not ( n273773 , n273772 );
not ( n273774 , n273773 );
not ( n273775 , n249610 );
or ( n273776 , n273774 , n273775 );
nand ( n273777 , n249600 , n273772 );
nand ( n273778 , n273776 , n273777 );
not ( n273779 , n273778 );
or ( n273780 , n273771 , n273779 );
or ( n273781 , n250234 , n273778 );
nand ( n273782 , n273780 , n273781 );
not ( n273783 , n273782 );
nand ( n273784 , n221272 , n273783 );
or ( n273785 , n273770 , n273784 );
not ( n273786 , n221272 );
not ( n273787 , n42442 );
or ( n273788 , n273786 , n273787 );
nor ( n273789 , n273783 , n35816 );
nand ( n273790 , n273788 , n273789 );
nand ( n273791 , n252711 , n34362 );
nand ( n273792 , n273785 , n273790 , n273791 );
buf ( n273793 , n273792 );
not ( n273794 , RI19acd808_2228);
or ( n273795 , n25328 , n273794 );
or ( n273796 , n25335 , n262667 );
nand ( n273797 , n273795 , n273796 );
buf ( n273798 , n273797 );
not ( n273799 , n30954 );
not ( n273800 , n246963 );
or ( n273801 , n273799 , n273800 );
not ( n273802 , n30954 );
nand ( n273803 , n273802 , n246968 );
nand ( n273804 , n273801 , n273803 );
and ( n273805 , n273804 , n247019 );
not ( n273806 , n273804 );
and ( n273807 , n273806 , n247014 );
nor ( n273808 , n273805 , n273807 );
not ( n273809 , n273808 );
not ( n273810 , n252964 );
not ( n273811 , n273810 );
not ( n273812 , n233271 );
or ( n273813 , n273811 , n273812 );
not ( n273814 , n273810 );
nand ( n273815 , n273814 , n233264 );
nand ( n273816 , n273813 , n273815 );
and ( n273817 , n273816 , n266838 );
not ( n273818 , n273816 );
and ( n273819 , n273818 , n266835 );
nor ( n273820 , n273817 , n273819 );
not ( n273821 , n273820 );
nand ( n273822 , n273809 , n273821 );
not ( n273823 , n247075 );
not ( n273824 , n273823 );
not ( n273825 , n253578 );
or ( n273826 , n273824 , n273825 );
or ( n273827 , n253464 , n273823 );
nand ( n273828 , n273826 , n273827 );
and ( n273829 , n273828 , n253475 );
not ( n273830 , n273828 );
and ( n273831 , n273830 , n253478 );
nor ( n273832 , n273829 , n273831 );
nand ( n273833 , n273832 , n245241 );
or ( n273834 , n273822 , n273833 );
nor ( n273835 , n273832 , n247698 );
nand ( n273836 , n273822 , n273835 );
nand ( n273837 , n246460 , n28324 );
nand ( n273838 , n273834 , n273836 , n273837 );
buf ( n273839 , n273838 );
buf ( n273840 , n29144 );
not ( n273841 , RI19a9aac0_2607);
or ( n273842 , n25328 , n273841 );
not ( n273843 , RI19a90a70_2678);
or ( n273844 , n25336 , n273843 );
nand ( n273845 , n273842 , n273844 );
buf ( n273846 , n273845 );
not ( n273847 , RI1754af90_50);
or ( n273848 , n249126 , n273847 );
not ( n273849 , n258658 );
not ( n273850 , n273849 );
nand ( n273851 , n259432 , RI1754a5b8_71);
not ( n273852 , n273851 );
and ( n273853 , n273850 , n273852 );
and ( n273854 , n244606 , n32818 );
nor ( n273855 , n273853 , n273854 );
nand ( n273856 , n273848 , n273855 );
buf ( n273857 , n273856 );
not ( n273858 , n245213 );
not ( n273859 , n272892 );
nand ( n273860 , n273858 , n273859 );
or ( n273861 , n270460 , n273860 );
not ( n273862 , n273859 );
not ( n273863 , n270459 );
or ( n273864 , n273862 , n273863 );
not ( n273865 , n270449 );
nand ( n273866 , n273864 , n273865 );
nand ( n273867 , n247744 , n32191 );
nand ( n273868 , n273861 , n273866 , n273867 );
buf ( n273869 , n273868 );
or ( n273870 , n233507 , n271870 );
not ( n273871 , RI19aa7090_2516);
or ( n273872 , n25335 , n273871 );
nand ( n273873 , n273870 , n273872 );
buf ( n273874 , n273873 );
buf ( n273875 , n37890 );
buf ( n273876 , n40547 );
buf ( n273877 , n35001 );
not ( n273878 , n230453 );
not ( n273879 , n258610 );
or ( n273880 , n273878 , n273879 );
not ( n273881 , n230453 );
nand ( n273882 , n273881 , n271722 );
nand ( n273883 , n273880 , n273882 );
and ( n273884 , n273883 , n258618 );
not ( n273885 , n273883 );
and ( n273886 , n273885 , n258622 );
nor ( n273887 , n273884 , n273886 );
nand ( n273888 , n273887 , n235051 );
nand ( n273889 , n264513 , n264523 );
or ( n273890 , n273888 , n273889 );
not ( n273891 , n264523 );
not ( n273892 , n273887 );
or ( n273893 , n273891 , n273892 );
nor ( n273894 , n264513 , n236795 );
nand ( n273895 , n273893 , n273894 );
nand ( n273896 , n256673 , n44128 );
nand ( n273897 , n273890 , n273895 , n273896 );
buf ( n273898 , n273897 );
not ( n273899 , n267987 );
nand ( n273900 , n267959 , n254528 );
not ( n273901 , n273900 );
or ( n273902 , n273899 , n273901 );
not ( n273903 , n242069 );
not ( n273904 , n239724 );
not ( n273905 , n239107 );
or ( n273906 , n273904 , n273905 );
nand ( n273907 , n239099 , n239723 );
nand ( n273908 , n273906 , n273907 );
not ( n273909 , n273908 );
or ( n273910 , n273903 , n273909 );
or ( n273911 , n242069 , n273908 );
nand ( n273912 , n273910 , n273911 );
nand ( n273913 , n273902 , n273912 );
nor ( n273914 , n267959 , n235732 );
nor ( n273915 , n267970 , n273912 );
and ( n273916 , n273914 , n273915 );
and ( n273917 , n251717 , n204732 );
nor ( n273918 , n273916 , n273917 );
nand ( n273919 , n273913 , n273918 );
buf ( n273920 , n273919 );
not ( n273921 , RI19acdcb8_2226);
or ( n273922 , n226819 , n273921 );
not ( n273923 , RI19ac5108_2291);
or ( n273924 , n25336 , n273923 );
nand ( n273925 , n273922 , n273924 );
buf ( n273926 , n273925 );
not ( n273927 , n232053 );
not ( n273928 , n51342 );
or ( n273929 , n273927 , n273928 );
not ( n273930 , n232053 );
nand ( n273931 , n273930 , n51336 );
nand ( n273932 , n273929 , n273931 );
and ( n273933 , n273932 , n251488 );
not ( n273934 , n273932 );
and ( n273935 , n273934 , n51349 );
nor ( n273936 , n273933 , n273935 );
nor ( n273937 , n266549 , n273936 );
nand ( n273938 , n272115 , n273937 );
not ( n273939 , n272114 );
not ( n273940 , n273936 );
nand ( n273941 , n273939 , n273940 );
nand ( n273942 , n273941 , n266549 , n245241 );
nand ( n273943 , n37728 , n29111 );
nand ( n273944 , n273938 , n273942 , n273943 );
buf ( n273945 , n273944 );
not ( n273946 , n54646 );
not ( n273947 , n257703 );
or ( n273948 , n273946 , n273947 );
not ( n273949 , n54646 );
nand ( n273950 , n273949 , n245517 );
nand ( n273951 , n273948 , n273950 );
and ( n273952 , n273951 , n245524 );
not ( n273953 , n273951 );
and ( n273954 , n273953 , n268159 );
nor ( n273955 , n273952 , n273954 );
not ( n273956 , n273955 );
not ( n273957 , n260594 );
nand ( n273958 , n273956 , n273957 );
or ( n273959 , n260584 , n273958 );
nor ( n273960 , n260583 , n40465 );
nand ( n273961 , n273960 , n273958 );
nand ( n273962 , n244840 , n28622 );
nand ( n273963 , n273959 , n273961 , n273962 );
buf ( n273964 , n273963 );
nand ( n273965 , n271457 , n205649 );
not ( n273966 , n252617 );
not ( n273967 , n253264 );
or ( n273968 , n273966 , n273967 );
not ( n273969 , n252617 );
nand ( n273970 , n273969 , n253271 );
nand ( n273971 , n273968 , n273970 );
and ( n273972 , n273971 , n232899 );
not ( n273973 , n273971 );
and ( n273974 , n273973 , n232900 );
nor ( n273975 , n273972 , n273974 );
not ( n273976 , n273975 );
nand ( n273977 , n271469 , n273976 );
or ( n273978 , n273965 , n273977 );
not ( n273979 , n271469 );
not ( n273980 , n271457 );
or ( n273981 , n273979 , n273980 );
nor ( n273982 , n273976 , n219702 );
nand ( n273983 , n273981 , n273982 );
nand ( n273984 , n51381 , n36514 );
nand ( n273985 , n273978 , n273983 , n273984 );
buf ( n273986 , n273985 );
not ( n273987 , RI19aaf448_2459);
or ( n273988 , n226819 , n273987 );
not ( n273989 , RI19a82b50_2775);
or ( n273990 , n25335 , n273989 );
nand ( n273991 , n273988 , n273990 );
buf ( n273992 , n273991 );
nand ( n273993 , n257822 , n257845 );
not ( n273994 , n263910 );
or ( n273995 , n273993 , n273994 );
nor ( n273996 , n263904 , n249531 );
nand ( n273997 , n273993 , n273996 );
nand ( n273998 , n31577 , n221738 );
nand ( n273999 , n273995 , n273997 , n273998 );
buf ( n274000 , n273999 );
not ( n274001 , n243331 );
not ( n274002 , n250811 );
or ( n274003 , n274001 , n274002 );
not ( n274004 , n250805 );
or ( n274005 , n274004 , n243331 );
nand ( n274006 , n274003 , n274005 );
and ( n274007 , n274006 , n257382 );
not ( n274008 , n274006 );
and ( n274009 , n274008 , n270150 );
nor ( n274010 , n274007 , n274009 );
buf ( n274011 , n45475 );
not ( n274012 , n274011 );
not ( n274013 , n248154 );
or ( n274014 , n274012 , n274013 );
not ( n274015 , n274011 );
nand ( n274016 , n274015 , n248161 );
nand ( n274017 , n274014 , n274016 );
and ( n274018 , n274017 , n248211 );
not ( n274019 , n274017 );
and ( n274020 , n274019 , n248220 );
nor ( n274021 , n274018 , n274020 );
nor ( n274022 , n274010 , n274021 );
or ( n274023 , n267122 , n274022 );
nor ( n274024 , n267121 , n221279 );
nand ( n274025 , n274024 , n274022 );
nand ( n274026 , n39766 , n204862 );
nand ( n274027 , n274023 , n274025 , n274026 );
buf ( n274028 , n274027 );
not ( n274029 , RI19a876c8_2742);
or ( n274030 , n25328 , n274029 );
or ( n274031 , n25335 , n256419 );
nand ( n274032 , n274030 , n274031 );
buf ( n274033 , n274032 );
not ( n274034 , RI19a82d30_2774);
or ( n274035 , n25328 , n274034 );
or ( n274036 , n25336 , n260901 );
nand ( n274037 , n274035 , n274036 );
buf ( n274038 , n274037 );
buf ( n274039 , n33131 );
not ( n274040 , RI19aae458_2466);
or ( n274041 , n25328 , n274040 );
not ( n274042 , RI19aa3ee0_2538);
or ( n274043 , n226822 , n274042 );
nand ( n274044 , n274041 , n274043 );
buf ( n274045 , n274044 );
buf ( n274046 , n220535 );
not ( n274047 , n273425 );
nand ( n274048 , n274047 , n251456 );
or ( n274049 , n273415 , n274048 );
not ( n274050 , n274047 );
not ( n274051 , n251379 );
or ( n274052 , n274050 , n274051 );
nor ( n274053 , n251456 , n49051 );
nand ( n274054 , n274052 , n274053 );
nand ( n274055 , n35431 , n25419 );
nand ( n274056 , n274049 , n274054 , n274055 );
buf ( n274057 , n274056 );
not ( n274058 , n248765 );
nand ( n274059 , n274058 , n255961 );
not ( n274060 , n270835 );
or ( n274061 , n274059 , n274060 );
nand ( n274062 , n274059 , n270939 );
nand ( n274063 , n39766 , n42738 );
nand ( n274064 , n274061 , n274062 , n274063 );
buf ( n274065 , n274064 );
not ( n274066 , n270900 );
not ( n274067 , n274066 );
not ( n274068 , n270916 );
or ( n274069 , n274067 , n274068 );
not ( n274070 , n268754 );
nor ( n274071 , n274070 , n234818 );
nand ( n274072 , n274069 , n274071 );
nor ( n274073 , n270900 , n268754 );
nand ( n274074 , n270913 , n274073 );
nand ( n274075 , n246460 , n208672 );
nand ( n274076 , n274072 , n274074 , n274075 );
buf ( n274077 , n274076 );
not ( n274078 , n272909 );
not ( n274079 , n244003 );
not ( n274080 , n274079 );
not ( n274081 , n252318 );
or ( n274082 , n274080 , n274081 );
or ( n274083 , n252321 , n274079 );
nand ( n274084 , n274082 , n274083 );
and ( n274085 , n274084 , n252324 );
not ( n274086 , n274084 );
and ( n274087 , n274086 , n252327 );
nor ( n274088 , n274085 , n274087 );
nor ( n274089 , n262438 , n274088 );
or ( n274090 , n274078 , n274089 );
nor ( n274091 , n272914 , n236795 );
nand ( n274092 , n274091 , n274089 );
nand ( n274093 , n234448 , n216717 );
nand ( n274094 , n274090 , n274092 , n274093 );
buf ( n274095 , n274094 );
not ( n274096 , n40538 );
not ( n274097 , n245701 );
or ( n274098 , n274096 , n274097 );
nand ( n274099 , n271112 , n257333 );
not ( n274100 , n274099 );
not ( n274101 , n251550 );
and ( n274102 , n274100 , n274101 );
and ( n274103 , n274099 , n251550 );
nor ( n274104 , n274102 , n274103 );
or ( n274105 , n274104 , n261009 );
nand ( n274106 , n274098 , n274105 );
buf ( n274107 , n274106 );
buf ( n274108 , n29043 );
buf ( n274109 , n25408 );
not ( n274110 , RI19abe2e0_2348);
or ( n274111 , n25328 , n274110 );
not ( n274112 , RI19a843b0_2764);
or ( n274113 , n226822 , n274112 );
nand ( n274114 , n274111 , n274113 );
buf ( n274115 , n274114 );
not ( n274116 , n36036 );
not ( n274117 , n234453 );
or ( n274118 , n274116 , n274117 );
not ( n274119 , n42200 );
not ( n274120 , n234305 );
or ( n274121 , n274119 , n274120 );
not ( n274122 , n42200 );
nand ( n274123 , n274122 , n234298 );
nand ( n274124 , n274121 , n274123 );
and ( n274125 , n274124 , n256932 );
not ( n274126 , n274124 );
and ( n274127 , n274126 , n256928 );
nor ( n274128 , n274125 , n274127 );
not ( n274129 , n274128 );
not ( n274130 , n251137 );
not ( n274131 , n242520 );
or ( n274132 , n274130 , n274131 );
not ( n274133 , n251137 );
nand ( n274134 , n274133 , n242527 );
nand ( n274135 , n274132 , n274134 );
and ( n274136 , n274135 , n242575 );
not ( n274137 , n274135 );
and ( n274138 , n274137 , n242571 );
nor ( n274139 , n274136 , n274138 );
nand ( n274140 , n274129 , n274139 );
buf ( n274141 , n236621 );
not ( n274142 , n274141 );
not ( n274143 , n43504 );
or ( n274144 , n274142 , n274143 );
or ( n274145 , n248066 , n274141 );
nand ( n274146 , n274144 , n274145 );
not ( n274147 , n274146 );
not ( n274148 , n268003 );
and ( n274149 , n274147 , n274148 );
and ( n274150 , n274146 , n268003 );
nor ( n274151 , n274149 , n274150 );
not ( n274152 , n274151 );
and ( n274153 , n274140 , n274152 );
not ( n274154 , n274140 );
and ( n274155 , n274154 , n274151 );
nor ( n274156 , n274153 , n274155 );
or ( n274157 , n274156 , n235052 );
nand ( n274158 , n274118 , n274157 );
buf ( n274159 , n274158 );
not ( n274160 , RI1754bda0_20);
or ( n274161 , n255977 , n274160 );
nand ( n274162 , n244606 , n35139 );
nand ( n274163 , n274161 , n274162 );
buf ( n274164 , n274163 );
or ( n274165 , n226819 , n273694 );
not ( n274166 , RI19a92bb8_2663);
or ( n274167 , n25335 , n274166 );
nand ( n274168 , n274165 , n274167 );
buf ( n274169 , n274168 );
not ( n274170 , n29811 );
not ( n274171 , n51381 );
or ( n274172 , n274170 , n274171 );
nand ( n274173 , n261310 , n261320 );
and ( n274174 , n274173 , n265309 );
not ( n274175 , n274173 );
and ( n274176 , n274175 , n265308 );
nor ( n274177 , n274174 , n274176 );
or ( n274178 , n274177 , n250068 );
nand ( n274179 , n274172 , n274178 );
buf ( n274180 , n274179 );
not ( n274181 , n47777 );
nor ( n274182 , n274181 , n245932 );
nand ( n274183 , n258419 , n274182 );
not ( n274184 , n245933 );
not ( n274185 , n48241 );
or ( n274186 , n274184 , n274185 );
nor ( n274187 , n47777 , n240080 );
nand ( n274188 , n274186 , n274187 );
nand ( n274189 , n245701 , n39836 );
nand ( n274190 , n274183 , n274188 , n274189 );
buf ( n274191 , n274190 );
or ( n274192 , n25328 , n269257 );
not ( n274193 , RI19ac1b98_2316);
or ( n274194 , n25335 , n274193 );
nand ( n274195 , n274192 , n274194 );
buf ( n274196 , n274195 );
not ( n274197 , n256799 );
nand ( n274198 , n256789 , n274197 );
or ( n274199 , n252874 , n274198 );
not ( n274200 , n252871 );
nand ( n274201 , n274200 , n254227 );
not ( n274202 , n274201 );
nand ( n274203 , n274202 , n274198 );
nand ( n274204 , n255116 , n205718 );
nand ( n274205 , n274199 , n274203 , n274204 );
buf ( n274206 , n274205 );
not ( n274207 , n25922 );
not ( n274208 , n234823 );
or ( n274209 , n274207 , n274208 );
nand ( n274210 , n35633 , n204518 , n245003 , n245839 );
not ( n274211 , n274210 );
not ( n274212 , n263055 );
or ( n274213 , n274211 , n274212 );
or ( n274214 , n263055 , n274210 );
nand ( n274215 , n274213 , n274214 );
not ( n274216 , n274215 );
not ( n274217 , n231945 );
not ( n274218 , n242380 );
or ( n274219 , n274217 , n274218 );
not ( n274220 , n231945 );
nand ( n274221 , n274220 , n242373 );
nand ( n274222 , n274219 , n274221 );
and ( n274223 , n274222 , n243660 );
not ( n274224 , n274222 );
and ( n274225 , n274224 , n243659 );
nor ( n274226 , n274223 , n274225 );
nor ( n274227 , n274226 , n263066 );
not ( n274228 , n274227 );
and ( n274229 , n274216 , n274228 );
and ( n274230 , n274215 , n274227 );
nor ( n274231 , n274229 , n274230 );
or ( n274232 , n274231 , n238223 );
nand ( n274233 , n274209 , n274232 );
buf ( n274234 , n274233 );
buf ( n274235 , n31192 );
not ( n274236 , n256272 );
nand ( n274237 , n274236 , n256284 );
or ( n274238 , n271523 , n274237 );
nand ( n274239 , n253720 , n274237 );
nand ( n274240 , n50615 , n37813 );
nand ( n274241 , n274238 , n274239 , n274240 );
buf ( n274242 , n274241 );
buf ( n274243 , n27903 );
not ( n274244 , n235469 );
not ( n274245 , n248135 );
or ( n274246 , n274244 , n274245 );
not ( n274247 , n235469 );
nand ( n274248 , n274247 , n248143 );
nand ( n274249 , n274246 , n274248 );
and ( n274250 , n274249 , n248146 );
not ( n274251 , n274249 );
and ( n274252 , n274251 , n248149 );
nor ( n274253 , n274250 , n274252 );
not ( n274254 , n274253 );
not ( n274255 , n274254 );
not ( n274256 , n252543 );
not ( n274257 , n249362 );
or ( n274258 , n274256 , n274257 );
not ( n274259 , n252543 );
nand ( n274260 , n274259 , n271683 );
nand ( n274261 , n274258 , n274260 );
and ( n274262 , n274261 , n261550 );
not ( n274263 , n274261 );
and ( n274264 , n274263 , n261547 );
nor ( n274265 , n274262 , n274264 );
nand ( n274266 , n274255 , n274265 );
or ( n274267 , n268400 , n274266 );
not ( n274268 , n274265 );
not ( n274269 , n268399 );
or ( n274270 , n274268 , n274269 );
nor ( n274271 , n274253 , n37725 );
nand ( n274272 , n274270 , n274271 );
nand ( n274273 , n35431 , n40393 );
nand ( n274274 , n274267 , n274272 , n274273 );
buf ( n274275 , n274274 );
buf ( n274276 , n30669 );
buf ( n274277 , n41384 );
or ( n274278 , n233507 , n268832 );
or ( n274279 , n25336 , n246464 );
nand ( n274280 , n274278 , n274279 );
buf ( n274281 , n274280 );
not ( n274282 , n249284 );
buf ( n274283 , n237581 );
not ( n274284 , n274283 );
not ( n274285 , n249276 );
or ( n274286 , n274284 , n274285 );
or ( n274287 , n263562 , n274283 );
nand ( n274288 , n274286 , n274287 );
not ( n274289 , n274288 );
or ( n274290 , n274282 , n274289 );
or ( n274291 , n274288 , n263568 );
nand ( n274292 , n274290 , n274291 );
nor ( n274293 , n274292 , n267386 );
nand ( n274294 , n267399 , n274293 );
not ( n274295 , n267386 );
nand ( n274296 , n274295 , n267397 );
not ( n274297 , n251190 );
nand ( n274298 , n274296 , n274292 , n274297 );
nand ( n274299 , n241068 , n28982 );
nand ( n274300 , n274294 , n274298 , n274299 );
buf ( n274301 , n274300 );
not ( n274302 , RI19a23150_2796);
or ( n274303 , n25328 , n274302 );
not ( n274304 , RI19a864f8_2750);
or ( n274305 , n226822 , n274304 );
nand ( n274306 , n274303 , n274305 );
buf ( n274307 , n274306 );
nand ( n274308 , n256403 , n252224 , n271922 );
not ( n274309 , n256397 );
nand ( n274310 , n274309 , n271922 );
not ( n274311 , n252358 );
nand ( n274312 , n274310 , n252225 , n274311 );
nand ( n274313 , n37728 , n34630 );
nand ( n274314 , n274308 , n274312 , n274313 );
buf ( n274315 , n274314 );
not ( n274316 , n267365 );
not ( n274317 , n238728 );
not ( n274318 , n247991 );
or ( n274319 , n274317 , n274318 );
not ( n274320 , n238728 );
nand ( n274321 , n274320 , n247999 );
nand ( n274322 , n274319 , n274321 );
and ( n274323 , n274322 , n261862 );
not ( n274324 , n274322 );
and ( n274325 , n274324 , n261859 );
nor ( n274326 , n274323 , n274325 );
nand ( n274327 , n262382 , n274326 );
or ( n274328 , n274316 , n274327 );
not ( n274329 , n262382 );
not ( n274330 , n262358 );
not ( n274331 , n274330 );
or ( n274332 , n274329 , n274331 );
buf ( n274333 , n40465 );
nor ( n274334 , n274326 , n274333 );
nand ( n274335 , n274332 , n274334 );
nand ( n274336 , n31577 , n28783 );
nand ( n274337 , n274328 , n274335 , n274336 );
buf ( n274338 , n274337 );
or ( n274339 , n25328 , n274042 );
not ( n274340 , RI19a9a868_2608);
or ( n274341 , n25336 , n274340 );
nand ( n274342 , n274339 , n274341 );
buf ( n274343 , n274342 );
not ( n274344 , RI19a94df0_2648);
or ( n274345 , n25328 , n274344 );
or ( n274346 , n25335 , n272731 );
nand ( n274347 , n274345 , n274346 );
buf ( n274348 , n274347 );
not ( n274349 , n241353 );
not ( n274350 , n245338 );
or ( n274351 , n274349 , n274350 );
or ( n274352 , n250708 , n241353 );
nand ( n274353 , n274351 , n274352 );
not ( n274354 , n274353 );
not ( n274355 , n245393 );
and ( n274356 , n274354 , n274355 );
and ( n274357 , n274353 , n253363 );
nor ( n274358 , n274356 , n274357 );
nor ( n274359 , n274358 , n50944 );
not ( n274360 , n274359 );
not ( n274361 , n236174 );
nand ( n274362 , n274361 , n236394 );
or ( n274363 , n274360 , n274362 );
not ( n274364 , n274361 );
not ( n274365 , n274358 );
not ( n274366 , n274365 );
or ( n274367 , n274364 , n274366 );
nand ( n274368 , n274367 , n265907 );
nand ( n274369 , n255116 , n32545 );
nand ( n274370 , n274363 , n274368 , n274369 );
buf ( n274371 , n274370 );
not ( n274372 , n38860 );
not ( n274373 , n51381 );
or ( n274374 , n274372 , n274373 );
not ( n274375 , n38636 );
nand ( n274376 , n274375 , n256102 );
and ( n274377 , n274376 , n55149 );
not ( n274378 , n274376 );
and ( n274379 , n274378 , n39757 );
nor ( n274380 , n274377 , n274379 );
or ( n274381 , n274380 , n238223 );
nand ( n274382 , n274374 , n274381 );
buf ( n274383 , n274382 );
not ( n274384 , n249665 );
not ( n274385 , n259590 );
or ( n274386 , n274384 , n274385 );
or ( n274387 , n248385 , n249665 );
nand ( n274388 , n274386 , n274387 );
and ( n274389 , n274388 , n255885 );
not ( n274390 , n274388 );
and ( n274391 , n274390 , n259595 );
nor ( n274392 , n274389 , n274391 );
not ( n274393 , n274392 );
nand ( n274394 , n274393 , n222532 );
not ( n274395 , n243835 );
not ( n274396 , n246705 );
or ( n274397 , n274395 , n274396 );
or ( n274398 , n246705 , n243835 );
nand ( n274399 , n274397 , n274398 );
not ( n274400 , n274399 );
not ( n274401 , n246768 );
or ( n274402 , n274400 , n274401 );
or ( n274403 , n246768 , n274399 );
nand ( n274404 , n274402 , n274403 );
not ( n274405 , n274404 );
not ( n274406 , n234405 );
not ( n274407 , n274406 );
not ( n274408 , n238106 );
or ( n274409 , n274407 , n274408 );
not ( n274410 , n274406 );
nand ( n274411 , n274410 , n238101 );
nand ( n274412 , n274409 , n274411 );
and ( n274413 , n274412 , n244390 );
not ( n274414 , n274412 );
and ( n274415 , n274414 , n244387 );
nor ( n274416 , n274413 , n274415 );
nand ( n274417 , n274405 , n274416 );
or ( n274418 , n274394 , n274417 );
not ( n274419 , n274405 );
not ( n274420 , n274393 );
or ( n274421 , n274419 , n274420 );
nor ( n274422 , n274416 , n221279 );
nand ( n274423 , n274421 , n274422 );
nand ( n274424 , n238638 , n204851 );
nand ( n274425 , n274418 , n274423 , n274424 );
buf ( n274426 , n274425 );
not ( n274427 , n34714 );
not ( n274428 , n234453 );
or ( n274429 , n274427 , n274428 );
nand ( n274430 , n244477 , n49193 );
and ( n274431 , n274430 , n260170 );
not ( n274432 , n274430 );
and ( n274433 , n274432 , n49629 );
nor ( n274434 , n274431 , n274433 );
or ( n274435 , n274434 , n244837 );
nand ( n274436 , n274429 , n274435 );
buf ( n274437 , n274436 );
not ( n274438 , n25857 );
not ( n274439 , n55760 );
or ( n274440 , n274438 , n274439 );
not ( n274441 , n256810 );
nand ( n274442 , n274441 , n252938 );
and ( n274443 , n274442 , n274197 );
not ( n274444 , n274442 );
and ( n274445 , n274444 , n256799 );
nor ( n274446 , n274443 , n274445 );
or ( n274447 , n274446 , n226003 );
nand ( n274448 , n274440 , n274447 );
buf ( n274449 , n274448 );
not ( n274450 , n249804 );
not ( n274451 , n272884 );
or ( n274452 , n274450 , n274451 );
nand ( n274453 , n51747 , n249805 );
nand ( n274454 , n274452 , n274453 );
and ( n274455 , n274454 , n51753 );
not ( n274456 , n274454 );
and ( n274457 , n274456 , n229518 );
nor ( n274458 , n274455 , n274457 );
nor ( n274459 , n273371 , n274458 );
nand ( n274460 , n273347 , n274459 );
not ( n274461 , n274458 );
nand ( n274462 , n273359 , n274461 );
nand ( n274463 , n274462 , n273371 , n246697 );
nand ( n274464 , n261585 , n34787 );
nand ( n274465 , n274460 , n274463 , n274464 );
buf ( n274466 , n274465 );
not ( n274467 , n45003 );
not ( n274468 , n274467 );
not ( n274469 , n244009 );
or ( n274470 , n274468 , n274469 );
or ( n274471 , n244459 , n274467 );
nand ( n274472 , n274470 , n274471 );
and ( n274473 , n274472 , n244056 );
not ( n274474 , n274472 );
and ( n274475 , n274474 , n257630 );
nor ( n274476 , n274473 , n274475 );
not ( n274477 , n274476 );
not ( n274478 , n254877 );
or ( n274479 , n274477 , n274478 );
not ( n274480 , n252603 );
not ( n274481 , n253264 );
or ( n274482 , n274480 , n274481 );
not ( n274483 , n252603 );
nand ( n274484 , n274483 , n253271 );
nand ( n274485 , n274482 , n274484 );
and ( n274486 , n274485 , n232900 );
not ( n274487 , n274485 );
not ( n274488 , n55135 );
and ( n274489 , n274487 , n274488 );
nor ( n274490 , n274486 , n274489 );
nor ( n274491 , n274490 , n234440 );
nand ( n274492 , n274479 , n274491 );
not ( n274493 , n274476 );
nor ( n274494 , n274493 , n52445 );
nand ( n274495 , n274494 , n254877 , n274490 );
nand ( n274496 , n245701 , n25463 );
nand ( n274497 , n274492 , n274495 , n274496 );
buf ( n274498 , n274497 );
not ( n274499 , n271332 );
nand ( n274500 , n274499 , n271352 );
not ( n274501 , n49908 );
not ( n274502 , n245862 );
or ( n274503 , n274501 , n274502 );
not ( n274504 , n49908 );
nand ( n274505 , n274504 , n245872 );
nand ( n274506 , n274503 , n274505 );
and ( n274507 , n274506 , n245920 );
not ( n274508 , n274506 );
and ( n274509 , n274508 , n245930 );
nor ( n274510 , n274507 , n274509 );
not ( n274511 , n274510 );
nor ( n274512 , n274511 , n244216 );
not ( n274513 , n274512 );
or ( n274514 , n274500 , n274513 );
nor ( n274515 , n274510 , n226004 );
nand ( n274516 , n274500 , n274515 );
nand ( n274517 , n41945 , n43611 );
nand ( n274518 , n274514 , n274516 , n274517 );
buf ( n274519 , n274518 );
not ( n274520 , n45207 );
not ( n274521 , n258213 );
or ( n274522 , n274520 , n274521 );
not ( n274523 , n244038 );
not ( n274524 , n54917 );
or ( n274525 , n274523 , n274524 );
not ( n274526 , n244038 );
nand ( n274527 , n274526 , n54926 );
nand ( n274528 , n274525 , n274527 );
and ( n274529 , n274528 , n240073 );
not ( n274530 , n274528 );
and ( n274531 , n274530 , n55068 );
nor ( n274532 , n274529 , n274531 );
nand ( n274533 , n274532 , n273808 );
not ( n274534 , n274533 );
not ( n274535 , n273820 );
and ( n274536 , n274534 , n274535 );
and ( n274537 , n274533 , n273820 );
nor ( n274538 , n274536 , n274537 );
or ( n274539 , n274538 , n39763 );
nand ( n274540 , n274522 , n274539 );
buf ( n274541 , n274540 );
not ( n274542 , RI19aa1618_2557);
or ( n274543 , n25328 , n274542 );
not ( n274544 , RI19a97b68_2628);
or ( n274545 , n25335 , n274544 );
nand ( n274546 , n274543 , n274545 );
buf ( n274547 , n274546 );
not ( n274548 , n266926 );
nand ( n274549 , n274548 , n257063 );
or ( n274550 , n257069 , n274549 );
not ( n274551 , n274548 );
not ( n274552 , n257037 );
or ( n274553 , n274551 , n274552 );
nor ( n274554 , n257063 , n242391 );
nand ( n274555 , n274553 , n274554 );
nand ( n274556 , n245701 , n28446 );
nand ( n274557 , n274550 , n274555 , n274556 );
buf ( n274558 , n274557 );
or ( n274559 , n25328 , n256298 );
or ( n274560 , n226822 , n266358 );
nand ( n274561 , n274559 , n274560 );
buf ( n274562 , n274561 );
not ( n274563 , n241105 );
not ( n274564 , n235580 );
or ( n274565 , n274563 , n274564 );
not ( n274566 , n241105 );
nand ( n274567 , n274566 , n235590 );
nand ( n274568 , n274565 , n274567 );
and ( n274569 , n274568 , n235720 );
not ( n274570 , n274568 );
and ( n274571 , n274570 , n243244 );
nor ( n274572 , n274569 , n274571 );
not ( n274573 , n274572 );
not ( n274574 , n252007 );
not ( n274575 , n49626 );
or ( n274576 , n274574 , n274575 );
or ( n274577 , n49626 , n252007 );
nand ( n274578 , n274576 , n274577 );
and ( n274579 , n274578 , n253265 );
not ( n274580 , n274578 );
and ( n274581 , n274580 , n253272 );
nor ( n274582 , n274579 , n274581 );
nand ( n274583 , n274573 , n274582 );
not ( n274584 , n33322 );
not ( n274585 , n233904 );
or ( n274586 , n274584 , n274585 );
or ( n274587 , n244207 , n33322 );
nand ( n274588 , n274586 , n274587 );
and ( n274589 , n274588 , n233968 );
not ( n274590 , n274588 );
and ( n274591 , n274590 , n233960 );
nor ( n274592 , n274589 , n274591 );
nand ( n274593 , n274592 , n226010 );
or ( n274594 , n274583 , n274593 );
nor ( n274595 , n274592 , n221279 );
nand ( n274596 , n274595 , n274583 );
nand ( n274597 , n245701 , n30908 );
nand ( n274598 , n274594 , n274596 , n274597 );
buf ( n274599 , n274598 );
not ( n274600 , n42791 );
not ( n274601 , n243215 );
or ( n274602 , n274600 , n274601 );
not ( n274603 , n42791 );
nand ( n274604 , n274603 , n243222 );
nand ( n274605 , n274602 , n274604 );
and ( n274606 , n274605 , n243226 );
not ( n274607 , n274605 );
and ( n274608 , n274607 , n243230 );
nor ( n274609 , n274606 , n274608 );
not ( n274610 , n274609 );
not ( n274611 , n274610 );
not ( n274612 , n274128 );
or ( n274613 , n274611 , n274612 );
nor ( n274614 , n274139 , n33254 );
nand ( n274615 , n274613 , n274614 );
nor ( n274616 , n274609 , n42443 );
nand ( n274617 , n274128 , n274616 , n274139 );
nand ( n274618 , n50615 , n34490 );
nand ( n274619 , n274615 , n274617 , n274618 );
buf ( n274620 , n274619 );
not ( n274621 , n231542 );
not ( n274622 , n238297 );
or ( n274623 , n274621 , n274622 );
or ( n274624 , n238297 , n231542 );
nand ( n274625 , n274623 , n274624 );
not ( n274626 , n274625 );
not ( n274627 , n238401 );
and ( n274628 , n274626 , n274627 );
and ( n274629 , n274625 , n238401 );
nor ( n274630 , n274628 , n274629 );
nand ( n274631 , n274630 , n237385 );
not ( n274632 , n245297 );
not ( n274633 , n254761 );
or ( n274634 , n274632 , n274633 );
or ( n274635 , n254761 , n245297 );
nand ( n274636 , n274634 , n274635 );
and ( n274637 , n274636 , n252242 );
not ( n274638 , n274636 );
and ( n274639 , n274638 , n252239 );
nor ( n274640 , n274637 , n274639 );
not ( n274641 , n274640 );
not ( n274642 , n226619 );
not ( n274643 , n274642 );
not ( n274644 , n44315 );
or ( n274645 , n274643 , n274644 );
not ( n274646 , n274642 );
nand ( n274647 , n274646 , n44324 );
nand ( n274648 , n274645 , n274647 );
and ( n274649 , n274648 , n254603 );
not ( n274650 , n274648 );
and ( n274651 , n274650 , n256460 );
nor ( n274652 , n274649 , n274651 );
nand ( n274653 , n274641 , n274652 );
or ( n274654 , n274631 , n274653 );
nor ( n274655 , n274630 , n221279 );
nand ( n274656 , n274653 , n274655 );
nand ( n274657 , n239240 , n224315 );
nand ( n274658 , n274654 , n274656 , n274657 );
buf ( n274659 , n274658 );
not ( n274660 , n233721 );
not ( n274661 , n251213 );
or ( n274662 , n274660 , n274661 );
not ( n274663 , n233721 );
nand ( n274664 , n274663 , n251217 );
nand ( n274665 , n274662 , n274664 );
and ( n274666 , n274665 , n251224 );
not ( n274667 , n274665 );
and ( n274668 , n274667 , n251220 );
nor ( n274669 , n274666 , n274668 );
not ( n274670 , n274669 );
nor ( n274671 , n274670 , n55146 );
not ( n274672 , n247457 );
not ( n274673 , n243510 );
or ( n274674 , n274672 , n274673 );
not ( n274675 , n247457 );
nand ( n274676 , n274675 , n243503 );
nand ( n274677 , n274674 , n274676 );
and ( n274678 , n274677 , n248481 );
not ( n274679 , n274677 );
and ( n274680 , n274679 , n248478 );
nor ( n274681 , n274678 , n274680 );
nand ( n274682 , n274671 , n252773 , n274681 );
nand ( n274683 , n274681 , n274669 );
nand ( n274684 , n274683 , n252774 , n241704 );
nand ( n274685 , n35431 , n206160 );
nand ( n274686 , n274682 , n274684 , n274685 );
buf ( n274687 , n274686 );
nor ( n274688 , n267165 , n43968 );
not ( n274689 , n274688 );
nand ( n274690 , n261411 , n261437 );
or ( n274691 , n274689 , n274690 );
not ( n274692 , n267166 );
not ( n274693 , n261411 );
or ( n274694 , n274692 , n274693 );
nor ( n274695 , n261437 , n234440 );
nand ( n274696 , n274694 , n274695 );
nand ( n274697 , n41945 , n205414 );
nand ( n274698 , n274691 , n274696 , n274697 );
buf ( n274699 , n274698 );
or ( n274700 , n25328 , n264639 );
or ( n274701 , n226822 , n258912 );
nand ( n274702 , n274700 , n274701 );
buf ( n274703 , n274702 );
or ( n274704 , n25328 , n264135 );
or ( n274705 , n25335 , n53009 );
nand ( n274706 , n274704 , n274705 );
buf ( n274707 , n274706 );
or ( n274708 , n25328 , n259430 );
not ( n274709 , RI19acd100_2231);
or ( n274710 , n226822 , n274709 );
nand ( n274711 , n274708 , n274710 );
buf ( n274712 , n274711 );
not ( n274713 , n249827 );
not ( n274714 , n274713 );
not ( n274715 , n272884 );
or ( n274716 , n274714 , n274715 );
or ( n274717 , n272884 , n274713 );
nand ( n274718 , n274716 , n274717 );
and ( n274719 , n274718 , n51753 );
not ( n274720 , n274718 );
and ( n274721 , n274720 , n229518 );
nor ( n274722 , n274719 , n274721 );
nand ( n274723 , n274722 , n205649 );
buf ( n274724 , n248372 );
not ( n274725 , n274724 );
not ( n274726 , n246321 );
or ( n274727 , n274725 , n274726 );
not ( n274728 , n274724 );
nand ( n274729 , n274728 , n246326 );
nand ( n274730 , n274727 , n274729 );
and ( n274731 , n274730 , n254483 );
not ( n274732 , n274730 );
and ( n274733 , n274732 , n246331 );
nor ( n274734 , n274731 , n274733 );
not ( n274735 , n274734 );
not ( n274736 , n251839 );
not ( n274737 , n258512 );
or ( n274738 , n274736 , n274737 );
not ( n274739 , n251839 );
nand ( n274740 , n274739 , n259214 );
nand ( n274741 , n274738 , n274740 );
and ( n274742 , n274741 , n260551 );
not ( n274743 , n274741 );
and ( n274744 , n274743 , n260558 );
nor ( n274745 , n274742 , n274744 );
nand ( n274746 , n274735 , n274745 );
or ( n274747 , n274723 , n274746 );
not ( n274748 , n274745 );
not ( n274749 , n274722 );
or ( n274750 , n274748 , n274749 );
nor ( n274751 , n274735 , n37725 );
nand ( n274752 , n274750 , n274751 );
nand ( n274753 , n31577 , n208196 );
nand ( n274754 , n274747 , n274752 , n274753 );
buf ( n274755 , n274754 );
not ( n274756 , n237897 );
not ( n274757 , n246759 );
or ( n274758 , n274756 , n274757 );
or ( n274759 , n246759 , n237897 );
nand ( n274760 , n274758 , n274759 );
and ( n274761 , n274760 , n254006 );
not ( n274762 , n274760 );
and ( n274763 , n274762 , n254010 );
nor ( n274764 , n274761 , n274763 );
not ( n274765 , n274764 );
nand ( n274766 , n274765 , n226010 );
not ( n274767 , n245727 );
not ( n274768 , n274767 );
not ( n274769 , n230367 );
or ( n274770 , n274768 , n274769 );
nand ( n274771 , n230374 , n245727 );
nand ( n274772 , n274770 , n274771 );
not ( n274773 , n274772 );
not ( n274774 , n52757 );
and ( n274775 , n274773 , n274774 );
and ( n274776 , n274772 , n52757 );
nor ( n274777 , n274775 , n274776 );
not ( n274778 , n274777 );
buf ( n274779 , n228439 );
not ( n274780 , n274779 );
not ( n274781 , n255503 );
or ( n274782 , n274780 , n274781 );
or ( n274783 , n255508 , n274779 );
nand ( n274784 , n274782 , n274783 );
and ( n274785 , n274784 , n265402 );
not ( n274786 , n274784 );
and ( n274787 , n274786 , n255515 );
nor ( n274788 , n274785 , n274787 );
not ( n274789 , n274788 );
nand ( n274790 , n274778 , n274789 );
or ( n274791 , n274766 , n274790 );
not ( n274792 , n274778 );
not ( n274793 , n274765 );
or ( n274794 , n274792 , n274793 );
nand ( n274795 , n274788 , n247275 );
not ( n274796 , n274795 );
nand ( n274797 , n274794 , n274796 );
nand ( n274798 , n31577 , n35990 );
nand ( n274799 , n274791 , n274797 , n274798 );
buf ( n274800 , n274799 );
not ( n274801 , n55492 );
not ( n274802 , n233967 );
or ( n274803 , n274801 , n274802 );
not ( n274804 , n55492 );
nand ( n274805 , n274804 , n233959 );
nand ( n274806 , n274803 , n274805 );
and ( n274807 , n274806 , n238621 );
not ( n274808 , n274806 );
and ( n274809 , n274808 , n238629 );
nor ( n274810 , n274807 , n274809 );
not ( n274811 , n274810 );
nor ( n274812 , n274811 , n256413 );
not ( n274813 , n225061 );
not ( n274814 , n245170 );
or ( n274815 , n274813 , n274814 );
or ( n274816 , n245170 , n225061 );
nand ( n274817 , n274815 , n274816 );
and ( n274818 , n274817 , n254080 );
not ( n274819 , n274817 );
and ( n274820 , n274819 , n254083 );
nor ( n274821 , n274818 , n274820 );
buf ( n274822 , n238926 );
not ( n274823 , n274822 );
not ( n274824 , n229763 );
or ( n274825 , n274823 , n274824 );
or ( n274826 , n229763 , n274822 );
nand ( n274827 , n274825 , n274826 );
not ( n274828 , n274827 );
not ( n274829 , n242890 );
and ( n274830 , n274828 , n274829 );
and ( n274831 , n274827 , n52223 );
nor ( n274832 , n274830 , n274831 );
not ( n274833 , n274832 );
nor ( n274834 , n274821 , n274833 );
nand ( n274835 , n274812 , n274834 );
nand ( n274836 , n274810 , n274832 );
nand ( n274837 , n274836 , n274821 , n274297 );
nand ( n274838 , n241068 , n32763 );
nand ( n274839 , n274835 , n274837 , n274838 );
buf ( n274840 , n274839 );
not ( n274841 , n242044 );
not ( n274842 , n51381 );
or ( n274843 , n274841 , n274842 );
not ( n274844 , n239841 );
not ( n274845 , n46708 );
or ( n274846 , n274844 , n274845 );
not ( n274847 , n239841 );
nand ( n274848 , n274847 , n46716 );
nand ( n274849 , n274846 , n274848 );
and ( n274850 , n274849 , n52439 );
not ( n274851 , n274849 );
and ( n274852 , n274851 , n256438 );
nor ( n274853 , n274850 , n274852 );
not ( n274854 , n236853 );
not ( n274855 , n242201 );
not ( n274856 , n274855 );
or ( n274857 , n274854 , n274856 );
not ( n274858 , n236853 );
nand ( n274859 , n274858 , n242205 );
nand ( n274860 , n274857 , n274859 );
and ( n274861 , n274860 , n255160 );
not ( n274862 , n274860 );
and ( n274863 , n274862 , n255163 );
nor ( n274864 , n274861 , n274863 );
nand ( n274865 , n274853 , n274864 );
and ( n274866 , n274865 , n274641 );
not ( n274867 , n274865 );
and ( n274868 , n274867 , n274640 );
nor ( n274869 , n274866 , n274868 );
or ( n274870 , n274869 , n258280 );
nand ( n274871 , n274843 , n274870 );
buf ( n274872 , n274871 );
not ( n274873 , n52597 );
not ( n274874 , n240053 );
or ( n274875 , n274873 , n274874 );
not ( n274876 , n52597 );
nand ( n274877 , n274876 , n240056 );
nand ( n274878 , n274875 , n274877 );
not ( n274879 , n272973 );
and ( n274880 , n274878 , n274879 );
not ( n274881 , n274878 );
and ( n274882 , n274881 , n269447 );
nor ( n274883 , n274880 , n274882 );
nand ( n274884 , n274883 , n253928 );
nand ( n274885 , n255296 , n255307 );
or ( n274886 , n274884 , n274885 );
not ( n274887 , n274883 );
not ( n274888 , n255307 );
or ( n274889 , n274887 , n274888 );
nor ( n274890 , n255296 , n55108 );
nand ( n274891 , n274889 , n274890 );
nand ( n274892 , n50615 , n38114 );
nand ( n274893 , n274886 , n274891 , n274892 );
buf ( n274894 , n274893 );
not ( n274895 , n37513 );
not ( n274896 , n258213 );
or ( n274897 , n274895 , n274896 );
not ( n274898 , n37281 );
not ( n274899 , n240799 );
or ( n274900 , n274898 , n274899 );
not ( n274901 , n37281 );
nand ( n274902 , n274901 , n240810 );
nand ( n274903 , n274900 , n274902 );
and ( n274904 , n274903 , n260011 );
not ( n274905 , n274903 );
and ( n274906 , n274905 , n252447 );
nor ( n274907 , n274904 , n274906 );
not ( n274908 , n274907 );
nand ( n274909 , n274908 , n273955 );
and ( n274910 , n274909 , n260594 );
not ( n274911 , n274909 );
and ( n274912 , n274911 , n273957 );
nor ( n274913 , n274910 , n274912 );
or ( n274914 , n274913 , n257174 );
nand ( n274915 , n274897 , n274914 );
buf ( n274916 , n274915 );
not ( n274917 , RI19a87b78_2740);
or ( n274918 , n25328 , n274917 );
or ( n274919 , n25336 , n273494 );
nand ( n274920 , n274918 , n274919 );
buf ( n274921 , n274920 );
buf ( n274922 , n26257 );
not ( n274923 , RI19acffe0_2211);
or ( n274924 , n25328 , n274923 );
or ( n274925 , n226822 , n268938 );
nand ( n274926 , n274924 , n274925 );
buf ( n274927 , n274926 );
nand ( n274928 , n262528 , n244515 );
not ( n274929 , n242577 );
nand ( n274930 , n262515 , n274929 );
or ( n274931 , n274928 , n274930 );
not ( n274932 , n262515 );
not ( n274933 , n262528 );
or ( n274934 , n274932 , n274933 );
nor ( n274935 , n274929 , n252070 );
nand ( n274936 , n274934 , n274935 );
nand ( n274937 , n234024 , n33880 );
nand ( n274938 , n274931 , n274936 , n274937 );
buf ( n274939 , n274938 );
not ( n274940 , RI19aad828_2471);
or ( n274941 , n25328 , n274940 );
not ( n274942 , RI19aa3580_2542);
or ( n274943 , n226822 , n274942 );
nand ( n274944 , n274941 , n274943 );
buf ( n274945 , n274944 );
buf ( n274946 , n37877 );
buf ( n274947 , n34162 );
not ( n274948 , n40535 );
not ( n274949 , n245702 );
or ( n274950 , n274948 , n274949 );
not ( n274951 , n237781 );
not ( n274952 , n245392 );
or ( n274953 , n274951 , n274952 );
not ( n274954 , n237781 );
nand ( n274955 , n274954 , n245402 );
nand ( n274956 , n274953 , n274955 );
and ( n274957 , n274956 , n255149 );
not ( n274958 , n274956 );
and ( n274959 , n274958 , n255146 );
nor ( n274960 , n274957 , n274959 );
nand ( n274961 , n265044 , n274960 );
and ( n274962 , n274961 , n265054 );
not ( n274963 , n274961 );
and ( n274964 , n274963 , n267004 );
nor ( n274965 , n274962 , n274964 );
or ( n274966 , n274965 , n257174 );
nand ( n274967 , n274950 , n274966 );
buf ( n274968 , n274967 );
not ( n274969 , n41710 );
not ( n274970 , n262000 );
or ( n274971 , n274969 , n274970 );
not ( n274972 , n253161 );
not ( n274973 , n223827 );
or ( n274974 , n274972 , n274973 );
not ( n274975 , n253161 );
nand ( n274976 , n274975 , n46074 );
nand ( n274977 , n274974 , n274976 );
and ( n274978 , n274977 , n244509 );
not ( n274979 , n274977 );
and ( n274980 , n274979 , n244508 );
nor ( n274981 , n274978 , n274980 );
not ( n274982 , n274981 );
not ( n274983 , n45434 );
not ( n274984 , n274983 );
not ( n274985 , n248154 );
or ( n274986 , n274984 , n274985 );
not ( n274987 , n274983 );
nand ( n274988 , n274987 , n248161 );
nand ( n274989 , n274986 , n274988 );
and ( n274990 , n274989 , n248211 );
not ( n274991 , n274989 );
and ( n274992 , n274991 , n248220 );
nor ( n274993 , n274990 , n274992 );
nand ( n274994 , n274982 , n274993 );
and ( n274995 , n274994 , n218985 );
not ( n274996 , n274994 );
and ( n274997 , n274996 , n218984 );
nor ( n274998 , n274995 , n274997 );
or ( n274999 , n274998 , n258179 );
nand ( n275000 , n274971 , n274999 );
buf ( n275001 , n275000 );
nand ( n275002 , n263572 , n266350 , n252703 );
not ( n275003 , n252678 );
not ( n275004 , n266350 );
or ( n275005 , n275003 , n275004 );
not ( n275006 , n265147 );
nand ( n275007 , n275005 , n275006 );
nand ( n275008 , n241378 , n30814 );
nand ( n275009 , n275002 , n275007 , n275008 );
buf ( n275010 , n275009 );
not ( n275011 , n274201 );
nand ( n275012 , n274441 , n252939 );
not ( n275013 , n275012 );
and ( n275014 , n275011 , n275013 );
nor ( n275015 , n256812 , n252939 );
nor ( n275016 , n275014 , n275015 );
not ( n275017 , n252874 );
nand ( n275018 , n275017 , n256810 );
nand ( n275019 , n50615 , n37186 );
nand ( n275020 , n275016 , n275018 , n275019 );
buf ( n275021 , n275020 );
not ( n275022 , n28388 );
not ( n275023 , n237361 );
or ( n275024 , n275022 , n275023 );
not ( n275025 , n254225 );
nand ( n275026 , n275025 , n260318 );
not ( n275027 , n254250 );
and ( n275028 , n275026 , n275027 );
not ( n275029 , n275026 );
and ( n275030 , n275029 , n254250 );
nor ( n275031 , n275028 , n275030 );
or ( n275032 , n275031 , n244217 );
nand ( n275033 , n275024 , n275032 );
buf ( n275034 , n275033 );
not ( n275035 , n55653 );
not ( n275036 , n251465 );
or ( n275037 , n275035 , n275036 );
not ( n275038 , n239043 );
not ( n275039 , n275038 );
not ( n275040 , n52221 );
or ( n275041 , n275039 , n275040 );
not ( n275042 , n275038 );
nand ( n275043 , n275042 , n52229 );
nand ( n275044 , n275041 , n275043 );
xor ( n275045 , n275044 , n264699 );
nand ( n275046 , n275045 , n264335 );
and ( n275047 , n265669 , n275046 );
not ( n275048 , n265669 );
not ( n275049 , n275046 );
and ( n275050 , n275048 , n275049 );
nor ( n275051 , n275047 , n275050 );
or ( n275052 , n275051 , n237358 );
nand ( n275053 , n275037 , n275052 );
buf ( n275054 , n275053 );
nor ( n275055 , n274265 , n235050 );
nand ( n275056 , n275055 , n274255 , n268416 );
not ( n275057 , n274265 );
not ( n275058 , n275057 );
not ( n275059 , n274253 );
or ( n275060 , n275058 , n275059 );
nor ( n275061 , n268416 , n250431 );
nand ( n275062 , n275060 , n275061 );
nand ( n275063 , n238638 , n29498 );
nand ( n275064 , n275056 , n275062 , n275063 );
buf ( n275065 , n275064 );
or ( n275066 , n25328 , n264141 );
or ( n275067 , n25335 , n244488 );
nand ( n275068 , n275066 , n275067 );
buf ( n275069 , n275068 );
not ( n275070 , n33988 );
not ( n275071 , n244606 );
or ( n275072 , n275070 , n275071 );
not ( n275073 , RI1754aea0_52);
or ( n275074 , n269544 , n275073 );
nand ( n275075 , n275072 , n275074 );
buf ( n275076 , n275075 );
not ( n275077 , n28307 );
not ( n275078 , n254441 );
or ( n275079 , n275077 , n275078 );
nand ( n275080 , n244534 , n244594 );
not ( n275081 , n259941 );
and ( n275082 , n275080 , n275081 );
not ( n275083 , n275080 );
and ( n275084 , n275083 , n259941 );
nor ( n275085 , n275082 , n275084 );
or ( n275086 , n275085 , n259425 );
nand ( n275087 , n275079 , n275086 );
buf ( n275088 , n275087 );
not ( n275089 , n255100 );
buf ( n275090 , n243538 );
not ( n275091 , n275090 );
and ( n275092 , n275089 , n275091 );
and ( n275093 , n258514 , n275090 );
nor ( n275094 , n275092 , n275093 );
and ( n275095 , n275094 , n259218 );
not ( n275096 , n275094 );
and ( n275097 , n275096 , n259215 );
nor ( n275098 , n275095 , n275097 );
nand ( n275099 , n275098 , n222531 );
not ( n275100 , n251207 );
nand ( n275101 , n275100 , n251226 );
or ( n275102 , n275099 , n275101 );
not ( n275103 , n275100 );
not ( n275104 , n275098 );
or ( n275105 , n275103 , n275104 );
nand ( n275106 , n275105 , n256324 );
nand ( n275107 , n236798 , n32660 );
nand ( n275108 , n275102 , n275106 , n275107 );
buf ( n275109 , n275108 );
buf ( n275110 , n205318 );
buf ( n275111 , n29558 );
nand ( n275112 , n250503 , n258206 );
buf ( n275113 , n237433 );
not ( n275114 , n275113 );
not ( n275115 , n247813 );
or ( n275116 , n275114 , n275115 );
not ( n275117 , n275113 );
nand ( n275118 , n275117 , n247822 );
nand ( n275119 , n275116 , n275118 );
and ( n275120 , n275119 , n247873 );
not ( n275121 , n275119 );
and ( n275122 , n275121 , n247872 );
nor ( n275123 , n275120 , n275122 );
not ( n275124 , n275123 );
buf ( n275125 , n245780 );
not ( n275126 , n275125 );
not ( n275127 , n245264 );
or ( n275128 , n275126 , n275127 );
or ( n275129 , n245264 , n275125 );
nand ( n275130 , n275128 , n275129 );
not ( n275131 , n275130 );
not ( n275132 , n251156 );
and ( n275133 , n275131 , n275132 );
and ( n275134 , n275130 , n251156 );
nor ( n275135 , n275133 , n275134 );
not ( n275136 , n275135 );
nand ( n275137 , n275124 , n275136 );
or ( n275138 , n275112 , n275137 );
nand ( n275139 , n250504 , n275137 );
nand ( n275140 , n251465 , n26197 );
nand ( n275141 , n275138 , n275139 , n275140 );
buf ( n275142 , n275141 );
not ( n275143 , n34284 );
not ( n275144 , n257764 );
or ( n275145 , n275143 , n275144 );
not ( n275146 , n253171 );
not ( n275147 , n223827 );
or ( n275148 , n275146 , n275147 );
not ( n275149 , n253171 );
nand ( n275150 , n275149 , n46074 );
nand ( n275151 , n275148 , n275150 );
and ( n275152 , n275151 , n244508 );
not ( n275153 , n275151 );
and ( n275154 , n275153 , n244509 );
nor ( n275155 , n275152 , n275154 );
nand ( n275156 , n275155 , n263354 );
not ( n275157 , n263365 );
and ( n275158 , n275156 , n275157 );
not ( n275159 , n275156 );
and ( n275160 , n275159 , n263365 );
nor ( n275161 , n275158 , n275160 );
or ( n275162 , n275161 , n258179 );
nand ( n275163 , n275145 , n275162 );
buf ( n275164 , n275163 );
not ( n275165 , RI19a983d8_2624);
or ( n275166 , n25328 , n275165 );
not ( n275167 , RI19a8e220_2696);
or ( n275168 , n25335 , n275167 );
nand ( n275169 , n275166 , n275168 );
buf ( n275170 , n275169 );
nand ( n275171 , n273389 , n258918 );
nor ( n275172 , n258977 , n273402 );
or ( n275173 , n275171 , n275172 );
nor ( n275174 , n273389 , n55146 );
nand ( n275175 , n275174 , n275172 );
nand ( n275176 , n254798 , n41058 );
nand ( n275177 , n275173 , n275175 , n275176 );
buf ( n275178 , n275177 );
not ( n275179 , RI1754b260_44);
or ( n275180 , n249126 , n275179 );
nand ( n275181 , n249131 , n28271 );
nand ( n275182 , n275180 , n275181 );
buf ( n275183 , n275182 );
not ( n275184 , n238638 );
not ( n275185 , n275184 );
not ( n275186 , n30089 );
and ( n275187 , n275185 , n275186 );
nor ( n275188 , n244629 , n221279 );
nor ( n275189 , n244780 , n269006 );
and ( n275190 , n275188 , n275189 );
nor ( n275191 , n275187 , n275190 );
not ( n275192 , n244630 );
nand ( n275193 , n275192 , n269006 );
nand ( n275194 , n269003 , n244780 );
nand ( n275195 , n275191 , n275193 , n275194 );
buf ( n275196 , n275195 );
or ( n275197 , n25328 , n271876 );
or ( n275198 , n25336 , n247223 );
nand ( n275199 , n275197 , n275198 );
buf ( n275200 , n275199 );
not ( n275201 , n274832 );
not ( n275202 , n274821 );
nand ( n275203 , n275201 , n275202 );
not ( n275204 , n231985 );
not ( n275205 , n275204 );
not ( n275206 , n252185 );
or ( n275207 , n275205 , n275206 );
not ( n275208 , n275204 );
nand ( n275209 , n275208 , n252192 );
nand ( n275210 , n275207 , n275209 );
and ( n275211 , n275210 , n268643 );
not ( n275212 , n275210 );
and ( n275213 , n275212 , n268640 );
nor ( n275214 , n275211 , n275213 );
nor ( n275215 , n275214 , n235732 );
not ( n275216 , n275215 );
or ( n275217 , n275203 , n275216 );
not ( n275218 , n275214 );
nor ( n275219 , n275218 , n235050 );
nand ( n275220 , n275203 , n275219 );
nand ( n275221 , n250916 , n35771 );
nand ( n275222 , n275217 , n275220 , n275221 );
buf ( n275223 , n275222 );
not ( n275224 , n224724 );
not ( n275225 , n262000 );
or ( n275226 , n275224 , n275225 );
nand ( n275227 , n266671 , n272341 );
not ( n275228 , n261507 );
and ( n275229 , n275227 , n275228 );
not ( n275230 , n275227 );
and ( n275231 , n275230 , n261507 );
nor ( n275232 , n275229 , n275231 );
or ( n275233 , n275232 , n49959 );
nand ( n275234 , n275226 , n275233 );
buf ( n275235 , n275234 );
or ( n275236 , n25328 , n273096 );
or ( n275237 , n25336 , n254428 );
nand ( n275238 , n275236 , n275237 );
buf ( n275239 , n275238 );
buf ( n275240 , n30491 );
buf ( n275241 , n30598 );
and ( n275242 , n27883 , n204520 );
buf ( n275243 , n275242 );
not ( n275244 , n272167 );
not ( n275245 , n253181 );
not ( n275246 , n223827 );
or ( n275247 , n275245 , n275246 );
not ( n275248 , n253181 );
nand ( n275249 , n275248 , n46074 );
nand ( n275250 , n275247 , n275249 );
and ( n275251 , n275250 , n244509 );
not ( n275252 , n275250 );
and ( n275253 , n275252 , n244508 );
nor ( n275254 , n275251 , n275253 );
not ( n275255 , n235869 );
not ( n275256 , n245793 );
or ( n275257 , n275255 , n275256 );
not ( n275258 , n235869 );
nand ( n275259 , n275258 , n245797 );
nand ( n275260 , n275257 , n275259 );
and ( n275261 , n275260 , n250808 );
not ( n275262 , n275260 );
and ( n275263 , n275262 , n250813 );
nor ( n275264 , n275261 , n275263 );
nand ( n275265 , n275254 , n275264 );
or ( n275266 , n275244 , n275265 );
not ( n275267 , n275264 );
not ( n275268 , n272163 );
or ( n275269 , n275267 , n275268 );
nor ( n275270 , n275254 , n52445 );
nand ( n275271 , n275269 , n275270 );
nand ( n275272 , n241976 , n31054 );
nand ( n275273 , n275266 , n275271 , n275272 );
buf ( n275274 , n275273 );
or ( n275275 , n226819 , n256421 );
or ( n275276 , n25335 , n271874 );
nand ( n275277 , n275275 , n275276 );
buf ( n275278 , n275277 );
buf ( n275279 , n217113 );
buf ( n275280 , n28539 );
nand ( n275281 , n266730 , n43969 );
nor ( n275282 , n253681 , n266733 );
or ( n275283 , n275281 , n275282 );
nor ( n275284 , n266730 , n40465 );
nand ( n275285 , n275284 , n275282 );
nand ( n275286 , n234453 , n26469 );
nand ( n275287 , n275283 , n275285 , n275286 );
buf ( n275288 , n275287 );
not ( n275289 , n29078 );
not ( n275290 , n51381 );
or ( n275291 , n275289 , n275290 );
not ( n275292 , n264275 );
not ( n275293 , n236220 );
not ( n275294 , n241256 );
or ( n275295 , n275293 , n275294 );
not ( n275296 , n236220 );
nand ( n275297 , n275296 , n241255 );
nand ( n275298 , n275295 , n275297 );
and ( n275299 , n275298 , n241370 );
not ( n275300 , n275298 );
and ( n275301 , n275300 , n241361 );
nor ( n275302 , n275299 , n275301 );
nand ( n275303 , n275292 , n275302 );
and ( n275304 , n275303 , n260972 );
not ( n275305 , n275303 );
and ( n275306 , n275305 , n260971 );
nor ( n275307 , n275304 , n275306 );
or ( n275308 , n275307 , n49959 );
nand ( n275309 , n275291 , n275308 );
buf ( n275310 , n275309 );
not ( n275311 , RI19a88be0_2733);
or ( n275312 , n25328 , n275311 );
or ( n275313 , n226822 , n262545 );
nand ( n275314 , n275312 , n275313 );
buf ( n275315 , n275314 );
buf ( n275316 , n38114 );
buf ( n275317 , n35057 );
not ( n275318 , n245526 );
not ( n275319 , n267895 );
not ( n275320 , n275319 );
or ( n275321 , n275318 , n275320 );
nor ( n275322 , n245683 , n46425 );
nand ( n275323 , n275321 , n275322 );
nand ( n275324 , n267897 , n275319 , n245683 );
nand ( n275325 , n234024 , n43257 );
nand ( n275326 , n275323 , n275324 , n275325 );
buf ( n275327 , n275326 );
not ( n275328 , n272839 );
nand ( n275329 , n275328 , n264905 );
not ( n275330 , n275329 );
nor ( n275331 , n272851 , n252358 );
not ( n275332 , n275331 );
or ( n275333 , n275330 , n275332 );
nor ( n275334 , n272839 , n252070 );
and ( n275335 , n275334 , n272851 , n264905 );
not ( n275336 , n35851 );
nor ( n275337 , n275336 , n263991 );
nor ( n275338 , n275335 , n275337 );
nand ( n275339 , n275333 , n275338 );
buf ( n275340 , n275339 );
not ( n275341 , RI19a88028_2738);
or ( n275342 , n25328 , n275341 );
not ( n275343 , RI19acc3e0_2237);
or ( n275344 , n25336 , n275343 );
nand ( n275345 , n275342 , n275344 );
buf ( n275346 , n275345 );
not ( n275347 , n254841 );
not ( n275348 , n55345 );
or ( n275349 , n275347 , n275348 );
not ( n275350 , n254841 );
nand ( n275351 , n275350 , n33708 );
nand ( n275352 , n275349 , n275351 );
and ( n275353 , n275352 , n233265 );
not ( n275354 , n275352 );
and ( n275355 , n275354 , n55511 );
nor ( n275356 , n275353 , n275355 );
not ( n275357 , n275356 );
nand ( n275358 , n275357 , n241459 );
not ( n275359 , n244740 );
not ( n275360 , n241877 );
or ( n275361 , n275359 , n275360 );
not ( n275362 , n244740 );
nand ( n275363 , n275362 , n241884 );
nand ( n275364 , n275361 , n275363 );
and ( n275365 , n275364 , n254238 );
not ( n275366 , n275364 );
and ( n275367 , n275366 , n254235 );
nor ( n275368 , n275365 , n275367 );
not ( n275369 , n275368 );
nand ( n275370 , n259557 , n275369 );
or ( n275371 , n275358 , n275370 );
not ( n275372 , n259557 );
not ( n275373 , n275357 );
or ( n275374 , n275372 , n275373 );
nor ( n275375 , n275369 , n40465 );
nand ( n275376 , n275374 , n275375 );
nand ( n275377 , n252711 , n33633 );
nand ( n275378 , n275371 , n275376 , n275377 );
buf ( n275379 , n275378 );
or ( n275380 , n226819 , n274193 );
or ( n275381 , n25336 , n262581 );
nand ( n275382 , n275380 , n275381 );
buf ( n275383 , n275382 );
nand ( n275384 , n265575 , n50945 );
not ( n275385 , n262746 );
nand ( n275386 , n262735 , n275385 );
or ( n275387 , n275384 , n275386 );
not ( n275388 , n275385 );
not ( n275389 , n265575 );
or ( n275390 , n275388 , n275389 );
nor ( n275391 , n262735 , n55152 );
nand ( n275392 , n275390 , n275391 );
nand ( n275393 , n37728 , n29969 );
nand ( n275394 , n275387 , n275392 , n275393 );
buf ( n275395 , n275394 );
or ( n275396 , n25328 , n274709 );
not ( n275397 , RI19ac4460_2297);
or ( n275398 , n25335 , n275397 );
nand ( n275399 , n275396 , n275398 );
buf ( n275400 , n275399 );
not ( n275401 , n29935 );
not ( n275402 , n234453 );
or ( n275403 , n275401 , n275402 );
nand ( n275404 , n266904 , n242082 );
and ( n275405 , n275404 , n48809 );
not ( n275406 , n275404 );
and ( n275407 , n275406 , n226569 );
nor ( n275408 , n275405 , n275407 );
or ( n275409 , n275408 , n52445 );
nand ( n275410 , n275403 , n275409 );
buf ( n275411 , n275410 );
not ( n275412 , RI19a88460_2736);
or ( n275413 , n226819 , n275412 );
not ( n275414 , RI19acc818_2235);
or ( n275415 , n226822 , n275414 );
nand ( n275416 , n275413 , n275415 );
buf ( n275417 , n275416 );
not ( n275418 , RI19aca298_2254);
or ( n275419 , n25328 , n275418 );
not ( n275420 , RI19ac0f68_2323);
or ( n275421 , n25336 , n275420 );
nand ( n275422 , n275419 , n275421 );
buf ( n275423 , n275422 );
nand ( n275424 , n273291 , n40466 );
not ( n275425 , n247138 );
not ( n275426 , n253474 );
or ( n275427 , n275425 , n275426 );
not ( n275428 , n247138 );
nand ( n275429 , n275428 , n248276 );
nand ( n275430 , n275427 , n275429 );
and ( n275431 , n275430 , n248281 );
not ( n275432 , n275430 );
and ( n275433 , n275432 , n248284 );
nor ( n275434 , n275431 , n275433 );
not ( n275435 , n275434 );
nand ( n275436 , n275435 , n273316 );
or ( n275437 , n275424 , n275436 );
not ( n275438 , n273316 );
not ( n275439 , n273291 );
or ( n275440 , n275438 , n275439 );
nor ( n275441 , n275435 , n47173 );
nand ( n275442 , n275440 , n275441 );
nand ( n275443 , n234453 , n35551 );
nand ( n275444 , n275437 , n275442 , n275443 );
buf ( n275445 , n275444 );
not ( n275446 , n37314 );
not ( n275447 , n51381 );
or ( n275448 , n275446 , n275447 );
nand ( n275449 , n258722 , n258733 );
not ( n275450 , n272234 );
and ( n275451 , n275449 , n275450 );
not ( n275452 , n275449 );
and ( n275453 , n275452 , n272234 );
nor ( n275454 , n275451 , n275453 );
or ( n275455 , n275454 , n251498 );
nand ( n275456 , n275448 , n275455 );
buf ( n275457 , n275456 );
buf ( n275458 , n34174 );
nand ( n275459 , n245405 , n234111 );
nand ( n275460 , n263996 , n263884 );
or ( n275461 , n275459 , n275460 );
not ( n275462 , n263996 );
not ( n275463 , n245405 );
or ( n275464 , n275462 , n275463 );
not ( n275465 , n205649 );
nor ( n275466 , n275465 , n263884 );
nand ( n275467 , n275464 , n275466 );
nand ( n275468 , n49054 , n37985 );
nand ( n275469 , n275461 , n275467 , n275468 );
buf ( n275470 , n275469 );
buf ( n275471 , n32591 );
buf ( n275472 , n34251 );
not ( n275473 , n242410 );
nor ( n275474 , n275473 , n242577 );
nand ( n275475 , n262535 , n275474 );
not ( n275476 , n274929 );
not ( n275477 , n262515 );
not ( n275478 , n275477 );
or ( n275479 , n275476 , n275478 );
nor ( n275480 , n242410 , n46425 );
nand ( n275481 , n275479 , n275480 );
nand ( n275482 , n31577 , n205210 );
nand ( n275483 , n275475 , n275481 , n275482 );
buf ( n275484 , n275483 );
nor ( n275485 , n274722 , n252872 );
not ( n275486 , n275485 );
not ( n275487 , n32464 );
not ( n275488 , n51269 );
not ( n275489 , n275488 );
or ( n275490 , n275487 , n275489 );
not ( n275491 , n32464 );
nand ( n275492 , n275491 , n51269 );
nand ( n275493 , n275490 , n275492 );
and ( n275494 , n275493 , n250746 );
not ( n275495 , n275493 );
and ( n275496 , n275495 , n269613 );
nor ( n275497 , n275494 , n275496 );
nor ( n275498 , n275497 , n274745 );
or ( n275499 , n275486 , n275498 );
not ( n275500 , n274722 );
nor ( n275501 , n275500 , n238900 );
nand ( n275502 , n275501 , n275498 );
nand ( n275503 , n41945 , n204289 );
nand ( n275504 , n275499 , n275502 , n275503 );
buf ( n275505 , n275504 );
not ( n275506 , n238316 );
not ( n275507 , n254337 );
or ( n275508 , n275506 , n275507 );
not ( n275509 , n238316 );
nand ( n275510 , n275509 , n254344 );
nand ( n275511 , n275508 , n275510 );
and ( n275512 , n275511 , n256646 );
not ( n275513 , n275511 );
and ( n275514 , n275513 , n256649 );
nor ( n275515 , n275512 , n275514 );
nor ( n275516 , n275515 , n248810 );
nand ( n275517 , n254736 , n275516 );
not ( n275518 , n248811 );
not ( n275519 , n254739 );
or ( n275520 , n275518 , n275519 );
not ( n275521 , n275515 );
nor ( n275522 , n275521 , n37725 );
nand ( n275523 , n275520 , n275522 );
nand ( n275524 , n39767 , n204277 );
nand ( n275525 , n275517 , n275523 , n275524 );
buf ( n275526 , n275525 );
buf ( n275527 , n234227 );
not ( n275528 , n275527 );
not ( n275529 , n41933 );
or ( n275530 , n275528 , n275529 );
or ( n275531 , n41933 , n275527 );
nand ( n275532 , n275530 , n275531 );
not ( n275533 , n275532 );
not ( n275534 , n262783 );
and ( n275535 , n275533 , n275534 );
and ( n275536 , n275532 , n261058 );
nor ( n275537 , n275535 , n275536 );
not ( n275538 , n250220 );
not ( n275539 , n249381 );
or ( n275540 , n275538 , n275539 );
not ( n275541 , n250220 );
nand ( n275542 , n275541 , n243197 );
nand ( n275543 , n275540 , n275542 );
and ( n275544 , n275543 , n249395 );
not ( n275545 , n275543 );
and ( n275546 , n275545 , n249398 );
nor ( n275547 , n275544 , n275546 );
not ( n275548 , n275547 );
nand ( n275549 , n275537 , n275548 );
or ( n275550 , n275549 , n263696 );
nand ( n275551 , n275549 , n263702 );
nand ( n275552 , n35431 , n29144 );
nand ( n275553 , n275550 , n275551 , n275552 );
buf ( n275554 , n275553 );
not ( n275555 , n33993 );
not ( n275556 , n234453 );
or ( n275557 , n275555 , n275556 );
not ( n275558 , n246313 );
not ( n275559 , n260985 );
or ( n275560 , n275558 , n275559 );
not ( n275561 , n246313 );
nand ( n275562 , n275561 , n244116 );
nand ( n275563 , n275560 , n275562 );
and ( n275564 , n275563 , n239654 );
not ( n275565 , n275563 );
and ( n275566 , n275565 , n244127 );
nor ( n275567 , n275564 , n275566 );
nand ( n275568 , n275567 , n271818 );
and ( n275569 , n275568 , n273217 );
not ( n275570 , n275568 );
and ( n275571 , n275570 , n273216 );
nor ( n275572 , n275569 , n275571 );
or ( n275573 , n275572 , n52445 );
nand ( n275574 , n275557 , n275573 );
buf ( n275575 , n275574 );
not ( n275576 , n30613 );
not ( n275577 , n234453 );
or ( n275578 , n275576 , n275577 );
nand ( n275579 , n273633 , n273647 );
not ( n275580 , n250093 );
not ( n275581 , n275580 );
not ( n275582 , n236063 );
not ( n275583 , n275582 );
or ( n275584 , n275581 , n275583 );
nand ( n275585 , n236063 , n250093 );
nand ( n275586 , n275584 , n275585 );
and ( n275587 , n275586 , n236167 );
not ( n275588 , n275586 );
and ( n275589 , n275588 , n236171 );
nor ( n275590 , n275587 , n275589 );
not ( n275591 , n275590 );
and ( n275592 , n275579 , n275591 );
not ( n275593 , n275579 );
and ( n275594 , n275593 , n275590 );
nor ( n275595 , n275592 , n275594 );
or ( n275596 , n275595 , n253544 );
nand ( n275597 , n275578 , n275596 );
buf ( n275598 , n275597 );
not ( n275599 , RI19acef78_2218);
or ( n275600 , n233507 , n275599 );
or ( n275601 , n25336 , n251565 );
nand ( n275602 , n275600 , n275601 );
buf ( n275603 , n275602 );
or ( n275604 , n25328 , n275420 );
not ( n275605 , RI19ab82c8_2394);
or ( n275606 , n25336 , n275605 );
nand ( n275607 , n275604 , n275606 );
buf ( n275608 , n275607 );
not ( n275609 , n261389 );
nand ( n275610 , n275609 , n270222 );
not ( n275611 , n261377 );
or ( n275612 , n275610 , n275611 );
nand ( n275613 , n275610 , n256030 );
nand ( n275614 , n50615 , n33869 );
nand ( n275615 , n275612 , n275613 , n275614 );
buf ( n275616 , n275615 );
buf ( n275617 , n36055 );
buf ( n275618 , n38995 );
not ( n275619 , RI19aa5740_2526);
or ( n275620 , n25328 , n275619 );
not ( n275621 , RI19a9c1b8_2597);
or ( n275622 , n25335 , n275621 );
nand ( n275623 , n275620 , n275622 );
buf ( n275624 , n275623 );
buf ( n275625 , n32985 );
buf ( n275626 , n35350 );
not ( n275627 , n259891 );
nand ( n275628 , n275627 , n259917 );
or ( n275629 , n263716 , n275628 );
nor ( n275630 , n263715 , n50944 );
nand ( n275631 , n275630 , n275628 );
nand ( n275632 , n246460 , n30920 );
nand ( n275633 , n275629 , n275631 , n275632 );
buf ( n275634 , n275633 );
not ( n275635 , n37080 );
not ( n275636 , n234453 );
or ( n275637 , n275635 , n275636 );
nand ( n275638 , n262788 , n262799 );
not ( n275639 , n268151 );
and ( n275640 , n275638 , n275639 );
not ( n275641 , n275638 );
and ( n275642 , n275641 , n268151 );
nor ( n275643 , n275640 , n275642 );
or ( n275644 , n275643 , n235052 );
nand ( n275645 , n275637 , n275644 );
buf ( n275646 , n275645 );
nand ( n275647 , n270496 , n270663 , n263441 );
nand ( n275648 , n270494 , n263441 );
nand ( n275649 , n275648 , n270664 , n254528 );
nand ( n275650 , n254798 , n226680 );
nand ( n275651 , n275647 , n275649 , n275650 );
buf ( n275652 , n275651 );
not ( n275653 , n34029 );
not ( n275654 , n51381 );
or ( n275655 , n275653 , n275654 );
not ( n275656 , n55467 );
not ( n275657 , n233967 );
or ( n275658 , n275656 , n275657 );
not ( n275659 , n55467 );
nand ( n275660 , n275659 , n233959 );
nand ( n275661 , n275658 , n275660 );
and ( n275662 , n275661 , n238621 );
not ( n275663 , n275661 );
and ( n275664 , n275663 , n238629 );
nor ( n275665 , n275662 , n275664 );
not ( n275666 , n252115 );
not ( n275667 , n47310 );
or ( n275668 , n275666 , n275667 );
not ( n275669 , n252115 );
nand ( n275670 , n275669 , n47319 );
nand ( n275671 , n275668 , n275670 );
and ( n275672 , n275671 , n225083 );
not ( n275673 , n275671 );
and ( n275674 , n275673 , n225086 );
nor ( n275675 , n275672 , n275674 );
nand ( n275676 , n275665 , n275675 );
not ( n275677 , n46499 );
not ( n275678 , n51606 );
or ( n275679 , n275677 , n275678 );
not ( n275680 , n46499 );
nand ( n275681 , n275680 , n51597 );
nand ( n275682 , n275679 , n275681 );
and ( n275683 , n275682 , n253197 );
not ( n275684 , n275682 );
and ( n275685 , n275684 , n253189 );
nor ( n275686 , n275683 , n275685 );
not ( n275687 , n275686 );
and ( n275688 , n275676 , n275687 );
not ( n275689 , n275676 );
and ( n275690 , n275689 , n275686 );
nor ( n275691 , n275688 , n275690 );
or ( n275692 , n275691 , n258280 );
nand ( n275693 , n275655 , n275692 );
buf ( n275694 , n275693 );
not ( n275695 , n247297 );
nand ( n275696 , n275695 , n241459 );
not ( n275697 , n235991 );
not ( n275698 , n260550 );
or ( n275699 , n275697 , n275698 );
not ( n275700 , n235991 );
nand ( n275701 , n275700 , n260557 );
nand ( n275702 , n275699 , n275701 );
and ( n275703 , n275702 , n262915 );
not ( n275704 , n275702 );
and ( n275705 , n275704 , n262914 );
nor ( n275706 , n275703 , n275705 );
nand ( n275707 , n247406 , n275706 );
or ( n275708 , n275696 , n275707 );
not ( n275709 , n247406 );
not ( n275710 , n275695 );
or ( n275711 , n275709 , n275710 );
nor ( n275712 , n275706 , n37724 );
nand ( n275713 , n275711 , n275712 );
nand ( n275714 , n244484 , n41716 );
nand ( n275715 , n275708 , n275713 , n275714 );
buf ( n275716 , n275715 );
nand ( n275717 , n267178 , n261423 );
not ( n275718 , n267167 );
or ( n275719 , n275717 , n275718 );
nand ( n275720 , n274688 , n275717 );
nand ( n275721 , n41944 , n30343 );
nand ( n275722 , n275719 , n275720 , n275721 );
buf ( n275723 , n275722 );
nor ( n275724 , n264937 , n264925 );
nand ( n275725 , n273040 , n275724 );
not ( n275726 , n264937 );
not ( n275727 , n275726 );
not ( n275728 , n273038 );
or ( n275729 , n275727 , n275728 );
nor ( n275730 , n264926 , n238635 );
nand ( n275731 , n275729 , n275730 );
nand ( n275732 , n261585 , n31337 );
nand ( n275733 , n275725 , n275731 , n275732 );
buf ( n275734 , n275733 );
not ( n275735 , n31646 );
not ( n275736 , n55760 );
or ( n275737 , n275735 , n275736 );
nand ( n275738 , n252244 , n256397 );
and ( n275739 , n275738 , n271923 );
not ( n275740 , n275738 );
and ( n275741 , n275740 , n271922 );
nor ( n275742 , n275739 , n275741 );
or ( n275743 , n275742 , n226003 );
nand ( n275744 , n275737 , n275743 );
buf ( n275745 , n275744 );
not ( n275746 , n32820 );
not ( n275747 , n234453 );
or ( n275748 , n275746 , n275747 );
nand ( n275749 , n266548 , n273936 );
and ( n275750 , n275749 , n272102 );
not ( n275751 , n275749 );
and ( n275752 , n275751 , n266560 );
nor ( n275753 , n275750 , n275752 );
or ( n275754 , n275753 , n244837 );
nand ( n275755 , n275748 , n275754 );
buf ( n275756 , n275755 );
not ( n275757 , n41887 );
not ( n275758 , n233090 );
or ( n275759 , n275757 , n275758 );
not ( n275760 , n41887 );
nand ( n275761 , n275760 , n55322 );
nand ( n275762 , n275759 , n275761 );
and ( n275763 , n275762 , n272687 );
not ( n275764 , n275762 );
and ( n275765 , n275764 , n242272 );
nor ( n275766 , n275763 , n275765 );
not ( n275767 , n275766 );
nand ( n275768 , n275687 , n275767 );
not ( n275769 , n275768 );
buf ( n275770 , n44446 );
not ( n275771 , n275770 );
not ( n275772 , n241360 );
or ( n275773 , n275771 , n275772 );
not ( n275774 , n275770 );
nand ( n275775 , n275774 , n241369 );
nand ( n275776 , n275773 , n275775 );
not ( n275777 , n275776 );
not ( n275778 , n258972 );
and ( n275779 , n275777 , n275778 );
and ( n275780 , n275776 , n258972 );
nor ( n275781 , n275779 , n275780 );
nor ( n275782 , n275781 , n255014 );
not ( n275783 , n275782 );
or ( n275784 , n275769 , n275783 );
nor ( n275785 , n275766 , n31572 );
and ( n275786 , n275785 , n275781 , n275687 );
not ( n275787 , n29699 );
not ( n275788 , n41944 );
nor ( n275789 , n275787 , n275788 );
nor ( n275790 , n275786 , n275789 );
nand ( n275791 , n275784 , n275790 );
buf ( n275792 , n275791 );
or ( n275793 , n25328 , n263814 );
or ( n275794 , n25335 , n262137 );
nand ( n275795 , n275793 , n275794 );
buf ( n275796 , n275795 );
not ( n275797 , n41772 );
not ( n275798 , n275797 );
not ( n275799 , n233090 );
or ( n275800 , n275798 , n275799 );
not ( n275801 , n275797 );
nand ( n275802 , n275801 , n55322 );
nand ( n275803 , n275800 , n275802 );
and ( n275804 , n275803 , n242272 );
not ( n275805 , n275803 );
and ( n275806 , n275805 , n272687 );
nor ( n275807 , n275804 , n275806 );
not ( n275808 , n275807 );
not ( n275809 , n239335 );
not ( n275810 , n252917 );
or ( n275811 , n275809 , n275810 );
not ( n275812 , n239335 );
nand ( n275813 , n275812 , n258055 );
nand ( n275814 , n275811 , n275813 );
and ( n275815 , n275814 , n258058 );
not ( n275816 , n275814 );
and ( n275817 , n275816 , n258061 );
nor ( n275818 , n275815 , n275817 );
not ( n275819 , n275818 );
not ( n275820 , n275819 );
or ( n275821 , n275808 , n275820 );
nand ( n275822 , n275821 , n263107 );
not ( n275823 , n275807 );
nor ( n275824 , n275823 , n31572 );
nand ( n275825 , n275824 , n263106 , n275819 );
nand ( n275826 , n244987 , n34804 );
nand ( n275827 , n275822 , n275825 , n275826 );
buf ( n275828 , n275827 );
nand ( n275829 , n272795 , n235051 );
not ( n275830 , n260532 );
not ( n275831 , n275830 );
not ( n275832 , n50274 );
or ( n275833 , n275831 , n275832 );
not ( n275834 , n275830 );
nand ( n275835 , n275834 , n228042 );
nand ( n275836 , n275833 , n275835 );
and ( n275837 , n275836 , n50483 );
not ( n275838 , n275836 );
and ( n275839 , n275838 , n50475 );
nor ( n275840 , n275837 , n275839 );
not ( n275841 , n275840 );
not ( n275842 , n253287 );
not ( n275843 , n243043 );
not ( n275844 , n273449 );
or ( n275845 , n275843 , n275844 );
nand ( n275846 , n248677 , n243042 );
nand ( n275847 , n275845 , n275846 );
not ( n275848 , n275847 );
or ( n275849 , n275842 , n275848 );
or ( n275850 , n253287 , n275847 );
nand ( n275851 , n275849 , n275850 );
not ( n275852 , n275851 );
nand ( n275853 , n275841 , n275852 );
or ( n275854 , n275829 , n275853 );
not ( n275855 , n275852 );
not ( n275856 , n272795 );
or ( n275857 , n275855 , n275856 );
nor ( n275858 , n275841 , n52445 );
nand ( n275859 , n275857 , n275858 );
nand ( n275860 , n31577 , n30193 );
nand ( n275861 , n275854 , n275859 , n275860 );
buf ( n275862 , n275861 );
not ( n275863 , n259324 );
not ( n275864 , n265952 );
or ( n275865 , n275863 , n275864 );
not ( n275866 , n55147 );
nor ( n275867 , n275866 , n268510 );
nand ( n275868 , n275865 , n275867 );
nor ( n275869 , n259310 , n265349 );
nand ( n275870 , n259321 , n275869 );
nand ( n275871 , n39767 , n36006 );
nand ( n275872 , n275868 , n275870 , n275871 );
buf ( n275873 , n275872 );
not ( n275874 , n274735 );
not ( n275875 , n275500 );
or ( n275876 , n275874 , n275875 );
not ( n275877 , n247374 );
not ( n275878 , n240504 );
or ( n275879 , n275877 , n275878 );
or ( n275880 , n240508 , n247374 );
nand ( n275881 , n275879 , n275880 );
not ( n275882 , n275881 );
not ( n275883 , n246173 );
and ( n275884 , n275882 , n275883 );
and ( n275885 , n275881 , n246173 );
nor ( n275886 , n275884 , n275885 );
nor ( n275887 , n275886 , n236795 );
nand ( n275888 , n275876 , n275887 );
not ( n275889 , n275886 );
nor ( n275890 , n275889 , n274734 );
nand ( n275891 , n275485 , n275890 );
nand ( n275892 , n31576 , n206723 );
nand ( n275893 , n275888 , n275891 , n275892 );
buf ( n275894 , n275893 );
not ( n275895 , n31170 );
not ( n275896 , n234823 );
or ( n275897 , n275895 , n275896 );
not ( n275898 , n247528 );
not ( n275899 , n243801 );
or ( n275900 , n275898 , n275899 );
not ( n275901 , n247528 );
nand ( n275902 , n275901 , n243810 );
nand ( n275903 , n275900 , n275902 );
and ( n275904 , n275903 , n243960 );
not ( n275905 , n275903 );
and ( n275906 , n275905 , n243954 );
nor ( n275907 , n275904 , n275906 );
not ( n275908 , n46121 );
not ( n275909 , n54195 );
or ( n275910 , n275908 , n275909 );
not ( n275911 , n46121 );
nand ( n275912 , n275911 , n231952 );
nand ( n275913 , n275910 , n275912 );
and ( n275914 , n275913 , n264882 );
not ( n275915 , n275913 );
and ( n275916 , n275915 , n264879 );
nor ( n275917 , n275914 , n275916 );
nand ( n275918 , n275907 , n275917 );
not ( n275919 , n49936 );
not ( n275920 , n275919 );
not ( n275921 , n245862 );
or ( n275922 , n275920 , n275921 );
not ( n275923 , n275919 );
nand ( n275924 , n275923 , n245872 );
nand ( n275925 , n275922 , n275924 );
and ( n275926 , n275925 , n245930 );
not ( n275927 , n275925 );
and ( n275928 , n275927 , n245920 );
nor ( n275929 , n275926 , n275928 );
and ( n275930 , n275918 , n275929 );
not ( n275931 , n275918 );
not ( n275932 , n275929 );
and ( n275933 , n275931 , n275932 );
nor ( n275934 , n275930 , n275933 );
or ( n275935 , n275934 , n251498 );
nand ( n275936 , n275897 , n275935 );
buf ( n275937 , n275936 );
buf ( n275938 , n251272 );
not ( n275939 , n275938 );
not ( n275940 , n249939 );
or ( n275941 , n275939 , n275940 );
or ( n275942 , n249006 , n275938 );
nand ( n275943 , n275941 , n275942 );
and ( n275944 , n275943 , n249929 );
not ( n275945 , n275943 );
and ( n275946 , n275945 , n267247 );
nor ( n275947 , n275944 , n275946 );
nor ( n275948 , n275947 , n35816 );
nand ( n275949 , n275948 , n271223 , n259958 );
not ( n275950 , n275947 );
not ( n275951 , n275950 );
not ( n275952 , n271223 );
or ( n275953 , n275951 , n275952 );
nand ( n275954 , n275953 , n259959 );
nand ( n275955 , n31577 , n31192 );
nand ( n275956 , n275949 , n275954 , n275955 );
buf ( n275957 , n275956 );
not ( n275958 , n252148 );
not ( n275959 , n220460 );
or ( n275960 , n275958 , n275959 );
not ( n275961 , n252148 );
nand ( n275962 , n275961 , n220467 );
nand ( n275963 , n275960 , n275962 );
and ( n275964 , n275963 , n43011 );
not ( n275965 , n275963 );
and ( n275966 , n275965 , n43006 );
nor ( n275967 , n275964 , n275966 );
and ( n275968 , n275967 , n254660 );
nor ( n275969 , n275968 , n43968 );
and ( n275970 , n275969 , n262955 );
not ( n275971 , n35431 );
nor ( n275972 , n275971 , n30868 );
nor ( n275973 , n275970 , n275972 );
not ( n275974 , n275967 );
nor ( n275975 , n275974 , n219702 );
not ( n275976 , n262955 );
nand ( n275977 , n275975 , n275976 , n254660 );
nand ( n275978 , n275973 , n275977 );
buf ( n275979 , n275978 );
not ( n275980 , n250771 );
not ( n275981 , n275980 );
not ( n275982 , n251154 );
or ( n275983 , n275981 , n275982 );
not ( n275984 , n275980 );
nand ( n275985 , n275984 , n251253 );
nand ( n275986 , n275983 , n275985 );
and ( n275987 , n275986 , n251314 );
not ( n275988 , n275986 );
and ( n275989 , n275988 , n251299 );
nor ( n275990 , n275987 , n275989 );
not ( n275991 , n275990 );
nand ( n275992 , n266858 , n275991 );
or ( n275993 , n265212 , n275992 );
not ( n275994 , n275991 );
not ( n275995 , n265211 );
or ( n275996 , n275994 , n275995 );
nor ( n275997 , n266858 , n55108 );
nand ( n275998 , n275996 , n275997 );
nand ( n275999 , n234448 , n29265 );
nand ( n276000 , n275993 , n275998 , n275999 );
buf ( n276001 , n276000 );
or ( n276002 , n25328 , n238229 );
or ( n276003 , n25336 , n272217 );
nand ( n276004 , n276002 , n276003 );
buf ( n276005 , n276004 );
buf ( n276006 , RI19ad0bb0_2206);
and ( n276007 , n25326 , n276006 );
buf ( n276008 , n276007 );
not ( n276009 , n250914 );
nand ( n276010 , n263158 , n270306 );
or ( n276011 , n276009 , n276010 );
not ( n276012 , n263158 );
not ( n276013 , n250908 );
or ( n276014 , n276012 , n276013 );
nor ( n276015 , n270306 , n52445 );
nand ( n276016 , n276014 , n276015 );
nand ( n276017 , n245414 , n28951 );
nand ( n276018 , n276011 , n276016 , n276017 );
buf ( n276019 , n276018 );
nand ( n276020 , n269088 , n257190 );
nand ( n276021 , n257201 , n50945 );
or ( n276022 , n276020 , n276021 );
nor ( n276023 , n257201 , n238635 );
nand ( n276024 , n276020 , n276023 );
nand ( n276025 , n39767 , n25355 );
nand ( n276026 , n276022 , n276024 , n276025 );
buf ( n276027 , n276026 );
not ( n276028 , n40854 );
not ( n276029 , n244789 );
or ( n276030 , n276028 , n276029 );
not ( n276031 , n245620 );
nand ( n276032 , n276031 , n267884 );
and ( n276033 , n276032 , n275319 );
not ( n276034 , n276032 );
and ( n276035 , n276034 , n267895 );
nor ( n276036 , n276033 , n276035 );
or ( n276037 , n276036 , n260861 );
nand ( n276038 , n276030 , n276037 );
buf ( n276039 , n276038 );
nor ( n276040 , n264776 , n254100 );
nand ( n276041 , n262866 , n276040 );
not ( n276042 , n262863 );
not ( n276043 , n276042 );
not ( n276044 , n264776 );
not ( n276045 , n276044 );
or ( n276046 , n276043 , n276045 );
nand ( n276047 , n276046 , n254066 );
nand ( n276048 , n246217 , n28522 );
nand ( n276049 , n276041 , n276047 , n276048 );
buf ( n276050 , n276049 );
not ( n276051 , n263000 );
nand ( n276052 , n276051 , n263021 );
not ( n276053 , n270115 );
or ( n276054 , n276052 , n276053 );
not ( n276055 , n270110 );
not ( n276056 , n276051 );
or ( n276057 , n276055 , n276056 );
nor ( n276058 , n263021 , n240080 );
nand ( n276059 , n276057 , n276058 );
nand ( n276060 , n255116 , n25998 );
nand ( n276061 , n276054 , n276059 , n276060 );
buf ( n276062 , n276061 );
not ( n276063 , n252015 );
not ( n276064 , n49617 );
or ( n276065 , n276063 , n276064 );
not ( n276066 , n252015 );
nand ( n276067 , n276066 , n49626 );
nand ( n276068 , n276065 , n276067 );
and ( n276069 , n276068 , n253265 );
not ( n276070 , n276068 );
and ( n276071 , n276070 , n253272 );
nor ( n276072 , n276069 , n276071 );
not ( n276073 , n276072 );
buf ( n276074 , n249891 );
and ( n276075 , n276074 , n242911 );
not ( n276076 , n276074 );
and ( n276077 , n276076 , n227707 );
nor ( n276078 , n276075 , n276077 );
and ( n276079 , n276078 , n242978 );
not ( n276080 , n276078 );
and ( n276081 , n276080 , n242970 );
nor ( n276082 , n276079 , n276081 );
nand ( n276083 , n276073 , n276082 );
not ( n276084 , n258077 );
not ( n276085 , n52890 );
not ( n276086 , n276085 );
not ( n276087 , n246882 );
or ( n276088 , n276086 , n276087 );
nand ( n276089 , n246891 , n52890 );
nand ( n276090 , n276088 , n276089 );
not ( n276091 , n276090 );
or ( n276092 , n276084 , n276091 );
or ( n276093 , n258077 , n276090 );
nand ( n276094 , n276092 , n276093 );
nor ( n276095 , n276094 , n249531 );
not ( n276096 , n276095 );
or ( n276097 , n276083 , n276096 );
not ( n276098 , n276094 );
nor ( n276099 , n276098 , n262719 );
nand ( n276100 , n276083 , n276099 );
nand ( n276101 , n245414 , n28333 );
nand ( n276102 , n276097 , n276100 , n276101 );
buf ( n276103 , n276102 );
buf ( n276104 , n54837 );
not ( n276105 , n276104 );
not ( n276106 , n237944 );
or ( n276107 , n276105 , n276106 );
or ( n276108 , n237944 , n276104 );
nand ( n276109 , n276107 , n276108 );
not ( n276110 , n276109 );
not ( n276111 , n256042 );
and ( n276112 , n276110 , n276111 );
and ( n276113 , n276109 , n237947 );
nor ( n276114 , n276112 , n276113 );
nor ( n276115 , n276114 , n252679 );
not ( n276116 , n276115 );
not ( n276117 , n250009 );
not ( n276118 , n276117 );
not ( n276119 , n228527 );
or ( n276120 , n276118 , n276119 );
not ( n276121 , n276117 );
nand ( n276122 , n276121 , n50776 );
nand ( n276123 , n276120 , n276122 );
and ( n276124 , n276123 , n50931 );
not ( n276125 , n276123 );
and ( n276126 , n276125 , n50941 );
nor ( n276127 , n276124 , n276126 );
not ( n276128 , n276127 );
nand ( n276129 , n274572 , n276128 );
or ( n276130 , n276116 , n276129 );
not ( n276131 , n276128 );
not ( n276132 , n276114 );
not ( n276133 , n276132 );
or ( n276134 , n276131 , n276133 );
nor ( n276135 , n274572 , n264469 );
nand ( n276136 , n276134 , n276135 );
nand ( n276137 , n234024 , n31359 );
nand ( n276138 , n276130 , n276136 , n276137 );
buf ( n276139 , n276138 );
buf ( n276140 , n30062 );
buf ( n276141 , n30482 );
buf ( n276142 , n25672 );
not ( n276143 , n266761 );
nand ( n276144 , n276143 , n258088 );
or ( n276145 , n266753 , n276144 );
not ( n276146 , n276143 );
not ( n276147 , n258063 );
or ( n276148 , n276146 , n276147 );
nand ( n276149 , n276148 , n266608 );
nand ( n276150 , n35431 , n36785 );
nand ( n276151 , n276145 , n276149 , n276150 );
buf ( n276152 , n276151 );
not ( n276153 , n31802 );
not ( n276154 , n39766 );
or ( n276155 , n276153 , n276154 );
nand ( n276156 , n259621 , n259353 );
not ( n276157 , n241201 );
and ( n276158 , n276156 , n276157 );
not ( n276159 , n276156 );
and ( n276160 , n276159 , n241201 );
nor ( n276161 , n276158 , n276160 );
or ( n276162 , n276161 , n253358 );
nand ( n276163 , n276155 , n276162 );
buf ( n276164 , n276163 );
not ( n276165 , RI19aa12d0_2559);
or ( n276166 , n25328 , n276165 );
or ( n276167 , n226822 , n273488 );
nand ( n276168 , n276166 , n276167 );
buf ( n276169 , n276168 );
not ( n276170 , n250236 );
not ( n276171 , n276170 );
not ( n276172 , n252658 );
or ( n276173 , n276171 , n276172 );
not ( n276174 , n52532 );
not ( n276175 , n240053 );
or ( n276176 , n276174 , n276175 );
not ( n276177 , n52532 );
nand ( n276178 , n276177 , n240056 );
nand ( n276179 , n276176 , n276178 );
and ( n276180 , n276179 , n274879 );
not ( n276181 , n276179 );
and ( n276182 , n276181 , n269447 );
nor ( n276183 , n276180 , n276182 );
not ( n276184 , n276183 );
nor ( n276185 , n276184 , n252872 );
nand ( n276186 , n276173 , n276185 );
nand ( n276187 , n276184 , n252658 , n250242 );
nand ( n276188 , n252711 , n25724 );
nand ( n276189 , n276186 , n276187 , n276188 );
buf ( n276190 , n276189 );
nand ( n276191 , n269191 , n255152 );
not ( n276192 , n37030 );
not ( n276193 , n240799 );
or ( n276194 , n276192 , n276193 );
not ( n276195 , n37030 );
nand ( n276196 , n276195 , n240810 );
nand ( n276197 , n276194 , n276196 );
and ( n276198 , n276197 , n252447 );
not ( n276199 , n276197 );
and ( n276200 , n276199 , n252444 );
nor ( n276201 , n276198 , n276200 );
not ( n276202 , n276201 );
nand ( n276203 , n268798 , n276202 );
or ( n276204 , n276191 , n276203 );
not ( n276205 , n276202 );
not ( n276206 , n269191 );
or ( n276207 , n276205 , n276206 );
nor ( n276208 , n268798 , n252070 );
nand ( n276209 , n276207 , n276208 );
nand ( n276210 , n50615 , n40383 );
nand ( n276211 , n276204 , n276209 , n276210 );
buf ( n276212 , n276211 );
not ( n276213 , n38486 );
not ( n276214 , n234513 );
or ( n276215 , n276213 , n276214 );
not ( n276216 , n38486 );
nand ( n276217 , n276216 , n234521 );
nand ( n276218 , n276215 , n276217 );
and ( n276219 , n276218 , n243427 );
not ( n276220 , n276218 );
and ( n276221 , n276220 , n243431 );
nor ( n276222 , n276219 , n276221 );
not ( n276223 , n276222 );
nand ( n276224 , n259268 , n276223 );
not ( n276225 , n259256 );
nand ( n276226 , n276224 , n276225 , n250111 );
nor ( n276227 , n276222 , n235050 );
nand ( n276228 , n276227 , n259256 , n259268 );
nand ( n276229 , n31577 , n36791 );
nand ( n276230 , n276226 , n276228 , n276229 );
buf ( n276231 , n276230 );
not ( n276232 , n269965 );
not ( n276233 , n47062 );
not ( n276234 , n252823 );
or ( n276235 , n276233 , n276234 );
not ( n276236 , n47062 );
nand ( n276237 , n276236 , n252831 );
nand ( n276238 , n276235 , n276237 );
and ( n276239 , n276238 , n252837 );
not ( n276240 , n276238 );
and ( n276241 , n276240 , n252834 );
nor ( n276242 , n276239 , n276241 );
not ( n276243 , n276242 );
not ( n276244 , n230818 );
not ( n276245 , n42149 );
or ( n276246 , n276244 , n276245 );
not ( n276247 , n230818 );
nand ( n276248 , n276247 , n42156 );
nand ( n276249 , n276246 , n276248 );
and ( n276250 , n276249 , n220201 );
not ( n276251 , n276249 );
and ( n276252 , n276251 , n259553 );
nor ( n276253 , n276250 , n276252 );
nor ( n276254 , n276243 , n276253 );
or ( n276255 , n276232 , n276254 );
nor ( n276256 , n269963 , n247212 );
nand ( n276257 , n276256 , n276254 );
nand ( n276258 , n234453 , n29271 );
nand ( n276259 , n276255 , n276257 , n276258 );
buf ( n276260 , n276259 );
not ( n276261 , n271550 );
nand ( n276262 , n276261 , n267923 );
or ( n276263 , n276262 , n271553 );
not ( n276264 , n271552 );
not ( n276265 , n276261 );
or ( n276266 , n276264 , n276265 );
nand ( n276267 , n276266 , n267924 );
nand ( n276268 , n246460 , n29308 );
nand ( n276269 , n276263 , n276267 , n276268 );
buf ( n276270 , n276269 );
not ( n276271 , n244838 );
nand ( n276272 , n262482 , n262496 );
or ( n276273 , n276271 , n276272 );
not ( n276274 , n244830 );
not ( n276275 , n276274 );
not ( n276276 , n262482 );
or ( n276277 , n276275 , n276276 );
nor ( n276278 , n262496 , n235050 );
nand ( n276279 , n276277 , n276278 );
nand ( n276280 , n35431 , n32375 );
nand ( n276281 , n276273 , n276279 , n276280 );
buf ( n276282 , n276281 );
not ( n276283 , n270430 );
nand ( n276284 , n276283 , n246177 );
nand ( n276285 , n273069 , n270420 );
or ( n276286 , n276284 , n276285 );
not ( n276287 , n270420 );
not ( n276288 , n276283 );
or ( n276289 , n276287 , n276288 );
nor ( n276290 , n273069 , n55104 );
nand ( n276291 , n276289 , n276290 );
nand ( n276292 , n245414 , n25672 );
nand ( n276293 , n276286 , n276291 , n276292 );
buf ( n276294 , n276293 );
nand ( n276295 , n257538 , n260879 );
buf ( n276296 , n246843 );
not ( n276297 , n276296 );
not ( n276298 , n242852 );
or ( n276299 , n276297 , n276298 );
or ( n276300 , n242860 , n276296 );
nand ( n276301 , n276299 , n276300 );
not ( n276302 , n276301 );
not ( n276303 , n261185 );
and ( n276304 , n276302 , n276303 );
and ( n276305 , n276301 , n242867 );
nor ( n276306 , n276304 , n276305 );
nand ( n276307 , n276306 , n257550 );
or ( n276308 , n276295 , n276307 );
not ( n276309 , n257550 );
not ( n276310 , n257538 );
or ( n276311 , n276309 , n276310 );
nor ( n276312 , n276306 , n233972 );
nand ( n276313 , n276311 , n276312 );
nand ( n276314 , n241068 , n34973 );
nand ( n276315 , n276308 , n276313 , n276314 );
buf ( n276316 , n276315 );
not ( n276317 , n262735 );
nand ( n276318 , n276317 , n262757 );
nand ( n276319 , n276318 , n265563 , n226010 );
nand ( n276320 , n265564 , n275391 , n262757 );
nand ( n276321 , n35431 , n204770 );
nand ( n276322 , n276319 , n276320 , n276321 );
buf ( n276323 , n276322 );
not ( n276324 , n33965 );
not ( n276325 , n244190 );
or ( n276326 , n276324 , n276325 );
not ( n276327 , n33965 );
nand ( n276328 , n276327 , n244199 );
nand ( n276329 , n276326 , n276328 );
and ( n276330 , n276329 , n244208 );
not ( n276331 , n276329 );
and ( n276332 , n276331 , n244204 );
nor ( n276333 , n276330 , n276332 );
nor ( n276334 , n276333 , n219702 );
not ( n276335 , n47990 );
not ( n276336 , n48676 );
or ( n276337 , n276335 , n276336 );
not ( n276338 , n47990 );
nand ( n276339 , n276338 , n48686 );
nand ( n276340 , n276337 , n276339 );
and ( n276341 , n276340 , n48797 );
not ( n276342 , n276340 );
and ( n276343 , n276342 , n48806 );
nor ( n276344 , n276341 , n276343 );
not ( n276345 , n276344 );
nor ( n276346 , n276345 , n275932 );
nand ( n276347 , n276334 , n276346 );
not ( n276348 , n275929 );
not ( n276349 , n276333 );
not ( n276350 , n276349 );
or ( n276351 , n276348 , n276350 );
nor ( n276352 , n276344 , n33254 );
nand ( n276353 , n276351 , n276352 );
nand ( n276354 , n35431 , n204797 );
nand ( n276355 , n276347 , n276353 , n276354 );
buf ( n276356 , n276355 );
not ( n276357 , n234871 );
not ( n276358 , n276357 );
not ( n276359 , n225525 );
or ( n276360 , n276358 , n276359 );
not ( n276361 , n276357 );
nand ( n276362 , n276361 , n47773 );
nand ( n276363 , n276360 , n276362 );
and ( n276364 , n276363 , n262494 );
not ( n276365 , n276363 );
and ( n276366 , n276365 , n246207 );
nor ( n276367 , n276364 , n276366 );
nor ( n276368 , n276367 , n234021 );
not ( n276369 , n274883 );
nand ( n276370 , n276368 , n276369 , n255307 );
not ( n276371 , n276367 );
not ( n276372 , n276371 );
not ( n276373 , n276369 );
or ( n276374 , n276372 , n276373 );
nor ( n276375 , n255307 , n251190 );
nand ( n276376 , n276374 , n276375 );
nand ( n276377 , n31577 , n37860 );
nand ( n276378 , n276370 , n276376 , n276377 );
buf ( n276379 , n276378 );
or ( n276380 , n25328 , n268940 );
or ( n276381 , n226822 , n260456 );
nand ( n276382 , n276380 , n276381 );
buf ( n276383 , n276382 );
nand ( n276384 , n251316 , n237385 );
not ( n276385 , n233875 );
not ( n276386 , n276385 );
not ( n276387 , n244282 );
or ( n276388 , n276386 , n276387 );
or ( n276389 , n244282 , n276385 );
nand ( n276390 , n276388 , n276389 );
and ( n276391 , n276390 , n244347 );
not ( n276392 , n276390 );
and ( n276393 , n276392 , n258153 );
nor ( n276394 , n276391 , n276393 );
nand ( n276395 , n276394 , n251355 );
or ( n276396 , n276384 , n276395 );
not ( n276397 , n276394 );
not ( n276398 , n251316 );
or ( n276399 , n276397 , n276398 );
nor ( n276400 , n251355 , n55104 );
nand ( n276401 , n276399 , n276400 );
nand ( n276402 , n234448 , n45199 );
nand ( n276403 , n276396 , n276401 , n276402 );
buf ( n276404 , n276403 );
nand ( n276405 , n276082 , n276072 );
not ( n276406 , n228471 );
not ( n276407 , n237867 );
or ( n276408 , n276406 , n276407 );
not ( n276409 , n228471 );
nand ( n276410 , n276409 , n255503 );
nand ( n276411 , n276408 , n276410 );
and ( n276412 , n276411 , n265402 );
not ( n276413 , n276411 );
and ( n276414 , n276413 , n255515 );
nor ( n276415 , n276412 , n276414 );
nand ( n276416 , n276415 , n250111 );
or ( n276417 , n276405 , n276416 );
not ( n276418 , n276415 );
not ( n276419 , n276072 );
or ( n276420 , n276418 , n276419 );
nor ( n276421 , n276082 , n260567 );
nand ( n276422 , n276420 , n276421 );
nand ( n276423 , n55760 , n28303 );
nand ( n276424 , n276417 , n276422 , n276423 );
buf ( n276425 , n276424 );
buf ( n276426 , RI19a24a28_2784);
not ( n276427 , n276426 );
not ( n276428 , n257347 );
or ( n276429 , n276427 , n276428 );
nand ( n276430 , n257351 , n268968 );
nand ( n276431 , n276429 , n276430 );
buf ( n276432 , n276431 );
not ( n276433 , n32221 );
not ( n276434 , n252711 );
or ( n276435 , n276433 , n276434 );
nand ( n276436 , n253735 , n253748 );
and ( n276437 , n276436 , n274236 );
not ( n276438 , n276436 );
and ( n276439 , n276438 , n256272 );
nor ( n276440 , n276437 , n276439 );
or ( n276441 , n276440 , n258759 );
nand ( n276442 , n276435 , n276441 );
buf ( n276443 , n276442 );
not ( n276444 , n55301 );
not ( n276445 , n53077 );
or ( n276446 , n276444 , n276445 );
or ( n276447 , n53081 , n55301 );
nand ( n276448 , n276446 , n276447 );
not ( n276449 , n276448 );
not ( n276450 , n230903 );
and ( n276451 , n276449 , n276450 );
and ( n276452 , n276448 , n230906 );
nor ( n276453 , n276451 , n276452 );
not ( n276454 , n273912 );
nand ( n276455 , n276453 , n276454 );
or ( n276456 , n267987 , n276455 );
not ( n276457 , n276454 );
not ( n276458 , n267970 );
or ( n276459 , n276457 , n276458 );
nor ( n276460 , n276453 , n234440 );
nand ( n276461 , n276459 , n276460 );
nand ( n276462 , n244987 , n26344 );
nand ( n276463 , n276456 , n276461 , n276462 );
buf ( n276464 , n276463 );
not ( n276465 , n247252 );
nand ( n276466 , n262108 , n276465 );
or ( n276467 , n247240 , n276466 );
not ( n276468 , n276465 );
not ( n276469 , n247239 );
or ( n276470 , n276468 , n276469 );
nor ( n276471 , n262108 , n50944 );
nand ( n276472 , n276470 , n276471 );
nand ( n276473 , n237361 , n28552 );
nand ( n276474 , n276467 , n276472 , n276473 );
buf ( n276475 , n276474 );
not ( n276476 , n238188 );
nand ( n276477 , n238217 , n276476 );
not ( n276478 , n271301 );
or ( n276479 , n276477 , n276478 );
not ( n276480 , n271298 );
nor ( n276481 , n276480 , n219702 );
nand ( n276482 , n276477 , n276481 );
nand ( n276483 , n253486 , n29929 );
nand ( n276484 , n276479 , n276482 , n276483 );
buf ( n276485 , n276484 );
buf ( n276486 , n36284 );
buf ( n276487 , n34132 );
not ( n276488 , n260959 );
not ( n276489 , n275302 );
nand ( n276490 , n276488 , n276489 );
or ( n276491 , n260947 , n276490 );
not ( n276492 , n276488 );
not ( n276493 , n260946 );
or ( n276494 , n276492 , n276493 );
nor ( n276495 , n276489 , n236795 );
nand ( n276496 , n276494 , n276495 );
nand ( n276497 , n247423 , n25907 );
nand ( n276498 , n276491 , n276496 , n276497 );
buf ( n276499 , n276498 );
buf ( n276500 , n29112 );
buf ( n276501 , n33880 );
not ( n276502 , n260236 );
not ( n276503 , n276502 );
not ( n276504 , n260219 );
or ( n276505 , n276503 , n276504 );
not ( n276506 , n246069 );
nand ( n276507 , n276505 , n276506 );
nor ( n276508 , n260218 , n254150 );
nor ( n276509 , n276506 , n246085 );
and ( n276510 , n276508 , n276509 );
and ( n276511 , n48251 , n38317 );
nor ( n276512 , n276510 , n276511 );
nand ( n276513 , n276507 , n276512 );
buf ( n276514 , n276513 );
not ( n276515 , RI19ac7250_2276);
or ( n276516 , n25328 , n276515 );
not ( n276517 , RI19abe4c0_2347);
or ( n276518 , n226822 , n276517 );
nand ( n276519 , n276516 , n276518 );
buf ( n276520 , n276519 );
not ( n276521 , n256980 );
not ( n276522 , n256955 );
or ( n276523 , n276521 , n276522 );
nand ( n276524 , n276523 , n260879 );
or ( n276525 , n276524 , n260994 );
nand ( n276526 , n256955 , n226010 );
nand ( n276527 , n260994 , n256980 );
or ( n276528 , n276526 , n276527 );
nand ( n276529 , n39766 , n30825 );
nand ( n276530 , n276525 , n276528 , n276529 );
buf ( n276531 , n276530 );
not ( n276532 , n260975 );
not ( n276533 , n264275 );
nand ( n276534 , n276489 , n276533 );
or ( n276535 , n276532 , n276534 );
not ( n276536 , n276489 );
not ( n276537 , n260946 );
not ( n276538 , n276537 );
or ( n276539 , n276536 , n276538 );
nor ( n276540 , n276533 , n226004 );
nand ( n276541 , n276539 , n276540 );
nand ( n276542 , n246460 , n209722 );
nand ( n276543 , n276535 , n276541 , n276542 );
buf ( n276544 , n276543 );
not ( n276545 , n27769 );
not ( n276546 , n244789 );
or ( n276547 , n276545 , n276546 );
nand ( n276548 , n269988 , n269985 );
not ( n276549 , n276253 );
and ( n276550 , n276548 , n276549 );
not ( n276551 , n276548 );
and ( n276552 , n276551 , n276253 );
nor ( n276553 , n276550 , n276552 );
or ( n276554 , n276553 , n255135 );
nand ( n276555 , n276547 , n276554 );
buf ( n276556 , n276555 );
not ( n276557 , RI19aaac18_2490);
or ( n276558 , n25328 , n276557 );
not ( n276559 , RI19aa0d30_2562);
or ( n276560 , n25336 , n276559 );
nand ( n276561 , n276558 , n276560 );
buf ( n276562 , n276561 );
not ( n276563 , n263695 );
not ( n276564 , n275537 );
not ( n276565 , n276564 );
or ( n276566 , n276563 , n276565 );
nor ( n276567 , n263682 , n250909 );
nand ( n276568 , n276566 , n276567 );
not ( n276569 , n263696 );
nand ( n276570 , n276564 , n276569 , n263682 );
nand ( n276571 , n256292 , n32514 );
nand ( n276572 , n276568 , n276570 , n276571 );
buf ( n276573 , n276572 );
not ( n276574 , n262294 );
nand ( n276575 , n276574 , n253928 );
not ( n276576 , n256355 );
nand ( n276577 , n256345 , n276576 );
or ( n276578 , n276575 , n276577 );
not ( n276579 , n276576 );
not ( n276580 , n276574 );
or ( n276581 , n276579 , n276580 );
nor ( n276582 , n256345 , n53680 );
nand ( n276583 , n276581 , n276582 );
nand ( n276584 , n39767 , n230663 );
nand ( n276585 , n276578 , n276583 , n276584 );
buf ( n276586 , n276585 );
nand ( n276587 , n272448 , n262712 );
or ( n276588 , n273479 , n276587 );
not ( n276589 , n272448 );
not ( n276590 , n262688 );
or ( n276591 , n276589 , n276590 );
not ( n276592 , n255152 );
nor ( n276593 , n262712 , n276592 );
nand ( n276594 , n276591 , n276593 );
nand ( n276595 , n241068 , n25646 );
nand ( n276596 , n276588 , n276594 , n276595 );
buf ( n276597 , n276596 );
buf ( n276598 , n46583 );
buf ( n276599 , n38428 );
buf ( n276600 , n26043 );
nand ( n276601 , n45264 , n250302 );
or ( n276602 , n223840 , n276601 );
not ( n276603 , n46077 );
not ( n276604 , n45264 );
or ( n276605 , n276603 , n276604 );
nand ( n276606 , n276605 , n250303 );
nand ( n276607 , n250916 , n27937 );
nand ( n276608 , n276602 , n276606 , n276607 );
buf ( n276609 , n276608 );
buf ( n276610 , n28103 );
not ( n276611 , n37446 );
not ( n276612 , n51381 );
or ( n276613 , n276611 , n276612 );
not ( n276614 , n250400 );
not ( n276615 , n42382 );
not ( n276616 , n234305 );
or ( n276617 , n276615 , n276616 );
not ( n276618 , n42382 );
nand ( n276619 , n276618 , n234298 );
nand ( n276620 , n276617 , n276619 );
and ( n276621 , n276620 , n256932 );
not ( n276622 , n276620 );
and ( n276623 , n276622 , n256928 );
nor ( n276624 , n276621 , n276623 );
not ( n276625 , n276624 );
nand ( n276626 , n276614 , n276625 );
and ( n276627 , n276626 , n269154 );
not ( n276628 , n276626 );
and ( n276629 , n276628 , n250414 );
nor ( n276630 , n276627 , n276629 );
or ( n276631 , n276630 , n256376 );
nand ( n276632 , n276613 , n276631 );
buf ( n276633 , n276632 );
not ( n276634 , RI19a9a3b8_2610);
or ( n276635 , n25328 , n276634 );
not ( n276636 , RI19a90188_2682);
or ( n276637 , n25336 , n276636 );
nand ( n276638 , n276635 , n276637 );
buf ( n276639 , n276638 );
not ( n276640 , n221883 );
not ( n276641 , n46083 );
or ( n276642 , n276640 , n276641 );
not ( n276643 , n258076 );
nand ( n276644 , n276643 , n266619 );
and ( n276645 , n276644 , n276143 );
not ( n276646 , n276644 );
and ( n276647 , n276646 , n266761 );
nor ( n276648 , n276645 , n276647 );
or ( n276649 , n276648 , n244217 );
nand ( n276650 , n276642 , n276649 );
buf ( n276651 , n276650 );
not ( n276652 , n261193 );
nor ( n276653 , n276652 , n252070 );
not ( n276654 , n276653 );
not ( n276655 , n261181 );
nand ( n276656 , n276655 , n270083 );
or ( n276657 , n276654 , n276656 );
not ( n276658 , n276655 );
not ( n276659 , n261193 );
or ( n276660 , n276658 , n276659 );
nor ( n276661 , n270083 , n54208 );
nand ( n276662 , n276660 , n276661 );
nand ( n276663 , n31577 , n29673 );
nand ( n276664 , n276657 , n276662 , n276663 );
buf ( n276665 , n276664 );
buf ( n276666 , n30017 );
buf ( n276667 , n26129 );
buf ( n276668 , n35150 );
or ( n276669 , n25328 , n261253 );
or ( n276670 , n25335 , n273094 );
nand ( n276671 , n276669 , n276670 );
buf ( n276672 , n276671 );
nand ( n276673 , n258044 , n265594 );
or ( n276674 , n272407 , n276673 );
nand ( n276675 , n249098 , n276673 );
nand ( n276676 , n247423 , n29582 );
nand ( n276677 , n276674 , n276675 , n276676 );
buf ( n276678 , n276677 );
buf ( n276679 , n29546 );
buf ( n276680 , n30193 );
buf ( n276681 , n205306 );
not ( n276682 , n235861 );
not ( n276683 , n245797 );
or ( n276684 , n276682 , n276683 );
or ( n276685 , n263379 , n235861 );
nand ( n276686 , n276684 , n276685 );
and ( n276687 , n276686 , n250813 );
not ( n276688 , n276686 );
and ( n276689 , n276688 , n263382 );
nor ( n276690 , n276687 , n276689 );
not ( n276691 , n276690 );
nand ( n276692 , n276691 , n252259 );
not ( n276693 , n247957 );
not ( n276694 , n239930 );
or ( n276695 , n276693 , n276694 );
not ( n276696 , n247957 );
nand ( n276697 , n276696 , n239922 );
nand ( n276698 , n276695 , n276697 );
and ( n276699 , n276698 , n243504 );
not ( n276700 , n276698 );
and ( n276701 , n276700 , n243511 );
nor ( n276702 , n276699 , n276701 );
not ( n276703 , n276702 );
nand ( n276704 , n268633 , n276703 );
or ( n276705 , n276692 , n276704 );
not ( n276706 , n268633 );
not ( n276707 , n276691 );
or ( n276708 , n276706 , n276707 );
nor ( n276709 , n276703 , n250909 );
nand ( n276710 , n276708 , n276709 );
nand ( n276711 , n50615 , n41736 );
nand ( n276712 , n276705 , n276710 , n276711 );
buf ( n276713 , n276712 );
not ( n276714 , n206513 );
not ( n276715 , n51381 );
or ( n276716 , n276714 , n276715 );
not ( n276717 , n272341 );
nand ( n276718 , n276717 , n261507 );
and ( n276719 , n276718 , n261518 );
not ( n276720 , n276718 );
and ( n276721 , n276720 , n261519 );
nor ( n276722 , n276719 , n276721 );
or ( n276723 , n276722 , n258280 );
nand ( n276724 , n276716 , n276723 );
buf ( n276725 , n276724 );
buf ( n276726 , n205372 );
not ( n276727 , n274582 );
nand ( n276728 , n276727 , n276114 );
or ( n276729 , n274593 , n276728 );
not ( n276730 , n276727 );
not ( n276731 , n274592 );
or ( n276732 , n276730 , n276731 );
nand ( n276733 , n276732 , n276115 );
nand ( n276734 , n231444 , n40873 );
nand ( n276735 , n276729 , n276733 , n276734 );
buf ( n276736 , n276735 );
not ( n276737 , n234036 );
not ( n276738 , n39766 );
or ( n276739 , n276737 , n276738 );
not ( n276740 , n228908 );
not ( n276741 , n276740 );
not ( n276742 , n257184 );
or ( n276743 , n276741 , n276742 );
nand ( n276744 , n255762 , n228908 );
nand ( n276745 , n276743 , n276744 );
not ( n276746 , n276745 );
not ( n276747 , n255814 );
and ( n276748 , n276746 , n276747 );
and ( n276749 , n276745 , n255810 );
nor ( n276750 , n276748 , n276749 );
buf ( n276751 , n245496 );
not ( n276752 , n276751 );
not ( n276753 , n276752 );
not ( n276754 , n55066 );
or ( n276755 , n276753 , n276754 );
nand ( n276756 , n241893 , n276751 );
nand ( n276757 , n276755 , n276756 );
not ( n276758 , n276757 );
not ( n276759 , n241963 );
or ( n276760 , n276758 , n276759 );
or ( n276761 , n261037 , n276757 );
nand ( n276762 , n276760 , n276761 );
nand ( n276763 , n276750 , n276762 );
not ( n276764 , n276763 );
buf ( n276765 , n254687 );
not ( n276766 , n276765 );
not ( n276767 , n249610 );
or ( n276768 , n276766 , n276767 );
or ( n276769 , n249610 , n276765 );
nand ( n276770 , n276768 , n276769 );
and ( n276771 , n276770 , n265476 );
not ( n276772 , n276770 );
and ( n276773 , n276772 , n250234 );
nor ( n276774 , n276771 , n276773 );
not ( n276775 , n276774 );
and ( n276776 , n276764 , n276775 );
and ( n276777 , n276763 , n276774 );
nor ( n276778 , n276776 , n276777 );
or ( n276779 , n276778 , n234818 );
nand ( n276780 , n276739 , n276779 );
buf ( n276781 , n276780 );
nand ( n276782 , n254162 , n258918 );
nand ( n276783 , n271134 , n254173 );
or ( n276784 , n276782 , n276783 );
not ( n276785 , n254173 );
not ( n276786 , n254162 );
or ( n276787 , n276785 , n276786 );
nor ( n276788 , n271134 , n251190 );
nand ( n276789 , n276787 , n276788 );
nand ( n276790 , n41945 , n235505 );
nand ( n276791 , n276784 , n276789 , n276790 );
buf ( n276792 , n276791 );
not ( n276793 , n25436 );
not ( n276794 , n234453 );
or ( n276795 , n276793 , n276794 );
not ( n276796 , n205228 );
not ( n276797 , n276796 );
not ( n276798 , n228364 );
or ( n276799 , n276797 , n276798 );
not ( n276800 , n276796 );
nand ( n276801 , n276800 , n50539 );
nand ( n276802 , n276799 , n276801 );
and ( n276803 , n276802 , n55726 );
not ( n276804 , n276802 );
and ( n276805 , n276804 , n55727 );
nor ( n276806 , n276803 , n276805 );
not ( n276807 , n276806 );
nand ( n276808 , n276807 , n272284 );
and ( n276809 , n276808 , n269148 );
not ( n276810 , n276808 );
and ( n276811 , n276810 , n269134 );
nor ( n276812 , n276809 , n276811 );
or ( n276813 , n276812 , n254882 );
nand ( n276814 , n276795 , n276813 );
buf ( n276815 , n276814 );
or ( n276816 , n226819 , n262552 );
not ( n276817 , RI19a93068_2661);
or ( n276818 , n25336 , n276817 );
nand ( n276819 , n276816 , n276818 );
buf ( n276820 , n276819 );
not ( n276821 , n34038 );
not ( n276822 , n51381 );
or ( n276823 , n276821 , n276822 );
buf ( n276824 , n251292 );
not ( n276825 , n276824 );
not ( n276826 , n249939 );
or ( n276827 , n276825 , n276826 );
or ( n276828 , n242574 , n276824 );
nand ( n276829 , n276827 , n276828 );
not ( n276830 , n276829 );
not ( n276831 , n276830 );
not ( n276832 , n267247 );
or ( n276833 , n276831 , n276832 );
nand ( n276834 , n249929 , n276829 );
nand ( n276835 , n276833 , n276834 );
not ( n276836 , n276835 );
nand ( n276837 , n276836 , n255934 );
not ( n276838 , n47758 );
not ( n276839 , n238033 );
or ( n276840 , n276838 , n276839 );
not ( n276841 , n47758 );
nand ( n276842 , n276841 , n238040 );
nand ( n276843 , n276840 , n276842 );
not ( n276844 , n276843 );
not ( n276845 , n238102 );
and ( n276846 , n276844 , n276845 );
and ( n276847 , n276843 , n238102 );
nor ( n276848 , n276846 , n276847 );
not ( n276849 , n276848 );
and ( n276850 , n276837 , n276849 );
not ( n276851 , n276837 );
and ( n276852 , n276851 , n276848 );
nor ( n276853 , n276850 , n276852 );
or ( n276854 , n276853 , n251498 );
nand ( n276855 , n276823 , n276854 );
buf ( n276856 , n276855 );
buf ( n276857 , n248644 );
not ( n276858 , n276857 );
not ( n276859 , n251855 );
or ( n276860 , n276858 , n276859 );
or ( n276861 , n251855 , n276857 );
nand ( n276862 , n276860 , n276861 );
and ( n276863 , n276862 , n267341 );
not ( n276864 , n276862 );
and ( n276865 , n276864 , n260967 );
nor ( n276866 , n276863 , n276865 );
nor ( n276867 , n276866 , n252679 );
not ( n276868 , n276774 );
not ( n276869 , n239270 );
not ( n276870 , n276869 );
not ( n276871 , n248755 );
or ( n276872 , n276870 , n276871 );
not ( n276873 , n276869 );
nand ( n276874 , n276873 , n248762 );
nand ( n276875 , n276872 , n276874 );
and ( n276876 , n276875 , n252919 );
not ( n276877 , n276875 );
and ( n276878 , n276877 , n252924 );
nor ( n276879 , n276876 , n276878 );
nor ( n276880 , n276868 , n276879 );
nand ( n276881 , n276867 , n276880 );
not ( n276882 , n276774 );
not ( n276883 , n276866 );
not ( n276884 , n276883 );
or ( n276885 , n276882 , n276884 );
not ( n276886 , n276879 );
nor ( n276887 , n276886 , n243434 );
nand ( n276888 , n276885 , n276887 );
nand ( n276889 , n55760 , n29245 );
nand ( n276890 , n276881 , n276888 , n276889 );
buf ( n276891 , n276890 );
nand ( n276892 , n254649 , n254661 );
not ( n276893 , n275975 );
or ( n276894 , n276892 , n276893 );
nor ( n276895 , n275967 , n35427 );
nand ( n276896 , n276892 , n276895 );
nand ( n276897 , n39767 , n38279 );
nand ( n276898 , n276894 , n276896 , n276897 );
buf ( n276899 , n276898 );
buf ( n276900 , n235193 );
not ( n276901 , n276900 );
not ( n276902 , n276901 );
not ( n276903 , n248446 );
or ( n276904 , n276902 , n276903 );
nand ( n276905 , n248455 , n276900 );
nand ( n276906 , n276904 , n276905 );
not ( n276907 , n276906 );
not ( n276908 , n248386 );
and ( n276909 , n276907 , n276908 );
and ( n276910 , n276906 , n248386 );
nor ( n276911 , n276909 , n276910 );
not ( n276912 , n251037 );
not ( n276913 , n50482 );
or ( n276914 , n276912 , n276913 );
or ( n276915 , n50482 , n251037 );
nand ( n276916 , n276914 , n276915 );
and ( n276917 , n276916 , n263851 );
not ( n276918 , n276916 );
and ( n276919 , n276918 , n263848 );
nor ( n276920 , n276917 , n276919 );
nand ( n276921 , n276911 , n276920 );
not ( n276922 , n260125 );
not ( n276923 , n239566 );
not ( n276924 , n260112 );
or ( n276925 , n276923 , n276924 );
not ( n276926 , n239566 );
nand ( n276927 , n276926 , n260122 );
nand ( n276928 , n276925 , n276927 );
not ( n276929 , n276928 );
or ( n276930 , n276922 , n276929 );
or ( n276931 , n276928 , n260125 );
nand ( n276932 , n276930 , n276931 );
nor ( n276933 , n276932 , n238635 );
not ( n276934 , n276933 );
or ( n276935 , n276921 , n276934 );
not ( n276936 , n276932 );
nor ( n276937 , n276936 , n234440 );
nand ( n276938 , n276921 , n276937 );
nand ( n276939 , n238114 , n29905 );
nand ( n276940 , n276935 , n276938 , n276939 );
buf ( n276941 , n276940 );
not ( n276942 , n37340 );
not ( n276943 , n234453 );
or ( n276944 , n276942 , n276943 );
nand ( n276945 , n262919 , n261576 );
not ( n276946 , n262931 );
and ( n276947 , n276945 , n276946 );
not ( n276948 , n276945 );
and ( n276949 , n276948 , n262931 );
nor ( n276950 , n276947 , n276949 );
or ( n276951 , n276950 , n253544 );
nand ( n276952 , n276944 , n276951 );
buf ( n276953 , n276952 );
or ( n276954 , n25328 , n266718 );
or ( n276955 , n25335 , n256085 );
nand ( n276956 , n276954 , n276955 );
buf ( n276957 , n276956 );
or ( n276958 , n226819 , n262139 );
or ( n276959 , n25335 , n268830 );
nand ( n276960 , n276958 , n276959 );
buf ( n276961 , n276960 );
not ( n276962 , RI19aa40c0_2537);
or ( n276963 , n25328 , n276962 );
not ( n276964 , RI19a87470_2743);
or ( n276965 , n226822 , n276964 );
nand ( n276966 , n276963 , n276965 );
buf ( n276967 , n276966 );
not ( n276968 , n241703 );
nand ( n276969 , n276968 , n241888 );
or ( n276970 , n267097 , n276969 );
not ( n276971 , n267096 );
not ( n276972 , n276968 );
or ( n276973 , n276971 , n276972 );
nor ( n276974 , n241888 , n52445 );
nand ( n276975 , n276973 , n276974 );
nand ( n276976 , n50615 , n35872 );
nand ( n276977 , n276970 , n276975 , n276976 );
buf ( n276978 , n276977 );
nand ( n276979 , n260582 , n55147 );
nand ( n276980 , n274907 , n260609 );
or ( n276981 , n276979 , n276980 );
not ( n276982 , n260609 );
not ( n276983 , n260582 );
or ( n276984 , n276982 , n276983 );
nor ( n276985 , n274907 , n49051 );
nand ( n276986 , n276984 , n276985 );
nand ( n276987 , n252711 , n32499 );
nand ( n276988 , n276981 , n276986 , n276987 );
buf ( n276989 , n276988 );
buf ( n276990 , n25886 );
or ( n276991 , n25328 , n259243 );
or ( n276992 , n25335 , n269855 );
nand ( n276993 , n276991 , n276992 );
buf ( n276994 , n276993 );
buf ( n276995 , n207202 );
nand ( n276996 , n253611 , n266742 );
or ( n276997 , n275281 , n276996 );
not ( n276998 , n266742 );
not ( n276999 , n266730 );
or ( n277000 , n276998 , n276999 );
nand ( n277001 , n277000 , n253612 );
nand ( n277002 , n244484 , n26391 );
nand ( n277003 , n276997 , n277001 , n277002 );
buf ( n277004 , n277003 );
not ( n277005 , n255544 );
not ( n277006 , n238628 );
or ( n277007 , n277005 , n277006 );
not ( n277008 , n255544 );
nand ( n277009 , n277008 , n238620 );
nand ( n277010 , n277007 , n277009 );
and ( n277011 , n277010 , n257188 );
not ( n277012 , n277010 );
and ( n277013 , n277012 , n257185 );
nor ( n277014 , n277011 , n277013 );
nor ( n277015 , n277014 , n55104 );
buf ( n277016 , n253798 );
not ( n277017 , n277016 );
not ( n277018 , n250576 );
or ( n277019 , n277017 , n277018 );
or ( n277020 , n250576 , n277016 );
nand ( n277021 , n277019 , n277020 );
and ( n277022 , n277021 , n252052 );
not ( n277023 , n277021 );
and ( n277024 , n277023 , n252037 );
nor ( n277025 , n277022 , n277024 );
nand ( n277026 , n277015 , n277025 , n266400 );
not ( n277027 , n277014 );
not ( n277028 , n277027 );
not ( n277029 , n277025 );
or ( n277030 , n277028 , n277029 );
nand ( n277031 , n277030 , n266404 );
nand ( n277032 , n237714 , n33359 );
nand ( n277033 , n277026 , n277031 , n277032 );
buf ( n277034 , n277033 );
buf ( n277035 , n242012 );
not ( n277036 , n277035 );
not ( n277037 , n255822 );
or ( n277038 , n277036 , n277037 );
or ( n277039 , n246389 , n277035 );
nand ( n277040 , n277038 , n277039 );
and ( n277041 , n277040 , n246449 );
not ( n277042 , n277040 );
and ( n277043 , n277042 , n246441 );
nor ( n277044 , n277041 , n277043 );
nor ( n277045 , n277044 , n43968 );
not ( n277046 , n277045 );
not ( n277047 , n265381 );
nand ( n277048 , n277047 , n265393 );
or ( n277049 , n277046 , n277048 );
not ( n277050 , n277047 );
not ( n277051 , n277044 );
not ( n277052 , n277051 );
or ( n277053 , n277050 , n277052 );
nor ( n277054 , n265393 , n234440 );
nand ( n277055 , n277053 , n277054 );
nand ( n277056 , n241068 , n29104 );
nand ( n277057 , n277049 , n277055 , n277056 );
buf ( n277058 , n277057 );
not ( n277059 , n205902 );
not ( n277060 , n258213 );
or ( n277061 , n277059 , n277060 );
not ( n277062 , n245176 );
nand ( n277063 , n277062 , n245192 );
and ( n277064 , n277063 , n273859 );
not ( n277065 , n277063 );
and ( n277066 , n277065 , n272892 );
nor ( n277067 , n277064 , n277066 );
or ( n277068 , n277067 , n257174 );
nand ( n277069 , n277061 , n277068 );
buf ( n277070 , n277069 );
not ( n277071 , n265886 );
not ( n277072 , n270114 );
or ( n277073 , n277071 , n277072 );
nor ( n277074 , n276051 , n233972 );
nand ( n277075 , n277073 , n277074 );
nand ( n277076 , n270111 , n276051 , n265886 );
nand ( n277077 , n39766 , n32955 );
nand ( n277078 , n277075 , n277076 , n277077 );
buf ( n277079 , n277078 );
not ( n277080 , n45720 );
not ( n277081 , n248210 );
or ( n277082 , n277080 , n277081 );
not ( n277083 , n45720 );
nand ( n277084 , n277083 , n248219 );
nand ( n277085 , n277082 , n277084 );
and ( n277086 , n277085 , n261434 );
not ( n277087 , n277085 );
and ( n277088 , n277087 , n261431 );
nor ( n277089 , n277086 , n277088 );
nor ( n277090 , n277089 , n40465 );
not ( n277091 , n277090 );
not ( n277092 , n264165 );
nand ( n277093 , n277092 , n261146 );
or ( n277094 , n277091 , n277093 );
not ( n277095 , n277089 );
not ( n277096 , n277095 );
not ( n277097 , n277092 );
or ( n277098 , n277096 , n277097 );
nor ( n277099 , n261146 , n31572 );
nand ( n277100 , n277098 , n277099 );
nand ( n277101 , n35431 , n39615 );
nand ( n277102 , n277094 , n277100 , n277101 );
buf ( n277103 , n277102 );
not ( n277104 , n266378 );
not ( n277105 , n277025 );
nand ( n277106 , n277104 , n277105 );
not ( n277107 , n277015 );
or ( n277108 , n277106 , n277107 );
nor ( n277109 , n277027 , n49959 );
nand ( n277110 , n277106 , n277109 );
nand ( n277111 , n31577 , n29283 );
nand ( n277112 , n277108 , n277110 , n277111 );
buf ( n277113 , n277112 );
not ( n277114 , RI19a85760_2756);
or ( n277115 , n233507 , n277114 );
or ( n277116 , n25335 , n275418 );
nand ( n277117 , n277115 , n277116 );
buf ( n277118 , n277117 );
buf ( n277119 , n35771 );
buf ( n277120 , n35082 );
buf ( n277121 , n30426 );
nand ( n277122 , n273543 , n270602 );
not ( n277123 , n243321 );
not ( n277124 , n250805 );
or ( n277125 , n277123 , n277124 );
not ( n277126 , n243321 );
nand ( n277127 , n277126 , n250806 );
nand ( n277128 , n277125 , n277127 );
and ( n277129 , n277128 , n257382 );
not ( n277130 , n277128 );
and ( n277131 , n277130 , n257379 );
nor ( n277132 , n277129 , n277131 );
nor ( n277133 , n277132 , n226003 );
not ( n277134 , n277133 );
or ( n277135 , n277122 , n277134 );
not ( n277136 , n277132 );
nor ( n277137 , n277136 , n50944 );
nand ( n277138 , n277122 , n277137 );
nand ( n277139 , n241976 , n31201 );
nand ( n277140 , n277135 , n277138 , n277139 );
buf ( n277141 , n277140 );
nand ( n277142 , n267131 , n235051 );
nand ( n277143 , n274021 , n267145 );
or ( n277144 , n277142 , n277143 );
not ( n277145 , n267145 );
not ( n277146 , n267131 );
or ( n277147 , n277145 , n277146 );
nor ( n277148 , n274021 , n236795 );
nand ( n277149 , n277147 , n277148 );
nand ( n277150 , n55760 , n37636 );
nand ( n277151 , n277144 , n277149 , n277150 );
buf ( n277152 , n277151 );
not ( n277153 , n34132 );
not ( n277154 , n37728 );
or ( n277155 , n277153 , n277154 );
not ( n277156 , n273069 );
nand ( n277157 , n277156 , n261865 );
not ( n277158 , n261840 );
and ( n277159 , n277157 , n277158 );
not ( n277160 , n277157 );
and ( n277161 , n277160 , n261840 );
nor ( n277162 , n277159 , n277161 );
or ( n277163 , n277162 , n49959 );
nand ( n277164 , n277155 , n277163 );
buf ( n277165 , n277164 );
nand ( n277166 , n267311 , n243233 );
nand ( n277167 , n263788 , n267324 );
or ( n277168 , n277166 , n277167 );
not ( n277169 , n267311 );
not ( n277170 , n263788 );
or ( n277171 , n277169 , n277170 );
nor ( n277172 , n267324 , n240080 );
nand ( n277173 , n277171 , n277172 );
nand ( n277174 , n236798 , n28482 );
nand ( n277175 , n277168 , n277173 , n277174 );
buf ( n277176 , n277175 );
or ( n277177 , n25328 , n258787 );
or ( n277178 , n25335 , n264961 );
nand ( n277179 , n277177 , n277178 );
buf ( n277180 , n277179 );
nand ( n277181 , n264239 , n247444 );
not ( n277182 , n252749 );
nand ( n277183 , n277182 , n264251 );
or ( n277184 , n277181 , n277183 );
not ( n277185 , n264251 );
not ( n277186 , n264239 );
or ( n277187 , n277185 , n277186 );
nor ( n277188 , n277182 , n247212 );
nand ( n277189 , n277187 , n277188 );
nand ( n277190 , n256292 , n37250 );
nand ( n277191 , n277184 , n277189 , n277190 );
buf ( n277192 , n277191 );
not ( n277193 , n28407 );
not ( n277194 , n244606 );
or ( n277195 , n277193 , n277194 );
not ( n277196 , RI1754ae28_53);
or ( n277197 , n269544 , n277196 );
nand ( n277198 , n277195 , n277197 );
buf ( n277199 , n277198 );
not ( n277200 , RI19aa4cf0_2531);
or ( n277201 , n25328 , n277200 );
not ( n277202 , RI19a9b678_2602);
or ( n277203 , n25336 , n277202 );
nand ( n277204 , n277201 , n277203 );
buf ( n277205 , n277204 );
not ( n277206 , RI19a83b40_2768);
or ( n277207 , n25328 , n277206 );
or ( n277208 , n226822 , n269255 );
nand ( n277209 , n277207 , n277208 );
buf ( n277210 , n277209 );
nor ( n277211 , n275155 , n263369 );
nand ( n277212 , n267828 , n277211 );
nand ( n277213 , n267824 , n263369 );
not ( n277214 , n275155 );
not ( n277215 , n277214 );
not ( n277216 , n263355 );
not ( n277217 , n277216 );
and ( n277218 , n277215 , n277217 );
and ( n277219 , n236798 , n31750 );
nor ( n277220 , n277218 , n277219 );
nand ( n277221 , n277212 , n277213 , n277220 );
buf ( n277222 , n277221 );
not ( n277223 , n28578 );
not ( n277224 , n237714 );
or ( n277225 , n277223 , n277224 );
nand ( n277226 , n272020 , n258643 );
and ( n277227 , n277226 , n254539 );
not ( n277228 , n277226 );
and ( n277229 , n277228 , n258645 );
nor ( n277230 , n277227 , n277229 );
or ( n277231 , n277230 , n254882 );
nand ( n277232 , n277225 , n277231 );
buf ( n277233 , n277232 );
nand ( n277234 , n253976 , n254227 );
not ( n277235 , n253991 );
nand ( n277236 , n249368 , n277235 );
or ( n277237 , n277234 , n277236 );
not ( n277238 , n253976 );
not ( n277239 , n249368 );
or ( n277240 , n277238 , n277239 );
nor ( n277241 , n277235 , n234021 );
nand ( n277242 , n277240 , n277241 );
nand ( n277243 , n35431 , n37831 );
nand ( n277244 , n277237 , n277242 , n277243 );
buf ( n277245 , n277244 );
buf ( n277246 , n34501 );
buf ( n277247 , n29245 );
buf ( n277248 , n35990 );
not ( n277249 , n30612 );
not ( n277250 , n55760 );
or ( n277251 , n277249 , n277250 );
nand ( n277252 , n263986 , n263884 );
and ( n277253 , n277252 , n245268 );
not ( n277254 , n277252 );
and ( n277255 , n277254 , n245267 );
nor ( n277256 , n277253 , n277255 );
or ( n277257 , n277256 , n39763 );
nand ( n277258 , n277251 , n277257 );
buf ( n277259 , n277258 );
not ( n277260 , n240986 );
not ( n277261 , n277260 );
not ( n277262 , n54134 );
or ( n277263 , n277261 , n277262 );
or ( n277264 , n54134 , n277260 );
nand ( n277265 , n277263 , n277264 );
and ( n277266 , n277265 , n54192 );
not ( n277267 , n277265 );
and ( n277268 , n277267 , n231958 );
nor ( n277269 , n277266 , n277268 );
nand ( n277270 , n256079 , n236999 , n277269 );
not ( n277271 , n256073 );
not ( n277272 , n277271 );
not ( n277273 , n277269 );
or ( n277274 , n277272 , n277273 );
nor ( n277275 , n236999 , n235732 );
nand ( n277276 , n277274 , n277275 );
nand ( n277277 , n246460 , n37164 );
nand ( n277278 , n277270 , n277276 , n277277 );
buf ( n277279 , n277278 );
buf ( n277280 , n35010 );
nand ( n277281 , n266974 , n239934 );
not ( n277282 , n270529 );
nand ( n277283 , n263934 , n277282 );
or ( n277284 , n277281 , n277283 );
not ( n277285 , n277282 );
not ( n277286 , n266974 );
or ( n277287 , n277285 , n277286 );
nor ( n277288 , n263934 , n254740 );
nand ( n277289 , n277287 , n277288 );
nand ( n277290 , n241976 , n32708 );
nand ( n277291 , n277284 , n277289 , n277290 );
buf ( n277292 , n277291 );
not ( n277293 , n266189 );
nand ( n277294 , n277293 , n205649 );
nand ( n277295 , n259058 , n266201 );
or ( n277296 , n277294 , n277295 );
not ( n277297 , n266201 );
not ( n277298 , n277293 );
or ( n277299 , n277297 , n277298 );
nor ( n277300 , n259058 , n226955 );
nand ( n277301 , n277299 , n277300 );
nand ( n277302 , n238114 , n25341 );
nand ( n277303 , n277296 , n277301 , n277302 );
buf ( n277304 , n277303 );
nand ( n277305 , n276333 , n254528 );
not ( n277306 , n275917 );
nand ( n277307 , n276344 , n277306 );
or ( n277308 , n277305 , n277307 );
not ( n277309 , n276333 );
not ( n277310 , n276344 );
or ( n277311 , n277309 , n277310 );
nor ( n277312 , n277306 , n234440 );
nand ( n277313 , n277311 , n277312 );
nand ( n277314 , n50615 , n205053 );
nand ( n277315 , n277308 , n277313 , n277314 );
buf ( n277316 , n277315 );
not ( n277317 , n246335 );
nand ( n277318 , n277317 , n246452 );
or ( n277319 , n271012 , n277318 );
not ( n277320 , n271011 );
nand ( n277321 , n277320 , n251859 );
not ( n277322 , n277321 );
nand ( n277323 , n277322 , n277318 );
nand ( n277324 , n31577 , n208904 );
nand ( n277325 , n277319 , n277323 , n277324 );
buf ( n277326 , n277325 );
buf ( n277327 , n206043 );
buf ( n277328 , n208883 );
buf ( n277329 , n28499 );
not ( n277330 , n40837 );
not ( n277331 , n245943 );
or ( n277332 , n277330 , n277331 );
buf ( n277333 , n239902 );
not ( n277334 , n277333 );
not ( n277335 , n277334 );
not ( n277336 , n247569 );
or ( n277337 , n277335 , n277336 );
nand ( n277338 , n230199 , n277333 );
nand ( n277339 , n277337 , n277338 );
and ( n277340 , n277339 , n242696 );
not ( n277341 , n277339 );
and ( n277342 , n277341 , n247575 );
nor ( n277343 , n277340 , n277342 );
not ( n277344 , n277343 );
nand ( n277345 , n256046 , n277344 );
and ( n277346 , n277345 , n234191 );
not ( n277347 , n277345 );
and ( n277348 , n277347 , n234190 );
nor ( n277349 , n277346 , n277348 );
or ( n277350 , n277349 , n226003 );
nand ( n277351 , n277332 , n277350 );
buf ( n277352 , n277351 );
or ( n277353 , n25328 , n273585 );
not ( n277354 , RI19a8f648_2687);
or ( n277355 , n25335 , n277354 );
nand ( n277356 , n277353 , n277355 );
buf ( n277357 , n277356 );
not ( n277358 , n274853 );
not ( n277359 , n274652 );
nand ( n277360 , n277358 , n277359 );
or ( n277361 , n274631 , n277360 );
not ( n277362 , n277359 );
not ( n277363 , n274630 );
or ( n277364 , n277362 , n277363 );
nor ( n277365 , n277358 , n265700 );
nand ( n277366 , n277364 , n277365 );
nand ( n277367 , n234024 , n35675 );
nand ( n277368 , n277361 , n277366 , n277367 );
buf ( n277369 , n277368 );
buf ( n277370 , n36918 );
not ( n277371 , RI1754a888_65);
or ( n277372 , n249125 , n277371 );
not ( n277373 , RI19ac1d78_2315);
or ( n277374 , n25335 , n277373 );
nand ( n277375 , n277372 , n277374 );
buf ( n277376 , n277375 );
not ( n277377 , n276911 );
not ( n277378 , n252567 );
not ( n277379 , n248883 );
not ( n277380 , n277379 );
not ( n277381 , n237340 );
or ( n277382 , n277380 , n277381 );
nand ( n277383 , n237350 , n248883 );
nand ( n277384 , n277382 , n277383 );
not ( n277385 , n277384 );
or ( n277386 , n277378 , n277385 );
or ( n277387 , n277384 , n256280 );
nand ( n277388 , n277386 , n277387 );
not ( n277389 , n277388 );
nand ( n277390 , n276933 , n277377 , n277389 );
not ( n277391 , n276936 );
not ( n277392 , n277377 );
or ( n277393 , n277391 , n277392 );
nor ( n277394 , n277389 , n40465 );
nand ( n277395 , n277393 , n277394 );
nand ( n277396 , n254441 , n32892 );
nand ( n277397 , n277390 , n277395 , n277396 );
buf ( n277398 , n277397 );
not ( n277399 , n258864 );
nor ( n277400 , n258853 , n277399 );
not ( n277401 , n277400 );
not ( n277402 , n273681 );
or ( n277403 , n277401 , n277402 );
nand ( n277404 , n237714 , n29759 );
nand ( n277405 , n277403 , n277404 );
not ( n277406 , n277405 );
not ( n277407 , n273667 );
nand ( n277408 , n277407 , n277399 );
nor ( n277409 , n258864 , n42443 );
nand ( n277410 , n277409 , n258853 );
nand ( n277411 , n277406 , n277408 , n277410 );
buf ( n277412 , n277411 );
not ( n277413 , n38232 );
and ( n277414 , n54307 , n51336 );
not ( n277415 , n54307 );
and ( n277416 , n277415 , n51335 );
nor ( n277417 , n277414 , n277416 );
not ( n277418 , n277417 );
or ( n277419 , n277413 , n277418 );
not ( n277420 , n277417 );
nand ( n277421 , n38222 , n277420 );
nand ( n277422 , n277419 , n277421 );
not ( n277423 , n277422 );
not ( n277424 , n277423 );
not ( n277425 , n258439 );
not ( n277426 , n277425 );
or ( n277427 , n277424 , n277426 );
nor ( n277428 , n248002 , n235732 );
nand ( n277429 , n277427 , n277428 );
nor ( n277430 , n277422 , n235050 );
nand ( n277431 , n277425 , n277430 , n248002 );
nand ( n277432 , n237714 , n33597 );
nand ( n277433 , n277429 , n277431 , n277432 );
buf ( n277434 , n277433 );
nand ( n277435 , n269123 , n276807 , n272283 );
not ( n277436 , n269122 );
not ( n277437 , n277436 );
not ( n277438 , n272283 );
or ( n277439 , n277437 , n277438 );
nor ( n277440 , n276807 , n253213 );
nand ( n277441 , n277439 , n277440 );
nand ( n277442 , n245701 , n27694 );
nand ( n277443 , n277435 , n277441 , n277442 );
buf ( n277444 , n277443 );
not ( n277445 , n267488 );
nand ( n277446 , n277445 , n253397 );
not ( n277447 , n264664 );
buf ( n277448 , n249453 );
not ( n277449 , n277448 );
not ( n277450 , n38633 );
or ( n277451 , n277449 , n277450 );
or ( n277452 , n38633 , n277448 );
nand ( n277453 , n277451 , n277452 );
and ( n277454 , n277453 , n49191 );
not ( n277455 , n277453 );
and ( n277456 , n277455 , n49182 );
nor ( n277457 , n277454 , n277456 );
not ( n277458 , n277457 );
nand ( n277459 , n277447 , n277458 );
or ( n277460 , n277446 , n277459 );
nor ( n277461 , n277445 , n226003 );
nand ( n277462 , n277461 , n277459 );
nand ( n277463 , n247585 , n32448 );
nand ( n277464 , n277460 , n277462 , n277463 );
buf ( n277465 , n277464 );
nand ( n277466 , n270046 , n246177 );
nand ( n277467 , n250032 , n250051 );
or ( n277468 , n277466 , n277467 );
not ( n277469 , n270046 );
not ( n277470 , n250032 );
or ( n277471 , n277469 , n277470 );
nor ( n277472 , n250051 , n40465 );
nand ( n277473 , n277471 , n277472 );
nand ( n277474 , n247744 , n34154 );
nand ( n277475 , n277468 , n277473 , n277474 );
buf ( n277476 , n277475 );
nor ( n277477 , n264755 , n252070 );
not ( n277478 , n277477 );
not ( n277479 , n230828 );
not ( n277480 , n42149 );
or ( n277481 , n277479 , n277480 );
not ( n277482 , n230828 );
nand ( n277483 , n277482 , n42156 );
nand ( n277484 , n277481 , n277483 );
and ( n277485 , n277484 , n220201 );
not ( n277486 , n277484 );
and ( n277487 , n277486 , n220198 );
nor ( n277488 , n277485 , n277487 );
nand ( n277489 , n260815 , n277488 );
or ( n277490 , n277478 , n277489 );
nand ( n277491 , n264750 , n277489 );
nand ( n277492 , n245701 , n45301 );
nand ( n277493 , n277490 , n277491 , n277492 );
buf ( n277494 , n277493 );
buf ( n277495 , n31201 );
buf ( n277496 , n31657 );
not ( n277497 , RI19ab4380_2422);
or ( n277498 , n226819 , n277497 );
not ( n277499 , RI19aaa330_2494);
or ( n277500 , n226822 , n277499 );
nand ( n277501 , n277498 , n277500 );
buf ( n277502 , n277501 );
not ( n277503 , n275974 );
not ( n277504 , n275976 );
or ( n277505 , n277503 , n277504 );
nand ( n277506 , n277505 , n254636 );
nand ( n277507 , n276895 , n254635 , n275976 );
nand ( n277508 , n241976 , n36095 );
nand ( n277509 , n277506 , n277507 , n277508 );
buf ( n277510 , n277509 );
not ( n277511 , n254409 );
nor ( n277512 , n260716 , n268986 );
or ( n277513 , n277511 , n277512 );
nor ( n277514 , n254390 , n55146 );
nand ( n277515 , n277514 , n277512 );
nand ( n277516 , n35431 , n30350 );
nand ( n277517 , n277513 , n277515 , n277516 );
buf ( n277518 , n277517 );
not ( n277519 , n46474 );
not ( n277520 , n51606 );
or ( n277521 , n277519 , n277520 );
not ( n277522 , n46474 );
nand ( n277523 , n277522 , n51597 );
nand ( n277524 , n277521 , n277523 );
and ( n277525 , n277524 , n253197 );
not ( n277526 , n277524 );
and ( n277527 , n277526 , n253189 );
nor ( n277528 , n277525 , n277527 );
not ( n277529 , n277528 );
nand ( n277530 , n274777 , n277529 );
or ( n277531 , n274766 , n277530 );
nor ( n277532 , n274765 , n40465 );
nand ( n277533 , n277532 , n277530 );
nand ( n277534 , n39766 , n204960 );
nand ( n277535 , n277531 , n277533 , n277534 );
buf ( n277536 , n277535 );
not ( n277537 , n250576 );
not ( n277538 , n253780 );
not ( n277539 , n277538 );
and ( n277540 , n277537 , n277539 );
and ( n277541 , n250576 , n277538 );
nor ( n277542 , n277540 , n277541 );
and ( n277543 , n277542 , n252037 );
not ( n277544 , n277542 );
and ( n277545 , n277544 , n252052 );
nor ( n277546 , n277543 , n277545 );
nor ( n277547 , n262571 , n277546 );
nand ( n277548 , n256512 , n277547 );
not ( n277549 , n262574 );
not ( n277550 , n256492 );
or ( n277551 , n277549 , n277550 );
not ( n277552 , n277546 );
nor ( n277553 , n277552 , n40465 );
nand ( n277554 , n277551 , n277553 );
nand ( n277555 , n39767 , n38408 );
nand ( n277556 , n277548 , n277554 , n277555 );
buf ( n277557 , n277556 );
nand ( n277558 , n273127 , n254035 );
or ( n277559 , n257462 , n277558 );
not ( n277560 , n254035 );
not ( n277561 , n254023 );
or ( n277562 , n277560 , n277561 );
nor ( n277563 , n273127 , n234440 );
nand ( n277564 , n277562 , n277563 );
nand ( n277565 , n244789 , n28612 );
nand ( n277566 , n277559 , n277564 , n277565 );
buf ( n277567 , n277566 );
not ( n277568 , n254827 );
nand ( n277569 , n254876 , n277568 );
not ( n277570 , n274494 );
or ( n277571 , n277569 , n277570 );
nor ( n277572 , n274476 , n234440 );
nand ( n277573 , n277569 , n277572 );
nand ( n277574 , n247585 , n27725 );
nand ( n277575 , n277571 , n277573 , n277574 );
buf ( n277576 , n277575 );
not ( n277577 , RI19aabcf8_2483);
or ( n277578 , n25328 , n277577 );
not ( n277579 , RI19aa1d20_2554);
or ( n277580 , n25335 , n277579 );
nand ( n277581 , n277578 , n277580 );
buf ( n277582 , n277581 );
not ( n277583 , n259756 );
not ( n277584 , n247625 );
not ( n277585 , n48233 );
or ( n277586 , n277584 , n277585 );
not ( n277587 , n247625 );
nand ( n277588 , n277587 , n48232 );
nand ( n277589 , n277586 , n277588 );
not ( n277590 , n277589 );
or ( n277591 , n277583 , n277590 );
or ( n277592 , n277589 , n253578 );
nand ( n277593 , n277591 , n277592 );
not ( n277594 , n277593 );
nand ( n277595 , n277594 , n272515 );
nand ( n277596 , n268206 , n241459 );
or ( n277597 , n277595 , n277596 );
nand ( n277598 , n277595 , n268210 );
nand ( n277599 , n49054 , n205100 );
nand ( n277600 , n277597 , n277598 , n277599 );
buf ( n277601 , n277600 );
buf ( n277602 , n25806 );
buf ( n277603 , n28836 );
nor ( n277604 , n252449 , n252462 );
not ( n277605 , n238692 );
not ( n277606 , n247991 );
or ( n277607 , n277605 , n277606 );
or ( n277608 , n247991 , n238692 );
nand ( n277609 , n277607 , n277608 );
and ( n277610 , n277609 , n261859 );
not ( n277611 , n277609 );
and ( n277612 , n277611 , n261862 );
nor ( n277613 , n277610 , n277612 );
nand ( n277614 , n277613 , n259783 );
or ( n277615 , n277604 , n277614 );
nor ( n277616 , n277613 , n244399 );
nand ( n277617 , n277616 , n277604 );
nand ( n277618 , n49054 , n225252 );
nand ( n277619 , n277615 , n277617 , n277618 );
buf ( n277620 , n277619 );
buf ( n277621 , n49741 );
buf ( n277622 , n29066 );
not ( n277623 , RI19ac3b00_2301);
or ( n277624 , n25328 , n277623 );
or ( n277625 , n25335 , n272172 );
nand ( n277626 , n277624 , n277625 );
buf ( n277627 , n277626 );
buf ( n277628 , n204851 );
buf ( n277629 , n26065 );
buf ( n277630 , n36064 );
buf ( n277631 , n36272 );
nand ( n277632 , n271202 , n261996 );
or ( n277633 , n262003 , n277632 );
not ( n277634 , n271202 );
not ( n277635 , n261972 );
or ( n277636 , n277634 , n277635 );
nor ( n277637 , n261996 , n249531 );
nand ( n277638 , n277636 , n277637 );
nand ( n277639 , n241378 , n26401 );
nand ( n277640 , n277633 , n277638 , n277639 );
buf ( n277641 , n277640 );
buf ( n277642 , n25718 );
or ( n277643 , n233507 , n276817 );
not ( n277644 , RI19a89018_2731);
or ( n277645 , n25335 , n277644 );
nand ( n277646 , n277643 , n277645 );
buf ( n277647 , n277646 );
buf ( n277648 , n41436 );
buf ( n277649 , n31412 );
or ( n277650 , n233507 , n265260 );
or ( n277651 , n25336 , n271705 );
nand ( n277652 , n277650 , n277651 );
buf ( n277653 , n277652 );
nand ( n277654 , n259280 , n255152 );
not ( n277655 , n47224 );
not ( n277656 , n277655 );
not ( n277657 , n254076 );
or ( n277658 , n277656 , n277657 );
nand ( n277659 , n254077 , n47224 );
nand ( n277660 , n277658 , n277659 );
and ( n277661 , n277660 , n237639 );
not ( n277662 , n277660 );
and ( n277663 , n277662 , n254080 );
nor ( n277664 , n277661 , n277663 );
nand ( n277665 , n277664 , n276222 );
or ( n277666 , n277654 , n277665 );
not ( n277667 , n277664 );
not ( n277668 , n259280 );
or ( n277669 , n277667 , n277668 );
nand ( n277670 , n277669 , n276227 );
nand ( n277671 , n31576 , n44121 );
nand ( n277672 , n277666 , n277670 , n277671 );
buf ( n277673 , n277672 );
not ( n277674 , n276835 );
or ( n277675 , n255912 , n277674 );
nor ( n277676 , n255911 , n242391 );
nor ( n277677 , n255934 , n276835 );
nand ( n277678 , n277676 , n277677 );
not ( n277679 , n255935 );
nand ( n277680 , n276835 , n243438 );
not ( n277681 , n277680 );
and ( n277682 , n277679 , n277681 );
and ( n277683 , n46083 , n204867 );
nor ( n277684 , n277682 , n277683 );
nand ( n277685 , n277675 , n277678 , n277684 );
buf ( n277686 , n277685 );
not ( n277687 , n27891 );
not ( n277688 , n251465 );
or ( n277689 , n277687 , n277688 );
nand ( n277690 , n240059 , n249212 );
and ( n277691 , n277690 , n240077 );
not ( n277692 , n277690 );
not ( n277693 , n240077 );
and ( n277694 , n277692 , n277693 );
nor ( n277695 , n277691 , n277694 );
or ( n277696 , n277695 , n256214 );
nand ( n277697 , n277689 , n277696 );
buf ( n277698 , n277697 );
nand ( n277699 , n273996 , n260774 , n257833 );
not ( n277700 , n263909 );
not ( n277701 , n260774 );
or ( n277702 , n277700 , n277701 );
nor ( n277703 , n257833 , n31572 );
nand ( n277704 , n277702 , n277703 );
nand ( n277705 , n234448 , n37877 );
nand ( n277706 , n277699 , n277704 , n277705 );
buf ( n277707 , n277706 );
nand ( n277708 , n272820 , n275852 );
or ( n277709 , n272797 , n277708 );
not ( n277710 , n272820 );
not ( n277711 , n272796 );
or ( n277712 , n277710 , n277711 );
nor ( n277713 , n275852 , n241065 );
nand ( n277714 , n277712 , n277713 );
nand ( n277715 , n238114 , n29209 );
nand ( n277716 , n277709 , n277714 , n277715 );
buf ( n277717 , n277716 );
nand ( n277718 , n270952 , n25321 , n266635 );
and ( n277719 , n277718 , n266633 );
nor ( n277720 , n251562 , RI1754c610_2);
not ( n277721 , n277720 );
nor ( n277722 , n277719 , n277721 );
buf ( n277723 , n277722 );
not ( n277724 , n263671 );
nand ( n277725 , n277724 , n241704 );
nand ( n277726 , n275537 , n275547 );
or ( n277727 , n277725 , n277726 );
not ( n277728 , n275547 );
not ( n277729 , n277724 );
or ( n277730 , n277728 , n277729 );
nor ( n277731 , n275537 , n250909 );
nand ( n277732 , n277730 , n277731 );
nand ( n277733 , n31577 , n26034 );
nand ( n277734 , n277727 , n277732 , n277733 );
buf ( n277735 , n277734 );
nand ( n277736 , n276866 , n222532 );
not ( n277737 , n276762 );
nand ( n277738 , n276886 , n277737 );
or ( n277739 , n277736 , n277738 );
not ( n277740 , n276886 );
not ( n277741 , n276866 );
or ( n277742 , n277740 , n277741 );
nor ( n277743 , n277737 , n256481 );
nand ( n277744 , n277742 , n277743 );
nand ( n277745 , n245414 , n240166 );
nand ( n277746 , n277739 , n277744 , n277745 );
buf ( n277747 , n277746 );
not ( n277748 , n272550 );
nand ( n277749 , n277748 , n272561 );
or ( n277750 , n262880 , n277749 );
not ( n277751 , n277748 );
not ( n277752 , n262879 );
or ( n277753 , n277751 , n277752 );
nor ( n277754 , n272561 , n219702 );
nand ( n277755 , n277753 , n277754 );
nand ( n277756 , n35431 , n223454 );
nand ( n277757 , n277750 , n277755 , n277756 );
buf ( n277758 , n277757 );
not ( n277759 , RI19ac9b90_2257);
or ( n277760 , n226819 , n277759 );
not ( n277761 , RI19ac0860_2327);
or ( n277762 , n25335 , n277761 );
nand ( n277763 , n277760 , n277762 );
buf ( n277764 , n277763 );
nand ( n277765 , n265563 , n275385 );
or ( n277766 , n277765 , n265577 );
not ( n277767 , n265576 );
not ( n277768 , n265563 );
or ( n277769 , n277767 , n277768 );
nor ( n277770 , n275385 , n234021 );
nand ( n277771 , n277769 , n277770 );
nand ( n277772 , n246217 , n28222 );
nand ( n277773 , n277766 , n277771 , n277772 );
buf ( n277774 , n277773 );
not ( n277775 , n277269 );
nand ( n277776 , n236999 , n277775 );
or ( n277777 , n236826 , n277776 );
nor ( n277778 , n236825 , n244216 );
nand ( n277779 , n277778 , n277776 );
nand ( n277780 , n41944 , n25806 );
nand ( n277781 , n277777 , n277779 , n277780 );
buf ( n277782 , n277781 );
or ( n277783 , n25328 , n276517 );
or ( n277784 , n226822 , n248829 );
nand ( n277785 , n277783 , n277784 );
buf ( n277786 , n277785 );
nand ( n277787 , n264324 , n249009 );
nand ( n277788 , n275045 , n264336 );
or ( n277789 , n277787 , n277788 );
not ( n277790 , n264336 );
not ( n277791 , n264324 );
or ( n277792 , n277790 , n277791 );
nor ( n277793 , n275045 , n55104 );
nand ( n277794 , n277792 , n277793 );
nand ( n277795 , n31577 , n33641 );
nand ( n277796 , n277789 , n277794 , n277795 );
buf ( n277797 , n277796 );
not ( n277798 , n204419 );
not ( n277799 , n234823 );
or ( n277800 , n277798 , n277799 );
not ( n277801 , n273166 );
nand ( n277802 , n277801 , n35815 );
and ( n277803 , n277802 , n269201 );
not ( n277804 , n277802 );
and ( n277805 , n277804 , n36734 );
nor ( n277806 , n277803 , n277805 );
or ( n277807 , n277806 , n238223 );
nand ( n277808 , n277800 , n277807 );
buf ( n277809 , n277808 );
not ( n277810 , n27881 );
not ( n277811 , n204518 );
or ( n277812 , n277810 , n277811 );
nand ( n277813 , n277812 , n204515 );
and ( n277814 , n27883 , n277813 );
buf ( n277815 , n277814 );
not ( n277816 , n26332 );
not ( n277817 , n245943 );
or ( n277818 , n277816 , n277817 );
not ( n277819 , n264615 );
not ( n277820 , n264629 );
nand ( n277821 , n277819 , n277820 );
and ( n277822 , n277821 , n270883 );
not ( n277823 , n277821 );
and ( n277824 , n277823 , n266426 );
nor ( n277825 , n277822 , n277824 );
or ( n277826 , n277825 , n244217 );
nand ( n277827 , n277818 , n277826 );
buf ( n277828 , n277827 );
not ( n277829 , n43712 );
not ( n277830 , n242270 );
or ( n277831 , n277829 , n277830 );
not ( n277832 , n43712 );
nand ( n277833 , n277832 , n252503 );
nand ( n277834 , n277831 , n277833 );
and ( n277835 , n277834 , n252553 );
not ( n277836 , n277834 );
and ( n277837 , n277836 , n252562 );
nor ( n277838 , n277835 , n277837 );
not ( n277839 , n277838 );
not ( n277840 , n254356 );
nand ( n277841 , n277839 , n277840 );
or ( n277842 , n277841 , n254271 );
not ( n277843 , n267561 );
nand ( n277844 , n277843 , n277841 );
nand ( n277845 , n246460 , n39635 );
nand ( n277846 , n277842 , n277844 , n277845 );
buf ( n277847 , n277846 );
not ( n277848 , n222471 );
not ( n277849 , n244073 );
or ( n277850 , n277848 , n277849 );
nand ( n277851 , n247405 , n275706 );
and ( n277852 , n277851 , n271619 );
not ( n277853 , n277851 );
not ( n277854 , n271619 );
and ( n277855 , n277853 , n277854 );
nor ( n277856 , n277852 , n277855 );
or ( n277857 , n277856 , n235052 );
nand ( n277858 , n277850 , n277857 );
buf ( n277859 , n277858 );
or ( n277860 , n25328 , n263874 );
or ( n277861 , n25336 , n270332 );
nand ( n277862 , n277860 , n277861 );
buf ( n277863 , n277862 );
buf ( n277864 , n257918 );
not ( n277865 , n277864 );
not ( n277866 , n250691 );
or ( n277867 , n277865 , n277866 );
or ( n277868 , n250691 , n277864 );
nand ( n277869 , n277867 , n277868 );
and ( n277870 , n277869 , n262217 );
not ( n277871 , n277869 );
and ( n277872 , n277871 , n262220 );
nor ( n277873 , n277870 , n277872 );
not ( n277874 , n277873 );
nand ( n277875 , n270733 , n277874 );
or ( n277876 , n242687 , n277875 );
not ( n277877 , n270733 );
not ( n277878 , n242686 );
or ( n277879 , n277877 , n277878 );
nor ( n277880 , n277874 , n40465 );
nand ( n277881 , n277879 , n277880 );
nand ( n277882 , n255116 , n25796 );
nand ( n277883 , n277876 , n277881 , n277882 );
buf ( n277884 , n277883 );
nand ( n277885 , n262007 , n271203 , n262339 );
nand ( n277886 , n262339 , n262005 );
nand ( n277887 , n277886 , n271202 , n205649 );
nand ( n277888 , n55760 , n26459 );
nand ( n277889 , n277885 , n277887 , n277888 );
buf ( n277890 , n277889 );
nor ( n277891 , n259580 , n39763 );
not ( n277892 , n27878 );
not ( n277893 , n242116 );
not ( n277894 , n277893 );
not ( n277895 , n204544 );
or ( n277896 , n277894 , n277895 );
nand ( n277897 , n204553 , n242116 );
nand ( n277898 , n277896 , n277897 );
not ( n277899 , n277898 );
or ( n277900 , n277892 , n277899 );
or ( n277901 , n277898 , n27878 );
nand ( n277902 , n277900 , n277901 );
not ( n277903 , n277902 );
nor ( n277904 , n265683 , n277903 );
nand ( n277905 , n277891 , n277904 );
not ( n277906 , n277902 );
not ( n277907 , n259580 );
not ( n277908 , n277907 );
or ( n277909 , n277906 , n277908 );
nor ( n277910 , n259597 , n226955 );
nand ( n277911 , n277909 , n277910 );
nand ( n277912 , n31577 , n25836 );
nand ( n277913 , n277905 , n277911 , n277912 );
buf ( n277914 , n277913 );
not ( n277915 , RI19a96e48_2634);
or ( n277916 , n25328 , n277915 );
not ( n277917 , RI19a8cb28_2706);
or ( n277918 , n226822 , n277917 );
nand ( n277919 , n277916 , n277918 );
buf ( n277920 , n277919 );
not ( n277921 , RI1754bbc0_24);
or ( n277922 , n255977 , n277921 );
nand ( n277923 , n258185 , n34282 );
nand ( n277924 , n277922 , n277923 );
buf ( n277925 , n277924 );
not ( n277926 , n29791 );
not ( n277927 , n245943 );
or ( n277928 , n277926 , n277927 );
nand ( n277929 , n275368 , n259533 );
not ( n277930 , n277929 );
not ( n277931 , n259545 );
and ( n277932 , n277930 , n277931 );
and ( n277933 , n277929 , n259545 );
nor ( n277934 , n277932 , n277933 );
or ( n277935 , n277934 , n240080 );
nand ( n277936 , n277928 , n277935 );
buf ( n277937 , n277936 );
not ( n277938 , n268574 );
not ( n277939 , n264079 );
or ( n277940 , n277938 , n277939 );
nor ( n277941 , n267448 , n235895 );
nand ( n277942 , n277940 , n277941 );
nand ( n277943 , n264079 , n272781 , n267448 );
nand ( n277944 , n35431 , n29492 );
nand ( n277945 , n277942 , n277943 , n277944 );
buf ( n277946 , n277945 );
not ( n277947 , RI19abf690_2337);
or ( n277948 , n226819 , n277947 );
or ( n277949 , n25335 , n264400 );
nand ( n277950 , n277948 , n277949 );
buf ( n277951 , n277950 );
not ( n277952 , n250526 );
not ( n277953 , n227174 );
or ( n277954 , n277952 , n277953 );
not ( n277955 , n250526 );
nand ( n277956 , n277955 , n49420 );
nand ( n277957 , n277954 , n277956 );
and ( n277958 , n277957 , n49618 );
not ( n277959 , n277957 );
and ( n277960 , n277959 , n49627 );
nor ( n277961 , n277958 , n277960 );
nor ( n277962 , n277961 , n37725 );
not ( n277963 , n253564 );
nand ( n277964 , n277963 , n253591 );
nand ( n277965 , n277962 , n277964 );
not ( n277966 , n277961 );
nor ( n277967 , n277966 , n253590 );
nand ( n277968 , n277967 , n265001 );
nand ( n277969 , n238114 , n29725 );
nand ( n277970 , n277965 , n277968 , n277969 );
buf ( n277971 , n277970 );
not ( n277972 , n35524 );
not ( n277973 , n258213 );
or ( n277974 , n277972 , n277973 );
nand ( n277975 , n251461 , n251453 );
and ( n277976 , n277975 , n273436 );
not ( n277977 , n277975 );
and ( n277978 , n277977 , n273435 );
nor ( n277979 , n277976 , n277978 );
or ( n277980 , n277979 , n255707 );
nand ( n277981 , n277974 , n277980 );
buf ( n277982 , n277981 );
not ( n277983 , n253199 );
nor ( n277984 , n269920 , n277983 );
nand ( n277985 , n253214 , n277984 );
not ( n277986 , n253199 );
not ( n277987 , n253138 );
not ( n277988 , n277987 );
or ( n277989 , n277986 , n277988 );
nor ( n277990 , n269919 , n237384 );
nand ( n277991 , n277989 , n277990 );
nand ( n277992 , n234453 , n29841 );
nand ( n277993 , n277985 , n277991 , n277992 );
buf ( n277994 , n277993 );
not ( n277995 , n31813 );
not ( n277996 , n258213 );
or ( n277997 , n277995 , n277996 );
nand ( n277998 , n258396 , n258406 );
not ( n277999 , n266957 );
and ( n278000 , n277998 , n277999 );
not ( n278001 , n277998 );
and ( n278002 , n278001 , n266957 );
nor ( n278003 , n278000 , n278002 );
or ( n278004 , n278003 , n255707 );
nand ( n278005 , n277997 , n278004 );
buf ( n278006 , n278005 );
not ( n278007 , n267044 );
not ( n278008 , n270476 );
or ( n278009 , n278007 , n278008 );
nor ( n278010 , n269022 , n236795 );
nand ( n278011 , n278009 , n278010 );
nand ( n278012 , n267046 , n269022 , n270476 );
nand ( n278013 , n51381 , n30715 );
nand ( n278014 , n278011 , n278012 , n278013 );
buf ( n278015 , n278014 );
not ( n278016 , n255754 );
not ( n278017 , n249541 );
or ( n278018 , n278016 , n278017 );
or ( n278019 , n249541 , n255754 );
nand ( n278020 , n278018 , n278019 );
and ( n278021 , n278020 , n249549 );
not ( n278022 , n278020 );
and ( n278023 , n278022 , n249546 );
nor ( n278024 , n278021 , n278023 );
nand ( n278025 , n278024 , n272711 );
not ( n278026 , n37363 );
not ( n278027 , n278026 );
not ( n278028 , n257724 );
or ( n278029 , n278027 , n278028 );
or ( n278030 , n258715 , n278026 );
nand ( n278031 , n278029 , n278030 );
and ( n278032 , n278031 , n257732 );
not ( n278033 , n278031 );
and ( n278034 , n278033 , n257729 );
nor ( n278035 , n278032 , n278034 );
not ( n278036 , n278035 );
nand ( n278037 , n253539 , n278036 );
or ( n278038 , n278025 , n278037 );
nor ( n278039 , n278024 , n40465 );
nand ( n278040 , n278039 , n278037 );
nand ( n278041 , n249622 , n28219 );
nand ( n278042 , n278038 , n278040 , n278041 );
buf ( n278043 , n278042 );
buf ( n278044 , RI19ad0e08_2205);
and ( n278045 , n25326 , n278044 );
buf ( n278046 , n278045 );
not ( n278047 , n269476 );
not ( n278048 , n254847 );
not ( n278049 , n55345 );
or ( n278050 , n278048 , n278049 );
not ( n278051 , n254847 );
nand ( n278052 , n278051 , n33708 );
nand ( n278053 , n278050 , n278052 );
and ( n278054 , n278053 , n55511 );
not ( n278055 , n278053 );
and ( n278056 , n278055 , n233265 );
nor ( n278057 , n278054 , n278056 );
nand ( n278058 , n278057 , n266088 );
or ( n278059 , n278047 , n278058 );
not ( n278060 , n269471 );
not ( n278061 , n278057 );
or ( n278062 , n278060 , n278061 );
nor ( n278063 , n266088 , n240080 );
nand ( n278064 , n278062 , n278063 );
nand ( n278065 , n41945 , n25619 );
nand ( n278066 , n278059 , n278064 , n278065 );
buf ( n278067 , n278066 );
not ( n278068 , n270917 );
nand ( n278069 , n274070 , n268775 );
or ( n278070 , n278068 , n278069 );
not ( n278071 , n274070 );
not ( n278072 , n270912 );
or ( n278073 , n278071 , n278072 );
nor ( n278074 , n268775 , n219702 );
nand ( n278075 , n278073 , n278074 );
nand ( n278076 , n263598 , n38640 );
nand ( n278077 , n278070 , n278075 , n278076 );
buf ( n278078 , n278077 );
nand ( n278079 , n265189 , n252873 );
not ( n278080 , n246984 );
not ( n278081 , n278080 );
not ( n278082 , n242148 );
or ( n278083 , n278081 , n278082 );
not ( n278084 , n278080 );
nand ( n278085 , n278084 , n242155 );
nand ( n278086 , n278083 , n278085 );
and ( n278087 , n278086 , n242206 );
not ( n278088 , n278086 );
and ( n278089 , n278088 , n242202 );
nor ( n278090 , n278087 , n278089 );
not ( n278091 , n278090 );
not ( n278092 , n246425 );
not ( n278093 , n256742 );
or ( n278094 , n278092 , n278093 );
not ( n278095 , n246425 );
nand ( n278096 , n278095 , n256738 );
nand ( n278097 , n278094 , n278096 );
and ( n278098 , n278097 , n256748 );
not ( n278099 , n278097 );
and ( n278100 , n278099 , n261630 );
nor ( n278101 , n278098 , n278100 );
nand ( n278102 , n278091 , n278101 );
or ( n278103 , n278079 , n278102 );
not ( n278104 , n278101 );
not ( n278105 , n265189 );
or ( n278106 , n278104 , n278105 );
nor ( n278107 , n278091 , n234021 );
nand ( n278108 , n278106 , n278107 );
nand ( n278109 , n31576 , n25447 );
nand ( n278110 , n278103 , n278108 , n278109 );
buf ( n278111 , n278110 );
not ( n278112 , n270234 );
nand ( n278113 , n278112 , n50945 );
not ( n278114 , n47429 );
not ( n278115 , n263900 );
or ( n278116 , n278114 , n278115 );
not ( n278117 , n47429 );
nand ( n278118 , n278117 , n250896 );
nand ( n278119 , n278116 , n278118 );
and ( n278120 , n278119 , n250903 );
not ( n278121 , n278119 );
and ( n278122 , n278121 , n250906 );
nor ( n278123 , n278120 , n278122 );
not ( n278124 , n278123 );
nand ( n278125 , n270245 , n278124 );
or ( n278126 , n278113 , n278125 );
not ( n278127 , n270245 );
not ( n278128 , n278112 );
or ( n278129 , n278127 , n278128 );
nor ( n278130 , n278124 , n55146 );
nand ( n278131 , n278129 , n278130 );
nand ( n278132 , n238114 , n32713 );
nand ( n278133 , n278126 , n278131 , n278132 );
buf ( n278134 , n278133 );
not ( n278135 , n251362 );
not ( n278136 , n276394 );
nand ( n278137 , n278136 , n259645 );
or ( n278138 , n278135 , n278137 );
not ( n278139 , n259645 );
not ( n278140 , n251335 );
or ( n278141 , n278139 , n278140 );
nor ( n278142 , n278136 , n253904 );
nand ( n278143 , n278141 , n278142 );
nand ( n278144 , n234024 , n31019 );
nand ( n278145 , n278138 , n278143 , n278144 );
buf ( n278146 , n278145 );
not ( n278147 , n261049 );
nand ( n278148 , n278147 , n261062 );
or ( n278149 , n269677 , n278148 );
nor ( n278150 , n269676 , n234021 );
nand ( n278151 , n278150 , n278148 );
nand ( n278152 , n35431 , n32625 );
nand ( n278153 , n278149 , n278151 , n278152 );
buf ( n278154 , n278153 );
not ( n278155 , n259174 );
not ( n278156 , n278155 );
not ( n278157 , n256209 );
or ( n278158 , n278156 , n278157 );
nor ( n278159 , n259158 , n247276 );
nand ( n278160 , n278158 , n278159 );
nor ( n278161 , n259174 , n39763 );
nand ( n278162 , n278161 , n256209 , n259158 );
nand ( n278163 , n234453 , n32746 );
nand ( n278164 , n278160 , n278162 , n278163 );
buf ( n278165 , n278164 );
nand ( n278166 , n257734 , n257747 );
not ( n278167 , n237992 );
not ( n278168 , n278167 );
not ( n278169 , n226319 );
or ( n278170 , n278168 , n278169 );
nand ( n278171 , n257110 , n237992 );
nand ( n278172 , n278170 , n278171 );
and ( n278173 , n278172 , n257116 );
not ( n278174 , n278172 );
and ( n278175 , n278174 , n258557 );
nor ( n278176 , n278173 , n278175 );
nand ( n278177 , n278176 , n257527 );
or ( n278178 , n278166 , n278177 );
not ( n278179 , n278176 );
not ( n278180 , n257734 );
or ( n278181 , n278179 , n278180 );
nor ( n278182 , n257747 , n244399 );
nand ( n278183 , n278181 , n278182 );
nand ( n278184 , n49054 , n31310 );
nand ( n278185 , n278178 , n278183 , n278184 );
buf ( n278186 , n278185 );
buf ( n278187 , n206401 );
not ( n278188 , n255563 );
not ( n278189 , n238628 );
or ( n278190 , n278188 , n278189 );
not ( n278191 , n255563 );
nand ( n278192 , n278191 , n238620 );
nand ( n278193 , n278190 , n278192 );
and ( n278194 , n278193 , n257185 );
not ( n278195 , n278193 );
and ( n278196 , n278195 , n257188 );
nor ( n278197 , n278194 , n278196 );
not ( n278198 , n248231 );
not ( n278199 , n240312 );
or ( n278200 , n278198 , n278199 );
not ( n278201 , n248231 );
nand ( n278202 , n278201 , n240316 );
nand ( n278203 , n278200 , n278202 );
and ( n278204 , n278203 , n240508 );
not ( n278205 , n278203 );
and ( n278206 , n278205 , n240505 );
nor ( n278207 , n278204 , n278206 );
nand ( n278208 , n268103 , n278197 , n278207 );
not ( n278209 , n268099 );
not ( n278210 , n278197 );
or ( n278211 , n278209 , n278210 );
nor ( n278212 , n278207 , n250909 );
nand ( n278213 , n278211 , n278212 );
nand ( n278214 , n35431 , n207997 );
nand ( n278215 , n278208 , n278213 , n278214 );
buf ( n278216 , n278215 );
nand ( n278217 , n276806 , n269134 );
not ( n278218 , n269147 );
or ( n278219 , n278217 , n278218 );
nand ( n278220 , n278217 , n272287 );
nand ( n278221 , n244789 , n215681 );
nand ( n278222 , n278219 , n278220 , n278221 );
buf ( n278223 , n278222 );
not ( n278224 , n275782 );
not ( n278225 , n275665 );
nand ( n278226 , n278225 , n275675 );
or ( n278227 , n278224 , n278226 );
not ( n278228 , n278225 );
not ( n278229 , n275781 );
not ( n278230 , n278229 );
or ( n278231 , n278228 , n278230 );
nor ( n278232 , n275675 , n37725 );
nand ( n278233 , n278231 , n278232 );
nand ( n278234 , n31577 , n47282 );
nand ( n278235 , n278227 , n278233 , n278234 );
buf ( n278236 , n278235 );
not ( n278237 , n255848 );
not ( n278238 , n278237 );
not ( n278239 , n229300 );
or ( n278240 , n278238 , n278239 );
not ( n278241 , n278237 );
nand ( n278242 , n278241 , n51549 );
nand ( n278243 , n278240 , n278242 );
and ( n278244 , n278243 , n51598 );
not ( n278245 , n278243 );
and ( n278246 , n278245 , n51607 );
nor ( n278247 , n278244 , n278246 );
nor ( n278248 , n278247 , n271667 );
nand ( n278249 , n257715 , n278248 );
not ( n278250 , n271666 );
not ( n278251 , n257696 );
not ( n278252 , n278251 );
or ( n278253 , n278250 , n278252 );
not ( n278254 , n278247 );
nor ( n278255 , n278254 , n252679 );
nand ( n278256 , n278253 , n278255 );
nand ( n278257 , n238638 , n32667 );
nand ( n278258 , n278249 , n278256 , n278257 );
buf ( n278259 , n278258 );
buf ( n278260 , n29236 );
nand ( n278261 , n275434 , n244515 );
buf ( n278262 , n35606 );
not ( n278263 , n278262 );
not ( n278264 , n236886 );
or ( n278265 , n278263 , n278264 );
or ( n278266 , n236886 , n278262 );
nand ( n278267 , n278265 , n278266 );
not ( n278268 , n278267 );
not ( n278269 , n258860 );
and ( n278270 , n278268 , n278269 );
and ( n278271 , n278267 , n258860 );
nor ( n278272 , n278270 , n278271 );
nand ( n278273 , n278272 , n273303 );
or ( n278274 , n278261 , n278273 );
not ( n278275 , n275434 );
not ( n278276 , n278272 );
or ( n278277 , n278275 , n278276 );
nor ( n278278 , n273303 , n244399 );
nand ( n278279 , n278277 , n278278 );
nand ( n278280 , n31577 , n33624 );
nand ( n278281 , n278274 , n278279 , n278280 );
buf ( n278282 , n278281 );
nand ( n278283 , n260615 , n273955 , n274907 );
not ( n278284 , n260609 );
nand ( n278285 , n278284 , n274907 );
nand ( n278286 , n278285 , n273956 , n259619 );
nand ( n278287 , n37728 , n25735 );
nand ( n278288 , n278283 , n278286 , n278287 );
buf ( n278289 , n278288 );
not ( n278290 , n205284 );
not ( n278291 , n245943 );
or ( n278292 , n278290 , n278291 );
not ( n278293 , n253878 );
nand ( n278294 , n278293 , n261239 );
and ( n278295 , n278294 , n264979 );
not ( n278296 , n278294 );
and ( n278297 , n278296 , n264978 );
nor ( n278298 , n278295 , n278297 );
or ( n278299 , n278298 , n258179 );
nand ( n278300 , n278292 , n278299 );
buf ( n278301 , n278300 );
nand ( n278302 , n47327 , n245802 );
not ( n278303 , n274187 );
or ( n278304 , n278302 , n278303 );
not ( n278305 , n274181 );
not ( n278306 , n47327 );
or ( n278307 , n278305 , n278306 );
nor ( n278308 , n245802 , n50944 );
nand ( n278309 , n278307 , n278308 );
nand ( n278310 , n247585 , n34066 );
nand ( n278311 , n278304 , n278309 , n278310 );
buf ( n278312 , n278311 );
buf ( n278313 , n225252 );
buf ( n278314 , n221006 );
buf ( n278315 , n25323 );
not ( n278316 , n258237 );
not ( n278317 , n251706 );
nand ( n278318 , n278316 , n278317 );
or ( n278319 , n251635 , n278318 );
not ( n278320 , n278317 );
not ( n278321 , n251634 );
or ( n278322 , n278320 , n278321 );
nor ( n278323 , n278316 , n251361 );
nand ( n278324 , n278322 , n278323 );
nand ( n278325 , n31577 , n204922 );
nand ( n278326 , n278319 , n278324 , n278325 );
buf ( n278327 , n278326 );
not ( n278328 , n29263 );
not ( n278329 , n31577 );
or ( n278330 , n278328 , n278329 );
not ( n278331 , n266389 );
nand ( n278332 , n278331 , n266378 );
and ( n278333 , n278332 , n277025 );
not ( n278334 , n278332 );
and ( n278335 , n278334 , n277105 );
nor ( n278336 , n278333 , n278335 );
or ( n278337 , n278336 , n254882 );
nand ( n278338 , n278330 , n278337 );
buf ( n278339 , n278338 );
nand ( n278340 , n265904 , n236509 );
nand ( n278341 , n274358 , n260375 );
or ( n278342 , n278340 , n278341 );
nand ( n278343 , n278340 , n274359 );
nand ( n278344 , n241378 , n209347 );
nand ( n278345 , n278342 , n278343 , n278344 );
buf ( n278346 , n278345 );
not ( n278347 , n205181 );
not ( n278348 , n51381 );
or ( n278349 , n278347 , n278348 );
nand ( n278350 , n271572 , n271177 );
not ( n278351 , n38053 );
not ( n278352 , n227795 );
or ( n278353 , n278351 , n278352 );
or ( n278354 , n227795 , n38053 );
nand ( n278355 , n278353 , n278354 );
and ( n278356 , n278355 , n234514 );
not ( n278357 , n278355 );
and ( n278358 , n278357 , n234522 );
nor ( n278359 , n278356 , n278358 );
not ( n278360 , n278359 );
and ( n278361 , n278350 , n278360 );
not ( n278362 , n278350 );
and ( n278363 , n278362 , n278359 );
nor ( n278364 , n278361 , n278363 );
or ( n278365 , n278364 , n237358 );
nand ( n278366 , n278349 , n278365 );
buf ( n278367 , n278366 );
not ( n278368 , n270646 );
nand ( n278369 , n256663 , n255701 );
or ( n278370 , n278368 , n278369 );
not ( n278371 , n255701 );
not ( n278372 , n255678 );
or ( n278373 , n278371 , n278372 );
nor ( n278374 , n256663 , n35427 );
nand ( n278375 , n278373 , n278374 );
nand ( n278376 , n234453 , n36177 );
nand ( n278377 , n278370 , n278375 , n278376 );
buf ( n278378 , n278377 );
or ( n278379 , n25328 , n261021 );
or ( n278380 , n25335 , n267843 );
nand ( n278381 , n278379 , n278380 );
buf ( n278382 , n278381 );
buf ( n278383 , n30030 );
buf ( n278384 , n32892 );
not ( n278385 , n272021 );
not ( n278386 , n254613 );
not ( n278387 , n278386 );
or ( n278388 , n278385 , n278387 );
nand ( n278389 , n278388 , n241459 );
or ( n278390 , n278389 , n258643 );
not ( n278391 , n254619 );
nand ( n278392 , n272021 , n258643 );
or ( n278393 , n278391 , n278392 );
nand ( n278394 , n247585 , n36181 );
nand ( n278395 , n278390 , n278393 , n278394 );
buf ( n278396 , n278395 );
not ( n278397 , n263323 );
nand ( n278398 , n278397 , n266840 );
not ( n278399 , n272775 );
or ( n278400 , n278398 , n278399 );
nor ( n278401 , n272767 , n39763 );
nand ( n278402 , n278398 , n278401 );
nand ( n278403 , n55760 , n208141 );
nand ( n278404 , n278400 , n278402 , n278403 );
buf ( n278405 , n278404 );
not ( n278406 , n253904 );
not ( n278407 , n273832 );
nand ( n278408 , n278406 , n278407 );
not ( n278409 , n249395 );
not ( n278410 , n250173 );
not ( n278411 , n249381 );
or ( n278412 , n278410 , n278411 );
not ( n278413 , n250173 );
nand ( n278414 , n278413 , n249388 );
nand ( n278415 , n278412 , n278414 );
not ( n278416 , n278415 );
or ( n278417 , n278409 , n278416 );
or ( n278418 , n278415 , n249395 );
nand ( n278419 , n278417 , n278418 );
not ( n278420 , n278419 );
not ( n278421 , n274532 );
nand ( n278422 , n278420 , n278421 );
or ( n278423 , n278408 , n278422 );
not ( n278424 , n278420 );
not ( n278425 , n278407 );
or ( n278426 , n278424 , n278425 );
nor ( n278427 , n278421 , n258327 );
nand ( n278428 , n278426 , n278427 );
nand ( n278429 , n37728 , n31030 );
nand ( n278430 , n278423 , n278428 , n278429 );
buf ( n278431 , n278430 );
not ( n278432 , n42995 );
not ( n278433 , n243222 );
or ( n278434 , n278432 , n278433 );
or ( n278435 , n243222 , n42995 );
nand ( n278436 , n278434 , n278435 );
not ( n278437 , n278436 );
not ( n278438 , n243226 );
or ( n278439 , n278437 , n278438 );
or ( n278440 , n243226 , n278436 );
nand ( n278441 , n278439 , n278440 );
nor ( n278442 , n278441 , n249531 );
not ( n278443 , n273566 );
nand ( n278444 , n278442 , n273249 , n278443 );
not ( n278445 , n278441 );
not ( n278446 , n278445 );
not ( n278447 , n273249 );
or ( n278448 , n278446 , n278447 );
nor ( n278449 , n278443 , n55152 );
nand ( n278450 , n278448 , n278449 );
nand ( n278451 , n252711 , n208085 );
nand ( n278452 , n278444 , n278450 , n278451 );
buf ( n278453 , n278452 );
not ( n278454 , n252462 );
not ( n278455 , n231413 );
not ( n278456 , n250496 );
or ( n278457 , n278455 , n278456 );
not ( n278458 , n231413 );
nand ( n278459 , n278458 , n255291 );
nand ( n278460 , n278457 , n278459 );
and ( n278461 , n278460 , n244190 );
not ( n278462 , n278460 );
and ( n278463 , n278462 , n260370 );
nor ( n278464 , n278461 , n278463 );
not ( n278465 , n278464 );
nor ( n278466 , n278454 , n278465 );
nand ( n278467 , n277616 , n278466 );
not ( n278468 , n252462 );
not ( n278469 , n277613 );
not ( n278470 , n278469 );
or ( n278471 , n278468 , n278470 );
nor ( n278472 , n278464 , n55152 );
nand ( n278473 , n278471 , n278472 );
nand ( n278474 , n231444 , n37063 );
nand ( n278475 , n278467 , n278473 , n278474 );
buf ( n278476 , n278475 );
or ( n278477 , n25328 , n259768 );
or ( n278478 , n226822 , n277200 );
nand ( n278479 , n278477 , n278478 );
buf ( n278480 , n278479 );
not ( n278481 , n270285 );
not ( n278482 , n270273 );
nand ( n278483 , n278481 , n278482 );
or ( n278484 , n268474 , n278483 );
nand ( n278485 , n268487 , n278483 );
nand ( n278486 , n239240 , n28697 );
nand ( n278487 , n278484 , n278485 , n278486 );
buf ( n278488 , n278487 );
buf ( n278489 , n39078 );
buf ( n278490 , n27742 );
nand ( n278491 , n273190 , n272711 );
nand ( n278492 , n266322 , n273198 );
or ( n278493 , n278491 , n278492 );
not ( n278494 , n273198 );
not ( n278495 , n273190 );
or ( n278496 , n278494 , n278495 );
nor ( n278497 , n266322 , n256413 );
nand ( n278498 , n278496 , n278497 );
nand ( n278499 , n49054 , n33969 );
nand ( n278500 , n278493 , n278498 , n278499 );
buf ( n278501 , n278500 );
not ( n278502 , n265866 );
not ( n278503 , n240031 );
not ( n278504 , n40194 );
or ( n278505 , n278503 , n278504 );
not ( n278506 , n240031 );
nand ( n278507 , n278506 , n40203 );
nand ( n278508 , n278505 , n278507 );
and ( n278509 , n278508 , n251346 );
not ( n278510 , n278508 );
and ( n278511 , n278510 , n251350 );
nor ( n278512 , n278509 , n278511 );
not ( n278513 , n278512 );
nand ( n278514 , n278513 , n268737 );
or ( n278515 , n278502 , n278514 );
not ( n278516 , n278513 );
not ( n278517 , n265847 );
or ( n278518 , n278516 , n278517 );
nor ( n278519 , n268737 , n234440 );
nand ( n278520 , n278518 , n278519 );
nand ( n278521 , n50615 , n30317 );
nand ( n278522 , n278515 , n278520 , n278521 );
buf ( n278523 , n278522 );
or ( n278524 , n25328 , n274544 );
not ( n278525 , RI19a8db18_2699);
or ( n278526 , n226822 , n278525 );
nand ( n278527 , n278524 , n278526 );
buf ( n278528 , n278527 );
xor ( n278529 , n51664 , n267305 );
xnor ( n278530 , n278529 , n260340 );
not ( n278531 , n278530 );
nand ( n278532 , n278531 , n262961 );
not ( n278533 , n248938 );
not ( n278534 , n278533 );
not ( n278535 , n250099 );
or ( n278536 , n278534 , n278535 );
or ( n278537 , n250102 , n278533 );
nand ( n278538 , n278536 , n278537 );
and ( n278539 , n278538 , n250105 );
not ( n278540 , n278538 );
and ( n278541 , n278540 , n250108 );
nor ( n278542 , n278539 , n278541 );
nor ( n278543 , n260649 , n278542 );
or ( n278544 , n278532 , n278543 );
nor ( n278545 , n278531 , n249531 );
nand ( n278546 , n278545 , n278543 );
nand ( n278547 , n234453 , n38068 );
nand ( n278548 , n278544 , n278546 , n278547 );
buf ( n278549 , n278548 );
not ( n278550 , n270693 );
not ( n278551 , n242618 );
not ( n278552 , n244939 );
or ( n278553 , n278551 , n278552 );
not ( n278554 , n242618 );
nand ( n278555 , n278554 , n244954 );
nand ( n278556 , n278553 , n278555 );
and ( n278557 , n278556 , n254867 );
not ( n278558 , n278556 );
and ( n278559 , n278558 , n254874 );
nor ( n278560 , n278557 , n278559 );
not ( n278561 , n278560 );
nand ( n278562 , n278550 , n278561 );
not ( n278563 , n270711 );
or ( n278564 , n278562 , n278563 );
nand ( n278565 , n278562 , n271847 );
nand ( n278566 , n234453 , n35504 );
nand ( n278567 , n278564 , n278565 , n278566 );
buf ( n278568 , n278567 );
or ( n278569 , n25328 , n269276 );
or ( n278570 , n25335 , n267289 );
nand ( n278571 , n278569 , n278570 );
buf ( n278572 , n278571 );
not ( n278573 , RI19a9af70_2605);
or ( n278574 , n25328 , n278573 );
not ( n278575 , RI19a90f20_2676);
or ( n278576 , n25335 , n278575 );
nand ( n278577 , n278574 , n278576 );
buf ( n278578 , n278577 );
not ( n278579 , n275766 );
not ( n278580 , n275781 );
or ( n278581 , n278579 , n278580 );
nor ( n278582 , n278225 , n226003 );
nand ( n278583 , n278581 , n278582 );
nor ( n278584 , n275767 , n234021 );
nand ( n278585 , n278584 , n275781 , n278225 );
nand ( n278586 , n256673 , n34667 );
nand ( n278587 , n278583 , n278585 , n278586 );
buf ( n278588 , n278587 );
not ( n278589 , n235749 );
not ( n278590 , n245743 );
or ( n278591 , n278589 , n278590 );
or ( n278592 , n245743 , n235749 );
nand ( n278593 , n278591 , n278592 );
and ( n278594 , n278593 , n245794 );
not ( n278595 , n278593 );
and ( n278596 , n278595 , n245799 );
nor ( n278597 , n278594 , n278596 );
not ( n278598 , n278597 );
nand ( n278599 , n278598 , n258918 );
nand ( n278600 , n274152 , n274609 );
or ( n278601 , n278599 , n278600 );
not ( n278602 , n274152 );
not ( n278603 , n278598 );
or ( n278604 , n278602 , n278603 );
nand ( n278605 , n278604 , n274616 );
nand ( n278606 , n251465 , n36822 );
nand ( n278607 , n278601 , n278605 , n278606 );
buf ( n278608 , n278607 );
not ( n278609 , RI19ab0c30_2448);
or ( n278610 , n25328 , n278609 );
or ( n278611 , n25335 , n274034 );
nand ( n278612 , n278610 , n278611 );
buf ( n278613 , n278612 );
not ( n278614 , RI19ad0238_2210);
or ( n278615 , n25335 , n278614 );
nand ( n278616 , RI1754a630_70 , RI1754a5b8_71);
or ( n278617 , n273849 , n278616 );
not ( n278618 , n249125 );
nand ( n278619 , n278618 , RI1754a810_66);
nand ( n278620 , n278615 , n278617 , n278619 );
buf ( n278621 , n278620 );
nor ( n278622 , n276774 , n276750 );
or ( n278623 , n277736 , n278622 );
nand ( n278624 , n276867 , n278622 );
nand ( n278625 , n247585 , n32000 );
nand ( n278626 , n278623 , n278624 , n278625 );
buf ( n278627 , n278626 );
buf ( n278628 , n204932 );
buf ( n278629 , n33057 );
not ( n278630 , RI19ac0d88_2324);
or ( n278631 , n25328 , n278630 );
not ( n278632 , RI19ab7f80_2395);
or ( n278633 , n25335 , n278632 );
nand ( n278634 , n278631 , n278633 );
buf ( n278635 , n278634 );
buf ( n278636 , n216999 );
not ( n278637 , n36936 );
not ( n278638 , n51381 );
or ( n278639 , n278637 , n278638 );
nand ( n278640 , n270165 , n271900 );
and ( n278641 , n278640 , n270175 );
not ( n278642 , n278640 );
not ( n278643 , n270175 );
and ( n278644 , n278642 , n278643 );
nor ( n278645 , n278641 , n278644 );
or ( n278646 , n278645 , n49959 );
nand ( n278647 , n278639 , n278646 );
buf ( n278648 , n278647 );
not ( n278649 , n33914 );
not ( n278650 , n37728 );
or ( n278651 , n278649 , n278650 );
nand ( n278652 , n268497 , n268485 );
not ( n278653 , n270285 );
and ( n278654 , n278652 , n278653 );
not ( n278655 , n278652 );
and ( n278656 , n278655 , n270285 );
nor ( n278657 , n278654 , n278656 );
or ( n278658 , n278657 , n251462 );
nand ( n278659 , n278651 , n278658 );
buf ( n278660 , n278659 );
not ( n278661 , n27827 );
not ( n278662 , n51381 );
or ( n278663 , n278661 , n278662 );
not ( n278664 , n237846 );
not ( n278665 , n254916 );
or ( n278666 , n278664 , n278665 );
not ( n278667 , n237846 );
nand ( n278668 , n278667 , n251684 );
nand ( n278669 , n278666 , n278668 );
and ( n278670 , n278669 , n260132 );
not ( n278671 , n278669 );
and ( n278672 , n278671 , n251692 );
nor ( n278673 , n278670 , n278672 );
not ( n278674 , n41622 );
not ( n278675 , n233026 );
or ( n278676 , n278674 , n278675 );
not ( n278677 , n41622 );
nand ( n278678 , n278677 , n233035 );
nand ( n278679 , n278676 , n278678 );
and ( n278680 , n278679 , n233084 );
not ( n278681 , n278679 );
and ( n278682 , n278681 , n233091 );
nor ( n278683 , n278680 , n278682 );
nand ( n278684 , n278673 , n278683 );
not ( n278685 , n278684 );
not ( n278686 , n256632 );
and ( n278687 , n278685 , n278686 );
and ( n278688 , n278684 , n256618 );
nor ( n278689 , n278687 , n278688 );
or ( n278690 , n278689 , n238223 );
nand ( n278691 , n278663 , n278690 );
buf ( n278692 , n278691 );
not ( n278693 , n210737 );
not ( n278694 , n244789 );
or ( n278695 , n278693 , n278694 );
nand ( n278696 , n276453 , n273912 );
and ( n278697 , n278696 , n267981 );
not ( n278698 , n278696 );
not ( n278699 , n267981 );
and ( n278700 , n278698 , n278699 );
nor ( n278701 , n278697 , n278700 );
or ( n278702 , n278701 , n260861 );
nand ( n278703 , n278695 , n278702 );
buf ( n278704 , n278703 );
not ( n278705 , n265467 );
not ( n278706 , n271134 );
nand ( n278707 , n278706 , n265478 );
or ( n278708 , n278705 , n278707 );
nand ( n278709 , n254151 , n278707 );
nand ( n278710 , n256673 , n34194 );
nand ( n278711 , n278708 , n278709 , n278710 );
buf ( n278712 , n278711 );
not ( n278713 , n33072 );
not ( n278714 , n255116 );
or ( n278715 , n278713 , n278714 );
not ( n278716 , n277664 );
nand ( n278717 , n278716 , n276222 );
and ( n278718 , n278717 , n259269 );
not ( n278719 , n278717 );
and ( n278720 , n278719 , n259268 );
nor ( n278721 , n278718 , n278720 );
or ( n278722 , n278721 , n251498 );
nand ( n278723 , n278715 , n278722 );
buf ( n278724 , n278723 );
nand ( n278725 , n259545 , n259558 );
or ( n278726 , n278725 , n275358 );
nor ( n278727 , n275357 , n234440 );
nand ( n278728 , n278727 , n278725 );
nand ( n278729 , n239240 , n40503 );
nand ( n278730 , n278726 , n278728 , n278729 );
buf ( n278731 , n278730 );
or ( n278732 , n25328 , n276559 );
not ( n278733 , RI19a97208_2632);
or ( n278734 , n25335 , n278733 );
nand ( n278735 , n278732 , n278734 );
buf ( n278736 , n278735 );
nand ( n278737 , n274981 , n41937 );
or ( n278738 , n40467 , n278737 );
not ( n278739 , n41937 );
not ( n278740 , n40464 );
or ( n278741 , n278739 , n278740 );
nor ( n278742 , n274981 , n250431 );
nand ( n278743 , n278741 , n278742 );
nand ( n278744 , n31576 , n32209 );
nand ( n278745 , n278738 , n278743 , n278744 );
buf ( n278746 , n278745 );
buf ( n278747 , n205559 );
buf ( n278748 , n242473 );
buf ( n278749 , n29639 );
nor ( n278750 , n257526 , n237384 );
not ( n278751 , n44050 );
not ( n278752 , n54325 );
or ( n278753 , n278751 , n278752 );
not ( n278754 , n44050 );
nand ( n278755 , n278754 , n255320 );
nand ( n278756 , n278753 , n278755 );
and ( n278757 , n278756 , n234098 );
not ( n278758 , n278756 );
and ( n278759 , n278758 , n234107 );
nor ( n278760 , n278757 , n278759 );
nor ( n278761 , n257538 , n278760 );
nand ( n278762 , n278750 , n278761 );
not ( n278763 , n278760 );
not ( n278764 , n278763 );
not ( n278765 , n257526 );
not ( n278766 , n278765 );
or ( n278767 , n278764 , n278766 );
nor ( n278768 , n257539 , n274333 );
nand ( n278769 , n278767 , n278768 );
nand ( n278770 , n35431 , n205157 );
nand ( n278771 , n278762 , n278769 , n278770 );
buf ( n278772 , n278771 );
buf ( n278773 , n28714 );
not ( n278774 , n257867 );
not ( n278775 , n278774 );
not ( n278776 , n248240 );
not ( n278777 , n240316 );
or ( n278778 , n278776 , n278777 );
or ( n278779 , n240316 , n248240 );
nand ( n278780 , n278778 , n278779 );
and ( n278781 , n278780 , n240505 );
not ( n278782 , n278780 );
and ( n278783 , n278782 , n240508 );
nor ( n278784 , n278781 , n278783 );
not ( n278785 , n278784 );
not ( n278786 , n278785 );
or ( n278787 , n278775 , n278786 );
not ( n278788 , n234524 );
nor ( n278789 , n278788 , n253358 );
nand ( n278790 , n278787 , n278789 );
nand ( n278791 , n278785 , n257870 , n278788 );
nand ( n278792 , n250916 , n41436 );
nand ( n278793 , n278790 , n278791 , n278792 );
buf ( n278794 , n278793 );
not ( n278795 , RI19aa7888_2513);
or ( n278796 , n25328 , n278795 );
not ( n278797 , RI19a9de50_2585);
or ( n278798 , n25335 , n278797 );
nand ( n278799 , n278796 , n278798 );
buf ( n278800 , n278799 );
not ( n278801 , n271998 );
not ( n278802 , n239600 );
not ( n278803 , n260122 );
or ( n278804 , n278802 , n278803 );
or ( n278805 , n260122 , n239600 );
nand ( n278806 , n278804 , n278805 );
and ( n278807 , n278806 , n237746 );
not ( n278808 , n278806 );
and ( n278809 , n278808 , n261776 );
nor ( n278810 , n278807 , n278809 );
not ( n278811 , n239357 );
not ( n278812 , n278811 );
not ( n278813 , n252917 );
or ( n278814 , n278812 , n278813 );
not ( n278815 , n278811 );
nand ( n278816 , n278815 , n252922 );
nand ( n278817 , n278814 , n278816 );
and ( n278818 , n278817 , n258058 );
not ( n278819 , n278817 );
and ( n278820 , n278819 , n258061 );
nor ( n278821 , n278818 , n278820 );
nand ( n278822 , n278810 , n278821 );
or ( n278823 , n278801 , n278822 );
not ( n278824 , n278821 );
not ( n278825 , n271979 );
or ( n278826 , n278824 , n278825 );
nor ( n278827 , n278810 , n247698 );
nand ( n278828 , n278826 , n278827 );
nand ( n278829 , n46083 , n42363 );
nand ( n278830 , n278823 , n278828 , n278829 );
buf ( n278831 , n278830 );
or ( n278832 , n25328 , n266944 );
or ( n278833 , n25335 , n264139 );
nand ( n278834 , n278832 , n278833 );
buf ( n278835 , n278834 );
or ( n278836 , n226819 , n268961 );
or ( n278837 , n25335 , n274029 );
nand ( n278838 , n278836 , n278837 );
buf ( n278839 , n278838 );
not ( n278840 , n27699 );
not ( n278841 , n51381 );
or ( n278842 , n278840 , n278841 );
nand ( n278843 , n275841 , n275851 );
not ( n278844 , n272808 );
and ( n278845 , n278843 , n278844 );
not ( n278846 , n278843 );
and ( n278847 , n278846 , n272808 );
nor ( n278848 , n278845 , n278847 );
or ( n278849 , n278848 , n251498 );
nand ( n278850 , n278842 , n278849 );
buf ( n278851 , n278850 );
not ( n278852 , n260507 );
not ( n278853 , n232996 );
not ( n278854 , n239398 );
or ( n278855 , n278853 , n278854 );
not ( n278856 , n232996 );
nand ( n278857 , n278856 , n239390 );
nand ( n278858 , n278855 , n278857 );
and ( n278859 , n278858 , n249021 );
not ( n278860 , n278858 );
not ( n278861 , n249021 );
and ( n278862 , n278860 , n278861 );
nor ( n278863 , n278859 , n278862 );
nand ( n278864 , n278852 , n278863 );
not ( n278865 , n259738 );
not ( n278866 , n227495 );
and ( n278867 , n278865 , n278866 );
and ( n278868 , n259738 , n227495 );
nor ( n278869 , n278867 , n278868 );
and ( n278870 , n278869 , n259744 );
not ( n278871 , n278869 );
and ( n278872 , n278871 , n259747 );
nor ( n278873 , n278870 , n278872 );
nand ( n278874 , n278873 , n241373 );
or ( n278875 , n278864 , n278874 );
not ( n278876 , n278873 );
not ( n278877 , n278863 );
or ( n278878 , n278876 , n278877 );
nand ( n278879 , n278878 , n233973 );
or ( n278880 , n278879 , n278852 );
nand ( n278881 , n252711 , n25586 );
nand ( n278882 , n278875 , n278880 , n278881 );
buf ( n278883 , n278882 );
not ( n278884 , n271400 );
not ( n278885 , n217056 );
and ( n278886 , n278884 , n278885 );
not ( n278887 , n244309 );
not ( n278888 , n278887 );
not ( n278889 , n29962 );
or ( n278890 , n278888 , n278889 );
or ( n278891 , n29962 , n278887 );
nand ( n278892 , n278890 , n278891 );
and ( n278893 , n278892 , n256366 );
not ( n278894 , n278892 );
and ( n278895 , n278894 , n263797 );
nor ( n278896 , n278893 , n278895 );
nor ( n278897 , n278896 , n221279 );
not ( n278898 , n270760 );
nor ( n278899 , n278898 , n270770 );
and ( n278900 , n278897 , n278899 );
nor ( n278901 , n278886 , n278900 );
nand ( n278902 , n278896 , n239934 );
not ( n278903 , n278902 );
nand ( n278904 , n278903 , n278898 );
nor ( n278905 , n270760 , n254150 );
nand ( n278906 , n278905 , n270770 );
nand ( n278907 , n278901 , n278904 , n278906 );
buf ( n278908 , n278907 );
not ( n278909 , n33251 );
nand ( n278910 , n278909 , n249009 );
not ( n278911 , n278910 );
not ( n278912 , n247654 );
not ( n278913 , n278912 );
not ( n278914 , n48015 );
or ( n278915 , n278913 , n278914 );
not ( n278916 , n278912 );
nand ( n278917 , n278916 , n48019 );
nand ( n278918 , n278915 , n278917 );
and ( n278919 , n278918 , n225998 );
not ( n278920 , n278918 );
and ( n278921 , n278920 , n48238 );
nor ( n278922 , n278919 , n278921 );
not ( n278923 , n278922 );
nand ( n278924 , n278923 , n34455 );
not ( n278925 , n278924 );
and ( n278926 , n278911 , n278925 );
and ( n278927 , n257764 , n31020 );
nor ( n278928 , n278926 , n278927 );
not ( n278929 , n33256 );
nand ( n278930 , n278929 , n278922 );
nand ( n278931 , n278922 , n244809 );
not ( n278932 , n278931 );
nand ( n278933 , n278932 , n34454 );
nand ( n278934 , n278928 , n278930 , n278933 );
buf ( n278935 , n278934 );
not ( n278936 , n253502 );
nand ( n278937 , n278035 , n278936 );
or ( n278938 , n278025 , n278937 );
not ( n278939 , n278035 );
not ( n278940 , n278024 );
or ( n278941 , n278939 , n278940 );
nor ( n278942 , n278936 , n37724 );
nand ( n278943 , n278941 , n278942 );
nand ( n278944 , n241976 , n36211 );
nand ( n278945 , n278938 , n278943 , n278944 );
buf ( n278946 , n278945 );
not ( n278947 , RI19a9e6c0_2581);
or ( n278948 , n25328 , n278947 );
or ( n278949 , n25335 , n275599 );
nand ( n278950 , n278948 , n278949 );
buf ( n278951 , n278950 );
not ( n278952 , n273055 );
nand ( n278953 , n275726 , n273052 );
or ( n278954 , n278952 , n278953 );
not ( n278955 , n273052 );
not ( n278956 , n273039 );
or ( n278957 , n278955 , n278956 );
nor ( n278958 , n275726 , n237384 );
nand ( n278959 , n278957 , n278958 );
nand ( n278960 , n246460 , n28458 );
nand ( n278961 , n278954 , n278959 , n278960 );
buf ( n278962 , n278961 );
nand ( n278963 , n270708 , n259009 );
nand ( n278964 , n278560 , n271844 );
or ( n278965 , n278963 , n278964 );
not ( n278966 , n271844 );
not ( n278967 , n270708 );
or ( n278968 , n278966 , n278967 );
nor ( n278969 , n278560 , n251361 );
nand ( n278970 , n278968 , n278969 );
nand ( n278971 , n245701 , n25402 );
nand ( n278972 , n278965 , n278970 , n278971 );
buf ( n278973 , n278972 );
or ( n278974 , n25328 , n273490 );
not ( n278975 , RI19abdbd8_2352);
or ( n278976 , n25336 , n278975 );
nand ( n278977 , n278974 , n278976 );
buf ( n278978 , n278977 );
nand ( n278979 , n265546 , n254988 );
or ( n278980 , n272042 , n278979 );
not ( n278981 , n272041 );
nand ( n278982 , n278981 , n237385 );
not ( n278983 , n278982 );
nand ( n278984 , n278983 , n278979 );
nand ( n278985 , n41945 , n36462 );
nand ( n278986 , n278980 , n278984 , n278985 );
buf ( n278987 , n278986 );
not ( n278988 , RI19ac1a30_2317);
or ( n278989 , n25328 , n278988 );
or ( n278990 , n25336 , n260289 );
nand ( n278991 , n278989 , n278990 );
buf ( n278992 , n278991 );
not ( n278993 , RI1754b440_40);
or ( n278994 , n249128 , n278993 );
nand ( n278995 , n249131 , n40554 );
nand ( n278996 , n278994 , n278995 );
buf ( n278997 , n278996 );
not ( n278998 , n33742 );
not ( n278999 , n239240 );
or ( n279000 , n278998 , n278999 );
nand ( n279001 , n265508 , n265518 );
not ( n279002 , n242636 );
not ( n279003 , n244939 );
or ( n279004 , n279002 , n279003 );
not ( n279005 , n242636 );
nand ( n279006 , n279005 , n244954 );
nand ( n279007 , n279004 , n279006 );
and ( n279008 , n279007 , n254867 );
not ( n279009 , n279007 );
and ( n279010 , n279009 , n254874 );
nor ( n279011 , n279008 , n279010 );
not ( n279012 , n279011 );
and ( n279013 , n279001 , n279012 );
not ( n279014 , n279001 );
and ( n279015 , n279014 , n279011 );
nor ( n279016 , n279013 , n279015 );
or ( n279017 , n279016 , n234110 );
nand ( n279018 , n279000 , n279017 );
buf ( n279019 , n279018 );
not ( n279020 , n34890 );
not ( n279021 , n245701 );
or ( n279022 , n279020 , n279021 );
nand ( n279023 , n250966 , n261369 );
not ( n279024 , n250946 );
and ( n279025 , n279023 , n279024 );
not ( n279026 , n279023 );
and ( n279027 , n279026 , n250946 );
nor ( n279028 , n279025 , n279027 );
or ( n279029 , n279028 , n260861 );
nand ( n279030 , n279022 , n279029 );
buf ( n279031 , n279030 );
not ( n279032 , n276352 );
nand ( n279033 , n275907 , n277306 );
or ( n279034 , n279032 , n279033 );
not ( n279035 , n277306 );
not ( n279036 , n276345 );
or ( n279037 , n279035 , n279036 );
nor ( n279038 , n275907 , n55152 );
nand ( n279039 , n279037 , n279038 );
nand ( n279040 , n31577 , n32066 );
nand ( n279041 , n279034 , n279039 , n279040 );
buf ( n279042 , n279041 );
nor ( n279043 , n256934 , n263278 );
nand ( n279044 , n231964 , n279043 );
nor ( n279045 , n263277 , n235732 );
not ( n279046 , n54199 );
nand ( n279047 , n279046 , n256935 );
nand ( n279048 , n279045 , n279047 );
nand ( n279049 , n244484 , n32289 );
nand ( n279050 , n279044 , n279048 , n279049 );
buf ( n279051 , n279050 );
not ( n279052 , n29354 );
not ( n279053 , n51381 );
or ( n279054 , n279052 , n279053 );
nand ( n279055 , n258112 , n240521 );
not ( n279056 , n258123 );
and ( n279057 , n279055 , n279056 );
not ( n279058 , n279055 );
and ( n279059 , n279058 , n258123 );
nor ( n279060 , n279057 , n279059 );
or ( n279061 , n279060 , n256214 );
nand ( n279062 , n279054 , n279061 );
buf ( n279063 , n279062 );
not ( n279064 , n260429 );
nand ( n279065 , n260065 , n269405 );
or ( n279066 , n279064 , n279065 );
not ( n279067 , n260065 );
not ( n279068 , n260043 );
not ( n279069 , n279068 );
or ( n279070 , n279067 , n279069 );
nor ( n279071 , n269405 , n256413 );
nand ( n279072 , n279070 , n279071 );
nand ( n279073 , n49054 , n41503 );
nand ( n279074 , n279066 , n279072 , n279073 );
buf ( n279075 , n279074 );
nand ( n279076 , n257684 , n235051 );
nand ( n279077 , n278247 , n257708 );
or ( n279078 , n279076 , n279077 );
not ( n279079 , n278247 );
not ( n279080 , n257684 );
or ( n279081 , n279079 , n279080 );
nor ( n279082 , n257708 , n53680 );
nand ( n279083 , n279081 , n279082 );
nand ( n279084 , n238114 , n30652 );
nand ( n279085 , n279078 , n279083 , n279084 );
buf ( n279086 , n279085 );
not ( n279087 , n29464 );
not ( n279088 , n244606 );
or ( n279089 , n279087 , n279088 );
not ( n279090 , RI1754adb0_54);
or ( n279091 , n269544 , n279090 );
nand ( n279092 , n279089 , n279091 );
buf ( n279093 , n279092 );
not ( n279094 , n255347 );
nand ( n279095 , n255369 , n279094 );
not ( n279096 , n233886 );
not ( n279097 , n279096 );
not ( n279098 , n244273 );
or ( n279099 , n279097 , n279098 );
not ( n279100 , n279096 );
nand ( n279101 , n279100 , n244282 );
nand ( n279102 , n279099 , n279101 );
and ( n279103 , n279102 , n258153 );
not ( n279104 , n279102 );
and ( n279105 , n279104 , n244347 );
nor ( n279106 , n279103 , n279105 );
not ( n279107 , n279106 );
nor ( n279108 , n279107 , n234818 );
not ( n279109 , n279108 );
or ( n279110 , n279095 , n279109 );
nor ( n279111 , n279106 , n55146 );
nand ( n279112 , n279095 , n279111 );
nand ( n279113 , n241378 , n30856 );
nand ( n279114 , n279110 , n279112 , n279113 );
buf ( n279115 , n279114 );
not ( n279116 , n37052 );
not ( n279117 , n244606 );
or ( n279118 , n279116 , n279117 );
not ( n279119 , RI1754c3b8_7);
or ( n279120 , n244611 , n279119 );
nand ( n279121 , n279118 , n279120 );
buf ( n279122 , n279121 );
not ( n279123 , n273145 );
not ( n279124 , n266740 );
not ( n279125 , n236079 );
not ( n279126 , n279125 );
not ( n279127 , n251082 );
not ( n279128 , n279127 );
or ( n279129 , n279126 , n279128 );
nand ( n279130 , n251082 , n236079 );
nand ( n279131 , n279129 , n279130 );
not ( n279132 , n279131 );
and ( n279133 , n279124 , n279132 );
and ( n279134 , n251029 , n279131 );
nor ( n279135 , n279133 , n279134 );
nand ( n279136 , n279123 , n279135 );
not ( n279137 , n272984 );
or ( n279138 , n279136 , n279137 );
nand ( n279139 , n279135 , n272977 );
nand ( n279140 , n279139 , n273145 , n260879 );
nand ( n279141 , n50615 , n30230 );
nand ( n279142 , n279138 , n279140 , n279141 );
buf ( n279143 , n279142 );
not ( n279144 , n255789 );
not ( n279145 , n246548 );
or ( n279146 , n279144 , n279145 );
not ( n279147 , n255789 );
nand ( n279148 , n279147 , n246553 );
nand ( n279149 , n279146 , n279148 );
and ( n279150 , n279149 , n246654 );
not ( n279151 , n279149 );
and ( n279152 , n279151 , n246661 );
nor ( n279153 , n279150 , n279152 );
nand ( n279154 , n279153 , n259619 );
not ( n279155 , n261634 );
nand ( n279156 , n256462 , n279155 );
or ( n279157 , n279154 , n279156 );
not ( n279158 , n279155 );
not ( n279159 , n279153 );
or ( n279160 , n279158 , n279159 );
nor ( n279161 , n256462 , n251361 );
nand ( n279162 , n279160 , n279161 );
nand ( n279163 , n31576 , n208643 );
nand ( n279164 , n279157 , n279162 , n279163 );
buf ( n279165 , n279164 );
not ( n279166 , n266113 );
not ( n279167 , n269475 );
or ( n279168 , n279166 , n279167 );
nor ( n279169 , n278057 , n47173 );
nand ( n279170 , n279168 , n279169 );
not ( n279171 , n278057 );
nor ( n279172 , n279171 , n266112 );
nand ( n279173 , n269472 , n279172 );
nand ( n279174 , n39767 , n28836 );
nand ( n279175 , n279170 , n279173 , n279174 );
buf ( n279176 , n279175 );
or ( n279177 , n25328 , n273025 );
or ( n279178 , n25335 , n264542 );
nand ( n279179 , n279177 , n279178 );
buf ( n279180 , n279179 );
nand ( n279181 , n276849 , n255921 );
or ( n279182 , n255912 , n279181 );
nand ( n279183 , n277676 , n279181 );
nand ( n279184 , n256292 , n29711 );
nand ( n279185 , n279182 , n279183 , n279184 );
buf ( n279186 , n279185 );
not ( n279187 , n253019 );
nand ( n279188 , n279187 , n257527 );
not ( n279189 , n279188 );
nand ( n279190 , n253031 , n255035 );
not ( n279191 , n279190 );
and ( n279192 , n279189 , n279191 );
and ( n279193 , n245702 , n204901 );
nor ( n279194 , n279192 , n279193 );
not ( n279195 , n253020 );
nand ( n279196 , n279195 , n255036 );
nand ( n279197 , n255052 , n253030 );
nand ( n279198 , n279194 , n279196 , n279197 );
buf ( n279199 , n279198 );
and ( n279200 , n275215 , n274810 );
and ( n279201 , n41945 , n35304 );
nor ( n279202 , n279200 , n279201 );
not ( n279203 , n260107 );
not ( n279204 , n251526 );
or ( n279205 , n279203 , n279204 );
or ( n279206 , n249693 , n260107 );
nand ( n279207 , n279205 , n279206 );
not ( n279208 , n279207 );
not ( n279209 , n279208 );
not ( n279210 , n249750 );
or ( n279211 , n279209 , n279210 );
nand ( n279212 , n249759 , n279207 );
nand ( n279213 , n279211 , n279212 );
nand ( n279214 , n274812 , n279213 );
not ( n279215 , n279213 );
nand ( n279216 , n275219 , n274811 , n279215 );
nand ( n279217 , n279202 , n279214 , n279216 );
buf ( n279218 , n279217 );
not ( n279219 , RI19a831e0_2772);
or ( n279220 , n25328 , n279219 );
not ( n279221 , RI19ac8330_2268);
or ( n279222 , n226822 , n279221 );
nand ( n279223 , n279220 , n279222 );
buf ( n279224 , n279223 );
or ( n279225 , n226819 , n259448 );
not ( n279226 , RI19a8c498_2709);
or ( n279227 , n25335 , n279226 );
nand ( n279228 , n279225 , n279227 );
buf ( n279229 , n279228 );
or ( n279230 , n233507 , n265417 );
not ( n279231 , RI19ac5bd0_2286);
or ( n279232 , n25336 , n279231 );
nand ( n279233 , n279230 , n279232 );
buf ( n279234 , n279233 );
not ( n279235 , n29314 );
not ( n279236 , n245702 );
or ( n279237 , n279235 , n279236 );
not ( n279238 , n47026 );
not ( n279239 , n252823 );
or ( n279240 , n279238 , n279239 );
not ( n279241 , n47026 );
nand ( n279242 , n279241 , n252831 );
nand ( n279243 , n279240 , n279242 );
and ( n279244 , n279243 , n252837 );
not ( n279245 , n279243 );
and ( n279246 , n279245 , n252834 );
nor ( n279247 , n279244 , n279246 );
nand ( n279248 , n274292 , n279247 );
and ( n279249 , n279248 , n267379 );
not ( n279250 , n279248 );
not ( n279251 , n267379 );
and ( n279252 , n279250 , n279251 );
nor ( n279253 , n279249 , n279252 );
or ( n279254 , n279253 , n253544 );
nand ( n279255 , n279237 , n279254 );
buf ( n279256 , n279255 );
or ( n279257 , n25328 , n277499 );
or ( n279258 , n25335 , n263544 );
nand ( n279259 , n279257 , n279258 );
buf ( n279260 , n279259 );
buf ( n279261 , n39120 );
nand ( n279262 , n277014 , n50945 );
nand ( n279263 , n266389 , n266400 );
or ( n279264 , n279262 , n279263 );
not ( n279265 , n266400 );
not ( n279266 , n277014 );
or ( n279267 , n279265 , n279266 );
nor ( n279268 , n266389 , n46425 );
nand ( n279269 , n279267 , n279268 );
nand ( n279270 , n252711 , n30576 );
nand ( n279271 , n279264 , n279269 , n279270 );
buf ( n279272 , n279271 );
buf ( n279273 , n36152 );
not ( n279274 , n273506 );
nand ( n279275 , n263644 , n260405 );
or ( n279276 , n279274 , n279275 );
not ( n279277 , n263644 );
not ( n279278 , n260374 );
not ( n279279 , n279278 );
or ( n279280 , n279277 , n279279 );
nor ( n279281 , n260405 , n234440 );
nand ( n279282 , n279280 , n279281 );
nand ( n279283 , n237361 , n33904 );
nand ( n279284 , n279276 , n279282 , n279283 );
buf ( n279285 , n279284 );
or ( n279286 , n226819 , n43526 );
not ( n279287 , RI19ab48a8_2419);
or ( n279288 , n25335 , n279287 );
nand ( n279289 , n279286 , n279288 );
buf ( n279290 , n279289 );
buf ( n279291 , n32100 );
not ( n279292 , n268419 );
nand ( n279293 , n268409 , n274265 );
or ( n279294 , n279292 , n279293 );
not ( n279295 , n268409 );
not ( n279296 , n268399 );
not ( n279297 , n279296 );
or ( n279298 , n279295 , n279297 );
nand ( n279299 , n279298 , n275055 );
nand ( n279300 , n41944 , n33592 );
nand ( n279301 , n279294 , n279299 , n279300 );
buf ( n279302 , n279301 );
not ( n279303 , n36199 );
not ( n279304 , n254441 );
or ( n279305 , n279303 , n279304 );
nand ( n279306 , n260891 , n237735 );
not ( n279307 , n237756 );
and ( n279308 , n279306 , n279307 );
not ( n279309 , n279306 );
and ( n279310 , n279309 , n237756 );
nor ( n279311 , n279308 , n279310 );
or ( n279312 , n279311 , n259425 );
nand ( n279313 , n279305 , n279312 );
buf ( n279314 , n279313 );
not ( n279315 , RI19ab7878_2398);
or ( n279316 , n226819 , n279315 );
not ( n279317 , RI19aadd50_2469);
or ( n279318 , n25335 , n279317 );
nand ( n279319 , n279316 , n279318 );
buf ( n279320 , n279319 );
buf ( n279321 , n35700 );
or ( n279322 , n25328 , n257408 );
or ( n279323 , n25335 , n266876 );
nand ( n279324 , n279322 , n279323 );
buf ( n279325 , n279324 );
not ( n279326 , n48113 );
not ( n279327 , n226557 );
or ( n279328 , n279326 , n279327 );
not ( n279329 , n48113 );
nand ( n279330 , n279329 , n48804 );
nand ( n279331 , n279328 , n279330 );
and ( n279332 , n279331 , n260471 );
not ( n279333 , n279331 );
and ( n279334 , n279333 , n259388 );
nor ( n279335 , n279332 , n279334 );
not ( n279336 , n258611 );
buf ( n279337 , n230305 );
not ( n279338 , n279337 );
not ( n279339 , n240052 );
or ( n279340 , n279338 , n279339 );
or ( n279341 , n240052 , n279337 );
nand ( n279342 , n279340 , n279341 );
not ( n279343 , n279342 );
not ( n279344 , n279343 );
or ( n279345 , n279336 , n279344 );
nand ( n279346 , n272973 , n279342 );
nand ( n279347 , n279345 , n279346 );
nor ( n279348 , n279335 , n279347 );
or ( n279349 , n274394 , n279348 );
nor ( n279350 , n274393 , n53680 );
nand ( n279351 , n279350 , n279348 );
nand ( n279352 , n241378 , n29681 );
nand ( n279353 , n279349 , n279351 , n279352 );
buf ( n279354 , n279353 );
nand ( n279355 , n272908 , n222531 );
nand ( n279356 , n274088 , n272912 );
or ( n279357 , n279355 , n279356 );
not ( n279358 , n274088 );
not ( n279359 , n272908 );
or ( n279360 , n279358 , n279359 );
nor ( n279361 , n272912 , n234021 );
nand ( n279362 , n279360 , n279361 );
nand ( n279363 , n256673 , n204932 );
nand ( n279364 , n279357 , n279362 , n279363 );
buf ( n279365 , n279364 );
buf ( n279366 , n31310 );
buf ( n279367 , n38968 );
buf ( n279368 , n29003 );
or ( n279369 , n25328 , n249040 );
or ( n279370 , n226822 , n274940 );
nand ( n279371 , n279369 , n279370 );
buf ( n279372 , n279371 );
or ( n279373 , n25328 , n271943 );
or ( n279374 , n25335 , n270716 );
nand ( n279375 , n279373 , n279374 );
buf ( n279376 , n279375 );
nand ( n279377 , n272529 , n269523 );
not ( n279378 , n269604 );
or ( n279379 , n279377 , n279378 );
nor ( n279380 , n269602 , n38637 );
nand ( n279381 , n279377 , n279380 );
nand ( n279382 , n224937 , n32855 );
nand ( n279383 , n279379 , n279381 , n279382 );
buf ( n279384 , n279383 );
not ( n279385 , n269767 );
nand ( n279386 , n279385 , n222532 );
nand ( n279387 , n269779 , n258018 );
not ( n279388 , n279387 );
or ( n279389 , n279386 , n279388 );
or ( n279390 , n269768 , n279387 );
nand ( n279391 , n35431 , n39078 );
nand ( n279392 , n279389 , n279390 , n279391 );
buf ( n279393 , n279392 );
or ( n279394 , n25328 , n272174 );
or ( n279395 , n25335 , n266446 );
nand ( n279396 , n279394 , n279395 );
buf ( n279397 , n279396 );
nand ( n279398 , n262460 , n273755 );
nand ( n279399 , n258466 , n235051 );
or ( n279400 , n279398 , n279399 );
not ( n279401 , n258466 );
not ( n279402 , n262460 );
or ( n279403 , n279401 , n279402 );
nor ( n279404 , n273755 , n243434 );
nand ( n279405 , n279403 , n279404 );
nand ( n279406 , n31577 , n33162 );
nand ( n279407 , n279400 , n279405 , n279406 );
buf ( n279408 , n279407 );
not ( n279409 , n274595 );
nand ( n279410 , n276114 , n276128 );
or ( n279411 , n279409 , n279410 );
not ( n279412 , n276114 );
not ( n279413 , n274592 );
not ( n279414 , n279413 );
or ( n279415 , n279412 , n279414 );
nor ( n279416 , n276128 , n226003 );
nand ( n279417 , n279415 , n279416 );
nand ( n279418 , n35431 , n38643 );
nand ( n279419 , n279411 , n279417 , n279418 );
buf ( n279420 , n279419 );
nand ( n279421 , n254085 , n276044 );
or ( n279422 , n262864 , n279421 );
not ( n279423 , n262863 );
not ( n279424 , n254085 );
or ( n279425 , n279423 , n279424 );
nor ( n279426 , n276044 , n35427 );
nand ( n279427 , n279425 , n279426 );
nand ( n279428 , n238638 , n33491 );
nand ( n279429 , n279422 , n279427 , n279428 );
buf ( n279430 , n279429 );
nand ( n279431 , n47169 , n223839 );
or ( n279432 , n279431 , n262030 );
not ( n279433 , n262033 );
not ( n279434 , n46424 );
and ( n279435 , n279433 , n279434 );
and ( n279436 , n31577 , n36205 );
nor ( n279437 , n279435 , n279436 );
nor ( n279438 , n262017 , n38637 );
nand ( n279439 , n262030 , n279438 , n46424 );
nand ( n279440 , n279432 , n279437 , n279439 );
buf ( n279441 , n279440 );
buf ( n279442 , n34906 );
not ( n279443 , n276835 );
not ( n279444 , n276848 );
or ( n279445 , n279443 , n279444 );
nand ( n279446 , n279445 , n226010 );
or ( n279447 , n279446 , n255921 );
not ( n279448 , n277680 );
nand ( n279449 , n279448 , n276848 , n255921 );
nand ( n279450 , n48251 , n216868 );
nand ( n279451 , n279447 , n279449 , n279450 );
buf ( n279452 , n279451 );
not ( n279453 , n261239 );
not ( n279454 , n279453 );
not ( n279455 , n264978 );
or ( n279456 , n279454 , n279455 );
nor ( n279457 , n264980 , n258369 );
nand ( n279458 , n279456 , n279457 );
nand ( n279459 , n264978 , n261246 , n264980 );
nand ( n279460 , n31577 , n205247 );
nand ( n279461 , n279458 , n279459 , n279460 );
buf ( n279462 , n279461 );
not ( n279463 , RI19acb300_2246);
or ( n279464 , n25328 , n279463 );
or ( n279465 , n25335 , n270611 );
nand ( n279466 , n279464 , n279465 );
buf ( n279467 , n279466 );
or ( n279468 , n226819 , n262679 );
or ( n279469 , n25335 , n235903 );
nand ( n279470 , n279468 , n279469 );
buf ( n279471 , n279470 );
buf ( n279472 , n34980 );
not ( n279473 , n249400 );
nand ( n279474 , n279473 , n249369 );
or ( n279475 , n277234 , n279474 );
nand ( n279476 , n279474 , n253994 );
nand ( n279477 , n237361 , n208419 );
nand ( n279478 , n279475 , n279476 , n279477 );
buf ( n279479 , n279478 );
not ( n279480 , n30229 );
not ( n279481 , n237361 );
or ( n279482 , n279480 , n279481 );
nand ( n279483 , n278560 , n271843 );
not ( n279484 , n279483 );
not ( n279485 , n270693 );
and ( n279486 , n279484 , n279485 );
and ( n279487 , n279483 , n270693 );
nor ( n279488 , n279486 , n279487 );
or ( n279489 , n279488 , n234818 );
nand ( n279490 , n279482 , n279489 );
buf ( n279491 , n279490 );
or ( n279492 , n25328 , n41957 );
or ( n279493 , n25335 , n276634 );
nand ( n279494 , n279492 , n279493 );
buf ( n279495 , n279494 );
buf ( n279496 , n32124 );
nand ( n279497 , n261694 , n55147 );
not ( n279498 , n265105 );
nand ( n279499 , n261717 , n279498 );
or ( n279500 , n279497 , n279499 );
not ( n279501 , n261717 );
not ( n279502 , n261694 );
or ( n279503 , n279501 , n279502 );
nor ( n279504 , n279498 , n221279 );
nand ( n279505 , n279503 , n279504 );
nand ( n279506 , n35431 , n27737 );
nand ( n279507 , n279500 , n279505 , n279506 );
buf ( n279508 , n279507 );
buf ( n279509 , n37969 );
not ( n279510 , RI19aa0100_2568);
or ( n279511 , n226819 , n279510 );
not ( n279512 , RI19a96290_2639);
or ( n279513 , n25336 , n279512 );
nand ( n279514 , n279511 , n279513 );
buf ( n279515 , n279514 );
not ( n279516 , n53919 );
not ( n279517 , n238400 );
or ( n279518 , n279516 , n279517 );
not ( n279519 , n53919 );
nand ( n279520 , n279519 , n238408 );
nand ( n279521 , n279518 , n279520 );
and ( n279522 , n279521 , n251451 );
not ( n279523 , n279521 );
and ( n279524 , n279523 , n251444 );
nor ( n279525 , n279522 , n279524 );
not ( n279526 , n279525 );
nor ( n279527 , n279526 , n264725 );
or ( n279528 , n268438 , n279527 );
nor ( n279529 , n268437 , n222533 );
nand ( n279530 , n279529 , n279527 );
nand ( n279531 , n238638 , n34702 );
nand ( n279532 , n279528 , n279530 , n279531 );
buf ( n279533 , n279532 );
not ( n279534 , n264600 );
nor ( n279535 , n249841 , n246913 );
not ( n279536 , n279535 );
not ( n279537 , n246914 );
nand ( n279538 , n279537 , n249841 );
nand ( n279539 , n279536 , n279538 );
not ( n279540 , n279539 );
or ( n279541 , n279534 , n279540 );
or ( n279542 , n279539 , n264600 );
nand ( n279543 , n279541 , n279542 );
nor ( n279544 , n279543 , n43968 );
not ( n279545 , n250746 );
not ( n279546 , n32092 );
not ( n279547 , n51269 );
or ( n279548 , n279546 , n279547 );
or ( n279549 , n51269 , n32092 );
nand ( n279550 , n279548 , n279549 );
not ( n279551 , n279550 );
or ( n279552 , n279545 , n279551 );
or ( n279553 , n279550 , n250746 );
nand ( n279554 , n279552 , n279553 );
not ( n279555 , n279554 );
nor ( n279556 , n279555 , n265434 );
nand ( n279557 , n279544 , n279556 );
not ( n279558 , n279543 );
not ( n279559 , n279558 );
not ( n279560 , n279554 );
or ( n279561 , n279559 , n279560 );
nor ( n279562 , n265433 , n252872 );
nand ( n279563 , n279561 , n279562 );
nand ( n279564 , n31577 , n205109 );
nand ( n279565 , n279557 , n279563 , n279564 );
buf ( n279566 , n279565 );
not ( n279567 , n251284 );
not ( n279568 , n279567 );
not ( n279569 , n249006 );
or ( n279570 , n279568 , n279569 );
or ( n279571 , n249939 , n279567 );
nand ( n279572 , n279570 , n279571 );
and ( n279573 , n279572 , n267247 );
not ( n279574 , n279572 );
and ( n279575 , n279574 , n249929 );
nor ( n279576 , n279573 , n279575 );
not ( n279577 , n279576 );
nand ( n279578 , n55732 , n279577 );
or ( n279579 , n261083 , n279578 );
not ( n279580 , n55513 );
not ( n279581 , n55732 );
or ( n279582 , n279580 , n279581 );
nor ( n279583 , n279577 , n234440 );
nand ( n279584 , n279582 , n279583 );
nand ( n279585 , n251712 , n34060 );
nand ( n279586 , n279579 , n279584 , n279585 );
buf ( n279587 , n279586 );
not ( n279588 , n278982 );
nand ( n279589 , n272043 , n265544 );
not ( n279590 , n279589 );
and ( n279591 , n279588 , n279590 );
and ( n279592 , n255116 , n37876 );
nor ( n279593 , n279591 , n279592 );
not ( n279594 , n272042 );
nand ( n279595 , n279594 , n254943 );
not ( n279596 , n254944 );
nand ( n279597 , n279596 , n265543 );
nand ( n279598 , n279593 , n279595 , n279597 );
buf ( n279599 , n279598 );
not ( n279600 , n257384 );
nand ( n279601 , n257395 , n279600 );
nand ( n279602 , n279601 , n265752 , n237385 );
not ( n279603 , n265752 );
nand ( n279604 , n279603 , n271863 , n257395 );
nand ( n279605 , n35431 , n34035 );
nand ( n279606 , n279602 , n279604 , n279605 );
buf ( n279607 , n279606 );
not ( n279608 , n26129 );
not ( n279609 , n245943 );
or ( n279610 , n279608 , n279609 );
nand ( n279611 , n274811 , n279213 );
and ( n279612 , n279611 , n274833 );
not ( n279613 , n279611 );
and ( n279614 , n279613 , n274832 );
nor ( n279615 , n279612 , n279614 );
or ( n279616 , n279615 , n262962 );
nand ( n279617 , n279610 , n279616 );
buf ( n279618 , n279617 );
or ( n279619 , n25328 , n256057 );
not ( n279620 , RI19aca748_2252);
or ( n279621 , n25335 , n279620 );
nand ( n279622 , n279619 , n279621 );
buf ( n279623 , n279622 );
buf ( n279624 , n33026 );
buf ( n279625 , n31633 );
or ( n279626 , n226819 , n267745 );
or ( n279627 , n25335 , n270874 );
nand ( n279628 , n279626 , n279627 );
buf ( n279629 , n279628 );
not ( n279630 , n267595 );
nand ( n279631 , n267592 , n253274 );
or ( n279632 , n279630 , n279631 );
not ( n279633 , n267592 );
not ( n279634 , n267581 );
not ( n279635 , n279634 );
or ( n279636 , n279633 , n279635 );
nand ( n279637 , n279636 , n253275 );
nand ( n279638 , n31577 , n39621 );
nand ( n279639 , n279632 , n279637 , n279638 );
buf ( n279640 , n279639 );
buf ( n279641 , n204839 );
buf ( n279642 , n32132 );
not ( n279643 , n265820 );
not ( n279644 , n268361 );
nand ( n279645 , n252492 , n279644 );
or ( n279646 , n279643 , n279645 );
not ( n279647 , n265818 );
not ( n279648 , n279644 );
or ( n279649 , n279647 , n279648 );
nor ( n279650 , n252492 , n256481 );
nand ( n279651 , n279649 , n279650 );
nand ( n279652 , n238638 , n41831 );
nand ( n279653 , n279646 , n279651 , n279652 );
buf ( n279654 , n279653 );
not ( n279655 , n279247 );
nor ( n279656 , n274292 , n279655 );
nand ( n279657 , n267402 , n279656 );
not ( n279658 , n267398 );
not ( n279659 , n274292 );
not ( n279660 , n279659 );
or ( n279661 , n279658 , n279660 );
nor ( n279662 , n279247 , n37725 );
nand ( n279663 , n279661 , n279662 );
nand ( n279664 , n247744 , n208100 );
nand ( n279665 , n279657 , n279663 , n279664 );
buf ( n279666 , n279665 );
not ( n279667 , n28979 );
not ( n279668 , n55760 );
or ( n279669 , n279667 , n279668 );
not ( n279670 , n267934 );
nand ( n279671 , n279670 , n267942 );
not ( n279672 , n279671 );
not ( n279673 , n276261 );
and ( n279674 , n279672 , n279673 );
and ( n279675 , n279671 , n276261 );
nor ( n279676 , n279674 , n279675 );
or ( n279677 , n279676 , n39763 );
nand ( n279678 , n279669 , n279677 );
buf ( n279679 , n279678 );
not ( n279680 , RI19a85508_2757);
or ( n279681 , n226819 , n279680 );
not ( n279682 , RI19a869a8_2748);
or ( n279683 , n25335 , n279682 );
nand ( n279684 , n279681 , n279683 );
buf ( n279685 , n279684 );
not ( n279686 , n37982 );
not ( n279687 , n239240 );
or ( n279688 , n279686 , n279687 );
nand ( n279689 , n262700 , n262711 );
and ( n279690 , n279689 , n273480 );
not ( n279691 , n279689 );
and ( n279692 , n279691 , n272438 );
nor ( n279693 , n279690 , n279692 );
or ( n279694 , n279693 , n234110 );
nand ( n279695 , n279688 , n279694 );
buf ( n279696 , n279695 );
buf ( n279697 , n238783 );
not ( n279698 , n279697 );
not ( n279699 , n279698 );
not ( n279700 , n247991 );
or ( n279701 , n279699 , n279700 );
nand ( n279702 , n247999 , n279697 );
nand ( n279703 , n279701 , n279702 );
not ( n279704 , n279703 );
not ( n279705 , n261862 );
and ( n279706 , n279704 , n279705 );
and ( n279707 , n279703 , n261862 );
nor ( n279708 , n279706 , n279707 );
not ( n279709 , n279708 );
not ( n279710 , n238946 );
not ( n279711 , n279710 );
not ( n279712 , n229763 );
or ( n279713 , n279711 , n279712 );
or ( n279714 , n229763 , n279710 );
nand ( n279715 , n279713 , n279714 );
and ( n279716 , n279715 , n52223 );
not ( n279717 , n279715 );
and ( n279718 , n279717 , n229991 );
nor ( n279719 , n279716 , n279718 );
nand ( n279720 , n279709 , n279719 );
or ( n279721 , n272712 , n279720 );
not ( n279722 , n272679 );
nand ( n279723 , n279722 , n279720 );
nand ( n279724 , n255116 , n30175 );
nand ( n279725 , n279721 , n279723 , n279724 );
buf ( n279726 , n279725 );
not ( n279727 , n263968 );
nand ( n279728 , n279727 , n246177 );
not ( n279729 , n279728 );
nand ( n279730 , n256529 , n256541 );
not ( n279731 , n279730 );
and ( n279732 , n279729 , n279731 );
and ( n279733 , n37728 , n35542 );
nor ( n279734 , n279732 , n279733 );
not ( n279735 , n263969 );
nand ( n279736 , n279735 , n256540 );
not ( n279737 , n257312 );
nand ( n279738 , n279737 , n256530 );
nand ( n279739 , n279734 , n279736 , n279738 );
buf ( n279740 , n279739 );
nand ( n279741 , n221271 , n235051 );
nand ( n279742 , n254201 , n273783 );
or ( n279743 , n279741 , n279742 );
not ( n279744 , n273783 );
not ( n279745 , n221271 );
or ( n279746 , n279744 , n279745 );
nor ( n279747 , n254201 , n37725 );
nand ( n279748 , n279746 , n279747 );
nand ( n279749 , n35431 , n37016 );
nand ( n279750 , n279743 , n279748 , n279749 );
buf ( n279751 , n279750 );
buf ( n279752 , n29209 );
buf ( n279753 , n40805 );
buf ( n279754 , n25952 );
buf ( n279755 , n38518 );
or ( n279756 , n271012 , n246237 );
not ( n279757 , n277321 );
nand ( n279758 , n271023 , n246237 );
not ( n279759 , n279758 );
and ( n279760 , n279757 , n279759 );
and ( n279761 , n244073 , n209153 );
nor ( n279762 , n279760 , n279761 );
nand ( n279763 , n246238 , n271022 );
nand ( n279764 , n279756 , n279762 , n279763 );
buf ( n279765 , n279764 );
buf ( n279766 , RI1753a460_587);
and ( n279767 , n27883 , n279766 );
buf ( n279768 , n279767 );
nor ( n279769 , n274669 , n55146 );
nand ( n279770 , n279769 , n252853 , n274681 );
not ( n279771 , n274670 );
not ( n279772 , n252853 );
or ( n279773 , n279771 , n279772 );
nor ( n279774 , n274681 , n234445 );
nand ( n279775 , n279773 , n279774 );
nand ( n279776 , n31577 , n216999 );
nand ( n279777 , n279770 , n279775 , n279776 );
buf ( n279778 , n279777 );
not ( n279779 , n40464 );
nand ( n279780 , n279779 , n254528 );
nand ( n279781 , n274981 , n274993 );
or ( n279782 , n279780 , n279781 );
not ( n279783 , n274981 );
not ( n279784 , n279779 );
or ( n279785 , n279783 , n279784 );
nor ( n279786 , n274993 , n252258 );
nand ( n279787 , n279785 , n279786 );
nand ( n279788 , n239240 , n42494 );
nand ( n279789 , n279782 , n279787 , n279788 );
buf ( n279790 , n279789 );
nand ( n279791 , n246175 , n259009 );
not ( n279792 , n245853 );
not ( n279793 , n39444 );
or ( n279794 , n279792 , n279793 );
not ( n279795 , n245853 );
nand ( n279796 , n279795 , n39434 );
nand ( n279797 , n279794 , n279796 );
and ( n279798 , n279797 , n250255 );
not ( n279799 , n279797 );
and ( n279800 , n279799 , n248795 );
nor ( n279801 , n279798 , n279800 );
not ( n279802 , n279801 );
nand ( n279803 , n279802 , n246209 );
or ( n279804 , n279791 , n279803 );
not ( n279805 , n246209 );
not ( n279806 , n246175 );
or ( n279807 , n279805 , n279806 );
nor ( n279808 , n279802 , n256413 );
nand ( n279809 , n279807 , n279808 );
nand ( n279810 , n31577 , n206887 );
nand ( n279811 , n279804 , n279809 , n279810 );
buf ( n279812 , n279811 );
nand ( n279813 , n275450 , n267249 );
not ( n279814 , n279813 );
not ( n279815 , n258709 );
or ( n279816 , n279814 , n279815 );
nor ( n279817 , n272237 , n272234 );
and ( n279818 , n279817 , n258708 );
not ( n279819 , n39767 );
nor ( n279820 , n279819 , n35244 );
nor ( n279821 , n279818 , n279820 );
nand ( n279822 , n279816 , n279821 );
buf ( n279823 , n279822 );
not ( n279824 , n28374 );
not ( n279825 , n37728 );
or ( n279826 , n279824 , n279825 );
nand ( n279827 , n255217 , n255205 );
and ( n279828 , n279827 , n271361 );
not ( n279829 , n279827 );
and ( n279830 , n279829 , n264483 );
nor ( n279831 , n279828 , n279830 );
or ( n279832 , n279831 , n254882 );
nand ( n279833 , n279826 , n279832 );
buf ( n279834 , n279833 );
not ( n279835 , n55733 );
nand ( n279836 , n261081 , n279577 );
or ( n279837 , n279835 , n279836 );
not ( n279838 , n279577 );
not ( n279839 , n55736 );
or ( n279840 , n279838 , n279839 );
nor ( n279841 , n261081 , n238635 );
nand ( n279842 , n279840 , n279841 );
nand ( n279843 , n253486 , n33409 );
nand ( n279844 , n279837 , n279842 , n279843 );
buf ( n279845 , n279844 );
or ( n279846 , n25328 , n279231 );
or ( n279847 , n25336 , n263188 );
nand ( n279848 , n279846 , n279847 );
buf ( n279849 , n279848 );
buf ( n279850 , n38184 );
not ( n279851 , n274960 );
nand ( n279852 , n267011 , n279851 );
or ( n279853 , n265034 , n279852 );
not ( n279854 , n267011 );
not ( n279855 , n265033 );
or ( n279856 , n279854 , n279855 );
nor ( n279857 , n279851 , n254882 );
nand ( n279858 , n279856 , n279857 );
nand ( n279859 , n35431 , n29827 );
nand ( n279860 , n279853 , n279858 , n279859 );
buf ( n279861 , n279860 );
not ( n279862 , n278197 );
nand ( n279863 , n279862 , n254528 );
nor ( n279864 , n268073 , n268099 );
or ( n279865 , n279863 , n279864 );
not ( n279866 , n268073 );
nand ( n279867 , n268100 , n278197 , n279866 );
nand ( n279868 , n246460 , n25396 );
nand ( n279869 , n279865 , n279867 , n279868 );
buf ( n279870 , n279869 );
not ( n279871 , n252317 );
not ( n279872 , n279871 );
buf ( n279873 , n243997 );
not ( n279874 , n279873 );
and ( n279875 , n279872 , n279874 );
and ( n279876 , n279871 , n279873 );
nor ( n279877 , n279875 , n279876 );
and ( n279878 , n279877 , n252327 );
not ( n279879 , n279877 );
and ( n279880 , n279879 , n252324 );
nor ( n279881 , n279878 , n279880 );
nand ( n279882 , n236768 , n279881 );
not ( n279883 , n236796 );
or ( n279884 , n279882 , n279883 );
nor ( n279885 , n236541 , n234818 );
nand ( n279886 , n279882 , n279885 );
nand ( n279887 , n234024 , n26183 );
nand ( n279888 , n279884 , n279886 , n279887 );
buf ( n279889 , n279888 );
not ( n279890 , n37908 );
not ( n279891 , n31577 );
or ( n279892 , n279890 , n279891 );
nand ( n279893 , n272691 , n272702 );
and ( n279894 , n279893 , n279709 );
not ( n279895 , n279893 );
and ( n279896 , n279895 , n279708 );
nor ( n279897 , n279894 , n279896 );
or ( n279898 , n279897 , n254882 );
nand ( n279899 , n279892 , n279898 );
buf ( n279900 , n279899 );
not ( n279901 , RI19a95de0_2641);
or ( n279902 , n25328 , n279901 );
not ( n279903 , RI19a8be08_2712);
or ( n279904 , n25335 , n279903 );
nand ( n279905 , n279902 , n279904 );
buf ( n279906 , n279905 );
not ( n279907 , RI19ac92a8_2261);
or ( n279908 , n25328 , n279907 );
or ( n279909 , n25335 , n264133 );
nand ( n279910 , n279908 , n279909 );
buf ( n279911 , n279910 );
buf ( n279912 , RI19ad1060_2204);
and ( n279913 , n25326 , n279912 );
buf ( n279914 , n279913 );
not ( n279915 , n278673 );
nand ( n279916 , n279915 , n256617 );
not ( n279917 , n256607 );
or ( n279918 , n279916 , n279917 );
nor ( n279919 , n256605 , n38637 );
nand ( n279920 , n279916 , n279919 );
nand ( n279921 , n39766 , n33194 );
nand ( n279922 , n279918 , n279920 , n279921 );
buf ( n279923 , n279922 );
not ( n279924 , n25994 );
not ( n279925 , n55760 );
or ( n279926 , n279924 , n279925 );
not ( n279927 , n265783 );
nand ( n279928 , n279927 , n265794 );
not ( n279929 , n249549 );
not ( n279930 , n255736 );
not ( n279931 , n279930 );
not ( n279932 , n256131 );
or ( n279933 , n279931 , n279932 );
nand ( n279934 , n256130 , n255736 );
nand ( n279935 , n279933 , n279934 );
not ( n279936 , n279935 );
and ( n279937 , n279929 , n279936 );
and ( n279938 , n249549 , n279935 );
nor ( n279939 , n279937 , n279938 );
not ( n279940 , n279939 );
and ( n279941 , n279928 , n279940 );
not ( n279942 , n279928 );
and ( n279943 , n279942 , n279939 );
nor ( n279944 , n279941 , n279943 );
or ( n279945 , n279944 , n257174 );
nand ( n279946 , n279926 , n279945 );
buf ( n279947 , n279946 );
or ( n279948 , n25328 , n274112 );
or ( n279949 , n25335 , n279907 );
nand ( n279950 , n279948 , n279949 );
buf ( n279951 , n279950 );
not ( n279952 , n41051 );
not ( n279953 , n255116 );
or ( n279954 , n279952 , n279953 );
nand ( n279955 , n253611 , n266741 );
not ( n279956 , n253681 );
and ( n279957 , n279955 , n279956 );
not ( n279958 , n279955 );
and ( n279959 , n279958 , n253681 );
nor ( n279960 , n279957 , n279959 );
or ( n279961 , n279960 , n251498 );
nand ( n279962 , n279954 , n279961 );
buf ( n279963 , n279962 );
not ( n279964 , n26138 );
not ( n279965 , n245701 );
or ( n279966 , n279964 , n279965 );
nand ( n279967 , n268668 , n271773 );
and ( n279968 , n279967 , n268691 );
not ( n279969 , n279967 );
and ( n279970 , n279969 , n268694 );
nor ( n279971 , n279968 , n279970 );
or ( n279972 , n279971 , n244217 );
nand ( n279973 , n279966 , n279972 );
buf ( n279974 , n279973 );
not ( n279975 , n46081 );
nand ( n279976 , n250377 , n250302 );
or ( n279977 , n279975 , n279976 );
not ( n279978 , n250302 );
not ( n279979 , n46077 );
not ( n279980 , n279979 );
or ( n279981 , n279978 , n279980 );
nor ( n279982 , n250377 , n50944 );
nand ( n279983 , n279981 , n279982 );
nand ( n279984 , n244484 , n33816 );
nand ( n279985 , n279977 , n279983 , n279984 );
buf ( n279986 , n279985 );
and ( n279987 , n248264 , n240316 );
not ( n279988 , n248264 );
and ( n279989 , n279988 , n240312 );
or ( n279990 , n279987 , n279989 );
and ( n279991 , n279990 , n240505 );
not ( n279992 , n279990 );
and ( n279993 , n279992 , n240508 );
nor ( n279994 , n279991 , n279993 );
nand ( n279995 , n279994 , n246177 );
not ( n279996 , n265641 );
nand ( n279997 , n265651 , n279996 );
or ( n279998 , n279995 , n279997 );
not ( n279999 , n279996 );
not ( n280000 , n279994 );
or ( n280001 , n279999 , n280000 );
nor ( n280002 , n265651 , n249531 );
nand ( n280003 , n280001 , n280002 );
nand ( n280004 , n41944 , n26168 );
nand ( n280005 , n279998 , n280003 , n280004 );
buf ( n280006 , n280005 );
not ( n280007 , n263119 );
nand ( n280008 , n275818 , n280007 );
not ( n280009 , n275824 );
or ( n280010 , n280008 , n280009 );
nor ( n280011 , n275807 , n244399 );
nand ( n280012 , n280008 , n280011 );
nand ( n280013 , n233501 , n33278 );
nand ( n280014 , n280010 , n280012 , n280013 );
buf ( n280015 , n280014 );
not ( n280016 , n252196 );
not ( n280017 , n252088 );
or ( n280018 , n280016 , n280017 );
not ( n280019 , n46468 );
not ( n280020 , n280019 );
not ( n280021 , n51597 );
or ( n280022 , n280020 , n280021 );
or ( n280023 , n51597 , n280019 );
nand ( n280024 , n280022 , n280023 );
and ( n280025 , n280024 , n253189 );
not ( n280026 , n280024 );
and ( n280027 , n280026 , n253197 );
nor ( n280028 , n280025 , n280027 );
nand ( n280029 , n280028 , n230207 );
not ( n280030 , n280029 );
nand ( n280031 , n280018 , n280030 );
not ( n280032 , n252089 );
nor ( n280033 , n280028 , n252197 );
nand ( n280034 , n280032 , n280033 );
nand ( n280035 , n239240 , n204910 );
nand ( n280036 , n280031 , n280034 , n280035 );
buf ( n280037 , n280036 );
buf ( n280038 , n38029 );
buf ( n280039 , n28659 );
buf ( n280040 , n204299 );
not ( n280041 , n272255 );
not ( n280042 , n38940 );
not ( n280043 , n251313 );
or ( n280044 , n280042 , n280043 );
or ( n280045 , n251313 , n38940 );
nand ( n280046 , n280044 , n280045 );
and ( n280047 , n280046 , n256008 );
not ( n280048 , n280046 );
and ( n280049 , n280048 , n256012 );
nor ( n280050 , n280047 , n280049 );
nand ( n280051 , n280041 , n280050 );
nor ( n280052 , n271052 , n37725 );
not ( n280053 , n280052 );
or ( n280054 , n280051 , n280053 );
nand ( n280055 , n280051 , n271054 );
nand ( n280056 , n255116 , n28231 );
nand ( n280057 , n280054 , n280055 , n280056 );
buf ( n280058 , n280057 );
nand ( n280059 , n247211 , n271417 );
or ( n280060 , n260326 , n280059 );
not ( n280061 , n247198 );
not ( n280062 , n247211 );
or ( n280063 , n280061 , n280062 );
nor ( n280064 , n271417 , n40465 );
nand ( n280065 , n280063 , n280064 );
nand ( n280066 , n239240 , n31452 );
nand ( n280067 , n280060 , n280065 , n280066 );
buf ( n280068 , n280067 );
not ( n280069 , n269683 );
not ( n280070 , n280069 );
not ( n280071 , n269677 );
or ( n280072 , n280070 , n280071 );
nand ( n280073 , n280072 , n261039 );
and ( n280074 , n278150 , n265719 , n265721 );
and ( n280075 , n33102 , n35431 );
nor ( n280076 , n280074 , n280075 );
nand ( n280077 , n280073 , n280076 );
buf ( n280078 , n280077 );
nor ( n280079 , n50037 , n256481 );
not ( n280080 , n248313 );
not ( n280081 , n246321 );
or ( n280082 , n280080 , n280081 );
not ( n280083 , n248313 );
nand ( n280084 , n280083 , n246326 );
nand ( n280085 , n280082 , n280084 );
and ( n280086 , n280085 , n254483 );
not ( n280087 , n280085 );
and ( n280088 , n280087 , n246331 );
nor ( n280089 , n280086 , n280088 );
nand ( n280090 , n280079 , n280089 , n50485 );
not ( n280091 , n50037 );
not ( n280092 , n280091 );
not ( n280093 , n280089 );
or ( n280094 , n280092 , n280093 );
nand ( n280095 , n280094 , n270385 );
nand ( n280096 , n237361 , n205253 );
nand ( n280097 , n280090 , n280095 , n280096 );
buf ( n280098 , n280097 );
or ( n280099 , n233507 , n273080 );
or ( n280100 , n25336 , n272003 );
nand ( n280101 , n280099 , n280100 );
buf ( n280102 , n280101 );
buf ( n280103 , n29319 );
buf ( n280104 , n30241 );
buf ( n280105 , n34723 );
buf ( n280106 , n26095 );
or ( n280107 , n25328 , n279221 );
not ( n280108 , RI19abf2d0_2339);
or ( n280109 , n25336 , n280108 );
nand ( n280110 , n280107 , n280109 );
buf ( n280111 , n280110 );
not ( n280112 , n249008 );
nand ( n280113 , n280112 , n50945 );
not ( n280114 , n280113 );
not ( n280115 , n244392 );
nand ( n280116 , n280115 , n249024 );
not ( n280117 , n280116 );
and ( n280118 , n280114 , n280117 );
and ( n280119 , n244073 , n34321 );
nor ( n280120 , n280118 , n280119 );
not ( n280121 , n249010 );
nand ( n280122 , n280121 , n244392 );
not ( n280123 , n244394 );
nand ( n280124 , n280123 , n249023 );
nand ( n280125 , n280120 , n280122 , n280124 );
buf ( n280126 , n280125 );
not ( n280127 , n268329 );
nand ( n280128 , n280127 , n241459 );
not ( n280129 , n237868 );
not ( n280130 , n44583 );
not ( n280131 , n280130 );
not ( n280132 , n237810 );
or ( n280133 , n280131 , n280132 );
nand ( n280134 , n237817 , n44583 );
nand ( n280135 , n280133 , n280134 );
not ( n280136 , n280135 );
or ( n280137 , n280129 , n280136 );
or ( n280138 , n280135 , n237868 );
nand ( n280139 , n280137 , n280138 );
not ( n280140 , n280139 );
nand ( n280141 , n268318 , n280140 );
or ( n280142 , n280128 , n280141 );
not ( n280143 , n268318 );
not ( n280144 , n280127 );
or ( n280145 , n280143 , n280144 );
nor ( n280146 , n280140 , n253213 );
nand ( n280147 , n280145 , n280146 );
nand ( n280148 , n31577 , n32298 );
nand ( n280149 , n280142 , n280147 , n280148 );
buf ( n280150 , n280149 );
not ( n280151 , n271298 );
not ( n280152 , n259781 );
or ( n280153 , n280151 , n280152 );
nand ( n280154 , n280153 , n226010 );
or ( n280155 , n280154 , n259785 );
nand ( n280156 , n259781 , n276481 , n259785 );
nand ( n280157 , n236798 , n31686 );
nand ( n280158 , n280155 , n280156 , n280157 );
buf ( n280159 , n280158 );
or ( n280160 , n25328 , n250977 );
not ( n280161 , RI19aa24a0_2550);
or ( n280162 , n25336 , n280161 );
nand ( n280163 , n280160 , n280162 );
buf ( n280164 , n280163 );
not ( n280165 , n252089 );
not ( n280166 , n280029 );
or ( n280167 , n280165 , n280166 );
not ( n280168 , n243772 );
not ( n280169 , n258257 );
or ( n280170 , n280168 , n280169 );
not ( n280171 , n243772 );
nand ( n280172 , n280171 , n246028 );
nand ( n280173 , n280170 , n280172 );
and ( n280174 , n280173 , n260422 );
not ( n280175 , n280173 );
and ( n280176 , n280175 , n246065 );
nor ( n280177 , n280174 , n280176 );
nand ( n280178 , n280167 , n280177 );
nor ( n280179 , n280028 , n280177 );
and ( n280180 , n252201 , n280179 );
and ( n280181 , n245702 , n33968 );
nor ( n280182 , n280180 , n280181 );
nand ( n280183 , n280178 , n280182 );
buf ( n280184 , n280183 );
nand ( n280185 , n265457 , n279555 );
not ( n280186 , n279544 );
or ( n280187 , n280185 , n280186 );
nor ( n280188 , n279558 , n37725 );
nand ( n280189 , n280185 , n280188 );
nand ( n280190 , n35431 , n31592 );
nand ( n280191 , n280187 , n280189 , n280190 );
buf ( n280192 , n280191 );
not ( n280193 , n240667 );
not ( n280194 , n247393 );
or ( n280195 , n280193 , n280194 );
not ( n280196 , n240667 );
nand ( n280197 , n280196 , n247399 );
nand ( n280198 , n280195 , n280197 );
and ( n280199 , n280198 , n267358 );
not ( n280200 , n280198 );
and ( n280201 , n280200 , n247349 );
nor ( n280202 , n280199 , n280201 );
not ( n280203 , n280202 );
nand ( n280204 , n280203 , n270783 );
or ( n280205 , n278902 , n280204 );
nand ( n280206 , n278897 , n280204 );
nand ( n280207 , n245221 , n31186 );
nand ( n280208 , n280205 , n280206 , n280207 );
buf ( n280209 , n280208 );
not ( n280210 , n54501 );
not ( n280211 , n237361 );
or ( n280212 , n280210 , n280211 );
not ( n280213 , n246198 );
not ( n280214 , n44169 );
not ( n280215 , n54325 );
or ( n280216 , n280214 , n280215 );
not ( n280217 , n44169 );
nand ( n280218 , n280217 , n255320 );
nand ( n280219 , n280216 , n280218 );
and ( n280220 , n280219 , n234098 );
not ( n280221 , n280219 );
and ( n280222 , n280221 , n234107 );
nor ( n280223 , n280220 , n280222 );
nand ( n280224 , n279801 , n280223 );
not ( n280225 , n280224 );
and ( n280226 , n280213 , n280225 );
and ( n280227 , n280224 , n246198 );
nor ( n280228 , n280226 , n280227 );
or ( n280229 , n280228 , n257851 );
nand ( n280230 , n280212 , n280229 );
buf ( n280231 , n280230 );
nand ( n280232 , n267804 , n269053 );
nand ( n280233 , n255165 , n258918 );
or ( n280234 , n280232 , n280233 );
not ( n280235 , n255165 );
not ( n280236 , n267804 );
or ( n280237 , n280235 , n280236 );
nor ( n280238 , n269053 , n221279 );
nand ( n280239 , n280237 , n280238 );
nand ( n280240 , n39766 , n37737 );
nand ( n280241 , n280234 , n280239 , n280240 );
buf ( n280242 , n280241 );
not ( n280243 , n33387 );
not ( n280244 , n245943 );
or ( n280245 , n280243 , n280244 );
not ( n280246 , n246663 );
nand ( n280247 , n280246 , n260141 );
and ( n280248 , n280247 , n246481 );
not ( n280249 , n280247 );
not ( n280250 , n246481 );
and ( n280251 , n280249 , n280250 );
nor ( n280252 , n280248 , n280251 );
or ( n280253 , n280252 , n258327 );
nand ( n280254 , n280245 , n280253 );
buf ( n280255 , n280254 );
or ( n280256 , n25328 , n272665 );
or ( n280257 , n226822 , n263258 );
nand ( n280258 , n280256 , n280257 );
buf ( n280259 , n280258 );
nand ( n280260 , n257599 , n267700 );
nor ( n280261 , n264826 , n55108 );
not ( n280262 , n280261 );
or ( n280263 , n280260 , n280262 );
nand ( n280264 , n280260 , n264828 );
nand ( n280265 , n255116 , n32029 );
nand ( n280266 , n280263 , n280264 , n280265 );
buf ( n280267 , n280266 );
or ( n280268 , n25328 , n251104 );
or ( n280269 , n25336 , n279901 );
nand ( n280270 , n280268 , n280269 );
buf ( n280271 , n280270 );
not ( n280272 , n33975 );
not ( n280273 , n245943 );
or ( n280274 , n280272 , n280273 );
nand ( n280275 , n253030 , n255035 );
not ( n280276 , n255046 );
and ( n280277 , n280275 , n280276 );
not ( n280278 , n280275 );
and ( n280279 , n280278 , n255046 );
nor ( n280280 , n280277 , n280279 );
or ( n280281 , n280280 , n258179 );
nand ( n280282 , n280274 , n280281 );
buf ( n280283 , n280282 );
not ( n280284 , n266441 );
nand ( n280285 , n264603 , n264629 );
or ( n280286 , n280284 , n280285 );
not ( n280287 , n264603 );
not ( n280288 , n266436 );
or ( n280289 , n280287 , n280288 );
nor ( n280290 , n264629 , n49051 );
nand ( n280291 , n280289 , n280290 );
nand ( n280292 , n245701 , n210628 );
nand ( n280293 , n280286 , n280291 , n280292 );
buf ( n280294 , n280293 );
or ( n280295 , n25328 , n269224 );
or ( n280296 , n25335 , n270927 );
nand ( n280297 , n280295 , n280296 );
buf ( n280298 , n280297 );
not ( n280299 , n240745 );
not ( n280300 , n247348 );
or ( n280301 , n280299 , n280300 );
not ( n280302 , n240745 );
nand ( n280303 , n280302 , n263230 );
nand ( n280304 , n280301 , n280303 );
and ( n280305 , n280304 , n263235 );
not ( n280306 , n280304 );
and ( n280307 , n280306 , n257952 );
nor ( n280308 , n280305 , n280307 );
not ( n280309 , n280308 );
not ( n280310 , n240299 );
not ( n280311 , n252051 );
or ( n280312 , n280310 , n280311 );
not ( n280313 , n240299 );
nand ( n280314 , n280313 , n252036 );
nand ( n280315 , n280312 , n280314 );
and ( n280316 , n280315 , n252644 );
not ( n280317 , n280315 );
and ( n280318 , n280317 , n256227 );
nor ( n280319 , n280316 , n280318 );
nand ( n280320 , n280309 , n280319 );
buf ( n280321 , n49097 );
not ( n280322 , n280321 );
not ( n280323 , n45506 );
or ( n280324 , n280322 , n280323 );
or ( n280325 , n243426 , n280321 );
nand ( n280326 , n280324 , n280325 );
not ( n280327 , n280326 );
not ( n280328 , n45727 );
and ( n280329 , n280327 , n280328 );
and ( n280330 , n280326 , n45728 );
nor ( n280331 , n280329 , n280330 );
not ( n280332 , n280331 );
nor ( n280333 , n280332 , n234440 );
not ( n280334 , n280333 );
or ( n280335 , n280320 , n280334 );
nor ( n280336 , n280331 , n236795 );
nand ( n280337 , n280336 , n280320 );
nand ( n280338 , n46083 , n29034 );
nand ( n280339 , n280335 , n280337 , n280338 );
buf ( n280340 , n280339 );
nor ( n280341 , n241703 , n261742 );
nand ( n280342 , n267100 , n280341 );
not ( n280343 , n261739 );
not ( n280344 , n267096 );
not ( n280345 , n280344 );
or ( n280346 , n280343 , n280345 );
nor ( n280347 , n276968 , n234021 );
nand ( n280348 , n280346 , n280347 );
nand ( n280349 , n237714 , n30006 );
nand ( n280350 , n280342 , n280348 , n280349 );
buf ( n280351 , n280350 );
not ( n280352 , RI1754ba58_27);
or ( n280353 , n229127 , n280352 );
or ( n280354 , n25335 , n272663 );
nand ( n280355 , n280353 , n280354 );
buf ( n280356 , n280355 );
not ( n280357 , n250899 );
not ( n280358 , n50835 );
not ( n280359 , n263897 );
or ( n280360 , n280358 , n280359 );
or ( n280361 , n256494 , n50835 );
nand ( n280362 , n280360 , n280361 );
not ( n280363 , n280362 );
or ( n280364 , n280357 , n280363 );
or ( n280365 , n280362 , n263900 );
nand ( n280366 , n280364 , n280365 );
not ( n280367 , n280366 );
nand ( n280368 , n280367 , n264011 );
not ( n280369 , n269243 );
nand ( n280370 , n280369 , n241459 );
or ( n280371 , n280368 , n280370 );
nor ( n280372 , n280369 , n33254 );
nand ( n280373 , n280372 , n280368 );
nand ( n280374 , n247744 , n36805 );
nand ( n280375 , n280371 , n280373 , n280374 );
buf ( n280376 , n280375 );
not ( n280377 , n256163 );
nand ( n280378 , n257236 , n257245 );
or ( n280379 , n280377 , n280378 );
not ( n280380 , n257245 );
not ( n280381 , n256141 );
or ( n280382 , n280380 , n280381 );
nor ( n280383 , n257236 , n43968 );
nand ( n280384 , n280382 , n280383 );
nand ( n280385 , n35431 , n40710 );
nand ( n280386 , n280379 , n280384 , n280385 );
buf ( n280387 , n280386 );
buf ( n280388 , n28990 );
buf ( n280389 , n39635 );
buf ( n280390 , n31301 );
buf ( n280391 , n237478 );
not ( n280392 , n280391 );
not ( n280393 , n263562 );
or ( n280394 , n280392 , n280393 );
or ( n280395 , n263562 , n280391 );
nand ( n280396 , n280394 , n280395 );
xnor ( n280397 , n280396 , n249285 );
nand ( n280398 , n280397 , n250111 );
not ( n280399 , n271742 );
nand ( n280400 , n271731 , n280399 );
or ( n280401 , n280398 , n280400 );
not ( n280402 , n280399 );
not ( n280403 , n280397 );
or ( n280404 , n280402 , n280403 );
nor ( n280405 , n271731 , n254150 );
nand ( n280406 , n280404 , n280405 );
nand ( n280407 , n244987 , n33397 );
nand ( n280408 , n280401 , n280406 , n280407 );
buf ( n280409 , n280408 );
nand ( n280410 , n267064 , n267074 );
or ( n280411 , n265999 , n280410 );
not ( n280412 , n267074 );
not ( n280413 , n265991 );
or ( n280414 , n280412 , n280413 );
nor ( n280415 , n267064 , n52445 );
nand ( n280416 , n280414 , n280415 );
nand ( n280417 , n37728 , n28573 );
nand ( n280418 , n280411 , n280416 , n280417 );
buf ( n280419 , n280418 );
nand ( n280420 , n258963 , n273401 );
or ( n280421 , n275171 , n280420 );
not ( n280422 , n273401 );
not ( n280423 , n273389 );
or ( n280424 , n280422 , n280423 );
nand ( n280425 , n280424 , n258964 );
nand ( n280426 , n234024 , n37867 );
nand ( n280427 , n280421 , n280425 , n280426 );
buf ( n280428 , n280427 );
not ( n280429 , RI19aa0970_2564);
or ( n280430 , n226819 , n280429 );
or ( n280431 , n25335 , n277915 );
nand ( n280432 , n280430 , n280431 );
buf ( n280433 , n280432 );
buf ( n280434 , n42272 );
buf ( n280435 , n30836 );
not ( n280436 , n31732 );
not ( n280437 , n51381 );
or ( n280438 , n280436 , n280437 );
not ( n280439 , n252781 );
not ( n280440 , n50940 );
or ( n280441 , n280439 , n280440 );
not ( n280442 , n252781 );
nand ( n280443 , n280442 , n50930 );
nand ( n280444 , n280441 , n280443 );
and ( n280445 , n280444 , n244529 );
not ( n280446 , n280444 );
and ( n280447 , n280446 , n244532 );
nor ( n280448 , n280445 , n280447 );
not ( n280449 , n280448 );
nand ( n280450 , n280449 , n267779 );
not ( n280451 , n244586 );
not ( n280452 , n236335 );
not ( n280453 , n244583 );
or ( n280454 , n280452 , n280453 );
or ( n280455 , n255121 , n236335 );
nand ( n280456 , n280454 , n280455 );
not ( n280457 , n280456 );
and ( n280458 , n280451 , n280457 );
and ( n280459 , n244591 , n280456 );
nor ( n280460 , n280458 , n280459 );
not ( n280461 , n280460 );
and ( n280462 , n280450 , n280461 );
not ( n280463 , n280450 );
and ( n280464 , n280463 , n280460 );
nor ( n280465 , n280462 , n280464 );
or ( n280466 , n280465 , n255533 );
nand ( n280467 , n280438 , n280466 );
buf ( n280468 , n280467 );
nand ( n280469 , n269296 , n277047 );
nand ( n280470 , n277044 , n241459 );
or ( n280471 , n280469 , n280470 );
not ( n280472 , n277044 );
not ( n280473 , n269296 );
or ( n280474 , n280472 , n280473 );
nor ( n280475 , n277047 , n243204 );
nand ( n280476 , n280474 , n280475 );
nand ( n280477 , n31577 , n29100 );
nand ( n280478 , n280471 , n280476 , n280477 );
buf ( n280479 , n280478 );
buf ( n280480 , n37552 );
not ( n280481 , n35512 );
not ( n280482 , n258213 );
or ( n280483 , n280481 , n280482 );
not ( n280484 , n278176 );
nand ( n280485 , n273598 , n280484 );
and ( n280486 , n280485 , n257735 );
not ( n280487 , n280485 );
and ( n280488 , n280487 , n257734 );
nor ( n280489 , n280486 , n280488 );
or ( n280490 , n280489 , n255707 );
nand ( n280491 , n280483 , n280490 );
buf ( n280492 , n280491 );
nand ( n280493 , n275356 , n222532 );
nand ( n280494 , n275369 , n259533 );
or ( n280495 , n280493 , n280494 );
not ( n280496 , n275369 );
not ( n280497 , n275356 );
or ( n280498 , n280496 , n280497 );
nand ( n280499 , n280498 , n259534 );
nand ( n280500 , n247744 , n26479 );
nand ( n280501 , n280495 , n280499 , n280500 );
buf ( n280502 , n280501 );
not ( n280503 , n246198 );
not ( n280504 , n280223 );
nand ( n280505 , n280503 , n280504 );
or ( n280506 , n280505 , n246178 );
nor ( n280507 , n246176 , n233972 );
nand ( n280508 , n280507 , n280505 );
nand ( n280509 , n255116 , n40702 );
nand ( n280510 , n280506 , n280508 , n280509 );
buf ( n280511 , n280510 );
not ( n280512 , n40834 );
not ( n280513 , n245701 );
or ( n280514 , n280512 , n280513 );
not ( n280515 , n245348 );
not ( n280516 , n235357 );
or ( n280517 , n280515 , n280516 );
not ( n280518 , n245348 );
nand ( n280519 , n280518 , n235366 );
nand ( n280520 , n280517 , n280519 );
and ( n280521 , n280520 , n235372 );
not ( n280522 , n280520 );
and ( n280523 , n280522 , n235369 );
nor ( n280524 , n280521 , n280523 );
not ( n280525 , n280524 );
nand ( n280526 , n280525 , n262179 );
and ( n280527 , n280526 , n267230 );
not ( n280528 , n280526 );
not ( n280529 , n267230 );
and ( n280530 , n280528 , n280529 );
nor ( n280531 , n280527 , n280530 );
or ( n280532 , n280531 , n254882 );
nand ( n280533 , n280514 , n280532 );
buf ( n280534 , n280533 );
not ( n280535 , n262496 );
nand ( n280536 , n262500 , n280535 );
or ( n280537 , n244810 , n280536 );
not ( n280538 , n244807 );
nor ( n280539 , n280538 , n249531 );
nand ( n280540 , n280539 , n280536 );
nand ( n280541 , n39766 , n28567 );
nand ( n280542 , n280537 , n280540 , n280541 );
buf ( n280543 , n280542 );
not ( n280544 , n267012 );
nand ( n280545 , n265044 , n279851 );
or ( n280546 , n280544 , n280545 );
not ( n280547 , n279851 );
not ( n280548 , n267003 );
or ( n280549 , n280547 , n280548 );
nor ( n280550 , n265044 , n236795 );
nand ( n280551 , n280549 , n280550 );
nand ( n280552 , n39767 , n35535 );
nand ( n280553 , n280546 , n280551 , n280552 );
buf ( n280554 , n280553 );
not ( n280555 , n277132 );
not ( n280556 , n270578 );
or ( n280557 , n280555 , n280556 );
nor ( n280558 , n270591 , n50944 );
nand ( n280559 , n280557 , n280558 );
nand ( n280560 , n277137 , n270591 , n270578 );
nand ( n280561 , n31577 , n217071 );
nand ( n280562 , n280559 , n280560 , n280561 );
buf ( n280563 , n280562 );
buf ( n280564 , n45301 );
or ( n280565 , n25328 , n263260 );
not ( n280566 , RI19ab4740_2420);
or ( n280567 , n25335 , n280566 );
nand ( n280568 , n280565 , n280567 );
buf ( n280569 , n280568 );
nand ( n280570 , n259220 , n274311 );
not ( n280571 , n206859 );
not ( n280572 , n256711 );
or ( n280573 , n280571 , n280572 );
not ( n280574 , n206859 );
nand ( n280575 , n280574 , n253009 );
nand ( n280576 , n280573 , n280575 );
and ( n280577 , n280576 , n253015 );
not ( n280578 , n280576 );
and ( n280579 , n280578 , n263207 );
nor ( n280580 , n280577 , n280579 );
nand ( n280581 , n280580 , n259230 );
or ( n280582 , n280570 , n280581 );
not ( n280583 , n259230 );
not ( n280584 , n259220 );
or ( n280585 , n280583 , n280584 );
nor ( n280586 , n280580 , n233971 );
nand ( n280587 , n280585 , n280586 );
nand ( n280588 , n49054 , n30116 );
nand ( n280589 , n280582 , n280587 , n280588 );
buf ( n280590 , n280589 );
buf ( n280591 , n35919 );
not ( n280592 , n267362 );
nand ( n280593 , n280592 , n274326 );
not ( n280594 , n262388 );
or ( n280595 , n280593 , n280594 );
nand ( n280596 , n262381 , n274326 );
nand ( n280597 , n280596 , n267362 , n241459 );
nand ( n280598 , n238638 , n34352 );
nand ( n280599 , n280595 , n280597 , n280598 );
buf ( n280600 , n280599 );
nor ( n280601 , n250582 , n235895 );
nor ( n280602 , n275136 , n250592 );
nand ( n280603 , n280601 , n280602 );
not ( n280604 , n250593 );
not ( n280605 , n250582 );
not ( n280606 , n280605 );
or ( n280607 , n280604 , n280606 );
nor ( n280608 , n275135 , n252258 );
nand ( n280609 , n280607 , n280608 );
nand ( n280610 , n41945 , n29639 );
nand ( n280611 , n280603 , n280609 , n280610 );
buf ( n280612 , n280611 );
not ( n280613 , n279994 );
nor ( n280614 , n280613 , n238635 );
not ( n280615 , n245462 );
not ( n280616 , n250439 );
or ( n280617 , n280615 , n280616 );
or ( n280618 , n261036 , n245462 );
nand ( n280619 , n280617 , n280618 );
not ( n280620 , n280619 );
not ( n280621 , n250501 );
and ( n280622 , n280620 , n280621 );
and ( n280623 , n280619 , n250501 );
nor ( n280624 , n280622 , n280623 );
nand ( n280625 , n280624 , n265629 );
nand ( n280626 , n280614 , n280625 );
not ( n280627 , n280624 );
nor ( n280628 , n280627 , n53680 );
nor ( n280629 , n279994 , n265628 );
nand ( n280630 , n280628 , n280629 );
nand ( n280631 , n256292 , n35350 );
nand ( n280632 , n280626 , n280630 , n280631 );
buf ( n280633 , n280632 );
not ( n280634 , n226260 );
not ( n280635 , n280634 );
not ( n280636 , n262629 );
or ( n280637 , n280635 , n280636 );
not ( n280638 , n262628 );
or ( n280639 , n280638 , n280634 );
nand ( n280640 , n280637 , n280639 );
and ( n280641 , n280640 , n262633 );
not ( n280642 , n280640 );
and ( n280643 , n280642 , n263297 );
nor ( n280644 , n280641 , n280643 );
not ( n280645 , n280644 );
nand ( n280646 , n280645 , n205649 );
not ( n280647 , n263479 );
not ( n280648 , n235798 );
not ( n280649 , n245738 );
or ( n280650 , n280648 , n280649 );
not ( n280651 , n235798 );
nand ( n280652 , n280651 , n245743 );
nand ( n280653 , n280650 , n280652 );
and ( n280654 , n280653 , n245794 );
not ( n280655 , n280653 );
and ( n280656 , n280655 , n245799 );
nor ( n280657 , n280654 , n280656 );
not ( n280658 , n280657 );
nand ( n280659 , n280647 , n280658 );
or ( n280660 , n280646 , n280659 );
not ( n280661 , n280658 );
not ( n280662 , n280645 );
or ( n280663 , n280661 , n280662 );
nor ( n280664 , n280647 , n27889 );
nand ( n280665 , n280663 , n280664 );
nand ( n280666 , n234024 , n30929 );
nand ( n280667 , n280660 , n280665 , n280666 );
buf ( n280668 , n280667 );
not ( n280669 , n29788 );
not ( n280670 , n37728 );
or ( n280671 , n280669 , n280670 );
nand ( n280672 , n251909 , n251906 );
not ( n280673 , n259693 );
and ( n280674 , n280672 , n280673 );
not ( n280675 , n280672 );
and ( n280676 , n280675 , n259693 );
nor ( n280677 , n280674 , n280676 );
or ( n280678 , n280677 , n261009 );
nand ( n280679 , n280671 , n280678 );
buf ( n280680 , n280679 );
not ( n280681 , n33080 );
not ( n280682 , n245221 );
or ( n280683 , n280681 , n280682 );
not ( n280684 , n264023 );
nand ( n280685 , n280684 , n264012 );
and ( n280686 , n280685 , n280366 );
not ( n280687 , n280685 );
not ( n280688 , n280366 );
and ( n280689 , n280687 , n280688 );
nor ( n280690 , n280686 , n280689 );
or ( n280691 , n280690 , n252859 );
nand ( n280692 , n280683 , n280691 );
buf ( n280693 , n280692 );
nand ( n280694 , n256911 , n269702 );
or ( n280695 , n258207 , n280694 );
not ( n280696 , n256911 );
not ( n280697 , n258205 );
or ( n280698 , n280696 , n280697 );
nand ( n280699 , n280698 , n270620 );
nand ( n280700 , n250916 , n237050 );
nand ( n280701 , n280695 , n280699 , n280700 );
buf ( n280702 , n280701 );
not ( n280703 , n31495 );
not ( n280704 , n249131 );
or ( n280705 , n280703 , n280704 );
not ( n280706 , RI1754c340_8);
or ( n280707 , n244611 , n280706 );
nand ( n280708 , n280705 , n280707 );
buf ( n280709 , n280708 );
not ( n280710 , n29558 );
not ( n280711 , n257764 );
or ( n280712 , n280710 , n280711 );
nand ( n280713 , n269393 , n269404 );
and ( n280714 , n280713 , n260055 );
not ( n280715 , n280713 );
and ( n280716 , n280715 , n260416 );
nor ( n280717 , n280714 , n280716 );
or ( n280718 , n280717 , n49959 );
nand ( n280719 , n280712 , n280718 );
buf ( n280720 , n280719 );
or ( n280721 , n25328 , n271707 );
or ( n280722 , n25335 , n258906 );
nand ( n280723 , n280721 , n280722 );
buf ( n280724 , n280723 );
or ( n280725 , n25328 , n260907 );
not ( n280726 , RI19ac7958_2273);
or ( n280727 , n25335 , n280726 );
nand ( n280728 , n280725 , n280727 );
buf ( n280729 , n280728 );
nand ( n280730 , n273166 , n37717 );
or ( n280731 , n269215 , n280730 );
not ( n280732 , n37717 );
not ( n280733 , n269214 );
or ( n280734 , n280732 , n280733 );
nor ( n280735 , n273166 , n37725 );
nand ( n280736 , n280734 , n280735 );
nand ( n280737 , n246217 , n30397 );
nand ( n280738 , n280731 , n280736 , n280737 );
buf ( n280739 , n280738 );
not ( n280740 , n257887 );
nand ( n280741 , n280740 , n230207 );
nand ( n280742 , n257900 , n270558 );
or ( n280743 , n280741 , n280742 );
not ( n280744 , n270558 );
not ( n280745 , n280740 );
or ( n280746 , n280744 , n280745 );
nor ( n280747 , n257900 , n237384 );
nand ( n280748 , n280746 , n280747 );
nand ( n280749 , n31577 , n25546 );
nand ( n280750 , n280743 , n280748 , n280749 );
buf ( n280751 , n280750 );
not ( n280752 , n247177 );
not ( n280753 , n253474 );
or ( n280754 , n280752 , n280753 );
not ( n280755 , n247177 );
nand ( n280756 , n280755 , n248276 );
nand ( n280757 , n280754 , n280756 );
and ( n280758 , n280757 , n248284 );
not ( n280759 , n280757 );
and ( n280760 , n280759 , n248281 );
nor ( n280761 , n280758 , n280760 );
nor ( n280762 , n280761 , n52445 );
nor ( n280763 , n236769 , n279881 );
nand ( n280764 , n280762 , n280763 );
not ( n280765 , n280761 );
not ( n280766 , n279881 );
nand ( n280767 , n280765 , n280766 );
nand ( n280768 , n280767 , n236769 , n40466 );
nand ( n280769 , n48251 , n36500 );
nand ( n280770 , n280764 , n280768 , n280769 );
buf ( n280771 , n280770 );
not ( n280772 , RI19a9f368_2575);
or ( n280773 , n25328 , n280772 );
not ( n280774 , RI19a954f8_2645);
or ( n280775 , n25335 , n280774 );
nand ( n280776 , n280773 , n280775 );
buf ( n280777 , n280776 );
not ( n280778 , n278863 );
nand ( n280779 , n280778 , n278852 );
or ( n280780 , n260497 , n280779 );
nor ( n280781 , n260496 , n252872 );
nand ( n280782 , n280781 , n280779 );
nand ( n280783 , n55760 , n36655 );
nand ( n280784 , n280780 , n280782 , n280783 );
buf ( n280785 , n280784 );
buf ( n280786 , n38365 );
buf ( n280787 , n35907 );
buf ( n280788 , n29802 );
not ( n280789 , n26358 );
not ( n280790 , n51381 );
or ( n280791 , n280789 , n280790 );
not ( n280792 , n247325 );
not ( n280793 , n246165 );
or ( n280794 , n280792 , n280793 );
or ( n280795 , n246166 , n247325 );
nand ( n280796 , n280794 , n280795 );
not ( n280797 , n280796 );
not ( n280798 , n250682 );
and ( n280799 , n280797 , n280798 );
and ( n280800 , n280796 , n250682 );
nor ( n280801 , n280799 , n280800 );
nand ( n280802 , n280801 , n277388 );
and ( n280803 , n280802 , n276920 );
not ( n280804 , n280802 );
not ( n280805 , n276920 );
and ( n280806 , n280804 , n280805 );
nor ( n280807 , n280803 , n280806 );
or ( n280808 , n280807 , n258327 );
nand ( n280809 , n280791 , n280808 );
buf ( n280810 , n280809 );
or ( n280811 , n25328 , n270792 );
not ( n280812 , RI19abfa50_2335);
or ( n280813 , n25336 , n280812 );
nand ( n280814 , n280811 , n280813 );
buf ( n280815 , n280814 );
or ( n280816 , n25328 , n261224 );
or ( n280817 , n25335 , n278573 );
nand ( n280818 , n280816 , n280817 );
buf ( n280819 , n280818 );
or ( n280820 , n25328 , n270929 );
not ( n280821 , RI19a8a2d8_2723);
or ( n280822 , n25335 , n280821 );
nand ( n280823 , n280820 , n280822 );
buf ( n280824 , n280823 );
not ( n280825 , RI1754aa68_61);
or ( n280826 , n249125 , n280825 );
or ( n280827 , n25335 , n271535 );
nand ( n280828 , n280826 , n280827 );
buf ( n280829 , n280828 );
nand ( n280830 , n264861 , n258825 );
or ( n280831 , n272627 , n280830 );
nor ( n280832 , n272626 , n235050 );
nand ( n280833 , n280832 , n280830 );
nand ( n280834 , n255116 , n26225 );
nand ( n280835 , n280831 , n280833 , n280834 );
buf ( n280836 , n280835 );
nand ( n280837 , n268502 , n270273 );
or ( n280838 , n268474 , n280837 );
nand ( n280839 , n268473 , n270273 );
nand ( n280840 , n280839 , n268497 , n254227 );
nand ( n280841 , n35431 , n32938 );
nand ( n280842 , n280838 , n280840 , n280841 );
buf ( n280843 , n280842 );
not ( n280844 , n275331 );
nand ( n280845 , n264884 , n272854 );
or ( n280846 , n280844 , n280845 );
not ( n280847 , n272854 );
not ( n280848 , n272851 );
not ( n280849 , n280848 );
or ( n280850 , n280847 , n280849 );
nor ( n280851 , n264884 , n247212 );
nand ( n280852 , n280850 , n280851 );
nand ( n280853 , n251712 , n32591 );
nand ( n280854 , n280846 , n280852 , n280853 );
buf ( n280855 , n280854 );
not ( n280856 , n266691 );
nand ( n280857 , n280856 , n233973 );
nand ( n280858 , n266504 , n266705 );
or ( n280859 , n280857 , n280858 );
not ( n280860 , n266705 );
not ( n280861 , n280856 );
or ( n280862 , n280860 , n280861 );
nand ( n280863 , n280862 , n269261 );
nand ( n280864 , n238114 , n42459 );
nand ( n280865 , n280859 , n280863 , n280864 );
buf ( n280866 , n280865 );
or ( n280867 , n25328 , n272651 );
or ( n280868 , n226822 , n273692 );
nand ( n280869 , n280867 , n280868 );
buf ( n280870 , n280869 );
or ( n280871 , n25328 , n266582 );
or ( n280872 , n25335 , n275619 );
nand ( n280873 , n280871 , n280872 );
buf ( n280874 , n280873 );
not ( n280875 , RI19aae7a0_2465);
or ( n280876 , n25328 , n280875 );
not ( n280877 , RI19aa44f8_2535);
or ( n280878 , n25335 , n280877 );
nand ( n280879 , n280876 , n280878 );
buf ( n280880 , n280879 );
nand ( n280881 , n267768 , n280461 );
or ( n280882 , n267758 , n280881 );
nor ( n280883 , n267757 , n256376 );
nand ( n280884 , n280883 , n280881 );
nand ( n280885 , n35431 , n26338 );
nand ( n280886 , n280882 , n280884 , n280885 );
buf ( n280887 , n280886 );
nand ( n280888 , n261163 , n277092 , n277089 );
not ( n280889 , n261159 );
not ( n280890 , n277089 );
or ( n280891 , n280889 , n280890 );
nor ( n280892 , n277092 , n219702 );
nand ( n280893 , n280891 , n280892 );
nand ( n280894 , n49054 , n205926 );
nand ( n280895 , n280888 , n280893 , n280894 );
buf ( n280896 , n280895 );
nand ( n280897 , n267860 , n267871 );
or ( n280898 , n261489 , n280897 );
not ( n280899 , n267871 );
not ( n280900 , n261473 );
or ( n280901 , n280899 , n280900 );
nor ( n280902 , n267860 , n252258 );
nand ( n280903 , n280901 , n280902 );
nand ( n280904 , n31577 , n29867 );
nand ( n280905 , n280898 , n280903 , n280904 );
buf ( n280906 , n280905 );
not ( n280907 , n25640 );
not ( n280908 , n263819 );
or ( n280909 , n280907 , n280908 );
not ( n280910 , n235173 );
not ( n280911 , n248446 );
or ( n280912 , n280910 , n280911 );
not ( n280913 , n235173 );
nand ( n280914 , n280913 , n248455 );
nand ( n280915 , n280912 , n280914 );
and ( n280916 , n280915 , n248386 );
not ( n280917 , n280915 );
and ( n280918 , n280917 , n255830 );
nor ( n280919 , n280916 , n280918 );
nand ( n280920 , n280919 , n275591 );
and ( n280921 , n280920 , n273622 );
not ( n280922 , n280920 );
not ( n280923 , n273622 );
and ( n280924 , n280922 , n280923 );
nor ( n280925 , n280921 , n280924 );
or ( n280926 , n280925 , n226003 );
nand ( n280927 , n280909 , n280926 );
buf ( n280928 , n280927 );
or ( n280929 , n25328 , n267106 );
not ( n280930 , RI19a89720_2728);
or ( n280931 , n25335 , n280930 );
nand ( n280932 , n280929 , n280931 );
buf ( n280933 , n280932 );
not ( n280934 , n29742 );
not ( n280935 , n253009 );
or ( n280936 , n280934 , n280935 );
or ( n280937 , n253009 , n29742 );
nand ( n280938 , n280936 , n280937 );
and ( n280939 , n280938 , n263207 );
not ( n280940 , n280938 );
and ( n280941 , n280940 , n253015 );
nor ( n280942 , n280939 , n280941 );
nand ( n280943 , n280942 , n205649 );
not ( n280944 , n260256 );
nand ( n280945 , n280944 , n260258 );
or ( n280946 , n280943 , n280945 );
not ( n280947 , n280942 );
not ( n280948 , n280944 );
or ( n280949 , n280947 , n280948 );
nor ( n280950 , n260258 , n54208 );
nand ( n280951 , n280949 , n280950 );
nand ( n280952 , n241068 , n33209 );
nand ( n280953 , n280946 , n280951 , n280952 );
buf ( n280954 , n280953 );
not ( n280955 , n256180 );
nand ( n280956 , n280955 , n256208 );
not ( n280957 , n278161 );
or ( n280958 , n280956 , n280957 );
not ( n280959 , n259175 );
nand ( n280960 , n280959 , n280956 );
nand ( n280961 , n35431 , n26124 );
nand ( n280962 , n280958 , n280960 , n280961 );
buf ( n280963 , n280962 );
or ( n280964 , n226819 , n277373 );
not ( n280965 , RI19a87920_2741);
or ( n280966 , n25335 , n280965 );
nand ( n280967 , n280964 , n280966 );
buf ( n280968 , n280967 );
not ( n280969 , n39120 );
not ( n280970 , n245943 );
or ( n280971 , n280969 , n280970 );
nand ( n280972 , n263671 , n263683 );
and ( n280973 , n280972 , n275548 );
not ( n280974 , n280972 );
and ( n280975 , n280974 , n275547 );
nor ( n280976 , n280973 , n280975 );
or ( n280977 , n280976 , n250068 );
nand ( n280978 , n280971 , n280977 );
buf ( n280979 , n280978 );
nor ( n280980 , n53676 , n268556 );
nand ( n280981 , n272494 , n280980 );
not ( n280982 , n268557 );
not ( n280983 , n270347 );
or ( n280984 , n280982 , n280983 );
nand ( n280985 , n280984 , n53148 );
nand ( n280986 , n31577 , n31857 );
nand ( n280987 , n280981 , n280985 , n280986 );
buf ( n280988 , n280987 );
not ( n280989 , n40852 );
not ( n280990 , n244606 );
or ( n280991 , n280989 , n280990 );
not ( n280992 , RI1754ad38_55);
or ( n280993 , n269544 , n280992 );
nand ( n280994 , n280991 , n280993 );
buf ( n280995 , n280994 );
nand ( n280996 , n263807 , n263800 );
or ( n280997 , n280996 , n277166 );
nand ( n280998 , n267312 , n280996 );
nand ( n280999 , n35431 , n32586 );
nand ( n281000 , n280997 , n280998 , n280999 );
buf ( n281001 , n281000 );
nand ( n281002 , n261311 , n267906 );
or ( n281003 , n261326 , n281002 );
not ( n281004 , n267906 );
not ( n281005 , n261297 );
or ( n281006 , n281004 , n281005 );
nor ( n281007 , n261311 , n240080 );
nand ( n281008 , n281006 , n281007 );
nand ( n281009 , n238638 , n33654 );
nand ( n281010 , n281003 , n281008 , n281009 );
buf ( n281011 , n281010 );
or ( n281012 , n259010 , n266231 );
nor ( n281013 , n260473 , n266230 );
nand ( n281014 , n259034 , n281013 );
nand ( n281015 , n266230 , n247444 );
not ( n281016 , n281015 );
not ( n281017 , n260474 );
and ( n281018 , n281016 , n281017 );
and ( n281019 , n35431 , n26209 );
nor ( n281020 , n281018 , n281019 );
nand ( n281021 , n281012 , n281014 , n281020 );
buf ( n281022 , n281021 );
not ( n281023 , n210564 );
not ( n281024 , n31577 );
or ( n281025 , n281023 , n281024 );
nand ( n281026 , n273374 , n273371 );
not ( n281027 , n35734 );
not ( n281028 , n236883 );
or ( n281029 , n281027 , n281028 );
or ( n281030 , n236883 , n35734 );
nand ( n281031 , n281029 , n281030 );
not ( n281032 , n281031 );
not ( n281033 , n236994 );
and ( n281034 , n281032 , n281033 );
and ( n281035 , n281031 , n236997 );
nor ( n281036 , n281034 , n281035 );
not ( n281037 , n281036 );
and ( n281038 , n281026 , n281037 );
not ( n281039 , n281026 );
and ( n281040 , n281039 , n281036 );
nor ( n281041 , n281038 , n281040 );
or ( n281042 , n281041 , n254515 );
nand ( n281043 , n281025 , n281042 );
buf ( n281044 , n281043 );
not ( n281045 , n28176 );
not ( n281046 , n245943 );
or ( n281047 , n281045 , n281046 );
not ( n281048 , n43013 );
nand ( n281049 , n254201 , n273782 );
not ( n281050 , n281049 );
and ( n281051 , n281048 , n281050 );
and ( n281052 , n43013 , n281049 );
nor ( n281053 , n281051 , n281052 );
or ( n281054 , n281053 , n260760 );
nand ( n281055 , n281047 , n281054 );
buf ( n281056 , n281055 );
not ( n281057 , n26157 );
not ( n281058 , n256877 );
or ( n281059 , n281057 , n281058 );
or ( n281060 , n267305 , n26157 );
nand ( n281061 , n281059 , n281060 );
and ( n281062 , n281061 , n50604 );
not ( n281063 , n281061 );
and ( n281064 , n281063 , n50540 );
nor ( n281065 , n281062 , n281064 );
not ( n281066 , n281065 );
nor ( n281067 , n271754 , n281066 );
or ( n281068 , n280398 , n281067 );
nor ( n281069 , n280397 , n222533 );
nand ( n281070 , n281069 , n281067 );
nand ( n281071 , n31576 , n31457 );
nand ( n281072 , n281068 , n281070 , n281071 );
buf ( n281073 , n281072 );
not ( n281074 , n25726 );
not ( n281075 , n245702 );
or ( n281076 , n281074 , n281075 );
not ( n281077 , n264677 );
nand ( n281078 , n264664 , n281077 );
not ( n281079 , n281078 );
not ( n281080 , n277457 );
and ( n281081 , n281079 , n281080 );
and ( n281082 , n281078 , n277457 );
nor ( n281083 , n281081 , n281082 );
or ( n281084 , n281083 , n259425 );
nand ( n281085 , n281076 , n281084 );
buf ( n281086 , n281085 );
not ( n281087 , n245713 );
not ( n281088 , n281087 );
not ( n281089 , n230367 );
or ( n281090 , n281088 , n281089 );
not ( n281091 , n281087 );
nand ( n281092 , n281091 , n230374 );
nand ( n281093 , n281090 , n281092 );
and ( n281094 , n281093 , n245265 );
not ( n281095 , n281093 );
and ( n281096 , n281095 , n52757 );
nor ( n281097 , n281094 , n281096 );
nor ( n281098 , n281097 , n226004 );
not ( n281099 , n251732 );
nor ( n281100 , n281099 , n268598 );
nand ( n281101 , n281098 , n281100 );
not ( n281102 , n281097 );
not ( n281103 , n281102 );
not ( n281104 , n251732 );
or ( n281105 , n281103 , n281104 );
not ( n281106 , n268598 );
nor ( n281107 , n281106 , n253358 );
nand ( n281108 , n281105 , n281107 );
nand ( n281109 , n237714 , n41848 );
nand ( n281110 , n281101 , n281108 , n281109 );
buf ( n281111 , n281110 );
not ( n281112 , n258897 );
not ( n281113 , n266787 );
not ( n281114 , n281113 );
or ( n281115 , n281112 , n281114 );
nand ( n281116 , n281115 , n251183 );
nand ( n281117 , n258901 , n251182 , n281113 );
nand ( n281118 , n41944 , n29219 );
nand ( n281119 , n281116 , n281117 , n281118 );
buf ( n281120 , n281119 );
not ( n281121 , n29292 );
not ( n281122 , n251717 );
or ( n281123 , n281121 , n281122 );
not ( n281124 , n266171 );
nand ( n281125 , n263222 , n263237 );
not ( n281126 , n281125 );
and ( n281127 , n281124 , n281126 );
and ( n281128 , n266171 , n281125 );
nor ( n281129 , n281127 , n281128 );
or ( n281130 , n281129 , n254882 );
nand ( n281131 , n281123 , n281130 );
buf ( n281132 , n281131 );
buf ( n281133 , n42616 );
not ( n281134 , n33328 );
not ( n281135 , n258213 );
or ( n281136 , n281134 , n281135 );
nand ( n281137 , n266858 , n275990 );
not ( n281138 , n265222 );
and ( n281139 , n281137 , n281138 );
not ( n281140 , n281137 );
and ( n281141 , n281140 , n265222 );
nor ( n281142 , n281139 , n281141 );
or ( n281143 , n281142 , n255707 );
nand ( n281144 , n281136 , n281143 );
buf ( n281145 , n281144 );
not ( n281146 , n248222 );
nand ( n281147 , n281146 , n248289 );
not ( n281148 , n250259 );
or ( n281149 , n281147 , n281148 );
nor ( n281150 , n250257 , n251361 );
nand ( n281151 , n281147 , n281150 );
nand ( n281152 , n31577 , n37732 );
nand ( n281153 , n281149 , n281151 , n281152 );
buf ( n281154 , n281153 );
buf ( n281155 , n42281 );
buf ( n281156 , n35455 );
nand ( n281157 , n259646 , n278136 );
or ( n281158 , n276384 , n281157 );
nand ( n281159 , n251317 , n281157 );
nand ( n281160 , n256673 , n28265 );
nand ( n281161 , n281158 , n281159 , n281160 );
buf ( n281162 , n281161 );
buf ( n281163 , n39199 );
not ( n281164 , n244477 );
nand ( n281165 , n281164 , n227713 );
or ( n281166 , n260172 , n281165 );
not ( n281167 , n227713 );
not ( n281168 , n244464 );
or ( n281169 , n281167 , n281168 );
nor ( n281170 , n281164 , n35428 );
nand ( n281171 , n281169 , n281170 );
nand ( n281172 , n241068 , n29658 );
nand ( n281173 , n281166 , n281171 , n281172 );
buf ( n281174 , n281173 );
not ( n281175 , n278810 );
nor ( n281176 , n281175 , n278821 );
or ( n281177 , n271968 , n281176 );
nor ( n281178 , n271967 , n252070 );
nand ( n281179 , n281178 , n281176 );
nand ( n281180 , n39767 , n37429 );
nand ( n281181 , n281177 , n281179 , n281180 );
buf ( n281182 , n281181 );
nor ( n281183 , n260832 , n277488 );
nand ( n281184 , n277477 , n281183 );
not ( n281185 , n277488 );
not ( n281186 , n281185 );
not ( n281187 , n264749 );
or ( n281188 , n281186 , n281187 );
nand ( n281189 , n281188 , n260803 );
nand ( n281190 , n244840 , n30669 );
nand ( n281191 , n281184 , n281189 , n281190 );
buf ( n281192 , n281191 );
not ( n281193 , RI19ab4560_2421);
or ( n281194 , n226819 , n281193 );
not ( n281195 , RI19aaa510_2493);
or ( n281196 , n226822 , n281195 );
nand ( n281197 , n281194 , n281196 );
buf ( n281198 , n281197 );
nor ( n281199 , n267731 , n52445 );
not ( n281200 , n281199 );
nand ( n281201 , n255502 , n267732 );
or ( n281202 , n281200 , n281201 );
not ( n281203 , n267732 );
not ( n281204 , n267731 );
not ( n281205 , n281204 );
or ( n281206 , n281203 , n281205 );
nor ( n281207 , n255502 , n243204 );
nand ( n281208 , n281206 , n281207 );
nand ( n281209 , n39766 , n227655 );
nand ( n281210 , n281202 , n281208 , n281209 );
buf ( n281211 , n281210 );
not ( n281212 , n33417 );
not ( n281213 , n51381 );
or ( n281214 , n281212 , n281213 );
nand ( n281215 , n261081 , n279576 );
and ( n281216 , n281215 , n55332 );
not ( n281217 , n281215 );
and ( n281218 , n281217 , n55737 );
nor ( n281219 , n281216 , n281218 );
or ( n281220 , n281219 , n258327 );
nand ( n281221 , n281214 , n281220 );
buf ( n281222 , n281221 );
not ( n281223 , n38284 );
not ( n281224 , n55760 );
or ( n281225 , n281223 , n281224 );
not ( n281226 , n279153 );
nand ( n281227 , n281226 , n256450 );
and ( n281228 , n281227 , n261634 );
not ( n281229 , n281227 );
and ( n281230 , n281229 , n279155 );
nor ( n281231 , n281228 , n281230 );
or ( n281232 , n281231 , n46425 );
nand ( n281233 , n281225 , n281232 );
buf ( n281234 , n281233 );
not ( n281235 , RI19ab7a58_2397);
or ( n281236 , n25328 , n281235 );
or ( n281237 , n25335 , n219716 );
nand ( n281238 , n281236 , n281237 );
buf ( n281239 , n281238 );
nand ( n281240 , n260892 , n237873 );
or ( n281241 , n260876 , n281240 );
not ( n281242 , n237873 );
not ( n281243 , n260875 );
or ( n281244 , n281242 , n281243 );
nor ( n281245 , n260892 , n276592 );
nand ( n281246 , n281244 , n281245 );
nand ( n281247 , n31577 , n48456 );
nand ( n281248 , n281241 , n281246 , n281247 );
buf ( n281249 , n281248 );
nand ( n281250 , n274226 , n263067 );
or ( n281251 , n268381 , n281250 );
not ( n281252 , n274226 );
not ( n281253 , n268380 );
or ( n281254 , n281252 , n281253 );
nor ( n281255 , n263067 , n247276 );
nand ( n281256 , n281254 , n281255 );
nand ( n281257 , n247744 , n25886 );
nand ( n281258 , n281251 , n281256 , n281257 );
buf ( n281259 , n281258 );
not ( n281260 , RI19a9b420_2603);
or ( n281261 , n25328 , n281260 );
or ( n281262 , n25335 , n266240 );
nand ( n281263 , n281261 , n281262 );
buf ( n281264 , n281263 );
or ( n281265 , n25328 , n256304 );
or ( n281266 , n25336 , n277577 );
nand ( n281267 , n281265 , n281266 );
buf ( n281268 , n281267 );
or ( n281269 , n226819 , n261613 );
or ( n281270 , n25335 , n279510 );
nand ( n281271 , n281269 , n281270 );
buf ( n281272 , n281271 );
or ( n281273 , n25328 , n256382 );
not ( n281274 , RI19a8d410_2702);
or ( n281275 , n25335 , n281274 );
nand ( n281276 , n281273 , n281275 );
buf ( n281277 , n281276 );
buf ( n281278 , n28860 );
nand ( n281279 , n278254 , n271667 );
or ( n281280 , n279076 , n281279 );
nand ( n281281 , n257685 , n281279 );
nand ( n281282 , n35431 , n45290 );
nand ( n281283 , n281280 , n281281 , n281282 );
buf ( n281284 , n281283 );
buf ( n281285 , n30184 );
buf ( n281286 , n207164 );
buf ( n281287 , n30741 );
not ( n281288 , n264462 );
nand ( n281289 , n264466 , n281288 );
not ( n281290 , n247582 );
or ( n281291 , n281289 , n281290 );
nand ( n281292 , n281289 , n272741 );
nand ( n281293 , n255116 , n38428 );
nand ( n281294 , n281291 , n281292 , n281293 );
buf ( n281295 , n281294 );
not ( n281296 , RI19ac0a40_2326);
or ( n281297 , n25328 , n281296 );
not ( n281298 , RI19a84950_2762);
or ( n281299 , n25335 , n281298 );
nand ( n281300 , n281297 , n281299 );
buf ( n281301 , n281300 );
buf ( n281302 , n30576 );
not ( n281303 , n32171 );
not ( n281304 , n234453 );
or ( n281305 , n281303 , n281304 );
not ( n281306 , n241667 );
nand ( n281307 , n281306 , n260277 );
and ( n281308 , n281307 , n262268 );
not ( n281309 , n281307 );
not ( n281310 , n262268 );
and ( n281311 , n281309 , n281310 );
nor ( n281312 , n281308 , n281311 );
or ( n281313 , n281312 , n244837 );
nand ( n281314 , n281305 , n281313 );
buf ( n281315 , n281314 );
nand ( n281316 , n269975 , n205649 );
nand ( n281317 , n276242 , n276253 );
or ( n281318 , n281316 , n281317 );
not ( n281319 , n276253 );
not ( n281320 , n269975 );
or ( n281321 , n281319 , n281320 );
nor ( n281322 , n276242 , n226003 );
nand ( n281323 , n281321 , n281322 );
nand ( n281324 , n246217 , n31244 );
nand ( n281325 , n281318 , n281323 , n281324 );
buf ( n281326 , n281325 );
buf ( n281327 , n209367 );
or ( n281328 , n25328 , n280161 );
or ( n281329 , n25335 , n260241 );
nand ( n281330 , n281328 , n281329 );
buf ( n281331 , n281330 );
buf ( n281332 , n208196 );
nor ( n281333 , n249144 , n55108 );
not ( n281334 , n281333 );
nand ( n281335 , n240059 , n249213 );
or ( n281336 , n281334 , n281335 );
not ( n281337 , n249213 );
not ( n281338 , n249144 );
not ( n281339 , n281338 );
or ( n281340 , n281337 , n281339 );
nor ( n281341 , n240059 , n35427 );
nand ( n281342 , n281340 , n281341 );
nand ( n281343 , n31577 , n204457 );
nand ( n281344 , n281336 , n281342 , n281343 );
buf ( n281345 , n281344 );
buf ( n281346 , n28324 );
not ( n281347 , n252738 );
not ( n281348 , n252725 );
not ( n281349 , n281348 );
or ( n281350 , n281347 , n281349 );
nor ( n281351 , n264240 , n249531 );
nand ( n281352 , n281350 , n281351 );
nor ( n281353 , n252725 , n242391 );
nor ( n281354 , n264239 , n252737 );
nand ( n281355 , n281353 , n281354 );
nand ( n281356 , n246460 , n38334 );
nand ( n281357 , n281352 , n281355 , n281356 );
buf ( n281358 , n281357 );
not ( n281359 , n30146 );
not ( n281360 , n234453 );
or ( n281361 , n281359 , n281360 );
not ( n281362 , n40016 );
not ( n281363 , n281362 );
not ( n281364 , n235807 );
or ( n281365 , n281363 , n281364 );
not ( n281366 , n281362 );
nand ( n281367 , n281366 , n235815 );
nand ( n281368 , n281365 , n281367 );
and ( n281369 , n281368 , n235879 );
not ( n281370 , n281368 );
and ( n281371 , n281370 , n235888 );
nor ( n281372 , n281369 , n281371 );
not ( n281373 , n281372 );
nand ( n281374 , n281373 , n242208 );
and ( n281375 , n281374 , n242277 );
not ( n281376 , n281374 );
and ( n281377 , n281376 , n242276 );
nor ( n281378 , n281375 , n281377 );
or ( n281379 , n281378 , n52445 );
nand ( n281380 , n281361 , n281379 );
buf ( n281381 , n281380 );
buf ( n281382 , n215143 );
buf ( n281383 , n29503 );
buf ( n281384 , n37851 );
buf ( n281385 , n35568 );
buf ( n281386 , n205210 );
buf ( n281387 , n39790 );
not ( n281388 , n251820 );
not ( n281389 , n258512 );
or ( n281390 , n281388 , n281389 );
not ( n281391 , n251820 );
nand ( n281392 , n281391 , n259214 );
nand ( n281393 , n281390 , n281392 );
and ( n281394 , n281393 , n260558 );
not ( n281395 , n281393 );
and ( n281396 , n281395 , n260551 );
nor ( n281397 , n281394 , n281396 );
nand ( n281398 , n279108 , n255370 , n281397 );
not ( n281399 , n279106 );
not ( n281400 , n255370 );
or ( n281401 , n281399 , n281400 );
nor ( n281402 , n281397 , n33254 );
nand ( n281403 , n281401 , n281402 );
nand ( n281404 , n250916 , n36425 );
nand ( n281405 , n281398 , n281403 , n281404 );
buf ( n281406 , n281405 );
or ( n281407 , n226819 , n280812 );
or ( n281408 , n25335 , n259714 );
nand ( n281409 , n281407 , n281408 );
buf ( n281410 , n281409 );
nand ( n281411 , n266171 , n268715 );
or ( n281412 , n266157 , n281411 );
not ( n281413 , n266171 );
not ( n281414 , n266156 );
or ( n281415 , n281413 , n281414 );
nor ( n281416 , n268715 , n222533 );
nand ( n281417 , n281415 , n281416 );
nand ( n281418 , n246217 , n30564 );
nand ( n281419 , n281412 , n281417 , n281418 );
buf ( n281420 , n281419 );
or ( n281421 , n25328 , n275397 );
or ( n281422 , n25335 , n273100 );
nand ( n281423 , n281421 , n281422 );
buf ( n281424 , n281423 );
not ( n281425 , n237873 );
nand ( n281426 , n281425 , n279307 );
or ( n281427 , n260876 , n281426 );
not ( n281428 , n260880 );
nand ( n281429 , n281428 , n281426 );
nand ( n281430 , n51381 , n204757 );
nand ( n281431 , n281427 , n281429 , n281430 );
buf ( n281432 , n281431 );
not ( n281433 , n32619 );
not ( n281434 , n237361 );
or ( n281435 , n281433 , n281434 );
nand ( n281436 , n246894 , n249761 );
and ( n281437 , n281436 , n246770 );
not ( n281438 , n281436 );
and ( n281439 , n281438 , n246771 );
nor ( n281440 , n281437 , n281439 );
or ( n281441 , n281440 , n257851 );
nand ( n281442 , n281435 , n281441 );
buf ( n281443 , n281442 );
nand ( n281444 , n264035 , n280366 );
or ( n281445 , n280370 , n281444 );
not ( n281446 , n280366 );
not ( n281447 , n280369 );
or ( n281448 , n281446 , n281447 );
nand ( n281449 , n281448 , n264036 );
nand ( n281450 , n247585 , n42616 );
nand ( n281451 , n281445 , n281449 , n281450 );
buf ( n281452 , n281451 );
nand ( n281453 , n269558 , n257792 );
not ( n281454 , n246718 );
not ( n281455 , n45261 );
or ( n281456 , n281454 , n281455 );
not ( n281457 , n246718 );
nand ( n281458 , n281457 , n45253 );
nand ( n281459 , n281456 , n281458 );
and ( n281460 , n281459 , n255248 );
not ( n281461 , n281459 );
and ( n281462 , n281461 , n255245 );
nor ( n281463 , n281460 , n281462 );
not ( n281464 , n281463 );
nand ( n281465 , n269565 , n281464 );
or ( n281466 , n281453 , n281465 );
not ( n281467 , n281464 );
not ( n281468 , n269558 );
or ( n281469 , n281467 , n281468 );
nor ( n281470 , n269565 , n221279 );
nand ( n281471 , n281469 , n281470 );
nand ( n281472 , n31576 , n25699 );
nand ( n281473 , n281466 , n281471 , n281472 );
buf ( n281474 , n281473 );
or ( n281475 , n25328 , n272733 );
not ( n281476 , RI19ac2840_2310);
or ( n281477 , n25335 , n281476 );
nand ( n281478 , n281475 , n281477 );
buf ( n281479 , n281478 );
buf ( n281480 , n39990 );
buf ( n281481 , n33742 );
nand ( n281482 , n265968 , n205649 );
nor ( n281483 , n265980 , n267064 );
or ( n281484 , n281482 , n281483 );
nand ( n281485 , n265969 , n281483 );
nand ( n281486 , n35431 , n39344 );
nand ( n281487 , n281484 , n281485 , n281486 );
buf ( n281488 , n281487 );
not ( n281489 , n36508 );
not ( n281490 , n245943 );
or ( n281491 , n281489 , n281490 );
nand ( n281492 , n275135 , n250592 );
and ( n281493 , n281492 , n275123 );
not ( n281494 , n281492 );
and ( n281495 , n281494 , n275124 );
nor ( n281496 , n281493 , n281495 );
or ( n281497 , n281496 , n262962 );
nand ( n281498 , n281491 , n281497 );
buf ( n281499 , n281498 );
not ( n281500 , RI19aa9688_2500);
or ( n281501 , n25328 , n281500 );
or ( n281502 , n25336 , n262143 );
nand ( n281503 , n281501 , n281502 );
buf ( n281504 , n281503 );
or ( n281505 , n226819 , n275621 );
not ( n281506 , RI19a920f0_2668);
or ( n281507 , n226822 , n281506 );
nand ( n281508 , n281505 , n281507 );
buf ( n281509 , n281508 );
buf ( n281510 , RI19ad12b8_2203);
and ( n281511 , n25326 , n281510 );
buf ( n281512 , n281511 );
nand ( n281513 , n269728 , n223839 );
nand ( n281514 , n272376 , n269750 );
or ( n281515 , n281513 , n281514 );
not ( n281516 , n269750 );
not ( n281517 , n269728 );
or ( n281518 , n281516 , n281517 );
nor ( n281519 , n272376 , n50944 );
nand ( n281520 , n281518 , n281519 );
nand ( n281521 , n41944 , n30147 );
nand ( n281522 , n281515 , n281520 , n281521 );
buf ( n281523 , n281522 );
nand ( n281524 , n269268 , n266527 );
or ( n281525 , n266692 , n281524 );
nor ( n281526 , n266691 , n33254 );
nand ( n281527 , n281526 , n281524 );
nand ( n281528 , n258743 , n33089 );
nand ( n281529 , n281525 , n281527 , n281528 );
buf ( n281530 , n281529 );
not ( n281531 , n252576 );
not ( n281532 , n265819 );
or ( n281533 , n281531 , n281532 );
nor ( n281534 , n279644 , n31571 );
nand ( n281535 , n281533 , n281534 );
nand ( n281536 , n252581 , n279644 , n265819 );
nand ( n281537 , n35431 , n43228 );
nand ( n281538 , n281535 , n281536 , n281537 );
buf ( n281539 , n281538 );
or ( n281540 , n25328 , n254424 );
not ( n281541 , RI19ab7da0_2396);
or ( n281542 , n25335 , n281541 );
nand ( n281543 , n281540 , n281542 );
buf ( n281544 , n281543 );
not ( n281545 , n278683 );
nand ( n281546 , n279919 , n256629 , n281545 );
not ( n281547 , n256629 );
not ( n281548 , n256606 );
or ( n281549 , n281547 , n281548 );
nor ( n281550 , n281545 , n47173 );
nand ( n281551 , n281549 , n281550 );
nand ( n281552 , n31577 , n25687 );
nand ( n281553 , n281546 , n281551 , n281552 );
buf ( n281554 , n281553 );
nand ( n281555 , n268798 , n276201 );
and ( n281556 , n281555 , n268809 , n253928 );
not ( n281557 , n29486 );
nor ( n281558 , n281557 , n275788 );
nor ( n281559 , n281556 , n281558 );
nor ( n281560 , n276202 , n236795 );
nand ( n281561 , n281560 , n268810 , n268798 );
nand ( n281562 , n281559 , n281561 );
buf ( n281563 , n281562 );
not ( n281564 , n32795 );
not ( n281565 , n51381 );
or ( n281566 , n281564 , n281565 );
not ( n281567 , n237706 );
nand ( n281568 , n281567 , n237596 );
not ( n281569 , n281568 );
not ( n281570 , n270132 );
and ( n281571 , n281569 , n281570 );
and ( n281572 , n281568 , n270132 );
nor ( n281573 , n281571 , n281572 );
or ( n281574 , n281573 , n258280 );
nand ( n281575 , n281566 , n281574 );
buf ( n281576 , n281575 );
not ( n281577 , n35384 );
not ( n281578 , n234453 );
or ( n281579 , n281577 , n281578 );
not ( n281580 , n240017 );
not ( n281581 , n281580 );
not ( n281582 , n40194 );
or ( n281583 , n281581 , n281582 );
not ( n281584 , n281580 );
nand ( n281585 , n281584 , n40203 );
nand ( n281586 , n281583 , n281585 );
and ( n281587 , n281586 , n251346 );
not ( n281588 , n281586 );
and ( n281589 , n281588 , n251350 );
nor ( n281590 , n281587 , n281589 );
nand ( n281591 , n271480 , n281590 );
and ( n281592 , n281591 , n271469 );
not ( n281593 , n281591 );
not ( n281594 , n271469 );
and ( n281595 , n281593 , n281594 );
nor ( n281596 , n281592 , n281595 );
or ( n281597 , n281596 , n264257 );
nand ( n281598 , n281579 , n281597 );
buf ( n281599 , n281598 );
nand ( n281600 , n262416 , n253397 );
not ( n281601 , n274088 );
nand ( n281602 , n281601 , n262438 );
or ( n281603 , n281600 , n281602 );
not ( n281604 , n262438 );
not ( n281605 , n262416 );
or ( n281606 , n281604 , n281605 );
nor ( n281607 , n281601 , n221279 );
nand ( n281608 , n281606 , n281607 );
nand ( n281609 , n35431 , n26282 );
nand ( n281610 , n281603 , n281608 , n281609 );
buf ( n281611 , n281610 );
not ( n281612 , n205193 );
not ( n281613 , n241068 );
or ( n281614 , n281612 , n281613 );
nand ( n281615 , n267673 , n267686 );
not ( n281616 , n238589 );
not ( n281617 , n241122 );
or ( n281618 , n281616 , n281617 );
not ( n281619 , n238589 );
nand ( n281620 , n281619 , n241131 );
nand ( n281621 , n281618 , n281620 );
and ( n281622 , n281621 , n241181 );
not ( n281623 , n281621 );
and ( n281624 , n281623 , n241180 );
nor ( n281625 , n281622 , n281624 );
and ( n281626 , n281615 , n281625 );
not ( n281627 , n281615 );
not ( n281628 , n281625 );
and ( n281629 , n281627 , n281628 );
nor ( n281630 , n281626 , n281629 );
or ( n281631 , n281630 , n261009 );
nand ( n281632 , n281614 , n281631 );
buf ( n281633 , n281632 );
nand ( n281634 , n258395 , n266957 );
not ( n281635 , n266961 );
or ( n281636 , n281634 , n281635 );
nand ( n281637 , n281634 , n262247 );
nand ( n281638 , n241378 , n27742 );
nand ( n281639 , n281636 , n281637 , n281638 );
buf ( n281640 , n281639 );
or ( n281641 , n233507 , n266988 );
or ( n281642 , n226822 , n270211 );
nand ( n281643 , n281641 , n281642 );
buf ( n281644 , n281643 );
or ( n281645 , n25328 , n272213 );
or ( n281646 , n25335 , n281193 );
nand ( n281647 , n281645 , n281646 );
buf ( n281648 , n281647 );
buf ( n281649 , n35238 );
buf ( n281650 , n220690 );
or ( n281651 , n25328 , n271712 );
or ( n281652 , n25336 , n273583 );
nand ( n281653 , n281651 , n281652 );
buf ( n281654 , n281653 );
not ( n281655 , n25830 );
not ( n281656 , n51381 );
or ( n281657 , n281655 , n281656 );
nand ( n281658 , n250376 , n45729 );
and ( n281659 , n281658 , n45264 );
not ( n281660 , n281658 );
and ( n281661 , n281660 , n223026 );
nor ( n281662 , n281659 , n281661 );
or ( n281663 , n281662 , n258280 );
nand ( n281664 , n281657 , n281663 );
buf ( n281665 , n281664 );
nand ( n281666 , n235374 , n235213 );
or ( n281667 , n268045 , n281666 );
not ( n281668 , n235213 );
not ( n281669 , n268044 );
or ( n281670 , n281668 , n281669 );
nor ( n281671 , n235374 , n33253 );
nand ( n281672 , n281670 , n281671 );
nand ( n281673 , n234024 , n38154 );
nand ( n281674 , n281667 , n281672 , n281673 );
buf ( n281675 , n281674 );
or ( n281676 , n25328 , n264289 );
or ( n281677 , n25336 , n281500 );
nand ( n281678 , n281676 , n281677 );
buf ( n281679 , n281678 );
or ( n281680 , n25328 , n270935 );
or ( n281681 , n25335 , n274542 );
nand ( n281682 , n281680 , n281681 );
buf ( n281683 , n281682 );
not ( n281684 , n276096 );
not ( n281685 , n276415 );
not ( n281686 , n281685 );
and ( n281687 , n281684 , n281686 );
and ( n281688 , n251712 , n226914 );
nor ( n281689 , n281687 , n281688 );
not ( n281690 , n249250 );
not ( n281691 , n244889 );
or ( n281692 , n281690 , n281691 );
not ( n281693 , n249250 );
nand ( n281694 , n281693 , n244899 );
nand ( n281695 , n281692 , n281694 );
and ( n281696 , n281695 , n244940 );
not ( n281697 , n281695 );
and ( n281698 , n281697 , n244955 );
nor ( n281699 , n281696 , n281698 );
nand ( n281700 , n276099 , n281699 , n281685 );
or ( n281701 , n276416 , n281699 );
nand ( n281702 , n281689 , n281700 , n281701 );
buf ( n281703 , n281702 );
not ( n281704 , n279801 );
nand ( n281705 , n281704 , n246215 );
or ( n281706 , n281705 , n280504 );
not ( n281707 , n246209 );
nand ( n281708 , n279802 , n281707 );
nand ( n281709 , n281708 , n280504 , n205649 );
nand ( n281710 , n241378 , n39381 );
nand ( n281711 , n281706 , n281709 , n281710 );
buf ( n281712 , n281711 );
nand ( n281713 , n276690 , n272711 );
nor ( n281714 , n268633 , n268645 );
or ( n281715 , n281713 , n281714 );
nor ( n281716 , n276690 , n247276 );
nand ( n281717 , n281716 , n281714 );
nand ( n281718 , n251465 , n37320 );
nand ( n281719 , n281715 , n281717 , n281718 );
buf ( n281720 , n281719 );
not ( n281721 , n271575 );
nor ( n281722 , n271167 , n278359 );
or ( n281723 , n281721 , n281722 );
nand ( n281724 , n271562 , n281722 );
nand ( n281725 , n246217 , n34992 );
nand ( n281726 , n281723 , n281724 , n281725 );
buf ( n281727 , n281726 );
buf ( n281728 , n25796 );
nand ( n281729 , n268821 , n276202 );
or ( n281730 , n269193 , n281729 );
not ( n281731 , n269192 );
not ( n281732 , n268821 );
or ( n281733 , n281731 , n281732 );
nand ( n281734 , n281733 , n281560 );
nand ( n281735 , n39767 , n33580 );
nand ( n281736 , n281730 , n281734 , n281735 );
buf ( n281737 , n281736 );
nand ( n281738 , n281037 , n274458 );
not ( n281739 , n273347 );
or ( n281740 , n281738 , n281739 );
nand ( n281741 , n273360 , n281738 );
nand ( n281742 , n247585 , n235477 );
nand ( n281743 , n281740 , n281741 , n281742 );
buf ( n281744 , n281743 );
nor ( n281745 , n218985 , n41937 );
nand ( n281746 , n279786 , n281745 );
not ( n281747 , n274993 );
not ( n281748 , n281747 );
not ( n281749 , n218984 );
or ( n281750 , n281748 , n281749 );
nor ( n281751 , n41938 , n35428 );
nand ( n281752 , n281750 , n281751 );
nand ( n281753 , n255116 , n28133 );
nand ( n281754 , n281746 , n281752 , n281753 );
buf ( n281755 , n281754 );
buf ( n281756 , RI175385e8_592);
and ( n281757 , n27883 , n281756 );
buf ( n281758 , n281757 );
not ( n281759 , n35365 );
not ( n281760 , n255116 );
or ( n281761 , n281759 , n281760 );
nand ( n281762 , n268240 , n272202 );
and ( n281763 , n281762 , n271242 );
not ( n281764 , n281762 );
not ( n281765 , n271242 );
and ( n281766 , n281764 , n281765 );
nor ( n281767 , n281763 , n281766 );
or ( n281768 , n281767 , n238223 );
nand ( n281769 , n281761 , n281768 );
buf ( n281770 , n281769 );
not ( n281771 , n33805 );
not ( n281772 , n245702 );
or ( n281773 , n281771 , n281772 );
not ( n281774 , n236950 );
not ( n281775 , n239298 );
or ( n281776 , n281774 , n281775 );
not ( n281777 , n236950 );
nand ( n281778 , n281777 , n239297 );
nand ( n281779 , n281776 , n281778 );
and ( n281780 , n281779 , n239391 );
not ( n281781 , n281779 );
and ( n281782 , n281781 , n239399 );
nor ( n281783 , n281780 , n281782 );
nand ( n281784 , n281783 , n280308 );
not ( n281785 , n281784 );
not ( n281786 , n280319 );
not ( n281787 , n281786 );
and ( n281788 , n281785 , n281787 );
and ( n281789 , n281784 , n281786 );
nor ( n281790 , n281788 , n281789 );
or ( n281791 , n281790 , n258328 );
nand ( n281792 , n281773 , n281791 );
buf ( n281793 , n281792 );
not ( n281794 , RI1754be90_18);
or ( n281795 , n51369 , n281794 );
not ( n281796 , n226822 );
not ( n281797 , n268836 );
and ( n281798 , n281796 , n281797 );
nor ( n281799 , n51365 , n273851 );
and ( n281800 , n51363 , n281799 );
nor ( n281801 , n281798 , n281800 );
nand ( n281802 , n281795 , n281801 );
buf ( n281803 , n281802 );
not ( n281804 , n25852 );
not ( n281805 , n244606 );
or ( n281806 , n281804 , n281805 );
not ( n281807 , RI1754c2c8_9);
or ( n281808 , n244611 , n281807 );
nand ( n281809 , n281806 , n281808 );
buf ( n281810 , n281809 );
or ( n281811 , n25328 , n279317 );
or ( n281812 , n25335 , n264734 );
nand ( n281813 , n281811 , n281812 );
buf ( n281814 , n281813 );
not ( n281815 , RI19a98888_2622);
or ( n281816 , n25328 , n281815 );
not ( n281817 , RI19a8e6d0_2694);
or ( n281818 , n25336 , n281817 );
nand ( n281819 , n281816 , n281818 );
buf ( n281820 , n281819 );
not ( n281821 , n221492 );
not ( n281822 , n245221 );
or ( n281823 , n281821 , n281822 );
not ( n281824 , n246019 );
nand ( n281825 , n281824 , n276506 );
and ( n281826 , n281825 , n260230 );
not ( n281827 , n281825 );
and ( n281828 , n281827 , n260229 );
nor ( n281829 , n281826 , n281828 );
or ( n281830 , n281829 , n252859 );
nand ( n281831 , n281823 , n281830 );
buf ( n281832 , n281831 );
nand ( n281833 , n257011 , n269864 );
or ( n281834 , n257001 , n281833 );
not ( n281835 , n257011 );
not ( n281836 , n257000 );
or ( n281837 , n281835 , n281836 );
nor ( n281838 , n269864 , n221279 );
nand ( n281839 , n281837 , n281838 );
nand ( n281840 , n39766 , n33466 );
nand ( n281841 , n281834 , n281839 , n281840 );
buf ( n281842 , n281841 );
not ( n281843 , RI1754c1d8_11);
or ( n281844 , n51369 , n281843 );
nand ( n281845 , n244606 , n36946 );
nand ( n281846 , n281844 , n281845 );
buf ( n281847 , n281846 );
not ( n281848 , RI19a86de0_2746);
or ( n281849 , n25328 , n281848 );
or ( n281850 , n25336 , n271039 );
nand ( n281851 , n281849 , n281850 );
buf ( n281852 , n281851 );
not ( n281853 , n279719 );
nand ( n281854 , n272692 , n281853 );
or ( n281855 , n272712 , n281854 );
not ( n281856 , n281853 );
not ( n281857 , n272677 );
or ( n281858 , n281856 , n281857 );
nor ( n281859 , n272692 , n249531 );
nand ( n281860 , n281858 , n281859 );
nand ( n281861 , n234448 , n25434 );
nand ( n281862 , n281855 , n281860 , n281861 );
buf ( n281863 , n281862 );
or ( n281864 , n233507 , n262967 );
or ( n281865 , n226822 , n271868 );
nand ( n281866 , n281864 , n281865 );
buf ( n281867 , n281866 );
not ( n281868 , n227097 );
not ( n281869 , n39766 );
or ( n281870 , n281868 , n281869 );
not ( n281871 , n254035 );
nand ( n281872 , n281871 , n273127 );
and ( n281873 , n281872 , n257455 );
not ( n281874 , n281872 );
not ( n281875 , n257455 );
and ( n281876 , n281874 , n281875 );
nor ( n281877 , n281873 , n281876 );
or ( n281878 , n281877 , n261009 );
nand ( n281879 , n281870 , n281878 );
buf ( n281880 , n281879 );
not ( n281881 , n30305 );
not ( n281882 , n233501 );
or ( n281883 , n281881 , n281882 );
nand ( n281884 , n275886 , n274734 );
not ( n281885 , n275497 );
and ( n281886 , n281884 , n281885 );
not ( n281887 , n281884 );
and ( n281888 , n281887 , n275497 );
nor ( n281889 , n281886 , n281888 );
or ( n281890 , n281889 , n234818 );
nand ( n281891 , n281883 , n281890 );
buf ( n281892 , n281891 );
nand ( n281893 , n265992 , n267074 );
or ( n281894 , n281482 , n281893 );
not ( n281895 , n265992 );
not ( n281896 , n265968 );
or ( n281897 , n281895 , n281896 );
nor ( n281898 , n267074 , n249531 );
nand ( n281899 , n281897 , n281898 );
nand ( n281900 , n35431 , n28559 );
nand ( n281901 , n281894 , n281899 , n281900 );
buf ( n281902 , n281901 );
nand ( n281903 , n239658 , n263867 );
not ( n281904 , n239402 );
or ( n281905 , n281903 , n281904 );
nor ( n281906 , n239783 , n234440 );
nand ( n281907 , n281903 , n281906 );
nand ( n281908 , n244987 , n31093 );
nand ( n281909 , n281905 , n281907 , n281908 );
buf ( n281910 , n281909 );
not ( n281911 , n239933 );
nand ( n281912 , n281911 , n252858 );
nand ( n281913 , n249144 , n240077 );
or ( n281914 , n281912 , n281913 );
not ( n281915 , n240077 );
not ( n281916 , n281911 );
or ( n281917 , n281915 , n281916 );
nand ( n281918 , n281917 , n281333 );
nand ( n281919 , n244484 , n206789 );
nand ( n281920 , n281914 , n281918 , n281919 );
buf ( n281921 , n281920 );
not ( n281922 , RI19ace168_2224);
or ( n281923 , n25328 , n281922 );
or ( n281924 , n226822 , n273499 );
nand ( n281925 , n281923 , n281924 );
buf ( n281926 , n281925 );
or ( n281927 , n25328 , n266413 );
or ( n281928 , n25336 , n273686 );
nand ( n281929 , n281927 , n281928 );
buf ( n281930 , n281929 );
nand ( n281931 , n266863 , n265210 , n275991 );
not ( n281932 , n265234 );
not ( n281933 , n265210 );
or ( n281934 , n281932 , n281933 );
nor ( n281935 , n275991 , n31572 );
nand ( n281936 , n281934 , n281935 );
nand ( n281937 , n46083 , n31241 );
nand ( n281938 , n281931 , n281936 , n281937 );
buf ( n281939 , n281938 );
not ( n281940 , n266032 );
not ( n281941 , n255066 );
nand ( n281942 , n281941 , n255092 );
or ( n281943 , n281940 , n281942 );
not ( n281944 , n281941 );
not ( n281945 , n266015 );
or ( n281946 , n281944 , n281945 );
nor ( n281947 , n255092 , n226955 );
nand ( n281948 , n281946 , n281947 );
nand ( n281949 , n246217 , n33793 );
nand ( n281950 , n281943 , n281948 , n281949 );
buf ( n281951 , n281950 );
nand ( n281952 , n235896 , n232864 , n264127 );
not ( n281953 , n55107 );
not ( n281954 , n232864 );
or ( n281955 , n281953 , n281954 );
nor ( n281956 , n264127 , n40465 );
nand ( n281957 , n281955 , n281956 );
nand ( n281958 , n245414 , n26217 );
nand ( n281959 , n281952 , n281957 , n281958 );
buf ( n281960 , n281959 );
nand ( n281961 , n268211 , n277593 );
or ( n281962 , n281961 , n277596 );
nand ( n281963 , n277593 , n268206 );
nand ( n281964 , n268195 , n281963 , n259847 );
nand ( n281965 , n256292 , n32539 );
nand ( n281966 , n281962 , n281964 , n281965 );
buf ( n281967 , n281966 );
nand ( n281968 , n273013 , n262201 );
not ( n281969 , n238110 );
or ( n281970 , n281968 , n281969 );
not ( n281971 , n238109 );
not ( n281972 , n281971 );
not ( n281973 , n273013 );
or ( n281974 , n281972 , n281973 );
nor ( n281975 , n262201 , n252872 );
nand ( n281976 , n281974 , n281975 );
nand ( n281977 , n41945 , n38871 );
nand ( n281978 , n281970 , n281976 , n281977 );
buf ( n281979 , n281978 );
not ( n281980 , n276256 );
nand ( n281981 , n276243 , n269990 );
or ( n281982 , n281980 , n281981 );
not ( n281983 , n276243 );
not ( n281984 , n269964 );
or ( n281985 , n281983 , n281984 );
nor ( n281986 , n269990 , n239237 );
nand ( n281987 , n281985 , n281986 );
nand ( n281988 , n35431 , n33334 );
nand ( n281989 , n281982 , n281987 , n281988 );
buf ( n281990 , n281989 );
not ( n281991 , n273755 );
nand ( n281992 , n281991 , n258527 );
or ( n281993 , n273757 , n281992 );
not ( n281994 , n281991 );
not ( n281995 , n258455 );
or ( n281996 , n281994 , n281995 );
nor ( n281997 , n258527 , n251361 );
nand ( n281998 , n281996 , n281997 );
nand ( n281999 , n35431 , n36234 );
nand ( n282000 , n281993 , n281998 , n281999 );
buf ( n282001 , n282000 );
or ( n282002 , n25328 , n268955 );
or ( n282003 , n25335 , n280772 );
nand ( n282004 , n282002 , n282003 );
buf ( n282005 , n282004 );
not ( n282006 , RI19aa8530_2507);
or ( n282007 , n233507 , n282006 );
not ( n282008 , RI19a9ed50_2578);
or ( n282009 , n25335 , n282008 );
nand ( n282010 , n282007 , n282009 );
buf ( n282011 , n282010 );
not ( n282012 , n33822 );
not ( n282013 , n51381 );
or ( n282014 , n282012 , n282013 );
nand ( n282015 , n265694 , n259607 );
and ( n282016 , n282015 , n277902 );
not ( n282017 , n282015 );
and ( n282018 , n282017 , n277903 );
nor ( n282019 , n282016 , n282018 );
or ( n282020 , n282019 , n253358 );
nand ( n282021 , n282014 , n282020 );
buf ( n282022 , n282021 );
not ( n282023 , RI19a94940_2650);
or ( n282024 , n25328 , n282023 );
not ( n282025 , RI19a8aad0_2720);
or ( n282026 , n226822 , n282025 );
nand ( n282027 , n282024 , n282026 );
buf ( n282028 , n282027 );
nand ( n282029 , n268622 , n276703 );
or ( n282030 , n281713 , n282029 );
not ( n282031 , n276703 );
not ( n282032 , n276690 );
or ( n282033 , n282031 , n282032 );
nand ( n282034 , n282033 , n268623 );
nand ( n282035 , n31577 , n35242 );
nand ( n282036 , n282030 , n282034 , n282035 );
buf ( n282037 , n282036 );
nand ( n282038 , n251547 , n254528 );
nand ( n282039 , n271112 , n257334 );
or ( n282040 , n282038 , n282039 );
not ( n282041 , n257334 );
not ( n282042 , n251547 );
or ( n282043 , n282041 , n282042 );
nor ( n282044 , n271112 , n55104 );
nand ( n282045 , n282043 , n282044 );
nand ( n282046 , n247585 , n44391 );
nand ( n282047 , n282040 , n282045 , n282046 );
buf ( n282048 , n282047 );
buf ( n282049 , n32946 );
not ( n282050 , n256436 );
not ( n282051 , n256451 );
or ( n282052 , n282050 , n282051 );
nor ( n282053 , n281226 , n33253 );
nand ( n282054 , n282052 , n282053 );
nand ( n282055 , n261637 , n281226 , n256451 );
nand ( n282056 , n261585 , n220535 );
nand ( n282057 , n282054 , n282055 , n282056 );
buf ( n282058 , n282057 );
buf ( n282059 , n39233 );
not ( n282060 , n259871 );
not ( n282061 , n282060 );
not ( n282062 , n259860 );
or ( n282063 , n282061 , n282062 );
nor ( n282064 , n261278 , n250431 );
nand ( n282065 , n282063 , n282064 );
nand ( n282066 , n259860 , n269881 , n261278 );
nand ( n282067 , n256292 , n27833 );
nand ( n282068 , n282065 , n282066 , n282067 );
buf ( n282069 , n282068 );
buf ( n282070 , n37099 );
buf ( n282071 , n28810 );
buf ( n282072 , n26197 );
buf ( n282073 , n32841 );
buf ( n282074 , n228982 );
buf ( n282075 , n35377 );
not ( n282076 , n40888 );
not ( n282077 , n51381 );
or ( n282078 , n282076 , n282077 );
nand ( n282079 , n280647 , n280657 );
not ( n282080 , n263489 );
and ( n282081 , n282079 , n282080 );
not ( n282082 , n282079 );
and ( n282083 , n282082 , n263489 );
nor ( n282084 , n282081 , n282083 );
or ( n282085 , n282084 , n256214 );
nand ( n282086 , n282078 , n282085 );
buf ( n282087 , n282086 );
buf ( n282088 , RI19a247d0_2785);
not ( n282089 , n282088 );
not ( n282090 , n257347 );
or ( n282091 , n282089 , n282090 );
nand ( n282092 , n257351 , n276426 );
nand ( n282093 , n282091 , n282092 );
buf ( n282094 , n282093 );
buf ( n282095 , n27712 );
buf ( n282096 , n38903 );
buf ( n282097 , n210118 );
nand ( n282098 , n280644 , n258918 );
nand ( n282099 , n263499 , n280658 );
or ( n282100 , n282098 , n282099 );
not ( n282101 , n263499 );
not ( n282102 , n280644 );
or ( n282103 , n282101 , n282102 );
nor ( n282104 , n280658 , n49959 );
nand ( n282105 , n282103 , n282104 );
nand ( n282106 , n35431 , n40045 );
nand ( n282107 , n282100 , n282105 , n282106 );
buf ( n282108 , n282107 );
or ( n282109 , n233507 , n261015 );
not ( n282110 , RI19a8efb8_2690);
or ( n282111 , n25335 , n282110 );
nand ( n282112 , n282109 , n282111 );
buf ( n282113 , n282112 );
xor ( n282114 , n51740 , n267305 );
xnor ( n282115 , n282114 , n260340 );
not ( n282116 , n282115 );
nand ( n282117 , n282116 , n241373 );
not ( n282118 , n247155 );
not ( n282119 , n253474 );
or ( n282120 , n282118 , n282119 );
not ( n282121 , n247155 );
nand ( n282122 , n282121 , n248276 );
nand ( n282123 , n282120 , n282122 );
and ( n282124 , n282123 , n248284 );
not ( n282125 , n282123 );
and ( n282126 , n282125 , n248281 );
nor ( n282127 , n282124 , n282126 );
not ( n282128 , n243660 );
not ( n282129 , n54145 );
not ( n282130 , n282129 );
not ( n282131 , n242380 );
or ( n282132 , n282130 , n282131 );
nand ( n282133 , n242373 , n54145 );
nand ( n282134 , n282132 , n282133 );
not ( n282135 , n282134 );
or ( n282136 , n282128 , n282135 );
or ( n282137 , n282134 , n243660 );
nand ( n282138 , n282136 , n282137 );
not ( n282139 , n282138 );
nand ( n282140 , n282127 , n282139 );
or ( n282141 , n282117 , n282140 );
not ( n282142 , n282139 );
not ( n282143 , n282116 );
or ( n282144 , n282142 , n282143 );
nor ( n282145 , n282127 , n254740 );
nand ( n282146 , n282144 , n282145 );
nand ( n282147 , n39767 , n39943 );
nand ( n282148 , n282141 , n282146 , n282147 );
buf ( n282149 , n282148 );
nand ( n282150 , n270412 , n244378 );
or ( n282151 , n249010 , n282150 );
nor ( n282152 , n249008 , n235895 );
nand ( n282153 , n282152 , n282150 );
nand ( n282154 , n35431 , n28630 );
nand ( n282155 , n282151 , n282153 , n282154 );
buf ( n282156 , n282155 );
nor ( n282157 , n254769 , n257168 );
nand ( n282158 , n263249 , n282157 );
not ( n282159 , n257169 );
not ( n282160 , n254757 );
or ( n282161 , n282159 , n282160 );
nor ( n282162 , n254770 , n35428 );
nand ( n282163 , n282161 , n282162 );
nand ( n282164 , n237361 , n29236 );
nand ( n282165 , n282158 , n282163 , n282164 );
buf ( n282166 , n282165 );
not ( n282167 , RI19aa8f80_2503);
or ( n282168 , n25328 , n282167 );
or ( n282169 , n25335 , n274923 );
nand ( n282170 , n282168 , n282169 );
buf ( n282171 , n282170 );
or ( n282172 , n25328 , n254187 );
or ( n282173 , n25335 , n262587 );
nand ( n282174 , n282172 , n282173 );
buf ( n282175 , n282174 );
not ( n282176 , RI19a9d9a0_2587);
or ( n282177 , n25328 , n282176 );
or ( n282178 , n25335 , n234028 );
nand ( n282179 , n282177 , n282178 );
buf ( n282180 , n282179 );
nand ( n282181 , n259123 , n241459 );
nand ( n282182 , n266883 , n261112 );
or ( n282183 , n282181 , n282182 );
not ( n282184 , n266883 );
not ( n282185 , n259123 );
or ( n282186 , n282184 , n282185 );
nor ( n282187 , n261112 , n55152 );
nand ( n282188 , n282186 , n282187 );
nand ( n282189 , n31577 , n33393 );
nand ( n282190 , n282183 , n282188 , n282189 );
buf ( n282191 , n282190 );
not ( n282192 , n29277 );
not ( n282193 , n245943 );
or ( n282194 , n282192 , n282193 );
nand ( n282195 , n254896 , n257089 );
and ( n282196 , n282195 , n261918 );
not ( n282197 , n282195 );
and ( n282198 , n282197 , n261919 );
nor ( n282199 , n282196 , n282198 );
or ( n282200 , n282199 , n258327 );
nand ( n282201 , n282194 , n282200 );
buf ( n282202 , n282201 );
nand ( n282203 , n272772 , n263313 );
not ( n282204 , n278401 );
or ( n282205 , n282203 , n282204 );
not ( n282206 , n272766 );
not ( n282207 , n272772 );
or ( n282208 , n282206 , n282207 );
nor ( n282209 , n263313 , n38637 );
nand ( n282210 , n282208 , n282209 );
nand ( n282211 , n246217 , n204411 );
nand ( n282212 , n282205 , n282210 , n282211 );
buf ( n282213 , n282212 );
not ( n282214 , n258896 );
not ( n282215 , n251173 );
not ( n282216 , n282215 );
or ( n282217 , n282214 , n282216 );
nor ( n282218 , n281113 , n264469 );
nand ( n282219 , n282217 , n282218 );
nand ( n282220 , n258898 , n282215 , n281113 );
nand ( n282221 , n241378 , n206978 );
nand ( n282222 , n282219 , n282220 , n282221 );
buf ( n282223 , n282222 );
not ( n282224 , n269426 );
nor ( n282225 , n282224 , n269436 );
nand ( n282226 , n271515 , n282225 );
not ( n282227 , n269436 );
not ( n282228 , n282227 );
not ( n282229 , n271517 );
or ( n282230 , n282228 , n282229 );
nor ( n282231 , n269426 , n49959 );
nand ( n282232 , n282230 , n282231 );
nand ( n282233 , n238114 , n55544 );
nand ( n282234 , n282226 , n282232 , n282233 );
buf ( n282235 , n282234 );
not ( n282236 , n33728 );
not ( n282237 , n50615 );
or ( n282238 , n282236 , n282237 );
not ( n282239 , n259860 );
nand ( n282240 , n282239 , n261278 );
and ( n282241 , n282240 , n261266 );
not ( n282242 , n282240 );
not ( n282243 , n261266 );
and ( n282244 , n282242 , n282243 );
nor ( n282245 , n282241 , n282244 );
or ( n282246 , n282245 , n245938 );
nand ( n282247 , n282238 , n282246 );
buf ( n282248 , n282247 );
or ( n282249 , n25328 , n277202 );
not ( n282250 , RI19a91358_2674);
or ( n282251 , n226822 , n282250 );
nand ( n282252 , n282249 , n282251 );
buf ( n282253 , n282252 );
not ( n282254 , n278873 );
or ( n282255 , n260497 , n282254 );
not ( n282256 , n278874 );
not ( n282257 , n260561 );
and ( n282258 , n282256 , n282257 );
and ( n282259 , n224937 , n31753 );
nor ( n282260 , n282258 , n282259 );
nor ( n282261 , n260560 , n278873 );
nand ( n282262 , n280781 , n282261 );
nand ( n282263 , n282255 , n282260 , n282262 );
buf ( n282264 , n282263 );
not ( n282265 , n278177 );
not ( n282266 , n273599 );
and ( n282267 , n282265 , n282266 );
and ( n282268 , n237361 , n30241 );
nor ( n282269 , n282267 , n282268 );
not ( n282270 , n257760 );
nand ( n282271 , n282270 , n278176 );
nand ( n282272 , n257762 , n273599 , n280484 );
nand ( n282273 , n282269 , n282271 , n282272 );
buf ( n282274 , n282273 );
not ( n282275 , n234856 );
not ( n282276 , n225525 );
or ( n282277 , n282275 , n282276 );
not ( n282278 , n234856 );
nand ( n282279 , n282278 , n47773 );
nand ( n282280 , n282277 , n282279 );
and ( n282281 , n282280 , n234437 );
not ( n282282 , n282280 );
and ( n282283 , n282282 , n246207 );
nor ( n282284 , n282281 , n282283 );
not ( n282285 , n282284 );
not ( n282286 , n282285 );
not ( n282287 , n268306 );
or ( n282288 , n282286 , n282287 );
nor ( n282289 , n268317 , n47173 );
nand ( n282290 , n282288 , n282289 );
nor ( n282291 , n282284 , n49051 );
nand ( n282292 , n268306 , n282291 , n268317 );
nand ( n282293 , n256292 , n36128 );
nand ( n282294 , n282290 , n282292 , n282293 );
buf ( n282295 , n282294 );
nand ( n282296 , n258127 , n279056 );
or ( n282297 , n282296 , n240158 );
nor ( n282298 , n240157 , n252070 );
nand ( n282299 , n282298 , n282296 );
nand ( n282300 , n41945 , n205232 );
nand ( n282301 , n282297 , n282299 , n282300 );
buf ( n282302 , n282301 );
not ( n282303 , n255502 );
nand ( n282304 , n282303 , n255528 );
nor ( n282305 , n267721 , n243434 );
not ( n282306 , n282305 );
or ( n282307 , n282304 , n282306 );
not ( n282308 , n254227 );
not ( n282309 , n267721 );
nor ( n282310 , n282308 , n282309 );
nand ( n282311 , n282304 , n282310 );
nand ( n282312 , n31577 , n31875 );
nand ( n282313 , n282307 , n282311 , n282312 );
buf ( n282314 , n282313 );
nand ( n282315 , n247715 , n272079 );
not ( n282316 , n247699 );
or ( n282317 , n282315 , n282316 );
nand ( n282318 , n282315 , n271692 );
nand ( n282319 , n39766 , n34162 );
nand ( n282320 , n282317 , n282318 , n282319 );
buf ( n282321 , n282320 );
buf ( n282322 , n30133 );
buf ( n282323 , n205718 );
not ( n282324 , n36907 );
not ( n282325 , n255116 );
or ( n282326 , n282324 , n282325 );
nand ( n282327 , n268622 , n276702 );
and ( n282328 , n282327 , n268646 );
not ( n282329 , n282327 );
and ( n282330 , n282329 , n268645 );
nor ( n282331 , n282328 , n282330 );
or ( n282332 , n282331 , n39763 );
nand ( n282333 , n282326 , n282332 );
buf ( n282334 , n282333 );
buf ( n282335 , n31161 );
buf ( n282336 , n232391 );
not ( n282337 , RI1754b170_46);
or ( n282338 , n249126 , n282337 );
nand ( n282339 , n244606 , n25377 );
nand ( n282340 , n282338 , n282339 );
buf ( n282341 , n282340 );
nand ( n282342 , n265846 , n278513 );
or ( n282343 , n268739 , n282342 );
not ( n282344 , n265835 );
not ( n282345 , n265846 );
or ( n282346 , n282344 , n282345 );
nor ( n282347 , n278513 , n236795 );
nand ( n282348 , n282346 , n282347 );
nand ( n282349 , n35431 , n232391 );
nand ( n282350 , n282343 , n282348 , n282349 );
buf ( n282351 , n282350 );
not ( n282352 , n272141 );
nor ( n282353 , n275264 , n235050 );
nand ( n282354 , n282352 , n282353 , n275254 );
not ( n282355 , n275264 );
nand ( n282356 , n275254 , n282355 );
nand ( n282357 , n282356 , n272141 , n205649 );
nand ( n282358 , n31577 , n204556 );
nand ( n282359 , n282354 , n282357 , n282358 );
buf ( n282360 , n282359 );
not ( n282361 , n275823 );
not ( n282362 , n263106 );
or ( n282363 , n282361 , n282362 );
nor ( n282364 , n263131 , n52445 );
nand ( n282365 , n282363 , n282364 );
nand ( n282366 , n280011 , n263106 , n263131 );
nand ( n282367 , n237714 , n29112 );
nand ( n282368 , n282365 , n282366 , n282367 );
buf ( n282369 , n282368 );
not ( n282370 , n276453 );
nand ( n282371 , n282370 , n278699 );
or ( n282372 , n267960 , n282371 );
nand ( n282373 , n273914 , n282371 );
nand ( n282374 , n255116 , n29887 );
nand ( n282375 , n282372 , n282373 , n282374 );
buf ( n282376 , n282375 );
not ( n282377 , n252054 );
not ( n282378 , n264103 );
nand ( n282379 , n282377 , n282378 );
not ( n282380 , n252071 );
or ( n282381 , n282379 , n282380 );
nor ( n282382 , n251980 , n252070 );
nand ( n282383 , n282379 , n282382 );
nand ( n282384 , n31577 , n28470 );
nand ( n282385 , n282381 , n282383 , n282384 );
buf ( n282386 , n282385 );
nand ( n282387 , n257286 , n264375 , n257272 );
nand ( n282388 , n257272 , n257289 );
not ( n282389 , n264375 );
nand ( n282390 , n282388 , n282389 , n254227 );
nand ( n282391 , n35431 , n31633 );
nand ( n282392 , n282387 , n282390 , n282391 );
buf ( n282393 , n282392 );
not ( n282394 , RI1754aae0_60);
or ( n282395 , n249125 , n282394 );
or ( n282396 , n25335 , n281848 );
nand ( n282397 , n282395 , n282396 );
buf ( n282398 , n282397 );
not ( n282399 , n31368 );
not ( n282400 , n244606 );
or ( n282401 , n282399 , n282400 );
not ( n282402 , RI1754acc0_56);
or ( n282403 , n269544 , n282402 );
nand ( n282404 , n282401 , n282403 );
buf ( n282405 , n282404 );
buf ( n282406 , n28446 );
buf ( n282407 , n209468 );
not ( n282408 , n270495 );
not ( n282409 , n270663 );
or ( n282410 , n282408 , n282409 );
nor ( n282411 , n263418 , n247698 );
nand ( n282412 , n282410 , n282411 );
nand ( n282413 , n270499 , n270663 , n263418 );
nand ( n282414 , n35431 , n36050 );
nand ( n282415 , n282412 , n282413 , n282414 );
buf ( n282416 , n282415 );
or ( n282417 , n25328 , n278614 );
or ( n282418 , n25335 , n274917 );
nand ( n282419 , n282417 , n282418 );
buf ( n282420 , n282419 );
not ( n282421 , RI19ab2508_2437);
or ( n282422 , n25328 , n282421 );
or ( n282423 , n25335 , n252364 );
nand ( n282424 , n282422 , n282423 );
buf ( n282425 , n282424 );
nand ( n282426 , n258875 , n277399 );
nand ( n282427 , n282426 , n273677 , n33255 );
nand ( n282428 , n277409 , n273678 , n258875 );
nand ( n282429 , n37728 , n205289 );
nand ( n282430 , n282427 , n282428 , n282429 );
buf ( n282431 , n282430 );
not ( n282432 , n32574 );
not ( n282433 , n263819 );
or ( n282434 , n282432 , n282433 );
not ( n282435 , n264113 );
nand ( n282436 , n282435 , n264103 );
and ( n282437 , n282436 , n252054 );
not ( n282438 , n282436 );
and ( n282439 , n282438 , n282377 );
nor ( n282440 , n282437 , n282439 );
or ( n282441 , n282440 , n238223 );
nand ( n282442 , n282434 , n282441 );
buf ( n282443 , n282442 );
not ( n282444 , n41136 );
not ( n282445 , n245702 );
or ( n282446 , n282444 , n282445 );
nand ( n282447 , n278512 , n268737 );
and ( n282448 , n282447 , n265858 );
not ( n282449 , n282447 );
and ( n282450 , n282449 , n265859 );
nor ( n282451 , n282448 , n282450 );
or ( n282452 , n282451 , n257174 );
nand ( n282453 , n282446 , n282452 );
buf ( n282454 , n282453 );
not ( n282455 , RI19acaf40_2248);
or ( n282456 , n25328 , n282455 );
or ( n282457 , n25336 , n278988 );
nand ( n282458 , n282456 , n282457 );
buf ( n282459 , n282458 );
or ( n282460 , n25328 , n271319 );
not ( n282461 , RI19a8faf8_2685);
or ( n282462 , n226822 , n282461 );
nand ( n282463 , n282460 , n282462 );
buf ( n282464 , n282463 );
buf ( n282465 , n204575 );
buf ( n282466 , n204419 );
not ( n282467 , n274493 );
not ( n282468 , n274490 );
or ( n282469 , n282467 , n282468 );
nor ( n282470 , n254815 , n251361 );
nand ( n282471 , n282469 , n282470 );
nand ( n282472 , n277572 , n254815 , n274490 );
nand ( n282473 , n237714 , n31838 );
nand ( n282474 , n282471 , n282472 , n282473 );
buf ( n282475 , n282474 );
buf ( n282476 , n40038 );
buf ( n282477 , n32191 );
nand ( n282478 , n264925 , n243233 );
nand ( n282479 , n273051 , n264947 );
or ( n282480 , n282478 , n282479 );
not ( n282481 , n264925 );
not ( n282482 , n264947 );
or ( n282483 , n282481 , n282482 );
nor ( n282484 , n273051 , n37725 );
nand ( n282485 , n282483 , n282484 );
nand ( n282486 , n39767 , n205117 );
nand ( n282487 , n282480 , n282485 , n282486 );
buf ( n282488 , n282487 );
not ( n282489 , n250425 );
nand ( n282490 , n282489 , n276624 );
or ( n282491 , n269166 , n282490 );
not ( n282492 , n269165 );
not ( n282493 , n282489 );
or ( n282494 , n282492 , n282493 );
nor ( n282495 , n276624 , n40465 );
nand ( n282496 , n282494 , n282495 );
nand ( n282497 , n234024 , n31657 );
nand ( n282498 , n282491 , n282496 , n282497 );
buf ( n282499 , n282498 );
not ( n282500 , RI19acbe40_2240);
or ( n282501 , n25328 , n282500 );
or ( n282502 , n25336 , n269997 );
nand ( n282503 , n282501 , n282502 );
buf ( n282504 , n282503 );
or ( n282505 , n25328 , n278975 );
or ( n282506 , n25336 , n277497 );
nand ( n282507 , n282505 , n282506 );
buf ( n282508 , n282507 );
nand ( n282509 , n281150 , n248151 , n250277 );
nand ( n282510 , n250258 , n250277 );
nand ( n282511 , n282510 , n248152 , n254528 );
nand ( n282512 , n245414 , n34696 );
nand ( n282513 , n282509 , n282511 , n282512 );
buf ( n282514 , n282513 );
not ( n282515 , n55152 );
nand ( n282516 , n282515 , n247238 );
nand ( n282517 , n262108 , n262119 );
or ( n282518 , n282516 , n282517 );
not ( n282519 , n262108 );
not ( n282520 , n247238 );
or ( n282521 , n282519 , n282520 );
nor ( n282522 , n262119 , n55146 );
nand ( n282523 , n282521 , n282522 );
nand ( n282524 , n31577 , n54785 );
nand ( n282525 , n282518 , n282523 , n282524 );
buf ( n282526 , n282525 );
not ( n282527 , n53331 );
not ( n282528 , n250359 );
or ( n282529 , n282527 , n282528 );
not ( n282530 , n53331 );
nand ( n282531 , n282530 , n250366 );
nand ( n282532 , n282529 , n282531 );
and ( n282533 , n282532 , n250374 );
not ( n282534 , n282532 );
and ( n282535 , n282534 , n250371 );
nor ( n282536 , n282533 , n282535 );
not ( n282537 , n282536 );
nand ( n282538 , n282537 , n35420 );
or ( n282539 , n33256 , n282538 );
nor ( n282540 , n33251 , n35427 );
nand ( n282541 , n282540 , n282538 );
nand ( n282542 , n51381 , n28313 );
nand ( n282543 , n282539 , n282541 , n282542 );
buf ( n282544 , n282543 );
nand ( n282545 , n260630 , n260658 );
or ( n282546 , n278532 , n282545 );
not ( n282547 , n260630 );
not ( n282548 , n278531 );
or ( n282549 , n282547 , n282548 );
nor ( n282550 , n260658 , n236795 );
nand ( n282551 , n282549 , n282550 );
nand ( n282552 , n234448 , n35866 );
nand ( n282553 , n282546 , n282551 , n282552 );
buf ( n282554 , n282553 );
buf ( n282555 , RI17536d88_596);
and ( n282556 , n27883 , n282555 );
buf ( n282557 , n282556 );
nand ( n282558 , n278207 , n268085 );
or ( n282559 , n279863 , n282558 );
not ( n282560 , n278207 );
not ( n282561 , n279862 );
or ( n282562 , n282560 , n282561 );
nor ( n282563 , n268085 , n46425 );
nand ( n282564 , n282562 , n282563 );
nand ( n282565 , n238638 , n35501 );
nand ( n282566 , n282559 , n282564 , n282565 );
buf ( n282567 , n282566 );
buf ( n282568 , n204797 );
buf ( n282569 , n204368 );
buf ( n282570 , n28303 );
buf ( n282571 , n25843 );
not ( n282572 , n278272 );
nand ( n282573 , n282572 , n273303 );
not ( n282574 , n282573 );
or ( n282575 , n275424 , n282574 );
or ( n282576 , n273293 , n282573 );
nand ( n282577 , n239240 , n26480 );
nand ( n282578 , n282575 , n282576 , n282577 );
buf ( n282579 , n282578 );
or ( n282580 , n25328 , n281541 );
or ( n282581 , n25335 , n264359 );
nand ( n282582 , n282580 , n282581 );
buf ( n282583 , n282582 );
nor ( n282584 , n271619 , n275706 );
or ( n282585 , n247416 , n282584 );
nand ( n282586 , n271626 , n282584 );
nand ( n282587 , n39766 , n39771 );
nand ( n282588 , n282585 , n282586 , n282587 );
buf ( n282589 , n282588 );
nand ( n282590 , n280448 , n260930 );
nand ( n282591 , n267768 , n280460 );
or ( n282592 , n282590 , n282591 );
not ( n282593 , n280460 );
not ( n282594 , n280448 );
or ( n282595 , n282593 , n282594 );
nor ( n282596 , n267768 , n252258 );
nand ( n282597 , n282595 , n282596 );
nand ( n282598 , n244987 , n204734 );
nand ( n282599 , n282592 , n282597 , n282598 );
buf ( n282600 , n282599 );
not ( n282601 , n37596 );
not ( n282602 , n241068 );
or ( n282603 , n282601 , n282602 );
not ( n282604 , n263863 );
nand ( n282605 , n282604 , n263853 );
and ( n282606 , n282605 , n239659 );
not ( n282607 , n282605 );
and ( n282608 , n282607 , n239658 );
nor ( n282609 , n282606 , n282608 );
or ( n282610 , n282609 , n256376 );
nand ( n282611 , n282603 , n282610 );
buf ( n282612 , n282611 );
nand ( n282613 , n265273 , n257792 );
nand ( n282614 , n258298 , n265288 );
or ( n282615 , n282613 , n282614 );
not ( n282616 , n265288 );
not ( n282617 , n265273 );
or ( n282618 , n282616 , n282617 );
nor ( n282619 , n258298 , n235050 );
nand ( n282620 , n282618 , n282619 );
nand ( n282621 , n237361 , n220347 );
nand ( n282622 , n282615 , n282620 , n282621 );
buf ( n282623 , n282622 );
buf ( n282624 , n36836 );
or ( n282625 , n25328 , n280566 );
or ( n282626 , n25335 , n265141 );
nand ( n282627 , n282625 , n282626 );
buf ( n282628 , n282627 );
nor ( n282629 , n259664 , n259676 );
nand ( n282630 , n259411 , n282629 );
nand ( n282631 , n259404 , n259675 );
nand ( n282632 , n282631 , n259664 , n233973 );
nand ( n282633 , n256292 , n32418 );
nand ( n282634 , n282630 , n282632 , n282633 );
buf ( n282635 , n282634 );
nand ( n282636 , n272376 , n269751 );
or ( n282637 , n272366 , n282636 );
nand ( n282638 , n272612 , n282636 );
nand ( n282639 , n41944 , n36973 );
nand ( n282640 , n282637 , n282638 , n282639 );
buf ( n282641 , n282640 );
nand ( n282642 , n279774 , n252773 , n252840 );
not ( n282643 , n274681 );
not ( n282644 , n282643 );
not ( n282645 , n252773 );
or ( n282646 , n282644 , n282645 );
nor ( n282647 , n252840 , n31572 );
nand ( n282648 , n282646 , n282647 );
nand ( n282649 , n238114 , n38995 );
nand ( n282650 , n282642 , n282648 , n282649 );
buf ( n282651 , n282650 );
not ( n282652 , n251979 );
not ( n282653 , n252067 );
or ( n282654 , n282652 , n282653 );
nor ( n282655 , n264113 , n258327 );
nand ( n282656 , n282654 , n282655 );
nand ( n282657 , n282382 , n252067 , n264113 );
nand ( n282658 , n37728 , n35831 );
nand ( n282659 , n282656 , n282657 , n282658 );
buf ( n282660 , n282659 );
not ( n282661 , n251858 );
nand ( n282662 , n282661 , n247444 );
nand ( n282663 , n273523 , n273511 );
or ( n282664 , n282662 , n282663 );
not ( n282665 , n273523 );
not ( n282666 , n282661 );
or ( n282667 , n282665 , n282666 );
nor ( n282668 , n273511 , n234110 );
nand ( n282669 , n282667 , n282668 );
nand ( n282670 , n252711 , n26177 );
nand ( n282671 , n282664 , n282669 , n282670 );
buf ( n282672 , n282671 );
not ( n282673 , n268437 );
nand ( n282674 , n282673 , n245241 );
nand ( n282675 , n279526 , n268439 );
or ( n282676 , n282674 , n282675 );
not ( n282677 , n279526 );
not ( n282678 , n282673 );
or ( n282679 , n282677 , n282678 );
nor ( n282680 , n268439 , n33253 );
nand ( n282681 , n282679 , n282680 );
nand ( n282682 , n247585 , n204833 );
nand ( n282683 , n282676 , n282681 , n282682 );
buf ( n282684 , n282683 );
not ( n282685 , RI1754a978_63);
or ( n282686 , n249125 , n282685 );
or ( n282687 , n25335 , n276962 );
nand ( n282688 , n282686 , n282687 );
buf ( n282689 , n282688 );
not ( n282690 , RI19a981f8_2625);
or ( n282691 , n25328 , n282690 );
or ( n282692 , n226822 , n241980 );
nand ( n282693 , n282691 , n282692 );
buf ( n282694 , n282693 );
buf ( n282695 , RI19ad1588_2202);
and ( n282696 , n25326 , n282695 );
buf ( n282697 , n282696 );
or ( n282698 , n25328 , n280774 );
not ( n282699 , RI19a8b250_2717);
or ( n282700 , n226822 , n282699 );
nand ( n282701 , n282698 , n282700 );
buf ( n282702 , n282701 );
nand ( n282703 , n282284 , n280140 );
or ( n282704 , n268330 , n282703 );
not ( n282705 , n280140 );
not ( n282706 , n268329 );
or ( n282707 , n282705 , n282706 );
nand ( n282708 , n282707 , n282291 );
nand ( n282709 , n49054 , n37244 );
nand ( n282710 , n282704 , n282708 , n282709 );
buf ( n282711 , n282710 );
nand ( n282712 , n280923 , n256751 );
not ( n282713 , n280919 );
nand ( n282714 , n282713 , n273634 );
or ( n282715 , n282712 , n282714 );
not ( n282716 , n282713 );
not ( n282717 , n280923 );
or ( n282718 , n282716 , n282717 );
nand ( n282719 , n282718 , n273635 );
nand ( n282720 , n256292 , n40103 );
nand ( n282721 , n282715 , n282719 , n282720 );
buf ( n282722 , n282721 );
not ( n282723 , n280628 );
not ( n282724 , n265651 );
nand ( n282725 , n282724 , n265628 );
or ( n282726 , n282723 , n282725 );
nor ( n282727 , n280624 , n255533 );
nand ( n282728 , n282727 , n282725 );
nand ( n282729 , n258213 , n33548 );
nand ( n282730 , n282726 , n282728 , n282729 );
buf ( n282731 , n282730 );
nor ( n282732 , n280942 , n52445 );
nor ( n282733 , n260256 , n259760 );
nand ( n282734 , n282732 , n282733 );
nor ( n282735 , n280944 , n255014 );
not ( n282736 , n280942 );
nand ( n282737 , n282736 , n259757 );
nand ( n282738 , n282735 , n282737 );
nand ( n282739 , n245414 , n33751 );
nand ( n282740 , n282734 , n282738 , n282739 );
buf ( n282741 , n282740 );
or ( n282742 , n25328 , n281298 );
or ( n282743 , n25335 , n259041 );
nand ( n282744 , n282742 , n282743 );
buf ( n282745 , n282744 );
not ( n282746 , n271480 );
nor ( n282747 , n282746 , n281590 );
nand ( n282748 , n273982 , n282747 );
not ( n282749 , n281590 );
nand ( n282750 , n273975 , n282749 );
nand ( n282751 , n282750 , n282746 , n254013 );
nand ( n282752 , n31577 , n35662 );
nand ( n282753 , n282748 , n282751 , n282752 );
buf ( n282754 , n282753 );
buf ( n282755 , n36646 );
buf ( n282756 , n37642 );
buf ( n282757 , n204787 );
or ( n282758 , n25328 , n242605 );
or ( n282759 , n25335 , n278630 );
nand ( n282760 , n282758 , n282759 );
buf ( n282761 , n282760 );
nor ( n282762 , n233999 , n272592 );
nand ( n282763 , n272595 , n282762 );
not ( n282764 , n234017 );
not ( n282765 , n272592 );
not ( n282766 , n282765 );
or ( n282767 , n282764 , n282766 );
not ( n282768 , n233999 );
nor ( n282769 , n282768 , n43517 );
nand ( n282770 , n282767 , n282769 );
nand ( n282771 , n239240 , n35842 );
nand ( n282772 , n282763 , n282770 , n282771 );
buf ( n282773 , n282772 );
nand ( n282774 , n278784 , n254013 );
nand ( n282775 , n234540 , n278788 );
or ( n282776 , n282774 , n282775 );
not ( n282777 , n278788 );
not ( n282778 , n278784 );
or ( n282779 , n282777 , n282778 );
nor ( n282780 , n234540 , n234110 );
nand ( n282781 , n282779 , n282780 );
nand ( n282782 , n31576 , n25755 );
nand ( n282783 , n282776 , n282781 , n282782 );
buf ( n282784 , n282783 );
nor ( n282785 , n280525 , n234021 );
nor ( n282786 , n262169 , n267230 );
nand ( n282787 , n282785 , n282786 );
not ( n282788 , n280524 );
not ( n282789 , n280529 );
or ( n282790 , n282788 , n282789 );
nor ( n282791 , n267220 , n219702 );
nand ( n282792 , n282790 , n282791 );
nand ( n282793 , n256673 , n42942 );
nand ( n282794 , n282787 , n282792 , n282793 );
buf ( n282795 , n282794 );
nand ( n282796 , n267824 , n263343 , n277214 );
not ( n282797 , n267827 );
not ( n282798 , n263343 );
or ( n282799 , n282797 , n282798 );
nor ( n282800 , n277214 , n37724 );
nand ( n282801 , n282799 , n282800 );
nand ( n282802 , n35431 , n205277 );
nand ( n282803 , n282796 , n282801 , n282802 );
buf ( n282804 , n282803 );
not ( n282805 , n232141 );
not ( n282806 , n237361 );
or ( n282807 , n282805 , n282806 );
nand ( n282808 , n274254 , n268416 );
and ( n282809 , n282808 , n268409 );
not ( n282810 , n282808 );
not ( n282811 , n268409 );
and ( n282812 , n282810 , n282811 );
nor ( n282813 , n282809 , n282812 );
or ( n282814 , n282813 , n245938 );
nand ( n282815 , n282807 , n282814 );
buf ( n282816 , n282815 );
not ( n282817 , RI1754b620_36);
or ( n282818 , n249128 , n282817 );
nand ( n282819 , n249131 , n33918 );
nand ( n282820 , n282818 , n282819 );
buf ( n282821 , n282820 );
not ( n282822 , RI1754bd28_21);
or ( n282823 , n255977 , n282822 );
nand ( n282824 , n258185 , n30303 );
nand ( n282825 , n282823 , n282824 );
buf ( n282826 , n282825 );
buf ( n282827 , n26469 );
buf ( n282828 , n204432 );
buf ( n282829 , n32438 );
nand ( n282830 , n251093 , n266599 , n243963 );
not ( n282831 , n251097 );
not ( n282832 , n266599 );
or ( n282833 , n282831 , n282832 );
nor ( n282834 , n243963 , n252070 );
nand ( n282835 , n282833 , n282834 );
nand ( n282836 , n251717 , n37394 );
nand ( n282837 , n282830 , n282835 , n282836 );
buf ( n282838 , n282837 );
not ( n282839 , n29622 );
not ( n282840 , n233501 );
or ( n282841 , n282839 , n282840 );
nand ( n282842 , n280761 , n236791 );
and ( n282843 , n282842 , n279881 );
not ( n282844 , n282842 );
and ( n282845 , n282844 , n280766 );
nor ( n282846 , n282843 , n282845 );
or ( n282847 , n282846 , n257851 );
nand ( n282848 , n282841 , n282847 );
buf ( n282849 , n282848 );
nand ( n282850 , n260229 , n246019 );
or ( n282851 , n260219 , n282850 );
nand ( n282852 , n282850 , n276508 );
nand ( n282853 , n241068 , n33026 );
nand ( n282854 , n282851 , n282852 , n282853 );
buf ( n282855 , n282854 );
nand ( n282856 , n234308 , n255152 );
nand ( n282857 , n256046 , n277343 );
or ( n282858 , n282856 , n282857 );
not ( n282859 , n277343 );
not ( n282860 , n234308 );
or ( n282861 , n282859 , n282860 );
nor ( n282862 , n256046 , n40465 );
nand ( n282863 , n282861 , n282862 );
nand ( n282864 , n238638 , n28888 );
nand ( n282865 , n282858 , n282863 , n282864 );
buf ( n282866 , n282865 );
buf ( n282867 , n36344 );
buf ( n282868 , n25707 );
buf ( n282869 , n30388 );
nand ( n282870 , n279939 , n265793 );
nor ( n282871 , n270864 , n43968 );
not ( n282872 , n282871 );
or ( n282873 , n282870 , n282872 );
nand ( n282874 , n282870 , n270862 );
nand ( n282875 , n245414 , n33920 );
nand ( n282876 , n282873 , n282874 , n282875 );
buf ( n282877 , n282876 );
not ( n282878 , n273543 );
nand ( n282879 , n277133 , n270578 , n282878 );
not ( n282880 , n277136 );
not ( n282881 , n282878 );
or ( n282882 , n282880 , n282881 );
nor ( n282883 , n270578 , n53680 );
nand ( n282884 , n282882 , n282883 );
nand ( n282885 , n237714 , n31412 );
nand ( n282886 , n282879 , n282884 , n282885 );
buf ( n282887 , n282886 );
not ( n282888 , RI19abf870_2336);
or ( n282889 , n25328 , n282888 );
or ( n282890 , n25335 , n250975 );
nand ( n282891 , n282889 , n282890 );
buf ( n282892 , n282891 );
nand ( n282893 , n269779 , n258017 );
nand ( n282894 , n258003 , n38638 );
or ( n282895 , n282893 , n282894 );
not ( n282896 , n258003 );
not ( n282897 , n258017 );
or ( n282898 , n282896 , n282897 );
nor ( n282899 , n269779 , n43968 );
nand ( n282900 , n282898 , n282899 );
nand ( n282901 , n237361 , n33437 );
nand ( n282902 , n282895 , n282900 , n282901 );
buf ( n282903 , n282902 );
not ( n282904 , n33780 );
not ( n282905 , n251465 );
or ( n282906 , n282904 , n282905 );
nand ( n282907 , n243203 , n242980 );
and ( n282908 , n282907 , n257505 );
not ( n282909 , n282907 );
and ( n282910 , n282909 , n269844 );
nor ( n282911 , n282908 , n282910 );
or ( n282912 , n282911 , n244837 );
nand ( n282913 , n282906 , n282912 );
buf ( n282914 , n282913 );
or ( n282915 , n25328 , n275343 );
not ( n282916 , RI19ac34e8_2304);
or ( n282917 , n25335 , n282916 );
nand ( n282918 , n282915 , n282917 );
buf ( n282919 , n282918 );
nand ( n282920 , n263157 , n253397 );
nand ( n282921 , n250847 , n270306 );
or ( n282922 , n282920 , n282921 );
not ( n282923 , n270306 );
not ( n282924 , n263157 );
or ( n282925 , n282923 , n282924 );
nor ( n282926 , n250847 , n237384 );
nand ( n282927 , n282925 , n282926 );
nand ( n282928 , n236798 , n30300 );
nand ( n282929 , n282922 , n282927 , n282928 );
buf ( n282930 , n282929 );
nor ( n282931 , n35632 , n204520 , n272603 );
xor ( n282932 , n282931 , n266028 );
nand ( n282933 , n255104 , n255091 );
xnor ( n282934 , n282932 , n282933 );
or ( n282935 , n282934 , n235732 );
nand ( n282936 , n241378 , n204452 );
nand ( n282937 , n282935 , n282936 );
buf ( n282938 , n282937 );
or ( n282939 , n25328 , n274304 );
or ( n282940 , n25335 , n282455 );
nand ( n282941 , n282939 , n282940 );
buf ( n282942 , n282941 );
or ( n282943 , n25328 , n263196 );
not ( n282944 , RI19ac8768_2266);
or ( n282945 , n25336 , n282944 );
nand ( n282946 , n282943 , n282945 );
buf ( n282947 , n282946 );
or ( n282948 , n25328 , n272489 );
or ( n282949 , n25335 , n278795 );
nand ( n282950 , n282948 , n282949 );
buf ( n282951 , n282950 );
not ( n282952 , n267121 );
nand ( n282953 , n282952 , n226010 );
nand ( n282954 , n267132 , n274010 );
or ( n282955 , n282953 , n282954 );
not ( n282956 , n274010 );
not ( n282957 , n282952 );
or ( n282958 , n282956 , n282957 );
nor ( n282959 , n267132 , n46425 );
nand ( n282960 , n282958 , n282959 );
nand ( n282961 , n241976 , n204828 );
nand ( n282962 , n282955 , n282960 , n282961 );
buf ( n282963 , n282962 );
nand ( n282964 , n252382 , n278464 );
or ( n282965 , n277614 , n282964 );
not ( n282966 , n277613 );
not ( n282967 , n278464 );
or ( n282968 , n282966 , n282967 );
nor ( n282969 , n252382 , n242391 );
nand ( n282970 , n282968 , n282969 );
nand ( n282971 , n238638 , n40805 );
nand ( n282972 , n282965 , n282970 , n282971 );
buf ( n282973 , n282972 );
not ( n282974 , RI1754b9e0_28);
or ( n282975 , n229127 , n282974 );
not ( n282976 , RI19aa5a88_2525);
or ( n282977 , n25335 , n282976 );
nand ( n282978 , n282975 , n282977 );
buf ( n282979 , n282978 );
nand ( n282980 , n255817 , n222532 );
nand ( n282981 , n255895 , n258942 );
or ( n282982 , n282980 , n282981 );
not ( n282983 , n255817 );
not ( n282984 , n255895 );
or ( n282985 , n282983 , n282984 );
nor ( n282986 , n258942 , n235050 );
nand ( n282987 , n282985 , n282986 );
nand ( n282988 , n239240 , n53517 );
nand ( n282989 , n282982 , n282987 , n282988 );
buf ( n282990 , n282989 );
not ( n282991 , n253082 );
nand ( n282992 , n282991 , n280276 );
or ( n282993 , n253020 , n282992 );
not ( n282994 , n279188 );
nand ( n282995 , n282994 , n282992 );
nand ( n282996 , n31576 , n26289 );
nand ( n282997 , n282993 , n282995 , n282996 );
buf ( n282998 , n282997 );
not ( n282999 , RI1754bb48_25);
or ( n283000 , n255977 , n282999 );
nand ( n283001 , n258185 , n28758 );
nand ( n283002 , n283000 , n283001 );
buf ( n283003 , n283002 );
nand ( n283004 , n268681 , n271774 );
or ( n283005 , n270378 , n283004 );
not ( n283006 , n270377 );
not ( n283007 , n268681 );
or ( n283008 , n283006 , n283007 );
nor ( n283009 , n271774 , n53680 );
nand ( n283010 , n283008 , n283009 );
nand ( n283011 , n39766 , n39476 );
nand ( n283012 , n283005 , n283010 , n283011 );
buf ( n283013 , n283012 );
nor ( n283014 , n255066 , n266029 );
nand ( n283015 , n266016 , n283014 );
not ( n283016 , n266028 );
not ( n283017 , n266014 );
or ( n283018 , n283016 , n283017 );
nor ( n283019 , n281941 , n238635 );
nand ( n283020 , n283018 , n283019 );
nand ( n283021 , n49054 , n27903 );
nand ( n283022 , n283015 , n283020 , n283021 );
buf ( n283023 , n283022 );
buf ( n283024 , n32636 );
buf ( n283025 , n208643 );
not ( n283026 , n276367 );
not ( n283027 , n255326 );
or ( n283028 , n283026 , n283027 );
not ( n283029 , n274883 );
nor ( n283030 , n283029 , n37725 );
nand ( n283031 , n283028 , n283030 );
nor ( n283032 , n276371 , n236795 );
nand ( n283033 , n283032 , n255326 , n283029 );
nand ( n283034 , n263598 , n30681 );
nand ( n283035 , n283031 , n283033 , n283034 );
buf ( n283036 , n283035 );
not ( n283037 , n268184 );
not ( n283038 , n277593 );
nand ( n283039 , n272518 , n283038 );
or ( n283040 , n283037 , n283039 );
not ( n283041 , n272518 );
not ( n283042 , n268182 );
or ( n283043 , n283041 , n283042 );
nor ( n283044 , n283038 , n251862 );
nand ( n283045 , n283043 , n283044 );
nand ( n283046 , n35431 , n205098 );
nand ( n283047 , n283040 , n283045 , n283046 );
buf ( n283048 , n283047 );
nand ( n283049 , n265075 , n257663 );
or ( n283050 , n283049 , n257669 );
nand ( n283051 , n283049 , n248994 );
nand ( n283052 , n31577 , n34857 );
nand ( n283053 , n283050 , n283051 , n283052 );
buf ( n283054 , n283053 );
or ( n283055 , n25335 , n279680 );
nand ( n283056 , n278618 , RI1754ab58_59);
nand ( n283057 , n25325 , n51362 );
or ( n283058 , n283057 , n249124 );
not ( n283059 , n25325 );
or ( n283060 , n283059 , n266632 );
nand ( n283061 , n283058 , n283060 );
nand ( n283062 , n283061 , n270952 );
nand ( n283063 , n283055 , n283056 , n283062 );
buf ( n283064 , n283063 );
nand ( n283065 , n269919 , n269934 );
or ( n283066 , n253139 , n283065 );
not ( n283067 , n269919 );
not ( n283068 , n253138 );
or ( n283069 , n283067 , n283068 );
nor ( n283070 , n269934 , n234021 );
nand ( n283071 , n283069 , n283070 );
nand ( n283072 , n247744 , n35543 );
nand ( n283073 , n283066 , n283071 , n283072 );
buf ( n283074 , n283073 );
not ( n283075 , n29366 );
not ( n283076 , n51381 );
or ( n283077 , n283075 , n283076 );
nand ( n283078 , n242869 , n277873 );
and ( n283079 , n283078 , n242703 );
not ( n283080 , n283078 );
not ( n283081 , n242703 );
and ( n283082 , n283080 , n283081 );
nor ( n283083 , n283079 , n283082 );
or ( n283084 , n283083 , n259651 );
nand ( n283085 , n283077 , n283084 );
buf ( n283086 , n283085 );
not ( n283087 , n250110 );
not ( n283088 , n258280 );
nand ( n283089 , n283087 , n283088 );
nand ( n283090 , n276183 , n250126 );
or ( n283091 , n283089 , n283090 );
not ( n283092 , n276183 );
not ( n283093 , n283087 );
or ( n283094 , n283092 , n283093 );
nor ( n283095 , n250126 , n250909 );
nand ( n283096 , n283094 , n283095 );
nand ( n283097 , n247744 , n38741 );
nand ( n283098 , n283091 , n283096 , n283097 );
buf ( n283099 , n283098 );
not ( n283100 , n261369 );
nand ( n283101 , n250966 , n283100 );
or ( n283102 , n261356 , n283101 );
not ( n283103 , n283100 );
not ( n283104 , n261355 );
or ( n283105 , n283103 , n283104 );
nor ( n283106 , n250966 , n52445 );
nand ( n283107 , n283105 , n283106 );
nand ( n283108 , n244987 , n31044 );
nand ( n283109 , n283102 , n283107 , n283108 );
buf ( n283110 , n283109 );
not ( n283111 , n255296 );
nand ( n283112 , n283111 , n255329 );
not ( n283113 , n283032 );
or ( n283114 , n283112 , n283113 );
nand ( n283115 , n283112 , n276368 );
nand ( n283116 , n39767 , n30647 );
nand ( n283117 , n283114 , n283115 , n283116 );
buf ( n283118 , n283117 );
not ( n283119 , n40024 );
not ( n283120 , n37728 );
or ( n283121 , n283119 , n283120 );
nand ( n283122 , n274572 , n276127 );
and ( n283123 , n283122 , n276727 );
not ( n283124 , n283122 );
and ( n283125 , n283124 , n274582 );
nor ( n283126 , n283123 , n283125 );
or ( n283127 , n283126 , n49959 );
nand ( n283128 , n283121 , n283127 );
buf ( n283129 , n283128 );
not ( n283130 , n265404 );
not ( n283131 , n269296 );
nand ( n283132 , n283130 , n283131 );
or ( n283133 , n283132 , n280470 );
nand ( n283134 , n283132 , n277045 );
nand ( n283135 , n237361 , n33292 );
nand ( n283136 , n283133 , n283134 , n283135 );
buf ( n283137 , n283136 );
not ( n283138 , n263387 );
not ( n283139 , n265130 );
nor ( n283140 , n235044 , n283139 );
or ( n283141 , n283138 , n283140 );
nand ( n283142 , n263391 , n283140 );
nand ( n283143 , n246460 , n35700 );
nand ( n283144 , n283141 , n283142 , n283143 );
buf ( n283145 , n283144 );
not ( n283146 , n251743 );
nand ( n283147 , n283146 , n281099 );
nand ( n283148 , n281102 , n226010 );
or ( n283149 , n283147 , n283148 );
nor ( n283150 , n281102 , n253904 );
nand ( n283151 , n283150 , n283147 );
nand ( n283152 , n41945 , n221006 );
nand ( n283153 , n283149 , n283151 , n283152 );
buf ( n283154 , n283153 );
or ( n283155 , n25328 , n273729 );
or ( n283156 , n25335 , n270506 );
nand ( n283157 , n283155 , n283156 );
buf ( n283158 , n283157 );
nand ( n283159 , n265286 , n258322 );
not ( n283160 , n283159 );
or ( n283161 , n282613 , n283160 );
or ( n283162 , n265275 , n283159 );
nand ( n283163 , n255116 , n36055 );
nand ( n283164 , n283161 , n283162 , n283163 );
buf ( n283165 , n283164 );
not ( n283166 , RI19abd9f8_2353);
or ( n283167 , n25328 , n283166 );
or ( n283168 , n25336 , n273089 );
nand ( n283169 , n283167 , n283168 );
buf ( n283170 , n283169 );
nand ( n283171 , n263043 , n268384 , n274226 );
not ( n283172 , n263041 );
not ( n283173 , n268384 );
or ( n283174 , n283172 , n283173 );
nor ( n283175 , n274226 , n243204 );
nand ( n283176 , n283174 , n283175 );
nand ( n283177 , n35431 , n27997 );
nand ( n283178 , n283171 , n283176 , n283177 );
buf ( n283179 , n283178 );
nand ( n283180 , n243435 , n257781 );
or ( n283181 , n283180 , n265938 );
nand ( n283182 , n257768 , n257781 );
nand ( n283183 , n283182 , n265938 , n246177 );
nand ( n283184 , n256673 , n204402 );
nand ( n283185 , n283181 , n283183 , n283184 );
buf ( n283186 , n283185 );
not ( n283187 , n256726 );
not ( n283188 , n256692 );
or ( n283189 , n283187 , n283188 );
nand ( n283190 , n283189 , n267468 );
nand ( n283191 , n267431 , n267469 );
not ( n283192 , n283191 );
not ( n283193 , n256691 );
and ( n283194 , n283192 , n283193 );
and ( n283195 , n234823 , n39221 );
nor ( n283196 , n283194 , n283195 );
nand ( n283197 , n283190 , n283196 );
buf ( n283198 , n283197 );
nor ( n283199 , n275907 , n275929 );
or ( n283200 , n277305 , n283199 );
nand ( n283201 , n276334 , n283199 );
nand ( n283202 , n31576 , n42281 );
nand ( n283203 , n283200 , n283201 , n283202 );
buf ( n283204 , n283203 );
nand ( n283205 , n269769 , n258004 );
or ( n283206 , n279386 , n283205 );
not ( n283207 , n269769 );
not ( n283208 , n279385 );
or ( n283209 , n283207 , n283208 );
not ( n283210 , n282894 );
nand ( n283211 , n283209 , n283210 );
nand ( n283212 , n239240 , n34071 );
nand ( n283213 , n283206 , n283211 , n283212 );
buf ( n283214 , n283213 );
or ( n283215 , n25328 , n274942 );
or ( n283216 , n226822 , n270362 );
nand ( n283217 , n283215 , n283216 );
buf ( n283218 , n283217 );
or ( n283219 , n25328 , n278797 );
or ( n283220 , n25335 , n271604 );
nand ( n283221 , n283219 , n283220 );
buf ( n283222 , n283221 );
not ( n283223 , n264884 );
not ( n283224 , n264905 );
nand ( n283225 , n283223 , n283224 );
not ( n283226 , n275334 );
or ( n283227 , n283225 , n283226 );
nand ( n283228 , n283225 , n272858 );
nand ( n283229 , n233501 , n32841 );
nand ( n283230 , n283227 , n283228 , n283229 );
buf ( n283231 , n283230 );
or ( n283232 , n25328 , n244996 );
not ( n283233 , RI19aac040_2482);
or ( n283234 , n25335 , n283233 );
nand ( n283235 , n283232 , n283234 );
buf ( n283236 , n283235 );
not ( n283237 , n262222 );
nand ( n283238 , n283237 , n223839 );
not ( n283239 , n266256 );
nand ( n283240 , n262224 , n283239 );
or ( n283241 , n283238 , n283240 );
not ( n283242 , n283239 );
not ( n283243 , n283237 );
or ( n283244 , n283242 , n283243 );
nor ( n283245 , n262224 , n242391 );
nand ( n283246 , n283244 , n283245 );
nand ( n283247 , n55760 , n38402 );
nand ( n283248 , n283241 , n283246 , n283247 );
buf ( n283249 , n283248 );
not ( n283250 , n268927 );
nand ( n283251 , n281625 , n283250 );
or ( n283252 , n283251 , n268917 );
nand ( n283253 , n283251 , n267663 );
nand ( n283254 , n39767 , n34933 );
nand ( n283255 , n283252 , n283253 , n283254 );
buf ( n283256 , n283255 );
not ( n283257 , n260451 );
not ( n283258 , n40599 );
not ( n283259 , n251450 );
or ( n283260 , n283258 , n283259 );
not ( n283261 , n40599 );
nand ( n283262 , n283261 , n251443 );
nand ( n283263 , n283260 , n283262 );
and ( n283264 , n283263 , n256965 );
not ( n283265 , n283263 );
and ( n283266 , n283265 , n253106 );
nor ( n283267 , n283264 , n283266 );
not ( n283268 , n283267 );
not ( n283269 , n254498 );
nand ( n283270 , n283268 , n283269 );
or ( n283271 , n283257 , n283270 );
not ( n283272 , n283268 );
not ( n283273 , n260447 );
or ( n283274 , n283272 , n283273 );
nor ( n283275 , n283269 , n237384 );
nand ( n283276 , n283274 , n283275 );
nand ( n283277 , n39766 , n32231 );
nand ( n283278 , n283271 , n283276 , n283277 );
buf ( n283279 , n283278 );
nor ( n283280 , n272152 , n282355 );
nand ( n283281 , n272164 , n283280 );
not ( n283282 , n272162 );
not ( n283283 , n272151 );
or ( n283284 , n283282 , n283283 );
nand ( n283285 , n283284 , n282353 );
nand ( n283286 , n39767 , n36324 );
nand ( n283287 , n283281 , n283285 , n283286 );
buf ( n283288 , n283287 );
not ( n283289 , n260013 );
nand ( n283290 , n283289 , n260024 );
nor ( n283291 , n266279 , n234445 );
not ( n283292 , n283291 );
or ( n283293 , n283290 , n283292 );
nand ( n283294 , n283290 , n266295 );
nand ( n283295 , n252711 , n38543 );
nand ( n283296 , n283293 , n283294 , n283295 );
buf ( n283297 , n283296 );
nand ( n283298 , n267694 , n281628 , n283250 );
not ( n283299 , n267674 );
not ( n283300 , n281628 );
or ( n283301 , n283299 , n283300 );
nor ( n283302 , n283250 , n40465 );
nand ( n283303 , n283301 , n283302 );
nand ( n283304 , n35431 , n204387 );
nand ( n283305 , n283298 , n283303 , n283304 );
buf ( n283306 , n283305 );
not ( n283307 , RI1754abd0_58);
or ( n283308 , n249126 , n283307 );
not ( n283309 , n273849 );
not ( n283310 , RI1754a5b8_71);
nand ( n283311 , n283310 , RI1754a630_70);
not ( n283312 , n283311 );
and ( n283313 , n283309 , n283312 );
and ( n283314 , n244606 , n31168 );
nor ( n283315 , n283313 , n283314 );
nand ( n283316 , n283308 , n283315 );
buf ( n283317 , n283316 );
nor ( n283318 , n262289 , n33254 );
nand ( n283319 , n283318 , n262294 , n276576 );
not ( n283320 , n262297 );
not ( n283321 , n262294 );
or ( n283322 , n283320 , n283321 );
nor ( n283323 , n276576 , n250909 );
nand ( n283324 , n283322 , n283323 );
nand ( n283325 , n31577 , n32696 );
nand ( n283326 , n283319 , n283324 , n283325 );
buf ( n283327 , n283326 );
not ( n283328 , n30415 );
not ( n283329 , n258213 );
or ( n283330 , n283328 , n283329 );
nand ( n283331 , n275521 , n248810 );
not ( n283332 , n254734 );
and ( n283333 , n283331 , n283332 );
not ( n283334 , n283331 );
and ( n283335 , n283334 , n254734 );
nor ( n283336 , n283333 , n283335 );
or ( n283337 , n283336 , n259651 );
nand ( n283338 , n283330 , n283337 );
buf ( n283339 , n283338 );
buf ( n283340 , n226914 );
buf ( n283341 , n25546 );
not ( n283342 , n25390 );
not ( n283343 , n244789 );
or ( n283344 , n283342 , n283343 );
not ( n283345 , n272966 );
nand ( n283346 , n283345 , n272978 );
not ( n283347 , n279135 );
and ( n283348 , n283346 , n283347 );
not ( n283349 , n283346 );
and ( n283350 , n283349 , n279135 );
nor ( n283351 , n283348 , n283350 );
or ( n283352 , n283351 , n255135 );
nand ( n283353 , n283344 , n283352 );
buf ( n283354 , n283353 );
buf ( n283355 , n28091 );
not ( n283356 , n275675 );
nand ( n283357 , n275686 , n283356 );
not ( n283358 , n275785 );
or ( n283359 , n283357 , n283358 );
nand ( n283360 , n283357 , n278584 );
nand ( n283361 , n247423 , n34587 );
nand ( n283362 , n283359 , n283360 , n283361 );
buf ( n283363 , n283362 );
not ( n283364 , RI1754b2d8_43);
or ( n283365 , n249126 , n283364 );
nand ( n283366 , n244606 , n204773 );
nand ( n283367 , n283365 , n283366 );
buf ( n283368 , n283367 );
not ( n283369 , RI19aa6988_2519);
or ( n283370 , n226819 , n283369 );
or ( n283371 , n25336 , n242883 );
nand ( n283372 , n283370 , n283371 );
buf ( n283373 , n283372 );
or ( n283374 , n25328 , n273923 );
or ( n283375 , n25336 , n267600 );
nand ( n283376 , n283374 , n283375 );
buf ( n283377 , n283376 );
nand ( n283378 , n274392 , n239934 );
nand ( n283379 , n274405 , n279347 );
or ( n283380 , n283378 , n283379 );
not ( n283381 , n279347 );
not ( n283382 , n274392 );
or ( n283383 , n283381 , n283382 );
nor ( n283384 , n274405 , n265700 );
nand ( n283385 , n283383 , n283384 );
nand ( n283386 , n237361 , n34723 );
nand ( n283387 , n283380 , n283385 , n283386 );
buf ( n283388 , n283387 );
buf ( n283389 , n32551 );
nand ( n283390 , n279662 , n279251 , n267386 );
not ( n283391 , n279655 );
not ( n283392 , n279251 );
or ( n283393 , n283391 , n283392 );
nor ( n283394 , n267386 , n221279 );
nand ( n283395 , n283393 , n283394 );
nand ( n283396 , n250916 , n205402 );
nand ( n283397 , n283390 , n283395 , n283396 );
buf ( n283398 , n283397 );
buf ( n283399 , n29292 );
nand ( n283400 , n270782 , n278898 );
nand ( n283401 , n283400 , n280202 , n254013 );
nand ( n283402 , n280203 , n278905 , n270782 );
nand ( n283403 , n237361 , n32023 );
nand ( n283404 , n283401 , n283402 , n283403 );
buf ( n283405 , n283404 );
not ( n283406 , n280883 );
nand ( n283407 , n280449 , n267780 );
or ( n283408 , n283406 , n283407 );
not ( n283409 , n267780 );
not ( n283410 , n267757 );
not ( n283411 , n283410 );
or ( n283412 , n283409 , n283411 );
nor ( n283413 , n280449 , n234818 );
nand ( n283414 , n283412 , n283413 );
nand ( n283415 , n41944 , n29881 );
nand ( n283416 , n283408 , n283414 , n283415 );
buf ( n283417 , n283416 );
nand ( n283418 , n273267 , n273259 );
not ( n283419 , n278442 );
or ( n283420 , n283418 , n283419 );
nor ( n283421 , n278445 , n238635 );
nand ( n283422 , n283418 , n283421 );
nand ( n283423 , n31577 , n28973 );
nand ( n283424 , n283420 , n283422 , n283423 );
buf ( n283425 , n283424 );
or ( n283426 , n25328 , n277761 );
or ( n283427 , n25335 , n281235 );
nand ( n283428 , n283426 , n283427 );
buf ( n283429 , n283428 );
or ( n283430 , n25328 , n266658 );
not ( n283431 , RI19a92528_2666);
or ( n283432 , n226822 , n283431 );
nand ( n283433 , n283430 , n283432 );
buf ( n283434 , n283433 );
not ( n283435 , n39293 );
not ( n283436 , n37728 );
or ( n283437 , n283435 , n283436 );
nand ( n283438 , n271022 , n246237 );
and ( n283439 , n283438 , n277317 );
not ( n283440 , n283438 );
and ( n283441 , n283440 , n246335 );
nor ( n283442 , n283439 , n283441 );
or ( n283443 , n283442 , n49959 );
nand ( n283444 , n283437 , n283443 );
buf ( n283445 , n283444 );
not ( n283446 , n26301 );
not ( n283447 , n234823 );
or ( n283448 , n283446 , n283447 );
nand ( n283449 , n280177 , n252099 );
not ( n283450 , n283449 );
not ( n283451 , n252196 );
and ( n283452 , n283450 , n283451 );
and ( n283453 , n283449 , n252196 );
nor ( n283454 , n283452 , n283453 );
or ( n283455 , n283454 , n251498 );
nand ( n283456 , n283448 , n283455 );
buf ( n283457 , n283456 );
nand ( n283458 , n282305 , n255527 , n267731 );
not ( n283459 , n282309 );
not ( n283460 , n255527 );
or ( n283461 , n283459 , n283460 );
nand ( n283462 , n283461 , n281199 );
nand ( n283463 , n245414 , n205355 );
nand ( n283464 , n283458 , n283462 , n283463 );
buf ( n283465 , n283464 );
nand ( n283466 , n273357 , n254528 );
nand ( n283467 , n281036 , n274458 );
or ( n283468 , n283466 , n283467 );
not ( n283469 , n273357 );
not ( n283470 , n281036 );
or ( n283471 , n283469 , n283470 );
nor ( n283472 , n274458 , n235050 );
nand ( n283473 , n283471 , n283472 );
nand ( n283474 , n31577 , n30054 );
nand ( n283475 , n283468 , n283473 , n283474 );
buf ( n283476 , n283475 );
or ( n283477 , n25328 , n262589 );
not ( n283478 , RI19aa4ed0_2530);
or ( n283479 , n226822 , n283478 );
nand ( n283480 , n283477 , n283479 );
buf ( n283481 , n283480 );
nand ( n283482 , n277457 , n267490 );
or ( n283483 , n277446 , n283482 );
not ( n283484 , n277457 );
not ( n283485 , n277445 );
or ( n283486 , n283484 , n283485 );
nand ( n283487 , n283486 , n264653 );
nand ( n283488 , n50615 , n28613 );
nand ( n283489 , n283483 , n283487 , n283488 );
buf ( n283490 , n283489 );
nand ( n283491 , n274764 , n259009 );
not ( n283492 , n240592 );
not ( n283493 , n247393 );
or ( n283494 , n283492 , n283493 );
not ( n283495 , n240592 );
nand ( n283496 , n283495 , n247399 );
nand ( n283497 , n283494 , n283496 );
and ( n283498 , n283497 , n247349 );
not ( n283499 , n283497 );
and ( n283500 , n283499 , n267358 );
nor ( n283501 , n283498 , n283500 );
nand ( n283502 , n283501 , n274789 );
or ( n283503 , n283491 , n283502 );
not ( n283504 , n274789 );
not ( n283505 , n274764 );
or ( n283506 , n283504 , n283505 );
nor ( n283507 , n283501 , n237384 );
nand ( n283508 , n283506 , n283507 );
nand ( n283509 , n245414 , n39233 );
nand ( n283510 , n283503 , n283508 , n283509 );
buf ( n283511 , n283510 );
or ( n283512 , n263532 , n248461 );
nor ( n283513 , n248470 , n49051 );
nand ( n283514 , n283512 , n283513 );
nand ( n283515 , n272401 , n248470 , n263539 );
nand ( n283516 , n41945 , n204667 );
nand ( n283517 , n283514 , n283515 , n283516 );
buf ( n283518 , n283517 );
not ( n283519 , n38984 );
not ( n283520 , n252711 );
or ( n283521 , n283519 , n283520 );
nand ( n283522 , n267458 , n267468 );
not ( n283523 , n256718 );
and ( n283524 , n283522 , n283523 );
not ( n283525 , n283522 );
and ( n283526 , n283525 , n256718 );
nor ( n283527 , n283524 , n283526 );
or ( n283528 , n283527 , n258759 );
nand ( n283529 , n283521 , n283528 );
buf ( n283530 , n283529 );
not ( n283531 , n34712 );
not ( n283532 , n244606 );
or ( n283533 , n283531 , n283532 );
not ( n283534 , RI1754c598_3);
or ( n283535 , n244611 , n283534 );
nand ( n283536 , n283533 , n283535 );
buf ( n283537 , n283536 );
or ( n283538 , n226819 , n259142 );
or ( n283539 , n25335 , n281815 );
nand ( n283540 , n283538 , n283539 );
buf ( n283541 , n283540 );
not ( n283542 , n32675 );
not ( n283543 , n245701 );
or ( n283544 , n283542 , n283543 );
nand ( n283545 , n260814 , n260827 );
and ( n283546 , n283545 , n281185 );
not ( n283547 , n283545 );
and ( n283548 , n283547 , n277488 );
nor ( n283549 , n283546 , n283548 );
or ( n283550 , n283549 , n260861 );
nand ( n283551 , n283544 , n283550 );
buf ( n283552 , n283551 );
not ( n283553 , n235633 );
not ( n283554 , n238461 );
or ( n283555 , n283553 , n283554 );
not ( n283556 , n235633 );
nand ( n283557 , n283556 , n238470 );
nand ( n283558 , n283555 , n283557 );
and ( n283559 , n283558 , n238476 );
not ( n283560 , n283558 );
and ( n283561 , n283560 , n238473 );
nor ( n283562 , n283559 , n283561 );
nand ( n283563 , n283562 , n226010 );
not ( n283564 , n271342 );
nand ( n283565 , n271332 , n283564 );
or ( n283566 , n283563 , n283565 );
not ( n283567 , n283564 );
not ( n283568 , n283562 );
or ( n283569 , n283567 , n283568 );
nor ( n283570 , n271332 , n254226 );
nand ( n283571 , n283569 , n283570 );
nand ( n283572 , n35431 , n34482 );
nand ( n283573 , n283566 , n283571 , n283572 );
buf ( n283574 , n283573 );
buf ( n283575 , n42505 );
nand ( n283576 , n248080 , n258439 );
not ( n283577 , n277430 );
or ( n283578 , n283576 , n283577 );
nor ( n283579 , n277423 , n219702 );
nand ( n283580 , n283576 , n283579 );
nand ( n283581 , n31577 , n32162 );
nand ( n283582 , n283578 , n283580 , n283581 );
buf ( n283583 , n283582 );
not ( n283584 , RI19ac1f58_2314);
or ( n283585 , n25328 , n283584 );
or ( n283586 , n25335 , n269837 );
nand ( n283587 , n283585 , n283586 );
buf ( n283588 , n283587 );
or ( n283589 , n233507 , n268710 );
or ( n283590 , n25335 , n282006 );
nand ( n283591 , n283589 , n283590 );
buf ( n283592 , n283591 );
not ( n283593 , n205912 );
not ( n283594 , n245701 );
or ( n283595 , n283593 , n283594 );
not ( n283596 , n254346 );
nand ( n283597 , n283596 , n267566 );
and ( n283598 , n283597 , n277839 );
not ( n283599 , n283597 );
and ( n283600 , n283599 , n277838 );
nor ( n283601 , n283598 , n283600 );
or ( n283602 , n283601 , n244217 );
nand ( n283603 , n283595 , n283602 );
buf ( n283604 , n283603 );
not ( n283605 , n282127 );
buf ( n283606 , n238141 );
not ( n283607 , n283606 );
not ( n283608 , n247727 );
or ( n283609 , n283607 , n283608 );
or ( n283610 , n247727 , n283606 );
nand ( n283611 , n283609 , n283610 );
not ( n283612 , n283611 );
not ( n283613 , n247733 );
and ( n283614 , n283612 , n283613 );
and ( n283615 , n283611 , n247733 );
nor ( n283616 , n283614 , n283615 );
nand ( n283617 , n283605 , n283616 );
not ( n283618 , n258502 );
not ( n283619 , n250230 );
or ( n283620 , n283618 , n283619 );
nand ( n283621 , n265774 , n258501 );
nand ( n283622 , n283620 , n283621 );
not ( n283623 , n283622 );
not ( n283624 , n250942 );
and ( n283625 , n283623 , n283624 );
and ( n283626 , n283622 , n250942 );
nor ( n283627 , n283625 , n283626 );
not ( n283628 , n283627 );
nor ( n283629 , n283628 , n234440 );
not ( n283630 , n283629 );
or ( n283631 , n283617 , n283630 );
nor ( n283632 , n283627 , n38637 );
nand ( n283633 , n283632 , n283617 );
nand ( n283634 , n261585 , n30506 );
nand ( n283635 , n283631 , n283633 , n283634 );
buf ( n283636 , n283635 );
nand ( n283637 , n274404 , n247444 );
nand ( n283638 , n274416 , n279335 );
or ( n283639 , n283637 , n283638 );
not ( n283640 , n274416 );
not ( n283641 , n274404 );
or ( n283642 , n283640 , n283641 );
nor ( n283643 , n279335 , n256481 );
nand ( n283644 , n283642 , n283643 );
nand ( n283645 , n251717 , n206630 );
nand ( n283646 , n283639 , n283644 , n283645 );
buf ( n283647 , n283646 );
not ( n283648 , n262775 );
nand ( n283649 , n283648 , n205649 );
nand ( n283650 , n268163 , n262800 );
or ( n283651 , n283649 , n283650 );
not ( n283652 , n268163 );
not ( n283653 , n283648 );
or ( n283654 , n283652 , n283653 );
nor ( n283655 , n262800 , n40465 );
nand ( n283656 , n283654 , n283655 );
nand ( n283657 , n35431 , n33712 );
nand ( n283658 , n283651 , n283656 , n283657 );
buf ( n283659 , n283658 );
not ( n283660 , n25562 );
not ( n283661 , n31577 );
or ( n283662 , n283660 , n283661 );
nand ( n283663 , n270396 , n228367 );
and ( n283664 , n283663 , n280089 );
not ( n283665 , n283663 );
not ( n283666 , n280089 );
and ( n283667 , n283665 , n283666 );
nor ( n283668 , n283664 , n283667 );
or ( n283669 , n283668 , n254515 );
nand ( n283670 , n283662 , n283669 );
buf ( n283671 , n283670 );
nand ( n283672 , n274640 , n274652 );
not ( n283673 , n274864 );
nand ( n283674 , n283673 , n247275 );
or ( n283675 , n283672 , n283674 );
not ( n283676 , n283673 );
not ( n283677 , n274640 );
or ( n283678 , n283676 , n283677 );
nor ( n283679 , n274652 , n244399 );
nand ( n283680 , n283678 , n283679 );
nand ( n283681 , n244840 , n30500 );
nand ( n283682 , n283675 , n283680 , n283681 );
buf ( n283683 , n283682 );
not ( n283684 , RI19a822e0_2779);
and ( n283685 , n283684 , n249124 );
nor ( n283686 , n283685 , RI1754c610_2);
buf ( n283687 , n283686 );
not ( n283688 , n204318 );
not ( n283689 , n234453 );
or ( n283690 , n283688 , n283689 );
not ( n283691 , n257550 );
nand ( n283692 , n283691 , n276306 );
and ( n283693 , n283692 , n278763 );
not ( n283694 , n283692 );
and ( n283695 , n283694 , n278760 );
nor ( n283696 , n283693 , n283695 );
or ( n283697 , n283696 , n35816 );
nand ( n283698 , n283690 , n283697 );
buf ( n283699 , n283698 );
or ( n283700 , n233507 , n248831 );
or ( n283701 , n25335 , n256380 );
nand ( n283702 , n283700 , n283701 );
buf ( n283703 , n283702 );
buf ( n283704 , n246739 );
not ( n283705 , n283704 );
not ( n283706 , n45253 );
or ( n283707 , n283705 , n283706 );
or ( n283708 , n45253 , n283704 );
nand ( n283709 , n283707 , n283708 );
and ( n283710 , n283709 , n255245 );
not ( n283711 , n283709 );
and ( n283712 , n283711 , n255248 );
nor ( n283713 , n283710 , n283712 );
not ( n283714 , n283713 );
nand ( n283715 , n283714 , n283088 );
not ( n283716 , n268906 );
nand ( n283717 , n272474 , n283716 );
or ( n283718 , n283715 , n283717 );
not ( n283719 , n272474 );
not ( n283720 , n283714 );
or ( n283721 , n283719 , n283720 );
not ( n283722 , n268907 );
nand ( n283723 , n283721 , n283722 );
nand ( n283724 , n31576 , n34084 );
nand ( n283725 , n283718 , n283723 , n283724 );
buf ( n283726 , n283725 );
not ( n283727 , n260679 );
nand ( n283728 , n272656 , n283727 , n249960 );
not ( n283729 , n249947 );
not ( n283730 , n283727 );
or ( n283731 , n283729 , n283730 );
nor ( n283732 , n249960 , n243204 );
nand ( n283733 , n283731 , n283732 );
nand ( n283734 , n245701 , n205062 );
nand ( n283735 , n283728 , n283733 , n283734 );
buf ( n283736 , n283735 );
not ( n283737 , n28055 );
not ( n283738 , n37728 );
or ( n283739 , n283737 , n283738 );
nand ( n283740 , n258351 , n258362 );
and ( n283741 , n283740 , n268005 );
not ( n283742 , n283740 );
and ( n283743 , n283742 , n268006 );
nor ( n283744 , n283741 , n283743 );
or ( n283745 , n283744 , n259425 );
nand ( n283746 , n283739 , n283745 );
buf ( n283747 , n283746 );
not ( n283748 , n270396 );
nand ( n283749 , n283748 , n283666 );
not ( n283750 , n280079 );
or ( n283751 , n283749 , n283750 );
not ( n283752 , n50038 );
nand ( n283753 , n283752 , n283749 );
nand ( n283754 , n261585 , n36635 );
nand ( n283755 , n283751 , n283753 , n283754 );
buf ( n283756 , n283755 );
not ( n283757 , n32722 );
not ( n283758 , n31577 );
or ( n283759 , n283757 , n283758 );
nand ( n283760 , n282389 , n264387 );
and ( n283761 , n283760 , n257262 );
not ( n283762 , n283760 );
and ( n283763 , n283762 , n266122 );
nor ( n283764 , n283761 , n283763 );
or ( n283765 , n283764 , n237358 );
nand ( n283766 , n283759 , n283765 );
buf ( n283767 , n283766 );
or ( n283768 , n25328 , n259136 );
or ( n283769 , n25336 , n283166 );
nand ( n283770 , n283768 , n283769 );
buf ( n283771 , n283770 );
buf ( n283772 , RI19ad1858_2201);
and ( n283773 , n25326 , n283772 );
buf ( n283774 , n283773 );
buf ( n283775 , n26217 );
not ( n283776 , n259403 );
nand ( n283777 , n259664 , n283776 );
or ( n283778 , n259378 , n283777 );
not ( n283779 , n259664 );
not ( n283780 , n259377 );
or ( n283781 , n283779 , n283780 );
nor ( n283782 , n283776 , n49959 );
nand ( n283783 , n283781 , n283782 );
nand ( n283784 , n237361 , n28531 );
nand ( n283785 , n283778 , n283783 , n283784 );
buf ( n283786 , n283785 );
buf ( n283787 , n32883 );
buf ( n283788 , n204960 );
nor ( n283789 , n273145 , n279135 );
or ( n283790 , n272954 , n283789 );
nor ( n283791 , n272953 , n54208 );
nand ( n283792 , n283791 , n283789 );
nand ( n283793 , n246460 , n31282 );
nand ( n283794 , n283790 , n283792 , n283793 );
buf ( n283795 , n283794 );
buf ( n283796 , n37737 );
not ( n283797 , n33012 );
not ( n283798 , n263819 );
or ( n283799 , n283797 , n283798 );
nand ( n283800 , n256934 , n263277 );
and ( n283801 , n283800 , n231460 );
not ( n283802 , n283800 );
and ( n283803 , n283802 , n231459 );
nor ( n283804 , n283801 , n283803 );
or ( n283805 , n283804 , n226003 );
nand ( n283806 , n283799 , n283805 );
buf ( n283807 , n283806 );
nand ( n283808 , n267616 , n264210 , n266478 );
not ( n283809 , n267614 );
not ( n283810 , n264210 );
or ( n283811 , n283809 , n283810 );
nor ( n283812 , n266478 , n253904 );
nand ( n283813 , n283811 , n283812 );
nand ( n283814 , n31577 , n42258 );
nand ( n283815 , n283808 , n283813 , n283814 );
buf ( n283816 , n283815 );
not ( n283817 , n39447 );
not ( n283818 , n256102 );
nand ( n283819 , n283817 , n283818 );
or ( n283820 , n55148 , n283819 );
not ( n283821 , n283817 );
not ( n283822 , n232906 );
or ( n283823 , n283821 , n283822 );
nor ( n283824 , n283818 , n233971 );
nand ( n283825 , n283823 , n283824 );
nand ( n283826 , n241378 , n28528 );
nand ( n283827 , n283820 , n283825 , n283826 );
buf ( n283828 , n283827 );
not ( n283829 , n257310 );
nand ( n283830 , n256529 , n283829 );
or ( n283831 , n263969 , n283830 );
not ( n283832 , n283829 );
not ( n283833 , n263968 );
or ( n283834 , n283832 , n283833 );
nor ( n283835 , n256529 , n27889 );
nand ( n283836 , n283834 , n283835 );
nand ( n283837 , n246460 , n29850 );
nand ( n283838 , n283831 , n283836 , n283837 );
buf ( n283839 , n283838 );
nand ( n283840 , n239401 , n241704 );
nand ( n283841 , n263863 , n239781 );
or ( n283842 , n283840 , n283841 );
not ( n283843 , n239781 );
not ( n283844 , n239401 );
or ( n283845 , n283843 , n283844 );
nor ( n283846 , n263863 , n250909 );
nand ( n283847 , n283845 , n283846 );
nand ( n283848 , n247744 , n45239 );
nand ( n283849 , n283842 , n283847 , n283848 );
buf ( n283850 , n283849 );
nand ( n283851 , n281097 , n244393 );
nand ( n283852 , n281106 , n268600 );
or ( n283853 , n283851 , n283852 );
not ( n283854 , n281097 );
not ( n283855 , n281106 );
or ( n283856 , n283854 , n283855 );
nor ( n283857 , n268600 , n252872 );
nand ( n283858 , n283856 , n283857 );
nand ( n283859 , n253486 , n28900 );
nand ( n283860 , n283853 , n283858 , n283859 );
buf ( n283861 , n283860 );
not ( n283862 , n28273 );
not ( n283863 , n37728 );
or ( n283864 , n283862 , n283863 );
nand ( n283865 , n278421 , n278419 );
not ( n283866 , n273808 );
and ( n283867 , n283865 , n283866 );
not ( n283868 , n283865 );
and ( n283869 , n283868 , n273808 );
nor ( n283870 , n283867 , n283869 );
or ( n283871 , n283870 , n259425 );
nand ( n283872 , n283864 , n283871 );
buf ( n283873 , n283872 );
nand ( n283874 , n278597 , n254528 );
not ( n283875 , n274139 );
nand ( n283876 , n274151 , n283875 );
not ( n283877 , n283876 );
or ( n283878 , n283874 , n283877 );
or ( n283879 , n278599 , n283876 );
nand ( n283880 , n255116 , n36044 );
nand ( n283881 , n283878 , n283879 , n283880 );
buf ( n283882 , n283881 );
nand ( n283883 , n269560 , n205649 );
nand ( n283884 , n262844 , n281463 );
or ( n283885 , n283883 , n283884 );
not ( n283886 , n269560 );
not ( n283887 , n262844 );
or ( n283888 , n283886 , n283887 );
nor ( n283889 , n281463 , n258369 );
nand ( n283890 , n283888 , n283889 );
nand ( n283891 , n250916 , n33731 );
nand ( n283892 , n283885 , n283890 , n283891 );
buf ( n283893 , n283892 );
nand ( n283894 , n255468 , n266256 );
not ( n283895 , n283894 );
or ( n283896 , n262223 , n283895 );
or ( n283897 , n283238 , n283894 );
nand ( n283898 , n263598 , n29529 );
nand ( n283899 , n283896 , n283897 , n283898 );
buf ( n283900 , n283899 );
nor ( n283901 , n263489 , n263499 );
or ( n283902 , n283901 , n280646 );
nor ( n283903 , n280645 , n274333 );
nand ( n283904 , n283903 , n283901 );
nand ( n283905 , n234453 , n31379 );
nand ( n283906 , n283902 , n283904 , n283905 );
buf ( n283907 , n283906 );
not ( n283908 , n278472 );
nand ( n283909 , n252382 , n252449 );
or ( n283910 , n283908 , n283909 );
not ( n283911 , n278465 );
not ( n283912 , n252382 );
or ( n283913 , n283911 , n283912 );
nor ( n283914 , n252449 , n233972 );
nand ( n283915 , n283913 , n283914 );
nand ( n283916 , n48251 , n31466 );
nand ( n283917 , n283910 , n283915 , n283916 );
buf ( n283918 , n283917 );
not ( n283919 , RI1754b4b8_39);
or ( n283920 , n249128 , n283919 );
nand ( n283921 , n249131 , n207567 );
nand ( n283922 , n283920 , n283921 );
buf ( n283923 , n283922 );
or ( n283924 , n226819 , n278632 );
or ( n283925 , n25335 , n274040 );
nand ( n283926 , n283924 , n283925 );
buf ( n283927 , n283926 );
not ( n283928 , n33171 );
not ( n283929 , n234453 );
or ( n283930 , n283928 , n283929 );
not ( n283931 , n271076 );
nand ( n283932 , n283931 , n272255 );
not ( n283933 , n280050 );
and ( n283934 , n283932 , n283933 );
not ( n283935 , n283932 );
and ( n283936 , n283935 , n280050 );
nor ( n283937 , n283934 , n283936 );
or ( n283938 , n283937 , n52445 );
nand ( n283939 , n283930 , n283938 );
buf ( n283940 , n283939 );
not ( n283941 , RI19a95048_2647);
or ( n283942 , n25328 , n283941 );
or ( n283943 , n25335 , n281922 );
nand ( n283944 , n283942 , n283943 );
buf ( n283945 , n283944 );
not ( n283946 , n39409 );
not ( n283947 , n251465 );
or ( n283948 , n283946 , n283947 );
nand ( n283949 , n258963 , n273400 );
not ( n283950 , n258977 );
and ( n283951 , n283949 , n283950 );
not ( n283952 , n283949 );
and ( n283953 , n283952 , n258977 );
nor ( n283954 , n283951 , n283953 );
or ( n283955 , n283954 , n256214 );
nand ( n283956 , n283948 , n283955 );
buf ( n283957 , n283956 );
nand ( n283958 , n279543 , n258918 );
nand ( n283959 , n265433 , n265444 );
or ( n283960 , n283958 , n283959 );
not ( n283961 , n265433 );
not ( n283962 , n279543 );
or ( n283963 , n283961 , n283962 );
nor ( n283964 , n265444 , n251361 );
nand ( n283965 , n283963 , n283964 );
nand ( n283966 , n237361 , n28427 );
nand ( n283967 , n283960 , n283965 , n283966 );
buf ( n283968 , n283967 );
nor ( n283969 , n265694 , n277902 );
or ( n283970 , n259581 , n283969 );
nand ( n283971 , n277891 , n283969 );
nand ( n283972 , n255116 , n31945 );
nand ( n283973 , n283970 , n283971 , n283972 );
buf ( n283974 , n283973 );
not ( n283975 , n261206 );
not ( n283976 , n270072 );
nand ( n283977 , n261203 , n283976 );
or ( n283978 , n283975 , n283977 );
nand ( n283979 , n276653 , n283977 );
nand ( n283980 , n262000 , n28849 );
nand ( n283981 , n283978 , n283979 , n283980 );
buf ( n283982 , n283981 );
or ( n283983 , n226819 , n233516 );
not ( n283984 , RI19ac4280_2298);
or ( n283985 , n25335 , n283984 );
nand ( n283986 , n283983 , n283985 );
buf ( n283987 , n283986 );
or ( n283988 , n233507 , n251567 );
or ( n283989 , n226822 , n268132 );
nand ( n283990 , n283988 , n283989 );
buf ( n283991 , n283990 );
not ( n283992 , RI19ab5f28_2409);
or ( n283993 , n25328 , n283992 );
or ( n283994 , n226822 , n259140 );
nand ( n283995 , n283993 , n283994 );
buf ( n283996 , n283995 );
nor ( n283997 , n279094 , n255358 );
nand ( n283998 , n281402 , n283997 );
not ( n283999 , n281397 );
not ( n284000 , n255358 );
nand ( n284001 , n283999 , n284000 );
nand ( n284002 , n284001 , n279094 , n253565 );
nand ( n284003 , n241378 , n220531 );
nand ( n284004 , n283998 , n284002 , n284003 );
buf ( n284005 , n284004 );
nand ( n284006 , n283713 , n257792 );
nand ( n284007 , n268894 , n283716 );
or ( n284008 , n284006 , n284007 );
not ( n284009 , n283716 );
not ( n284010 , n283713 );
or ( n284011 , n284009 , n284010 );
nor ( n284012 , n268894 , n237384 );
nand ( n284013 , n284011 , n284012 );
nand ( n284014 , n247423 , n41252 );
nand ( n284015 , n284008 , n284013 , n284014 );
buf ( n284016 , n284015 );
nand ( n284017 , n277838 , n277840 );
or ( n284018 , n284017 , n267557 );
not ( n284019 , n267556 );
not ( n284020 , n277838 );
or ( n284021 , n284019 , n284020 );
nor ( n284022 , n277840 , n55152 );
nand ( n284023 , n284021 , n284022 );
nand ( n284024 , n31577 , n28181 );
nand ( n284025 , n284018 , n284023 , n284024 );
buf ( n284026 , n284025 );
nor ( n284027 , n276934 , n280801 );
not ( n284028 , n284027 );
nand ( n284029 , n276937 , n280801 , n277389 );
nor ( n284030 , n280801 , n235732 );
nand ( n284031 , n284030 , n277388 );
nand ( n284032 , n246217 , n26329 );
nand ( n284033 , n284028 , n284029 , n284031 , n284032 );
buf ( n284034 , n284033 );
not ( n284035 , n31365 );
not ( n284036 , n244073 );
or ( n284037 , n284035 , n284036 );
not ( n284038 , n268775 );
nand ( n284039 , n284038 , n268765 );
and ( n284040 , n284039 , n274066 );
not ( n284041 , n284039 );
and ( n284042 , n284041 , n270900 );
nor ( n284043 , n284040 , n284042 );
or ( n284044 , n284043 , n235052 );
nand ( n284045 , n284037 , n284044 );
buf ( n284046 , n284045 );
not ( n284047 , n36995 );
not ( n284048 , n237361 );
or ( n284049 , n284047 , n284048 );
not ( n284050 , n274326 );
nand ( n284051 , n280592 , n284050 );
and ( n284052 , n284051 , n262370 );
not ( n284053 , n284051 );
and ( n284054 , n284053 , n262369 );
nor ( n284055 , n284052 , n284054 );
or ( n284056 , n284055 , n255967 );
nand ( n284057 , n284049 , n284056 );
buf ( n284058 , n284057 );
not ( n284059 , n274630 );
nor ( n284060 , n284059 , n254226 );
nand ( n284061 , n284060 , n283673 );
nor ( n284062 , n274853 , n283673 );
nand ( n284063 , n274655 , n284062 );
nor ( n284064 , n274864 , n253904 );
nand ( n284065 , n284064 , n274853 );
nand ( n284066 , n256673 , n39937 );
nand ( n284067 , n284061 , n284063 , n284065 , n284066 );
buf ( n284068 , n284067 );
not ( n284069 , n283616 );
not ( n284070 , n284069 );
not ( n284071 , n283627 );
or ( n284072 , n284070 , n284071 );
nor ( n284073 , n282115 , n52445 );
nand ( n284074 , n284072 , n284073 );
nand ( n284075 , n283629 , n282115 , n284069 );
nand ( n284076 , n255116 , n46560 );
nand ( n284077 , n284074 , n284075 , n284076 );
buf ( n284078 , n284077 );
not ( n284079 , n280405 );
nand ( n284080 , n271754 , n281065 );
or ( n284081 , n284079 , n284080 );
not ( n284082 , n271754 );
not ( n284083 , n271731 );
not ( n284084 , n284083 );
or ( n284085 , n284082 , n284084 );
nor ( n284086 , n281065 , n55146 );
nand ( n284087 , n284085 , n284086 );
nand ( n284088 , n251712 , n40793 );
nand ( n284089 , n284081 , n284087 , n284088 );
buf ( n284090 , n284089 );
nor ( n284091 , n253513 , n54208 );
nand ( n284092 , n284091 , n253538 , n278036 );
not ( n284093 , n253513 );
not ( n284094 , n284093 );
not ( n284095 , n253538 );
or ( n284096 , n284094 , n284095 );
nor ( n284097 , n278036 , n55104 );
nand ( n284098 , n284096 , n284097 );
nand ( n284099 , n31577 , n33147 );
nand ( n284100 , n284092 , n284098 , n284099 );
buf ( n284101 , n284100 );
nand ( n284102 , n270036 , n250062 );
nand ( n284103 , n250050 , n253393 );
or ( n284104 , n284102 , n284103 );
nand ( n284105 , n250050 , n250062 );
nand ( n284106 , n284105 , n270035 , n259847 );
nand ( n284107 , n233501 , n25608 );
nand ( n284108 , n284104 , n284106 , n284107 );
buf ( n284109 , n284108 );
or ( n284110 , n25328 , n241982 );
or ( n284111 , n25335 , n264287 );
nand ( n284112 , n284110 , n284111 );
buf ( n284113 , n284112 );
or ( n284114 , n233507 , n283233 );
or ( n284115 , n226822 , n271087 );
nand ( n284116 , n284114 , n284115 );
buf ( n284117 , n284116 );
nand ( n284118 , n244807 , n235051 );
nand ( n284119 , n262482 , n244830 );
or ( n284120 , n284118 , n284119 );
not ( n284121 , n244830 );
not ( n284122 , n244807 );
or ( n284123 , n284121 , n284122 );
nor ( n284124 , n262482 , n47173 );
nand ( n284125 , n284123 , n284124 );
nand ( n284126 , n41944 , n32367 );
nand ( n284127 , n284120 , n284125 , n284126 );
buf ( n284128 , n284127 );
nand ( n284129 , n251239 , n256322 );
not ( n284130 , n275098 );
nand ( n284131 , n284130 , n54200 );
or ( n284132 , n284129 , n284131 );
nor ( n284133 , n284130 , n49959 );
nand ( n284134 , n284129 , n284133 );
nand ( n284135 , n247744 , n37843 );
nand ( n284136 , n284132 , n284134 , n284135 );
buf ( n284137 , n284136 );
or ( n284138 , n226819 , n280726 );
or ( n284139 , n25335 , n272352 );
nand ( n284140 , n284138 , n284139 );
buf ( n284141 , n284140 );
not ( n284142 , n271378 );
nand ( n284143 , n284142 , n270018 );
not ( n284144 , n284143 );
nor ( n284145 , n271380 , n31572 );
not ( n284146 , n284145 );
or ( n284147 , n284144 , n284146 );
nor ( n284148 , n271378 , n252070 );
and ( n284149 , n284148 , n271380 , n270018 );
and ( n284150 , n204271 , n239240 );
nor ( n284151 , n284149 , n284150 );
nand ( n284152 , n284147 , n284151 );
buf ( n284153 , n284152 );
not ( n284154 , n29394 );
not ( n284155 , n257764 );
or ( n284156 , n284154 , n284155 );
nand ( n284157 , n266292 , n266288 );
and ( n284158 , n284157 , n283289 );
not ( n284159 , n284157 );
and ( n284160 , n284159 , n260013 );
nor ( n284161 , n284158 , n284160 );
or ( n284162 , n284161 , n258179 );
nand ( n284163 , n284156 , n284162 );
buf ( n284164 , n284163 );
not ( n284165 , n29466 );
not ( n284166 , n39766 );
or ( n284167 , n284165 , n284166 );
not ( n284168 , n283501 );
nand ( n284169 , n284168 , n277528 );
and ( n284170 , n284169 , n274778 );
not ( n284171 , n284169 );
and ( n284172 , n284171 , n274777 );
nor ( n284173 , n284170 , n284172 );
or ( n284174 , n284173 , n261009 );
nand ( n284175 , n284167 , n284174 );
buf ( n284176 , n284175 );
nand ( n284177 , n264211 , n266478 );
or ( n284178 , n266468 , n284177 );
not ( n284179 , n226010 );
nor ( n284180 , n284179 , n266467 );
nand ( n284181 , n284180 , n284177 );
nand ( n284182 , n245221 , n204815 );
nand ( n284183 , n284178 , n284181 , n284182 );
buf ( n284184 , n284183 );
nand ( n284185 , n264557 , n254013 );
nand ( n284186 , n264569 , n241062 );
or ( n284187 , n284185 , n284186 );
not ( n284188 , n264569 );
not ( n284189 , n264557 );
or ( n284190 , n284188 , n284189 );
nor ( n284191 , n241062 , n52445 );
nand ( n284192 , n284190 , n284191 );
nand ( n284193 , n39766 , n31970 );
nand ( n284194 , n284187 , n284192 , n284193 );
buf ( n284195 , n284194 );
not ( n284196 , n268048 );
nand ( n284197 , n267639 , n235213 );
or ( n284198 , n284196 , n284197 );
not ( n284199 , n267639 );
not ( n284200 , n268044 );
not ( n284201 , n284200 );
or ( n284202 , n284199 , n284201 );
nand ( n284203 , n284202 , n235733 );
nand ( n284204 , n256673 , n217588 );
nand ( n284205 , n284198 , n284203 , n284204 );
buf ( n284206 , n284205 );
or ( n284207 , n25328 , n279682 );
or ( n284208 , n226822 , n279463 );
nand ( n284209 , n284207 , n284208 );
buf ( n284210 , n284209 );
or ( n284211 , n25328 , n269839 );
not ( n284212 , RI19ac0680_2328);
or ( n284213 , n25336 , n284212 );
nand ( n284214 , n284211 , n284213 );
buf ( n284215 , n284214 );
not ( n284216 , n29666 );
not ( n284217 , n245702 );
or ( n284218 , n284216 , n284217 );
nand ( n284219 , n274021 , n267144 );
and ( n284220 , n284219 , n274010 );
not ( n284221 , n284219 );
not ( n284222 , n274010 );
and ( n284223 , n284221 , n284222 );
nor ( n284224 , n284220 , n284223 );
or ( n284225 , n284224 , n259425 );
nand ( n284226 , n284218 , n284225 );
buf ( n284227 , n284226 );
or ( n284228 , n25328 , n269075 );
or ( n284229 , n226822 , n236802 );
nand ( n284230 , n284228 , n284229 );
buf ( n284231 , n284230 );
not ( n284232 , n29196 );
not ( n284233 , n245702 );
or ( n284234 , n284232 , n284233 );
nand ( n284235 , n265166 , n278090 );
not ( n284236 , n284235 );
not ( n284237 , n265176 );
and ( n284238 , n284236 , n284237 );
and ( n284239 , n284235 , n265176 );
nor ( n284240 , n284238 , n284239 );
or ( n284241 , n284240 , n49959 );
nand ( n284242 , n284234 , n284241 );
buf ( n284243 , n284242 );
nand ( n284244 , n262845 , n281463 );
or ( n284245 , n281453 , n284244 );
nand ( n284246 , n269559 , n284244 );
nand ( n284247 , n251465 , n247098 );
nand ( n284248 , n284245 , n284246 , n284247 );
buf ( n284249 , n284248 );
nand ( n284250 , n273976 , n282749 );
or ( n284251 , n271459 , n284250 );
not ( n284252 , n273976 );
not ( n284253 , n271458 );
or ( n284254 , n284252 , n284253 );
nor ( n284255 , n282749 , n55146 );
nand ( n284256 , n284254 , n284255 );
nand ( n284257 , n245414 , n26188 );
nand ( n284258 , n284251 , n284256 , n284257 );
buf ( n284259 , n284258 );
not ( n284260 , RI1754b0f8_47);
or ( n284261 , n249126 , n284260 );
nand ( n284262 , n249131 , n35519 );
nand ( n284263 , n284261 , n284262 );
buf ( n284264 , n284263 );
not ( n284265 , n35837 );
not ( n284266 , n258213 );
or ( n284267 , n284265 , n284266 );
nand ( n284268 , n263775 , n267321 );
and ( n284269 , n284268 , n263800 );
not ( n284270 , n284268 );
and ( n284271 , n284270 , n263799 );
nor ( n284272 , n284269 , n284271 );
or ( n284273 , n284272 , n226003 );
nand ( n284274 , n284267 , n284273 );
buf ( n284275 , n284274 );
nand ( n284276 , n257118 , n249613 );
or ( n284277 , n267296 , n284276 );
not ( n284278 , n249613 );
not ( n284279 , n249530 );
or ( n284280 , n284278 , n284279 );
nor ( n284281 , n257118 , n247698 );
nand ( n284282 , n284280 , n284281 );
nand ( n284283 , n35431 , n207761 );
nand ( n284284 , n284277 , n284282 , n284283 );
buf ( n284285 , n284284 );
not ( n284286 , n255273 );
nand ( n284287 , n260200 , n284286 );
nand ( n284288 , n284287 , n259466 , n251859 );
not ( n284289 , n259466 );
nand ( n284290 , n284289 , n255279 , n260200 );
nand ( n284291 , n237714 , n37496 );
nand ( n284292 , n284288 , n284290 , n284291 );
buf ( n284293 , n284292 );
nand ( n284294 , n271226 , n259981 );
not ( n284295 , n265700 );
nand ( n284296 , n284295 , n275947 );
or ( n284297 , n284294 , n284296 );
nand ( n284298 , n284294 , n275948 );
nand ( n284299 , n246217 , n205012 );
nand ( n284300 , n284297 , n284298 , n284299 );
buf ( n284301 , n284300 );
not ( n284302 , n265660 );
not ( n284303 , n275045 );
nand ( n284304 , n284303 , n265666 );
or ( n284305 , n284302 , n284304 );
nand ( n284306 , n264313 , n284304 );
nand ( n284307 , n31576 , n29802 );
nand ( n284308 , n284305 , n284306 , n284307 );
buf ( n284309 , n284308 );
or ( n284310 , n25328 , n275414 );
or ( n284311 , n25336 , n277623 );
nand ( n284312 , n284310 , n284311 );
buf ( n284313 , n284312 );
buf ( n284314 , n37331 );
buf ( n284315 , n43257 );
buf ( n284316 , n36655 );
not ( n284317 , RI1754c0e8_13);
or ( n284318 , n51369 , n284317 );
nand ( n284319 , n249131 , n34508 );
nand ( n284320 , n284318 , n284319 );
buf ( n284321 , n284320 );
nand ( n284322 , n282536 , n35420 );
or ( n284323 , n284322 , n278931 );
not ( n284324 , n278922 );
not ( n284325 , n282536 );
or ( n284326 , n284324 , n284325 );
nor ( n284327 , n35420 , n35427 );
nand ( n284328 , n284326 , n284327 );
nand ( n284329 , n252711 , n227247 );
nand ( n284330 , n284323 , n284328 , n284329 );
buf ( n284331 , n284330 );
nand ( n284332 , n283267 , n254227 );
nand ( n284333 , n254488 , n283269 );
or ( n284334 , n284332 , n284333 );
not ( n284335 , n283269 );
not ( n284336 , n283267 );
or ( n284337 , n284335 , n284336 );
nor ( n284338 , n254488 , n39763 );
nand ( n284339 , n284337 , n284338 );
nand ( n284340 , n241378 , n37331 );
nand ( n284341 , n284334 , n284339 , n284340 );
buf ( n284342 , n284341 );
nand ( n284343 , n273110 , n47167 );
or ( n284344 , n284343 , n262033 );
nand ( n284345 , n284343 , n279438 );
nand ( n284346 , n237361 , n33153 );
nand ( n284347 , n284344 , n284345 , n284346 );
buf ( n284348 , n284347 );
nand ( n284349 , n238631 , n246177 );
nand ( n284350 , n260852 , n263177 );
or ( n284351 , n284349 , n284350 );
not ( n284352 , n263177 );
not ( n284353 , n238631 );
or ( n284354 , n284352 , n284353 );
nor ( n284355 , n260852 , n226003 );
nand ( n284356 , n284354 , n284355 );
nand ( n284357 , n261585 , n205256 );
nand ( n284358 , n284351 , n284356 , n284357 );
buf ( n284359 , n284358 );
not ( n284360 , n283562 );
nand ( n284361 , n274515 , n284360 , n283564 );
not ( n284362 , n274511 );
not ( n284363 , n284360 );
or ( n284364 , n284362 , n284363 );
nor ( n284365 , n283564 , n50944 );
nand ( n284366 , n284364 , n284365 );
nand ( n284367 , n245414 , n36816 );
nand ( n284368 , n284361 , n284366 , n284367 );
buf ( n284369 , n284368 );
not ( n284370 , n205045 );
not ( n284371 , n233501 );
or ( n284372 , n284370 , n284371 );
nand ( n284373 , n271514 , n271498 );
and ( n284374 , n284373 , n269436 );
not ( n284375 , n284373 );
and ( n284376 , n284375 , n282227 );
nor ( n284377 , n284374 , n284376 );
or ( n284378 , n284377 , n258759 );
nand ( n284379 , n284372 , n284378 );
buf ( n284380 , n284379 );
nand ( n284381 , n276879 , n256957 );
nand ( n284382 , n276750 , n277737 );
or ( n284383 , n284381 , n284382 );
not ( n284384 , n277737 );
not ( n284385 , n276879 );
or ( n284386 , n284384 , n284385 );
nor ( n284387 , n276750 , n247212 );
nand ( n284388 , n284386 , n284387 );
nand ( n284389 , n234024 , n41350 );
nand ( n284390 , n284383 , n284388 , n284389 );
buf ( n284391 , n284390 );
or ( n284392 , n25328 , n271144 );
not ( n284393 , RI19a8dfc8_2697);
or ( n284394 , n25336 , n284393 );
nand ( n284395 , n284392 , n284394 );
buf ( n284396 , n284395 );
nor ( n284397 , n259356 , n55146 );
nand ( n284398 , n284397 , n259342 , n276157 );
not ( n284399 , n276157 );
not ( n284400 , n241372 );
or ( n284401 , n284399 , n284400 );
nor ( n284402 , n259342 , n274333 );
nand ( n284403 , n284401 , n284402 );
nand ( n284404 , n234024 , n25469 );
nand ( n284405 , n284398 , n284403 , n284404 );
buf ( n284406 , n284405 );
buf ( n284407 , n223314 );
buf ( n284408 , n34404 );
nor ( n284409 , n268163 , n268151 );
or ( n284410 , n262776 , n284409 );
nor ( n284411 , n262775 , n52445 );
nand ( n284412 , n284411 , n284409 );
nand ( n284413 , n39766 , n31486 );
nand ( n284414 , n284410 , n284412 , n284413 );
buf ( n284415 , n284414 );
nand ( n284416 , n258173 , n269381 );
or ( n284417 , n267210 , n284416 );
not ( n284418 , n258150 );
not ( n284419 , n258173 );
or ( n284420 , n284418 , n284419 );
nor ( n284421 , n269381 , n27889 );
nand ( n284422 , n284420 , n284421 );
nand ( n284423 , n48251 , n36321 );
nand ( n284424 , n284417 , n284422 , n284423 );
buf ( n284425 , n284424 );
or ( n284426 , n25328 , n272484 );
not ( n284427 , RI19ab6090_2408);
or ( n284428 , n25336 , n284427 );
nand ( n284429 , n284426 , n284428 );
buf ( n284430 , n284429 );
nor ( n284431 , n268005 , n258351 );
or ( n284432 , n258773 , n284431 );
nand ( n284433 , n267993 , n284431 );
nand ( n284434 , n31577 , n25343 );
nand ( n284435 , n284432 , n284433 , n284434 );
buf ( n284436 , n284435 );
or ( n284437 , n233507 , n282976 );
or ( n284438 , n25336 , n266937 );
nand ( n284439 , n284437 , n284438 );
buf ( n284440 , n284439 );
or ( n284441 , n25328 , n273989 );
or ( n284442 , n25335 , n271313 );
nand ( n284443 , n284441 , n284442 );
buf ( n284444 , n284443 );
buf ( n284445 , n33557 );
buf ( n284446 , n205414 );
buf ( n284447 , n25419 );
buf ( n284448 , n29893 );
not ( n284449 , RI19a23330_2795);
or ( n284450 , n25328 , n284449 );
or ( n284451 , n25335 , n277114 );
nand ( n284452 , n284450 , n284451 );
buf ( n284453 , n284452 );
buf ( n284454 , n29984 );
nor ( n284455 , n264998 , n253577 );
nand ( n284456 , n277962 , n284455 );
not ( n284457 , n277966 );
not ( n284458 , n264998 );
not ( n284459 , n284458 );
or ( n284460 , n284457 , n284459 );
not ( n284461 , n253577 );
nor ( n284462 , n284461 , n234440 );
nand ( n284463 , n284460 , n284462 );
nand ( n284464 , n31577 , n204880 );
nand ( n284465 , n284456 , n284463 , n284464 );
buf ( n284466 , n284465 );
buf ( n284467 , n205277 );
nor ( n284468 , n259195 , n236795 );
not ( n284469 , n49308 );
not ( n284470 , n247126 );
or ( n284471 , n284469 , n284470 );
or ( n284472 , n247126 , n49308 );
nand ( n284473 , n284471 , n284472 );
and ( n284474 , n284473 , n247250 );
not ( n284475 , n284473 );
and ( n284476 , n284475 , n247196 );
nor ( n284477 , n284474 , n284476 );
nand ( n284478 , n284468 , n284477 , n259221 );
not ( n284479 , n259195 );
not ( n284480 , n284479 );
not ( n284481 , n284477 );
or ( n284482 , n284480 , n284481 );
nor ( n284483 , n259221 , n239237 );
nand ( n284484 , n284482 , n284483 );
nand ( n284485 , n41944 , n30255 );
nand ( n284486 , n284478 , n284484 , n284485 );
buf ( n284487 , n284486 );
not ( n284488 , n26450 );
not ( n284489 , n234823 );
or ( n284490 , n284488 , n284489 );
not ( n284491 , n272561 );
nand ( n284492 , n262900 , n284491 );
and ( n284493 , n284492 , n262890 );
not ( n284494 , n284492 );
not ( n284495 , n262890 );
and ( n284496 , n284494 , n284495 );
nor ( n284497 , n284493 , n284496 );
or ( n284498 , n284497 , n235052 );
nand ( n284499 , n284490 , n284498 );
buf ( n284500 , n284499 );
not ( n284501 , n34531 );
not ( n284502 , n55760 );
or ( n284503 , n284501 , n284502 );
not ( n284504 , n273887 );
nand ( n284505 , n284504 , n270985 );
and ( n284506 , n284505 , n264524 );
not ( n284507 , n284505 );
and ( n284508 , n284507 , n264523 );
nor ( n284509 , n284506 , n284508 );
or ( n284510 , n284509 , n246091 );
nand ( n284511 , n284503 , n284510 );
buf ( n284512 , n284511 );
not ( n284513 , n267537 );
nand ( n284514 , n269800 , n270202 );
or ( n284515 , n284513 , n284514 );
not ( n284516 , n270202 );
not ( n284517 , n267511 );
or ( n284518 , n284516 , n284517 );
nor ( n284519 , n269800 , n40465 );
nand ( n284520 , n284518 , n284519 );
nand ( n284521 , n234024 , n31480 );
nand ( n284522 , n284515 , n284520 , n284521 );
buf ( n284523 , n284522 );
buf ( n284524 , n26401 );
buf ( n284525 , n30564 );
nor ( n284526 , n275567 , n237384 );
nand ( n284527 , n284526 , n273216 , n271806 );
not ( n284528 , n275567 );
nand ( n284529 , n273216 , n284528 );
nand ( n284530 , n284529 , n271807 , n246697 );
nand ( n284531 , n255116 , n30876 );
nand ( n284532 , n284527 , n284530 , n284531 );
buf ( n284533 , n284532 );
not ( n284534 , n271053 );
not ( n284535 , n283933 );
or ( n284536 , n284534 , n284535 );
nor ( n284537 , n271065 , n33254 );
nand ( n284538 , n284536 , n284537 );
nand ( n284539 , n280052 , n283933 , n271065 );
nand ( n284540 , n258743 , n36221 );
nand ( n284541 , n284538 , n284539 , n284540 );
buf ( n284542 , n284541 );
not ( n284543 , RI1754bff8_15);
or ( n284544 , n51369 , n284543 );
nand ( n284545 , n258185 , n44922 );
nand ( n284546 , n284544 , n284545 );
buf ( n284547 , n284546 );
or ( n284548 , n25328 , n270213 );
or ( n284549 , n25336 , n259766 );
nand ( n284550 , n284548 , n284549 );
buf ( n284551 , n284550 );
or ( n284552 , n233507 , n263190 );
or ( n284553 , n25335 , n251102 );
nand ( n284554 , n284552 , n284553 );
buf ( n284555 , n284554 );
or ( n284556 , n233507 , n274340 );
not ( n284557 , RI19a90818_2679);
or ( n284558 , n226822 , n284557 );
nand ( n284559 , n284556 , n284558 );
buf ( n284560 , n284559 );
not ( n284561 , n277720 );
not ( n284562 , n257352 );
or ( n284563 , n284561 , n284562 );
nand ( n284564 , n284563 , n257350 );
buf ( n284565 , n284564 );
buf ( n284566 , n27808 );
buf ( n284567 , n37446 );
buf ( n284568 , n207477 );
buf ( n284569 , n28630 );
not ( n284570 , n269165 );
nor ( n284571 , n284570 , n37725 );
nand ( n284572 , n284571 , n250400 );
nor ( n284573 , n250400 , n276625 );
nand ( n284574 , n284573 , n269168 );
nor ( n284575 , n276614 , n235895 );
nand ( n284576 , n284575 , n276625 );
nand ( n284577 , n31577 , n34638 );
nand ( n284578 , n284572 , n284574 , n284576 , n284577 );
buf ( n284579 , n284578 );
not ( n284580 , n32600 );
not ( n284581 , n237361 );
or ( n284582 , n284580 , n284581 );
not ( n284583 , n233970 );
nand ( n284584 , n284583 , n233999 );
and ( n284585 , n284584 , n272582 );
not ( n284586 , n284584 );
and ( n284587 , n284586 , n272581 );
nor ( n284588 , n284585 , n284587 );
or ( n284589 , n284588 , n244217 );
nand ( n284590 , n284582 , n284589 );
buf ( n284591 , n284590 );
not ( n284592 , n31290 );
not ( n284593 , n39766 );
or ( n284594 , n284592 , n284593 );
not ( n284595 , n278207 );
nand ( n284596 , n284595 , n268085 );
and ( n284597 , n284596 , n279866 );
not ( n284598 , n284596 );
and ( n284599 , n284598 , n268073 );
nor ( n284600 , n284597 , n284599 );
or ( n284601 , n284600 , n261009 );
nand ( n284602 , n284594 , n284601 );
buf ( n284603 , n284602 );
nand ( n284604 , n265905 , n274361 );
or ( n284605 , n278341 , n284604 );
not ( n284606 , n274358 );
not ( n284607 , n265904 );
not ( n284608 , n284607 );
or ( n284609 , n284606 , n284608 );
nor ( n284610 , n274361 , n39763 );
nand ( n284611 , n284609 , n284610 );
nand ( n284612 , n239240 , n205106 );
nand ( n284613 , n284605 , n284611 , n284612 );
buf ( n284614 , n284613 );
or ( n284615 , n25328 , n53011 );
or ( n284616 , n25335 , n261819 );
nand ( n284617 , n284615 , n284616 );
buf ( n284618 , n284617 );
or ( n284619 , n25328 , n278733 );
not ( n284620 , RI19a8cfd8_2704);
or ( n284621 , n25336 , n284620 );
nand ( n284622 , n284619 , n284621 );
buf ( n284623 , n284622 );
not ( n284624 , n270152 );
not ( n284625 , n271888 );
or ( n284626 , n284624 , n284625 );
nor ( n284627 , n271901 , n247276 );
nand ( n284628 , n284626 , n284627 );
nand ( n284629 , n271888 , n270154 , n271901 );
nand ( n284630 , n256673 , n36091 );
nand ( n284631 , n284628 , n284629 , n284630 );
buf ( n284632 , n284631 );
not ( n284633 , n261158 );
not ( n284634 , n264167 );
or ( n284635 , n284633 , n284634 );
nand ( n284636 , n284635 , n277090 );
nand ( n284637 , n261160 , n264167 , n277089 );
nand ( n284638 , n253486 , n37001 );
nand ( n284639 , n284636 , n284637 , n284638 );
buf ( n284640 , n284639 );
nor ( n284641 , n259816 , n268452 );
or ( n284642 , n259487 , n284641 );
nand ( n284643 , n268450 , n284641 );
nand ( n284644 , n255116 , n204689 );
nand ( n284645 , n284642 , n284643 , n284644 );
buf ( n284646 , n284645 );
or ( n284647 , n25328 , n280877 );
or ( n284648 , n226822 , n273841 );
nand ( n284649 , n284647 , n284648 );
buf ( n284650 , n284649 );
not ( n284651 , n29538 );
not ( n284652 , n51381 );
or ( n284653 , n284651 , n284652 );
nand ( n284654 , n258930 , n258941 );
and ( n284655 , n284654 , n255887 );
not ( n284656 , n284654 );
and ( n284657 , n284656 , n255888 );
nor ( n284658 , n284655 , n284657 );
or ( n284659 , n284658 , n256214 );
nand ( n284660 , n284653 , n284659 );
buf ( n284661 , n284660 );
nand ( n284662 , n273708 , n278124 );
or ( n284663 , n270235 , n284662 );
not ( n284664 , n278124 );
not ( n284665 , n270234 );
or ( n284666 , n284664 , n284665 );
nand ( n284667 , n284666 , n273709 );
nand ( n284668 , n251712 , n39703 );
nand ( n284669 , n284663 , n284667 , n284668 );
buf ( n284670 , n284669 );
nand ( n284671 , n278530 , n258206 );
nand ( n284672 , n260630 , n278542 );
or ( n284673 , n284671 , n284672 );
not ( n284674 , n278542 );
not ( n284675 , n278530 );
or ( n284676 , n284674 , n284675 );
nand ( n284677 , n284676 , n260631 );
nand ( n284678 , n241068 , n30012 );
nand ( n284679 , n284673 , n284677 , n284678 );
buf ( n284680 , n284679 );
not ( n284681 , n277422 );
not ( n284682 , n248002 );
or ( n284683 , n284681 , n284682 );
nand ( n284684 , n284683 , n258441 );
nand ( n284685 , n283579 , n248002 , n248069 );
nand ( n284686 , n50615 , n40410 );
nand ( n284687 , n284684 , n284685 , n284686 );
buf ( n284688 , n284687 );
not ( n284689 , n33845 );
not ( n284690 , n245702 );
or ( n284691 , n284689 , n284690 );
nand ( n284692 , n249867 , n262079 );
not ( n284693 , n284692 );
and ( n284694 , n204515 , n204516 , n245839 );
and ( n284695 , n284694 , n245003 , n204523 );
and ( n284696 , n284695 , n271935 );
not ( n284697 , n284695 );
and ( n284698 , n284697 , n249851 );
nor ( n284699 , n284696 , n284698 );
not ( n284700 , n284699 );
and ( n284701 , n284693 , n284700 );
and ( n284702 , n284692 , n284699 );
nor ( n284703 , n284701 , n284702 );
or ( n284704 , n284703 , n257174 );
nand ( n284705 , n284691 , n284704 );
buf ( n284706 , n284705 );
not ( n284707 , n34684 );
not ( n284708 , n245701 );
or ( n284709 , n284707 , n284708 );
nand ( n284710 , n277961 , n253590 );
and ( n284711 , n284710 , n264998 );
not ( n284712 , n284710 );
and ( n284713 , n284712 , n284458 );
nor ( n284714 , n284711 , n284713 );
or ( n284715 , n284714 , n244217 );
nand ( n284716 , n284709 , n284715 );
buf ( n284717 , n284716 );
or ( n284718 , n25328 , n268950 );
or ( n284719 , n226822 , n276515 );
nand ( n284720 , n284718 , n284719 );
buf ( n284721 , n284720 );
buf ( n284722 , n32231 );
not ( n284723 , n260157 );
nand ( n284724 , n284723 , n254013 );
nand ( n284725 , n260159 , n243667 );
or ( n284726 , n284724 , n284725 );
not ( n284727 , n260159 );
not ( n284728 , n284723 );
or ( n284729 , n284727 , n284728 );
nor ( n284730 , n243667 , n226003 );
nand ( n284731 , n284729 , n284730 );
nand ( n284732 , n241068 , n34260 );
nand ( n284733 , n284726 , n284731 , n284732 );
buf ( n284734 , n284733 );
nor ( n284735 , n271352 , n274511 );
or ( n284736 , n283563 , n284735 );
nand ( n284737 , n274512 , n284360 , n271353 );
nand ( n284738 , n261585 , n36038 );
nand ( n284739 , n284736 , n284737 , n284738 );
buf ( n284740 , n284739 );
buf ( n284741 , n214640 );
or ( n284742 , n25328 , n268344 );
not ( n284743 , RI19aa5dd0_2524);
or ( n284744 , n25336 , n284743 );
nand ( n284745 , n284742 , n284744 );
buf ( n284746 , n284745 );
nand ( n284747 , n277182 , n264252 );
or ( n284748 , n252726 , n284747 );
nand ( n284749 , n281353 , n284747 );
nand ( n284750 , n241068 , n33016 );
nand ( n284751 , n284748 , n284749 , n284750 );
buf ( n284752 , n284751 );
nand ( n284753 , n271695 , n247715 , n272078 );
nand ( n284754 , n272078 , n271690 );
nand ( n284755 , n284754 , n247716 , n253397 );
nand ( n284756 , n224937 , n208883 );
nand ( n284757 , n284753 , n284755 , n284756 );
buf ( n284758 , n284757 );
or ( n284759 , n233507 , n261750 );
or ( n284760 , n25335 , n265678 );
nand ( n284761 , n284759 , n284760 );
buf ( n284762 , n284761 );
nor ( n284763 , n255887 , n258930 );
or ( n284764 , n282980 , n284763 );
nand ( n284765 , n255818 , n284763 );
nand ( n284766 , n255116 , n38411 );
nand ( n284767 , n284764 , n284765 , n284766 );
buf ( n284768 , n284767 );
nand ( n284769 , n274128 , n274609 );
or ( n284770 , n283874 , n284769 );
not ( n284771 , n274609 );
not ( n284772 , n278597 );
or ( n284773 , n284771 , n284772 );
nor ( n284774 , n274128 , n31572 );
nand ( n284775 , n284773 , n284774 );
nand ( n284776 , n31577 , n220343 );
nand ( n284777 , n284770 , n284775 , n284776 );
buf ( n284778 , n284777 );
nand ( n284779 , n282871 , n279940 , n265770 );
not ( n284780 , n270861 );
not ( n284781 , n279940 );
or ( n284782 , n284780 , n284781 );
nand ( n284783 , n284782 , n265771 );
nand ( n284784 , n31577 , n204708 );
nand ( n284785 , n284779 , n284783 , n284784 );
buf ( n284786 , n284785 );
not ( n284787 , n28990 );
not ( n284788 , n233501 );
or ( n284789 , n284787 , n284788 );
nand ( n284790 , n261424 , n261436 );
and ( n284791 , n284790 , n267179 );
not ( n284792 , n284790 );
and ( n284793 , n284792 , n267178 );
nor ( n284794 , n284791 , n284793 );
or ( n284795 , n284794 , n258280 );
nand ( n284796 , n284789 , n284795 );
buf ( n284797 , n284796 );
not ( n284798 , RI1754b698_35);
or ( n284799 , n249128 , n284798 );
nand ( n284800 , n249131 , n40716 );
nand ( n284801 , n284799 , n284800 );
buf ( n284802 , n284801 );
or ( n284803 , n25328 , n283984 );
or ( n284804 , n226822 , n273084 );
nand ( n284805 , n284803 , n284804 );
buf ( n284806 , n284805 );
or ( n284807 , n233507 , n273608 );
or ( n284808 , n25336 , n283369 );
nand ( n284809 , n284807 , n284808 );
buf ( n284810 , n284809 );
not ( n284811 , n33455 );
not ( n284812 , n245943 );
or ( n284813 , n284811 , n284812 );
nand ( n284814 , n252339 , n254134 );
and ( n284815 , n284814 , n272866 );
not ( n284816 , n284814 );
and ( n284817 , n284816 , n263831 );
nor ( n284818 , n284815 , n284817 );
or ( n284819 , n284818 , n244217 );
nand ( n284820 , n284813 , n284819 );
buf ( n284821 , n284820 );
buf ( n284822 , n28702 );
or ( n284823 , n25328 , n269948 );
not ( n284824 , RI19a91808_2672);
or ( n284825 , n25335 , n284824 );
nand ( n284826 , n284823 , n284825 );
buf ( n284827 , n284826 );
not ( n284828 , n229112 );
nand ( n284829 , n284828 , n261606 );
nor ( n284830 , n270805 , n31571 );
not ( n284831 , n284830 );
or ( n284832 , n284829 , n284831 );
nand ( n284833 , n284829 , n270807 );
nand ( n284834 , n31577 , n40144 );
nand ( n284835 , n284832 , n284833 , n284834 );
buf ( n284836 , n284835 );
not ( n284837 , n237596 );
nand ( n284838 , n284837 , n270131 );
not ( n284839 , n270120 );
or ( n284840 , n284838 , n284839 );
nand ( n284841 , n284838 , n266048 );
nand ( n284842 , n31576 , n30045 );
nand ( n284843 , n284840 , n284841 , n284842 );
buf ( n284844 , n284843 );
nor ( n284845 , n262268 , n260277 );
or ( n284846 , n241460 , n284845 );
nand ( n284847 , n262258 , n284845 );
nand ( n284848 , n251465 , n33606 );
nand ( n284849 , n284846 , n284847 , n284848 );
buf ( n284850 , n284849 );
or ( n284851 , n25328 , n284743 );
or ( n284852 , n226822 , n266807 );
nand ( n284853 , n284851 , n284852 );
buf ( n284854 , n284853 );
nand ( n284855 , n279111 , n281397 , n284000 );
not ( n284856 , n279107 );
not ( n284857 , n281397 );
or ( n284858 , n284856 , n284857 );
nor ( n284859 , n284000 , n252070 );
nand ( n284860 , n284858 , n284859 );
nand ( n284861 , n245701 , n26227 );
nand ( n284862 , n284855 , n284860 , n284861 );
buf ( n284863 , n284862 );
nand ( n284864 , n257493 , n259847 );
nand ( n284865 , n242981 , n242897 );
or ( n284866 , n284864 , n284865 );
not ( n284867 , n242897 );
not ( n284868 , n257493 );
or ( n284869 , n284867 , n284868 );
nor ( n284870 , n242981 , n39763 );
nand ( n284871 , n284869 , n284870 );
nand ( n284872 , n35431 , n204467 );
nand ( n284873 , n284866 , n284871 , n284872 );
buf ( n284874 , n284873 );
nor ( n284875 , n266337 , n240080 );
nor ( n284876 , n273190 , n273192 );
nand ( n284877 , n284875 , n284876 );
not ( n284878 , n266333 );
not ( n284879 , n266310 );
or ( n284880 , n284878 , n284879 );
nor ( n284881 , n273191 , n38637 );
nand ( n284882 , n284880 , n284881 );
nand ( n284883 , n39767 , n204899 );
nand ( n284884 , n284877 , n284882 , n284883 );
buf ( n284885 , n284884 );
buf ( n284886 , RI19ad1c18_2200);
and ( n284887 , n25326 , n284886 );
buf ( n284888 , n284887 );
not ( n284889 , n280336 );
not ( n284890 , n52996 );
not ( n284891 , n245906 );
not ( n284892 , n284891 );
not ( n284893 , n52982 );
or ( n284894 , n284892 , n284893 );
not ( n284895 , n284891 );
nand ( n284896 , n284895 , n52989 );
nand ( n284897 , n284894 , n284896 );
not ( n284898 , n284897 );
or ( n284899 , n284890 , n284898 );
or ( n284900 , n284897 , n52996 );
nand ( n284901 , n284899 , n284900 );
not ( n284902 , n284901 );
not ( n284903 , n281783 );
nand ( n284904 , n284902 , n284903 );
or ( n284905 , n284889 , n284904 );
not ( n284906 , n284902 );
not ( n284907 , n280332 );
or ( n284908 , n284906 , n284907 );
nor ( n284909 , n284903 , n253544 );
nand ( n284910 , n284908 , n284909 );
nand ( n284911 , n244987 , n204456 );
nand ( n284912 , n284905 , n284910 , n284911 );
buf ( n284913 , n284912 );
not ( n284914 , n31161 );
not ( n284915 , n234823 );
or ( n284916 , n284914 , n284915 );
not ( n284917 , n249960 );
nand ( n284918 , n284917 , n249972 );
and ( n284919 , n284918 , n260689 );
not ( n284920 , n284918 );
and ( n284921 , n284920 , n260690 );
nor ( n284922 , n284919 , n284921 );
or ( n284923 , n284922 , n238223 );
nand ( n284924 , n284916 , n284923 );
buf ( n284925 , n284924 );
not ( n284926 , n34008 );
not ( n284927 , n244606 );
or ( n284928 , n284926 , n284927 );
not ( n284929 , RI1754c520_4);
or ( n284930 , n244611 , n284929 );
nand ( n284931 , n284928 , n284930 );
buf ( n284932 , n284931 );
or ( n284933 , n25328 , n282916 );
or ( n284934 , n25335 , n271189 );
nand ( n284935 , n284933 , n284934 );
buf ( n284936 , n284935 );
nor ( n284937 , n262931 , n261566 );
or ( n284938 , n269625 , n284937 );
nor ( n284939 , n261552 , n254226 );
nand ( n284940 , n284939 , n284937 );
nand ( n284941 , n249622 , n35271 );
nand ( n284942 , n284938 , n284940 , n284941 );
buf ( n284943 , n284942 );
nand ( n284944 , n263951 , n266975 , n277282 );
not ( n284945 , n263947 );
not ( n284946 , n266975 );
or ( n284947 , n284945 , n284946 );
nor ( n284948 , n277282 , n52445 );
nand ( n284949 , n284947 , n284948 );
nand ( n284950 , n244484 , n26081 );
nand ( n284951 , n284944 , n284949 , n284950 );
buf ( n284952 , n284951 );
not ( n284953 , n28262 );
not ( n284954 , n233501 );
or ( n284955 , n284953 , n284954 );
nand ( n284956 , n278923 , n34454 );
and ( n284957 , n284956 , n282537 );
not ( n284958 , n284956 );
and ( n284959 , n284958 , n282536 );
nor ( n284960 , n284957 , n284959 );
or ( n284961 , n284960 , n258280 );
nand ( n284962 , n284955 , n284961 );
buf ( n284963 , n284962 );
nor ( n284964 , n278101 , n256481 );
not ( n284965 , n265166 );
nor ( n284966 , n284965 , n278090 );
nand ( n284967 , n284964 , n284966 );
not ( n284968 , n278101 );
not ( n284969 , n284968 );
not ( n284970 , n278091 );
or ( n284971 , n284969 , n284970 );
nor ( n284972 , n265166 , n31571 );
nand ( n284973 , n284971 , n284972 );
nand ( n284974 , n239240 , n37925 );
nand ( n284975 , n284967 , n284973 , n284974 );
buf ( n284976 , n284975 );
not ( n284977 , RI1754b968_29);
or ( n284978 , n229127 , n284977 );
or ( n284979 , n25335 , n268948 );
nand ( n284980 , n284978 , n284979 );
buf ( n284981 , n284980 );
not ( n284982 , RI19a91c40_2670);
or ( n284983 , n233507 , n284982 );
or ( n284984 , n25336 , n273921 );
nand ( n284985 , n284983 , n284984 );
buf ( n284986 , n284985 );
or ( n284987 , n25328 , n254430 );
or ( n284988 , n25335 , n270946 );
nand ( n284989 , n284987 , n284988 );
buf ( n284990 , n284989 );
buf ( n284991 , n28487 );
not ( n284992 , n236540 );
not ( n284993 , n236792 );
or ( n284994 , n284992 , n284993 );
nand ( n284995 , n284994 , n280762 );
nand ( n284996 , n279885 , n236792 , n280761 );
nand ( n284997 , n237361 , n38821 );
nand ( n284998 , n284995 , n284996 , n284997 );
buf ( n284999 , n284998 );
buf ( n285000 , n31110 );
buf ( n285001 , n27699 );
nand ( n285002 , n251773 , n273523 );
or ( n285003 , n251860 , n285002 );
not ( n285004 , n251773 );
not ( n285005 , n251858 );
or ( n285006 , n285004 , n285005 );
nand ( n285007 , n285006 , n273524 );
nand ( n285008 , n35431 , n36494 );
nand ( n285009 , n285003 , n285007 , n285008 );
buf ( n285010 , n285009 );
not ( n285011 , n260024 );
nand ( n285012 , n283291 , n266296 , n285011 );
not ( n285013 , n266289 );
nand ( n285014 , n285011 , n266278 );
nand ( n285015 , n285013 , n285014 , n245241 );
nand ( n285016 , n37728 , n32344 );
nand ( n285017 , n285012 , n285015 , n285016 );
buf ( n285018 , n285017 );
nand ( n285019 , n269313 , n239934 );
nand ( n285020 , n281372 , n242208 );
or ( n285021 , n285019 , n285020 );
not ( n285022 , n281372 );
not ( n285023 , n269313 );
or ( n285024 , n285022 , n285023 );
nand ( n285025 , n285024 , n242209 );
nand ( n285026 , n234024 , n29228 );
nand ( n285027 , n285021 , n285025 , n285026 );
buf ( n285028 , n285027 );
not ( n285029 , n270438 );
not ( n285030 , n244085 );
nand ( n285031 , n285030 , n244210 );
or ( n285032 , n285029 , n285031 );
nand ( n285033 , n263740 , n285031 );
nand ( n285034 , n31577 , n29059 );
nand ( n285035 , n285032 , n285033 , n285034 );
buf ( n285036 , n285035 );
nand ( n285037 , n221727 , n226010 );
not ( n285038 , n273458 );
nand ( n285039 , n285038 , n255008 );
or ( n285040 , n285037 , n285039 );
not ( n285041 , n255008 );
not ( n285042 , n221727 );
or ( n285043 , n285041 , n285042 );
nor ( n285044 , n285038 , n55146 );
nand ( n285045 , n285043 , n285044 );
nand ( n285046 , n241068 , n28140 );
nand ( n285047 , n285040 , n285045 , n285046 );
buf ( n285048 , n285047 );
nand ( n285049 , n242594 , n275473 );
or ( n285050 , n285049 , n262530 );
nor ( n285051 , n262529 , n55152 );
nand ( n285052 , n285049 , n285051 );
nand ( n285053 , n35431 , n35001 );
nand ( n285054 , n285050 , n285052 , n285053 );
buf ( n285055 , n285054 );
buf ( n285056 , n38284 );
not ( n285057 , n282298 );
nand ( n285058 , n258112 , n240522 );
or ( n285059 , n285057 , n285058 );
not ( n285060 , n240522 );
not ( n285061 , n240157 );
not ( n285062 , n285061 );
or ( n285063 , n285060 , n285062 );
nor ( n285064 , n258112 , n251361 );
nand ( n285065 , n285063 , n285064 );
nand ( n285066 , n35431 , n35290 );
nand ( n285067 , n285059 , n285065 , n285066 );
buf ( n285068 , n285067 );
nor ( n285069 , n272550 , n284495 );
nand ( n285070 , n262903 , n285069 );
not ( n285071 , n262890 );
not ( n285072 , n262879 );
not ( n285073 , n285072 );
or ( n285074 , n285071 , n285073 );
nor ( n285075 , n277748 , n252872 );
nand ( n285076 , n285074 , n285075 );
nand ( n285077 , n55760 , n26386 );
nand ( n285078 , n285070 , n285076 , n285077 );
buf ( n285079 , n285078 );
buf ( n285080 , n36462 );
not ( n285081 , n271167 );
nand ( n285082 , n285081 , n271578 , n278359 );
nand ( n285083 , n278359 , n271573 );
nand ( n285084 , n285083 , n271167 , n223839 );
nand ( n285085 , n31577 , n204375 );
nand ( n285086 , n285082 , n285084 , n285085 );
buf ( n285087 , n285086 );
buf ( n285088 , n31069 );
not ( n285089 , RI19a84e00_2760);
or ( n285090 , n25328 , n285089 );
or ( n285091 , n25336 , n277759 );
nand ( n285092 , n285090 , n285091 );
buf ( n285093 , n285092 );
nand ( n285094 , n282522 , n247271 , n247252 );
not ( n285095 , n262119 );
not ( n285096 , n285095 );
not ( n285097 , n247271 );
or ( n285098 , n285096 , n285097 );
nor ( n285099 , n247252 , n31572 );
nand ( n285100 , n285098 , n285099 );
nand ( n285101 , n31576 , n32426 );
nand ( n285102 , n285094 , n285100 , n285101 );
buf ( n285103 , n285102 );
not ( n285104 , n31652 );
not ( n285105 , n234453 );
or ( n285106 , n285104 , n285105 );
nand ( n285107 , n271980 , n271991 );
not ( n285108 , n278821 );
and ( n285109 , n285107 , n285108 );
not ( n285110 , n285107 );
and ( n285111 , n285110 , n278821 );
nor ( n285112 , n285109 , n285111 );
or ( n285113 , n285112 , n52445 );
nand ( n285114 , n285106 , n285113 );
buf ( n285115 , n285114 );
not ( n285116 , n44182 );
not ( n285117 , n51381 );
or ( n285118 , n285116 , n285117 );
not ( n285119 , n266648 );
nand ( n285120 , n285119 , n266652 );
and ( n285121 , n285120 , n262303 );
not ( n285122 , n285120 );
and ( n285123 , n285122 , n52761 );
nor ( n285124 , n285121 , n285123 );
or ( n285125 , n285124 , n264257 );
nand ( n285126 , n285118 , n285125 );
buf ( n285127 , n285126 );
not ( n285128 , n250928 );
not ( n285129 , n279024 );
or ( n285130 , n285128 , n285129 );
not ( n285131 , n261356 );
nand ( n285132 , n285130 , n285131 );
not ( n285133 , n250930 );
nor ( n285134 , n250946 , n261355 );
nand ( n285135 , n285133 , n285134 );
nand ( n285136 , n35431 , n28348 );
nand ( n285137 , n285132 , n285135 , n285136 );
buf ( n285138 , n285137 );
or ( n285139 , n233507 , n279287 );
or ( n285140 , n25336 , n276557 );
nand ( n285141 , n285139 , n285140 );
buf ( n285142 , n285141 );
buf ( n285143 , n41245 );
buf ( n285144 , n31866 );
not ( n285145 , n39896 );
not ( n285146 , n251465 );
or ( n285147 , n285145 , n285146 );
nand ( n285148 , n273646 , n275590 );
and ( n285149 , n285148 , n282713 );
not ( n285150 , n285148 );
and ( n285151 , n285150 , n280919 );
nor ( n285152 , n285149 , n285151 );
or ( n285153 , n285152 , n55108 );
nand ( n285154 , n285147 , n285153 );
buf ( n285155 , n285154 );
buf ( n285156 , n205062 );
nand ( n285157 , n275215 , n274821 , n279215 );
not ( n285158 , n275218 );
not ( n285159 , n274821 );
or ( n285160 , n285158 , n285159 );
nor ( n285161 , n279215 , n226003 );
nand ( n285162 , n285160 , n285161 );
nand ( n285163 , n238114 , n39464 );
nand ( n285164 , n285157 , n285162 , n285163 );
buf ( n285165 , n285164 );
nand ( n285166 , n268445 , n279525 , n264725 );
not ( n285167 , n264702 );
not ( n285168 , n285167 );
not ( n285169 , n264725 );
or ( n285170 , n285168 , n285169 );
nor ( n285171 , n279525 , n252872 );
nand ( n285172 , n285170 , n285171 );
nand ( n285173 , n237714 , n29667 );
nand ( n285174 , n285166 , n285172 , n285173 );
buf ( n285175 , n285174 );
nand ( n285176 , n279380 , n269615 , n269501 );
not ( n285177 , n269603 );
not ( n285178 , n269615 );
or ( n285179 , n285177 , n285178 );
nand ( n285180 , n285179 , n269502 );
nand ( n285181 , n31577 , n205085 );
nand ( n285182 , n285176 , n285180 , n285181 );
buf ( n285183 , n285182 );
not ( n285184 , n35428 );
not ( n285185 , n256750 );
nand ( n285186 , n285184 , n285185 );
nand ( n285187 , n268054 , n261778 );
or ( n285188 , n285186 , n285187 );
not ( n285189 , n268054 );
not ( n285190 , n285185 );
or ( n285191 , n285189 , n285190 );
nand ( n285192 , n285191 , n266802 );
nand ( n285193 , n244789 , n32702 );
nand ( n285194 , n285188 , n285192 , n285193 );
buf ( n285195 , n285194 );
not ( n285196 , n40995 );
not ( n285197 , n55760 );
or ( n285198 , n285196 , n285197 );
nand ( n285199 , n262571 , n277552 );
and ( n285200 , n285199 , n256507 );
not ( n285201 , n285199 );
and ( n285202 , n285201 , n256504 );
nor ( n285203 , n285200 , n285202 );
or ( n285204 , n285203 , n46425 );
nand ( n285205 , n285198 , n285204 );
buf ( n285206 , n285205 );
or ( n285207 , n25328 , n275605 );
or ( n285208 , n25336 , n280875 );
nand ( n285209 , n285207 , n285208 );
buf ( n285210 , n285209 );
nand ( n285211 , n263386 , n259619 );
not ( n285212 , n235024 );
nand ( n285213 , n285212 , n283139 );
or ( n285214 , n285211 , n285213 );
not ( n285215 , n283139 );
not ( n285216 , n263386 );
or ( n285217 , n285215 , n285216 );
nor ( n285218 , n285212 , n38637 );
nand ( n285219 , n285217 , n285218 );
nand ( n285220 , n234024 , n39965 );
nand ( n285221 , n285214 , n285219 , n285220 );
buf ( n285222 , n285221 );
not ( n285223 , n270770 );
nand ( n285224 , n280202 , n285223 );
or ( n285225 , n278902 , n285224 );
not ( n285226 , n280202 );
not ( n285227 , n278896 );
or ( n285228 , n285226 , n285227 );
nor ( n285229 , n285223 , n254740 );
nand ( n285230 , n285228 , n285229 );
nand ( n285231 , n258213 , n31398 );
nand ( n285232 , n285225 , n285230 , n285231 );
buf ( n285233 , n285232 );
or ( n285234 , n25328 , n271537 );
or ( n285235 , n25336 , n249626 );
nand ( n285236 , n285234 , n285235 );
buf ( n285237 , n285236 );
nand ( n285238 , n276225 , n277664 );
or ( n285239 , n259282 , n285238 );
not ( n285240 , n259281 );
not ( n285241 , n276225 );
or ( n285242 , n285240 , n285241 );
nor ( n285243 , n277664 , n31572 );
nand ( n285244 , n285242 , n285243 );
nand ( n285245 , n234453 , n34534 );
nand ( n285246 , n285239 , n285244 , n285245 );
buf ( n285247 , n285246 );
nand ( n285248 , n283632 , n282115 , n282139 );
not ( n285249 , n283628 );
not ( n285250 , n282115 );
or ( n285251 , n285249 , n285250 );
nor ( n285252 , n282139 , n234021 );
nand ( n285253 , n285251 , n285252 );
nand ( n285254 , n258213 , n35681 );
nand ( n285255 , n285248 , n285253 , n285254 );
buf ( n285256 , n285255 );
not ( n285257 , n35077 );
not ( n285258 , n37728 );
or ( n285259 , n285257 , n285258 );
not ( n285260 , n260658 );
nand ( n285261 , n260649 , n285260 );
and ( n285262 , n285261 , n278542 );
not ( n285263 , n285261 );
not ( n285264 , n278542 );
and ( n285265 , n285263 , n285264 );
nor ( n285266 , n285262 , n285265 );
or ( n285267 , n285266 , n251462 );
nand ( n285268 , n285259 , n285267 );
buf ( n285269 , n285268 );
not ( n285270 , n263176 );
not ( n285271 , n260852 );
or ( n285272 , n285270 , n285271 );
nor ( n285273 , n238411 , n235895 );
nand ( n285274 , n285272 , n285273 );
nand ( n285275 , n238411 , n263183 , n260852 );
nand ( n285276 , n39767 , n50639 );
nand ( n285277 , n285274 , n285275 , n285276 );
buf ( n285278 , n285277 );
or ( n285279 , n25328 , n273871 );
or ( n285280 , n226822 , n282176 );
nand ( n285281 , n285279 , n285280 );
buf ( n285282 , n285281 );
buf ( n285283 , n204717 );
buf ( n285284 , n205912 );
not ( n285285 , n233863 );
not ( n285286 , n285285 );
not ( n285287 , n244273 );
or ( n285288 , n285286 , n285287 );
not ( n285289 , n285285 );
nand ( n285290 , n285289 , n244282 );
nand ( n285291 , n285288 , n285290 );
and ( n285292 , n285291 , n244337 );
not ( n285293 , n285291 );
and ( n285294 , n285293 , n244347 );
nor ( n285295 , n285292 , n285294 );
nor ( n285296 , n285295 , n226003 );
not ( n285297 , n265500 );
nand ( n285298 , n285296 , n285297 , n265519 );
not ( n285299 , n285295 );
not ( n285300 , n285299 );
not ( n285301 , n285297 );
or ( n285302 , n285300 , n285301 );
nor ( n285303 , n265519 , n250909 );
nand ( n285304 , n285302 , n285303 );
nand ( n285305 , n39766 , n30598 );
nand ( n285306 , n285298 , n285304 , n285305 );
buf ( n285307 , n285306 );
not ( n285308 , n271443 );
nand ( n285309 , n261947 , n239231 );
or ( n285310 , n285308 , n285309 );
not ( n285311 , n239231 );
not ( n285312 , n239110 );
or ( n285313 , n285311 , n285312 );
nor ( n285314 , n261947 , n49051 );
nand ( n285315 , n285313 , n285314 );
nand ( n285316 , n37728 , n35876 );
nand ( n285317 , n285310 , n285315 , n285316 );
buf ( n285318 , n285317 );
not ( n285319 , n37004 );
not ( n285320 , n51381 );
or ( n285321 , n285319 , n285320 );
nand ( n285322 , n253285 , n253304 );
and ( n285323 , n285322 , n267592 );
not ( n285324 , n285322 );
not ( n285325 , n267592 );
and ( n285326 , n285324 , n285325 );
nor ( n285327 , n285323 , n285326 );
or ( n285328 , n285327 , n49959 );
nand ( n285329 , n285321 , n285328 );
buf ( n285330 , n285329 );
not ( n285331 , n205198 );
not ( n285332 , n244073 );
or ( n285333 , n285331 , n285332 );
nand ( n285334 , n257899 , n257967 );
not ( n285335 , n270548 );
and ( n285336 , n285334 , n285335 );
not ( n285337 , n285334 );
and ( n285338 , n285337 , n270548 );
nor ( n285339 , n285336 , n285338 );
or ( n285340 , n285339 , n254515 );
nand ( n285341 , n285333 , n285340 );
buf ( n285342 , n285341 );
buf ( n285343 , n40398 );
buf ( n285344 , n36514 );
not ( n285345 , n34211 );
not ( n285346 , n234453 );
or ( n285347 , n285345 , n285346 );
nand ( n285348 , n253210 , n269933 );
and ( n285349 , n285348 , n253199 );
not ( n285350 , n285348 );
and ( n285351 , n285350 , n277983 );
nor ( n285352 , n285349 , n285351 );
or ( n285353 , n285352 , n234110 );
nand ( n285354 , n285347 , n285353 );
buf ( n285355 , n285354 );
not ( n285356 , n30062 );
not ( n285357 , n239240 );
or ( n285358 , n285356 , n285357 );
nand ( n285359 , n263119 , n263130 );
and ( n285360 , n285359 , n275819 );
not ( n285361 , n285359 );
and ( n285362 , n285361 , n275818 );
nor ( n285363 , n285360 , n285362 );
or ( n285364 , n285363 , n234110 );
nand ( n285365 , n285358 , n285364 );
buf ( n285366 , n285365 );
not ( n285367 , RI19ab3c00_2425);
or ( n285368 , n25328 , n285367 );
or ( n285369 , n25335 , n279219 );
nand ( n285370 , n285368 , n285369 );
buf ( n285371 , n285370 );
or ( n285372 , n25328 , n252366 );
or ( n285373 , n25336 , n244994 );
nand ( n285374 , n285372 , n285373 );
buf ( n285375 , n285374 );
not ( n285376 , n269898 );
nor ( n285377 , n261717 , n265105 );
or ( n285378 , n285376 , n285377 );
nand ( n285379 , n265095 , n285377 );
nand ( n285380 , n37728 , n25472 );
nand ( n285381 , n285378 , n285379 , n285380 );
buf ( n285382 , n285381 );
nand ( n285383 , n272203 , n281765 , n271243 );
not ( n285384 , n272197 );
not ( n285385 , n281765 );
or ( n285386 , n285384 , n285385 );
nor ( n285387 , n271243 , n234440 );
nand ( n285388 , n285386 , n285387 );
nand ( n285389 , n255116 , n29613 );
nand ( n285390 , n285383 , n285388 , n285389 );
buf ( n285391 , n285390 );
buf ( n285392 , n32722 );
buf ( n285393 , n33517 );
not ( n285394 , n30275 );
not ( n285395 , n252711 );
or ( n285396 , n285394 , n285395 );
not ( n285397 , n261808 );
nand ( n285398 , n285397 , n261798 );
and ( n285399 , n285398 , n31563 );
not ( n285400 , n285398 );
and ( n285401 , n285400 , n31564 );
nor ( n285402 , n285399 , n285401 );
or ( n285403 , n285402 , n258759 );
nand ( n285404 , n285396 , n285403 );
buf ( n285405 , n285404 );
not ( n285406 , n276082 );
nand ( n285407 , n276095 , n285406 , n281699 );
not ( n285408 , n276098 );
not ( n285409 , n285406 );
or ( n285410 , n285408 , n285409 );
nor ( n285411 , n281699 , n27889 );
nand ( n285412 , n285410 , n285411 );
nand ( n285413 , n256292 , n36272 );
nand ( n285414 , n285407 , n285412 , n285413 );
buf ( n285415 , n285414 );
nor ( n285416 , n280319 , n284901 );
nand ( n285417 , n280333 , n285416 );
nor ( n285418 , n284902 , n47173 );
nand ( n285419 , n280331 , n281786 );
nand ( n285420 , n285418 , n285419 );
nand ( n285421 , n241976 , n28015 );
nand ( n285422 , n285417 , n285420 , n285421 );
buf ( n285423 , n285422 );
not ( n285424 , n33023 );
not ( n285425 , n255116 );
or ( n285426 , n285424 , n285425 );
not ( n285427 , n268306 );
not ( n285428 , n285427 );
nand ( n285429 , n282284 , n280139 );
not ( n285430 , n285429 );
and ( n285431 , n285428 , n285430 );
and ( n285432 , n285427 , n285429 );
nor ( n285433 , n285431 , n285432 );
or ( n285434 , n285433 , n238223 );
nand ( n285435 , n285426 , n285434 );
buf ( n285436 , n285435 );
not ( n285437 , n265508 );
nand ( n285438 , n285437 , n279011 );
nor ( n285439 , n285299 , n31571 );
not ( n285440 , n285439 );
or ( n285441 , n285438 , n285440 );
nand ( n285442 , n285438 , n285296 );
nand ( n285443 , n245414 , n33218 );
nand ( n285444 , n285441 , n285442 , n285443 );
buf ( n285445 , n285444 );
nand ( n285446 , n270072 , n270083 );
or ( n285447 , n261182 , n285446 );
not ( n285448 , n270083 );
not ( n285449 , n261181 );
or ( n285450 , n285448 , n285449 );
nor ( n285451 , n270072 , n52445 );
nand ( n285452 , n285450 , n285451 );
nand ( n285453 , n244987 , n34708 );
nand ( n285454 , n285447 , n285452 , n285453 );
buf ( n285455 , n285454 );
not ( n285456 , n280177 );
nand ( n285457 , n285456 , n252099 );
or ( n285458 , n280029 , n285457 );
not ( n285459 , n285456 );
not ( n285460 , n280028 );
or ( n285461 , n285459 , n285460 );
nor ( n285462 , n252099 , n235050 );
nand ( n285463 , n285461 , n285462 );
nand ( n285464 , n234448 , n216952 );
nand ( n285465 , n285458 , n285463 , n285464 );
buf ( n285466 , n285465 );
not ( n285467 , n229370 );
nand ( n285468 , n54331 , n285467 );
or ( n285469 , n267344 , n285468 );
not ( n285470 , n267343 );
not ( n285471 , n232090 );
not ( n285472 , n285471 );
or ( n285473 , n285470 , n285472 );
nor ( n285474 , n285467 , n250431 );
nand ( n285475 , n285473 , n285474 );
nand ( n285476 , n31577 , n29573 );
nand ( n285477 , n285469 , n285475 , n285476 );
buf ( n285478 , n285477 );
nor ( n285479 , n260129 , n42443 );
nand ( n285480 , n285479 , n280246 , n260140 );
not ( n285481 , n260129 );
nand ( n285482 , n285481 , n260140 );
nand ( n285483 , n246663 , n285482 , n244393 );
nand ( n285484 , n246217 , n29420 );
nand ( n285485 , n285480 , n285483 , n285484 );
buf ( n285486 , n285485 );
nand ( n285487 , n281372 , n242383 );
or ( n285488 , n269315 , n285487 );
and ( n285489 , n269314 , n242383 );
and ( n285490 , n285489 , n281373 , n255152 );
and ( n285491 , n244484 , n31225 );
and ( n285492 , n285488 , n285490 , n285491 );
buf ( n285493 , n285492 );
nand ( n285494 , n273820 , n278420 );
or ( n285495 , n285494 , n273833 );
not ( n285496 , n273832 );
not ( n285497 , n273820 );
or ( n285498 , n285496 , n285497 );
nor ( n285499 , n278420 , n37725 );
nand ( n285500 , n285498 , n285499 );
nand ( n285501 , n245701 , n36284 );
nand ( n285502 , n285495 , n285500 , n285501 );
buf ( n285503 , n285502 );
not ( n285504 , n270964 );
nand ( n285505 , n261673 , n266868 );
or ( n285506 , n285504 , n285505 );
not ( n285507 , n261662 );
not ( n285508 , n285507 );
not ( n285509 , n261673 );
or ( n285510 , n285508 , n285509 );
nor ( n285511 , n266868 , n40465 );
nand ( n285512 , n285510 , n285511 );
nand ( n285513 , n241976 , n42750 );
nand ( n285514 , n285506 , n285512 , n285513 );
buf ( n285515 , n285514 );
not ( n285516 , n265938 );
nand ( n285517 , n257786 , n265928 , n285516 );
not ( n285518 , n257781 );
nand ( n285519 , n285518 , n285516 );
nand ( n285520 , n285519 , n243284 , n257792 );
nand ( n285521 , n50615 , n34976 );
nand ( n285522 , n285517 , n285520 , n285521 );
buf ( n285523 , n285522 );
not ( n285524 , n221279 );
not ( n285525 , n265740 );
nand ( n285526 , n285524 , n285525 );
nand ( n285527 , n265752 , n271857 );
or ( n285528 , n285526 , n285527 );
not ( n285529 , n265752 );
not ( n285530 , n285525 );
or ( n285531 , n285529 , n285530 );
nor ( n285532 , n271857 , n247698 );
nand ( n285533 , n285531 , n285532 );
nand ( n285534 , n254798 , n207466 );
nand ( n285535 , n285528 , n285533 , n285534 );
buf ( n285536 , n285535 );
nand ( n285537 , n267805 , n269053 );
or ( n285538 , n285537 , n255153 );
nand ( n285539 , n285537 , n255169 );
nand ( n285540 , n263598 , n36064 );
nand ( n285541 , n285538 , n285539 , n285540 );
buf ( n285542 , n285541 );
nand ( n285543 , n285439 , n279012 , n285297 );
not ( n285544 , n285295 );
not ( n285545 , n279012 );
or ( n285546 , n285544 , n285545 );
nor ( n285547 , n285297 , n31572 );
nand ( n285548 , n285546 , n285547 );
nand ( n285549 , n241976 , n25707 );
nand ( n285550 , n285543 , n285548 , n285549 );
buf ( n285551 , n285550 );
or ( n285552 , n25328 , n256564 );
or ( n285553 , n25335 , n268337 );
nand ( n285554 , n285552 , n285553 );
buf ( n285555 , n285554 );
nand ( n285556 , n279171 , n235051 );
nand ( n285557 , n266101 , n266088 );
or ( n285558 , n285556 , n285557 );
not ( n285559 , n266088 );
not ( n285560 , n279171 );
or ( n285561 , n285559 , n285560 );
nor ( n285562 , n266101 , n37725 );
nand ( n285563 , n285561 , n285562 );
nand ( n285564 , n39767 , n35471 );
nand ( n285565 , n285558 , n285563 , n285564 );
buf ( n285566 , n285565 );
buf ( n285567 , n32648 );
buf ( n285568 , n25586 );
buf ( n285569 , n26431 );
buf ( n285570 , n35512 );
buf ( n285571 , n30350 );
buf ( n285572 , n33508 );
nand ( n285573 , n270035 , n250032 );
or ( n285574 , n270048 , n285573 );
not ( n285575 , n270035 );
not ( n285576 , n270047 );
or ( n285577 , n285575 , n285576 );
nor ( n285578 , n250032 , n254150 );
nand ( n285579 , n285577 , n285578 );
nand ( n285580 , n254798 , n31105 );
nand ( n285581 , n285574 , n285579 , n285580 );
buf ( n285582 , n285581 );
buf ( n285583 , n33162 );
buf ( n285584 , n30876 );
not ( n285585 , n280801 );
not ( n285586 , n285585 );
not ( n285587 , n280805 );
or ( n285588 , n285586 , n285587 );
nor ( n285589 , n276911 , n42443 );
nand ( n285590 , n285588 , n285589 );
nand ( n285591 , n284030 , n280805 , n276911 );
nand ( n285592 , n247585 , n32985 );
nand ( n285593 , n285590 , n285591 , n285592 );
buf ( n285594 , n285593 );
or ( n285595 , n226819 , n282008 );
or ( n285596 , n25335 , n282023 );
nand ( n285597 , n285595 , n285596 );
buf ( n285598 , n285597 );
or ( n285599 , n226819 , n247225 );
not ( n285600 , RI19a92960_2664);
or ( n285601 , n226822 , n285600 );
nand ( n285602 , n285599 , n285601 );
buf ( n285603 , n285602 );
nand ( n285604 , n246676 , n246481 , n260129 );
not ( n285605 , n246679 );
not ( n285606 , n246481 );
or ( n285607 , n285605 , n285606 );
nand ( n285608 , n285607 , n285479 );
nand ( n285609 , n256292 , n40780 );
nand ( n285610 , n285604 , n285608 , n285609 );
buf ( n285611 , n285610 );
not ( n285612 , n28651 );
not ( n285613 , n31577 );
or ( n285614 , n285612 , n285613 );
nand ( n285615 , n282127 , n282138 );
and ( n285616 , n285615 , n284069 );
not ( n285617 , n285615 );
and ( n285618 , n285617 , n283616 );
nor ( n285619 , n285616 , n285618 );
or ( n285620 , n285619 , n251498 );
nand ( n285621 , n285614 , n285620 );
buf ( n285622 , n285621 );
not ( n285623 , RI19aae980_2464);
or ( n285624 , n25328 , n285623 );
or ( n285625 , n226822 , n267215 );
nand ( n285626 , n285624 , n285625 );
buf ( n285627 , n285626 );
nor ( n285628 , n272474 , n268884 );
or ( n285629 , n284006 , n285628 );
nor ( n285630 , n283713 , n221279 );
nand ( n285631 , n285630 , n285628 );
nand ( n285632 , n233501 , n38171 );
nand ( n285633 , n285629 , n285631 , n285632 );
buf ( n285634 , n285633 );
not ( n285635 , n280832 );
not ( n285636 , n285635 );
nand ( n285637 , n272629 , n258814 );
not ( n285638 , n285637 );
and ( n285639 , n285636 , n285638 );
and ( n285640 , n263819 , n42764 );
nor ( n285641 , n285639 , n285640 );
not ( n285642 , n272627 );
nand ( n285643 , n285642 , n264850 );
nand ( n285644 , n264864 , n258803 );
nand ( n285645 , n285641 , n285643 , n285644 );
buf ( n285646 , n285645 );
not ( n285647 , n275887 );
not ( n285648 , n274745 );
nand ( n285649 , n275497 , n285648 );
or ( n285650 , n285647 , n285649 );
not ( n285651 , n275497 );
not ( n285652 , n275889 );
or ( n285653 , n285651 , n285652 );
nor ( n285654 , n285648 , n234110 );
nand ( n285655 , n285653 , n285654 );
nand ( n285656 , n247744 , n41145 );
nand ( n285657 , n285650 , n285655 , n285656 );
buf ( n285658 , n285657 );
not ( n285659 , n273221 );
nand ( n285660 , n275567 , n271819 );
not ( n285661 , n285660 );
and ( n285662 , n285659 , n285661 );
and ( n285663 , n233501 , n38265 );
nor ( n285664 , n285662 , n285663 );
not ( n285665 , n271797 );
nand ( n285666 , n285665 , n284528 );
nand ( n285667 , n284526 , n271818 );
nand ( n285668 , n285664 , n285666 , n285667 );
buf ( n285669 , n285668 );
or ( n285670 , n25328 , n284212 );
or ( n285671 , n25336 , n279315 );
nand ( n285672 , n285670 , n285671 );
buf ( n285673 , n285672 );
not ( n285674 , n264827 );
not ( n285675 , n257596 );
or ( n285676 , n285674 , n285675 );
nand ( n285677 , n285676 , n267699 );
nand ( n285678 , n280261 , n257596 , n264835 );
nand ( n285679 , n35431 , n31179 );
nand ( n285680 , n285677 , n285678 , n285679 );
buf ( n285681 , n285680 );
nand ( n285682 , n252852 , n252839 );
not ( n285683 , n279769 );
or ( n285684 , n285682 , n285683 );
nand ( n285685 , n285682 , n274671 );
nand ( n285686 , n31577 , n35978 );
nand ( n285687 , n285684 , n285685 , n285686 );
buf ( n285688 , n285687 );
not ( n285689 , n263715 );
nand ( n285690 , n285689 , n205649 );
nand ( n285691 , n259901 , n263717 );
or ( n285692 , n285690 , n285691 );
not ( n285693 , n263717 );
not ( n285694 , n285689 );
or ( n285695 , n285693 , n285694 );
nand ( n285696 , n285695 , n259916 );
nand ( n285697 , n247744 , n38650 );
nand ( n285698 , n285692 , n285696 , n285697 );
buf ( n285699 , n285698 );
buf ( n285700 , n33597 );
buf ( n285701 , n30801 );
buf ( n285702 , n26391 );
buf ( n285703 , n28176 );
or ( n285704 , n25328 , n244490 );
or ( n285705 , n25335 , n265252 );
nand ( n285706 , n285704 , n285705 );
buf ( n285707 , n285706 );
not ( n285708 , n262634 );
nand ( n285709 , n285708 , n270017 );
not ( n285710 , n284148 );
or ( n285711 , n285709 , n285710 );
nand ( n285712 , n285709 , n271386 );
nand ( n285713 , n46083 , n41117 );
nand ( n285714 , n285711 , n285712 , n285713 );
buf ( n285715 , n285714 );
nand ( n285716 , n247880 , n272645 );
not ( n285717 , n271599 );
or ( n285718 , n285716 , n285717 );
nand ( n285719 , n285716 , n261887 );
nand ( n285720 , n35431 , n27979 );
nand ( n285721 , n285718 , n285719 , n285720 );
buf ( n285722 , n285721 );
not ( n285723 , n270986 );
not ( n285724 , n264534 );
not ( n285725 , n285724 );
or ( n285726 , n285723 , n285725 );
nor ( n285727 , n284504 , n247276 );
nand ( n285728 , n285726 , n285727 );
nor ( n285729 , n273887 , n270985 );
nand ( n285730 , n264537 , n285729 );
nand ( n285731 , n39766 , n42604 );
nand ( n285732 , n285728 , n285730 , n285731 );
buf ( n285733 , n285732 );
nand ( n285734 , n277528 , n283501 );
or ( n285735 , n285734 , n274795 );
not ( n285736 , n274788 );
not ( n285737 , n283501 );
or ( n285738 , n285736 , n285737 );
nor ( n285739 , n277528 , n37725 );
nand ( n285740 , n285738 , n285739 );
nand ( n285741 , n37728 , n28398 );
nand ( n285742 , n285735 , n285740 , n285741 );
buf ( n285743 , n285742 );
nor ( n285744 , n265287 , n258322 );
nand ( n285745 , n285744 , n282619 );
not ( n285746 , n258321 );
not ( n285747 , n258298 );
not ( n285748 , n285747 );
or ( n285749 , n285746 , n285748 );
nor ( n285750 , n265286 , n236795 );
nand ( n285751 , n285749 , n285750 );
nand ( n285752 , n49054 , n43628 );
nand ( n285753 , n285745 , n285751 , n285752 );
buf ( n285754 , n285753 );
buf ( n285755 , n41506 );
buf ( n285756 , n34260 );
not ( n285757 , n37178 );
not ( n285758 , n252711 );
or ( n285759 , n285757 , n285758 );
not ( n285760 , n269582 );
nand ( n285761 , n285760 , n253328 );
not ( n285762 , n253340 );
and ( n285763 , n285761 , n285762 );
not ( n285764 , n285761 );
and ( n285765 , n285764 , n253340 );
nor ( n285766 , n285763 , n285765 );
or ( n285767 , n285766 , n35816 );
nand ( n285768 , n285759 , n285767 );
buf ( n285769 , n285768 );
buf ( n285770 , n41848 );
or ( n285771 , n25328 , n279620 );
or ( n285772 , n25335 , n258133 );
nand ( n285773 , n285771 , n285772 );
buf ( n285774 , n285773 );
nor ( n285775 , n261606 , n50943 );
nand ( n285776 , n284830 , n285775 );
nor ( n285777 , n270809 , n221279 );
nand ( n285778 , n261603 , n270806 );
nand ( n285779 , n285777 , n285778 );
nand ( n285780 , n31576 , n38532 );
nand ( n285781 , n285776 , n285779 , n285780 );
buf ( n285782 , n285781 );
not ( n285783 , n206043 );
not ( n285784 , n252711 );
or ( n285785 , n285783 , n285784 );
not ( n285786 , n281699 );
nand ( n285787 , n285786 , n281685 );
and ( n285788 , n285787 , n276073 );
not ( n285789 , n285787 );
and ( n285790 , n285789 , n276072 );
nor ( n285791 , n285788 , n285790 );
or ( n285792 , n285791 , n258759 );
nand ( n285793 , n285785 , n285792 );
buf ( n285794 , n285793 );
or ( n285795 , n25328 , n259716 );
or ( n285796 , n25336 , n261013 );
nand ( n285797 , n285795 , n285796 );
buf ( n285798 , n285797 );
or ( n285799 , n25328 , n277579 );
or ( n285800 , n226822 , n275165 );
nand ( n285801 , n285799 , n285800 );
buf ( n285802 , n285801 );
not ( n285803 , n256345 );
nand ( n285804 , n285803 , n256370 );
not ( n285805 , n262298 );
or ( n285806 , n285804 , n285805 );
nand ( n285807 , n285804 , n283318 );
nand ( n285808 , n245414 , n31616 );
nand ( n285809 , n285806 , n285807 , n285808 );
buf ( n285810 , n285809 );
not ( n285811 , n31500 );
not ( n285812 , n237361 );
or ( n285813 , n285811 , n285812 );
not ( n285814 , n237352 );
nand ( n285815 , n285814 , n256073 );
and ( n285816 , n285815 , n277775 );
not ( n285817 , n285815 );
not ( n285818 , n277775 );
and ( n285819 , n285817 , n285818 );
nor ( n285820 , n285816 , n285819 );
or ( n285821 , n285820 , n257174 );
nand ( n285822 , n285813 , n285821 );
buf ( n285823 , n285822 );
nand ( n285824 , n275515 , n256584 );
nand ( n285825 , n248799 , n254734 );
or ( n285826 , n285824 , n285825 );
not ( n285827 , n254734 );
not ( n285828 , n275515 );
or ( n285829 , n285827 , n285828 );
nor ( n285830 , n248799 , n252872 );
nand ( n285831 , n285829 , n285830 );
nand ( n285832 , n31576 , n28958 );
nand ( n285833 , n285826 , n285831 , n285832 );
buf ( n285834 , n285833 );
not ( n285835 , n256482 );
nand ( n285836 , n277546 , n256504 );
or ( n285837 , n285835 , n285836 );
nand ( n285838 , n262561 , n285836 );
nand ( n285839 , n245414 , n41498 );
nand ( n285840 , n285837 , n285838 , n285839 );
buf ( n285841 , n285840 );
not ( n285842 , RI19a8eb08_2692);
or ( n285843 , n25328 , n285842 );
or ( n285844 , n25336 , n273794 );
nand ( n285845 , n285843 , n285844 );
buf ( n285846 , n285845 );
or ( n285847 , n226819 , n281195 );
or ( n285848 , n226822 , n280429 );
nand ( n285849 , n285847 , n285848 );
buf ( n285850 , n285849 );
not ( n285851 , n265444 );
not ( n285852 , n285851 );
not ( n285853 , n265456 );
or ( n285854 , n285852 , n285853 );
nor ( n285855 , n279555 , n253213 );
nand ( n285856 , n285854 , n285855 );
nand ( n285857 , n265456 , n279555 , n283964 );
nand ( n285858 , n234024 , n31326 );
nand ( n285859 , n285856 , n285857 , n285858 );
buf ( n285860 , n285859 );
not ( n285861 , n25382 );
not ( n285862 , n245702 );
or ( n285863 , n285861 , n285862 );
nand ( n285864 , n259058 , n266200 );
not ( n285865 , n259069 );
and ( n285866 , n285864 , n285865 );
not ( n285867 , n285864 );
and ( n285868 , n285867 , n259069 );
nor ( n285869 , n285866 , n285868 );
or ( n285870 , n285869 , n46425 );
nand ( n285871 , n285863 , n285870 );
buf ( n285872 , n285871 );
not ( n285873 , n266230 );
not ( n285874 , n259020 );
or ( n285875 , n285873 , n285874 );
nor ( n285876 , n259031 , n46425 );
nand ( n285877 , n285875 , n285876 );
not ( n285878 , n281015 );
nand ( n285879 , n285878 , n259020 , n259031 );
nand ( n285880 , n35431 , n35330 );
nand ( n285881 , n285877 , n285879 , n285880 );
buf ( n285882 , n285881 );
or ( n285883 , n25328 , n263546 );
not ( n285884 , RI19a8c948_2707);
or ( n285885 , n226822 , n285884 );
nand ( n285886 , n285883 , n285885 );
buf ( n285887 , n285886 );
not ( n285888 , n278774 );
nand ( n285889 , n285888 , n234813 );
not ( n285890 , n285889 );
not ( n285891 , n245241 );
nor ( n285892 , n285891 , n278785 );
not ( n285893 , n285892 );
or ( n285894 , n285890 , n285893 );
nor ( n285895 , n257855 , n257868 );
and ( n285896 , n285895 , n278785 );
and ( n285897 , n30482 , n237361 );
nor ( n285898 , n285896 , n285897 );
nand ( n285899 , n285894 , n285898 );
buf ( n285900 , n285899 );
or ( n285901 , n25328 , n282944 );
or ( n285902 , n25335 , n282888 );
nand ( n285903 , n285901 , n285902 );
buf ( n285904 , n285903 );
buf ( n285905 , n205026 );
not ( n285906 , n280397 );
nand ( n285907 , n285906 , n223839 );
nand ( n285908 , n280399 , n281066 );
or ( n285909 , n285907 , n285908 );
not ( n285910 , n281066 );
not ( n285911 , n280397 );
not ( n285912 , n285911 );
or ( n285913 , n285910 , n285912 );
nor ( n285914 , n280399 , n222533 );
nand ( n285915 , n285913 , n285914 );
nand ( n285916 , n246217 , n29450 );
nand ( n285917 , n285909 , n285915 , n285916 );
buf ( n285918 , n285917 );
buf ( n285919 , n205795 );
nor ( n285920 , n259113 , n261112 );
or ( n285921 , n266882 , n285920 );
nor ( n285922 , n259100 , n226955 );
nand ( n285923 , n285922 , n285920 );
nand ( n285924 , n41945 , n40786 );
nand ( n285925 , n285921 , n285923 , n285924 );
buf ( n285926 , n285925 );
not ( n285927 , n258853 );
nand ( n285928 , n273677 , n285927 );
or ( n285929 , n273667 , n285928 );
not ( n285930 , n273677 );
not ( n285931 , n273666 );
or ( n285932 , n285930 , n285931 );
nor ( n285933 , n285927 , n239237 );
nand ( n285934 , n285932 , n285933 );
nand ( n285935 , n50615 , n34237 );
nand ( n285936 , n285929 , n285934 , n285935 );
buf ( n285937 , n285936 );
not ( n285938 , n28061 );
not ( n285939 , n255116 );
or ( n285940 , n285938 , n285939 );
not ( n285941 , n259230 );
nand ( n285942 , n280580 , n285941 );
and ( n285943 , n285942 , n284477 );
not ( n285944 , n285942 );
not ( n285945 , n284477 );
and ( n285946 , n285944 , n285945 );
nor ( n285947 , n285943 , n285946 );
or ( n285948 , n285947 , n31572 );
nand ( n285949 , n285940 , n285948 );
buf ( n285950 , n285949 );
not ( n285951 , n264420 );
nand ( n285952 , n285951 , n253941 );
or ( n285953 , n264409 , n285952 );
not ( n285954 , n285951 );
not ( n285955 , n264408 );
or ( n285956 , n285954 , n285955 );
nor ( n285957 , n253941 , n39763 );
nand ( n285958 , n285956 , n285957 );
nand ( n285959 , n244987 , n34840 );
nand ( n285960 , n285953 , n285958 , n285959 );
buf ( n285961 , n285960 );
nand ( n285962 , n266576 , n272114 , n273940 );
not ( n285963 , n266572 );
not ( n285964 , n272114 );
or ( n285965 , n285963 , n285964 );
nor ( n285966 , n273940 , n35428 );
nand ( n285967 , n285965 , n285966 );
nand ( n285968 , n48251 , n34792 );
nand ( n285969 , n285962 , n285967 , n285968 );
buf ( n285970 , n285969 );
nor ( n285971 , n284477 , n280580 );
or ( n285972 , n285971 , n259196 );
nand ( n285973 , n285971 , n284468 );
nand ( n285974 , n35431 , n25349 );
nand ( n285975 , n285972 , n285973 , n285974 );
buf ( n285976 , n285975 );
not ( n285977 , n270444 );
nand ( n285978 , n263753 , n244085 );
or ( n285979 , n285977 , n285978 );
not ( n285980 , n263753 );
not ( n285981 , n263751 );
or ( n285982 , n285980 , n285981 );
nor ( n285983 , n244085 , n251361 );
nand ( n285984 , n285982 , n285983 );
nand ( n285985 , n246217 , n25890 );
nand ( n285986 , n285979 , n285984 , n285985 );
buf ( n285987 , n285986 );
or ( n285988 , n25328 , n280108 );
or ( n285989 , n25335 , n283992 );
nand ( n285990 , n285988 , n285989 );
buf ( n285991 , n285990 );
or ( n285992 , n25328 , n284427 );
or ( n285993 , n25335 , n271852 );
nand ( n285994 , n285992 , n285993 );
buf ( n285995 , n285994 );
buf ( n285996 , RI19ad1ee8_2199);
and ( n285997 , n25326 , n285996 );
buf ( n285998 , n285997 );
or ( n285999 , n25328 , n276964 );
or ( n286000 , n25336 , n271941 );
nand ( n286001 , n285999 , n286000 );
buf ( n286002 , n286001 );
not ( n286003 , n255233 );
not ( n286004 , n264495 );
or ( n286005 , n286003 , n286004 );
nor ( n286006 , n255235 , n27889 );
nand ( n286007 , n286005 , n286006 );
nand ( n286008 , n255230 , n264495 , n255235 );
nand ( n286009 , n50615 , n34404 );
nand ( n286010 , n286007 , n286008 , n286009 );
buf ( n286011 , n286010 );
nand ( n286012 , n276023 , n269100 , n257215 );
not ( n286013 , n257202 );
not ( n286014 , n257215 );
or ( n286015 , n286013 , n286014 );
nor ( n286016 , n269100 , n250431 );
nand ( n286017 , n286015 , n286016 );
nand ( n286018 , n245701 , n204591 );
nand ( n286019 , n286012 , n286017 , n286018 );
buf ( n286020 , n286019 );
not ( n286021 , n33038 );
not ( n286022 , n39766 );
or ( n286023 , n286021 , n286022 );
nand ( n286024 , n258675 , n258686 );
and ( n286025 , n286024 , n257633 );
not ( n286026 , n286024 );
and ( n286027 , n286026 , n257632 );
nor ( n286028 , n286025 , n286027 );
or ( n286029 , n286028 , n251498 );
nand ( n286030 , n286023 , n286029 );
buf ( n286031 , n286030 );
not ( n286032 , n251463 );
nand ( n286033 , n273425 , n273435 );
or ( n286034 , n286032 , n286033 );
not ( n286035 , n273435 );
not ( n286036 , n251389 );
or ( n286037 , n286035 , n286036 );
nor ( n286038 , n273425 , n31572 );
nand ( n286039 , n286037 , n286038 );
nand ( n286040 , n247744 , n31301 );
nand ( n286041 , n286034 , n286039 , n286040 );
buf ( n286042 , n286041 );
not ( n286043 , RI19ac36c8_2303);
or ( n286044 , n25328 , n286043 );
or ( n286045 , n25335 , n285089 );
nand ( n286046 , n286044 , n286045 );
buf ( n286047 , n286046 );
or ( n286048 , n25328 , n255191 );
or ( n286049 , n25336 , n273023 );
nand ( n286050 , n286048 , n286049 );
buf ( n286051 , n286050 );
buf ( n286052 , n206630 );
nor ( n286053 , n255129 , n243664 );
or ( n286054 , n284724 , n286053 );
nor ( n286055 , n284723 , n236795 );
nand ( n286056 , n286055 , n286053 );
nand ( n286057 , n241976 , n205306 );
nand ( n286058 , n286054 , n286056 , n286057 );
buf ( n286059 , n286058 );
buf ( n286060 , n33845 );
not ( n286061 , n34293 );
not ( n286062 , n245221 );
or ( n286063 , n286061 , n286062 );
nand ( n286064 , n260560 , n282254 );
not ( n286065 , n278863 );
and ( n286066 , n286064 , n286065 );
not ( n286067 , n286064 );
and ( n286068 , n286067 , n278863 );
nor ( n286069 , n286066 , n286068 );
or ( n286070 , n286069 , n39763 );
nand ( n286071 , n286063 , n286070 );
buf ( n286072 , n286071 );
nand ( n286073 , n258174 , n269381 );
or ( n286074 , n267207 , n286073 );
not ( n286075 , n267199 );
nand ( n286076 , n286075 , n286073 );
nand ( n286077 , n238638 , n31050 );
nand ( n286078 , n286074 , n286076 , n286077 );
buf ( n286079 , n286078 );
nand ( n286080 , n269800 , n270203 );
or ( n286081 , n267541 , n286080 );
nand ( n286082 , n267533 , n286080 );
nand ( n286083 , n233501 , n37148 );
nand ( n286084 , n286081 , n286082 , n286083 );
buf ( n286085 , n286084 );
not ( n286086 , n28685 );
not ( n286087 , n234453 );
or ( n286088 , n286086 , n286087 );
nand ( n286089 , n260404 , n260394 );
not ( n286090 , n263655 );
and ( n286091 , n286089 , n286090 );
not ( n286092 , n286089 );
and ( n286093 , n286092 , n263655 );
nor ( n286094 , n286091 , n286093 );
xor ( n286095 , n286094 , n234818 );
nand ( n286096 , n286088 , n286095 );
buf ( n286097 , n286096 );
not ( n286098 , n234109 );
nand ( n286099 , n286098 , n260930 );
nand ( n286100 , n234309 , n277343 );
xor ( n286101 , n286099 , n286100 );
not ( n286102 , n234309 );
not ( n286103 , n286098 );
xor ( n286104 , n286102 , n286103 );
nor ( n286105 , n277343 , n243204 );
nand ( n286106 , n286104 , n286105 );
nand ( n286107 , n50615 , n41840 );
nand ( n286108 , n286101 , n286106 , n286107 );
buf ( n286109 , n286108 );
not ( n286110 , RI1754b008_49);
xor ( n286111 , n249126 , n286110 );
nand ( n286112 , n249131 , n32598 );
nand ( n286113 , n286111 , n286112 );
buf ( n286114 , n286113 );
xor ( n286115 , n233507 , n264736 );
not ( n286116 , RI19a8ffa8_2683);
xor ( n286117 , n25336 , n286116 );
nand ( n286118 , n286115 , n286117 );
buf ( n286119 , n286118 );
buf ( n286120 , n42459 );
buf ( n286121 , n36508 );
buf ( n286122 , n204708 );
not ( n286123 , n37642 );
not ( n286124 , n245221 );
or ( n286125 , n286123 , n286124 );
not ( n286126 , n279347 );
nand ( n286127 , n204515 , n245840 , n35627 , n35630 );
not ( n286128 , n286127 );
and ( n286129 , n286126 , n286128 );
and ( n286130 , n279347 , n286127 );
nor ( n286131 , n286129 , n286130 );
not ( n286132 , n274416 );
nand ( n286133 , n286132 , n279335 );
and ( n286134 , n286131 , n286133 );
not ( n286135 , n286131 );
not ( n286136 , n286133 );
and ( n286137 , n286135 , n286136 );
nor ( n286138 , n286134 , n286137 );
or ( n286139 , n286138 , n39763 );
nand ( n286140 , n286125 , n286139 );
buf ( n286141 , n286140 );
nand ( n286142 , n259943 , n244535 );
or ( n286143 , n265243 , n286142 );
not ( n286144 , n259943 );
not ( n286145 , n244513 );
or ( n286146 , n286144 , n286145 );
nor ( n286147 , n244535 , n54208 );
nand ( n286148 , n286146 , n286147 );
nand ( n286149 , n234024 , n28256 );
nand ( n286150 , n286143 , n286148 , n286149 );
buf ( n286151 , n286150 );
not ( n286152 , n33426 );
not ( n286153 , n244606 );
or ( n286154 , n286152 , n286153 );
not ( n286155 , RI1754c4a8_5);
or ( n286156 , n244611 , n286155 );
nand ( n286157 , n286154 , n286156 );
buf ( n286158 , n286157 );
nand ( n286159 , n279708 , n279719 );
or ( n286160 , n272708 , n286159 );
not ( n286161 , n279708 );
not ( n286162 , n272707 );
or ( n286163 , n286161 , n286162 );
nor ( n286164 , n279719 , n31571 );
nand ( n286165 , n286163 , n286164 );
nand ( n286166 , n49054 , n29185 );
nand ( n286167 , n286160 , n286165 , n286166 );
buf ( n286168 , n286167 );
not ( n286169 , n274490 );
nand ( n286170 , n286169 , n243438 );
nand ( n286171 , n254815 , n254827 );
or ( n286172 , n286170 , n286171 );
not ( n286173 , n286169 );
not ( n286174 , n254815 );
or ( n286175 , n286173 , n286174 );
nor ( n286176 , n254827 , n40465 );
nand ( n286177 , n286175 , n286176 );
nand ( n286178 , n31577 , n205339 );
nand ( n286179 , n286172 , n286177 , n286178 );
buf ( n286180 , n286179 );
not ( n286181 , n264430 );
nand ( n286182 , n253962 , n264420 , n286181 );
nand ( n286183 , n286181 , n253960 );
nand ( n286184 , n286183 , n285951 , n226010 );
nand ( n286185 , n241976 , n28743 );
nand ( n286186 , n286182 , n286184 , n286185 );
buf ( n286187 , n286186 );
or ( n286188 , n25328 , n283478 );
or ( n286189 , n226822 , n269173 );
nand ( n286190 , n286188 , n286189 );
buf ( n286191 , n286190 );
not ( n286192 , n32661 );
not ( n286193 , n51381 );
or ( n286194 , n286192 , n286193 );
nand ( n286195 , n253980 , n253991 );
and ( n286196 , n286195 , n279473 );
not ( n286197 , n286195 );
and ( n286198 , n286197 , n249400 );
nor ( n286199 , n286196 , n286198 );
or ( n286200 , n286199 , n256376 );
nand ( n286201 , n286194 , n286200 );
buf ( n286202 , n286201 );
not ( n286203 , n40492 );
not ( n286204 , n37728 );
or ( n286205 , n286203 , n286204 );
nand ( n286206 , n275435 , n273315 );
and ( n286207 , n286206 , n282572 );
not ( n286208 , n286206 );
and ( n286209 , n286208 , n278272 );
nor ( n286210 , n286207 , n286209 );
or ( n286211 , n286210 , n260861 );
nand ( n286212 , n286205 , n286211 );
buf ( n286213 , n286212 );
or ( n286214 , n278025 , n253513 );
nor ( n286215 , n253502 , n284093 );
nand ( n286216 , n278039 , n286215 );
and ( n286217 , n284091 , n253502 );
and ( n286218 , n31577 , n29979 );
nor ( n286219 , n286217 , n286218 );
nand ( n286220 , n286214 , n286216 , n286219 );
buf ( n286221 , n286220 );
or ( n286222 , n25335 , n273987 );
or ( n286223 , n255976 , n51365 );
nand ( n286224 , n258655 , RI1754b710_34);
nand ( n286225 , n286222 , n286223 , n286224 );
buf ( n286226 , n286225 );
nor ( n286227 , n259757 , n259733 );
or ( n286228 , n280943 , n286227 );
nand ( n286229 , n282732 , n286227 );
nand ( n286230 , n31577 , n27820 );
nand ( n286231 , n286228 , n286229 , n286230 );
buf ( n286232 , n286231 );
not ( n286233 , n29753 );
not ( n286234 , n46083 );
or ( n286235 , n286233 , n286234 );
nand ( n286236 , n253940 , n253953 );
and ( n286237 , n286236 , n264430 );
not ( n286238 , n286236 );
and ( n286239 , n286238 , n286181 );
nor ( n286240 , n286237 , n286239 );
or ( n286241 , n286240 , n255707 );
nand ( n286242 , n286235 , n286241 );
buf ( n286243 , n286242 );
nand ( n286244 , n282224 , n271499 );
or ( n286245 , n269452 , n286244 );
not ( n286246 , n269451 );
not ( n286247 , n282224 );
or ( n286248 , n286246 , n286247 );
nor ( n286249 , n271499 , n249531 );
nand ( n286250 , n286248 , n286249 );
nand ( n286251 , n254798 , n42261 );
nand ( n286252 , n286245 , n286250 , n286251 );
buf ( n286253 , n286252 );
nand ( n286254 , n266926 , n262659 );
or ( n286255 , n257069 , n286254 );
nand ( n286256 , n257038 , n286254 );
nand ( n286257 , n238638 , n32560 );
nand ( n286258 , n286255 , n286256 , n286257 );
buf ( n286259 , n286258 );
not ( n286260 , n268283 );
nand ( n286261 , n286260 , n269345 );
or ( n286262 , n268272 , n286261 );
not ( n286263 , n286260 );
not ( n286264 , n268271 );
or ( n286265 , n286263 , n286264 );
nor ( n286266 , n269345 , n259801 );
nand ( n286267 , n286265 , n286266 );
nand ( n286268 , n239240 , n39953 );
nand ( n286269 , n286262 , n286267 , n286268 );
buf ( n286270 , n286269 );
not ( n286271 , RI1754a9f0_62);
or ( n286272 , n249125 , n286271 );
or ( n286273 , n25335 , n274344 );
nand ( n286274 , n286272 , n286273 );
buf ( n286275 , n286274 );
not ( n286276 , n262043 );
not ( n286277 , n257347 );
or ( n286278 , n286276 , n286277 );
nand ( n286279 , n257351 , n282088 );
nand ( n286280 , n286278 , n286279 );
buf ( n286281 , n286280 );
nand ( n286282 , n254240 , n275027 );
or ( n286283 , n271391 , n286282 );
nand ( n286284 , n260306 , n286282 );
nand ( n286285 , n246460 , n204943 );
nand ( n286286 , n286283 , n286284 , n286285 );
buf ( n286287 , n286286 );
nand ( n286288 , n278765 , n205649 );
not ( n286289 , n276306 );
nand ( n286290 , n286289 , n278760 );
or ( n286291 , n286288 , n286290 );
nor ( n286292 , n278765 , n234110 );
nand ( n286293 , n286292 , n286290 );
nand ( n286294 , n238114 , n30377 );
nand ( n286295 , n286291 , n286293 , n286294 );
buf ( n286296 , n286295 );
not ( n286297 , RI1754b8f0_30);
or ( n286298 , n229127 , n286297 );
or ( n286299 , n226822 , n282167 );
nand ( n286300 , n286298 , n286299 );
buf ( n286301 , n286300 );
or ( n286302 , n226819 , n281476 );
or ( n286303 , n25335 , n269635 );
nand ( n286304 , n286302 , n286303 );
buf ( n286305 , n286304 );
or ( n286306 , n25328 , n246466 );
not ( n286307 , RI19a8f3f0_2688);
or ( n286308 , n25336 , n286307 );
nand ( n286309 , n286306 , n286308 );
buf ( n286310 , n286309 );
not ( n286311 , n281178 );
nand ( n286312 , n281175 , n271992 );
or ( n286313 , n286311 , n286312 );
not ( n286314 , n281175 );
not ( n286315 , n271967 );
not ( n286316 , n286315 );
or ( n286317 , n286314 , n286316 );
nor ( n286318 , n271992 , n257769 );
nand ( n286319 , n286317 , n286318 );
nand ( n286320 , n31577 , n31884 );
nand ( n286321 , n286313 , n286319 , n286320 );
buf ( n286322 , n286321 );
nor ( n286323 , n283419 , n273238 );
not ( n286324 , n286323 );
nand ( n286325 , n273239 , n273566 );
nand ( n286326 , n283421 , n273238 , n278443 );
nand ( n286327 , n251712 , n205423 );
nand ( n286328 , n286324 , n286325 , n286326 , n286327 );
buf ( n286329 , n286328 );
buf ( n286330 , RI17538c00_591);
and ( n286331 , n27883 , n286330 );
buf ( n286332 , n286331 );
or ( n286333 , n25328 , n271701 );
or ( n286334 , n226822 , n285623 );
nand ( n286335 , n286333 , n286334 );
buf ( n286336 , n286335 );
nand ( n286337 , n253274 , n253307 );
or ( n286338 , n267582 , n286337 );
not ( n286339 , n253274 );
not ( n286340 , n267581 );
or ( n286341 , n286339 , n286340 );
nor ( n286342 , n253307 , n226003 );
nand ( n286343 , n286341 , n286342 );
nand ( n286344 , n238638 , n28795 );
nand ( n286345 , n286338 , n286343 , n286344 );
buf ( n286346 , n286345 );
nand ( n286347 , n265176 , n278101 );
or ( n286348 , n265191 , n286347 );
not ( n286349 , n265176 );
not ( n286350 , n265194 );
or ( n286351 , n286349 , n286350 );
nand ( n286352 , n286351 , n284964 );
nand ( n286353 , n31576 , n27712 );
nand ( n286354 , n286348 , n286352 , n286353 );
buf ( n286355 , n286354 );
not ( n286356 , n262157 );
nand ( n286357 , n286356 , n280524 );
nand ( n286358 , n280524 , n283088 );
not ( n286359 , n286358 );
not ( n286360 , n262180 );
and ( n286361 , n286359 , n286360 );
and ( n286362 , n51381 , n206656 );
nor ( n286363 , n286361 , n286362 );
nor ( n286364 , n280524 , n262179 );
nand ( n286365 , n267233 , n286364 );
nand ( n286366 , n286357 , n286363 , n286365 );
buf ( n286367 , n286366 );
nand ( n286368 , n259802 , n246894 , n249762 );
not ( n286369 , n249772 );
not ( n286370 , n286369 );
not ( n286371 , n249762 );
or ( n286372 , n286370 , n286371 );
nor ( n286373 , n246894 , n238635 );
nand ( n286374 , n286372 , n286373 );
nand ( n286375 , n237714 , n44915 );
nand ( n286376 , n286368 , n286374 , n286375 );
buf ( n286377 , n286376 );
nand ( n286378 , n270732 , n259847 );
nand ( n286379 , n242869 , n277874 );
or ( n286380 , n286378 , n286379 );
not ( n286381 , n277874 );
not ( n286382 , n270732 );
or ( n286383 , n286381 , n286382 );
nor ( n286384 , n242869 , n54208 );
nand ( n286385 , n286383 , n286384 );
nand ( n286386 , n237361 , n37099 );
nand ( n286387 , n286380 , n286385 , n286386 );
buf ( n286388 , n286387 );
nor ( n286389 , n283267 , n254509 );
nand ( n286390 , n260448 , n286389 );
nor ( n286391 , n283268 , n247276 );
and ( n286392 , n260446 , n254510 );
and ( n286393 , n286391 , n286392 );
and ( n286394 , n258743 , n36918 );
and ( n286395 , n286390 , n286393 , n286394 );
buf ( n286396 , n286395 );
not ( n286397 , n243234 );
and ( n286398 , n286397 , n243269 , n263588 );
and ( n286399 , n263588 , n243232 );
and ( n286400 , n286399 , n243267 , n253393 );
and ( n286401 , n39767 , n30030 );
and ( n286402 , n286398 , n286400 , n286401 );
buf ( n286403 , n286402 );
not ( n286404 , RI19a8b958_2714);
or ( n286405 , n25328 , n286404 );
or ( n286406 , n25335 , n261251 );
nand ( n286407 , n286405 , n286406 );
buf ( n286408 , n286407 );
nand ( n286409 , n284901 , n239934 );
nand ( n286410 , n284903 , n280308 );
or ( n286411 , n286409 , n286410 );
not ( n286412 , n284903 );
not ( n286413 , n284901 );
or ( n286414 , n286412 , n286413 );
nor ( n286415 , n280308 , n238900 );
nand ( n286416 , n286414 , n286415 );
nand ( n286417 , n254798 , n205663 );
nand ( n286418 , n286411 , n286416 , n286417 );
buf ( n286419 , n286418 );
nand ( n286420 , n269004 , n254465 );
or ( n286421 , n286420 , n244630 );
nand ( n286422 , n286420 , n275188 );
nand ( n286423 , n31577 , n29132 );
nand ( n286424 , n286421 , n286422 , n286423 );
buf ( n286425 , n286424 );
buf ( n286426 , RI19ad0958_2207);
and ( n286427 , n25326 , n286426 );
buf ( n286428 , n286427 );
nor ( n286429 , n229370 , n54332 );
not ( n286430 , n286429 );
not ( n286431 , n267347 );
or ( n286432 , n286430 , n286431 );
nand ( n286433 , n54209 , n229370 );
nand ( n286434 , n286432 , n286433 );
not ( n286435 , n286434 );
not ( n286436 , n267343 );
nor ( n286437 , n286436 , n258369 );
nand ( n286438 , n286437 , n54332 );
nand ( n286439 , n247585 , n38883 );
nand ( n286440 , n286435 , n286438 , n286439 );
buf ( n286441 , n286440 );
nand ( n286442 , n256628 , n244393 );
nand ( n286443 , n278673 , n281545 );
or ( n286444 , n286442 , n286443 );
not ( n286445 , n281545 );
not ( n286446 , n256628 );
or ( n286447 , n286445 , n286446 );
nor ( n286448 , n278673 , n258327 );
nand ( n286449 , n286447 , n286448 );
nand ( n286450 , n37728 , n46900 );
nand ( n286451 , n286444 , n286449 , n286450 );
buf ( n286452 , n286451 );
nor ( n286453 , n276183 , n252658 );
or ( n286454 , n250112 , n286453 );
nor ( n286455 , n250110 , n40465 );
nand ( n286456 , n286455 , n286453 );
nand ( n286457 , n35431 , n25732 );
nand ( n286458 , n286454 , n286456 , n286457 );
buf ( n286459 , n286458 );
not ( n286460 , n30753 );
not ( n286461 , n255116 );
or ( n286462 , n286460 , n286461 );
nand ( n286463 , n273708 , n278123 );
not ( n286464 , n270256 );
and ( n286465 , n286463 , n286464 );
not ( n286466 , n286463 );
and ( n286467 , n286466 , n270256 );
nor ( n286468 , n286465 , n286467 );
or ( n286469 , n286468 , n31572 );
nand ( n286470 , n286462 , n286469 );
buf ( n286471 , n286470 );
buf ( n286472 , n34684 );
buf ( n286473 , n32615 );
nand ( n286474 , n272821 , n272808 );
not ( n286475 , n275858 );
or ( n286476 , n286474 , n286475 );
not ( n286477 , n272808 );
not ( n286478 , n275840 );
or ( n286479 , n286477 , n286478 );
nand ( n286480 , n286479 , n248981 );
or ( n286481 , n286480 , n272821 );
nand ( n286482 , n46083 , n240635 );
nand ( n286483 , n286476 , n286481 , n286482 );
buf ( n286484 , n286483 );
buf ( n286485 , n36440 );
not ( n286486 , n34412 );
not ( n286487 , n234453 );
or ( n286488 , n286486 , n286487 );
not ( n286489 , n272141 );
not ( n286490 , n275254 );
nand ( n286491 , n286489 , n286490 );
and ( n286492 , n286491 , n272151 );
not ( n286493 , n286491 );
and ( n286494 , n286493 , n272152 );
nor ( n286495 , n286492 , n286494 );
or ( n286496 , n286495 , n264257 );
nand ( n286497 , n286488 , n286496 );
buf ( n286498 , n286497 );
not ( n286499 , RI19aa7a68_2512);
or ( n286500 , n25328 , n286499 );
or ( n286501 , n25336 , n269534 );
nand ( n286502 , n286500 , n286501 );
buf ( n286503 , n286502 );
nand ( n286504 , n275947 , n259980 );
and ( n286505 , n286504 , n271224 , n226010 );
not ( n286506 , n209798 );
nor ( n286507 , n286506 , n263991 );
nor ( n286508 , n286505 , n286507 );
nor ( n286509 , n275950 , n244399 );
nand ( n286510 , n286509 , n271223 , n259980 );
nand ( n286511 , n286508 , n286510 );
buf ( n286512 , n286511 );
nand ( n286513 , n280613 , n279996 );
not ( n286514 , n282727 );
or ( n286515 , n286513 , n286514 );
not ( n286516 , n280627 );
not ( n286517 , n280613 );
or ( n286518 , n286516 , n286517 );
nor ( n286519 , n279996 , n251862 );
nand ( n286520 , n286518 , n286519 );
nand ( n286521 , n51381 , n29590 );
nand ( n286522 , n286515 , n286520 , n286521 );
buf ( n286523 , n286522 );
not ( n286524 , n256322 );
nand ( n286525 , n286524 , n275100 );
or ( n286526 , n284131 , n286525 );
not ( n286527 , n284130 );
not ( n286528 , n286524 );
or ( n286529 , n286527 , n286528 );
nor ( n286530 , n275100 , n55152 );
nand ( n286531 , n286529 , n286530 );
nand ( n286532 , n241976 , n38109 );
nand ( n286533 , n286526 , n286531 , n286532 );
buf ( n286534 , n286533 );
not ( n286535 , n28012 );
not ( n286536 , n37728 );
or ( n286537 , n286535 , n286536 );
nand ( n286538 , n244969 , n268537 );
and ( n286539 , n286538 , n268119 );
not ( n286540 , n286538 );
and ( n286541 , n286540 , n268120 );
nor ( n286542 , n286539 , n286541 );
or ( n286543 , n286542 , n254882 );
nand ( n286544 , n286537 , n286543 );
buf ( n286545 , n286544 );
or ( n286546 , n25328 , n280965 );
or ( n286547 , n25335 , n282500 );
nand ( n286548 , n286546 , n286547 );
buf ( n286549 , n286548 );
or ( n286550 , n226819 , n272874 );
or ( n286551 , n226822 , n286499 );
nand ( n286552 , n286550 , n286551 );
buf ( n286553 , n286552 );
not ( n286554 , n284875 );
nor ( n286555 , n266323 , n273198 );
or ( n286556 , n286554 , n286555 );
nand ( n286557 , n266311 , n286555 );
nand ( n286558 , n31577 , n216949 );
nand ( n286559 , n286556 , n286557 , n286558 );
buf ( n286560 , n286559 );
nand ( n286561 , n275123 , n250582 );
or ( n286562 , n275112 , n286561 );
not ( n286563 , n275123 );
not ( n286564 , n250503 );
or ( n286565 , n286563 , n286564 );
nand ( n286566 , n286565 , n280601 );
nand ( n286567 , n250916 , n36614 );
nand ( n286568 , n286562 , n286566 , n286567 );
buf ( n286569 , n286568 );
nand ( n286570 , n285038 , n255007 );
nand ( n286571 , n286570 , n44767 , n205649 );
nand ( n286572 , n255015 , n44766 , n285038 );
nand ( n286573 , n234024 , n36948 );
nand ( n286574 , n286571 , n286572 , n286573 );
buf ( n286575 , n286574 );
or ( n286576 , n25328 , n279512 );
not ( n286577 , RI19a8c240_2710);
or ( n286578 , n25335 , n286577 );
nand ( n286579 , n286576 , n286578 );
buf ( n286580 , n286579 );
endmodule

