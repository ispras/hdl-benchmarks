//NOTE: no-implementation module stub

module IDEBN (
    input wire ICK,
    input wire nSTBx,
    output reg nSTB
);

endmodule
