//
// Conformal-LEC Version 15.10-d003 ( 23-Apr-2015) ( 64 bit executable)
//
module top ( 
    n0 , 
    n1 , 
    n2 , 
    n3 , 
    n4 , 
    n5 , 
    n6 , 
    n7 , 
    n8 , 
    n9 , 
    n10 , 
    n11 , 
    n12 , 
    n13 , 
    n14 , 
    n15 , 
    n16 , 
    n17 , 
    n18 , 
    n19 , 
    n20 , 
    n21 , 
    n22 , 
    n23 , 
    n24 , 
    n25 , 
    n26 , 
    n27 , 
    n28 , 
    n29 , 
    n30 , 
    n31 , 
    n32 , 
    n33 , 
    n34 , 
    n35 , 
    n36 , 
    n37 , 
    n38 , 
    n39 , 
    n40 , 
    n41 , 
    n42 , 
    n43 , 
    n44 , 
    n45 , 
    n46 , 
    n47 , 
    n48 , 
    n49 , 
    n50 , 
    n51 , 
    n52 , 
    n53 , 
    n54 , 
    n55 , 
    n56 , 
    n57 , 
    n58 , 
    n59 , 
    n60 , 
    n61 , 
    n62 , 
    n63 , 
    n64 , 
    n65 , 
    n66 , 
    n67 , 
    n68 , 
    n69 , 
    n70 , 
    n71 , 
    n72 , 
    n73 , 
    n74 , 
    n75 , 
    n76 , 
    n77 , 
    n78 , 
    n79 , 
    n80 , 
    n81 , 
    n82 , 
    n83 , 
    n84 , 
    n85 , 
    n86 , 
    n87 , 
    n88 , 
    n89 , 
    n90 , 
    n91 , 
    n92 , 
    n93 , 
    n94 , 
    n95 , 
    n96 , 
    n97 , 
    n98 , 
    n99 , 
    n100 , 
    n101 , 
    n102 , 
    n103 , 
    n104 , 
    n105 , 
    n106 , 
    n107 , 
    n108 , 
    n109 , 
    n110 , 
    n111 , 
    n112 , 
    n113 , 
    n114 , 
    n115 , 
    n116 , 
    n117 , 
    n118 , 
    n119 , 
    n120 , 
    n121 , 
    n122 , 
    n123 , 
    n124 , 
    n125 , 
    n126 , 
    n127 , 
    n128 , 
    n129 , 
    n130 , 
    n131 , 
    n132 , 
    n133 , 
    n134 , 
    n135 , 
    n136 , 
    n137 , 
    n138 , 
    n139 , 
    n140 , 
    n141 , 
    n142 , 
    n143 , 
    n144 , 
    n145 , 
    n146 , 
    n147 , 
    n148 , 
    n149 , 
    n150 , 
    n151 , 
    n152 , 
    n153 , 
    n154 , 
    n155 , 
    n156 , 
    n157 , 
    n158 , 
    n159 , 
    n160 , 
    n161 , 
    n162 , 
    n163 , 
    n164 , 
    n165 , 
    n166 , 
    n167 , 
    n168 , 
    n169 , 
    n170 , 
    n171 , 
    n172 , 
    n173 , 
    n174 , 
    n175 , 
    n176 , 
    n177 , 
    n178 , 
    n179 , 
    n180 , 
    n181 , 
    n182 , 
    n183 , 
    n184 , 
    n185 , 
    n186 , 
    n187 , 
    n188 , 
    n189 , 
    n190 , 
    n191 , 
    n192 , 
    n193 , 
    n194 , 
    n195 , 
    n196 , 
    n197 , 
    n198 , 
    n199 , 
    n200 , 
    n201 , 
    n202 , 
    n203 , 
    n204 , 
    n205 , 
    n206 , 
    n207 , 
    n208 , 
    n209 , 
    n210 , 
    n211 , 
    n212 , 
    n213 , 
    n214 , 
    n215 , 
    n216 , 
    n217 , 
    n218 , 
    n219 , 
    n220 , 
    n221 , 
    n222 , 
    n223 , 
    n224 , 
    n225 , 
    n226 , 
    n227 , 
    n228 , 
    n229 , 
    n230 , 
    n231 , 
    n232 , 
    n233 , 
    n234 , 
    n235 , 
    n236 , 
    n237 , 
    n238 , 
    n239 , 
    n240 , 
    n241 , 
    n242 , 
    n243 , 
    n244 , 
    n245 , 
    n246 , 
    n247 , 
    n248 , 
    n249 , 
    n250 , 
    n251 , 
    n252 , 
    n253 , 
    n254 , 
    n255 , 
    n256 , 
    n257 , 
    n258 , 
    n259 , 
    n260 , 
    n261 , 
    n262 , 
    n263 , 
    n264 , 
    n265 , 
    n266 , 
    n267 , 
    n268 , 
    n269 , 
    n270 , 
    n271 , 
    n272 , 
    n273 , 
    n274 , 
    n275 , 
    n276 , 
    n277 , 
    n278 , 
    n279 , 
    n280 , 
    n281 , 
    n282 , 
    n283 , 
    n284 , 
    n285 , 
    n286 , 
    n287 , 
    n288 , 
    n289 , 
    n290 , 
    n291 , 
    n292 , 
    n293 , 
    n294 , 
    n295 , 
    n296 , 
    n297 , 
    n298 , 
    n299 , 
    n300 , 
    n301 , 
    n302 , 
    n303 , 
    n304 , 
    n305 , 
    n306 , 
    n307 , 
    n308 , 
    n309 , 
    n310 , 
    n311 , 
    n312 , 
    n313 , 
    n314 , 
    n315 , 
    n316 , 
    n317 , 
    n318 , 
    n319 , 
    n320 , 
    n321 , 
    n322 , 
    n323 , 
    n324 , 
    n325 , 
    n326 , 
    n327 , 
    n328 , 
    n329 , 
    n330 , 
    n331 , 
    n332 , 
    n333 , 
    n334 , 
    n335 , 
    n336 , 
    n337 , 
    n338 , 
    n339 , 
    n340 , 
    n341 , 
    n342 , 
    n343 , 
    n344 , 
    n345 , 
    n346 , 
    n347 , 
    n348 , 
    n349 , 
    n350 , 
    n351 , 
    n352 , 
    n353 , 
    n354 , 
    n355 , 
    n356 , 
    n357 , 
    n358 , 
    n359 , 
    n360 , 
    n361 , 
    n362 , 
    n363 , 
    n364 , 
    n365 , 
    n366 , 
    n367 , 
    n368 , 
    n369 , 
    n370 , 
    n371 , 
    n372 , 
    n373 , 
    n374 , 
    n375 , 
    n376 , 
    n377 , 
    n378 , 
    n379 , 
    n380 , 
    n381 , 
    n382 , 
    n383 , 
    n384 , 
    n385 , 
    n386 , 
    n387 , 
    n388 , 
    n389 , 
    n390 , 
    n391 , 
    n392 , 
    n393 , 
    n394 , 
    n395 , 
    n396 , 
    n397 , 
    n398 , 
    n399 , 
    n400 , 
    n401 , 
    n402 , 
    n403 , 
    n404 , 
    n405 , 
    n406 , 
    n407 , 
    n408 , 
    n409 , 
    n410 , 
    n411 , 
    n412 , 
    n413 , 
    n414 , 
    n415 , 
    n416 , 
    n417 , 
    n418 , 
    n419 , 
    n420 , 
    n421 , 
    n422 , 
    n423 , 
    n424 , 
    n425 , 
    n426 , 
    n427 , 
    n428 , 
    n429 , 
    n430 , 
    n431 , 
    n432 , 
    n433 , 
    n434 , 
    n435 , 
    n436 , 
    n437 , 
    n438 , 
    n439 , 
    n440 , 
    n441 , 
    n442 , 
    n443 , 
    n444 , 
    n445 , 
    n446 , 
    n447 , 
    n448 , 
    n449 , 
    n450 , 
    n451 , 
    n452 , 
    n453 , 
    n454 , 
    n455 , 
    n456 , 
    n457 , 
    n458 , 
    n459 , 
    n460 , 
    n461 , 
    n462 , 
    n463 , 
    n464 , 
    n465 , 
    n466 , 
    n467 , 
    n468 , 
    n469 , 
    n470 , 
    n471 , 
    n472 , 
    n473 , 
    n474 , 
    n475 , 
    n476 , 
    n477 , 
    n478 , 
    n479 , 
    n480 , 
    n481 , 
    n482 , 
    n483 , 
    n484 , 
    n485 , 
    n486 , 
    n487 , 
    n488 , 
    n489 , 
    n490 , 
    n491 , 
    n492 , 
    n493 , 
    n494 , 
    n495 , 
    n496 , 
    n497 , 
    n498 , 
    n499 , 
    n500 , 
    n501 , 
    n502 , 
    n503 , 
    n504 , 
    n505 , 
    n506 , 
    n507 , 
    n508 , 
    n509 , 
    n510 , 
    n511 , 
    n512 , 
    n513 , 
    n514 , 
    n515 , 
    n516 , 
    n517 , 
    n518 , 
    n519 , 
    n520 , 
    n521 , 
    n522 , 
    n523 , 
    n524 , 
    n525 , 
    n526 , 
    n527 , 
    n528 , 
    n529 , 
    n530 , 
    n531 , 
    n532 , 
    n533 , 
    n534 , 
    n535 , 
    n536 , 
    n537 , 
    n538 , 
    n539 , 
    n540 , 
    n541 , 
    n542 , 
    n543 , 
    n544 , 
    n545 , 
    n546 , 
    n547 , 
    n548 , 
    n549 , 
    n550 , 
    n551 , 
    n552 , 
    n553 , 
    n554 , 
    n555 , 
    n556 , 
    n557 , 
    n558 , 
    n559 , 
    n560 , 
    n561 , 
    n562 , 
    n563 , 
    n564 , 
    n565 , 
    n566 , 
    n567 , 
    n568 , 
    n569 , 
    n570 , 
    n571 , 
    n572 , 
    n573 , 
    n574 , 
    n575 , 
    n576 , 
    n577 , 
    n578 , 
    n579 , 
    n580 , 
    n581 , 
    n582 , 
    n583 , 
    n584 , 
    n585 , 
    n586 , 
    n587 , 
    n588 , 
    n589 , 
    n590 , 
    n591 , 
    n592 , 
    n593 , 
    n594 , 
    n595 , 
    n596 , 
    n597 , 
    n598 , 
    n599 , 
    n600 , 
    n601 , 
    n602 , 
    n603 , 
    n604 , 
    n605 , 
    n606 , 
    n607 , 
    n608 , 
    n609 , 
    n610 , 
    n611 , 
    n612 , 
    n613 , 
    n614 , 
    n615 , 
    n616 , 
    n617 , 
    n618 , 
    n619 , 
    n620 , 
    n621 , 
    n622 , 
    n623 , 
    n624 , 
    n625 , 
    n626 , 
    n627 , 
    n628 , 
    n629 , 
    n630 , 
    n631 , 
    n632 , 
    n633 , 
    n634 , 
    n635 , 
    n636 , 
    n637 , 
    n638 , 
    n639 , 
    n640 , 
    n641 , 
    n642 , 
    n643 , 
    n644 , 
    n645 , 
    n646 , 
    n647 , 
    n648 , 
    n649 , 
    n650 , 
    n651 , 
    n652 , 
    n653 , 
    n654 , 
    n655 , 
    n656 , 
    n657 , 
    n658 , 
    n659 , 
    n660 , 
    n661 , 
    n662 , 
    n663 , 
    n664 , 
    n665 , 
    n666 , 
    n667 , 
    n668 , 
    n669 , 
    n670 , 
    n671 , 
    n672 , 
    n673 , 
    n674 , 
    n675 , 
    n676 , 
    n677 , 
    n678 , 
    n679 , 
    n680 , 
    n681 , 
    n682 , 
    n683 , 
    n684 , 
    n685 , 
    n686 , 
    n687 , 
    n688 , 
    n689 , 
    n690 , 
    n691 , 
    n692 , 
    n693 , 
    n694 , 
    n695 , 
    n696 , 
    n697 , 
    n698 , 
    n699 , 
    n700 , 
    n701 , 
    n702 , 
    n703 , 
    n704 , 
    n705 , 
    n706 , 
    n707 , 
    n708 , 
    n709 , 
    n710 , 
    n711 , 
    n712 , 
    n713 , 
    n714 , 
    n715 , 
    n716 , 
    n717 , 
    n718 , 
    n719 , 
    n720 , 
    n721 , 
    n722 , 
    n723 , 
    n724 , 
    n725 , 
    n726 , 
    n727 , 
    n728 , 
    n729 , 
    n730 , 
    n731 , 
    n732 , 
    n733 , 
    n734 , 
    n735 , 
    n736 , 
    n737 , 
    n738 , 
    n739 , 
    n740 , 
    n741 , 
    n742 , 
    n743 , 
    n744 , 
    n745 , 
    n746 , 
    n747 , 
    n748 , 
    n749 , 
    n750 , 
    n751 , 
    n752 , 
    n753 , 
    n754 , 
    n755 , 
    n756 , 
    n757 , 
    n758 , 
    n759 , 
    n760 , 
    n761 , 
    n762 , 
    n763 , 
    n764 , 
    n765 , 
    n766 , 
    n767 , 
    n768 , 
    n769 , 
    n770 , 
    n771 , 
    n772 , 
    n773 , 
    n774 , 
    n775 , 
    n776 , 
    n777 , 
    n778 , 
    n779 , 
    n780 , 
    n781 , 
    n782 , 
    n783 , 
    n784 , 
    n785 , 
    n786 , 
    n787 , 
    n788 , 
    n789 , 
    n790 , 
    n791 , 
    n792 , 
    n793 , 
    n794 , 
    n795 , 
    n796 , 
    n797 , 
    n798 , 
    n799 , 
    n800 , 
    n801 , 
    n802 , 
    n803 , 
    n804 , 
    n805 , 
    n806 , 
    n807 , 
    n808 , 
    n809 , 
    n810 , 
    n811 , 
    n812 , 
    n813 , 
    n814 , 
    n815 , 
    n816 , 
    n817 , 
    n818 , 
    n819 , 
    n820 , 
    n821 , 
    n822 , 
    n823 , 
    n824 , 
    n825 , 
    n826 , 
    n827 , 
    n828 , 
    n829 , 
    n830 , 
    n831 , 
    n832 , 
    n833 , 
    n834 , 
    n835 , 
    n836 , 
    n837 , 
    n838 , 
    n839 , 
    n840 , 
    n841 , 
    n842 , 
    n843 , 
    n844 , 
    n845 , 
    n846 , 
    n847 , 
    n848 , 
    n849 , 
    n850 , 
    n851 , 
    n852 , 
    n853 , 
    n854 , 
    n855 , 
    n856 , 
    n857 , 
    n858 , 
    n859 , 
    n860 , 
    n861 , 
    n862 , 
    n863 , 
    n864 , 
    n865 , 
    n866 , 
    n867 , 
    n868 , 
    n869 , 
    n870 , 
    n871 , 
    n872 , 
    n873 , 
    n874 , 
    n875 , 
    n876 , 
    n877 , 
    n878 , 
    n879 , 
    n880 , 
    n881 , 
    n882 , 
    n883 , 
    n884 , 
    n885 , 
    n886 , 
    n887 , 
    n888 , 
    n889 , 
    n890 , 
    n891 , 
    n892 , 
    n893 , 
    n894 , 
    n895 , 
    n896 , 
    n897 , 
    n898 , 
    n899 , 
    n900 , 
    n901 , 
    n902 , 
    n903 , 
    n904 , 
    n905 , 
    n906 , 
    n907 , 
    n908 , 
    n909 , 
    n910 , 
    n911 , 
    n912 , 
    n913 , 
    n914 , 
    n915 , 
    n916 , 
    n917 , 
    n918 , 
    n919 , 
    n920 , 
    n921 , 
    n922 , 
    n923 , 
    n924 , 
    n925 , 
    n926 , 
    n927 , 
    n928 , 
    n929 , 
    n930 , 
    n931 , 
    n932 , 
    n933 , 
    n934 , 
    n935 , 
    n936 , 
    n937 , 
    n938 , 
    n939 , 
    n940 , 
    n941 , 
    n942 , 
    n943 , 
    n944 , 
    n945 , 
    n946 , 
    n947 , 
    n948 , 
    n949 , 
    n950 , 
    n951 , 
    n952 , 
    n953 , 
    n954 , 
    n955 , 
    n956 , 
    n957 , 
    n958 , 
    n959 , 
    n960 , 
    n961 , 
    n962 , 
    n963 , 
    n964 , 
    n965 , 
    n966 , 
    n967 , 
    n968 , 
    n969 , 
    n970 , 
    n971 , 
    n972 , 
    n973 , 
    n974 , 
    n975 , 
    n976 , 
    n977 , 
    n978 , 
    n979 , 
    n980 , 
    n981 , 
    n982 , 
    n983 , 
    n984 , 
    n985 , 
    n986 , 
    n987 , 
    n988 , 
    n989 , 
    n990 , 
    n991 , 
    n992 , 
    n993 , 
    n994 , 
    n995 , 
    n996 , 
    n997 , 
    n998 , 
    n999 , 
    n1000 , 
    n1001 , 
    n1002 , 
    n1003 , 
    n1004 , 
    n1005 , 
    n1006 , 
    n1007 , 
    n1008 , 
    n1009 , 
    n1010 , 
    n1011 , 
    n1012 , 
    n1013 , 
    n1014 , 
    n1015 , 
    n1016 , 
    n1017 , 
    n1018 , 
    n1019 , 
    n1020 , 
    n1021 , 
    n1022 , 
    n1023 , 
    n1024 , 
    n1025 , 
    n1026 , 
    n1027 , 
    n1028 , 
    n1029 , 
    n1030 , 
    n1031 , 
    n1032 , 
    n1033 , 
    n1034 , 
    n1035 , 
    n1036 , 
    n1037 , 
    n1038 , 
    n1039 , 
    n1040 , 
    n1041 , 
    n1042 , 
    n1043 , 
    n1044 , 
    n1045 , 
    n1046 , 
    n1047 , 
    n1048 , 
    n1049 , 
    n1050 , 
    n1051 , 
    n1052 , 
    n1053 , 
    n1054 , 
    n1055 , 
    n1056 , 
    n1057 , 
    n1058 , 
    n1059 , 
    n1060 , 
    n1061 , 
    n1062 , 
    n1063 , 
    n1064 , 
    n1065 , 
    n1066 , 
    n1067 , 
    n1068 , 
    n1069 , 
    n1070 , 
    n1071 , 
    n1072 , 
    n1073 , 
    n1074 , 
    n1075 , 
    n1076 , 
    n1077 , 
    n1078 , 
    n1079 , 
    n1080 , 
    n1081 , 
    n1082 , 
    n1083 , 
    n1084 , 
    n1085 , 
    n1086 , 
    n1087 , 
    n1088 , 
    n1089 , 
    n1090 , 
    n1091 , 
    n1092 , 
    n1093 , 
    n1094 , 
    n1095 , 
    n1096 , 
    n1097 , 
    n1098 , 
    n1099 , 
    n1100 , 
    n1101 , 
    n1102 , 
    n1103 , 
    n1104 , 
    n1105 , 
    n1106 , 
    n1107 , 
    n1108 , 
    n1109 , 
    n1110 , 
    n1111 , 
    n1112 , 
    n1113 , 
    n1114 , 
    n1115 , 
    n1116 , 
    n1117 , 
    n1118 , 
    n1119 , 
    n1120 , 
    n1121 , 
    n1122 , 
    n1123 , 
    n1124 , 
    n1125 , 
    n1126 , 
    n1127 , 
    n1128 , 
    n1129 , 
    n1130 , 
    n1131 , 
    n1132 , 
    n1133 , 
    n1134 , 
    n1135 , 
    n1136 , 
    n1137 , 
    n1138 , 
    n1139 , 
    n1140 , 
    n1141 , 
    n1142 , 
    n1143 , 
    n1144 , 
    n1145 , 
    n1146 , 
    n1147 , 
    n1148 , 
    n1149 , 
    n1150 , 
    n1151 , 
    n1152 , 
    n1153 , 
    n1154 , 
    n1155 , 
    n1156 , 
    n1157 , 
    n1158 , 
    n1159 , 
    n1160 , 
    n1161 , 
    n1162 , 
    n1163 , 
    n1164 , 
    n1165 , 
    n1166 , 
    n1167 , 
    n1168 , 
    n1169 , 
    n1170 , 
    n1171 , 
    n1172 , 
    n1173 , 
    n1174 , 
    n1175 , 
    n1176 , 
    n1177 , 
    n1178 , 
    n1179 , 
    n1180 , 
    n1181 , 
    n1182 , 
    n1183 , 
    n1184 , 
    n1185 , 
    n1186 , 
    n1187 , 
    n1188 , 
    n1189 , 
    n1190 , 
    n1191 , 
    n1192 , 
    n1193 , 
    n1194 , 
    n1195 , 
    n1196 , 
    n1197 , 
    n1198 , 
    n1199 , 
    n1200 , 
    n1201 , 
    n1202 , 
    n1203 , 
    n1204 , 
    n1205 , 
    n1206 , 
    n1207 , 
    n1208 , 
    n1209 , 
    n1210 , 
    n1211 , 
    n1212 , 
    n1213 , 
    n1214 , 
    n1215 , 
    n1216 , 
    n1217 , 
    n1218 , 
    n1219 , 
    n1220 , 
    n1221 , 
    n1222 , 
    n1223 , 
    n1224 , 
    n1225 , 
    n1226 , 
    n1227 , 
    n1228 , 
    n1229 , 
    n1230 , 
    n1231 , 
    n1232 , 
    n1233 , 
    n1234 , 
    n1235 , 
    n1236 , 
    n1237 , 
    n1238 , 
    n1239 , 
    n1240 , 
    n1241 , 
    n1242 , 
    n1243 , 
    n1244 , 
    n1245 , 
    n1246 , 
    n1247 , 
    n1248 , 
    n1249 , 
    n1250 , 
    n1251 , 
    n1252 , 
    n1253 , 
    n1254 , 
    n1255 , 
    n1256 , 
    n1257 , 
    n1258 , 
    n1259 , 
    n1260 , 
    n1261 , 
    n1262 , 
    n1263 , 
    n1264 , 
    n1265 , 
    n1266 , 
    n1267 , 
    n1268 , 
    n1269 , 
    n1270 , 
    n1271 , 
    n1272 , 
    n1273 , 
    n1274 , 
    n1275 , 
    n1276 , 
    n1277 , 
    n1278 , 
    n1279 , 
    n1280 , 
    n1281 , 
    n1282 , 
    n1283 , 
    n1284 , 
    n1285 , 
    n1286 , 
    n1287 , 
    n1288 , 
    n1289 , 
    n1290 , 
    n1291 , 
    n1292 , 
    n1293 , 
    n1294 , 
    n1295 , 
    n1296 , 
    n1297 , 
    n1298 , 
    n1299 , 
    n1300 , 
    n1301 , 
    n1302 , 
    n1303 , 
    n1304 , 
    n1305 , 
    n1306 , 
    n1307 , 
    n1308 , 
    n1309 , 
    n1310 , 
    n1311 , 
    n1312 , 
    n1313 , 
    n1314 , 
    n1315 , 
    n1316 , 
    n1317 , 
    n1318 , 
    n1319 , 
    n1320 , 
    n1321 , 
    n1322 , 
    n1323 , 
    n1324 , 
    n1325 , 
    n1326 , 
    n1327 , 
    n1328 , 
    n1329 , 
    n1330 , 
    n1331 , 
    n1332 , 
    n1333 , 
    n1334 , 
    n1335 , 
    n1336 , 
    n1337 , 
    n1338 , 
    n1339 , 
    n1340 , 
    n1341 , 
    n1342 , 
    n1343 , 
    n1344 , 
    n1345 , 
    n1346 , 
    n1347 , 
    n1348 , 
    n1349 , 
    n1350 , 
    n1351 , 
    n1352 , 
    n1353 , 
    n1354 , 
    n1355 , 
    n1356 , 
    n1357 , 
    n1358 , 
    n1359 , 
    n1360 , 
    n1361 , 
    n1362 , 
    n1363 , 
    n1364 , 
    n1365 , 
    n1366 , 
    n1367 , 
    n1368 , 
    n1369 , 
    n1370 , 
    n1371 , 
    n1372 , 
    n1373 , 
    n1374 , 
    n1375 , 
    n1376 , 
    n1377 , 
    n1378 , 
    n1379 , 
    n1380 , 
    n1381 , 
    n1382 , 
    n1383 , 
    n1384 , 
    n1385 , 
    n1386 , 
    n1387 , 
    n1388 , 
    n1389 , 
    n1390 , 
    n1391 , 
    n1392 , 
    n1393 , 
    n1394 , 
    n1395 , 
    n1396 , 
    n1397 , 
    n1398 , 
    n1399 , 
    n1400 , 
    n1401 , 
    n1402 , 
    n1403 , 
    n1404 , 
    n1405 , 
    n1406 , 
    n1407 , 
    n1408 , 
    n1409 , 
    n1410 , 
    n1411 , 
    n1412 , 
    n1413 , 
    n1414 , 
    n1415 , 
    n1416 , 
    n1417 , 
    n1418 , 
    n1419 , 
    n1420 , 
    n1421 , 
    n1422 , 
    n1423 , 
    n1424 , 
    n1425 , 
    n1426 , 
    n1427 , 
    n1428 , 
    n1429 , 
    n1430 , 
    n1431 , 
    n1432 , 
    n1433 , 
    n1434 , 
    n1435 , 
    n1436 , 
    n1437 , 
    n1438 , 
    n1439 , 
    n1440 , 
    n1441 , 
    n1442 , 
    n1443 , 
    n1444 , 
    n1445 , 
    n1446 , 
    n1447 , 
    n1448 , 
    n1449 , 
    n1450 , 
    n1451 , 
    n1452 , 
    n1453 , 
    n1454 , 
    n1455 , 
    n1456 , 
    n1457 , 
    n1458 , 
    n1459 , 
    n1460 , 
    n1461 , 
    n1462 , 
    n1463 , 
    n1464 , 
    n1465 , 
    n1466 , 
    n1467 , 
    n1468 , 
    n1469 , 
    n1470 , 
    n1471 , 
    n1472 , 
    n1473 , 
    n1474 , 
    n1475 , 
    n1476 , 
    n1477 , 
    n1478 , 
    n1479 , 
    n1480 , 
    n1481 , 
    n1482 , 
    n1483 , 
    n1484 , 
    n1485 , 
    n1486 , 
    n1487 , 
    n1488 , 
    n1489 , 
    n1490 , 
    n1491 , 
    n1492 , 
    n1493 , 
    n1494 , 
    n1495 , 
    n1496 , 
    n1497 , 
    n1498 , 
    n1499 , 
    n1500 , 
    n1501 , 
    n1502 , 
    n1503 , 
    n1504 , 
    n1505 , 
    n1506 , 
    n1507 , 
    n1508 , 
    n1509 , 
    n1510 , 
    n1511 , 
    n1512 , 
    n1513 , 
    n1514 , 
    n1515 , 
    n1516 , 
    n1517 , 
    n1518 , 
    n1519 , 
    n1520 , 
    n1521 , 
    n1522 , 
    n1523 , 
    n1524 , 
    n1525 , 
    n1526 , 
    n1527 , 
    n1528 , 
    n1529 , 
    n1530 , 
    n1531 , 
    n1532 , 
    n1533 , 
    n1534 , 
    n1535 , 
    n1536 , 
    n1537 , 
    n1538 , 
    n1539 , 
    n1540 , 
    n1541 , 
    n1542 , 
    n1543 , 
    n1544 , 
    n1545 , 
    n1546 , 
    n1547 , 
    n1548 , 
    n1549 , 
    n1550 , 
    n1551 , 
    n1552 , 
    n1553 , 
    n1554 , 
    n1555 , 
    n1556 , 
    n1557 , 
    n1558 , 
    n1559 , 
    n1560 , 
    n1561 , 
    n1562 , 
    n1563 , 
    n1564 , 
    n1565 , 
    n1566 , 
    n1567 , 
    n1568 , 
    n1569 , 
    n1570 , 
    n1571 , 
    n1572 , 
    n1573 , 
    n1574 , 
    n1575 , 
    n1576 , 
    n1577 , 
    n1578 , 
    n1579 , 
    n1580 , 
    n1581 , 
    n1582 , 
    n1583 , 
    n1584 , 
    n1585 , 
    n1586 , 
    n1587 , 
    n1588 , 
    n1589 , 
    n1590 , 
    n1591 , 
    n1592 , 
    n1593 , 
    n1594 , 
    n1595 , 
    n1596 , 
    n1597 , 
    n1598 , 
    n1599 , 
    n1600 , 
    n1601 , 
    n1602 , 
    n1603 , 
    n1604 , 
    n1605 , 
    n1606 , 
    n1607 , 
    n1608 , 
    n1609 , 
    n1610 , 
    n1611 , 
    n1612 , 
    n1613 , 
    n1614 , 
    n1615 , 
    n1616 , 
    n1617 , 
    n1618 , 
    n1619 , 
    n1620 , 
    n1621 , 
    n1622 , 
    n1623 , 
    n1624 , 
    n1625 , 
    n1626 , 
    n1627 , 
    n1628 , 
    n1629 , 
    n1630 , 
    n1631 , 
    n1632 , 
    n1633 , 
    n1634 , 
    n1635 , 
    n1636 , 
    n1637 , 
    n1638 , 
    n1639 , 
    n1640 , 
    n1641 , 
    n1642 , 
    n1643 , 
    n1644 , 
    n1645 , 
    n1646 , 
    n1647 , 
    n1648 , 
    n1649 , 
    n1650 , 
    n1651 , 
    n1652 , 
    n1653 , 
    n1654 , 
    n1655 , 
    n1656 , 
    n1657 , 
    n1658 , 
    n1659 , 
    n1660 , 
    n1661 , 
    n1662 , 
    n1663 , 
    n1664 , 
    n1665 , 
    n1666 , 
    n1667 , 
    n1668 , 
    n1669 , 
    n1670 , 
    n1671 , 
    n1672 , 
    n1673 , 
    n1674 , 
    n1675 , 
    n1676 , 
    n1677 , 
    n1678 , 
    n1679 , 
    n1680 , 
    n1681 , 
    n1682 , 
    n1683 , 
    n1684 , 
    n1685 , 
    n1686 , 
    n1687 , 
    n1688 , 
    n1689 , 
    n1690 , 
    n1691 , 
    n1692 , 
    n1693 , 
    n1694 , 
    n1695 , 
    n1696 , 
    n1697 , 
    n1698 , 
    n1699 , 
    n1700 , 
    n1701 , 
    n1702 , 
    n1703 , 
    n1704 , 
    n1705 , 
    n1706 , 
    n1707 , 
    n1708 , 
    n1709 , 
    n1710 , 
    n1711 , 
    n1712 , 
    n1713 , 
    n1714 , 
    n1715 , 
    n1716 , 
    n1717 , 
    n1718 , 
    n1719 , 
    n1720 , 
    n1721 , 
    n1722 , 
    n1723 , 
    n1724 , 
    n1725 , 
    n1726 , 
    n1727 , 
    n1728 , 
    n1729 , 
    n1730 , 
    n1731 , 
    n1732 , 
    n1733 , 
    n1734 , 
    n1735 , 
    n1736 , 
    n1737 , 
    n1738 , 
    n1739 , 
    n1740 , 
    n1741 , 
    n1742 , 
    n1743 , 
    n1744 , 
    n1745 , 
    n1746 , 
    n1747 , 
    n1748 , 
    n1749 , 
    n1750 , 
    n1751 , 
    n1752 , 
    n1753 , 
    n1754 , 
    n1755 , 
    n1756 , 
    n1757 , 
    n1758 , 
    n1759 , 
    n1760 , 
    n1761 , 
    n1762 , 
    n1763 , 
    n1764 , 
    n1765 , 
    n1766 , 
    n1767 , 
    n1768 , 
    n1769 , 
    n1770 , 
    n1771 , 
    n1772 , 
    n1773 , 
    n1774 , 
    n1775 , 
    n1776 , 
    n1777 , 
    n1778 , 
    n1779 , 
    n1780 , 
    n1781 , 
    n1782 , 
    n1783 , 
    n1784 , 
    n1785 , 
    n1786 , 
    n1787 , 
    n1788 , 
    n1789 , 
    n1790 , 
    n1791 , 
    n1792 , 
    n1793 , 
    n1794 , 
    n1795 , 
    n1796 , 
    n1797 , 
    n1798 , 
    n1799 , 
    n1800 , 
    n1801 , 
    n1802 , 
    n1803 , 
    n1804 , 
    n1805 , 
    n1806 , 
    n1807 , 
    n1808 , 
    n1809 , 
    n1810 , 
    n1811 , 
    n1812 , 
    n1813 , 
    n1814 , 
    n1815 , 
    n1816 , 
    n1817 , 
    n1818 , 
    n1819 , 
    n1820 , 
    n1821 , 
    n1822 , 
    n1823 , 
    n1824 , 
    n1825 , 
    n1826 , 
    n1827 , 
    n1828 , 
    n1829 , 
    n1830 , 
    n1831 , 
    n1832 , 
    n1833 , 
    n1834 , 
    n1835 , 
    n1836 , 
    n1837 , 
    n1838 , 
    n1839 , 
    n1840 , 
    n1841 , 
    n1842 , 
    n1843 , 
    n1844 , 
    n1845 , 
    n1846 , 
    n1847 , 
    n1848 , 
    n1849 , 
    n1850 , 
    n1851 , 
    n1852 , 
    n1853 , 
    n1854 , 
    n1855 , 
    n1856 , 
    n1857 , 
    n1858 , 
    n1859 , 
    n1860 , 
    n1861 , 
    n1862 , 
    n1863 , 
    n1864 , 
    n1865 , 
    n1866 , 
    n1867 , 
    n1868 , 
    n1869 , 
    n1870 , 
    n1871 , 
    n1872 , 
    n1873 , 
    n1874 , 
    n1875 , 
    n1876 , 
    n1877 , 
    n1878 , 
    n1879 , 
    n1880 , 
    n1881 , 
    n1882 , 
    n1883 , 
    n1884 , 
    n1885 , 
    n1886 , 
    n1887 , 
    n1888 , 
    n1889 , 
    n1890 , 
    n1891 , 
    n1892 , 
    n1893 , 
    n1894 , 
    n1895 , 
    n1896 , 
    n1897 , 
    n1898 , 
    n1899 , 
    n1900 , 
    n1901 , 
    n1902 , 
    n1903 , 
    n1904 , 
    n1905 , 
    n1906 , 
    n1907 , 
    n1908 , 
    n1909 , 
    n1910 , 
    n1911 , 
    n1912 , 
    n1913 , 
    n1914 , 
    n1915 , 
    n1916 , 
    n1917 , 
    n1918 , 
    n1919 , 
    n1920 , 
    n1921 , 
    n1922 , 
    n1923 , 
    n1924 , 
    n1925 , 
    n1926 , 
    n1927 , 
    n1928 , 
    n1929 , 
    n1930 , 
    n1931 , 
    n1932 , 
    n1933 , 
    n1934 , 
    n1935 , 
    n1936 , 
    n1937 , 
    n1938 , 
    n1939 , 
    n1940 , 
    n1941 , 
    n1942 , 
    n1943 , 
    n1944 , 
    n1945 , 
    n1946 , 
    n1947 , 
    n1948 , 
    n1949 , 
    n1950 , 
    n1951 , 
    n1952 , 
    n1953 , 
    n1954 , 
    n1955 , 
    n1956 , 
    n1957 , 
    n1958 , 
    n1959 , 
    n1960 , 
    n1961 , 
    n1962 , 
    n1963 , 
    n1964 , 
    n1965 , 
    n1966 , 
    n1967 , 
    n1968 , 
    n1969 , 
    n1970 , 
    n1971 , 
    n1972 , 
    n1973 , 
    n1974 , 
    n1975 , 
    n1976 , 
    n1977 , 
    n1978 , 
    n1979 , 
    n1980 , 
    n1981 , 
    n1982 , 
    n1983 , 
    n1984 , 
    n1985 , 
    n1986 , 
    n1987 , 
    n1988 , 
    n1989 , 
    n1990 , 
    n1991 , 
    n1992 , 
    n1993 , 
    n1994 , 
    n1995 , 
    n1996 , 
    n1997 , 
    n1998 , 
    n1999 , 
    n2000 , 
    n2001 , 
    n2002 , 
    n2003 , 
    n2004 , 
    n2005 , 
    n2006 , 
    n2007 , 
    n2008 , 
    n2009 , 
    n2010 , 
    n2011 , 
    n2012 , 
    n2013 , 
    n2014 , 
    n2015 , 
    n2016 , 
    n2017 , 
    n2018 , 
    n2019 , 
    n2020 , 
    n2021 , 
    n2022 , 
    n2023 , 
    n2024 , 
    n2025 , 
    n2026 , 
    n2027 , 
    n2028 , 
    n2029 , 
    n2030 , 
    n2031 , 
    n2032 , 
    n2033 , 
    n2034 , 
    n2035 , 
    n2036 , 
    n2037 , 
    n2038 , 
    n2039 , 
    n2040 , 
    n2041 , 
    n2042 , 
    n2043 , 
    n2044 , 
    n2045 , 
    n2046 , 
    n2047 , 
    n2048 , 
    n2049 , 
    n2050 , 
    n2051 , 
    n2052 , 
    n2053 , 
    n2054 , 
    n2055 , 
    n2056 , 
    n2057 , 
    n2058 , 
    n2059 , 
    n2060 , 
    n2061 , 
    n2062 , 
    n2063 , 
    n2064 , 
    n2065 , 
    n2066 , 
    n2067 , 
    n2068 , 
    n2069 , 
    n2070 , 
    n2071 , 
    n2072 , 
    n2073 , 
    n2074 , 
    n2075 , 
    n2076 , 
    n2077 , 
    n2078 , 
    n2079 , 
    n2080 , 
    n2081 , 
    n2082 , 
    n2083 , 
    n2084 , 
    n2085 , 
    n2086 , 
    n2087 , 
    n2088 , 
    n2089 , 
    n2090 , 
    n2091 , 
    n2092 , 
    n2093 , 
    n2094 , 
    n2095 , 
    n2096 , 
    n2097 , 
    n2098 , 
    n2099 , 
    n2100 , 
    n2101 , 
    n2102 , 
    n2103 , 
    n2104 , 
    n2105 , 
    n2106 , 
    n2107 , 
    n2108 , 
    n2109 , 
    n2110 , 
    n2111 , 
    n2112 , 
    n2113 , 
    n2114 , 
    n2115 , 
    n2116 , 
    n2117 , 
    n2118 , 
    n2119 , 
    n2120 , 
    n2121 , 
    n2122 , 
    n2123 , 
    n2124 , 
    n2125 , 
    n2126 , 
    n2127 , 
    n2128 , 
    n2129 , 
    n2130 , 
    n2131 , 
    n2132 , 
    n2133 , 
    n2134 , 
    n2135 , 
    n2136 , 
    n2137 , 
    n2138 , 
    n2139 , 
    n2140 , 
    n2141 , 
    n2142 , 
    n2143 , 
    n2144 , 
    n2145 , 
    n2146 , 
    n2147 , 
    n2148 , 
    n2149 , 
    n2150 , 
    n2151 , 
    n2152 , 
    n2153 , 
    n2154 , 
    n2155 , 
    n2156 , 
    n2157 , 
    n2158 , 
    n2159 , 
    n2160 , 
    n2161 , 
    n2162 , 
    n2163 , 
    n2164 , 
    n2165 , 
    n2166 , 
    n2167 , 
    n2168 , 
    n2169 , 
    n2170 , 
    n2171 , 
    n2172 , 
    n2173 , 
    n2174 , 
    n2175 , 
    n2176 , 
    n2177 , 
    n2178 , 
    n2179 , 
    n2180 , 
    n2181 , 
    n2182 , 
    n2183 , 
    n2184 , 
    n2185 , 
    n2186 , 
    n2187 , 
    n2188 , 
    n2189 , 
    n2190 , 
    n2191 , 
    n2192 , 
    n2193 , 
    n2194 , 
    n2195 , 
    n2196 , 
    n2197 , 
    n2198 , 
    n2199 , 
    n2200 , 
    n2201 , 
    n2202 , 
    n2203 , 
    n2204 , 
    n2205 , 
    n2206 , 
    n2207 , 
    n2208 , 
    n2209 , 
    n2210 , 
    n2211 , 
    n2212 , 
    n2213 , 
    n2214 , 
    n2215 , 
    n2216 , 
    n2217 , 
    n2218 , 
    n2219 , 
    n2220 , 
    n2221 , 
    n2222 , 
    n2223 , 
    n2224 , 
    n2225 , 
    n2226 , 
    n2227 , 
    n2228 , 
    n2229 , 
    n2230 , 
    n2231 , 
    n2232 , 
    n2233 , 
    n2234 , 
    n2235 , 
    n2236 , 
    n2237 , 
    n2238 , 
    n2239 , 
    n2240 , 
    n2241 , 
    n2242 , 
    n2243 , 
    n2244 , 
    n2245 , 
    n2246 , 
    n2247 , 
    n2248 , 
    n2249 , 
    n2250 , 
    n2251 , 
    n2252 , 
    n2253 , 
    n2254 , 
    n2255 , 
    n2256 , 
    n2257 , 
    n2258 , 
    n2259 , 
    n2260 , 
    n2261 , 
    n2262 , 
    n2263 , 
    n2264 , 
    n2265 , 
    n2266 , 
    n2267 , 
    n2268 , 
    n2269 , 
    n2270 , 
    n2271 , 
    n2272 , 
    n2273 , 
    n2274 , 
    n2275 , 
    n2276 , 
    n2277 , 
    n2278 , 
    n2279 , 
    n2280 , 
    n2281 , 
    n2282 , 
    n2283 , 
    n2284 , 
    n2285 , 
    n2286 , 
    n2287 , 
    n2288 , 
    n2289 , 
    n2290 , 
    n2291 , 
    n2292 , 
    n2293 , 
    n2294 , 
    n2295 , 
    n2296 , 
    n2297 , 
    n2298 , 
    n2299 , 
    n2300 , 
    n2301 , 
    n2302 , 
    n2303 , 
    n2304 , 
    n2305 , 
    n2306 , 
    n2307 , 
    n2308 , 
    n2309 , 
    n2310 , 
    n2311 , 
    n2312 , 
    n2313 , 
    n2314 , 
    n2315 , 
    n2316 , 
    n2317 , 
    n2318 , 
    n2319 , 
    n2320 , 
    n2321 , 
    n2322 , 
    n2323 , 
    n2324 , 
    n2325 , 
    n2326 , 
    n2327 , 
    n2328 , 
    n2329 , 
    n2330 , 
    n2331 , 
    n2332 , 
    n2333 , 
    n2334 , 
    n2335 , 
    n2336 , 
    n2337 , 
    n2338 , 
    n2339 , 
    n2340 , 
    n2341 , 
    n2342 , 
    n2343 , 
    n2344 , 
    n2345 , 
    n2346 , 
    n2347 , 
    n2348 , 
    n2349 , 
    n2350 , 
    n2351 , 
    n2352 , 
    n2353 , 
    n2354 , 
    n2355 , 
    n2356 , 
    n2357 , 
    n2358 , 
    n2359 , 
    n2360 , 
    n2361 , 
    n2362 , 
    n2363 , 
    n2364 , 
    n2365 , 
    n2366 , 
    n2367 , 
    n2368 , 
    n2369 , 
    n2370 , 
    n2371 , 
    n2372 , 
    n2373 , 
    n2374 , 
    n2375 , 
    n2376 , 
    n2377 , 
    n2378 , 
    n2379 , 
    n2380 , 
    n2381 , 
    n2382 , 
    n2383 , 
    n2384 , 
    n2385 , 
    n2386 , 
    n2387 , 
    n2388 , 
    n2389 , 
    n2390 , 
    n2391 , 
    n2392 , 
    n2393 , 
    n2394 , 
    n2395 , 
    n2396 , 
    n2397 , 
    n2398 , 
    n2399 , 
    n2400 , 
    n2401 , 
    n2402 , 
    n2403 , 
    n2404 , 
    n2405 , 
    n2406 , 
    n2407 , 
    n2408 , 
    n2409 , 
    n2410 , 
    n2411 , 
    n2412 , 
    n2413 , 
    n2414 , 
    n2415 , 
    n2416 , 
    n2417 , 
    n2418 , 
    n2419 , 
    n2420 , 
    n2421 , 
    n2422 , 
    n2423 , 
    n2424 , 
    n2425 , 
    n2426 , 
    n2427 , 
    n2428 , 
    n2429 , 
    n2430 , 
    n2431 , 
    n2432 , 
    n2433 , 
    n2434 , 
    n2435 , 
    n2436 , 
    n2437 , 
    n2438 , 
    n2439 , 
    n2440 , 
    n2441 , 
    n2442 , 
    n2443 , 
    n2444 , 
    n2445 , 
    n2446 , 
    n2447 , 
    n2448 , 
    n2449 , 
    n2450 , 
    n2451 , 
    n2452 , 
    n2453 , 
    n2454 , 
    n2455 , 
    n2456 , 
    n2457 , 
    n2458 , 
    n2459 , 
    n2460 , 
    n2461 , 
    n2462 , 
    n2463 , 
    n2464 , 
    n2465 , 
    n2466 , 
    n2467 , 
    n2468 , 
    n2469 , 
    n2470 , 
    n2471 , 
    n2472 , 
    n2473 , 
    n2474 , 
    n2475 , 
    n2476 , 
    n2477 , 
    n2478 , 
    n2479 , 
    n2480 , 
    n2481 , 
    n2482 , 
    n2483 , 
    n2484 , 
    n2485 , 
    n2486 , 
    n2487 , 
    n2488 , 
    n2489 , 
    n2490 , 
    n2491 , 
    n2492 , 
    n2493 , 
    n2494 , 
    n2495 , 
    n2496 , 
    n2497 , 
    n2498 , 
    n2499 , 
    n2500 , 
    n2501 , 
    n2502 , 
    n2503 , 
    n2504 , 
    n2505 , 
    n2506 , 
    n2507 , 
    n2508 , 
    n2509 , 
    n2510 , 
    n2511 , 
    n2512 , 
    n2513 , 
    n2514 , 
    n2515 , 
    n2516 , 
    n2517 , 
    n2518 , 
    n2519 , 
    n2520 , 
    n2521 , 
    n2522 , 
    n2523 , 
    n2524 , 
    n2525 , 
    n2526 , 
    n2527 , 
    n2528 , 
    n2529 , 
    n2530 , 
    n2531 , 
    n2532 , 
    n2533 , 
    n2534 , 
    n2535 , 
    n2536 , 
    n2537 , 
    n2538 , 
    n2539 , 
    n2540 , 
    n2541 , 
    n2542 , 
    n2543 , 
    n2544 , 
    n2545 , 
    n2546 , 
    n2547 , 
    n2548 , 
    n2549 , 
    n2550 , 
    n2551 , 
    n2552 , 
    n2553 , 
    n2554 , 
    n2555 , 
    n2556 , 
    n2557 , 
    n2558 , 
    n2559 , 
    n2560 , 
    n2561 , 
    n2562 , 
    n2563 , 
    n2564 , 
    n2565 , 
    n2566 , 
    n2567 , 
    n2568 , 
    n2569 , 
    n2570 , 
    n2571 , 
    n2572 , 
    n2573 , 
    n2574 , 
    n2575 , 
    n2576 , 
    n2577 , 
    n2578 , 
    n2579 , 
    n2580 , 
    n2581 , 
    n2582 , 
    n2583 , 
    n2584 , 
    n2585 , 
    n2586 , 
    n2587 , 
    n2588 , 
    n2589 , 
    n2590 , 
    n2591 , 
    n2592 , 
    n2593 , 
    n2594 , 
    n2595 , 
    n2596 , 
    n2597 , 
    n2598 , 
    n2599 , 
    n2600 , 
    n2601 , 
    n2602 , 
    n2603 , 
    n2604 , 
    n2605 , 
    n2606 , 
    n2607 , 
    n2608 , 
    n2609 , 
    n2610 , 
    n2611 , 
    n2612 , 
    n2613 , 
    n2614 , 
    n2615 , 
    n2616 , 
    n2617 , 
    n2618 , 
    n2619 , 
    n2620 , 
    n2621 , 
    n2622 , 
    n2623 , 
    n2624 , 
    n2625 , 
    n2626 , 
    n2627 , 
    n2628 , 
    n2629 , 
    n2630 , 
    n2631 , 
    n2632 , 
    n2633 , 
    n2634 , 
    n2635 , 
    n2636 , 
    n2637 , 
    n2638 , 
    n2639 , 
    n2640 , 
    n2641 , 
    n2642 , 
    n2643 , 
    n2644 , 
    n2645 , 
    n2646 , 
    n2647 , 
    n2648 , 
    n2649 , 
    n2650 , 
    n2651 , 
    n2652 , 
    n2653 , 
    n2654 , 
    n2655 , 
    n2656 , 
    n2657 , 
    n2658 , 
    n2659 , 
    n2660 , 
    n2661 , 
    n2662 , 
    n2663 , 
    n2664 , 
    n2665 , 
    n2666 , 
    n2667 , 
    n2668 , 
    n2669 , 
    n2670 , 
    n2671 , 
    n2672 , 
    n2673 , 
    n2674 , 
    n2675 , 
    n2676 , 
    n2677 , 
    n2678 , 
    n2679 , 
    n2680 , 
    n2681 , 
    n2682 , 
    n2683 , 
    n2684 , 
    n2685 , 
    n2686 , 
    n2687 , 
    n2688 , 
    n2689 , 
    n2690 , 
    n2691 , 
    n2692 , 
    n2693 , 
    n2694 , 
    n2695 , 
    n2696 , 
    n2697 , 
    n2698 , 
    n2699 , 
    n2700 , 
    n2701 , 
    n2702 , 
    n2703 , 
    n2704 , 
    n2705 , 
    n2706 , 
    n2707 , 
    n2708 , 
    n2709 , 
    n2710 , 
    n2711 , 
    n2712 , 
    n2713 , 
    n2714 , 
    n2715 , 
    n2716 , 
    n2717 , 
    n2718 , 
    n2719 , 
    n2720 , 
    n2721 , 
    n2722 , 
    n2723 , 
    n2724 , 
    n2725 , 
    n2726 , 
    n2727 , 
    n2728 , 
    n2729 , 
    n2730 , 
    n2731 , 
    n2732 , 
    n2733 , 
    n2734 , 
    n2735 , 
    n2736 , 
    n2737 , 
    n2738 , 
    n2739 , 
    n2740 , 
    n2741 , 
    n2742 , 
    n2743 , 
    n2744 , 
    n2745 , 
    n2746 , 
    n2747 , 
    n2748 , 
    n2749 , 
    n2750 , 
    n2751 , 
    n2752 , 
    n2753 , 
    n2754 , 
    n2755 , 
    n2756 , 
    n2757 , 
    n2758 , 
    n2759 , 
    n2760 , 
    n2761 , 
    n2762 , 
    n2763 , 
    n2764 , 
    n2765 , 
    n2766 , 
    n2767 , 
    n2768 , 
    n2769 , 
    n2770 , 
    n2771 , 
    n2772 , 
    n2773 , 
    n2774 , 
    n2775 , 
    n2776 , 
    n2777 , 
    n2778 , 
    n2779 , 
    n2780 , 
    n2781 , 
    n2782 , 
    n2783 , 
    n2784 , 
    n2785 , 
    n2786 , 
    n2787 , 
    n2788 , 
    n2789 , 
    n2790 , 
    n2791 , 
    n2792 , 
    n2793 , 
    n2794 , 
    n2795 , 
    n2796 , 
    n2797 , 
    n2798 , 
    n2799 , 
    n2800 , 
    n2801 , 
    n2802 , 
    n2803 , 
    n2804 , 
    n2805 , 
    n2806 , 
    n2807 , 
    n2808 , 
    n2809 , 
    n2810 , 
    n2811 , 
    n2812 , 
    n2813 , 
    n2814 , 
    n2815 , 
    n2816 , 
    n2817 , 
    n2818 , 
    n2819 , 
    n2820 , 
    n2821 , 
    n2822 , 
    n2823 , 
    n2824 , 
    n2825 , 
    n2826 , 
    n2827 , 
    n2828 , 
    n2829 , 
    n2830 , 
    n2831 , 
    n2832 , 
    n2833 , 
    n2834 , 
    n2835 , 
    n2836 , 
    n2837 , 
    n2838 , 
    n2839 , 
    n2840 , 
    n2841 , 
    n2842 , 
    n2843 , 
    n2844 , 
    n2845 , 
    n2846 , 
    n2847 , 
    n2848 , 
    n2849 , 
    n2850 , 
    n2851 , 
    n2852 , 
    n2853 , 
    n2854 , 
    n2855 , 
    n2856 , 
    n2857 , 
    n2858 , 
    n2859 , 
    n2860 , 
    n2861 , 
    n2862 , 
    n2863 , 
    n2864 , 
    n2865 , 
    n2866 , 
    n2867 , 
    n2868 , 
    n2869 , 
    n2870 , 
    n2871 , 
    n2872 , 
    n2873 , 
    n2874 , 
    n2875 , 
    n2876 , 
    n2877 , 
    n2878 , 
    n2879 , 
    n2880 , 
    n2881 , 
    n2882 , 
    n2883 , 
    n2884 , 
    n2885 , 
    n2886 , 
    n2887 , 
    n2888 , 
    n2889 , 
    n2890 , 
    n2891 , 
    n2892 , 
    n2893 , 
    n2894 , 
    n2895 , 
    n2896 , 
    n2897 , 
    n2898 , 
    n2899 , 
    n2900 , 
    n2901 , 
    n2902 , 
    n2903 , 
    n2904 , 
    n2905 , 
    n2906 , 
    n2907 , 
    n2908 , 
    n2909 , 
    n2910 , 
    n2911 , 
    n2912 , 
    n2913 , 
    n2914 , 
    n2915 , 
    n2916 , 
    n2917 , 
    n2918 , 
    n2919 , 
    n2920 , 
    n2921 , 
    n2922 , 
    n2923 , 
    n2924 , 
    n2925 , 
    n2926 , 
    n2927 , 
    n2928 , 
    n2929 , 
    n2930 , 
    n2931 , 
    n2932 , 
    n2933 , 
    n2934 , 
    n2935 , 
    n2936 , 
    n2937 , 
    n2938 , 
    n2939 , 
    n2940 , 
    n2941 , 
    n2942 , 
    n2943 , 
    n2944 , 
    n2945 , 
    n2946 , 
    n2947 , 
    n2948 , 
    n2949 , 
    n2950 , 
    n2951 , 
    n2952 , 
    n2953 , 
    n2954 , 
    n2955 , 
    n2956 , 
    n2957 , 
    n2958 , 
    n2959 , 
    n2960 , 
    n2961 , 
    n2962 , 
    n2963 , 
    n2964 , 
    n2965 , 
    n2966 , 
    n2967 , 
    n2968 , 
    n2969 , 
    n2970 , 
    n2971 , 
    n2972 , 
    n2973 , 
    n2974 , 
    n2975 , 
    n2976 , 
    n2977 , 
    n2978 , 
    n2979 , 
    n2980 , 
    n2981 , 
    n2982 , 
    n2983 , 
    n2984 , 
    n2985 , 
    n2986 , 
    n2987 , 
    n2988 , 
    n2989 , 
    n2990 , 
    n2991 , 
    n2992 , 
    n2993 , 
    n2994 , 
    n2995 , 
    n2996 , 
    n2997 , 
    n2998 , 
    n2999 , 
    n3000 , 
    n3001 , 
    n3002 , 
    n3003 , 
    n3004 , 
    n3005 , 
    n3006 , 
    n3007 , 
    n3008 , 
    n3009 , 
    n3010 , 
    n3011 , 
    n3012 , 
    n3013 , 
    n3014 , 
    n3015 , 
    n3016 , 
    n3017 , 
    n3018 , 
    n3019 , 
    n3020 , 
    n3021 , 
    n3022 , 
    n3023 , 
    n3024 , 
    n3025 , 
    n3026 , 
    n3027 , 
    n3028 , 
    n3029 , 
    n3030 , 
    n3031 , 
    n3032 , 
    n3033 , 
    n3034 , 
    n3035 , 
    n3036 , 
    n3037 , 
    n3038 , 
    n3039 , 
    n3040 , 
    n3041 , 
    n3042 , 
    n3043 , 
    n3044 , 
    n3045 , 
    n3046 , 
    n3047 , 
    n3048 , 
    n3049 , 
    n3050 , 
    n3051 , 
    n3052 , 
    n3053 , 
    n3054 , 
    n3055 , 
    n3056 , 
    n3057 , 
    n3058 , 
    n3059 , 
    n3060 , 
    n3061 , 
    n3062 , 
    n3063 , 
    n3064 , 
    n3065 , 
    n3066 , 
    n3067 , 
    n3068 , 
    n3069 , 
    n3070 , 
    n3071 , 
    n3072 , 
    n3073 , 
    n3074 , 
    n3075 , 
    n3076 , 
    n3077 , 
    n3078 , 
    n3079 , 
    n3080 , 
    n3081 , 
    n3082 , 
    n3083 , 
    n3084 , 
    n3085 , 
    n3086 , 
    n3087 , 
    n3088 , 
    n3089 , 
    n3090 , 
    n3091 , 
    n3092 , 
    n3093 , 
    n3094 , 
    n3095 , 
    n3096 , 
    n3097 , 
    n3098 , 
    n3099 , 
    n3100 , 
    n3101 , 
    n3102 , 
    n3103 , 
    n3104 , 
    n3105 , 
    n3106 , 
    n3107 , 
    n3108 , 
    n3109 , 
    n3110 , 
    n3111 , 
    n3112 , 
    n3113 , 
    n3114 , 
    n3115 , 
    n3116 , 
    n3117 , 
    n3118 , 
    n3119 , 
    n3120 , 
    n3121 , 
    n3122 , 
    n3123 );
input  n0 , 
    n1 , 
    n2 , 
    n3 , 
    n4 , 
    n5 , 
    n6 , 
    n7 , 
    n8 , 
    n9 , 
    n10 , 
    n11 , 
    n12 , 
    n13 , 
    n14 , 
    n15 , 
    n16 , 
    n17 , 
    n18 , 
    n19 , 
    n20 , 
    n21 , 
    n22 , 
    n23 , 
    n24 , 
    n25 , 
    n26 , 
    n27 , 
    n28 , 
    n29 , 
    n30 , 
    n31 , 
    n32 , 
    n33 , 
    n34 , 
    n35 , 
    n36 , 
    n37 , 
    n38 , 
    n39 , 
    n40 , 
    n41 , 
    n42 , 
    n43 , 
    n44 , 
    n45 , 
    n46 , 
    n47 , 
    n48 , 
    n49 , 
    n50 , 
    n51 , 
    n52 , 
    n53 , 
    n54 , 
    n55 , 
    n56 , 
    n57 , 
    n58 , 
    n59 , 
    n60 , 
    n61 , 
    n62 , 
    n63 , 
    n64 , 
    n65 , 
    n66 , 
    n67 , 
    n68 , 
    n69 , 
    n70 , 
    n71 , 
    n72 , 
    n73 , 
    n74 , 
    n75 , 
    n76 , 
    n77 , 
    n78 , 
    n79 , 
    n80 , 
    n81 , 
    n82 , 
    n83 , 
    n84 , 
    n85 , 
    n86 , 
    n87 , 
    n88 , 
    n89 , 
    n90 , 
    n91 , 
    n92 , 
    n93 , 
    n94 , 
    n95 , 
    n96 , 
    n97 , 
    n98 , 
    n99 , 
    n100 , 
    n101 , 
    n102 , 
    n103 , 
    n104 , 
    n105 , 
    n106 , 
    n107 , 
    n108 , 
    n109 , 
    n110 , 
    n111 , 
    n112 , 
    n113 , 
    n114 , 
    n115 , 
    n116 , 
    n117 , 
    n118 , 
    n119 , 
    n120 , 
    n121 , 
    n122 , 
    n123 , 
    n124 , 
    n125 , 
    n126 , 
    n127 , 
    n128 , 
    n129 , 
    n130 , 
    n131 , 
    n132 , 
    n133 , 
    n134 , 
    n135 , 
    n136 , 
    n137 , 
    n138 , 
    n139 , 
    n140 , 
    n141 , 
    n142 , 
    n143 , 
    n144 , 
    n145 , 
    n146 , 
    n147 , 
    n148 , 
    n149 , 
    n150 , 
    n151 , 
    n152 , 
    n153 , 
    n154 , 
    n155 , 
    n156 , 
    n157 , 
    n158 , 
    n159 , 
    n160 , 
    n161 , 
    n162 , 
    n163 , 
    n164 , 
    n165 , 
    n166 , 
    n167 , 
    n168 , 
    n169 , 
    n170 , 
    n171 , 
    n172 , 
    n173 , 
    n174 , 
    n175 , 
    n176 , 
    n177 , 
    n178 , 
    n179 , 
    n180 , 
    n181 , 
    n182 , 
    n183 , 
    n184 , 
    n185 , 
    n186 , 
    n187 , 
    n188 , 
    n189 , 
    n190 , 
    n191 , 
    n192 , 
    n193 , 
    n194 , 
    n195 , 
    n196 , 
    n197 , 
    n198 , 
    n199 , 
    n200 , 
    n201 , 
    n202 , 
    n203 , 
    n204 , 
    n205 , 
    n206 , 
    n207 , 
    n208 , 
    n209 , 
    n210 , 
    n211 , 
    n212 , 
    n213 , 
    n214 , 
    n215 , 
    n216 , 
    n217 , 
    n218 , 
    n219 , 
    n220 , 
    n221 , 
    n222 , 
    n223 , 
    n224 , 
    n225 , 
    n226 , 
    n227 , 
    n228 , 
    n229 , 
    n230 , 
    n231 , 
    n232 , 
    n233 , 
    n234 , 
    n235 , 
    n236 , 
    n237 , 
    n238 , 
    n239 , 
    n240 , 
    n241 , 
    n242 , 
    n243 , 
    n244 , 
    n245 , 
    n246 , 
    n247 , 
    n248 , 
    n249 , 
    n250 , 
    n251 , 
    n252 , 
    n253 , 
    n254 , 
    n255 , 
    n256 , 
    n257 , 
    n258 , 
    n259 , 
    n260 , 
    n261 , 
    n262 , 
    n263 , 
    n264 , 
    n265 , 
    n266 , 
    n267 , 
    n268 , 
    n269 , 
    n270 , 
    n271 , 
    n272 , 
    n273 , 
    n274 , 
    n275 , 
    n276 , 
    n277 , 
    n278 , 
    n279 , 
    n280 , 
    n281 , 
    n282 , 
    n283 , 
    n284 , 
    n285 , 
    n286 , 
    n287 , 
    n288 , 
    n289 , 
    n290 , 
    n291 , 
    n292 , 
    n293 , 
    n294 , 
    n295 , 
    n296 , 
    n297 , 
    n298 , 
    n299 , 
    n300 , 
    n301 , 
    n302 , 
    n303 , 
    n304 , 
    n305 , 
    n306 , 
    n307 , 
    n308 , 
    n309 , 
    n310 , 
    n311 , 
    n312 , 
    n313 , 
    n314 , 
    n315 , 
    n316 , 
    n317 , 
    n318 , 
    n319 , 
    n320 , 
    n321 , 
    n322 , 
    n323 , 
    n324 , 
    n325 , 
    n326 , 
    n327 , 
    n328 , 
    n329 , 
    n330 , 
    n331 , 
    n332 , 
    n333 , 
    n334 , 
    n335 , 
    n336 , 
    n337 , 
    n338 , 
    n339 , 
    n340 , 
    n341 , 
    n342 , 
    n343 , 
    n344 , 
    n345 , 
    n346 , 
    n347 , 
    n348 , 
    n349 , 
    n350 , 
    n351 , 
    n352 , 
    n353 , 
    n354 , 
    n355 , 
    n356 , 
    n357 , 
    n358 , 
    n359 , 
    n360 , 
    n361 , 
    n362 , 
    n363 , 
    n364 , 
    n365 , 
    n366 , 
    n367 , 
    n368 , 
    n369 , 
    n370 , 
    n371 , 
    n372 , 
    n373 , 
    n374 , 
    n375 , 
    n376 , 
    n377 , 
    n378 , 
    n379 , 
    n380 , 
    n381 , 
    n382 , 
    n383 , 
    n384 , 
    n385 , 
    n386 , 
    n387 , 
    n388 , 
    n389 , 
    n390 , 
    n391 , 
    n392 , 
    n393 , 
    n394 , 
    n395 , 
    n396 , 
    n397 , 
    n398 , 
    n399 , 
    n400 , 
    n401 , 
    n402 , 
    n403 , 
    n404 , 
    n405 , 
    n406 , 
    n407 , 
    n408 , 
    n409 , 
    n410 , 
    n411 , 
    n412 , 
    n413 , 
    n414 , 
    n415 , 
    n416 , 
    n417 , 
    n418 , 
    n419 , 
    n420 , 
    n421 , 
    n422 , 
    n423 , 
    n424 , 
    n425 , 
    n426 , 
    n427 , 
    n428 , 
    n429 , 
    n430 , 
    n431 , 
    n432 , 
    n433 , 
    n434 , 
    n435 , 
    n436 , 
    n437 , 
    n438 , 
    n439 , 
    n440 , 
    n441 , 
    n442 , 
    n443 , 
    n444 , 
    n445 , 
    n446 , 
    n447 , 
    n448 , 
    n449 , 
    n450 , 
    n451 , 
    n452 , 
    n453 , 
    n454 , 
    n455 , 
    n456 , 
    n457 , 
    n458 , 
    n459 , 
    n460 , 
    n461 , 
    n462 , 
    n463 , 
    n464 , 
    n465 , 
    n466 , 
    n467 , 
    n468 , 
    n469 , 
    n470 , 
    n471 , 
    n472 , 
    n473 , 
    n474 , 
    n475 , 
    n476 , 
    n477 , 
    n478 , 
    n479 , 
    n480 , 
    n481 , 
    n482 , 
    n483 , 
    n484 , 
    n485 , 
    n486 , 
    n487 , 
    n488 , 
    n489 , 
    n490 , 
    n491 , 
    n492 , 
    n493 , 
    n494 , 
    n495 , 
    n496 , 
    n497 , 
    n498 , 
    n499 , 
    n500 , 
    n501 , 
    n502 , 
    n503 , 
    n504 , 
    n505 , 
    n506 , 
    n507 , 
    n508 , 
    n509 , 
    n510 , 
    n511 , 
    n512 , 
    n513 , 
    n514 , 
    n515 , 
    n516 , 
    n517 , 
    n518 , 
    n519 , 
    n520 , 
    n521 , 
    n522 , 
    n523 , 
    n524 , 
    n525 , 
    n526 , 
    n527 , 
    n528 , 
    n529 , 
    n530 , 
    n531 , 
    n532 , 
    n533 , 
    n534 , 
    n535 , 
    n536 , 
    n537 , 
    n538 , 
    n539 , 
    n540 , 
    n541 , 
    n542 , 
    n543 , 
    n544 , 
    n545 , 
    n546 , 
    n547 , 
    n548 , 
    n549 , 
    n550 , 
    n551 , 
    n552 , 
    n553 , 
    n554 , 
    n555 , 
    n556 , 
    n557 , 
    n558 , 
    n559 , 
    n560 , 
    n561 , 
    n562 , 
    n563 , 
    n564 , 
    n565 , 
    n566 , 
    n567 , 
    n568 , 
    n569 , 
    n570 , 
    n571 , 
    n572 , 
    n573 , 
    n574 , 
    n575 , 
    n576 , 
    n577 , 
    n578 , 
    n579 , 
    n580 , 
    n581 , 
    n582 , 
    n583 , 
    n584 , 
    n585 , 
    n586 , 
    n587 , 
    n588 , 
    n589 , 
    n590 , 
    n591 , 
    n592 , 
    n593 , 
    n594 , 
    n595 , 
    n596 , 
    n597 , 
    n598 , 
    n599 , 
    n600 , 
    n601 , 
    n602 , 
    n603 , 
    n604 , 
    n605 , 
    n606 , 
    n607 , 
    n608 , 
    n609 , 
    n610 , 
    n611 , 
    n612 , 
    n613 , 
    n614 , 
    n615 , 
    n616 , 
    n617 , 
    n618 , 
    n619 , 
    n620 , 
    n621 , 
    n622 , 
    n623 , 
    n624 , 
    n625 , 
    n626 , 
    n627 , 
    n628 , 
    n629 , 
    n630 , 
    n631 , 
    n632 , 
    n633 , 
    n634 , 
    n635 , 
    n636 , 
    n637 , 
    n638 , 
    n639 , 
    n640 , 
    n641 , 
    n642 , 
    n643 , 
    n644 , 
    n645 , 
    n646 , 
    n647 , 
    n648 , 
    n649 ;
output 
    n650 , 
    n651 , 
    n652 , 
    n653 , 
    n654 , 
    n655 , 
    n656 , 
    n657 , 
    n658 , 
    n659 , 
    n660 , 
    n661 , 
    n662 , 
    n663 , 
    n664 , 
    n665 , 
    n666 , 
    n667 , 
    n668 , 
    n669 , 
    n670 , 
    n671 , 
    n672 , 
    n673 , 
    n674 , 
    n675 , 
    n676 , 
    n677 , 
    n678 , 
    n679 , 
    n680 , 
    n681 , 
    n682 , 
    n683 , 
    n684 , 
    n685 , 
    n686 , 
    n687 , 
    n688 , 
    n689 , 
    n690 , 
    n691 , 
    n692 , 
    n693 , 
    n694 , 
    n695 , 
    n696 , 
    n697 , 
    n698 , 
    n699 , 
    n700 , 
    n701 , 
    n702 , 
    n703 , 
    n704 , 
    n705 , 
    n706 , 
    n707 , 
    n708 , 
    n709 , 
    n710 , 
    n711 , 
    n712 , 
    n713 , 
    n714 , 
    n715 , 
    n716 , 
    n717 , 
    n718 , 
    n719 , 
    n720 , 
    n721 , 
    n722 , 
    n723 , 
    n724 , 
    n725 , 
    n726 , 
    n727 , 
    n728 , 
    n729 , 
    n730 , 
    n731 , 
    n732 , 
    n733 , 
    n734 , 
    n735 , 
    n736 , 
    n737 , 
    n738 , 
    n739 , 
    n740 , 
    n741 , 
    n742 , 
    n743 , 
    n744 , 
    n745 , 
    n746 , 
    n747 , 
    n748 , 
    n749 , 
    n750 , 
    n751 , 
    n752 , 
    n753 , 
    n754 , 
    n755 , 
    n756 , 
    n757 , 
    n758 , 
    n759 , 
    n760 , 
    n761 , 
    n762 , 
    n763 , 
    n764 , 
    n765 , 
    n766 , 
    n767 , 
    n768 , 
    n769 , 
    n770 , 
    n771 , 
    n772 , 
    n773 , 
    n774 , 
    n775 , 
    n776 , 
    n777 , 
    n778 , 
    n779 , 
    n780 , 
    n781 , 
    n782 , 
    n783 , 
    n784 , 
    n785 , 
    n786 , 
    n787 , 
    n788 , 
    n789 , 
    n790 , 
    n791 , 
    n792 , 
    n793 , 
    n794 , 
    n795 , 
    n796 , 
    n797 , 
    n798 , 
    n799 , 
    n800 , 
    n801 , 
    n802 , 
    n803 , 
    n804 , 
    n805 , 
    n806 , 
    n807 , 
    n808 , 
    n809 , 
    n810 , 
    n811 , 
    n812 , 
    n813 , 
    n814 , 
    n815 , 
    n816 , 
    n817 , 
    n818 , 
    n819 , 
    n820 , 
    n821 , 
    n822 , 
    n823 , 
    n824 , 
    n825 , 
    n826 , 
    n827 , 
    n828 , 
    n829 , 
    n830 , 
    n831 , 
    n832 , 
    n833 , 
    n834 , 
    n835 , 
    n836 , 
    n837 , 
    n838 , 
    n839 , 
    n840 , 
    n841 , 
    n842 , 
    n843 , 
    n844 , 
    n845 , 
    n846 , 
    n847 , 
    n848 , 
    n849 , 
    n850 , 
    n851 , 
    n852 , 
    n853 , 
    n854 , 
    n855 , 
    n856 , 
    n857 , 
    n858 , 
    n859 , 
    n860 , 
    n861 , 
    n862 , 
    n863 , 
    n864 , 
    n865 , 
    n866 , 
    n867 , 
    n868 , 
    n869 , 
    n870 , 
    n871 , 
    n872 , 
    n873 , 
    n874 , 
    n875 , 
    n876 , 
    n877 , 
    n878 , 
    n879 , 
    n880 , 
    n881 , 
    n882 , 
    n883 , 
    n884 , 
    n885 , 
    n886 , 
    n887 , 
    n888 , 
    n889 , 
    n890 , 
    n891 , 
    n892 , 
    n893 , 
    n894 , 
    n895 , 
    n896 , 
    n897 , 
    n898 , 
    n899 , 
    n900 , 
    n901 , 
    n902 , 
    n903 , 
    n904 , 
    n905 , 
    n906 , 
    n907 , 
    n908 , 
    n909 , 
    n910 , 
    n911 , 
    n912 , 
    n913 , 
    n914 , 
    n915 , 
    n916 , 
    n917 , 
    n918 , 
    n919 , 
    n920 , 
    n921 , 
    n922 , 
    n923 , 
    n924 , 
    n925 , 
    n926 , 
    n927 , 
    n928 , 
    n929 , 
    n930 , 
    n931 , 
    n932 , 
    n933 , 
    n934 , 
    n935 , 
    n936 , 
    n937 , 
    n938 , 
    n939 , 
    n940 , 
    n941 , 
    n942 , 
    n943 , 
    n944 , 
    n945 , 
    n946 , 
    n947 , 
    n948 , 
    n949 , 
    n950 , 
    n951 , 
    n952 , 
    n953 , 
    n954 , 
    n955 , 
    n956 , 
    n957 , 
    n958 , 
    n959 , 
    n960 , 
    n961 , 
    n962 , 
    n963 , 
    n964 , 
    n965 , 
    n966 , 
    n967 , 
    n968 , 
    n969 , 
    n970 , 
    n971 , 
    n972 , 
    n973 , 
    n974 , 
    n975 , 
    n976 , 
    n977 , 
    n978 , 
    n979 , 
    n980 , 
    n981 , 
    n982 , 
    n983 , 
    n984 , 
    n985 , 
    n986 , 
    n987 , 
    n988 , 
    n989 , 
    n990 , 
    n991 , 
    n992 , 
    n993 , 
    n994 , 
    n995 , 
    n996 , 
    n997 , 
    n998 , 
    n999 , 
    n1000 , 
    n1001 , 
    n1002 , 
    n1003 , 
    n1004 , 
    n1005 , 
    n1006 , 
    n1007 , 
    n1008 , 
    n1009 , 
    n1010 , 
    n1011 , 
    n1012 , 
    n1013 , 
    n1014 , 
    n1015 , 
    n1016 , 
    n1017 , 
    n1018 , 
    n1019 , 
    n1020 , 
    n1021 , 
    n1022 , 
    n1023 , 
    n1024 , 
    n1025 , 
    n1026 , 
    n1027 , 
    n1028 , 
    n1029 , 
    n1030 , 
    n1031 , 
    n1032 , 
    n1033 , 
    n1034 , 
    n1035 , 
    n1036 , 
    n1037 , 
    n1038 , 
    n1039 , 
    n1040 , 
    n1041 , 
    n1042 , 
    n1043 , 
    n1044 , 
    n1045 , 
    n1046 , 
    n1047 , 
    n1048 , 
    n1049 , 
    n1050 , 
    n1051 , 
    n1052 , 
    n1053 , 
    n1054 , 
    n1055 , 
    n1056 , 
    n1057 , 
    n1058 , 
    n1059 , 
    n1060 , 
    n1061 , 
    n1062 , 
    n1063 , 
    n1064 , 
    n1065 , 
    n1066 , 
    n1067 , 
    n1068 , 
    n1069 , 
    n1070 , 
    n1071 , 
    n1072 , 
    n1073 , 
    n1074 , 
    n1075 , 
    n1076 , 
    n1077 , 
    n1078 , 
    n1079 , 
    n1080 , 
    n1081 , 
    n1082 , 
    n1083 , 
    n1084 , 
    n1085 , 
    n1086 , 
    n1087 , 
    n1088 , 
    n1089 , 
    n1090 , 
    n1091 , 
    n1092 , 
    n1093 , 
    n1094 , 
    n1095 , 
    n1096 , 
    n1097 , 
    n1098 , 
    n1099 , 
    n1100 , 
    n1101 , 
    n1102 , 
    n1103 , 
    n1104 , 
    n1105 , 
    n1106 , 
    n1107 , 
    n1108 , 
    n1109 , 
    n1110 , 
    n1111 , 
    n1112 , 
    n1113 , 
    n1114 , 
    n1115 , 
    n1116 , 
    n1117 , 
    n1118 , 
    n1119 , 
    n1120 , 
    n1121 , 
    n1122 , 
    n1123 , 
    n1124 , 
    n1125 , 
    n1126 , 
    n1127 , 
    n1128 , 
    n1129 , 
    n1130 , 
    n1131 , 
    n1132 , 
    n1133 , 
    n1134 , 
    n1135 , 
    n1136 , 
    n1137 , 
    n1138 , 
    n1139 , 
    n1140 , 
    n1141 , 
    n1142 , 
    n1143 , 
    n1144 , 
    n1145 , 
    n1146 , 
    n1147 , 
    n1148 , 
    n1149 , 
    n1150 , 
    n1151 , 
    n1152 , 
    n1153 , 
    n1154 , 
    n1155 , 
    n1156 , 
    n1157 , 
    n1158 , 
    n1159 , 
    n1160 , 
    n1161 , 
    n1162 , 
    n1163 , 
    n1164 , 
    n1165 , 
    n1166 , 
    n1167 , 
    n1168 , 
    n1169 , 
    n1170 , 
    n1171 , 
    n1172 , 
    n1173 , 
    n1174 , 
    n1175 , 
    n1176 , 
    n1177 , 
    n1178 , 
    n1179 , 
    n1180 , 
    n1181 , 
    n1182 , 
    n1183 , 
    n1184 , 
    n1185 , 
    n1186 , 
    n1187 , 
    n1188 , 
    n1189 , 
    n1190 , 
    n1191 , 
    n1192 , 
    n1193 , 
    n1194 , 
    n1195 , 
    n1196 , 
    n1197 , 
    n1198 , 
    n1199 , 
    n1200 , 
    n1201 , 
    n1202 , 
    n1203 , 
    n1204 , 
    n1205 , 
    n1206 , 
    n1207 , 
    n1208 , 
    n1209 , 
    n1210 , 
    n1211 , 
    n1212 , 
    n1213 , 
    n1214 , 
    n1215 , 
    n1216 , 
    n1217 , 
    n1218 , 
    n1219 , 
    n1220 , 
    n1221 , 
    n1222 , 
    n1223 , 
    n1224 , 
    n1225 , 
    n1226 , 
    n1227 , 
    n1228 , 
    n1229 , 
    n1230 , 
    n1231 , 
    n1232 , 
    n1233 , 
    n1234 , 
    n1235 , 
    n1236 , 
    n1237 , 
    n1238 , 
    n1239 , 
    n1240 , 
    n1241 , 
    n1242 , 
    n1243 , 
    n1244 , 
    n1245 , 
    n1246 , 
    n1247 , 
    n1248 , 
    n1249 , 
    n1250 , 
    n1251 , 
    n1252 , 
    n1253 , 
    n1254 , 
    n1255 , 
    n1256 , 
    n1257 , 
    n1258 , 
    n1259 , 
    n1260 , 
    n1261 , 
    n1262 , 
    n1263 , 
    n1264 , 
    n1265 , 
    n1266 , 
    n1267 , 
    n1268 , 
    n1269 , 
    n1270 , 
    n1271 , 
    n1272 , 
    n1273 , 
    n1274 , 
    n1275 , 
    n1276 , 
    n1277 , 
    n1278 , 
    n1279 , 
    n1280 , 
    n1281 , 
    n1282 , 
    n1283 , 
    n1284 , 
    n1285 , 
    n1286 , 
    n1287 , 
    n1288 , 
    n1289 , 
    n1290 , 
    n1291 , 
    n1292 , 
    n1293 , 
    n1294 , 
    n1295 , 
    n1296 , 
    n1297 , 
    n1298 , 
    n1299 , 
    n1300 , 
    n1301 , 
    n1302 , 
    n1303 , 
    n1304 , 
    n1305 , 
    n1306 , 
    n1307 , 
    n1308 , 
    n1309 , 
    n1310 , 
    n1311 , 
    n1312 , 
    n1313 , 
    n1314 , 
    n1315 , 
    n1316 , 
    n1317 , 
    n1318 , 
    n1319 , 
    n1320 , 
    n1321 , 
    n1322 , 
    n1323 , 
    n1324 , 
    n1325 , 
    n1326 , 
    n1327 , 
    n1328 , 
    n1329 , 
    n1330 , 
    n1331 , 
    n1332 , 
    n1333 , 
    n1334 , 
    n1335 , 
    n1336 , 
    n1337 , 
    n1338 , 
    n1339 , 
    n1340 , 
    n1341 , 
    n1342 , 
    n1343 , 
    n1344 , 
    n1345 , 
    n1346 , 
    n1347 , 
    n1348 , 
    n1349 , 
    n1350 , 
    n1351 , 
    n1352 , 
    n1353 , 
    n1354 , 
    n1355 , 
    n1356 , 
    n1357 , 
    n1358 , 
    n1359 , 
    n1360 , 
    n1361 , 
    n1362 , 
    n1363 , 
    n1364 , 
    n1365 , 
    n1366 , 
    n1367 , 
    n1368 , 
    n1369 , 
    n1370 , 
    n1371 , 
    n1372 , 
    n1373 , 
    n1374 , 
    n1375 , 
    n1376 , 
    n1377 , 
    n1378 , 
    n1379 , 
    n1380 , 
    n1381 , 
    n1382 , 
    n1383 , 
    n1384 , 
    n1385 , 
    n1386 , 
    n1387 , 
    n1388 , 
    n1389 , 
    n1390 , 
    n1391 , 
    n1392 , 
    n1393 , 
    n1394 , 
    n1395 , 
    n1396 , 
    n1397 , 
    n1398 , 
    n1399 , 
    n1400 , 
    n1401 , 
    n1402 , 
    n1403 , 
    n1404 , 
    n1405 , 
    n1406 , 
    n1407 , 
    n1408 , 
    n1409 , 
    n1410 , 
    n1411 , 
    n1412 , 
    n1413 , 
    n1414 , 
    n1415 , 
    n1416 , 
    n1417 , 
    n1418 , 
    n1419 , 
    n1420 , 
    n1421 , 
    n1422 , 
    n1423 , 
    n1424 , 
    n1425 , 
    n1426 , 
    n1427 , 
    n1428 , 
    n1429 , 
    n1430 , 
    n1431 , 
    n1432 , 
    n1433 , 
    n1434 , 
    n1435 , 
    n1436 , 
    n1437 , 
    n1438 , 
    n1439 , 
    n1440 , 
    n1441 , 
    n1442 , 
    n1443 , 
    n1444 , 
    n1445 , 
    n1446 , 
    n1447 , 
    n1448 , 
    n1449 , 
    n1450 , 
    n1451 , 
    n1452 , 
    n1453 , 
    n1454 , 
    n1455 , 
    n1456 , 
    n1457 , 
    n1458 , 
    n1459 , 
    n1460 , 
    n1461 , 
    n1462 , 
    n1463 , 
    n1464 , 
    n1465 , 
    n1466 , 
    n1467 , 
    n1468 , 
    n1469 , 
    n1470 , 
    n1471 , 
    n1472 , 
    n1473 , 
    n1474 , 
    n1475 , 
    n1476 , 
    n1477 , 
    n1478 , 
    n1479 , 
    n1480 , 
    n1481 , 
    n1482 , 
    n1483 , 
    n1484 , 
    n1485 , 
    n1486 , 
    n1487 , 
    n1488 , 
    n1489 , 
    n1490 , 
    n1491 , 
    n1492 , 
    n1493 , 
    n1494 , 
    n1495 , 
    n1496 , 
    n1497 , 
    n1498 , 
    n1499 , 
    n1500 , 
    n1501 , 
    n1502 , 
    n1503 , 
    n1504 , 
    n1505 , 
    n1506 , 
    n1507 , 
    n1508 , 
    n1509 , 
    n1510 , 
    n1511 , 
    n1512 , 
    n1513 , 
    n1514 , 
    n1515 , 
    n1516 , 
    n1517 , 
    n1518 , 
    n1519 , 
    n1520 , 
    n1521 , 
    n1522 , 
    n1523 , 
    n1524 , 
    n1525 , 
    n1526 , 
    n1527 , 
    n1528 , 
    n1529 , 
    n1530 , 
    n1531 , 
    n1532 , 
    n1533 , 
    n1534 , 
    n1535 , 
    n1536 , 
    n1537 , 
    n1538 , 
    n1539 , 
    n1540 , 
    n1541 , 
    n1542 , 
    n1543 , 
    n1544 , 
    n1545 , 
    n1546 , 
    n1547 , 
    n1548 , 
    n1549 , 
    n1550 , 
    n1551 , 
    n1552 , 
    n1553 , 
    n1554 , 
    n1555 , 
    n1556 , 
    n1557 , 
    n1558 , 
    n1559 , 
    n1560 , 
    n1561 , 
    n1562 , 
    n1563 , 
    n1564 , 
    n1565 , 
    n1566 , 
    n1567 , 
    n1568 , 
    n1569 , 
    n1570 , 
    n1571 , 
    n1572 , 
    n1573 , 
    n1574 , 
    n1575 , 
    n1576 , 
    n1577 , 
    n1578 , 
    n1579 , 
    n1580 , 
    n1581 , 
    n1582 , 
    n1583 , 
    n1584 , 
    n1585 , 
    n1586 , 
    n1587 , 
    n1588 , 
    n1589 , 
    n1590 , 
    n1591 , 
    n1592 , 
    n1593 , 
    n1594 , 
    n1595 , 
    n1596 , 
    n1597 , 
    n1598 , 
    n1599 , 
    n1600 , 
    n1601 , 
    n1602 , 
    n1603 , 
    n1604 , 
    n1605 , 
    n1606 , 
    n1607 , 
    n1608 , 
    n1609 , 
    n1610 , 
    n1611 , 
    n1612 , 
    n1613 , 
    n1614 , 
    n1615 , 
    n1616 , 
    n1617 , 
    n1618 , 
    n1619 , 
    n1620 , 
    n1621 , 
    n1622 , 
    n1623 , 
    n1624 , 
    n1625 , 
    n1626 , 
    n1627 , 
    n1628 , 
    n1629 , 
    n1630 , 
    n1631 , 
    n1632 , 
    n1633 , 
    n1634 , 
    n1635 , 
    n1636 , 
    n1637 , 
    n1638 , 
    n1639 , 
    n1640 , 
    n1641 , 
    n1642 , 
    n1643 , 
    n1644 , 
    n1645 , 
    n1646 , 
    n1647 , 
    n1648 , 
    n1649 , 
    n1650 , 
    n1651 , 
    n1652 , 
    n1653 , 
    n1654 , 
    n1655 , 
    n1656 , 
    n1657 , 
    n1658 , 
    n1659 , 
    n1660 , 
    n1661 , 
    n1662 , 
    n1663 , 
    n1664 , 
    n1665 , 
    n1666 , 
    n1667 , 
    n1668 , 
    n1669 , 
    n1670 , 
    n1671 , 
    n1672 , 
    n1673 , 
    n1674 , 
    n1675 , 
    n1676 , 
    n1677 , 
    n1678 , 
    n1679 , 
    n1680 , 
    n1681 , 
    n1682 , 
    n1683 , 
    n1684 , 
    n1685 , 
    n1686 , 
    n1687 , 
    n1688 , 
    n1689 , 
    n1690 , 
    n1691 , 
    n1692 , 
    n1693 , 
    n1694 , 
    n1695 , 
    n1696 , 
    n1697 , 
    n1698 , 
    n1699 , 
    n1700 , 
    n1701 , 
    n1702 , 
    n1703 , 
    n1704 , 
    n1705 , 
    n1706 , 
    n1707 , 
    n1708 , 
    n1709 , 
    n1710 , 
    n1711 , 
    n1712 , 
    n1713 , 
    n1714 , 
    n1715 , 
    n1716 , 
    n1717 , 
    n1718 , 
    n1719 , 
    n1720 , 
    n1721 , 
    n1722 , 
    n1723 , 
    n1724 , 
    n1725 , 
    n1726 , 
    n1727 , 
    n1728 , 
    n1729 , 
    n1730 , 
    n1731 , 
    n1732 , 
    n1733 , 
    n1734 , 
    n1735 , 
    n1736 , 
    n1737 , 
    n1738 , 
    n1739 , 
    n1740 , 
    n1741 , 
    n1742 , 
    n1743 , 
    n1744 , 
    n1745 , 
    n1746 , 
    n1747 , 
    n1748 , 
    n1749 , 
    n1750 , 
    n1751 , 
    n1752 , 
    n1753 , 
    n1754 , 
    n1755 , 
    n1756 , 
    n1757 , 
    n1758 , 
    n1759 , 
    n1760 , 
    n1761 , 
    n1762 , 
    n1763 , 
    n1764 , 
    n1765 , 
    n1766 , 
    n1767 , 
    n1768 , 
    n1769 , 
    n1770 , 
    n1771 , 
    n1772 , 
    n1773 , 
    n1774 , 
    n1775 , 
    n1776 , 
    n1777 , 
    n1778 , 
    n1779 , 
    n1780 , 
    n1781 , 
    n1782 , 
    n1783 , 
    n1784 , 
    n1785 , 
    n1786 , 
    n1787 , 
    n1788 , 
    n1789 , 
    n1790 , 
    n1791 , 
    n1792 , 
    n1793 , 
    n1794 , 
    n1795 , 
    n1796 , 
    n1797 , 
    n1798 , 
    n1799 , 
    n1800 , 
    n1801 , 
    n1802 , 
    n1803 , 
    n1804 , 
    n1805 , 
    n1806 , 
    n1807 , 
    n1808 , 
    n1809 , 
    n1810 , 
    n1811 , 
    n1812 , 
    n1813 , 
    n1814 , 
    n1815 , 
    n1816 , 
    n1817 , 
    n1818 , 
    n1819 , 
    n1820 , 
    n1821 , 
    n1822 , 
    n1823 , 
    n1824 , 
    n1825 , 
    n1826 , 
    n1827 , 
    n1828 , 
    n1829 , 
    n1830 , 
    n1831 , 
    n1832 , 
    n1833 , 
    n1834 , 
    n1835 , 
    n1836 , 
    n1837 , 
    n1838 , 
    n1839 , 
    n1840 , 
    n1841 , 
    n1842 , 
    n1843 , 
    n1844 , 
    n1845 , 
    n1846 , 
    n1847 , 
    n1848 , 
    n1849 , 
    n1850 , 
    n1851 , 
    n1852 , 
    n1853 , 
    n1854 , 
    n1855 , 
    n1856 , 
    n1857 , 
    n1858 , 
    n1859 , 
    n1860 , 
    n1861 , 
    n1862 , 
    n1863 , 
    n1864 , 
    n1865 , 
    n1866 , 
    n1867 , 
    n1868 , 
    n1869 , 
    n1870 , 
    n1871 , 
    n1872 , 
    n1873 , 
    n1874 , 
    n1875 , 
    n1876 , 
    n1877 , 
    n1878 , 
    n1879 , 
    n1880 , 
    n1881 , 
    n1882 , 
    n1883 , 
    n1884 , 
    n1885 , 
    n1886 , 
    n1887 , 
    n1888 , 
    n1889 , 
    n1890 , 
    n1891 , 
    n1892 , 
    n1893 , 
    n1894 , 
    n1895 , 
    n1896 , 
    n1897 , 
    n1898 , 
    n1899 , 
    n1900 , 
    n1901 , 
    n1902 , 
    n1903 , 
    n1904 , 
    n1905 , 
    n1906 , 
    n1907 , 
    n1908 , 
    n1909 , 
    n1910 , 
    n1911 , 
    n1912 , 
    n1913 , 
    n1914 , 
    n1915 , 
    n1916 , 
    n1917 , 
    n1918 , 
    n1919 , 
    n1920 , 
    n1921 , 
    n1922 , 
    n1923 , 
    n1924 , 
    n1925 , 
    n1926 , 
    n1927 , 
    n1928 , 
    n1929 , 
    n1930 , 
    n1931 , 
    n1932 , 
    n1933 , 
    n1934 , 
    n1935 , 
    n1936 , 
    n1937 , 
    n1938 , 
    n1939 , 
    n1940 , 
    n1941 , 
    n1942 , 
    n1943 , 
    n1944 , 
    n1945 , 
    n1946 , 
    n1947 , 
    n1948 , 
    n1949 , 
    n1950 , 
    n1951 , 
    n1952 , 
    n1953 , 
    n1954 , 
    n1955 , 
    n1956 , 
    n1957 , 
    n1958 , 
    n1959 , 
    n1960 , 
    n1961 , 
    n1962 , 
    n1963 , 
    n1964 , 
    n1965 , 
    n1966 , 
    n1967 , 
    n1968 , 
    n1969 , 
    n1970 , 
    n1971 , 
    n1972 , 
    n1973 , 
    n1974 , 
    n1975 , 
    n1976 , 
    n1977 , 
    n1978 , 
    n1979 , 
    n1980 , 
    n1981 , 
    n1982 , 
    n1983 , 
    n1984 , 
    n1985 , 
    n1986 , 
    n1987 , 
    n1988 , 
    n1989 , 
    n1990 , 
    n1991 , 
    n1992 , 
    n1993 , 
    n1994 , 
    n1995 , 
    n1996 , 
    n1997 , 
    n1998 , 
    n1999 , 
    n2000 , 
    n2001 , 
    n2002 , 
    n2003 , 
    n2004 , 
    n2005 , 
    n2006 , 
    n2007 , 
    n2008 , 
    n2009 , 
    n2010 , 
    n2011 , 
    n2012 , 
    n2013 , 
    n2014 , 
    n2015 , 
    n2016 , 
    n2017 , 
    n2018 , 
    n2019 , 
    n2020 , 
    n2021 , 
    n2022 , 
    n2023 , 
    n2024 , 
    n2025 , 
    n2026 , 
    n2027 , 
    n2028 , 
    n2029 , 
    n2030 , 
    n2031 , 
    n2032 , 
    n2033 , 
    n2034 , 
    n2035 , 
    n2036 , 
    n2037 , 
    n2038 , 
    n2039 , 
    n2040 , 
    n2041 , 
    n2042 , 
    n2043 , 
    n2044 , 
    n2045 , 
    n2046 , 
    n2047 , 
    n2048 , 
    n2049 , 
    n2050 , 
    n2051 , 
    n2052 , 
    n2053 , 
    n2054 , 
    n2055 , 
    n2056 , 
    n2057 , 
    n2058 , 
    n2059 , 
    n2060 , 
    n2061 , 
    n2062 , 
    n2063 , 
    n2064 , 
    n2065 , 
    n2066 , 
    n2067 , 
    n2068 , 
    n2069 , 
    n2070 , 
    n2071 , 
    n2072 , 
    n2073 , 
    n2074 , 
    n2075 , 
    n2076 , 
    n2077 , 
    n2078 , 
    n2079 , 
    n2080 , 
    n2081 , 
    n2082 , 
    n2083 , 
    n2084 , 
    n2085 , 
    n2086 , 
    n2087 , 
    n2088 , 
    n2089 , 
    n2090 , 
    n2091 , 
    n2092 , 
    n2093 , 
    n2094 , 
    n2095 , 
    n2096 , 
    n2097 , 
    n2098 , 
    n2099 , 
    n2100 , 
    n2101 , 
    n2102 , 
    n2103 , 
    n2104 , 
    n2105 , 
    n2106 , 
    n2107 , 
    n2108 , 
    n2109 , 
    n2110 , 
    n2111 , 
    n2112 , 
    n2113 , 
    n2114 , 
    n2115 , 
    n2116 , 
    n2117 , 
    n2118 , 
    n2119 , 
    n2120 , 
    n2121 , 
    n2122 , 
    n2123 , 
    n2124 , 
    n2125 , 
    n2126 , 
    n2127 , 
    n2128 , 
    n2129 , 
    n2130 , 
    n2131 , 
    n2132 , 
    n2133 , 
    n2134 , 
    n2135 , 
    n2136 , 
    n2137 , 
    n2138 , 
    n2139 , 
    n2140 , 
    n2141 , 
    n2142 , 
    n2143 , 
    n2144 , 
    n2145 , 
    n2146 , 
    n2147 , 
    n2148 , 
    n2149 , 
    n2150 , 
    n2151 , 
    n2152 , 
    n2153 , 
    n2154 , 
    n2155 , 
    n2156 , 
    n2157 , 
    n2158 , 
    n2159 , 
    n2160 , 
    n2161 , 
    n2162 , 
    n2163 , 
    n2164 , 
    n2165 , 
    n2166 , 
    n2167 , 
    n2168 , 
    n2169 , 
    n2170 , 
    n2171 , 
    n2172 , 
    n2173 , 
    n2174 , 
    n2175 , 
    n2176 , 
    n2177 , 
    n2178 , 
    n2179 , 
    n2180 , 
    n2181 , 
    n2182 , 
    n2183 , 
    n2184 , 
    n2185 , 
    n2186 , 
    n2187 , 
    n2188 , 
    n2189 , 
    n2190 , 
    n2191 , 
    n2192 , 
    n2193 , 
    n2194 , 
    n2195 , 
    n2196 , 
    n2197 , 
    n2198 , 
    n2199 , 
    n2200 , 
    n2201 , 
    n2202 , 
    n2203 , 
    n2204 , 
    n2205 , 
    n2206 , 
    n2207 , 
    n2208 , 
    n2209 , 
    n2210 , 
    n2211 , 
    n2212 , 
    n2213 , 
    n2214 , 
    n2215 , 
    n2216 , 
    n2217 , 
    n2218 , 
    n2219 , 
    n2220 , 
    n2221 , 
    n2222 , 
    n2223 , 
    n2224 , 
    n2225 , 
    n2226 , 
    n2227 , 
    n2228 , 
    n2229 , 
    n2230 , 
    n2231 , 
    n2232 , 
    n2233 , 
    n2234 , 
    n2235 , 
    n2236 , 
    n2237 , 
    n2238 , 
    n2239 , 
    n2240 , 
    n2241 , 
    n2242 , 
    n2243 , 
    n2244 , 
    n2245 , 
    n2246 , 
    n2247 , 
    n2248 , 
    n2249 , 
    n2250 , 
    n2251 , 
    n2252 , 
    n2253 , 
    n2254 , 
    n2255 , 
    n2256 , 
    n2257 , 
    n2258 , 
    n2259 , 
    n2260 , 
    n2261 , 
    n2262 , 
    n2263 , 
    n2264 , 
    n2265 , 
    n2266 , 
    n2267 , 
    n2268 , 
    n2269 , 
    n2270 , 
    n2271 , 
    n2272 , 
    n2273 , 
    n2274 , 
    n2275 , 
    n2276 , 
    n2277 , 
    n2278 , 
    n2279 , 
    n2280 , 
    n2281 , 
    n2282 , 
    n2283 , 
    n2284 , 
    n2285 , 
    n2286 , 
    n2287 , 
    n2288 , 
    n2289 , 
    n2290 , 
    n2291 , 
    n2292 , 
    n2293 , 
    n2294 , 
    n2295 , 
    n2296 , 
    n2297 , 
    n2298 , 
    n2299 , 
    n2300 , 
    n2301 , 
    n2302 , 
    n2303 , 
    n2304 , 
    n2305 , 
    n2306 , 
    n2307 , 
    n2308 , 
    n2309 , 
    n2310 , 
    n2311 , 
    n2312 , 
    n2313 , 
    n2314 , 
    n2315 , 
    n2316 , 
    n2317 , 
    n2318 , 
    n2319 , 
    n2320 , 
    n2321 , 
    n2322 , 
    n2323 , 
    n2324 , 
    n2325 , 
    n2326 , 
    n2327 , 
    n2328 , 
    n2329 , 
    n2330 , 
    n2331 , 
    n2332 , 
    n2333 , 
    n2334 , 
    n2335 , 
    n2336 , 
    n2337 , 
    n2338 , 
    n2339 , 
    n2340 , 
    n2341 , 
    n2342 , 
    n2343 , 
    n2344 , 
    n2345 , 
    n2346 , 
    n2347 , 
    n2348 , 
    n2349 , 
    n2350 , 
    n2351 , 
    n2352 , 
    n2353 , 
    n2354 , 
    n2355 , 
    n2356 , 
    n2357 , 
    n2358 , 
    n2359 , 
    n2360 , 
    n2361 , 
    n2362 , 
    n2363 , 
    n2364 , 
    n2365 , 
    n2366 , 
    n2367 , 
    n2368 , 
    n2369 , 
    n2370 , 
    n2371 , 
    n2372 , 
    n2373 , 
    n2374 , 
    n2375 , 
    n2376 , 
    n2377 , 
    n2378 , 
    n2379 , 
    n2380 , 
    n2381 , 
    n2382 , 
    n2383 , 
    n2384 , 
    n2385 , 
    n2386 , 
    n2387 , 
    n2388 , 
    n2389 , 
    n2390 , 
    n2391 , 
    n2392 , 
    n2393 , 
    n2394 , 
    n2395 , 
    n2396 , 
    n2397 , 
    n2398 , 
    n2399 , 
    n2400 , 
    n2401 , 
    n2402 , 
    n2403 , 
    n2404 , 
    n2405 , 
    n2406 , 
    n2407 , 
    n2408 , 
    n2409 , 
    n2410 , 
    n2411 , 
    n2412 , 
    n2413 , 
    n2414 , 
    n2415 , 
    n2416 , 
    n2417 , 
    n2418 , 
    n2419 , 
    n2420 , 
    n2421 , 
    n2422 , 
    n2423 , 
    n2424 , 
    n2425 , 
    n2426 , 
    n2427 , 
    n2428 , 
    n2429 , 
    n2430 , 
    n2431 , 
    n2432 , 
    n2433 , 
    n2434 , 
    n2435 , 
    n2436 , 
    n2437 , 
    n2438 , 
    n2439 , 
    n2440 , 
    n2441 , 
    n2442 , 
    n2443 , 
    n2444 , 
    n2445 , 
    n2446 , 
    n2447 , 
    n2448 , 
    n2449 , 
    n2450 , 
    n2451 , 
    n2452 , 
    n2453 , 
    n2454 , 
    n2455 , 
    n2456 , 
    n2457 , 
    n2458 , 
    n2459 , 
    n2460 , 
    n2461 , 
    n2462 , 
    n2463 , 
    n2464 , 
    n2465 , 
    n2466 , 
    n2467 , 
    n2468 , 
    n2469 , 
    n2470 , 
    n2471 , 
    n2472 , 
    n2473 , 
    n2474 , 
    n2475 , 
    n2476 , 
    n2477 , 
    n2478 , 
    n2479 , 
    n2480 , 
    n2481 , 
    n2482 , 
    n2483 , 
    n2484 , 
    n2485 , 
    n2486 , 
    n2487 , 
    n2488 , 
    n2489 , 
    n2490 , 
    n2491 , 
    n2492 , 
    n2493 , 
    n2494 , 
    n2495 , 
    n2496 , 
    n2497 , 
    n2498 , 
    n2499 , 
    n2500 , 
    n2501 , 
    n2502 , 
    n2503 , 
    n2504 , 
    n2505 , 
    n2506 , 
    n2507 , 
    n2508 , 
    n2509 , 
    n2510 , 
    n2511 , 
    n2512 , 
    n2513 , 
    n2514 , 
    n2515 , 
    n2516 , 
    n2517 , 
    n2518 , 
    n2519 , 
    n2520 , 
    n2521 , 
    n2522 , 
    n2523 , 
    n2524 , 
    n2525 , 
    n2526 , 
    n2527 , 
    n2528 , 
    n2529 , 
    n2530 , 
    n2531 , 
    n2532 , 
    n2533 , 
    n2534 , 
    n2535 , 
    n2536 , 
    n2537 , 
    n2538 , 
    n2539 , 
    n2540 , 
    n2541 , 
    n2542 , 
    n2543 , 
    n2544 , 
    n2545 , 
    n2546 , 
    n2547 , 
    n2548 , 
    n2549 , 
    n2550 , 
    n2551 , 
    n2552 , 
    n2553 , 
    n2554 , 
    n2555 , 
    n2556 , 
    n2557 , 
    n2558 , 
    n2559 , 
    n2560 , 
    n2561 , 
    n2562 , 
    n2563 , 
    n2564 , 
    n2565 , 
    n2566 , 
    n2567 , 
    n2568 , 
    n2569 , 
    n2570 , 
    n2571 , 
    n2572 , 
    n2573 , 
    n2574 , 
    n2575 , 
    n2576 , 
    n2577 , 
    n2578 , 
    n2579 , 
    n2580 , 
    n2581 , 
    n2582 , 
    n2583 , 
    n2584 , 
    n2585 , 
    n2586 , 
    n2587 , 
    n2588 , 
    n2589 , 
    n2590 , 
    n2591 , 
    n2592 , 
    n2593 , 
    n2594 , 
    n2595 , 
    n2596 , 
    n2597 , 
    n2598 , 
    n2599 , 
    n2600 , 
    n2601 , 
    n2602 , 
    n2603 , 
    n2604 , 
    n2605 , 
    n2606 , 
    n2607 , 
    n2608 , 
    n2609 , 
    n2610 , 
    n2611 , 
    n2612 , 
    n2613 , 
    n2614 , 
    n2615 , 
    n2616 , 
    n2617 , 
    n2618 , 
    n2619 , 
    n2620 , 
    n2621 , 
    n2622 , 
    n2623 , 
    n2624 , 
    n2625 , 
    n2626 , 
    n2627 , 
    n2628 , 
    n2629 , 
    n2630 , 
    n2631 , 
    n2632 , 
    n2633 , 
    n2634 , 
    n2635 , 
    n2636 , 
    n2637 , 
    n2638 , 
    n2639 , 
    n2640 , 
    n2641 , 
    n2642 , 
    n2643 , 
    n2644 , 
    n2645 , 
    n2646 , 
    n2647 , 
    n2648 , 
    n2649 , 
    n2650 , 
    n2651 , 
    n2652 , 
    n2653 , 
    n2654 , 
    n2655 , 
    n2656 , 
    n2657 , 
    n2658 , 
    n2659 , 
    n2660 , 
    n2661 , 
    n2662 , 
    n2663 , 
    n2664 , 
    n2665 , 
    n2666 , 
    n2667 , 
    n2668 , 
    n2669 , 
    n2670 , 
    n2671 , 
    n2672 , 
    n2673 , 
    n2674 , 
    n2675 , 
    n2676 , 
    n2677 , 
    n2678 , 
    n2679 , 
    n2680 , 
    n2681 , 
    n2682 , 
    n2683 , 
    n2684 , 
    n2685 , 
    n2686 , 
    n2687 , 
    n2688 , 
    n2689 , 
    n2690 , 
    n2691 , 
    n2692 , 
    n2693 , 
    n2694 , 
    n2695 , 
    n2696 , 
    n2697 , 
    n2698 , 
    n2699 , 
    n2700 , 
    n2701 , 
    n2702 , 
    n2703 , 
    n2704 , 
    n2705 , 
    n2706 , 
    n2707 , 
    n2708 , 
    n2709 , 
    n2710 , 
    n2711 , 
    n2712 , 
    n2713 , 
    n2714 , 
    n2715 , 
    n2716 , 
    n2717 , 
    n2718 , 
    n2719 , 
    n2720 , 
    n2721 , 
    n2722 , 
    n2723 , 
    n2724 , 
    n2725 , 
    n2726 , 
    n2727 , 
    n2728 , 
    n2729 , 
    n2730 , 
    n2731 , 
    n2732 , 
    n2733 , 
    n2734 , 
    n2735 , 
    n2736 , 
    n2737 , 
    n2738 , 
    n2739 , 
    n2740 , 
    n2741 , 
    n2742 , 
    n2743 , 
    n2744 , 
    n2745 , 
    n2746 , 
    n2747 , 
    n2748 , 
    n2749 , 
    n2750 , 
    n2751 , 
    n2752 , 
    n2753 , 
    n2754 , 
    n2755 , 
    n2756 , 
    n2757 , 
    n2758 , 
    n2759 , 
    n2760 , 
    n2761 , 
    n2762 , 
    n2763 , 
    n2764 , 
    n2765 , 
    n2766 , 
    n2767 , 
    n2768 , 
    n2769 , 
    n2770 , 
    n2771 , 
    n2772 , 
    n2773 , 
    n2774 , 
    n2775 , 
    n2776 , 
    n2777 , 
    n2778 , 
    n2779 , 
    n2780 , 
    n2781 , 
    n2782 , 
    n2783 , 
    n2784 , 
    n2785 , 
    n2786 , 
    n2787 , 
    n2788 , 
    n2789 , 
    n2790 , 
    n2791 , 
    n2792 , 
    n2793 , 
    n2794 , 
    n2795 , 
    n2796 , 
    n2797 , 
    n2798 , 
    n2799 , 
    n2800 , 
    n2801 , 
    n2802 , 
    n2803 , 
    n2804 , 
    n2805 , 
    n2806 , 
    n2807 , 
    n2808 , 
    n2809 , 
    n2810 , 
    n2811 , 
    n2812 , 
    n2813 , 
    n2814 , 
    n2815 , 
    n2816 , 
    n2817 , 
    n2818 , 
    n2819 , 
    n2820 , 
    n2821 , 
    n2822 , 
    n2823 , 
    n2824 , 
    n2825 , 
    n2826 , 
    n2827 , 
    n2828 , 
    n2829 , 
    n2830 , 
    n2831 , 
    n2832 , 
    n2833 , 
    n2834 , 
    n2835 , 
    n2836 , 
    n2837 , 
    n2838 , 
    n2839 , 
    n2840 , 
    n2841 , 
    n2842 , 
    n2843 , 
    n2844 , 
    n2845 , 
    n2846 , 
    n2847 , 
    n2848 , 
    n2849 , 
    n2850 , 
    n2851 , 
    n2852 , 
    n2853 , 
    n2854 , 
    n2855 , 
    n2856 , 
    n2857 , 
    n2858 , 
    n2859 , 
    n2860 , 
    n2861 , 
    n2862 , 
    n2863 , 
    n2864 , 
    n2865 , 
    n2866 , 
    n2867 , 
    n2868 , 
    n2869 , 
    n2870 , 
    n2871 , 
    n2872 , 
    n2873 , 
    n2874 , 
    n2875 , 
    n2876 , 
    n2877 , 
    n2878 , 
    n2879 , 
    n2880 , 
    n2881 , 
    n2882 , 
    n2883 , 
    n2884 , 
    n2885 , 
    n2886 , 
    n2887 , 
    n2888 , 
    n2889 , 
    n2890 , 
    n2891 , 
    n2892 , 
    n2893 , 
    n2894 , 
    n2895 , 
    n2896 , 
    n2897 , 
    n2898 , 
    n2899 , 
    n2900 , 
    n2901 , 
    n2902 , 
    n2903 , 
    n2904 , 
    n2905 , 
    n2906 , 
    n2907 , 
    n2908 , 
    n2909 , 
    n2910 , 
    n2911 , 
    n2912 , 
    n2913 , 
    n2914 , 
    n2915 , 
    n2916 , 
    n2917 , 
    n2918 , 
    n2919 , 
    n2920 , 
    n2921 , 
    n2922 , 
    n2923 , 
    n2924 , 
    n2925 , 
    n2926 , 
    n2927 , 
    n2928 , 
    n2929 , 
    n2930 , 
    n2931 , 
    n2932 , 
    n2933 , 
    n2934 , 
    n2935 , 
    n2936 , 
    n2937 , 
    n2938 , 
    n2939 , 
    n2940 , 
    n2941 , 
    n2942 , 
    n2943 , 
    n2944 , 
    n2945 , 
    n2946 , 
    n2947 , 
    n2948 , 
    n2949 , 
    n2950 , 
    n2951 , 
    n2952 , 
    n2953 , 
    n2954 , 
    n2955 , 
    n2956 , 
    n2957 , 
    n2958 , 
    n2959 , 
    n2960 , 
    n2961 , 
    n2962 , 
    n2963 , 
    n2964 , 
    n2965 , 
    n2966 , 
    n2967 , 
    n2968 , 
    n2969 , 
    n2970 , 
    n2971 , 
    n2972 , 
    n2973 , 
    n2974 , 
    n2975 , 
    n2976 , 
    n2977 , 
    n2978 , 
    n2979 , 
    n2980 , 
    n2981 , 
    n2982 , 
    n2983 , 
    n2984 , 
    n2985 , 
    n2986 , 
    n2987 , 
    n2988 , 
    n2989 , 
    n2990 , 
    n2991 , 
    n2992 , 
    n2993 , 
    n2994 , 
    n2995 , 
    n2996 , 
    n2997 , 
    n2998 , 
    n2999 , 
    n3000 , 
    n3001 , 
    n3002 , 
    n3003 , 
    n3004 , 
    n3005 , 
    n3006 , 
    n3007 , 
    n3008 , 
    n3009 , 
    n3010 , 
    n3011 , 
    n3012 , 
    n3013 , 
    n3014 , 
    n3015 , 
    n3016 , 
    n3017 , 
    n3018 , 
    n3019 , 
    n3020 , 
    n3021 , 
    n3022 , 
    n3023 , 
    n3024 , 
    n3025 , 
    n3026 , 
    n3027 , 
    n3028 , 
    n3029 , 
    n3030 , 
    n3031 , 
    n3032 , 
    n3033 , 
    n3034 , 
    n3035 , 
    n3036 , 
    n3037 , 
    n3038 , 
    n3039 , 
    n3040 , 
    n3041 , 
    n3042 , 
    n3043 , 
    n3044 , 
    n3045 , 
    n3046 , 
    n3047 , 
    n3048 , 
    n3049 , 
    n3050 , 
    n3051 , 
    n3052 , 
    n3053 , 
    n3054 , 
    n3055 , 
    n3056 , 
    n3057 , 
    n3058 , 
    n3059 , 
    n3060 , 
    n3061 , 
    n3062 , 
    n3063 , 
    n3064 , 
    n3065 , 
    n3066 , 
    n3067 , 
    n3068 , 
    n3069 , 
    n3070 , 
    n3071 , 
    n3072 , 
    n3073 , 
    n3074 , 
    n3075 , 
    n3076 , 
    n3077 , 
    n3078 , 
    n3079 , 
    n3080 , 
    n3081 , 
    n3082 , 
    n3083 , 
    n3084 , 
    n3085 , 
    n3086 , 
    n3087 , 
    n3088 , 
    n3089 , 
    n3090 , 
    n3091 , 
    n3092 , 
    n3093 , 
    n3094 , 
    n3095 , 
    n3096 , 
    n3097 , 
    n3098 , 
    n3099 , 
    n3100 , 
    n3101 , 
    n3102 , 
    n3103 , 
    n3104 , 
    n3105 , 
    n3106 , 
    n3107 , 
    n3108 , 
    n3109 , 
    n3110 , 
    n3111 , 
    n3112 , 
    n3113 , 
    n3114 , 
    n3115 , 
    n3116 , 
    n3117 , 
    n3118 , 
    n3119 , 
    n3120 , 
    n3121 , 
    n3122 , 
    n3123 ;

wire  C0 , RI21a19c60_2 , 
    RI21a5daf0_1 , 
    RI2107e620_463 , 
    RI210bf4e0_288 , 
    RI21078b30_503 , 
    RI21a13090_74 , 
    RI210bf558_287 , 
    RI21078ba8_502 , 
    RI21a13108_73 , 
    RI21a116c8_87 , 
    RI210bd6e0_301 , 
    RI21077078_516 , 
    RI21a11dd0_86 , 
    RI210bd758_300 , 
    RI210770f0_515 , 
    RI21a11e48_85 , 
    RI210bd7d0_299 , 
    RI21077168_514 , 
    RI21a132e8_69 , 
    RI210bff30_283 , 
    RI210797d8_498 , 
    RI210bfeb8_284 , 
    RI21079760_499 , 
    RI21a13270_70 , 
    RI210be1a8_295 , 
    RI21077d98_510 , 
    RI21a12028_81 , 
    RI21a12730_80 , 
    RI210bea18_294 , 
    RI21077e10_509 , 
    RI21a127a8_79 , 
    RI210bea90_293 , 
    RI21077e88_508 , 
    RI21079850_497 , 
    RI21a139f0_68 , 
    RI21084368_418 , 
    RI21a11f38_83 , 
    RI210be0b8_297 , 
    RI21077258_512 , 
    RI21a11fb0_82 , 
    RI210be130_296 , 
    RI21077d20_511 , 
    RI210be040_298 , 
    RI210771e0_513 , 
    RI21a11ec0_84 , 
    RI21a13180_72 , 
    RI210bfdc8_286 , 
    RI21078c20_501 , 
    RI21a131f8_71 , 
    RI210bfe40_285 , 
    RI21078c98_500 , 
    RI2107a660_489 , 
    RI2107cd48_472 , 
    RI2106bde0_608 , 
    RI2107c118_476 , 
    RI2107a570_491 , 
    RI21079940_495 , 
    RI2107a5e8_490 , 
    RI2107d900_469 , 
    RI2107b1a0_487 , 
    RI2107d978_468 , 
    RI2107a480_493 , 
    RI2107da68_466 , 
    RI210799b8_494 , 
    RI2107d9f0_467 , 
    RI2107a4f8_492 , 
    RI210798c8_496 , 
    RI2107ce38_470 , 
    RI2107cdc0_471 , 
    RI2107ccd0_473 , 
    RI2107cc58_474 , 
    RI2107c028_478 , 
    RI2107cbe0_475 , 
    RI2107c0a0_477 , 
    RI2107bfb0_479 , 
    RI2107b3f8_482 , 
    RI2107bf38_480 , 
    RI2107bec0_481 , 
    RI2107b380_483 , 
    RI2107b308_484 , 
    RI2107b218_486 , 
    RI2107b290_485 , 
    RI2107a6d8_488 , 
    RI2106be58_607 , 
    RI2107dae0_465 , 
    RI2106ddc0_566 , 
    RI210730b8_542 , 
    RI2106cc68_590 , 
    RI2106a2b0_640 , 
    RI21069ab8_644 , 
    RI2106bfc0_604 , 
    RI2106c038_603 , 
    RI2106a148_643 , 
    RI2106bf48_605 , 
    RI21069a40_645 , 
    RI2106a760_630 , 
    RI2106a5f8_633 , 
    RI2106a670_632 , 
    RI2106bed0_606 , 
    RI2106a7d8_629 , 
    RI2106c308_597 , 
    RI2106ae68_628 , 
    RI2106a6e8_631 , 
    RI2106a580_634 , 
    RI2106a508_635 , 
    RI2106a490_636 , 
    RI2106a3a0_638 , 
    RI2106a328_639 , 
    RI2106a238_641 , 
    RI2106c290_598 , 
    RI2106c218_599 , 
    RI2106c1a0_600 , 
    RI2106c128_601 , 
    RI2106c0b0_602 , 
    RI2106dd48_567 , 
    RI21073040_543 , 
    RI2106cbf0_591 , 
    RI21a12820_78 , 
    RI210beb08_292 , 
    RI21a0e608_121 , 
    RI21077f00_507 , 
    RI210b87a8_334 , 
    RI21a11560_90 , 
    RI210bcd80_304 , 
    RI210cfcc8_237 , 
    RI210842f0_419 , 
    RI21a0efe0_114 , 
    RI210b92e8_327 , 
    RI21a0f148_111 , 
    RI21084278_420 , 
    RI21a0ef68_115 , 
    RI210b9270_328 , 
    RI21a0eef0_116 , 
    RI210b91f8_329 , 
    RI21a0e680_120 , 
    RI210b8820_333 , 
    RI21a0e6f8_119 , 
    RI210b8898_332 , 
    RI21a10c00_96 , 
    RI210bc2b8_310 , 
    RI21a11470_92 , 
    RI210bcc90_306 , 
    RI21a10cf0_94 , 
    RI210bc3a8_308 , 
    RI21a0e770_118 , 
    RI210b8910_331 , 
    RI21a10c78_95 , 
    RI210bc330_309 , 
    RI21a114e8_91 , 
    RI210bcd08_305 , 
    RI21a10d68_93 , 
    RI210bc420_307 , 
    RI21a0e7e8_117 , 
    RI210b9180_330 , 
    RI21a102a0_102 , 
    RI210baff8_316 , 
    RI21a10318_101 , 
    RI210bb070_315 , 
    RI21a101b0_104 , 
    RI210baf08_318 , 
    RI21a10228_103 , 
    RI210baf80_317 , 
    RI21a10390_100 , 
    RI210bb8e0_314 , 
    RI21a10408_99 , 
    RI210bb958_313 , 
    RI21a10b10_98 , 
    RI210bb9d0_312 , 
    RI21a10b88_97 , 
    RI210bba48_311 , 
    RI21a0f940_108 , 
    RI210ba530_322 , 
    RI21a0f9b8_107 , 
    RI210ba5a8_321 , 
    RI21a0fa30_106 , 
    RI210ba620_320 , 
    RI21a0faa8_105 , 
    RI210ba698_319 , 
    RI21a0f850_110 , 
    RI210b9c48_324 , 
    RI21a0f8c8_109 , 
    RI210b9cc0_323 , 
    RI21a0f0d0_112 , 
    RI210b9bd0_325 , 
    RI21a19990_4 , 
    RI2106cd58_588 , 
    RI2106deb0_564 , 
    RI21073c70_539 , 
    RI21a198a0_6 , 
    RI2106de38_565 , 
    RI21073bf8_540 , 
    RI2106cce0_589 , 
    RI21a19918_5 , 
    RI21a0f058_113 , 
    RI210b9b58_326 , 
    RI21a19a08_3 , 
    RI21a197b0_8 , 
    RI2106ce48_586 , 
    RI21073d60_537 , 
    RI2106dfa0_562 , 
    RI2106df28_563 , 
    RI2106cdd0_587 , 
    RI21073ce8_538 , 
    RI21a19828_7 , 
    RI2106cec0_585 , 
    RI21073dd8_536 , 
    RI2106e018_561 , 
    RI21a190a8_9 , 
    RI210748a0_535 , 
    RI2106e090_560 , 
    RI2106cf38_584 , 
    RI21a19030_10 , 
    RI2106cfb0_583 , 
    RI21074918_534 , 
    RI2106e108_559 , 
    RI21a18fb8_11 , 
    RI21074990_533 , 
    RI21070a48_558 , 
    RI2106d028_582 , 
    RI21a18f40_12 , 
    RI21a18e50_14 , 
    RI2106d118_580 , 
    RI21074a80_531 , 
    RI21071588_556 , 
    RI21070ac0_557 , 
    RI2106d0a0_581 , 
    RI21074a08_532 , 
    RI21a18ec8_13 , 
    RI21a186d0_16 , 
    RI2106b1b0_621 , 
    RI21075638_528 , 
    RI2106b570_613 , 
    RI2106b4f8_614 , 
    RI2106b138_622 , 
    RI210755c0_529 , 
    RI21a18748_15 , 
    RI2106bc00_612 , 
    RI210756b0_527 , 
    RI2106b228_620 , 
    RI21a18658_17 , 
    RI2106d190_579 , 
    RI21075728_526 , 
    RI21071600_555 , 
    RI21a185e0_18 , 
    RI21a17410_28 , 
    RI21072e60_547 , 
    RI2106af58_626 , 
    RI2106dcd0_568 , 
    RI2106dc58_569 , 
    RI21072398_548 , 
    RI2106aee0_627 , 
    RI21a17488_27 , 
    RI21a17320_30 , 
    RI21072f50_545 , 
    RI2106afd0_625 , 
    RI2106b318_618 , 
    RI2106cb00_593 , 
    RI2106b2a0_619 , 
    RI21072ed8_546 , 
    RI21a17398_29 , 
    RI21a16b28_33 , 
    RI2106b0c0_623 , 
    RI2106b480_615 , 
    RI21074af8_530 , 
    RI2106a418_637 , 
    RI21072230_551 , 
    RI210764c0_519 , 
    RI2106c380_596 , 
    RI2106daf0_572 , 
    RI21a16ab0_34 , 
    RI2106cb78_592 , 
    RI21072fc8_544 , 
    RI2106b390_617 , 
    RI21a172a8_31 , 
    RI2106b048_624 , 
    RI2106b408_616 , 
    RI21073b80_541 , 
    RI2106a1c0_642 , 
    RI21a17230_32 , 
    RI21a184f0_20 , 
    RI2106d898_577 , 
    RI2106bc78_611 , 
    RI21075818_524 , 
    RI210757a0_525 , 
    RI2106d208_578 , 
    RI21071678_554 , 
    RI21a18568_19 , 
    RI21a17d70_22 , 
    RI210716f0_553 , 
    RI2106d988_575 , 
    RI21076358_522 , 
    RI2106d910_576 , 
    RI2106bcf0_610 , 
    RI210762e0_523 , 
    RI21a17de8_21 , 
    RI210721b8_552 , 
    RI2106da00_574 , 
    RI210763d0_521 , 
    RI21a17cf8_23 , 
    RI2106da78_573 , 
    RI21076448_520 , 
    RI2106bd68_609 , 
    RI21a17c80_24 , 
    RI21a17b90_26 , 
    RI2106ca88_594 , 
    RI21072320_549 , 
    RI2106dbe0_570 , 
    RI2106ca10_595 , 
    RI210722a8_550 , 
    RI2106db68_571 , 
    RI21a17c08_25 , 
    RI21a14440_60 , 
    RI21a15f70_44 , 
    RI21a14350_62 , 
    RI21a13ae0_66 , 
    RI21a13b58_65 , 
    RI21a168d0_38 , 
    RI21a13bd0_64 , 
    RI21a16948_37 , 
    RI21a169c0_36 , 
    RI21a15778_47 , 
    RI21a15fe8_43 , 
    RI21a16150_40 , 
    RI21a143c8_61 , 
    RI21a161c8_39 , 
    RI21a14530_58 , 
    RI21a16060_42 , 
    RI21a160d8_41 , 
    RI21a13a68_67 , 
    RI21a13c48_63 , 
    RI21a15868_45 , 
    RI21a15688_49 , 
    RI21a15700_48 , 
    RI21a157f0_46 , 
    RI21a15610_50 , 
    RI21a14f08_51 , 
    RI21a14e90_52 , 
    RI21a14e18_53 , 
    RI21a14da0_54 , 
    RI21a14d28_55 , 
    RI21a145a8_57 , 
    RI21a14cb0_56 , 
    RI21a144b8_59 , 
    RI210d8710_180 , 
    RI21a0b6b0_152 , 
    RI210d41b0_209 , 
    RI21a0de10_124 , 
    RI210d8788_179 , 
    RI21a0b728_151 , 
    RI210d4228_208 , 
    RI21a0de88_123 , 
    RI210d37d8_213 , 
    RI210d7d38_184 , 
    RI21a0ae40_156 , 
    RI21a0dc30_128 , 
    RI21a0aeb8_155 , 
    RI210d7db0_183 , 
    RI210d3850_212 , 
    RI21a0dca8_127 , 
    RI210d5560_201 , 
    RI210d9b38_171 , 
    RI210d1078_229 , 
    RI21a0c100_144 , 
    RI210d9160_175 , 
    RI210d4b88_205 , 
    RI210d06a0_233 , 
    RI21a0b908_147 , 
    RI210d4c00_204 , 
    RI210d99d0_174 , 
    RI210d0718_232 , 
    RI21a0c010_146 , 
    RI210d42a0_207 , 
    RI210d9070_177 , 
    RI210cfdb8_235 , 
    RI21a0b818_149 , 
    RI210d4b10_206 , 
    RI210d90e8_176 , 
    RI210d0628_234 , 
    RI21a0b890_148 , 
    RI210d54e8_202 , 
    RI210d9ac0_172 , 
    RI210d1000_230 , 
    RI210cf2f0_241 , 
    RI210d4c78_203 , 
    RI210d9a48_173 , 
    RI210d0790_231 , 
    RI21a0c088_145 , 
    RI21a0af30_154 , 
    RI210d8620_182 , 
    RI210d38c8_211 , 
    RI21a0dd20_126 , 
    RI210d4138_210 , 
    RI210d8698_181 , 
    RI21a0dd98_125 , 
    RI21a0afa8_153 , 
    RI210d2ef0_215 , 
    RI210cea08_243 , 
    RI210d7cc0_185 , 
    RI210cfc50_238 , 
    RI210d3760_214 , 
    RI210cf278_242 , 
    RI210ce8a0_246 , 
    RI21a0d528_129 , 
    RI210d23b0_222 , 
    RI21a0a558_161 , 
    RI210d6a00_191 , 
    RI21a0d2d0_134 , 
    RI21a0a648_159 , 
    RI210d72e8_189 , 
    RI210d24a0_220 , 
    RI21a0d3c0_132 , 
    RI210ce030_247 , 
    RI21a0adc8_157 , 
    RI21a0d4b0_130 , 
    RI210d2e78_216 , 
    RI21a0a5d0_160 , 
    RI210d7270_190 , 
    RI21a0d348_133 , 
    RI210d2428_221 , 
    RI210ce990_244 , 
    RI210d7c48_186 , 
    RI210d2e00_217 , 
    RI210cf3e0_239 , 
    RI210d2518_219 , 
    RI210ce918_245 , 
    RI210d7360_188 , 
    RI210cf368_240 , 
    RI21a09e50_162 , 
    RI210d1b40_223 , 
    RI21a0cbc8_135 , 
    RI210d6988_192 , 
    RI21a09dd8_163 , 
    RI210d6910_193 , 
    RI21a0cb50_136 , 
    RI210d1ac8_224 , 
    RI21a09478_164 , 
    RI210d6898_194 , 
    RI210d1a50_225 , 
    RI21a0cad8_137 , 
    RI210d2d88_218 , 
    RI21a0d438_131 , 
    RI21a0a6c0_158 , 
    RI210d73d8_187 , 
    RI210d10f0_228 , 
    RI210d5ec0_198 , 
    RI210da498_168 , 
    RI21a0c268_141 , 
    RI210d5fb0_196 , 
    RI210dad80_166 , 
    RI210d1168_227 , 
    RI21a0c9e8_139 , 
    RI210d5f38_197 , 
    RI210da510_167 , 
    RI21a0c970_140 , 
    RI210da420_169 , 
    RI210d5650_199 , 
    RI21a0c1f0_142 , 
    RI210d6028_195 , 
    RI210dadf8_165 , 
    RI21a0ca60_138 , 
    RI210d19d8_226 , 
    RI210da3a8_170 , 
    RI210d55d8_200 , 
    RI21a0c178_143 , 
    RI210cdfb8_248 , 
    RI21a0e590_122 , 
    RI21a0b7a0_150 , 
    RI210d8ff8_178 , 
    RI210cfd40_236 , 
    RI21a16a38_35 , 
    RI21a115d8_89 , 
    RI21a11650_88 , 
    RI210ccb90_257 , 
    RI210c9b48_275 , 
    RI210cd658_251 , 
    RI210cc140_262 , 
    RI210ca430_273 , 
    RI210c9ad0_276 , 
    RI210c91e8_278 , 
    RI210c9a58_277 , 
    RI210c2078_280 , 
    RI210c9170_279 , 
    RI210c07a0_282 , 
    RI210c0818_281 , 
    RI210cd568_253 , 
    RI210cd5e0_252 , 
    RI210ccc80_255 , 
    RI210cd4f0_254 , 
    RI210ccc08_256 , 
    RI210cc2a8_259 , 
    RI210ccb18_258 , 
    RI210cc230_260 , 
    RI210cb8d0_263 , 
    RI210cb858_264 , 
    RI210cc1b8_261 , 
    RI210cb7e0_265 , 
    RI210cb768_266 , 
    RI210caef8_267 , 
    RI210cae80_268 , 
    RI210cae08_269 , 
    RI210cad90_270 , 
    RI210ca4a8_272 , 
    RI210ca520_271 , 
    RI210ca3b8_274 , 
    RI210aeb90_395 , 
    RI210b43b0_360 , 
    RI210b7f38_335 , 
    RI210b2538_374 , 
    RI210b5670_354 , 
    RI21081aa0_439 , 
    RI2107e878_458 , 
    RI210b07b0_386 , 
    RI210af478_393 , 
    RI21080d80_445 , 
    RI2107e698_462 , 
    RI210834e0_427 , 
    RI2107f3b8_456 , 
    RI21080f60_441 , 
    RI210835d0_425 , 
    RI21084458_416 , 
    RI210afdd8_390 , 
    RI21080ee8_442 , 
    RI2107e800_459 , 
    RI210b4d10_357 , 
    RI210aec08_394 , 
    RI210b25b0_373 , 
    RI210843e0_417 , 
    RI210b4428_359 , 
    RI210b08a0_384 , 
    RI210b2f88_369 , 
    RI210b5760_352 , 
    RI21084f98_414 , 
    RI210b2f10_370 , 
    RI210b0828_385 , 
    RI210b56e8_353 , 
    RI210b3078_367 , 
    RI210b1188_382 , 
    RI210b6048_350 , 
    RI21085088_412 , 
    RI210b3000_368 , 
    RI210b0918_383 , 
    RI21085010_413 , 
    RI210b57d8_351 , 
    RI21085c40_409 , 
    RI210b61b0_347 , 
    RI210b12f0_379 , 
    RI210b39d8_364 , 
    RI21085cb8_408 , 
    RI210b6a20_346 , 
    RI210b1b60_378 , 
    RI210b3a50_363 , 
    RI210b73f8_342 , 
    RI21085e20_405 , 
    RI2107f520_453 , 
    RI21081b90_437 , 
    RI210836c0_423 , 
    RI21085e98_404 , 
    RI21081c08_436 , 
    RI210b1c50_376 , 
    RI210b1200_381 , 
    RI210b38e8_366 , 
    RI210b60c0_349 , 
    RI21085100_411 , 
    RI210b6b10_344 , 
    RI21085da8_406 , 
    RI210b4338_361 , 
    RI2107f430_455 , 
    RI210b7470_341 , 
    RI21086a50_401 , 
    RI210800d8_450 , 
    RI210827c0_433 , 
    RI210b74e8_340 , 
    RI21086ac8_400 , 
    RI21082838_432 , 
    RI21080150_449 , 
    RI210802b8_446 , 
    RI210829a0_429 , 
    RI21086e10_397 , 
    RI210b7e48_337 , 
    RI210b1cc8_375 , 
    RI21082a18_428 , 
    RI210a63a0_396 , 
    RI210b7ec0_336 , 
    RI21085178_410 , 
    RI210b6138_348 , 
    RI210b1278_380 , 
    RI210b3960_365 , 
    RI210b6a98_345 , 
    RI21085d30_407 , 
    RI210b42c0_362 , 
    RI210b1bd8_377 , 
    RI210b26a0_371 , 
    RI210b4e00_355 , 
    RI210aff40_387 , 
    RI21083648_424 , 
    RI21084f20_415 , 
    RI210afe50_389 , 
    RI21080fd8_440 , 
    RI210af4f0_392 , 
    RI21080df8_444 , 
    RI2107e710_461 , 
    RI21083558_426 , 
    RI2107e788_460 , 
    RI210b4c98_358 , 
    RI210af568_391 , 
    RI21080e70_443 , 
    RI21083738_422 , 
    RI21086960_403 , 
    RI21081c80_435 , 
    RI2107f598_452 , 
    RI21084200_421 , 
    RI210869d8_402 , 
    RI21081cf8_434 , 
    RI21080060_451 , 
    RI210828b0_431 , 
    RI210801c8_448 , 
    RI21086b40_399 , 
    RI210b7560_339 , 
    RI21082928_430 , 
    RI21080240_447 , 
    RI210b7dd0_338 , 
    RI21086bb8_398 , 
    RI210b2628_372 , 
    RI210afec8_388 , 
    RI210b4d88_356 , 
    RI210b6b88_343 , 
    RI21081b18_438 , 
    RI2107f4a8_454 , 
    RI2107f340_457 , 
    RI210cdec8_250 , 
    RI210bcdf8_303 , 
    RI210bd668_302 , 
    RI21077000_517 , 
    RI21076538_518 , 
    RI21a12988_75 , 
    RI210bf468_289 , 
    RI21078ab8_504 , 
    RI21a12910_76 , 
    RI210bf3f0_290 , 
    RI21078a40_505 , 
    RI21a12898_77 , 
    RI210beb80_291 , 
    RI21077f78_506 , 
    RI210cdf40_249 , 
    RI2107db58_464 , 
    RI21069950_647 , 
    RI210699c8_646 , 
    R_61e_1dfaf3c8 , 
    R_8f7_1e09b6c8 , 
    R_714_1dfb8888 , 
    R_951_1e17ef68 , 
    R_28c_1d9fb268 , 
    R_9be_1e183888 , 
    R_9ab_1e1827a8 , 
    R_30f_1d9d04a8 , 
    R_959_1e17f468 , 
    R_b13_1e6b0908 , 
    R_519_1dda4b48 , 
    R_92d_1e09d888 , 
    R_c06_1e6bafe8 , 
    R_8c6_1e099d28 , 
    R_845_1e094788 , 
    R_414_1d9da7c8 , 
    R_313_1d9d0728 , 
    R_518_1dda4aa8 , 
    R_9d9_1e184468 , 
    R_4dd_1dda25c8 , 
    R_59f_1dda9f08 , 
    R_517_1dda4a08 , 
    R_509_1dda4148 , 
    R_508_1dda40a8 , 
    R_401_1d9d9be8 , 
    R_5f9_1ddad748 , 
    R_6ef_1dfb7168 , 
    R_a30_1e187ac8 , 
    R_2b0_1d9fc8e8 , 
    R_77c_1dfbc988 , 
    R_8f1_1e09b308 , 
    R_36a_1d9d4288 , 
    R_507_1dda4008 , 
    R_516_1dda4e68 , 
    R_98e_1e181a88 , 
    R_8d5_1e09a188 , 
    R_498_1dd9faa8 , 
    R_68b_1dfb32e8 , 
    R_773_1dfbc3e8 , 
    R_45b_1d9dd428 , 
    R_48d_1dd9f3c8 , 
    R_5ff_1ddadb08 , 
    R_705_1dfb7f28 , 
    R_644_1dfb0688 , 
    R_63a_1dfb0548 , 
    R_ac7_1e18d928 , 
    R_320_1d9d0f48 , 
    R_737_1dfb9e68 , 
    R_506_1dda4468 , 
    R_647_1dfb0868 , 
    R_b86_1e6bb4e8 , 
    R_883_1e096e48 , 
    R_6a8_1dfb4508 , 
    R_aa5_1e18c3e8 , 
    R_440_1d9dc348 , 
    R_2f9_1d9cf6e8 , 
    R_69c_1dfb3d88 , 
    R_65d_1dfb1628 , 
    R_b0c_1e6b04a8 , 
    R_b20_1e6b1128 , 
    R_a2e_1e189788 , 
    R_905_1e09bf88 , 
    R_a57_1e189328 , 
    R_5f8_1ddad6a8 , 
    R_54c_1dda6b28 , 
    R_bd2_1e6b32e8 , 
    R_aca_1e6ae068 , 
    R_58b_1dda9288 , 
    R_2e3_1d9ce928 , 
    R_3e2_1d9d8d88 , 
    R_8f6_1e09bb28 , 
    R_331_1d9d19e8 , 
    R_97d_1e180ae8 , 
    R_5cd_1ddabbc8 , 
    R_45c_1d9dd4c8 , 
    R_999_1e181c68 , 
    R_b99_1e6b5cc8 , 
    R_948_1e17e9c8 , 
    R_97e_1e181308 , 
    R_ab0_1e18cac8 , 
    R_bb8_1e6b7028 , 
    R_489_1dd9f148 , 
    R_4b6_1dda1268 , 
    R_63f_1dfb0368 , 
    R_3e7_1d9d8ba8 , 
    R_2bd_1d9fd108 , 
    R_81b_1e092d48 , 
    R_b54_1e6b31a8 , 
    R_4df_1dda2708 , 
    R_bab_1e6b6808 , 
    R_431_1d9db9e8 , 
    R_2f2_1d9cf788 , 
    R_601_1ddadc48 , 
    R_6e7_1dfb6c68 , 
    R_bdf_1e6b8888 , 
    R_656_1dfb1bc8 , 
    R_4e0_1dda27a8 , 
    R_4de_1dda2b68 , 
    R_a4e_1e189288 , 
    R_8e1_1e09a908 , 
    R_8f0_1e09b268 , 
    R_299_1d9fba88 , 
    R_292_1d9fb628 , 
    R_4e1_1dda2848 , 
    R_a7f_1e18ac28 , 
    R_c04_1e6b9fa8 , 
    R_3ef_1d9d90a8 , 
    R_5de_1dd9f1e8 , 
    R_878_1e096768 , 
    R_720_1dfb9008 , 
    R_ad6_1e6ae7e8 , 
    R_9a2_1e182708 , 
    R_630_1dfafa08 , 
    R_52f_1dda5908 , 
    R_7a9_1e08e608 , 
    R_976_1e180b88 , 
    R_439_1d9dbee8 , 
    R_604_1ddade28 , 
    R_530_1dda59a8 , 
    R_52e_1dda5d68 , 
    R_7ed_1e091088 , 
    R_3f2_1d9d4c88 , 
    R_3d4_1d9d7fc8 , 
    R_84a_1e094fa8 , 
    R_2de_1d9ceb08 , 
    R_690_1dfb3608 , 
    R_4cd_1dda1bc8 , 
    R_531_1dda5a48 , 
    R_b34_1e6b1da8 , 
    R_5f7_1ddad608 , 
    R_806_1e092528 , 
    R_a5b_1e1895a8 , 
    R_718_1dfb8b08 , 
    R_695_1dfb3928 , 
    R_7af_1e08e9c8 , 
    R_62b_1dfaf6e8 , 
    R_904_1e09bee8 , 
    R_501_1dda3c48 , 
    R_585_1dda8ec8 , 
    R_9cd_1e183ce8 , 
    R_78c_1dfbd388 , 
    R_392_1d9d5b88 , 
    R_4b4_1dda0c28 , 
    R_b44_1e6b27a8 , 
    R_969_1e17fe68 , 
    R_40d_1d9da368 , 
    R_627_1dfaf468 , 
    R_67a_1dfadfc8 , 
    R_45d_1d9dd568 , 
    R_7c1_1e08f508 , 
    R_552_1dda73e8 , 
    R_2bf_1d9fd248 , 
    R_5d4_1ddac028 , 
    R_b77_1e6b4788 , 
    R_3fa_1d9db088 , 
    R_6aa_1dfb4b48 , 
    R_82a_1e093ba8 , 
    R_3aa_1d9d6a88 , 
    R_300_1d9cfb48 , 
    R_405_1d9d9e68 , 
    R_953_1e17f0a8 , 
    R_3cf_1d9d7ca8 , 
    R_ac1_1e18d568 , 
    R_61c_1dfaed88 , 
    R_a99_1e18bc68 , 
    R_4ae_1dda0fe8 , 
    R_aec_1e6af0a8 , 
    R_af8_1e6af828 , 
    R_762_1dfbbe48 , 
    R_3a8_1d9d6448 , 
    R_4ca_1dda1ee8 , 
    R_6b7_1dfb4e68 , 
    R_57c_1dda8928 , 
    R_52b_1dda5688 , 
    R_8ef_1e09b1c8 , 
    R_8c5_1e099788 , 
    R_8ab_1e098748 , 
    R_71c_1dfb8d88 , 
    R_388_1d9d5048 , 
    R_b6e_1e6b46e8 , 
    R_9cc_1e183c48 , 
    R_65b_1dfb14e8 , 
    R_bbd_1e6b7348 , 
    R_3b2_1d9d6f88 , 
    R_862_1e095ea8 , 
    R_4a5_1dda02c8 , 
    R_90f_1e09c5c8 , 
    R_702_1dfb8248 , 
    R_29f_1d9fbe48 , 
    R_72b_1dfb96e8 , 
    R_6f4_1dfb7488 , 
    R_5f2_1dda8a68 , 
    R_a64_1e189b48 , 
    R_2e9_1d9cece8 , 
    R_683_1dfb2de8 , 
    R_2fd_1d9cf968 , 
    R_8b2_1e0990a8 , 
    R_5f0_1ddad1a8 , 
    R_bac_1e6b68a8 , 
    R_642_1dfb0a48 , 
    R_5f6_1d9fbda8 , 
    R_568_1dda7ca8 , 
    R_409_1d9da0e8 , 
    R_5a8_1ddaa4a8 , 
    R_5e3_1ddac988 , 
    R_96b_1e17ffa8 , 
    R_bca_1e6b14e8 , 
    R_3b8_1d9d6e48 , 
    R_789_1dfbd1a8 , 
    R_86a_1e0963a8 , 
    R_416_1ddabc68 , 
    R_903_1e09be48 , 
    R_a2d_1e1878e8 , 
    R_9cb_1e183ba8 , 
    R_59b_1dda9c88 , 
    R_a4c_1e188c48 , 
    R_79c_1dfbdd88 , 
    R_888_1e097168 , 
    R_2a7_1d9fc348 , 
    R_7f3_1e091448 , 
    R_73c_1dfba188 , 
    R_bd1_1e6b7fc8 , 
    R_4a6_1dda0868 , 
    R_3dd_1d9d8568 , 
    R_346_1d9d2c08 , 
    R_4c4_1dda1628 , 
    R_b15_1e6b0a48 , 
    R_5ec_1ddacf28 , 
    R_bb4_1e6b6da8 , 
    R_bed_1e6b9148 , 
    R_7bf_1e08f3c8 , 
    R_344_1d9d25c8 , 
    R_c0b_1e6ba408 , 
    R_6a5_1dfb4328 , 
    R_b8c_1e6b54a8 , 
    R_3a1_1d9d5fe8 , 
    R_7ea_1e09d928 , 
    R_46e_1dd9e568 , 
    R_8ee_1e09b628 , 
    R_697_1dfb3a68 , 
    R_77f_1dfbcb68 , 
    R_391_1d9d55e8 , 
    R_746_1dfb6448 , 
    R_b3b_1e6b2208 , 
    R_7f1_1e091308 , 
    R_410_1d9da548 , 
    R_700_1dfb7c08 , 
    R_58f_1dda9508 , 
    R_582_1dda91e8 , 
    R_793_1dfbd7e8 , 
    R_847_1e0948c8 , 
    R_95e_1e17fc88 , 
    R_560_1dda77a8 , 
    R_9ca_1e184008 , 
    R_397_1d9d59a8 , 
    R_46b_1d9dde28 , 
    R_44e_1d9fc028 , 
    R_6cc_1dfb5b88 , 
    R_62e_1dfafdc8 , 
    R_2b1_1d9fc988 , 
    R_6f9_1dfb77a8 , 
    R_af5_1e6af648 , 
    R_b81_1e6b4dc8 , 
    R_427_1d9db3a8 , 
    R_547_1dda6808 , 
    R_c1d_1e6baf48 , 
    R_a2c_1e187848 , 
    R_355_1d9d3068 , 
    R_857_1e0952c8 , 
    R_413_1d9da728 , 
    R_afa_1e6afe68 , 
    R_adc_1e6ae6a8 , 
    R_5fc_1ddad928 , 
    R_c24_1e6bb3a8 , 
    R_421_1d9dafe8 , 
    R_892_1e17e608 , 
    R_70b_1dfb82e8 , 
    R_aad_1e18c8e8 , 
    R_3ca_1d9d8108 , 
    R_7ac_1e08e7e8 , 
    R_8da_1e09a9a8 , 
    R_400_1d9d9b48 , 
    R_bb0_1e6b6b28 , 
    R_893_1e097848 , 
    R_902_1e09c2a8 , 
    R_a93_1e18b8a8 , 
    R_8cd_1e099c88 , 
    R_861_1e095908 , 
    R_3ea_1d9d9288 , 
    R_915_1e09c988 , 
    R_844_1e0946e8 , 
    R_677_1dfb2668 , 
    R_602_1dfae248 , 
    R_39c_1d9d5cc8 , 
    R_be3_1e6b8b08 , 
    R_bea_1e6b9468 , 
    R_993_1e1818a8 , 
    R_bad_1e6b6948 , 
    R_88d_1e097488 , 
    R_5a2_1ddaa5e8 , 
    R_655_1dfb1128 , 
    R_4ad_1dda07c8 , 
    R_493_1dd9f788 , 
    R_894_1e0978e8 , 
    R_668_1dfb1d08 , 
    R_730_1dfb9a08 , 
    R_7dc_1e0905e8 , 
    R_abd_1e18d2e8 , 
    R_662_1dfb1e48 , 
    R_a7c_1e18aa48 , 
    R_5cf_1ddabd08 , 
    R_328_1d9d1448 , 
    R_741_1dfba4a8 , 
    R_9a6_1e182988 , 
    R_36d_1d9d3f68 , 
    R_308_1d9d0048 , 
    R_95b_1e17f5a8 , 
    R_b63_1e6b3b08 , 
    R_2da_1d9ce888 , 
    R_5dc_1ddac528 , 
    R_49f_1dd9ff08 , 
    R_895_1e097988 , 
    R_761_1dfbb8a8 , 
    R_2e4_1d9ce9c8 , 
    R_ab5_1e18cde8 , 
    R_c28_1e6bb628 , 
    R_8d4_1e09a0e8 , 
    R_a8c_1e18b448 , 
    R_597_1dda9a08 , 
    R_5c4_1ddab628 , 
    R_384_1d9d4dc8 , 
    R_31c_1d9d0cc8 , 
    R_987_1e181128 , 
    R_b2e_1e6b1ee8 , 
    R_2f3_1d9cf328 , 
    R_6cf_1dfb5d68 , 
    R_6e4_1dfb6a88 , 
    R_357_1d9d31a8 , 
    R_3c1_1d9d73e8 , 
    R_5e7_1ddacc08 , 
    R_974_1e180548 , 
    R_61a_1dfaf148 , 
    R_3f8_1d9d9648 , 
    R_802_1e0922a8 , 
    R_593_1dda9788 , 
    R_a69_1e189e68 , 
    R_a87_1e18b128 , 
    R_a5d_1e1896e8 , 
    R_a2b_1e1877a8 , 
    R_671_1dfb22a8 , 
    R_4cf_1dda1d08 , 
    R_420_1d9daf48 , 
    R_6bc_1dfb5188 , 
    R_43f_1d9dc2a8 , 
    R_692_1dfb3c48 , 
    R_80b_1e092348 , 
    R_882_1e0972a8 , 
    R_871_1e096308 , 
    R_2c2_1d9fd928 , 
    R_2ce_1d9cfa08 , 
    R_a9c_1e18be48 , 
    R_768_1dfbbd08 , 
    R_56d_1dda7fc8 , 
    R_34c_1d9d2ac8 , 
    R_b8f_1e6b5688 , 
    R_b07_1e6b0188 , 
    R_6b5_1dfb4d28 , 
    R_5ae_1ddaad68 , 
    R_2df_1d9ce6a8 , 
    R_674_1dfb2488 , 
    R_608_1dfae108 , 
    R_ad3_1e6ae108 , 
    R_505_1dda3ec8 , 
    R_8bf_1e0993c8 , 
    R_542_1dda69e8 , 
    R_7f6_1e091b28 , 
    R_504_1dda3e28 , 
    R_8a7_1e0984c8 , 
    R_76a_1dfbc5c8 , 
    R_937_1e09dec8 , 
    R_6fb_1dfb78e8 , 
    R_3b0_1d9d6948 , 
    R_2c0_1d9fd2e8 , 
    R_37c_1d9d48c8 , 
    R_782_1dfbd248 , 
    R_503_1dda3d88 , 
    R_82e_1e093e28 , 
    R_8bb_1e099148 , 
    R_430_1d9db948 , 
    R_5cb_1ddaba88 , 
    R_ae6_1e6af1e8 , 
    R_7a3_1e08e248 , 
    R_b78_1e6b4828 , 
    R_bc9_1e6b7ac8 , 
    R_380_1d9d4b48 , 
    R_33d_1d9d2168 , 
    R_8e0_1e09a868 , 
    R_3c7_1d9d77a8 , 
    R_2b2_1d9fcf28 , 
    R_618_1dfaeb08 , 
    R_823_1e093248 , 
    R_89e_1e098428 , 
    R_502_1dda41e8 , 
    R_b6f_1e6b4288 , 
    R_c00_1e6b9d28 , 
    R_98d_1e1814e8 , 
    R_28b_1d9fb1c8 , 
    R_a55_1e1891e8 , 
    R_3c4_1d9d75c8 , 
    R_40c_1d9da2c8 , 
    R_2d2_1d9ce388 , 
    R_c21_1e6bb1c8 , 
    R_b3d_1e6b2348 , 
    R_877_1e0966c8 , 
    R_855_1e095188 , 
    R_41d_1d9dad68 , 
    R_438_1d9dbe48 , 
    R_2d6_1d9ce608 , 
    R_7da_1e0909a8 , 
    R_6f6_1dfb7ac8 , 
    R_9aa_1e182e88 , 
    R_b47_1e6b2988 , 
    R_a2a_1e6b3ce8 , 
    R_41f_1d9daea8 , 
    R_ae4_1e6aeba8 , 
    R_a79_1e18a868 , 
    R_3a3_1d9d6128 , 
    R_5bd_1ddab1c8 , 
    R_301_1d9cfbe8 , 
    R_298_1d9fb9e8 , 
    R_bb9_1e6b70c8 , 
    R_82d_1e093888 , 
    R_404_1d9d9dc8 , 
    R_a62_1e189f08 , 
    R_93c_1e17e248 , 
    R_62d_1dfaf828 , 
    R_579_1dda8748 , 
    R_452_1ddac3e8 , 
    R_54d_1dda6bc8 , 
    R_4d9_1dda2348 , 
    R_4d4_1dda2028 , 
    R_6c1_1dfb54a8 , 
    R_379_1d9d46e8 , 
    R_34e_1d9d3108 , 
    R_94a_1e097ca8 , 
    R_74b_1dfbaae8 , 
    R_ade_1e6aece8 , 
    R_79f_1e08dfc8 , 
    R_797_1dfbda68 , 
    R_943_1e17e6a8 , 
    R_653_1dfb0fe8 , 
    R_3d8_1d9d8248 , 
    R_b61_1e6b39c8 , 
    R_bc4_1e6b77a8 , 
    R_a02_1e186308 , 
    R_368_1d9d3c48 , 
    R_35e_1d9d3b08 , 
    R_7fe_1e092028 , 
    R_499_1dd9fb48 , 
    R_680_1dfb2c08 , 
    R_2a8_1d9fc3e8 , 
    R_6ec_1dfb6f88 , 
    R_776_1dfbcac8 , 
    R_b5e_1e6b0368 , 
    R_635_1dfafd28 , 
    R_7fa_1e091da8 , 
    R_af7_1e6af788 , 
    R_8c4_1e0996e8 , 
    R_408_1d9da048 , 
    R_ab9_1e18d068 , 
    R_6a2_1dfb61c8 , 
    R_291_1d9fb588 , 
    R_7b8_1e08ef68 , 
    R_8b6_1e08e6a8 , 
    R_48a_1dda0d68 , 
    R_6c7_1dfb5868 , 
    R_c10_1e6ba728 , 
    R_bf1_1e6b93c8 , 
    R_4d6_1dd9e2e8 , 
    R_5b3_1ddaab88 , 
    R_771_1dfbc2a8 , 
    R_af1_1e6af3c8 , 
    R_6e1_1dfb68a8 , 
    R_a9f_1e18c028 , 
    R_b17_1e6b0b88 , 
    R_b30_1e6b1b28 , 
    R_bde_1e6b37e8 , 
    R_998_1e181bc8 , 
    R_a4a_1e189008 , 
    R_48e_1dd9f968 , 
    R_688_1dfb3108 , 
    R_810_1e092668 , 
    R_75c_1dfbb588 , 
    R_3bb_1d9d7028 , 
    R_c2e_1e17f008 , 
    R_5d2_1d9db308 , 
    R_32e_1d9d1d08 , 
    R_580_1dda8ba8 , 
    R_453_1d9dcf28 , 
    R_83a_1e0913a8 , 
    R_41e_1d9dc988 , 
    R_97c_1e180a48 , 
    R_5b8_1ddaaea8 , 
    R_363_1d9d3928 , 
    R_94e_1ddadce8 , 
    R_7c4_1e08f6e8 , 
    R_52c_1dda5728 , 
    R_aa2_1e18c708 , 
    R_625_1dfaf328 , 
    R_4b7_1dda0e08 , 
    R_55d_1dda75c8 , 
    R_b0e_1e6b0ae8 , 
    R_425_1d9db268 , 
    R_30c_1d9d02c8 , 
    R_3db_1d9d8428 , 
    R_a48_1e1889c8 , 
    R_aaf_1e18ca28 , 
    R_5ad_1ddaa7c8 , 
    R_589_1dda9148 , 
    R_338_1d9d1e48 , 
    R_832_1e0940a8 , 
    R_790_1dfbd608 , 
    R_318_1d9d0a48 , 
    R_869_1e095e08 , 
    R_6d3_1dfb5fe8 , 
    R_60c_1dfae388 , 
    R_56a_1dda82e8 , 
    R_887_1e0970c8 , 
    R_815_1e092988 , 
    R_66b_1dfb1ee8 , 
    R_a34_1e187d48 , 
    R_40f_1d9da4a8 , 
    R_ac3_1e18d6a8 , 
    R_324_1d9d11c8 , 
    R_614_1dfae888 , 
    R_752_1dfbb448 , 
    R_4c0_1dda13a8 , 
    R_7d9_1e090408 , 
    R_ad0_1e18dec8 , 
    R_bee_1e6b96e8 , 
    R_736_1dfba2c8 , 
    R_727_1dfb9468 , 
    R_a8a_1e18b808 , 
    R_933_1e09dc48 , 
    R_8b1_1e098b08 , 
    R_606_1dfae4c8 , 
    R_927_1e09d4c8 , 
    R_a7a_1e18ae08 , 
    R_333_1d9d1b28 , 
    R_968_1e17fdc8 , 
    R_574_1dda8428 , 
    R_836_1e094328 , 
    R_757_1dfbb268 , 
    R_2db_1d9ce428 , 
    R_af4_1e6af5a8 , 
    R_454_1d9dcfc8 , 
    R_412_1d9dab88 , 
    R_709_1dfb81a8 , 
    R_8a4_1e0982e8 , 
    R_c1b_1e6bae08 , 
    R_846_1e094d28 , 
    R_3ff_1d9d9aa8 , 
    R_76e_1dfbdec8 , 
    R_33f_1d9d22a8 , 
    R_4af_1dda0908 , 
    R_a67_1e189d28 , 
    R_616_1dfaeec8 , 
    R_b49_1e6b2ac8 , 
    R_2f4_1d9cf3c8 , 
    R_426_1d9db808 , 
    R_2e5_1d9cea68 , 
    R_bb5_1e6b6e48 , 
    R_7b6_1e08f328 , 
    R_751_1dfbaea8 , 
    R_bd0_1e6b7f28 , 
    R_610_1dfae608 , 
    R_918_1e09cb68 , 
    R_35c_1d9d34c8 , 
    R_924_1e09d2e8 , 
    R_912_1e09cca8 , 
    R_77d_1dfbca28 , 
    R_774_1dfbc488 , 
    R_a71_1e18a368 , 
    R_32d_1d9d1768 , 
    R_99d_1e181ee8 , 
    R_87d_1e096a88 , 
    R_472_1dd9e7e8 , 
    R_b2a_1e6b1c68 , 
    R_56f_1dda8108 , 
    R_b87_1e6b5188 , 
    R_921_1e09d108 , 
    R_375_1d9d4468 , 
    R_576_1dda8ce8 , 
    R_b82_1e6b5368 , 
    R_39e_1d9d6308 , 
    R_856_1e095728 , 
    R_6c2_1dfb5a48 , 
    R_2c3_1d9fd4c8 , 
    R_90b_1e09c348 , 
    R_92f_1e09d9c8 , 
    R_38e_1d9d5908 , 
    R_b9e_1e18d388 , 
    R_8cc_1e099be8 , 
    R_860_1e095868 , 
    R_c09_1e6ba2c8 , 
    R_b09_1e6b02c8 , 
    R_521_1dda5048 , 
    R_b4a_1e6b3068 , 
    R_88c_1e0973e8 , 
    R_520_1dda4fa8 , 
    R_8b5_1e098d88 , 
    R_b5d_1e6b3748 , 
    R_843_1e094648 , 
    R_633_1dfafbe8 , 
    R_7c2_1e08faa8 , 
    R_6d8_1dfb6308 , 
    R_38d_1d9d5368 , 
    R_7e7_1e090cc8 , 
    R_bfc_1e6b9aa8 , 
    R_841_1e094508 , 
    R_a96_1e18bf88 , 
    R_7e5_1e090b88 , 
    R_51f_1dda4f08 , 
    R_949_1e17ea68 , 
    R_b5a_1e6b3a68 , 
    R_2e0_1d9ce748 , 
    R_acd_1e18dce8 , 
    R_70f_1dfb8568 , 
    R_c15_1e6baa48 , 
    R_310_1d9d0548 , 
    R_bf5_1e6b9648 , 
    R_314_1d9d07c8 , 
    R_6af_1dfb4968 , 
    R_445_1d9dc668 , 
    R_658_1dfb1308 , 
    R_a6c_1e18a048 , 
    R_2c1_1d9fd388 , 
    R_2b3_1d9fcac8 , 
    R_6de_1dfb6bc8 , 
    R_9b9_1e183068 , 
    R_6ad_1dfb4828 , 
    R_548_1dda68a8 , 
    R_4c9_1dda1948 , 
    R_51e_1dda5368 , 
    R_96a_1e180408 , 
    R_455_1d9dd068 , 
    R_8d3_1e09a048 , 
    R_bb1_1e6b6bc8 , 
    R_7d7_1e0902c8 , 
    R_6a0_1dfb4008 , 
    R_b79_1e6b48c8 , 
    R_565_1dda7ac8 , 
    R_586_1dda9468 , 
    R_4a7_1dda0408 , 
    R_b70_1e6b4328 , 
    R_661_1dfb18a8 , 
    R_2d3_1d9fdec8 , 
    R_ad9_1e6ae4c8 , 
    R_a85_1e18afe8 , 
    R_a77_1e18a728 , 
    R_2d7_1d9ce1a8 , 
    R_7b3_1e08ec48 , 
    R_870_1e096268 , 
    R_43e_1d9dc708 , 
    R_6db_1dfb64e8 , 
    R_807_1e0920c8 , 
    R_a74_1e18a548 , 
    R_bf9_1e6b98c8 , 
    R_321_1d9d0fe8 , 
    R_a53_1e1890a8 , 
    R_4e3_1dda2988 , 
    R_831_1e093b08 , 
    R_66e_1dfb25c8 , 
    R_ac6_1e18dd88 , 
    R_55a_1dda78e8 , 
    R_4c6_1dda1c68 , 
    R_4e4_1dda2a28 , 
    R_4e2_1dda2de8 , 
    R_c22_1e6b55e8 , 
    R_92c_1e09d7e8 , 
    R_7c9_1e08fa08 , 
    R_623_1dfaf1e8 , 
    R_b58_1e6b3428 , 
    R_370_1d9d4148 , 
    R_3be_1d9d7708 , 
    R_4e5_1dda2ac8 , 
    R_a03_1e185ea8 , 
    R_c12_1e6bad68 , 
    R_456_1d9dd608 , 
    R_bf2_1e6b9968 , 
    R_6a7_1dfb4468 , 
    R_c30_1e6bbb28 , 
    R_40b_1d9da228 , 
    R_42f_1d9db8a8 , 
    R_68d_1dfb3428 , 
    R_735_1dfb9d28 , 
    R_78d_1dfbd428 , 
    R_8df_1e09a7c8 , 
    R_41c_1d9dacc8 , 
    R_46f_1dd9e108 , 
    R_2a9_1d9fc488 , 
    R_81e_1e093428 , 
    R_5e0_1ddac7a8 , 
    R_462_1d9ddd88 , 
    R_60a_1dfae748 , 
    R_5a7_1ddaa408 , 
    R_403_1d9d9d28 , 
    R_2c6_1d9fdba8 , 
    R_7e3_1e090a48 , 
    R_7ee_1e09c528 , 
    R_706_1dfb84c8 , 
    R_c17_1e6bab88 , 
    R_c1f_1e6bb088 , 
    R_b93_1e6b5908 , 
    R_854_1e0950e8 , 
    R_b9f_1e6b6088 , 
    R_8e5_1e09ab88 , 
    R_437_1d9dbda8 , 
    R_612_1dfaec48 , 
    R_816_1e0931a8 , 
    R_b19_1e6b0cc8 , 
    R_73b_1dfba0e8 , 
    R_a44_1e188748 , 
    R_93e_1e17e888 , 
    R_67c_1dfb2988 , 
    R_992_1e181d08 , 
    R_494_1dd9f828 , 
    R_3e0_1d9d8748 , 
    R_7a7_1e08e4c8 , 
    R_876_1e096b28 , 
    R_543_1dda6588 , 
    R_8ae_1dfbc0c8 , 
    R_351_1d9d2de8 , 
    R_457_1d9dd1a8 , 
    R_bf6_1e6b3f68 , 
    R_a38_1e187fc8 , 
    R_6f1_1dfb72a8 , 
    R_b3e_1e6b28e8 , 
    R_53e_1dda6768 , 
    R_ac0_1e18d4c8 , 
    R_763_1dfbb9e8 , 
    R_c26_1e6b8ce8 , 
    R_650_1dfb0e08 , 
    R_361_1d9d37e8 , 
    R_aaa_1e187e88 , 
    R_b10_1e6b0728 , 
    R_b2c_1e6b18a8 , 
    R_5a1_1ddaa048 , 
    R_be7_1e6b8d88 , 
    R_b26_1e6b19e8 , 
    R_4a0_1dd9ffa8 , 
    R_95a_1e17fa08 , 
    R_909_1e09c208 , 
    R_463_1d9dd928 , 
    R_407_1d9d9fa8 , 
    R_5c5_1ddab6c8 , 
    R_986_1e181588 , 
    R_515_1dda48c8 , 
    R_5c1_1ddab448 , 
    R_297_1d9fb948 , 
    R_514_1dda4828 , 
    R_b4c_1e6b2ca8 , 
    R_973_1e1804a8 , 
    R_60e_1dfae9c8 , 
    R_7d4_1e0900e8 , 
    R_7c7_1e08f8c8 , 
    R_513_1dda4788 , 
    R_65f_1dfb1768 , 
    R_9b5_1e182de8 , 
    R_2ee_1d9cf508 , 
    R_91b_1e09cd48 , 
    R_af6_1e6afbe8 , 
    R_83d_1e094288 , 
    R_8c3_1e099648 , 
    R_458_1d9dd248 , 
    R_512_1dda4be8 , 
    R_ba6_1e6b69e8 , 
    R_5e5_1ddacac8 , 
    R_57b_1dda8888 , 
    R_aeb_1e6af008 , 
    R_7f4_1e0914e8 , 
    R_a46_1e188d88 , 
    R_b8d_1e6b5548 , 
    R_562_1dda7de8 , 
    R_745_1dfba728 , 
    R_557_1dda7208 , 
    R_464_1d9dd9c8 , 
    R_835_1e093d88 , 
    R_49a_1dda00e8 , 
    R_7d1_1e08ff08 , 
    R_911_1e09c708 , 
    R_6e9_1dfb6da8 , 
    R_723_1dfb91e8 , 
    R_a95_1e18b9e8 , 
    R_58d_1dda93c8 , 
    R_a89_1e18b268 , 
    R_780_1dfbcc08 , 
    R_740_1dfba408 , 
    R_72f_1dfb9968 , 
    R_828_1e093568 , 
    R_89c_1e097de8 , 
    R_a32_1e188108 , 
    R_840_1e094468 , 
    R_b37_1e6b1f88 , 
    R_9db_1e1845a8 , 
    R_b22_1e6b1768 , 
    R_9dc_1e184648 , 
    R_9da_1e184a08 , 
    R_794_1dfbd888 , 
    R_33a_1d9d2488 , 
    R_424_1d9db1c8 , 
    R_2dc_1d9ce4c8 , 
    R_a6f_1e18a228 , 
    R_98c_1e181448 , 
    R_6b6_1dfb52c8 , 
    R_908_1e09c168 , 
    R_9dd_1e1846e8 , 
    R_965_1e17fbe8 , 
    R_28a_1d9fb128 , 
    R_529_1dda5548 , 
    R_40e_1d9da908 , 
    R_bcd_1e6b7d48 , 
    R_476_1dd9ea68 , 
    R_393_1d9d5728 , 
    R_a40_1e1884c8 , 
    R_528_1dda54a8 , 
    R_2fa_1d9d0188 , 
    R_a3c_1e188248 , 
    R_868_1e095d68 , 
    R_2cf_1d9fdc48 , 
    R_2c4_1d9fd568 , 
    R_7cc_1e08fbe8 , 
    R_8fd_1e09ba88 , 
    R_3d5_1d9d8068 , 
    R_b64_1e6b3ba8 , 
    R_527_1dda5408 , 
    R_9d1_1e183f68 , 
    R_46c_1d9ddec8 , 
    R_2f5_1d9cf468 , 
    R_839_1e094008 , 
    R_554_1dda7028 , 
    R_3ab_1d9d6628 , 
    R_459_1d9dd2e8 , 
    R_b4f_1e6b2e88 , 
    R_886_1e097528 , 
    R_3e5_1d9d8a68 , 
    R_52d_1dda57c8 , 
    R_290_1d9fb4e8 , 
    R_b7a_1e18cc08 , 
    R_526_1dda5ae8 , 
    R_79a_1e098e28 , 
    R_ba0_1e6b6128 , 
    R_6d1_1dfb5ea8 , 
    R_713_1dfb87e8 , 
    R_685_1dfb2f28 , 
    R_3fe_1d9d9f08 , 
    R_638_1dfaff08 , 
    R_465_1d9dda68 , 
    R_b91_1e6b57c8 , 
    R_b53_1e6b3108 , 
    R_8ad_1e098888 , 
    R_59e_1dd9e068 , 
    R_9c5_1e1837e8 , 
    R_3a9_1d9d64e8 , 
    R_3b3_1d9d6b28 , 
    R_2b4_1d9fcb68 , 
    R_af3_1e6af508 , 
    R_4f9_1dda3748 , 
    R_a90_1e18b6c8 , 
    R_389_1d9d50e8 , 
    R_a6a_1e18a408 , 
    R_b1b_1e6b0e08 , 
    R_4f8_1dda36a8 , 
    R_b66_1e6b9be8 , 
    R_9d0_1e183ec8 , 
    R_2e1_1d9ce7e8 , 
    R_7d2_1e0904a8 , 
    R_803_1e091e48 , 
    R_91e_1e09d428 , 
    R_4f7_1dda3608 , 
    R_ab4_1e18cd48 , 
    R_6ee_1dfb75c8 , 
    R_c05_1e6ba048 , 
    R_704_1dfb7e88 , 
    R_353_1d9d2f28 , 
    R_ba7_1e6b6588 , 
    R_87c_1e0969e8 , 
    R_3f5_1d9d9468 , 
    R_abc_1e18d248 , 
    R_a83_1e18aea8 , 
    R_b40_1e6b2528 , 
    R_a06_1e186588 , 
    R_907_1e09c0c8 , 
    R_664_1dfb1a88 , 
    R_b71_1e6b43c8 , 
    R_4f6_1ddad2e8 , 
    R_8b9_1e099008 , 
    R_971_1e180368 , 
    R_64e_1dfb11c8 , 
    R_679_1dfb27a8 , 
    R_80c_1e0923e8 , 
    R_347_1d9d27a8 , 
    R_b28_1e6b1628 , 
    R_7cf_1e08fdc8 , 
    R_8fc_1e09b9e8 , 
    R_72d_1dfb9828 , 
    R_9c4_1e183748 , 
    R_997_1e181b28 , 
    R_85f_1e0957c8 , 
    R_2d4_1d9cdfc8 , 
    R_48f_1dd9f508 , 
    R_adb_1e6ae608 , 
    R_3b9_1d9d6ee8 , 
    R_a51_1e188f68 , 
    R_8cb_1e099b48 , 
    R_2d8_1d9ce248 , 
    R_a72_1e18a908 , 
    R_7f7_1e0916c8 , 
    R_4b5_1dda0cc8 , 
    R_88b_1e097348 , 
    R_aa7_1e18c528 , 
    R_699_1dfb3ba8 , 
    R_68a_1dfb3748 , 
    R_9cf_1e183e28 , 
    R_345_1d9d2668 , 
    R_76b_1dfbbee8 , 
    R_7aa_1e099328 , 
    R_5e9_1ddacd48 , 
    R_a04_1e185f48 , 
    R_36b_1d9d3e28 , 
    R_444_1d9dc5c8 , 
    R_842_1e094aa8 , 
    R_58a_1dda96e8 , 
    R_97b_1e1809a8 , 
    R_5bc_1ddab128 , 
    R_ae9_1e6aeec8 , 
    R_74e_1dfbc348 , 
    R_69b_1dfb3ce8 , 
    R_783_1dfbcde8 , 
    R_64d_1dfb0c28 , 
    R_938_1e17dfc8 , 
    R_7bd_1e08f288 , 
    R_7ca_1e08ffa8 , 
    R_482_1ddac668 , 
    R_2c7_1d9fd748 , 
    R_621_1dfaf0a8 , 
    R_9c3_1e1836a8 , 
    R_309_1d9d00e8 , 
    R_5f1_1ddad248 , 
    R_4b8_1dda0ea8 , 
    R_bcf_1e6b7e88 , 
    R_824_1e0932e8 , 
    R_6e6_1dfb70c8 , 
    R_7a4_1e08e2e8 , 
    R_59d_1dda9dc8 , 
    R_769_1dfbbda8 , 
    R_38a_1d9d5688 , 
    R_4cb_1dda1a88 , 
    R_8d9_1e09a408 , 
    R_8d2_1e09a4a8 , 
    R_b24_1e6b13a8 , 
    R_4ba_1d9d9a08 , 
    R_bdd_1e6b8748 , 
    R_398_1d9d5a48 , 
    R_31d_1d9d0d68 , 
    R_47a_1dd9ece8 , 
    R_2ca_1d9ce108 , 
    R_b03_1e6aff08 , 
    R_2a0_1d9fbee8 , 
    R_71f_1dfb8f68 , 
    R_950_1e17eec8 , 
    R_9ce_1e184288 , 
    R_aae_1e6b6c68 , 
    R_b39_1e6b20c8 , 
    R_906_1e090ea8 , 
    R_786_1dfbd4c8 , 
    R_81c_1e092de8 , 
    R_94b_1e17eba8 , 
    R_8fb_1e09b948 , 
    R_3cb_1d9d7a28 , 
    R_86f_1e0961c8 , 
    R_584_1dda8e28 , 
    R_40a_1d9da688 , 
    R_954_1e17f148 , 
    R_944_1e17e748 , 
    R_bc8_1e6b7a28 , 
    R_9a1_1e182168 , 
    R_c02_1e6ba5e8 , 
    R_967_1e17fd28 , 
    R_7ff_1e091bc8 , 
    R_329_1d9d14e8 , 
    R_ba1_1e6b61c8 , 
    R_717_1dfb8a68 , 
    R_aa1_1e18c168 , 
    R_591_1dda9648 , 
    R_99c_1e181e48 , 
    R_a42_1e188b08 , 
    R_ba8_1e6b6628 , 
    R_ae1_1e6ae9c8 , 
    R_9c2_1e183b08 , 
    R_6bb_1dfb50e8 , 
    R_41b_1d9dac28 , 
    R_93d_1e17e2e8 , 
    R_5b2_1ddaafe8 , 
    R_5d6_1d9dd388 , 
    R_402_1d9da188 , 
    R_4b0_1dda09a8 , 
    R_549_1dda6948 , 
    R_53a_1dda64e8 , 
    R_70d_1dfb8428 , 
    R_aa4_1e18c348 , 
    R_798_1dfbdb08 , 
    R_7fb_1e091948 , 
    R_32a_1d9d1a88 , 
    R_a36_1e188388 , 
    R_5ed_1ddacfc8 , 
    R_b9a_1e6b6268 , 
    R_c07_1e6ba188 , 
    R_47e_1dd9ef68 , 
    R_ad2_1e6ae568 , 
    R_39d_1d9d5d68 , 
    R_83f_1e0943c8 , 
    R_7eb_1e090f48 , 
    R_42e_1d9dbd08 , 
    R_b51_1e6b2fc8 , 
    R_6b4_1dfb4c88 , 
    R_694_1dfb3888 , 
    R_68f_1dfb3568 , 
    R_777_1dfbc668 , 
    R_7b0_1e08ea68 , 
    R_7a0_1e08e068 , 
    R_75e_1dfbbbc8 , 
    R_5b7_1ddaae08 , 
    R_63d_1dfb0228 , 
    R_636_1dfb02c8 , 
    R_8de_1e09ac28 , 
    R_2ef_1d9cf0a8 , 
    R_302_1d9d4508 , 
    R_9b8_1e182fc8 , 
    R_4b2_1dda14e8 , 
    R_8e4_1e09aae8 , 
    R_3de_1d9d8b08 , 
    R_ab8_1e18cfc8 , 
    R_71b_1dfb8ce8 , 
    R_c0c_1e6ba4a8 , 
    R_c2b_1e6bb808 , 
    R_5ac_1ddaa728 , 
    R_853_1e095048 , 
    R_2aa_1d9fca28 , 
    R_385_1d9d4e68 , 
    R_436_1d9dc208 , 
    R_a60_1e1898c8 , 
    R_7bb_1e08f148 , 
    R_811_1e092708 , 
    R_4c5_1dda16c8 , 
    R_406_1d9da408 , 
    R_473_1dd9e388 , 
    R_8aa_1e098ba8 , 
    R_b7e_1e6b50e8 , 
    R_7b5_1e08ed88 , 
    R_5fb_1ddad888 , 
    R_34d_1d9d2b68 , 
    R_ae3_1e6aeb08 , 
    R_6f3_1dfb73e8 , 
    R_82b_1e093748 , 
    R_72a_1dfbacc8 , 
    R_bc3_1e6b7708 , 
    R_8fa_1e09bda8 , 
    R_567_1dda7c08 , 
    R_89f_1e097fc8 , 
    R_3ed_1d9d8f68 , 
    R_599_1dda9b48 , 
    R_851_1e094f08 , 
    R_2dd_1d9ce568 , 
    R_4a8_1dda04a8 , 
    R_8a9_1e098608 , 
    R_366_1d9d4008 , 
    R_376_1ddad568 , 
    R_75d_1dfbb628 , 
    R_59a_1ddaa0e8 , 
    R_4c2_1dda19e8 , 
    R_8be_1e08eba8 , 
    R_2c5_1d9fd608 , 
    R_595_1dda98c8 , 
    R_446_1d9dd108 , 
    R_6c5_1dfb5728 , 
    R_5d8_1ddac2a8 , 
    R_682_1dfb3248 , 
    R_64b_1dfb0ae8 , 
    R_791_1dfbd6a8 , 
    R_b7b_1e6b4a08 , 
    R_3b1_1d9d69e8 , 
    R_7e9_1e090e08 , 
    R_beb_1e6b9008 , 
    R_6c0_1dfb5408 , 
    R_8ba_1e0995a8 , 
    R_a8e_1e17f508 , 
    R_3c8_1d9d7848 , 
    R_be4_1e6b8ba8 , 
    R_544_1dda6628 , 
    R_53f_1dda6308 , 
    R_90e_1e09ca28 , 
    R_381_1d9d4be8 , 
    R_a3e_1e188888 , 
    R_6fd_1dfb7a28 , 
    R_a3a_1e188608 , 
    R_8c2_1e099aa8 , 
    R_af0_1e6af328 , 
    R_296_1d9fb8a8 , 
    R_b12_1e6b0d68 , 
    R_ba9_1e6b66c8 , 
    R_b1d_1e6b0f48 , 
    R_2b5_1d9fcc08 , 
    R_6ff_1dfb7b68 , 
    R_a98_1e18bbc8 , 
    R_58e_1dda9968 , 
    R_753_1dfbafe8 , 
    R_3c5_1d9d7668 , 
    R_447_1d9dc7a8 , 
    R_61f_1dfaef68 , 
    R_54e_1dda28e8 , 
    R_6f8_1dfb7708 , 
    R_3a4_1d9d61c8 , 
    R_423_1d9db128 , 
    R_6a4_1dfb4288 , 
    R_b9b_1e6b5e08 , 
    R_a07_1e186128 , 
    R_55f_1dda7708 , 
    R_79d_1dfbde28 , 
    R_66d_1dfb2028 , 
    R_5e2_1ddacde8 , 
    R_48b_1dd9f288 , 
    R_5ee_1dda3a68 , 
    R_6c6_1dfb2d48 , 
    R_3e3_1d9d8928 , 
    R_b83_1e6b4f08 , 
    R_533_1dda5b88 , 
    R_42d_1d9db768 , 
    R_7e0_1e090868 , 
    R_696_1dfb3ec8 , 
    R_3f9_1d9d96e8 , 
    R_b88_1e6b5228 , 
    R_758_1dfbb308 , 
    R_3d2_1d9d8388 , 
    R_534_1dda5c28 , 
    R_532_1d9d1308 , 
    R_867_1e095cc8 , 
    R_2b6_1d9fd1a8 , 
    R_775_1dfbc528 , 
    R_3e8_1d9d8c48 , 
    R_4d0_1dda1da8 , 
    R_30d_1d9d0368 , 
    R_4e7_1dda2c08 , 
    R_70a_1dfb8748 , 
    R_a58_1e1893c8 , 
    R_4e8_1dda2ca8 , 
    R_4e6_1dda3068 , 
    R_535_1dda5cc8 , 
    R_5ea_1dda37e8 , 
    R_929_1e09d608 , 
    R_448_1d9dc848 , 
    R_b0b_1e6b0408 , 
    R_319_1d9d0ae8 , 
    R_985_1e180fe8 , 
    R_32f_1d9d18a8 , 
    R_4e9_1dda2d48 , 
    R_b1f_1e6b1088 , 
    R_495_1dd9f8c8 , 
    R_63b_1dfb00e8 , 
    R_536_1dda6268 , 
    R_3d9_1d9d82e8 , 
    R_a4f_1e188e28 , 
    R_470_1dd9e1a8 , 
    R_2d5_1d9ce068 , 
    R_3f0_1d9d9148 , 
    R_acf_1e18de28 , 
    R_ac2_1e18db08 , 
    R_9b4_1e182d48 , 
    R_a05_1e185fe8 , 
    R_2d9_1d9ce2e8 , 
    R_8ed_1e09b088 , 
    R_3f3_1d9d9328 , 
    R_af2_1e6af968 , 
    R_44d_1d9dcb68 , 
    R_645_1dfb0728 , 
    R_648_1dfb0908 , 
    R_4a1_1dda0048 , 
    R_749_1dfba9a8 , 
    R_2c8_1d9fd7e8 , 
    R_3bc_1d9d70c8 , 
    R_3f6_1ddad7e8 , 
    R_596_1dda9e68 , 
    R_c01_1e6b9dc8 , 
    R_734_1dfb9c88 , 
    R_5a5_1ddaa2c8 , 
    R_6e3_1dfb69e8 , 
    R_914_1e09c8e8 , 
    R_43d_1d9dc168 , 
    R_2cb_1d9fd9c8 , 
    R_3d0_1d9d7d48 , 
    R_b67_1e6b3d88 , 
    R_b01_1e6afdc8 , 
    R_37d_1d9d4968 , 
    R_a80_1e18acc8 , 
    R_9bd_1e1832e8 , 
    R_339_1d9d1ee8 , 
    R_7ad_1e08e888 , 
    R_972_1e180908 , 
    R_a22_1e184788 , 
    R_486_1ddacb68 , 
    R_5d5_1ddac0c8 , 
    R_592_1dda9be8 , 
    R_449_1d9dc8e8 , 
    R_87b_1e096948 , 
    R_8f5_1e09b588 , 
    R_35a_1d9d3888 , 
    R_37a_1ddab9e8 , 
    R_991_1e181768 , 
    R_62a_1dfb1448 , 
    R_808_1e092168 , 
    R_3a6_1d9d6808 , 
    R_b95_1e6b5a48 , 
    R_83e_1e17e108 , 
    R_386_1d9d5408 , 
    R_90d_1e09c488 , 
    R_931_1e09db08 , 
    R_ac9_1e18da68 , 
    R_a31_1e187b68 , 
    R_640_1dfb0408 , 
    R_667_1dfb1c68 , 
    R_6cb_1dfb5ae8 , 
    R_74a_1e17f288 , 
    R_676_1dfb2ac8 , 
    R_372_1d9d4788 , 
    R_56c_1dda7f28 , 
    R_334_1d9d1bc8 , 
    R_31e_1d9fc528 , 
    R_981_1e180d68 , 
    R_8ca_1e099fa8 , 
    R_85e_1e095c28 , 
    R_bbe_1e6af6e8 , 
    R_49b_1dd9fc88 , 
    R_73a_1dfba548 , 
    R_5fe_1dfaf8c8 , 
    R_98b_1e1813a8 , 
    R_88e_1e097a28 , 
    R_28f_1d9fb448 , 
    R_9bc_1e183248 , 
    R_5db_1ddac488 , 
    R_88a_1e08ee28 , 
    R_5a6_1ddaa868 , 
    R_443_1d9dc528 , 
    R_a0a_1e186808 , 
    R_358_1d9d3248 , 
    R_88f_1e0975c8 , 
    R_acc_1e18dc48 , 
    R_aac_1e18c848 , 
    R_2a2_1d9fde28 , 
    R_8a5_1e098388 , 
    R_8ec_1e09afe8 , 
    R_289_1d9fb088 , 
    R_340_1d9d2348 , 
    R_c2d_1e6bb948 , 
    R_964_1e17fb48 , 
    R_85d_1e095688 , 
    R_6fa_1dfb7d48 , 
    R_4d5_1dda20c8 , 
    R_a5a_1e18b308 , 
    R_7de_1e090c28 , 
    R_605_1ddadec8 , 
    R_311_1d9d05e8 , 
    R_8a6_1e098928 , 
    R_a2f_1e187a28 , 
    R_81f_1e092fc8 , 
    R_3b6_1d9d7208 , 
    R_315_1d9d0868 , 
    R_93f_1e17e428 , 
    R_5b1_1ddaaa48 , 
    R_631_1dfafaa8 , 
    R_890_1e097668 , 
    R_670_1dfb2208 , 
    R_b9c_1e6b5ea8 , 
    R_8e9_1e09ae08 , 
    R_932_1e093928 , 
    R_817_1e092ac8 , 
    R_b60_1e6b3928 , 
    R_979_1e180868 , 
    R_8d8_1e09a368 , 
    R_628_1dfaf508 , 
    R_729_1dfb95a8 , 
    R_a92_1e18bd08 , 
    R_b33_1e6b1d08 , 
    R_2ab_1d9fc5c8 , 
    R_5e6_1dd9f6e8 , 
    R_5c0_1ddab3a8 , 
    R_600_1ddadba8 , 
    R_8f4_1e09b4e8 , 
    R_29d_1d9fbd08 , 
    R_c11_1e6ba7c8 , 
    R_4d7_1dda2208 , 
    R_b43_1e6b2708 , 
    R_881_1e096d08 , 
    R_891_1e097708 , 
    R_8b4_1e098ce8 , 
    R_6ac_1dfb4788 , 
    R_2f0_1d9cf148 , 
    R_ad8_1e6ae428 , 
    R_9bb_1e1831a8 , 
    R_bd9_1e6b84c8 , 
    R_39f_1d9d5ea8 , 
    R_a5e_1e189c88 , 
    R_303_1d9cfd28 , 
    R_6ae_1dfb4dc8 , 
    R_477_1dd9e608 , 
    R_6d2_1e0981a8 , 
    R_38f_1d9d54a8 , 
    R_4d2_1dda23e8 , 
    R_82f_1e0939c8 , 
    R_61d_1dfaee28 , 
    R_673_1dfb23e8 , 
    R_578_1dda86a8 , 
    R_a65_1e189be8 , 
    R_9a5_1e1823e8 , 
    R_744_1dfba688 , 
    R_bfe_1e6ba0e8 , 
    R_86e_1e096628 , 
    R_6ce_1e0945a8 , 
    R_9df_1e184828 , 
    R_571_1dda8248 , 
    R_9e0_1e1848c8 , 
    R_9de_1e184c88 , 
    R_41a_1ddabee8 , 
    R_36e_1d9d1588 , 
    R_6b9_1dfb4fa8 , 
    R_b72_1e6b4968 , 
    R_73f_1dfba368 , 
    R_a4d_1e188ce8 , 
    R_9e1_1e184968 , 
    R_2d0_1d9fdce8 , 
    R_72e_1dfb9dc8 , 
    R_c25_1e6bb448 , 
    R_8eb_1e09af48 , 
    R_6eb_1dfb6ee8 , 
    R_764_1dfbba88 , 
    R_9b1_1e182b68 , 
    R_970_1e1802c8 , 
    R_bce_1e6b82e8 , 
    R_325_1d9d1268 , 
    R_65c_1dfb1588 , 
    R_643_1dfb05e8 , 
    R_abf_1e18d428 , 
    R_a9b_1e18bda8 , 
    R_b7c_1e6b4aa8 , 
    R_9ba_1e183608 , 
    R_bef_1e6b9288 , 
    R_b14_1e6b09a8 , 
    R_996_1e181f88 , 
    R_812_1e092ca8 , 
    R_4a2_1dda05e8 , 
    R_6e0_1dfb6808 , 
    R_490_1dd9f5a8 , 
    R_711_1dfb86a8 , 
    R_a86_1e18ba88 , 
    R_342_1d9d2988 , 
    R_c0e_1e6baae8 , 
    R_8e3_1e09aa48 , 
    R_646_1dfb0cc8 , 
    R_74d_1dfbac28 , 
    R_67f_1dfb2b68 , 
    R_34f_1d9d2ca8 , 
    R_8f3_1e09b448 , 
    R_bdc_1e6b86a8 , 
    R_57f_1dda8b08 , 
    R_77a_1dfbcd48 , 
    R_4c1_1dda1448 , 
    R_b8e_1e6b5ae8 , 
    R_c29_1e6bb6c8 , 
    R_875_1e096588 , 
    R_852_1e0954a8 , 
    R_6a6_1dfb48c8 , 
    R_76f_1dfbc168 , 
    R_984_1e180f48 , 
    R_39a_1d9d6088 , 
    R_35f_1d9d36a8 , 
    R_5d0_1ddabda8 , 
    R_b65_1e6b3c48 , 
    R_92b_1e09d748 , 
    R_3eb_1d9d8e28 , 
    R_53b_1dda6088 , 
    R_97a_1e180e08 , 
    R_369_1d9d3ce8 , 
    R_7f5_1e091588 , 
    R_588_1dda90a8 , 
    R_b6a_1e6b4468 , 
    R_435_1d9dbc68 , 
    R_a08_1e1861c8 , 
    R_7ef_1e0911c8 , 
    R_781_1dfbcca8 , 
    R_55c_1dda7528 , 
    R_3bf_1d9d72a8 , 
    R_850_1e094e68 , 
    R_2ea_1d9cf288 , 
    R_687_1dfb3068 , 
    R_795_1dfbd928 , 
    R_382_1d9d5188 , 
    R_63e_1dfb07c8 , 
    R_2b7_1d9fcd48 , 
    R_9b0_1e182ac8 , 
    R_6dd_1dfb6628 , 
    R_4be_1dda1768 , 
    R_bfd_1e6b9b48 , 
    R_b0d_1e6b0548 , 
    R_b9d_1e6b5f48 , 
    R_b3a_1e6b2668 , 
    R_4b9_1dda0f48 , 
    R_4bb_1dda1088 , 
    R_9a0_1e1820c8 , 
    R_83b_1e094148 , 
    R_8ea_1e09b3a8 , 
    R_b21_1e6b11c8 , 
    R_62f_1dfaf968 , 
    R_91d_1e09ce88 , 
    R_483_1dd9ed88 , 
    R_7c0_1e08f468 , 
    R_bd5_1e6b8248 , 
    R_364_1d9d39c8 , 
    R_322_1d9d2e88 , 
    R_326_1d9d1808 , 
    R_99b_1e181da8 , 
    R_961_1e17f968 , 
    R_726_1dfb98c8 , 
    R_a7d_1e18aae8 , 
    R_826_1e09de28 , 
    R_89a_1dfb4648 , 
    R_511_1dda4648 , 
    R_2fb_1d9cf828 , 
    R_b5c_1e6b36a8 , 
    R_8b0_1e098a68 , 
    R_708_1dfb8108 , 
    R_603_1ddadd88 , 
    R_804_1e091ee8 , 
    R_573_1dda8388 , 
    R_a56_1e189a08 , 
    R_510_1dda45a8 , 
    R_833_1e093c48 , 
    R_8c1_1e099508 , 
    R_966_1e180188 , 
    R_46d_1dd9dfc8 , 
    R_bcc_1e6b7ca8 , 
    R_47b_1dd9e888 , 
    R_aea_1e6af468 , 
    R_8d1_1e099f08 , 
    R_57a_1ddaa368 , 
    R_8f2_1e09b8a8 , 
    R_b35_1e6b1e48 , 
    R_b05_1e6b0048 , 
    R_aa9_1e18c668 , 
    R_9b7_1e182f28 , 
    R_3ae_1d9d6d08 , 
    R_50f_1dda4508 , 
    R_a23_1e1872a8 , 
    R_2c9_1d9fd888 , 
    R_5c6_1d9d7e88 , 
    R_8bd_1e099288 , 
    R_4b1_1dda0a48 , 
    R_b45_1e6b2848 , 
    R_422_1d9db588 , 
    R_2cc_1d9fda68 , 
    R_9d5_1e1841e8 , 
    R_37e_1d9d4f08 , 
    R_42c_1d9db6c8 , 
    R_a7e_1e18b088 , 
    R_a8d_1e18b4e8 , 
    R_50e_1dda4968 , 
    R_626_1dfafb48 , 
    R_5cc_1ddabb28 , 
    R_295_1d9fb808 , 
    R_a9e_1e18c488 , 
    R_80d_1e092488 , 
    R_9af_1e182a28 , 
    R_946_1e17ed88 , 
    R_a5c_1e189648 , 
    R_5bb_1ddab088 , 
    R_3e6_1d9d9008 , 
    R_ab3_1e18cca8 , 
    R_a1e_1e187488 , 
    R_66a_1dfb2348 , 
    R_7f8_1e091768 , 
    R_56e_1dda8568 , 
    R_3c2_1d9d7988 , 
    R_837_1e093ec8 , 
    R_866_1e096128 , 
    R_65a_1dfb1948 , 
    R_4aa_1dda0ae8 , 
    R_540_1dda63a8 , 
    R_61b_1dfaece8 , 
    R_78a_1dfbd748 , 
    R_76c_1dfbbf88 , 
    R_4c7_1dda1808 , 
    R_47f_1dd9eb08 , 
    R_34a_1d9d4a08 , 
    R_b57_1e6b3388 , 
    R_545_1dda66c8 , 
    R_c13_1e6ba908 , 
    R_44c_1d9dcac8 , 
    R_a0b_1e1863a8 , 
    R_6d5_1dfb6128 , 
    R_bf3_1e6b9508 , 
    R_3ee_1d9d9508 , 
    R_6d7_1dfb6268 , 
    R_3d6_1d9d9788 , 
    R_b06_1e6b05e8 , 
    R_9d4_1e184148 , 
    R_33b_1d9d2028 , 
    R_739_1dfb9fa8 , 
    R_a0e_1e186a88 , 
    R_7dd_1e090688 , 
    R_54f_1dda6d08 , 
    R_926_1e09dba8 , 
    R_abb_1e18d1a8 , 
    R_70e_1dfb89c8 , 
    R_ba2_1e6b6768 , 
    R_917_1e09cac8 , 
    R_923_1e09d248 , 
    R_784_1dfbce88 , 
    R_920_1e09d068 , 
    R_564_1dda7a28 , 
    R_9a9_1e182668 , 
    R_bfa_1e6b9e68 , 
    R_62c_1dfaf788 , 
    R_8c9_1e099a08 , 
    R_43c_1d9dc0c8 , 
    R_b00_1e6afd28 , 
    R_35d_1d9d3568 , 
    R_c18_1e6bac28 , 
    R_306_1d9d0408 , 
    R_939_1e17e068 , 
    R_474_1dd9e428 , 
    R_4a9_1dda0548 , 
    R_2ac_1d9fc668 , 
    R_609_1dfae1a8 , 
    R_94c_1e17ec48 , 
    R_90a_1e09c7a8 , 
    R_92e_1e0918a8 , 
    R_7be_1e08f828 , 
    R_825_1e093388 , 
    R_559_1dda7348 , 
    R_bf7_1e6b9788 , 
    R_87a_1e096da8 , 
    R_9d3_1e1840a8 , 
    R_394_1d9d57c8 , 
    R_31a_1d9d1088 , 
    R_69f_1dfb3f68 , 
    R_787_1dfbd068 , 
    R_a63_1e189aa8 , 
    R_9ae_1e183388 , 
    R_945_1e17e7e8 , 
    R_537_1dda5e08 , 
    R_725_1dfb9328 , 
    R_b68_1e6b3e28 , 
    R_7a5_1e08e388 , 
    R_4eb_1dda2e88 , 
    R_619_1dfaeba8 , 
    R_800_1e091c68 , 
    R_be8_1e6b8e28 , 
    R_4ec_1dda2f28 , 
    R_4ea_1dda32e8 , 
    R_2f1_1d9cf1e8 , 
    R_5d3_1ddabf88 , 
    R_6da_1dfb6948 , 
    R_5b6_1ddab268 , 
    R_3ac_1d9d66c8 , 
    R_983_1e180ea8 , 
    R_b73_1e6b4508 , 
    R_4ed_1dda2fc8 , 
    R_ada_1e6aea68 , 
    R_7fc_1e0919e8 , 
    R_b3c_1e6b22a8 , 
    R_304_1d9cfdc8 , 
    R_5ab_1ddaa688 , 
    R_85c_1e0955e8 , 
    R_442_1d9dcc08 , 
    R_3ce_1d9d8608 , 
    R_ad5_1e6ae248 , 
    R_ae8_1e6aee28 , 
    R_3b4_1d9d6bc8 , 
    R_8b8_1e098f68 , 
    R_b46_1e6b2de8 , 
    R_8e8_1e09ad68 , 
    R_bbf_1e6b7488 , 
    R_799_1dfbdba8 , 
    R_778_1dfbc708 , 
    R_a4b_1e188ba8 , 
    R_51d_1dda4dc8 , 
    R_657_1dfb1268 , 
    R_9d2_1e17f788 , 
    R_348_1d9d2848 , 
    R_51c_1dda4d28 , 
    R_8d7_1e09a2c8 , 
    R_9b3_1e182ca8 , 
    R_7db_1e090548 , 
    R_715_1dfb8928 , 
    R_68c_1dfb3388 , 
    R_880_1e096c68 , 
    R_29c_1d9fbc68 , 
    R_b7d_1e6b4b48 , 
    R_51b_1dda4c88 , 
    R_bba_1e6b7668 , 
    R_3dc_1d9d84c8 , 
    R_5a0_1dda9fa8 , 
    R_75f_1dfbb768 , 
    R_b7f_1e6b4c88 , 
    R_b16_1e6b0fe8 , 
    R_ba3_1e6b6308 , 
    R_654_1dfb1088 , 
    R_bc7_1e6b7988 , 
    R_2a3_1d9fc0c8 , 
    R_6f0_1dfb7208 , 
    R_7a1_1e08e108 , 
    R_371_1d9d41e8 , 
    R_51a_1dda50e8 , 
    R_ab7_1e18cf28 , 
    R_7e6_1e099828 , 
    R_b6b_1e6b4008 , 
    R_9ad_1e1828e8 , 
    R_935_1e09dd88 , 
    R_b8a_1e6bb768 , 
    R_69d_1dfb3e28 , 
    R_45e_1d9ddb08 , 
    R_a1a_1e187208 , 
    R_a49_1e188a68 , 
    R_a09_1e186268 , 
    R_496_1dd9fe68 , 
    R_336_1d9d2208 , 
    R_5df_1ddac708 , 
    R_5c7_1ddab808 , 
    R_990_1e1816c8 , 
    R_6c9_1dfb59a8 , 
    R_2eb_1d9cee28 , 
    R_2b8_1d9fcde8 , 
    R_ae0_1e6ae928 , 
    R_b2f_1e6b1a88 , 
    R_84d_1e094c88 , 
    R_a12_1e186d08 , 
    R_74f_1dfbad68 , 
    R_a35_1e187de8 , 
    R_28e_1d9fb3a8 , 
    R_81a_1e0936a8 , 
    R_487_1dd9f008 , 
    R_c1c_1e6baea8 , 
    R_7a8_1e08e568 , 
    R_471_1dd9e248 , 
    R_766_1e0986a8 , 
    R_38b_1d9d5228 , 
    R_a7b_1e18a9a8 , 
    R_b52_1e6b8568 , 
    R_9ff_1e185c28 , 
    R_7b9_1e08f008 , 
    R_67b_1dfb28e8 , 
    R_a00_1e185cc8 , 
    R_9fe_1e6bb9e8 , 
    R_980_1e180cc8 , 
    R_874_1e0964e8 , 
    R_49c_1dd9fd28 , 
    R_58c_1dda9328 , 
    R_45f_1d9dd6a8 , 
    R_98a_1e181808 , 
    R_8e2_1e09aea8 , 
    R_6ba_1dfb5548 , 
    R_bd8_1e6b8428 , 
    R_a8b_1e18b3a8 , 
    R_a01_1e185d68 , 
    R_6b3_1dfb4be8 , 
    R_60d_1dfae428 , 
    R_6e8_1dfb6d08 , 
    R_399_1d9d5ae8 , 
    R_a16_1e186f88 , 
    R_bc2_1e6b7b68 , 
    R_32b_1d9d1628 , 
    R_434_1d9dbbc8 , 
    R_a24_1e187348 , 
    R_377_1d9d45a8 , 
    R_3cc_1d9d7ac8 , 
    R_a68_1e189dc8 , 
    R_963_1e17faa8 , 
    R_7c5_1e08f788 , 
    R_615_1dfae928 , 
    R_8a2_1dfb9b48 , 
    R_722_1dfb9648 , 
    R_288_1d9f96e8 , 
    R_556_1dda7668 , 
    R_748_1dfba908 , 
    R_865_1e095b88 , 
    R_607_1dfae068 , 
    R_691_1dfb36a8 , 
    R_978_1e1807c8 , 
    R_84f_1e094dc8 , 
    R_2cd_1d9fdb08 , 
    R_ae2_1e6aef68 , 
    R_a1f_1e187028 , 
    R_721_1dfb90a8 , 
    R_733_1dfb9be8 , 
    R_9e3_1e184aa8 , 
    R_9e4_1e184b48 , 
    R_c23_1e6bb308 , 
    R_9e2_1e184f08 , 
    R_7ae_1dfbb1c8 , 
    R_91a_1e09d1a8 , 
    R_b84_1e6b4fa8 , 
    R_b92_1e181088 , 
    R_ba4_1e6b63a8 , 
    R_754_1dfbb088 , 
    R_5a4_1ddaa228 , 
    R_9a4_1e182348 , 
    R_b08_1e6b0228 , 
    R_9e5_1e184be8 , 
    R_617_1dfaea68 , 
    R_5ce_1ddac168 , 
    R_b89_1e6b52c8 , 
    R_7b2_1e09b128 , 
    R_460_1d9dd748 , 
    R_5e4_1ddaca28 , 
    R_30a_1d9d0688 , 
    R_a0c_1e186448 , 
    R_910_1e09c668 , 
    R_553_1dda6f88 , 
    R_86d_1e096088 , 
    R_a0f_1e186628 , 
    R_719_1dfb8ba8 , 
    R_b48_1e6b2a28 , 
    R_316_1d9d0e08 , 
    R_901_1e09bd08 , 
    R_611_1dfae6a8 , 
    R_ac5_1e18d7e8 , 
    R_6c4_1dfb5688 , 
    R_53c_1dda6128 , 
    R_712_1dfb8c48 , 
    R_2f6_1d9cfc88 , 
    R_829_1e093608 , 
    R_89d_1e097e88 , 
    R_8d0_1e099e68 , 
    R_8ac_1e0987e8 , 
    R_8a0_1e098068 , 
    R_aef_1e6af288 , 
    R_759_1dfbb3a8 , 
    R_a6d_1e18a0e8 , 
    R_6bf_1dfb5368 , 
    R_982_1e182c08 , 
    R_bdb_1e6b8608 , 
    R_684_1dfb2e88 , 
    R_7b7_1e08eec8 , 
    R_478_1dd9e6a8 , 
    R_be1_1e6b89c8 , 
    R_b55_1e6b3248 , 
    R_79b_1dfbdce8 , 
    R_c27_1e6bb588 , 
    R_96f_1e180228 , 
    R_42b_1d9db628 , 
    R_6cd_1dfb5c28 , 
    R_652_1dfb16c8 , 
    R_71d_1dfb8e28 , 
    R_703_1dfb7de8 , 
    R_a54_1e189148 , 
    R_4a3_1dda0188 , 
    R_634_1dfafc88 , 
    R_2ad_1d9fc708 , 
    R_4cc_1dda1b28 , 
    R_2a1_1d9fbf88 , 
    R_93a_1e0977a8 , 
    R_a78_1e18a7c8 , 
    R_c03_1e6b9f08 , 
    R_72c_1dfb9788 , 
    R_809_1e092208 , 
    R_5b0_1ddaa9a8 , 
    R_44b_1d9dca28 , 
    R_952_1ddab768 , 
    R_899_1e097c08 , 
    R_bd4_1e6b81a8 , 
    R_a94_1e18b948 , 
    R_6b1_1dfb4aa8 , 
    R_491_1dd9f648 , 
    R_5ca_1d9dae08 , 
    R_6f5_1dfb7528 , 
    R_9c9_1e183a68 , 
    R_75a_1dfbb948 , 
    R_461_1d9dd7e8 , 
    R_7c3_1e08f648 , 
    R_569_1dda7d48 , 
    R_a75_1e18a5e8 , 
    R_7ec_1e090fe8 , 
    R_c20_1e6bb128 , 
    R_96d_1e1800e8 , 
    R_54a_1dda6ee8 , 
    R_b31_1e6b1bc8 , 
    R_5bf_1ddab308 , 
    R_900_1e09bc68 , 
    R_b74_1e6b45a8 , 
    R_940_1e17e4c8 , 
    R_8dd_1e09a688 , 
    R_a88_1e18b1c8 , 
    R_743_1dfba5e8 , 
    R_2d1_1d9fdd88 , 
    R_4b3_1dda0b88 , 
    R_48c_1dd9f328 , 
    R_419_1d9daae8 , 
    R_2ba_1d9fd428 , 
    R_898_1e097b68 , 
    R_354_1d9d2fc8 , 
    R_3c9_1d9d78e8 , 
    R_afd_1e6afb48 , 
    R_698_1dfb3b08 , 
    R_8c8_1e099968 , 
    R_aff_1e6afc88 , 
    R_59c_1dda9d28 , 
    R_43b_1d9dc028 , 
    R_3e1_1d9d87e8 , 
    R_7d8_1e090368 , 
    R_624_1dfaf288 , 
    R_ace_1e6ae2e8 , 
    R_294_1d9fb768 , 
    R_818_1e092b68 , 
    R_9c8_1e1839c8 , 
    R_5c8_1ddab8a8 , 
    R_c2f_1e6bba88 , 
    R_ba5_1e6b6448 , 
    R_6d0_1dfb5e08 , 
    R_820_1e093068 , 
    R_30e_1d9d0908 , 
    R_99f_1e182028 , 
    R_73e_1dfba7c8 , 
    R_4ef_1dda3108 , 
    R_451_1d9dcde8 , 
    R_678_1dfb2708 , 
    R_663_1dfb19e8 , 
    R_5fa_1e091128 , 
    R_312_1d9d0b88 , 
    R_a45_1e1887e8 , 
    R_b18_1e6b0c28 , 
    R_4f0_1dda31a8 , 
    R_4ee_1dda3568 , 
    R_7ab_1e08e748 , 
    R_305_1d9cfe68 , 
    R_955_1e17f1e8 , 
    R_373_1d9d4328 , 
    R_a39_1e188068 , 
    R_669_1dfb1da8 , 
    R_3a5_1d9d6268 , 
    R_c0d_1e6ba548 , 
    R_4f1_1dda3248 , 
    R_541_1dda6448 , 
    R_69a_1dfb4148 , 
    R_b90_1e6b5728 , 
    R_99a_1e182208 , 
    R_960_1e17f8c8 , 
    R_6a9_1dfb45a8 , 
    R_4bc_1dda1128 , 
    R_897_1e097ac8 , 
    R_701_1dfb7ca8 , 
    R_36c_1d9d3ec8 , 
    R_60b_1dfae2e8 , 
    R_583_1dda8d88 , 
    R_330_1d9d1948 , 
    R_bb6_1e6b73e8 , 
    R_71e_1dfb93c8 , 
    R_590_1dda95a8 , 
    R_29e_1dda2668 , 
    R_b0f_1e6b0688 , 
    R_a1b_1e186da8 , 
    R_550_1dda6da8 , 
    R_ac8_1e18d9c8 , 
    R_a9d_1e18bee8 , 
    R_561_1dda7848 , 
    R_80e_1e092a28 , 
    R_9b6_1e187708 , 
    R_5e8_1ddacca8 , 
    R_613_1dfae7e8 , 
    R_b6c_1e6b40a8 , 
    R_3d3_1d9d7f28 , 
    R_31f_1d9d0ea8 , 
    R_9c7_1e183928 , 
    R_5dd_1ddac5c8 , 
    R_78e_1dfbd9c8 , 
    R_a13_1e1868a8 , 
    R_70c_1dfb8388 , 
    R_885_1e096f88 , 
    R_85b_1e095548 , 
    R_8ff_1e09bbc8 , 
    R_716_1dfb8ec8 , 
    R_2b9_1d9fce88 , 
    R_b69_1e6b3ec8 , 
    R_356_1d9d3608 , 
    R_2e6_1d9cf008 , 
    R_484_1dd9ee28 , 
    R_2ec_1d9ceec8 , 
    R_acb_1e18dba8 , 
    R_813_1e092848 , 
    R_4c3_1dda1588 , 
    R_a47_1e188928 , 
    R_81d_1e092e88 , 
    R_8e7_1e09acc8 , 
    R_5ef_1ddad108 , 
    R_896_1e094828 , 
    R_bec_1e6b90a8 , 
    R_b2b_1e6b1808 , 
    R_4ab_1dda0688 , 
    R_7e4_1e090ae8 , 
    R_a33_1e187ca8 , 
    R_47c_1dd9e928 , 
    R_8d6_1e09a728 , 
    R_87f_1e096bc8 , 
    R_5b5_1ddaacc8 , 
    R_651_1dfb0ea8 , 
    R_3da_1d9d8888 , 
    R_538_1dda5ea8 , 
    R_675_1dfb2528 , 
    R_60f_1dfae568 , 
    R_29b_1d9fbbc8 , 
    R_aa6_1e18c988 , 
    R_3bd_1d9d7168 , 
    R_be5_1e6b8c48 , 
    R_c0a_1e6ba868 , 
    R_5f5_1ddad4c8 , 
    R_b4b_1e6b2c08 , 
    R_7b1_1e08eb08 , 
    R_95d_1e17f6e8 , 
    R_a17_1e186b28 , 
    R_a29_1e187668 , 
    R_71a_1dfb9148 , 
    R_693_1dfb37e8 , 
    R_77b_1dfbc8e8 , 
    R_9c6_1e183d88 , 
    R_3a7_1d9d63a8 , 
    R_bc0_1e6b7528 , 
    R_68e_1dfb39c8 , 
    R_335_1d9d1c68 , 
    R_5eb_1ddace88 , 
    R_ad7_1e6ae388 , 
    R_765_1dfbbb28 , 
    R_387_1d9d4fa8 , 
    R_9a8_1e1825c8 , 
    R_632_1dfb0048 , 
    R_6e5_1dfb6b28 , 
    R_772_1dfbc848 , 
    R_995_1e1819e8 , 
    R_7d6_1e090728 , 
    R_598_1dda9aa8 , 
    R_a70_1e18a2c8 , 
    R_a25_1e1873e8 , 
    R_bbb_1e6b7208 , 
    R_6f2_1dfb7848 , 
    R_a41_1e188568 , 
    R_a66_1e18a188 , 
    R_a3d_1e1882e8 , 
    R_341_1d9d23e8 , 
    R_594_1dda9828 , 
    R_4fe_1dda5868 , 
    R_480_1dd9eba8 , 
    R_6ab_1dfb46e8 , 
    R_84c_1e094be8 , 
    R_660_1dfb1808 , 
    R_a20_1e1870c8 , 
    R_abe_1e6b64e8 , 
    R_566_1dda8068 , 
    R_7c8_1e08f968 , 
    R_5c2_1d9fc2a8 , 
    R_989_1e181268 , 
    R_8a8_1e098568 , 
    R_2a4_1d9fc168 , 
    R_7d5_1e090188 , 
    R_8fe_1e09c028 , 
    R_3b7_1d9d6da8 , 
    R_6b8_1dfb4f08 , 
    R_8b3_1e098c48 , 
    R_94f_1e17ee28 , 
    R_9fb_1e1859a8 , 
    R_a10_1e1866c8 , 
    R_b36_1e6b23e8 , 
    R_aa0_1e18c0c8 , 
    R_c1a_1e6bb268 , 
    R_82c_1e0937e8 , 
    R_4d1_1dda1e48 , 
    R_6fc_1dfb7988 , 
    R_9fa_1e185e08 , 
    R_9fc_1e185a48 , 
    R_a0d_1e1864e8 , 
    R_be2_1e6b8f68 , 
    R_b02_1e6b8068 , 
    R_a28_1e1875c8 , 
    R_4fd_1dda39c8 , 
    R_5fd_1ddad9c8 , 
    R_873_1e096448 , 
    R_9fd_1e185ae8 , 
    R_a6b_1e189fa8 , 
    R_aa3_1e18c2a8 , 
    R_738_1dfb9f08 , 
    R_805_1e091f88 , 
    R_2f7_1d9cf5a8 , 
    R_5ba_1ddab4e8 , 
    R_57d_1dda89c8 , 
    R_475_1dd9e4c8 , 
    R_433_1d9dbb28 , 
    R_aed_1e6af148 , 
    R_4fc_1dda3928 , 
    R_3a0_1d9d5f48 , 
    R_3f7_1d9d95a8 , 
    R_367_1d9d3ba8 , 
    R_947_1e17e928 , 
    R_b1a_1e6b1268 , 
    R_525_1dda52c8 , 
    R_50d_1dda43c8 , 
    R_390_1d9d5548 , 
    R_6fe_1dfb7fc8 , 
    R_6f7_1dfb7668 , 
    R_2ae_1d9fcca8 , 
    R_864_1e095ae8 , 
    R_9e7_1e184d28 , 
    R_524_1dda5228 , 
    R_50c_1dda4328 , 
    R_9e6_1e185188 , 
    R_9e8_1e184dc8 , 
    R_9b2_1e183108 , 
    R_7e2_1dfbaf48 , 
    R_622_1dfaf648 , 
    R_b4e_1e184508 , 
    R_a91_1e18b768 , 
    R_a84_1e18af48 , 
    R_4ce_1dda2168 , 
    R_bb2_1e6b7168 , 
    R_523_1dda5188 , 
    R_50b_1dda4288 , 
    R_9e9_1e184e68 , 
    R_4f3_1dda3388 , 
    R_4fb_1dda3888 , 
    R_4f2_1ddad068 , 
    R_4f4_1dda3428 , 
    R_55e_1dda7b68 , 
    R_84e_1e095228 , 
    R_a76_1e18ab88 , 
    R_5c9_1ddab948 , 
    R_343_1d9d2528 , 
    R_a73_1e18a4a8 , 
    R_7cd_1e08fc88 , 
    R_522_1dda55e8 , 
    R_50a_1dda46e8 , 
    R_4f5_1dda34c8 , 
    R_396_1d9d5e08 , 
    R_7f9_1e091808 , 
    R_681_1dfb2ca8 , 
    R_37b_1d9d4828 , 
    R_639_1dfaffa8 , 
    R_76d_1dfbc028 , 
    R_78b_1dfbd2e8 , 
    R_6a3_1dfb41e8 , 
    R_9ac_1e182848 , 
    R_86c_1e095fe8 , 
    R_c08_1e6ba228 , 
    R_2fc_1d9cf8c8 , 
    R_7f0_1e091268 , 
    R_c31_1e6bbbc8 , 
    R_a52_1e189508 , 
    R_ab2_1e18d108 , 
    R_28d_1d9fb308 , 
    R_bcb_1e6b7c08 , 
    R_4fa_1dda3f68 , 
    R_2bb_1d9fcfc8 , 
    R_b3f_1e6b2488 , 
    R_a27_1e187528 , 
    R_362_1d9d3d88 , 
    R_497_1dd9fa08 , 
    R_64f_1dfb0d68 , 
    R_bd7_1e6b8388 , 
    R_b75_1e6b4648 , 
    R_98f_1e181628 , 
    R_6ed_1dfb7028 , 
    R_7d3_1e090048 , 
    R_b27_1e6b1588 , 
    R_39b_1d9d5c28 , 
    R_8cf_1e099dc8 , 
    R_689_1dfb31a8 , 
    R_7c6_1e08fd28 , 
    R_b2d_1e6b1948 , 
    R_92a_1e092f28 , 
    R_66c_1dfb1f88 , 
    R_956_1e6b00e8 , 
    R_b96_1e18ce88 , 
    R_bae_1e6b6ee8 , 
    R_94d_1e17ece8 , 
    R_785_1dfbcf28 , 
    R_6e2_1dfb6e48 , 
    R_65e_1dfb5cc8 , 
    R_42a_1d9dba88 , 
    R_7e8_1e090d68 , 
    R_b4d_1e6b2d48 , 
    R_bff_1e6b9c88 , 
    R_3c0_1d9d7348 , 
    R_44a_1d9dce88 , 
    R_2fe_1d9cff08 , 
    R_383_1d9d4d28 , 
    R_928_1e09d568 , 
    R_488_1dd9f0a8 , 
    R_5aa_1ddaaae8 , 
    R_3fd_1d9d9968 , 
    R_7d0_1e08fe68 , 
    R_7b4_1e08ece8 , 
    R_4d8_1dda22a8 , 
    R_418_1d9daa48 , 
    R_a43_1e1886a8 , 
    R_327_1d9d13a8 , 
    R_849_1e094a08 , 
    R_b5f_1e6b3888 , 
    R_4d3_1dda1f88 , 
    R_a97_1e18bb28 , 
    R_aba_1e18d608 , 
    R_ab1_1e18cb68 , 
    R_97f_1e180c28 , 
    R_788_1dfbd108 , 
    R_a1c_1e186e48 , 
    R_b11_1e6b07c8 , 
    R_a37_1e187f28 , 
    R_801_1e091d08 , 
    R_581_1dda8c48 , 
    R_49d_1dd9fdc8 , 
    R_56b_1dda7e88 , 
    R_4da_1dda3ce8 , 
    R_7f2_1e09d6a8 , 
    R_53d_1dda61c8 , 
    R_3df_1d9d86a8 , 
    R_429_1d9db4e8 , 
    R_8dc_1e09a5e8 , 
    R_a14_1e186948 , 
    R_9d6_1e186088 , 
    R_add_1e6ae748 , 
    R_b6d_1e6b4148 , 
    R_c1e_1e6b4e68 , 
    R_7fd_1e091a88 , 
    R_859_1e095408 , 
    R_b23_1e6b1308 , 
    R_afc_1e6afaa8 , 
    R_913_1e09c848 , 
    R_450_1d9dcd48 , 
    R_7cb_1e08fb48 , 
    R_b38_1e6b2028 , 
    R_a26_1e187988 , 
    R_74c_1dfbab88 , 
    R_35b_1d9d3428 , 
    R_962_1e17ff08 , 
    R_2e7_1d9ceba8 , 
    R_8c0_1e099468 , 
    R_8c7_1e0998c8 , 
    R_afe_1e6b5d68 , 
    R_977_1e180728 , 
    R_925_1e09d388 , 
    R_919_1e09cc08 , 
    R_728_1dfb9508 , 
    R_43a_1d9dc488 , 
    R_bf0_1e6b9328 , 
    R_9a3_1e1822a8 , 
    R_3af_1d9d68a8 , 
    R_930_1e09da68 , 
    R_90c_1e09c3e8 , 
    R_5a9_1ddaa548 , 
    R_659_1dfb13a8 , 
    R_c0f_1e6ba688 , 
    R_307_1d9cffa8 , 
    R_8bc_1e0991e8 , 
    R_2ed_1d9cef68 , 
    R_770_1dfbc208 , 
    R_34b_1d9d2a28 , 
    R_37f_1d9d4aa8 , 
    R_5f4_1ddad428 , 
    R_779_1dfbc7a8 , 
    R_46a_1dd9f468 , 
    R_be0_1e6b8928 , 
    R_bd3_1e6b8108 , 
    R_466_1d9d9c88 , 
    R_77e_1dfbcfc8 , 
    R_575_1dda84c8 , 
    R_4ff_1dda3b08 , 
    R_a18_1e186bc8 , 
    R_bda_1e6b8a68 , 
    R_31b_1d9d0c28 , 
    R_3c6_1d9d7c08 , 
    R_792_1dfbdc48 , 
    R_54b_1dda6a88 , 
    R_6bd_1dfb5228 , 
    R_b50_1e6b2f28 , 
    R_a61_1e189968 , 
    R_b8b_1e6b5408 , 
    R_b80_1e6b4d28 , 
    R_33c_1d9d20c8 , 
    R_3c3_1d9d7528 , 
    R_666_1dfb20c8 , 
    R_c2a_1e6bbc68 , 
    R_359_1d9d32e8 , 
    R_415_1d9da868 , 
    R_5da_1ddac8e8 , 
    R_577_1dda8608 , 
    R_637_1dfafe68 , 
    R_9f7_1e185728 , 
    R_570_1dda81a8 , 
    R_9f6_1e185b88 , 
    R_9f8_1e1857c8 , 
    R_a6e_1e18a688 , 
    R_73d_1dfba228 , 
    R_293_1d9fb6c8 , 
    R_884_1e096ee8 , 
    R_3a2_1d9d6588 , 
    R_9f9_1e185868 , 
    R_957_1e17f328 , 
    R_ab6_1e6b5fe8 , 
    R_760_1dfbb808 , 
    R_a21_1e187168 , 
    R_bb7_1e6b6f88 , 
    R_9eb_1e184fa8 , 
    R_a3f_1e188428 , 
    R_747_1dfba868 , 
    R_4bf_1dda1308 , 
    R_3d7_1d9d81a8 , 
    R_4a4_1dda0228 , 
    R_441_1d9dc3e8 , 
    R_7ce_1e090228 , 
    R_85a_1e0959a8 , 
    R_66f_1dfb2168 , 
    R_9ea_1e185408 , 
    R_9ec_1e185048 , 
    R_a3b_1e1881a8 , 
    R_ad4_1e6ae1a8 , 
    R_b94_1e6b59a8 , 
    R_467_1d9ddba8 , 
    R_96e_1e180688 , 
    R_323_1d9d1128 , 
    R_6ea_1dfb7348 , 
    R_6ca_1dfb5f48 , 
    R_9ed_1e1850e8 , 
    R_ae7_1e6aed88 , 
    R_830_1e093a68 , 
    R_6d9_1dfb63a8 , 
    R_8e6_1e08f0a8 , 
    R_6a1_1dfb40a8 , 
    R_710_1dfb8608 , 
    R_b41_1e6b25c8 , 
    R_732_1dfba048 , 
    R_6df_1dfb6768 , 
    R_a11_1e186768 , 
    R_a8f_1e18b628 , 
    R_b97_1e6b5b88 , 
    R_bc6_1e6b7de8 , 
    R_4db_1dda2488 , 
    R_9d7_1e184328 , 
    R_b29_1e6b16c8 , 
    R_57e_1dda8f68 , 
    R_29a_1d9fbb28 , 
    R_36f_1d9d40a8 , 
    R_3e4_1d9d89c8 , 
    R_7bc_1e08f1e8 , 
    R_87e_1e097028 , 
    R_b1c_1e6b0ea8 , 
    R_aab_1e18c7a8 , 
    R_96c_1e180048 , 
    R_551_1dda6e48 , 
    R_6d4_1dfb6088 , 
    R_2af_1d9fc848 , 
    R_479_1dd9e748 , 
    R_5a3_1ddaa188 , 
    R_672_1dfb2848 , 
    R_587_1dda9008 , 
    R_767_1dfbbc68 , 
    R_395_1d9d5868 , 
    R_3e9_1d9d8ce8 , 
    R_2f8_1d9cf648 , 
    R_64c_1dfb0b88 , 
    R_5e1_1ddac848 , 
    R_3fc_1d9d98c8 , 
    R_468_1d9ddc48 , 
    R_3ba_1d9d7488 , 
    R_55b_1dda7488 , 
    R_67e_1dfb2fc8 , 
    R_8b7_1e098ec8 , 
    R_879_1e096808 , 
    R_b5b_1e6b3608 , 
    R_a82_1e18b588 , 
    R_ae5_1e6aec48 , 
    R_84b_1e094b48 , 
    R_99e_1e182488 , 
    R_6dc_1dfb6588 , 
    R_3ad_1d9d6768 , 
    R_a59_1e189468 , 
    R_b62_1e6ba368 , 
    R_731_1dfb9aa8 , 
    R_3f1_1d9d91e8 , 
    R_620_1dfaf008 , 
    R_67d_1dfb2a28 , 
    R_adf_1e6ae888 , 
    R_349_1d9d28e8 , 
    R_3d1_1d9d7de8 , 
    R_3f4_1d9d93c8 , 
    R_80a_1e0927a8 , 
    R_350_1d9d2d48 , 
    R_a50_1e188ec8 , 
    R_bc1_1e6b75c8 , 
    R_b85_1e6b5048 , 
    R_5d7_1ddac208 , 
    R_7a2_1ddada68 , 
    R_539_1dda5f48 , 
    R_bbc_1e6b72a8 , 
    R_c14_1e6ba9a8 , 
    R_6c8_1dfb5908 , 
    R_4c8_1dda18a8 , 
    R_360_1d9d3748 , 
    R_2e2_1d9ced88 , 
    R_936_1e17e388 , 
    R_9f3_1e1854a8 , 
    R_b25_1e6b1448 , 
    R_b0a_1e6b0868 , 
    R_b56_1e6b87e8 , 
    R_bf4_1e6b95a8 , 
    R_95f_1e17f828 , 
    R_3b5_1d9d6c68 , 
    R_52a_1dda5fe8 , 
    R_9f2_1e185908 , 
    R_9f4_1e185548 , 
    R_686_1dfb34c8 , 
    R_2bc_1d9fd068 , 
    R_7a6_1e08e928 , 
    R_9ef_1e185228 , 
    R_b1e_1e6b78e8 , 
    R_bfb_1e6b9a08 , 
    R_378_1d9d4648 , 
    R_9ee_1e185688 , 
    R_9f0_1e1852c8 , 
    R_9f5_1e1855e8 , 
    R_4bd_1dda11c8 , 
    R_5af_1ddaa908 , 
    R_822_1e097f28 , 
    R_872_1e0968a8 , 
    R_9f1_1e185368 , 
    R_337_1d9d1da8 , 
    R_707_1dfb8068 , 
    R_755_1dfbb128 , 
    R_8f9_1e09b808 , 
    R_432_1d9dbf88 , 
    R_8af_1e0989c8 , 
    R_bc5_1e6b7848 , 
    R_934_1e09dce8 , 
    R_469_1d9ddce8 , 
    R_572_1dda87e8 , 
    R_863_1e095a48 , 
    R_958_1e17f3c8 , 
    R_742_1dfbaa48 , 
    R_2a5_1d9fc208 , 
    R_a9a_1e18c208 , 
    R_af9_1e6af8c8 , 
    R_9c1_1e183568 , 
    R_83c_1e0941e8 , 
    R_a81_1e18ad68 , 
    R_c19_1e6bacc8 , 
    R_91c_1e09cde8 , 
    R_4ac_1dda0728 , 
    R_bf8_1e6b9828 , 
    R_5be_1dda7168 , 
    R_93b_1e17e1a8 , 
    R_63c_1dfb0188 , 
    R_7e1_1e090908 , 
    R_7ba_1e08f5a8 , 
    R_6b2_1dfb5048 , 
    R_4dc_1dda2528 , 
    R_79e_1e08e428 , 
    R_492_1dd9fbe8 , 
    R_750_1dfbae08 , 
    R_9d8_1e1843c8 , 
    R_365_1d9d3a68 , 
    R_994_1e181948 , 
    R_95c_1e17f648 , 
    R_2ff_1d9cfaa8 , 
    R_89b_1e097d48 , 
    R_827_1e0934c8 , 
    R_332_1d9d1f88 , 
    R_9a7_1e182528 , 
    R_834_1e093ce8 , 
    R_30b_1d9d0228 , 
    R_86b_1e095f48 , 
    R_649_1dfb09a8 , 
    R_a1d_1e186ee8 , 
    R_b59_1e6b34c8 , 
    R_bb3_1e6b6d08 , 
    R_796_1e08e1a8 , 
    R_941_1e17e568 , 
    R_be9_1e6b8ec8 , 
    R_485_1dd9eec8 , 
    R_317_1d9d09a8 , 
    R_8a3_1e098248 , 
    R_49e_1dda0368 , 
    R_9c0_1e1834c8 , 
    R_32c_1d9d16c8 , 
    R_6d6_1dfb66c8 , 
    R_a15_1e1869e8 , 
    R_33e_1d9d2708 , 
    R_38c_1d9d52c8 , 
    R_75b_1dfbb4e8 , 
    R_ac4_1e18d748 , 
    R_5d9_1ddac348 , 
    R_546_1dda6c68 , 
    R_2be_1d9fd6a8 , 
    R_b76_1e6b4be8 , 
    R_975_1e1805e8 , 
    R_5c3_1ddab588 , 
    R_500_1dda3ba8 , 
    R_889_1e097208 , 
    R_988_1e1811c8 , 
    R_c2c_1e6bb8a8 , 
    R_b98_1e6b5c28 , 
    R_47d_1dd9e9c8 , 
    R_417_1d9da9a8 , 
    R_819_1e092c08 , 
    R_8f8_1e09b768 , 
    R_942_1e17eb08 , 
    R_ad1_1e6adfc8 , 
    R_8ce_1e09a228 , 
    R_563_1dda7988 , 
    R_2e8_1d9cec48 , 
    R_838_1e093f68 , 
    R_aee_1e187c08 , 
    R_641_1dfb04a8 , 
    R_c16_1e6b41e8 , 
    R_6c3_1dfb55e8 , 
    R_5f3_1ddad388 , 
    R_558_1dda72a8 , 
    R_821_1e093108 , 
    R_a5f_1e189828 , 
    R_3cd_1d9d7b68 , 
    R_80f_1e0925c8 , 
    R_724_1dfb9288 , 
    R_848_1e094968 , 
    R_9bf_1e183428 , 
    R_a19_1e186c68 , 
    R_baf_1e6b6a88 , 
    R_64a_1dfb0f48 , 
    R_aa8_1e18c5c8 , 
    R_6be_1dfb57c8 , 
    R_481_1dd9ec48 , 
    R_428_1d9db448 , 
    R_be6_1e6b91e8 , 
    R_44f_1d9dcca8 , 
    R_5b4_1ddaac28 , 
    R_629_1dfaf5a8 , 
    R_78f_1dfbd568 , 
    R_91f_1e09cfc8 , 
    R_858_1e095368 , 
    R_afb_1e6afa08 , 
    R_3fb_1d9d9828 , 
    R_922_1e091628 , 
    R_916_1e09cf28 , 
    R_8a1_1e098108 , 
    R_8db_1e09a548 , 
    R_b32_1e6b2168 , 
    R_411_1d9da5e8 , 
    R_6b0_1dfb4a08 , 
    R_5d1_1ddabe48 , 
    R_7df_1e0907c8 , 
    R_b04_1e6affa8 , 
    R_45a_1d9dd888 , 
    R_814_1e0928e8 , 
    R_665_1dfb1b28 , 
    R_69e_1dfb43c8 , 
    R_b42_1e6b2b68 , 
    R_555_1dda70c8 , 
    R_374_1d9d43c8 , 
    R_352_1d9d3388 , 
    R_2a6_1d9fc7a8 , 
    R_756_1dfbb6c8 , 
    R_bd6_1e6b3568 , 
    R_baa_1e18d888 , 
    R_5b9_1ddaaf48 , 
    R_3ec_1d9d8ec8;
wire n273708 , n273709 , n273710 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , 
     n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , 
     n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , 
     n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , 
     n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , 
     n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , 
     n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , 
     n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , 
     n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , 
     n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , 
     n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , 
     n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , 
     n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , 
     n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , 
     n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , 
     n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , 
     n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , 
     n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , 
     n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , 
     n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , 
     n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , 
     n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , 
     n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , 
     n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , 
     n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , 
     n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , 
     n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , 
     n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , 
     n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , 
     n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , 
     n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , 
     n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , 
     n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , 
     n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , 
     n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , 
     n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , 
     n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , 
     n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , 
     n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , 
     n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , 
     n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , 
     n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , 
     n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , 
     n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , 
     n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , 
     n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , 
     n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , 
     n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , 
     n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , 
     n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , 
     n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , 
     n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , 
     n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , 
     n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , 
     n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , 
     n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , 
     n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , 
     n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , 
     n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , 
     n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , 
     n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , 
     n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , 
     n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , 
     n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , 
     n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , 
     n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , 
     n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , 
     n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , 
     n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , 
     n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , 
     n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , 
     n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , 
     n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , 
     n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , 
     n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , 
     n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , 
     n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , 
     n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , 
     n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , 
     n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , 
     n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , 
     n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , 
     n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , 
     n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , 
     n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , 
     n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , 
     n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , 
     n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , 
     n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , 
     n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , 
     n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , 
     n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , 
     n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , 
     n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , 
     n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , 
     n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , 
     n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , 
     n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , 
     n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , 
     n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , 
     n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , 
     n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , 
     n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , 
     n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , 
     n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , 
     n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , 
     n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , 
     n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , 
     n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , 
     n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , 
     n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , 
     n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , 
     n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , 
     n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , 
     n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , 
     n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , 
     n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , 
     n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , 
     n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , 
     n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , 
     n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , 
     n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , 
     n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n274934 , n274935 , n274936 , 
     n274937 , n274938 , n274939 , n274940 , n274941 , n274942 , n274943 , n274944 , n274945 , n274946 , 
     n274947 , n274948 , n274949 , n274950 , n274951 , n274952 , n274953 , n274954 , n274955 , n274956 , 
     n274957 , n274958 , n274959 , n274960 , n274961 , n274962 , n274963 , n274964 , n274965 , n274966 , 
     n274967 , n274968 , n274969 , n274970 , n274971 , n274972 , n274973 , n274974 , n274975 , n274976 , 
     n274977 , n274978 , n274979 , n274980 , n274981 , n274982 , n274983 , n274984 , n274985 , n274986 , 
     n274987 , n274988 , n274989 , n274990 , n274991 , n274992 , n274993 , n274994 , n274995 , n274996 , 
     n274997 , n274998 , n274999 , n275000 , n275001 , n275002 , n275003 , n275004 , n275005 , n275006 , 
     n275007 , n275008 , n275009 , n275010 , n275011 , n275012 , n275013 , n275014 , n275015 , n275016 , 
     n275017 , n275018 , n275019 , n275020 , n275021 , n275022 , n275023 , n275024 , n275025 , n275026 , 
     n275027 , n275028 , n275029 , n275030 , n275031 , n275032 , n275033 , n275034 , n275035 , n275036 , 
     n275037 , n275038 , n275039 , n275040 , n275041 , n275042 , n275043 , n275044 , n275045 , n275046 , 
     n275047 , n275048 , n275049 , n275050 , n275051 , n275052 , n275053 , n275054 , n275055 , n275056 , 
     n275057 , n275058 , n275059 , n275060 , n275061 , n275062 , n275063 , n275064 , n275065 , n275066 , 
     n275067 , n275068 , n275069 , n275070 , n275071 , n275072 , n275073 , n275074 , n275075 , n275076 , 
     n275077 , n275078 , n275079 , n275080 , n275081 , n275082 , n275083 , n275084 , n275085 , n275086 , 
     n275087 , n275088 , n275089 , n275090 , n275091 , n275092 , n275093 , n275094 , n275095 , n275096 , 
     n275097 , n275098 , n275099 , n275100 , n275101 , n275102 , n275103 , n275104 , n275105 , n275106 , 
     n275107 , n275108 , n275109 , n275110 , n275111 , n275112 , n275113 , n275114 , n275115 , n275116 , 
     n275117 , n275118 , n275119 , n275120 , n275121 , n275122 , n275123 , n275124 , n275125 , n275126 , 
     n275127 , n275128 , n275129 , n275130 , n275131 , n275132 , n275133 , n275134 , n275135 , n275136 , 
     n275137 , n275138 , n275139 , n275140 , n275141 , n275142 , n275143 , n275144 , n275145 , n275146 , 
     n275147 , n275148 , n275149 , n275150 , n275151 , n275152 , n275153 , n275154 , n275155 , n275156 , 
     n275157 , n275158 , n275159 , n275160 , n275161 , n275162 , n275163 , n275164 , n275165 , n275166 , 
     n275167 , n275168 , n275169 , n275170 , n275171 , n275172 , n275173 , n275174 , n275175 , n275176 , 
     n275177 , n275178 , n275179 , n275180 , n275181 , n275182 , n275183 , n275184 , n275185 , n275186 , 
     n275187 , n275188 , n275189 , n275190 , n275191 , n275192 , n275193 , n275194 , n275195 , n275196 , 
     n275197 , n275198 , n275199 , n275200 , n275201 , n275202 , n275203 , n275204 , n275205 , n275206 , 
     n275207 , n275208 , n275209 , n275210 , n275211 , n275212 , n275213 , n275214 , n275215 , n275216 , 
     n275217 , n275218 , n275219 , n275220 , n275221 , n275222 , n275223 , n275224 , n275225 , n275226 , 
     n275227 , n275228 , n275229 , n275230 , n275231 , n275232 , n275233 , n275234 , n275235 , n275236 , 
     n275237 , n275238 , n275239 , n275240 , n275241 , n275242 , n275243 , n275244 , n275245 , n275246 , 
     n275247 , n275248 , n275249 , n275250 , n275251 , n275252 , n275253 , n275254 , n275255 , n275256 , 
     n275257 , n275258 , n275259 , n275260 , n275261 , n275262 , n275263 , n275264 , n275265 , n275266 , 
     n275267 , n275268 , n275269 , n275270 , n275271 , n275272 , n275273 , n275274 , n275275 , n275276 , 
     n275277 , n275278 , n275279 , n275280 , n275281 , n275282 , n275283 , n275284 , n275285 , n275286 , 
     n275287 , n275288 , n275289 , n275290 , n275291 , n275292 , n275293 , n275294 , n275295 , n275296 , 
     n275297 , n275298 , n275299 , n275300 , n275301 , n275302 , n275303 , n275304 , n275305 , n275306 , 
     n275307 , n275308 , n275309 , n275310 , n275311 , n275312 , n275313 , n275314 , n275315 , n275316 , 
     n275317 , n275318 , n275319 , n275320 , n275321 , n275322 , n275323 , n275324 , n275325 , n275326 , 
     n275327 , n275328 , n275329 , n275330 , n275331 , n275332 , n275333 , n275334 , n275335 , n275336 , 
     n275337 , n275338 , n275339 , n275340 , n275341 , n275342 , n275343 , n275344 , n275345 , n275346 , 
     n275347 , n275348 , n275349 , n275350 , n275351 , n275352 , n275353 , n275354 , n275355 , n275356 , 
     n275357 , n275358 , n275359 , n275360 , n275361 , n275362 , n275363 , n275364 , n275365 , n275366 , 
     n275367 , n275368 , n275369 , n275370 , n275371 , n275372 , n275373 , n275374 , n275375 , n275376 , 
     n275377 , n275378 , n275379 , n275380 , n275381 , n275382 , n275383 , n275384 , n275385 , n275386 , 
     n275387 , n275388 , n275389 , n275390 , n275391 , n275392 , n275393 , n275394 , n275395 , n275396 , 
     n275397 , n275398 , n275399 , n275400 , n275401 , n275402 , n275403 , n275404 , n275405 , n275406 , 
     n275407 , n275408 , n275409 , n275410 , n275411 , n275412 , n275413 , n275414 , n275415 , n275416 , 
     n275417 , n275418 , n275419 , n275420 , n275421 , n275422 , n275423 , n275424 , n275425 , n275426 , 
     n275427 , n275428 , n275429 , n275430 , n275431 , n275432 , n275433 , n275434 , n275435 , n275436 , 
     n275437 , n275438 , n275439 , n275440 , n275441 , n275442 , n275443 , n275444 , n275445 , n275446 , 
     n275447 , n275448 , n275449 , n275450 , n275451 , n275452 , n275453 , n275454 , n275455 , n275456 , 
     n275457 , n275458 , n275459 , n275460 , n275461 , n275462 , n275463 , n275464 , n275465 , n275466 , 
     n275467 , n275468 , n275469 , n275470 , n275471 , n275472 , n275473 , n275474 , n275475 , n275476 , 
     n275477 , n275478 , n275479 , n275480 , n275481 , n275482 , n275483 , n275484 , n275485 , n275486 , 
     n275487 , n275488 , n275489 , n275490 , n275491 , n275492 , n275493 , n275494 , n275495 , n275496 , 
     n275497 , n275498 , n275499 , n275500 , n275501 , n275502 , n275503 , n275504 , n275505 , n275506 , 
     n275507 , n275508 , n275509 , n275510 , n275511 , n275512 , n275513 , n275514 , n275515 , n275516 , 
     n275517 , n275518 , n275519 , n275520 , n275521 , n275522 , n275523 , n275524 , n275525 , n275526 , 
     n275527 , n275528 , n275529 , n275530 , n275531 , n275532 , n275533 , n275534 , n275535 , n275536 , 
     n275537 , n275538 , n275539 , n275540 , n275541 , n275542 , n275543 , n275544 , n275545 , n275546 , 
     n275547 , n275548 , n275549 , n275550 , n275551 , n275552 , n275553 , n275554 , n275555 , n275556 , 
     n275557 , n275558 , n275559 , n275560 , n275561 , n275562 , n275563 , n275564 , n275565 , n275566 , 
     n275567 , n275568 , n275569 , n275570 , n275571 , n275572 , n275573 , n275574 , n275575 , n275576 , 
     n275577 , n275578 , n275579 , n275580 , n275581 , n275582 , n275583 , n275584 , n275585 , n275586 , 
     n275587 , n275588 , n275589 , n275590 , n275591 , n275592 , n275593 , n275594 , n275595 , n275596 , 
     n275597 , n275598 , n275599 , n275600 , n275601 , n275602 , n275603 , n275604 , n275605 , n275606 , 
     n275607 , n275608 , n275609 , n275610 , n275611 , n275612 , n275613 , n275614 , n275615 , n275616 , 
     n275617 , n275618 , n275619 , n275620 , n275621 , n275622 , n275623 , n275624 , n275625 , n275626 , 
     n275627 , n275628 , n275629 , n275630 , n275631 , n275632 , n275633 , n275634 , n275635 , n275636 , 
     n275637 , n275638 , n275639 , n275640 , n275641 , n275642 , n275643 , n275644 , n275645 , n275646 , 
     n275647 , n275648 , n275649 , n275650 , n275651 , n275652 , n275653 , n275654 , n275655 , n275656 , 
     n275657 , n275658 , n275659 , n275660 , n275661 , n275662 , n275663 , n275664 , n275665 , n275666 , 
     n275667 , n275668 , n275669 , n275670 , n275671 , n275672 , n275673 , n275674 , n275675 , n275676 , 
     n275677 , n275678 , n275679 , n275680 , n275681 , n275682 , n275683 , n275684 , n275685 , n275686 , 
     n275687 , n275688 , n275689 , n275690 , n275691 , n275692 , n275693 , n275694 , n275695 , n275696 , 
     n275697 , n275698 , n275699 , n275700 , n275701 , n275702 , n275703 , n275704 , n275705 , n275706 , 
     n275707 , n275708 , n275709 , n275710 , n275711 , n275712 , n275713 , n275714 , n275715 , n275716 , 
     n275717 , n275718 , n275719 , n275720 , n275721 , n275722 , n275723 , n275724 , n275725 , n275726 , 
     n275727 , n275728 , n275729 , n275730 , n275731 , n275732 , n275733 , n275734 , n275735 , n275736 , 
     n275737 , n275738 , n275739 , n275740 , n275741 , n275742 , n275743 , n275744 , n275745 , n275746 , 
     n275747 , n275748 , n275749 , n275750 , n275751 , n275752 , n275753 , n275754 , n275755 , n275756 , 
     n275757 , n275758 , n275759 , n275760 , n275761 , n275762 , n275763 , n275764 , n275765 , n275766 , 
     n275767 , n275768 , n275769 , n275770 , n275771 , n275772 , n275773 , n275774 , n275775 , n275776 , 
     n275777 , n275778 , n275779 , n275780 , n275781 , n275782 , n275783 , n275784 , n275785 , n275786 , 
     n275787 , n275788 , n275789 , n275790 , n275791 , n275792 , n275793 , n275794 , n275795 , n275796 , 
     n275797 , n275798 , n275799 , n275800 , n275801 , n275802 , n275803 , n275804 , n275805 , n275806 , 
     n275807 , n275808 , n275809 , n275810 , n275811 , n275812 , n275813 , n275814 , n275815 , n275816 , 
     n275817 , n275818 , n275819 , n275820 , n275821 , n275822 , n275823 , n275824 , n275825 , n275826 , 
     n275827 , n275828 , n275829 , n275830 , n275831 , n275832 , n275833 , n275834 , n275835 , n275836 , 
     n275837 , n275838 , n275839 , n275840 , n275841 , n275842 , n275843 , n275844 , n275845 , n275846 , 
     n275847 , n275848 , n275849 , n275850 , n275851 , n275852 , n275853 , n275854 , n275855 , n275856 , 
     n275857 , n275858 , n275859 , n275860 , n275861 , n275862 , n275863 , n275864 , n275865 , n275866 , 
     n275867 , n275868 , n275869 , n275870 , n275871 , n275872 , n275873 , n275874 , n275875 , n275876 , 
     n275877 , n275878 , n275879 , n275880 , n275881 , n275882 , n275883 , n275884 , n275885 , n275886 , 
     n275887 , n275888 , n275889 , n275890 , n275891 , n275892 , n275893 , n275894 , n275895 , n275896 , 
     n275897 , n275898 , n275899 , n275900 , n275901 , n275902 , n275903 , n275904 , n275905 , n275906 , 
     n275907 , n275908 , n275909 , n275910 , n275911 , n275912 , n275913 , n275914 , n275915 , n275916 , 
     n275917 , n275918 , n275919 , n275920 , n275921 , n275922 , n275923 , n275924 , n275925 , n275926 , 
     n275927 , n275928 , n275929 , n275930 , n275931 , n275932 , n275933 , n275934 , n275935 , n275936 , 
     n275937 , n275938 , n275939 , n275940 , n275941 , n275942 , n275943 , n275944 , n275945 , n275946 , 
     n275947 , n275948 , n275949 , n275950 , n275951 , n275952 , n275953 , n275954 , n275955 , n275956 , 
     n275957 , n275958 , n275959 , n275960 , n275961 , n275962 , n275963 , n275964 , n275965 , n275966 , 
     n275967 , n275968 , n275969 , n275970 , n275971 , n275972 , n275973 , n275974 , n275975 , n275976 , 
     n275977 , n275978 , n275979 , n275980 , n275981 , n275982 , n275983 , n275984 , n275985 , n275986 , 
     n275987 , n275988 , n275989 , n275990 , n275991 , n275992 , n275993 , n275994 , n275995 , n275996 , 
     n275997 , n275998 , n275999 , n276000 , n276001 , n276002 , n276003 , n276004 , n276005 , n276006 , 
     n276007 , n276008 , n276009 , n276010 , n276011 , n276012 , n276013 , n276014 , n276015 , n276016 , 
     n276017 , n276018 , n276019 , n276020 , n276021 , n276022 , n276023 , n276024 , n276025 , n276026 , 
     n276027 , n276028 , n276029 , n276030 , n276031 , n276032 , n276033 , n276034 , n276035 , n276036 , 
     n276037 , n276038 , n276039 , n276040 , n276041 , n276042 , n276043 , n276044 , n276045 , n276046 , 
     n276047 , n276048 , n276049 , n276050 , n276051 , n276052 , n276053 , n276054 , n276055 , n276056 , 
     n276057 , n276058 , n276059 , n276060 , n276061 , n276062 , n276063 , n276064 , n276065 , n276066 , 
     n276067 , n276068 , n276069 , n276070 , n276071 , n276072 , n276073 , n276074 , n276075 , n276076 , 
     n276077 , n276078 , n276079 , n276080 , n276081 , n276082 , n276083 , n276084 , n276085 , n276086 , 
     n276087 , n276088 , n276089 , n276090 , n276091 , n276092 , n276093 , n276094 , n276095 , n276096 , 
     n276097 , n276098 , n276099 , n276100 , n276101 , n276102 , n276103 , n276104 , n276105 , n276106 , 
     n276107 , n276108 , n276109 , n276110 , n276111 , n276112 , n276113 , n276114 , n276115 , n276116 , 
     n276117 , n276118 , n276119 , n276120 , n276121 , n276122 , n276123 , n276124 , n276125 , n276126 , 
     n276127 , n276128 , n276129 , n276130 , n276131 , n276132 , n276133 , n276134 , n276135 , n276136 , 
     n276137 , n276138 , n276139 , n276140 , n276141 , n276142 , n276143 , n276144 , n276145 , n276146 , 
     n276147 , n276148 , n276149 , n276150 , n276151 , n276152 , n276153 , n276154 , n276155 , n276156 , 
     n276157 , n276158 , n276159 , n276160 , n276161 , n276162 , n276163 , n276164 , n276165 , n276166 , 
     n276167 , n276168 , n276169 , n276170 , n276171 , n276172 , n276173 , n276174 , n276175 , n276176 , 
     n276177 , n276178 , n276179 , n276180 , n276181 , n276182 , n276183 , n276184 , n276185 , n276186 , 
     n276187 , n276188 , n276189 , n276190 , n276191 , n276192 , n276193 , n276194 , n276195 , n276196 , 
     n276197 , n276198 , n276199 , n276200 , n276201 , n276202 , n276203 , n276204 , n276205 , n276206 , 
     n276207 , n276208 , n276209 , n276210 , n276211 , n276212 , n276213 , n276214 , n276215 , n276216 , 
     n276217 , n276218 , n276219 , n276220 , n276221 , n276222 , n276223 , n276224 , n276225 , n276226 , 
     n276227 , n276228 , n276229 , n276230 , n276231 , n276232 , n276233 , n276234 , n276235 , n276236 , 
     n276237 , n276238 , n276239 , n276240 , n276241 , n276242 , n276243 , n276244 , n276245 , n276246 , 
     n276247 , n276248 , n276249 , n276250 , n276251 , n276252 , n276253 , n276254 , n276255 , n276256 , 
     n276257 , n276258 , n276259 , n276260 , n276261 , n276262 , n276263 , n276264 , n276265 , n276266 , 
     n276267 , n276268 , n276269 , n276270 , n276271 , n276272 , n276273 , n276274 , n276275 , n276276 , 
     n276277 , n276278 , n276279 , n276280 , n276281 , n276282 , n276283 , n276284 , n276285 , n276286 , 
     n276287 , n276288 , n276289 , n276290 , n276291 , n276292 , n276293 , n276294 , n276295 , n276296 , 
     n276297 , n276298 , n276299 , n276300 , n276301 , n276302 , n276303 , n276304 , n276305 , n276306 , 
     n276307 , n276308 , n276309 , n276310 , n276311 , n276312 , n276313 , n276314 , n276315 , n276316 , 
     n276317 , n276318 , n276319 , n276320 , n276321 , n276322 , n276323 , n276324 , n276325 , n276326 , 
     n276327 , n276328 , n276329 , n276330 , n276331 , n276332 , n276333 , n276334 , n276335 , n276336 , 
     n276337 , n276338 , n276339 , n276340 , n276341 , n276342 , n276343 , n276344 , n276345 , n276346 , 
     n276347 , n276348 , n276349 , n276350 , n276351 , n276352 , n276353 , n276354 , n276355 , n276356 , 
     n276357 , n276358 , n276359 , n276360 , n276361 , n276362 , n276363 , n276364 , n276365 , n276366 , 
     n276367 , n276368 , n276369 , n276370 , n276371 , n276372 , n276373 , n276374 , n276375 , n276376 , 
     n276377 , n276378 , n276379 , n276380 , n276381 , n276382 , n276383 , n276384 , n276385 , n276386 , 
     n276387 , n276388 , n276389 , n276390 , n276391 , n276392 , n276393 , n276394 , n276395 , n276396 , 
     n276397 , n276398 , n276399 , n276400 , n276401 , n276402 , n276403 , n276404 , n276405 , n276406 , 
     n276407 , n276408 , n276409 , n276410 , n276411 , n276412 , n276413 , n276414 , n276415 , n276416 , 
     n276417 , n276418 , n276419 , n276420 , n276421 , n276422 , n276423 , n276424 , n276425 , n276426 , 
     n276427 , n276428 , n276429 , n276430 , n276431 , n276432 , n276433 , n276434 , n276435 , n276436 , 
     n276437 , n276438 , n276439 , n276440 , n276441 , n276442 , n276443 , n276444 , n276445 , n276446 , 
     n276447 , n276448 , n276449 , n276450 , n276451 , n276452 , n276453 , n276454 , n276455 , n276456 , 
     n276457 , n276458 , n276459 , n276460 , n276461 , n276462 , n276463 , n276464 , n276465 , n276466 , 
     n276467 , n276468 , n276469 , n276470 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , 
     n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , 
     n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , 
     n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , 
     n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , 
     n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , 
     n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , 
     n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , 
     n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , 
     n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , 
     n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , 
     n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , 
     n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , 
     n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , 
     n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , 
     n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , 
     n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , 
     n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , 
     n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , 
     n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , 
     n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , 
     n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , 
     n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , 
     n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , 
     n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , 
     n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , 
     n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , 
     n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , 
     n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , 
     n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , 
     n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , 
     n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , 
     n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , 
     n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , 
     n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , 
     n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , 
     n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , 
     n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , 
     n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , 
     n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , 
     n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , 
     n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , 
     n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , 
     n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , 
     n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , 
     n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , 
     n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , 
     n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , 
     n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , 
     n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , 
     n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , 
     n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , 
     n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , 
     n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , 
     n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , 
     n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , 
     n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , 
     n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , 
     n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , 
     n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , 
     n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , 
     n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , 
     n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , 
     n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , 
     n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , 
     n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , 
     n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , 
     n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , 
     n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , 
     n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , 
     n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , 
     n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , 
     n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , 
     n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , 
     n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , 
     n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , 
     n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , 
     n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , 
     n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , 
     n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , 
     n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n277273 , n277274 , n277275 , n277276 , 
     n277277 , n277278 , n277279 , n277280 , n277281 , n277282 , n277283 , n277284 , n277285 , n277286 , 
     n277287 , n277288 , n277289 , n277290 , n277291 , n277292 , n277293 , n277294 , n277295 , n277296 , 
     n277297 , n277298 , n277299 , n277300 , n277301 , n277302 , n277303 , n277304 , n277305 , n277306 , 
     n277307 , n277308 , n277309 , n277310 , n277311 , n277312 , n277313 , n277314 , n277315 , n277316 , 
     n277317 , n277318 , n277319 , n277320 , n277321 , n277322 , n277323 , n277324 , n277325 , n277326 , 
     n277327 , n277328 , n277329 , n277330 , n277331 , n277332 , n277333 , n277334 , n277335 , n277336 , 
     n277337 , n277338 , n277339 , n277340 , n277341 , n277342 , n277343 , n277344 , n277345 , n277346 , 
     n277347 , n277348 , n277349 , n277350 , n277351 , n277352 , n277353 , n277354 , n277355 , n277356 , 
     n277357 , n277358 , n277359 , n277360 , n277361 , n277362 , n277363 , n277364 , n277365 , n277366 , 
     n277367 , n277368 , n277369 , n277370 , n277371 , n277372 , n277373 , n277374 , n277375 , n277376 , 
     n277377 , n277378 , n277379 , n277380 , n277381 , n277382 , n277383 , n277384 , n277385 , n277386 , 
     n277387 , n277388 , n277389 , n277390 , n277391 , n277392 , n277393 , n277394 , n277395 , n277396 , 
     n277397 , n277398 , n277399 , n277400 , n277401 , n277402 , n277403 , n277404 , n277405 , n277406 , 
     n277407 , n277408 , n277409 , n277410 , n277411 , n277412 , n277413 , n277414 , n277415 , n277416 , 
     n277417 , n277418 , n277419 , n277420 , n277421 , n277422 , n277423 , n277424 , n277425 , n277426 , 
     n277427 , n277428 , n277429 , n277430 , n277431 , n277432 , n277433 , n277434 , n277435 , n277436 , 
     n277437 , n277438 , n277439 , n277440 , n277441 , n277442 , n277443 , n277444 , n277445 , n277446 , 
     n277447 , n277448 , n277449 , n277450 , n277451 , n277452 , n277453 , n277454 , n277455 , n277456 , 
     n277457 , n277458 , n277459 , n277460 , n277461 , n277462 , n277463 , n277464 , n277465 , n277466 , 
     n277467 , n277468 , n277469 , n277470 , n277471 , n277472 , n277473 , n277474 , n277475 , n277476 , 
     n277477 , n277478 , n277479 , n277480 , n277481 , n277482 , n277483 , n277484 , n277485 , n277486 , 
     n277487 , n277488 , n277489 , n277490 , n277491 , n277492 , n277493 , n277494 , n277495 , n277496 , 
     n277497 , n277498 , n277499 , n277500 , n277501 , n277502 , n277503 , n277504 , n277505 , n277506 , 
     n277507 , n277508 , n277509 , n277510 , n277511 , n277512 , n277513 , n277514 , n277515 , n277516 , 
     n277517 , n277518 , n277519 , n277520 , n277521 , n277522 , n277523 , n277524 , n277525 , n277526 , 
     n277527 , n277528 , n277529 , n277530 , n277531 , n277532 , n277533 , n277534 , n277535 , n277536 , 
     n277537 , n277538 , n277539 , n277540 , n277541 , n277542 , n277543 , n277544 , n277545 , n277546 , 
     n277547 , n277548 , n277549 , n277550 , n277551 , n277552 , n277553 , n277554 , n277555 , n277556 , 
     n277557 , n277558 , n277559 , n277560 , n277561 , n277562 , n277563 , n277564 , n277565 , n277566 , 
     n277567 , n277568 , n277569 , n277570 , n277571 , n277572 , n277573 , n277574 , n277575 , n277576 , 
     n277577 , n277578 , n277579 , n277580 , n277581 , n277582 , n277583 , n277584 , n277585 , n277586 , 
     n277587 , n277588 , n277589 , n277590 , n277591 , n277592 , n277593 , n277594 , n277595 , n277596 , 
     n277597 , n277598 , n277599 , n277600 , n277601 , n277602 , n277603 , n277604 , n277605 , n277606 , 
     n277607 , n277608 , n277609 , n277610 , n277611 , n277612 , n277613 , n277614 , n277615 , n277616 , 
     n277617 , n277618 , n277619 , n277620 , n277621 , n277622 , n277623 , n277624 , n277625 , n277626 , 
     n277627 , n277628 , n277629 , n277630 , n277631 , n277632 , n277633 , n277634 , n277635 , n277636 , 
     n277637 , n277638 , n277639 , n277640 , n277641 , n277642 , n277643 , n277644 , n277645 , n277646 , 
     n277647 , n277648 , n277649 , n277650 , n277651 , n277652 , n277653 , n277654 , n277655 , n277656 , 
     n277657 , n277658 , n277659 , n277660 , n277661 , n277662 , n277663 , n277664 , n277665 , n277666 , 
     n277667 , n277668 , n277669 , n277670 , n277671 , n277672 , n277673 , n277674 , n277675 , n277676 , 
     n277677 , n277678 , n277679 , n277680 , n277681 , n277682 , n277683 , n277684 , n277685 , n277686 , 
     n277687 , n277688 , n277689 , n277690 , n277691 , n277692 , n277693 , n277694 , n277695 , n277696 , 
     n277697 , n277698 , n277699 , n277700 , n277701 , n277702 , n277703 , n277704 , n277705 , n277706 , 
     n277707 , n277708 , n277709 , n277710 , n277711 , n277712 , n277713 , n277714 , n277715 , n277716 , 
     n277717 , n277718 , n277719 , n277720 , n277721 , n277722 , n277723 , n277724 , n277725 , n277726 , 
     n277727 , n277728 , n277729 , n277730 , n277731 , n277732 , n277733 , n277734 , n277735 , n277736 , 
     n277737 , n277738 , n277739 , n277740 , n277741 , n277742 , n277743 , n277744 , n277745 , n277746 , 
     n277747 , n277748 , n277749 , n277750 , n277751 , n277752 , n277753 , n277754 , n277755 , n277756 , 
     n277757 , n277758 , n277759 , n277760 , n277761 , n277762 , n277763 , n277764 , n277765 , n277766 , 
     n277767 , n277768 , n277769 , n277770 , n277771 , n277772 , n277773 , n277774 , n277775 , n277776 , 
     n277777 , n277778 , n277779 , n277780 , n277781 , n277782 , n277783 , n277784 , n277785 , n277786 , 
     n277787 , n277788 , n277789 , n277790 , n277791 , n277792 , n277793 , n277794 , n277795 , n277796 , 
     n277797 , n277798 , n277799 , n277800 , n277801 , n277802 , n277803 , n277804 , n277805 , n277806 , 
     n277807 , n277808 , n277809 , n277810 , n277811 , n277812 , n277813 , n277814 , n277815 , n277816 , 
     n277817 , n277818 , n277819 , n277820 , n277821 , n277822 , n277823 , n277824 , n277825 , n277826 , 
     n277827 , n277828 , n277829 , n277830 , n277831 , n277832 , n277833 , n277834 , n277835 , n277836 , 
     n277837 , n277838 , n277839 , n277840 , n277841 , n277842 , n277843 , n277844 , n277845 , n277846 , 
     n277847 , n277848 , n277849 , n277850 , n277851 , n277852 , n277853 , n277854 , n277855 , n277856 , 
     n277857 , n277858 , n277859 , n277860 , n277861 , n277862 , n277863 , n277864 , n277865 , n277866 , 
     n277867 , n277868 , n277869 , n277870 , n277871 , n277872 , n277873 , n277874 , n277875 , n277876 , 
     n277877 , n277878 , n277879 , n277880 , n277881 , n277882 , n277883 , n277884 , n277885 , n277886 , 
     n277887 , n277888 , n277889 , n277890 , n277891 , n277892 , n277893 , n277894 , n277895 , n277896 , 
     n277897 , n277898 , n277899 , n277900 , n277901 , n277902 , n277903 , n277904 , n277905 , n277906 , 
     n277907 , n277908 , n277909 , n277910 , n277911 , n277912 , n277913 , n277914 , n277915 , n277916 , 
     n277917 , n277918 , n277919 , n277920 , n277921 , n277922 , n277923 , n277924 , n277925 , n277926 , 
     n277927 , n277928 , n277929 , n277930 , n277931 , n277932 , n277933 , n277934 , n277935 , n277936 , 
     n277937 , n277938 , n277939 , n277940 , n277941 , n277942 , n277943 , n277944 , n277945 , n277946 , 
     n277947 , n277948 , n277949 , n277950 , n277951 , n277952 , n277953 , n277954 , n277955 , n277956 , 
     n277957 , n277958 , n277959 , n277960 , n277961 , n277962 , n277963 , n277964 , n277965 , n277966 , 
     n277967 , n277968 , n277969 , n277970 , n277971 , n277972 , n277973 , n277974 , n277975 , n277976 , 
     n277977 , n277978 , n277979 , n277980 , n277981 , n277982 , n277983 , n277984 , n277985 , n277986 , 
     n277987 , n277988 , n277989 , n277990 , n277991 , n277992 , n277993 , n277994 , n277995 , n277996 , 
     n277997 , n277998 , n277999 , n278000 , n278001 , n278002 , n278003 , n278004 , n278005 , n278006 , 
     n278007 , n278008 , n278009 , n278010 , n278011 , n278012 , n278013 , n278014 , n278015 , n278016 , 
     n278017 , n278018 , n278019 , n278020 , n278021 , n278022 , n278023 , n278024 , n278025 , n278026 , 
     n278027 , n278028 , n278029 , n278030 , n278031 , n278032 , n278033 , n278034 , n278035 , n278036 , 
     n278037 , n278038 , n278039 , n278040 , n278041 , n278042 , n278043 , n278044 , n278045 , n278046 , 
     n278047 , n278048 , n278049 , n278050 , n278051 , n278052 , n278053 , n278054 , n278055 , n278056 , 
     n278057 , n278058 , n278059 , n278060 , n278061 , n278062 , n278063 , n278064 , n278065 , n278066 , 
     n278067 , n278068 , n278069 , n278070 , n278071 , n278072 , n278073 , n278074 , n278075 , n10613 , 
     n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , 
     n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , 
     n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , 
     n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , 
     n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , 
     n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , 
     n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , 
     n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , 
     n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , 
     n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , 
     n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , 
     n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , 
     n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , 
     n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , 
     n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , 
     n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , 
     n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , 
     n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , 
     n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , 
     n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , 
     n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , 
     n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , 
     n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , 
     n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , 
     n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , 
     n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , 
     n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , 
     n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , 
     n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , 
     n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , 
     n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , 
     n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , 
     n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , 
     n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , 
     n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , 
     n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , 
     n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , 
     n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , 
     n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , 
     n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , 
     n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , 
     n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , 
     n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , 
     n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , 
     n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , 
     n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , 
     n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , 
     n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , 
     n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , 
     n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , 
     n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , 
     n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , 
     n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , 
     n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , 
     n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , 
     n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , 
     n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , 
     n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , 
     n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , 
     n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , 
     n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , 
     n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , 
     n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , 
     n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , 
     n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , 
     n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , 
     n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , 
     n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , 
     n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , 
     n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , 
     n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , 
     n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , 
     n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , 
     n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , 
     n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , 
     n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , 
     n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , 
     n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , 
     n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , 
     n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , 
     n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , 
     n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , 
     n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , 
     n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , 
     n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , 
     n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , 
     n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , 
     n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , 
     n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , 
     n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , 
     n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , 
     n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , 
     n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , 
     n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , 
     n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , 
     n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , 
     n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , 
     n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , 
     n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , 
     n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , 
     n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , 
     n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , 
     n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , 
     n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , 
     n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , 
     n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , 
     n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , 
     n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , 
     n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , 
     n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , 
     n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , 
     n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , 
     n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , 
     n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , 
     n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , 
     n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , 
     n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , 
     n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , 
     n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , 
     n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , 
     n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , 
     n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , 
     n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , 
     n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , 
     n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , 
     n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , 
     n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , 
     n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , 
     n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , 
     n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , 
     n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , 
     n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , 
     n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , 
     n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , 
     n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , 
     n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , 
     n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , 
     n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , 
     n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , 
     n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , 
     n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , 
     n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , 
     n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , 
     n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , 
     n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , 
     n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , 
     n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , 
     n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , 
     n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , 
     n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , 
     n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , 
     n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , 
     n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , 
     n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , 
     n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , 
     n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , 
     n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , 
     n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , 
     n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , 
     n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , 
     n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , 
     n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , 
     n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , 
     n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , 
     n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , 
     n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , 
     n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , 
     n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , 
     n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , 
     n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , 
     n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , 
     n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , 
     n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , 
     n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , 
     n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , 
     n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , 
     n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , 
     n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , 
     n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , 
     n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , 
     n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , 
     n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , 
     n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , 
     n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , 
     n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , 
     n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , 
     n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , 
     n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , 
     n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , 
     n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , 
     n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , 
     n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , 
     n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , 
     n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , 
     n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , 
     n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , 
     n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , 
     n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , 
     n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , 
     n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , 
     n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , 
     n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , 
     n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , 
     n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , 
     n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , 
     n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , 
     n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , 
     n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , 
     n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , 
     n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , 
     n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , 
     n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , 
     n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , 
     n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , 
     n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , 
     n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , 
     n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , 
     n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , 
     n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , 
     n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , 
     n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , 
     n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , 
     n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , 
     n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , 
     n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , 
     n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , 
     n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , 
     n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , 
     n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , 
     n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , 
     n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , 
     n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , 
     n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , 
     n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , 
     n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , 
     n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , 
     n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , 
     n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , 
     n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , 
     n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , 
     n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , 
     n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , 
     n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , 
     n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , 
     n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , 
     n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , 
     n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , 
     n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , 
     n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , 
     n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , 
     n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , 
     n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , 
     n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , 
     n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , 
     n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , 
     n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , 
     n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , 
     n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , 
     n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , 
     n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , 
     n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , 
     n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , 
     n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , 
     n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , 
     n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , 
     n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , 
     n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , 
     n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , 
     n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , 
     n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , 
     n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , 
     n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , 
     n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , 
     n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , 
     n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , 
     n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , 
     n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , 
     n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , 
     n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , 
     n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , 
     n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , 
     n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , 
     n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , 
     n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , 
     n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , 
     n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , 
     n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , 
     n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , 
     n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , 
     n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , 
     n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , 
     n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , 
     n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , 
     n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , 
     n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , 
     n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , 
     n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , 
     n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , 
     n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , 
     n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , 
     n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , 
     n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , 
     n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , 
     n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , 
     n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , 
     n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , 
     n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , 
     n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , 
     n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , 
     n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , 
     n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , 
     n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , 
     n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , 
     n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , 
     n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , 
     n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , 
     n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , 
     n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , 
     n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , 
     n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , 
     n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , 
     n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , 
     n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , 
     n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , 
     n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , 
     n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , 
     n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , 
     n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , 
     n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , 
     n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , 
     n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , 
     n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , 
     n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , 
     n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , 
     n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , 
     n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , 
     n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , 
     n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , 
     n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , 
     n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , 
     n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , 
     n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , 
     n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , 
     n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , 
     n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , 
     n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , 
     n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , 
     n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , 
     n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , 
     n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , 
     n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , 
     n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , 
     n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , 
     n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , 
     n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , 
     n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , 
     n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , 
     n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , 
     n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , 
     n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , 
     n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , 
     n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , 
     n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , 
     n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , 
     n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , 
     n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , 
     n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , 
     n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , 
     n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , 
     n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , 
     n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , 
     n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , 
     n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , 
     n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , 
     n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , 
     n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , 
     n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , 
     n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , 
     n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , 
     n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , 
     n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , 
     n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , 
     n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , 
     n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , 
     n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , 
     n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , 
     n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , 
     n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , 
     n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , 
     n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , 
     n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , 
     n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , 
     n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , 
     n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , 
     n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , 
     n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , 
     n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , 
     n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , 
     n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , 
     n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , 
     n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , 
     n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , 
     n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , 
     n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , 
     n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , 
     n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , 
     n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , 
     n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , 
     n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , 
     n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , 
     n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , 
     n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , 
     n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , 
     n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , 
     n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , 
     n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , 
     n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , 
     n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , 
     n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , 
     n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , 
     n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , 
     n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , 
     n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , 
     n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , 
     n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , 
     n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , 
     n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , 
     n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , 
     n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , 
     n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , 
     n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , 
     n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , 
     n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , 
     n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , 
     n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , 
     n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , 
     n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , 
     n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , 
     n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , 
     n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , 
     n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , 
     n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , 
     n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , 
     n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , 
     n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , 
     n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , 
     n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , 
     n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , 
     n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , 
     n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , 
     n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , 
     n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , 
     n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , 
     n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , 
     n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , 
     n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , 
     n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , 
     n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , 
     n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , 
     n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , 
     n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , 
     n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , 
     n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , 
     n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , 
     n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , 
     n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , 
     n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , 
     n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , 
     n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , 
     n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , 
     n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , 
     n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , 
     n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , 
     n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , 
     n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , 
     n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , 
     n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , 
     n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , 
     n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , 
     n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , 
     n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , 
     n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , 
     n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , 
     n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , 
     n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , 
     n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , 
     n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , 
     n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , 
     n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , 
     n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , 
     n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , 
     n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , 
     n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , 
     n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , 
     n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , 
     n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , 
     n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , 
     n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , 
     n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , 
     n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , 
     n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , 
     n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , 
     n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , 
     n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , 
     n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , 
     n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , 
     n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , 
     n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , 
     n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , 
     n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , 
     n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , 
     n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , 
     n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , 
     n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , 
     n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , 
     n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , 
     n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , 
     n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , 
     n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , 
     n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , 
     n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , 
     n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , 
     n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , 
     n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , 
     n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , 
     n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , 
     n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , 
     n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , 
     n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , 
     n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , 
     n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , 
     n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , 
     n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , 
     n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , 
     n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , 
     n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , 
     n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , 
     n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , 
     n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , 
     n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , 
     n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , 
     n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , 
     n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , 
     n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , 
     n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , 
     n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , 
     n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , 
     n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , 
     n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , 
     n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , 
     n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , 
     n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , 
     n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , 
     n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , 
     n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , 
     n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , 
     n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , 
     n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , 
     n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , 
     n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , 
     n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , 
     n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , 
     n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , 
     n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , 
     n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , 
     n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , 
     n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , 
     n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , 
     n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , 
     n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , 
     n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , 
     n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , 
     n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , 
     n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , 
     n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , 
     n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , 
     n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , 
     n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , 
     n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , 
     n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , 
     n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , 
     n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , 
     n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , 
     n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , 
     n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , 
     n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , 
     n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , 
     n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , 
     n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , 
     n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , 
     n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , 
     n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , 
     n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , 
     n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , 
     n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , 
     n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , 
     n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , 
     n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , 
     n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , 
     n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , 
     n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , 
     n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , 
     n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , 
     n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , 
     n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , 
     n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , 
     n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , 
     n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , 
     n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , 
     n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , 
     n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , 
     n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , 
     n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , 
     n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , 
     n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , 
     n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , 
     n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , 
     n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , 
     n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , 
     n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , 
     n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , 
     n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , 
     n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , 
     n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , 
     n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , 
     n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , 
     n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , 
     n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , 
     n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , 
     n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , 
     n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , 
     n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , 
     n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , 
     n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , 
     n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , 
     n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , 
     n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , 
     n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , 
     n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , 
     n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , 
     n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , 
     n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , 
     n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , 
     n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , 
     n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , 
     n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , 
     n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , 
     n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , 
     n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , 
     n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , 
     n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , 
     n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , 
     n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , 
     n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , 
     n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , 
     n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , 
     n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , 
     n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , 
     n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , 
     n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , 
     n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , 
     n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , 
     n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , 
     n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , 
     n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , 
     n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , 
     n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , 
     n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , 
     n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , 
     n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , 
     n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , 
     n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , 
     n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , 
     n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , 
     n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , 
     n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , 
     n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , 
     n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , 
     n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , 
     n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , 
     n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , 
     n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , 
     n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , 
     n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , 
     n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , 
     n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , 
     n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , 
     n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , 
     n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , 
     n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , 
     n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , 
     n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , 
     n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , 
     n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , 
     n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , 
     n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , 
     n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , 
     n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , 
     n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , 
     n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , 
     n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , 
     n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , 
     n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , 
     n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , 
     n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , 
     n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , 
     n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , 
     n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , 
     n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , 
     n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , 
     n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , 
     n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , 
     n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , 
     n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , 
     n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , 
     n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , 
     n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , 
     n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , 
     n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , 
     n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , 
     n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , 
     n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , 
     n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , 
     n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , 
     n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , 
     n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , 
     n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , 
     n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , 
     n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , 
     n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , 
     n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , 
     n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , 
     n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , 
     n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , 
     n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , 
     n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , 
     n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , 
     n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , 
     n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , 
     n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , 
     n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , 
     n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , 
     n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , 
     n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , 
     n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , 
     n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , 
     n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , 
     n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , 
     n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , 
     n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , 
     n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , 
     n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , 
     n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , 
     n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , 
     n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , 
     n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , 
     n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , 
     n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , 
     n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , 
     n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , 
     n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , 
     n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , 
     n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , 
     n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , 
     n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , 
     n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , 
     n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , 
     n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , 
     n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , 
     n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , 
     n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , 
     n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , 
     n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , 
     n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , 
     n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , 
     n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , 
     n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , 
     n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , 
     n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , 
     n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , 
     n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , 
     n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , 
     n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , 
     n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , 
     n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , 
     n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , 
     n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , 
     n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , 
     n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , 
     n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , 
     n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , 
     n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , 
     n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , 
     n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , 
     n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , 
     n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , 
     n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , 
     n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , 
     n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , 
     n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , 
     n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , 
     n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , 
     n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , 
     n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , 
     n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , 
     n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , 
     n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , 
     n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , 
     n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , 
     n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , 
     n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , 
     n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , 
     n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , 
     n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , 
     n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , 
     n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , 
     n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , 
     n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , 
     n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , 
     n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , 
     n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , 
     n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , 
     n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , 
     n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , 
     n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , 
     n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , 
     n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , 
     n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , 
     n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , 
     n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , 
     n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , 
     n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , 
     n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , 
     n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , 
     n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , 
     n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , 
     n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , 
     n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , 
     n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , 
     n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , 
     n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , 
     n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , 
     n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , 
     n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , 
     n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , 
     n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , 
     n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , 
     n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , 
     n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , 
     n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , 
     n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , 
     n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , 
     n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , 
     n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , 
     n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , 
     n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , 
     n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , 
     n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , 
     n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , 
     n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , 
     n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , 
     n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , 
     n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , 
     n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , 
     n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , 
     n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , 
     n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , 
     n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , 
     n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , 
     n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , 
     n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , 
     n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , 
     n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , 
     n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , 
     n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , 
     n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , 
     n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , 
     n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , 
     n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , 
     n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , 
     n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , 
     n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , 
     n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , 
     n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , 
     n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , 
     n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , 
     n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , 
     n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , 
     n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , 
     n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , 
     n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , 
     n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , 
     n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , 
     n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , 
     n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , 
     n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , 
     n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , 
     n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , 
     n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , 
     n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , 
     n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , 
     n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , 
     n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , 
     n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , 
     n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , 
     n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , 
     n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , 
     n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , 
     n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , 
     n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , 
     n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , 
     n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , 
     n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , 
     n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , 
     n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , 
     n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , 
     n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , 
     n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , 
     n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , 
     n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , 
     n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , 
     n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , 
     n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , 
     n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , 
     n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , 
     n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , 
     n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , 
     n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , 
     n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , 
     n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , 
     n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , 
     n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , 
     n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , 
     n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , 
     n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , 
     n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , 
     n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , 
     n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , 
     n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , 
     n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , 
     n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , 
     n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , 
     n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , 
     n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , 
     n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , 
     n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , 
     n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , 
     n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , 
     n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , 
     n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , 
     n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , 
     n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , 
     n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , 
     n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , 
     n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , 
     n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , 
     n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , 
     n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , 
     n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , 
     n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , 
     n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , 
     n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , 
     n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , 
     n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , 
     n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , 
     n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , 
     n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , 
     n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , 
     n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , 
     n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , 
     n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , 
     n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , 
     n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , 
     n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , 
     n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , 
     n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , 
     n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , 
     n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , 
     n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , 
     n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , 
     n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , 
     n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , 
     n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , 
     n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , 
     n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , 
     n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , 
     n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , 
     n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , 
     n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , 
     n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , 
     n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , 
     n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , 
     n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , 
     n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , 
     n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , 
     n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , 
     n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , 
     n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , 
     n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , 
     n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , 
     n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , 
     n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , 
     n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , 
     n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , 
     n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , 
     n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , 
     n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , 
     n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , 
     n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , 
     n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , 
     n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , 
     n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , 
     n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , 
     n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , 
     n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , 
     n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , 
     n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , 
     n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , 
     n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , 
     n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , 
     n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , 
     n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , 
     n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , 
     n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , 
     n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , 
     n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , 
     n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , 
     n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , 
     n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , 
     n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , 
     n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , 
     n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , 
     n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , 
     n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , 
     n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , 
     n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , 
     n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , 
     n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , 
     n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , 
     n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , 
     n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , 
     n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , 
     n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , 
     n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , 
     n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , 
     n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , 
     n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , 
     n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , 
     n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , 
     n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , 
     n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , 
     n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , 
     n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , 
     n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , 
     n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , 
     n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , 
     n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , 
     n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , 
     n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , 
     n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , 
     n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , 
     n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , 
     n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , 
     n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , 
     n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , 
     n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , 
     n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , 
     n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , 
     n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , 
     n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , 
     n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , 
     n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , 
     n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , 
     n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , 
     n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , 
     n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , 
     n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , 
     n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , 
     n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , 
     n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , 
     n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , 
     n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , 
     n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , 
     n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , 
     n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , 
     n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , 
     n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , 
     n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , 
     n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , 
     n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , 
     n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , 
     n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , 
     n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , 
     n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , 
     n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , 
     n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , 
     n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , 
     n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , 
     n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , 
     n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , 
     n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , 
     n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , 
     n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , 
     n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , 
     n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , 
     n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , 
     n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , 
     n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , 
     n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , 
     n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , 
     n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , 
     n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , 
     n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , 
     n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , 
     n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , 
     n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , 
     n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , 
     n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , 
     n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , 
     n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , 
     n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , 
     n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , 
     n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , 
     n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , 
     n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , 
     n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , 
     n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , 
     n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , 
     n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , 
     n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , 
     n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , 
     n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , 
     n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , 
     n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , 
     n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , 
     n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , 
     n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , 
     n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , 
     n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , 
     n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , 
     n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , 
     n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , 
     n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , 
     n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , 
     n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , 
     n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , 
     n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , 
     n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , 
     n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , 
     n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , 
     n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , 
     n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , 
     n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , 
     n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , 
     n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , 
     n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , 
     n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , 
     n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , 
     n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , 
     n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , 
     n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , 
     n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , 
     n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , 
     n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , 
     n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , 
     n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , 
     n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , 
     n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , 
     n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , 
     n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , 
     n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , 
     n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , 
     n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , 
     n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , 
     n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , 
     n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , 
     n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , 
     n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , 
     n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , 
     n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , 
     n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , 
     n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , 
     n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , 
     n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , 
     n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , 
     n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , 
     n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , 
     n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , 
     n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , 
     n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , 
     n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , 
     n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , 
     n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , 
     n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , 
     n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , 
     n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , 
     n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , 
     n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , 
     n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , 
     n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , 
     n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , 
     n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , 
     n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , 
     n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , 
     n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , 
     n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , 
     n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , 
     n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , 
     n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , 
     n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , 
     n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , 
     n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , 
     n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , 
     n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , 
     n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , 
     n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , 
     n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , 
     n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , 
     n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , 
     n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , 
     n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , 
     n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , 
     n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , 
     n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , 
     n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , 
     n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , 
     n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , 
     n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , 
     n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , 
     n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , 
     n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , 
     n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , 
     n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , 
     n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , 
     n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , 
     n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , 
     n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , 
     n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , 
     n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , 
     n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , 
     n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , 
     n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , 
     n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , 
     n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , 
     n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , 
     n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , 
     n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , 
     n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , 
     n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , 
     n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , 
     n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , 
     n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , 
     n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , 
     n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , 
     n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , 
     n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , 
     n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , 
     n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , 
     n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , 
     n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , 
     n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , 
     n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , 
     n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , 
     n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , 
     n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , 
     n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , 
     n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , 
     n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , 
     n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , 
     n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , 
     n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , 
     n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , 
     n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , 
     n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , 
     n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , 
     n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , 
     n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , 
     n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , 
     n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , 
     n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , 
     n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , 
     n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , 
     n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , 
     n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , 
     n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , 
     n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , 
     n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , 
     n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , 
     n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , 
     n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , 
     n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , 
     n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , 
     n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , 
     n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , 
     n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , 
     n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , 
     n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , 
     n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , 
     n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , 
     n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , 
     n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , 
     n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , 
     n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , 
     n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , 
     n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , 
     n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , 
     n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , 
     n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , 
     n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , 
     n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , 
     n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , 
     n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , 
     n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , 
     n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , 
     n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , 
     n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , 
     n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , 
     n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , 
     n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , 
     n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , 
     n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , 
     n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , 
     n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , 
     n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , 
     n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , 
     n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , 
     n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , 
     n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , 
     n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , 
     n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , 
     n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , 
     n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , 
     n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , 
     n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , 
     n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , 
     n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , 
     n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , 
     n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , 
     n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , 
     n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , 
     n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , 
     n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , 
     n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , 
     n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , 
     n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , 
     n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , 
     n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , 
     n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , 
     n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , 
     n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , 
     n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , 
     n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , 
     n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , 
     n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , 
     n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , 
     n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , 
     n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , 
     n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , 
     n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , 
     n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , 
     n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , 
     n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , 
     n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , 
     n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , 
     n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , 
     n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , 
     n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , 
     n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , 
     n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , 
     n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , 
     n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , 
     n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , 
     n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , 
     n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , 
     n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , 
     n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , 
     n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , 
     n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , 
     n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , 
     n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , 
     n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , 
     n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , 
     n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , 
     n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , 
     n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , 
     n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , 
     n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , 
     n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , 
     n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , 
     n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , 
     n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , 
     n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , 
     n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , 
     n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , 
     n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , 
     n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , 
     n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , 
     n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , 
     n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , 
     n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , 
     n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , 
     n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , 
     n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , 
     n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , 
     n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , 
     n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , 
     n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , 
     n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , 
     n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , 
     n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , 
     n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , 
     n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , 
     n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , 
     n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , 
     n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , 
     n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , 
     n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , 
     n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , 
     n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , 
     n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , 
     n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , 
     n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , 
     n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , 
     n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , 
     n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , 
     n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , 
     n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , 
     n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , 
     n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , 
     n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , 
     n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , 
     n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , 
     n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , 
     n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , 
     n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , 
     n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , 
     n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , 
     n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , 
     n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , 
     n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , 
     n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , 
     n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , 
     n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , 
     n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , 
     n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , 
     n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , 
     n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , 
     n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , 
     n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , 
     n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , 
     n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , 
     n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , 
     n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , 
     n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , 
     n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , 
     n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , 
     n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , 
     n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , 
     n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , 
     n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , 
     n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , 
     n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , 
     n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , 
     n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , 
     n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , 
     n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , 
     n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , 
     n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , 
     n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , 
     n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , 
     n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , 
     n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , 
     n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , 
     n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , 
     n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , 
     n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , 
     n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , 
     n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , 
     n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , 
     n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , 
     n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , 
     n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , 
     n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , 
     n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , 
     n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , 
     n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , 
     n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , 
     n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , 
     n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , 
     n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , 
     n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , 
     n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , 
     n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , 
     n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , 
     n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , 
     n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , 
     n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , 
     n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , 
     n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , 
     n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , 
     n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , 
     n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , 
     n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , 
     n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , 
     n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , 
     n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , 
     n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , 
     n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , 
     n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , 
     n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , 
     n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , 
     n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , 
     n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , 
     n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , 
     n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , 
     n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , 
     n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , 
     n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , 
     n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , 
     n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , 
     n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , 
     n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , 
     n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , 
     n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , 
     n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , 
     n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , 
     n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , 
     n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , 
     n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , 
     n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , 
     n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , 
     n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , 
     n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , 
     n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , 
     n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , 
     n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , 
     n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , 
     n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , 
     n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , 
     n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , 
     n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , 
     n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , 
     n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , 
     n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , 
     n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , 
     n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , 
     n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , 
     n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , 
     n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , 
     n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , 
     n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , 
     n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , 
     n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , 
     n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , 
     n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , 
     n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , 
     n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , 
     n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , 
     n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , 
     n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , 
     n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , 
     n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , 
     n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , 
     n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , 
     n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , 
     n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , 
     n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , 
     n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , 
     n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , 
     n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , 
     n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , 
     n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , 
     n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , 
     n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , 
     n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , 
     n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , 
     n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , 
     n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , 
     n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , 
     n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , 
     n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , 
     n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , 
     n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , 
     n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , 
     n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , 
     n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , 
     n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , 
     n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , 
     n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , 
     n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , 
     n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , 
     n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , 
     n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , 
     n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , 
     n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , 
     n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , 
     n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , 
     n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , 
     n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , 
     n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , 
     n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , 
     n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , 
     n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , 
     n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , 
     n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , 
     n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , 
     n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , 
     n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , 
     n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , 
     n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , 
     n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , 
     n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , 
     n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , 
     n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , 
     n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , 
     n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , 
     n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , 
     n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , 
     n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , 
     n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , 
     n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , 
     n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , 
     n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , 
     n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , 
     n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , 
     n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , 
     n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , 
     n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , 
     n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , 
     n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , 
     n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , 
     n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , 
     n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , 
     n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , 
     n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , 
     n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , 
     n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , 
     n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , 
     n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , 
     n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , 
     n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , 
     n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , 
     n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , 
     n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , 
     n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , 
     n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , 
     n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , 
     n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , 
     n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , 
     n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , 
     n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , 
     n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , 
     n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , 
     n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , 
     n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , 
     n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , 
     n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , 
     n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , 
     n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , 
     n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , 
     n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , 
     n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , 
     n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , 
     n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , 
     n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , 
     n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , 
     n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , 
     n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , 
     n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , 
     n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , 
     n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , 
     n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , 
     n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , 
     n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , 
     n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , 
     n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , 
     n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , 
     n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , 
     n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , 
     n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , 
     n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , 
     n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , 
     n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , 
     n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , 
     n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , 
     n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , 
     n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , 
     n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , 
     n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , 
     n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , 
     n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , 
     n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , 
     n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , 
     n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , 
     n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , 
     n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , 
     n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , 
     n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , 
     n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , 
     n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , 
     n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , 
     n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , 
     n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , 
     n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , 
     n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , 
     n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , 
     n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , 
     n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , 
     n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , 
     n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , 
     n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , 
     n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , 
     n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , 
     n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , 
     n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , 
     n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , 
     n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , 
     n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , 
     n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , 
     n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , 
     n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , 
     n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , 
     n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , 
     n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , 
     n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , 
     n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , 
     n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , 
     n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , 
     n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , 
     n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , 
     n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , 
     n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , 
     n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , 
     n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , 
     n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , 
     n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , 
     n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , 
     n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , 
     n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , 
     n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , 
     n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , 
     n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , 
     n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , 
     n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , 
     n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , 
     n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , 
     n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , 
     n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , 
     n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , 
     n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , 
     n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , 
     n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , 
     n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , 
     n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , 
     n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , 
     n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , 
     n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , 
     n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , 
     n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , 
     n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , 
     n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , 
     n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , 
     n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , 
     n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , 
     n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , 
     n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , 
     n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , 
     n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , 
     n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , 
     n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , 
     n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , 
     n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , 
     n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , 
     n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , 
     n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , 
     n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , 
     n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , 
     n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , 
     n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , 
     n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , 
     n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , 
     n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , 
     n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , 
     n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , 
     n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , 
     n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , 
     n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , 
     n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , 
     n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , 
     n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , 
     n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , 
     n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , 
     n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , 
     n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , 
     n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , 
     n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , 
     n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , 
     n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , 
     n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , 
     n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , 
     n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , 
     n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , 
     n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , 
     n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , 
     n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , 
     n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , 
     n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , 
     n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , 
     n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , 
     n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , 
     n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , 
     n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , 
     n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , 
     n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , 
     n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , 
     n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , 
     n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , 
     n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , 
     n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , 
     n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , 
     n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , 
     n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , 
     n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , 
     n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , 
     n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , 
     n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , 
     n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , 
     n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , 
     n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , 
     n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , 
     n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , 
     n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , 
     n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , 
     n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , 
     n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , 
     n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , 
     n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , 
     n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , 
     n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , 
     n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , 
     n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , 
     n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , 
     n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , 
     n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , 
     n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , 
     n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , 
     n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , 
     n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , 
     n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , 
     n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , 
     n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , 
     n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , 
     n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , 
     n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , 
     n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , 
     n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , 
     n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , 
     n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , 
     n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , 
     n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , 
     n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , 
     n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , 
     n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , 
     n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , 
     n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , 
     n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , 
     n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , 
     n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , 
     n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , 
     n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , 
     n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , 
     n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , 
     n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , 
     n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , 
     n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , 
     n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , 
     n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , 
     n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , 
     n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , 
     n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , 
     n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , 
     n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , 
     n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , 
     n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , 
     n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , 
     n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , 
     n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , 
     n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , 
     n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , 
     n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , 
     n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , 
     n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , 
     n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , 
     n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , 
     n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , 
     n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , 
     n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , 
     n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , 
     n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , 
     n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , 
     n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , 
     n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , 
     n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , 
     n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , 
     n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , 
     n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , 
     n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , 
     n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , 
     n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , 
     n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , 
     n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , 
     n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , 
     n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , 
     n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , 
     n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , 
     n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , 
     n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , 
     n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , 
     n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , 
     n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , 
     n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , 
     n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , 
     n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , 
     n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , 
     n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , 
     n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , 
     n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , 
     n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , 
     n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , 
     n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , 
     n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , 
     n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , 
     n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , 
     n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , 
     n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , 
     n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , 
     n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , 
     n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , 
     n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , 
     n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , 
     n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , 
     n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , 
     n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , 
     n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , 
     n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , 
     n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , 
     n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , 
     n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , 
     n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , 
     n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , 
     n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , 
     n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , 
     n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , 
     n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , 
     n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , 
     n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , 
     n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , 
     n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , 
     n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , 
     n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , 
     n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , 
     n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , 
     n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , 
     n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , 
     n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , 
     n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , 
     n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , 
     n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , 
     n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , 
     n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , 
     n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , 
     n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , 
     n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , 
     n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , 
     n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , 
     n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , 
     n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , 
     n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , 
     n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , 
     n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , 
     n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , 
     n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , 
     n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , 
     n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , 
     n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , 
     n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , 
     n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , 
     n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , 
     n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , 
     n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , 
     n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , 
     n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , 
     n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , 
     n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , 
     n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , 
     n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , 
     n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , 
     n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , 
     n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , 
     n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , 
     n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , 
     n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , 
     n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , 
     n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , 
     n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , 
     n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , 
     n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , 
     n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , 
     n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , 
     n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , 
     n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , 
     n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , 
     n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , 
     n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , 
     n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , 
     n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , 
     n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , 
     n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , 
     n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , 
     n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , 
     n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , 
     n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , 
     n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , 
     n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , 
     n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , 
     n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , 
     n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , 
     n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , 
     n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , 
     n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , 
     n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , 
     n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , 
     n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , 
     n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , 
     n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , 
     n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , 
     n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , 
     n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , 
     n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , 
     n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , 
     n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , 
     n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , 
     n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , 
     n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , 
     n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , 
     n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , 
     n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , 
     n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , 
     n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , 
     n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , 
     n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , 
     n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , 
     n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , 
     n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , 
     n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , 
     n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , 
     n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , 
     n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , 
     n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , 
     n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , 
     n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , 
     n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , 
     n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , 
     n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , 
     n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , 
     n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , 
     n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , 
     n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , 
     n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , 
     n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , 
     n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , 
     n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , 
     n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , 
     n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , 
     n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , 
     n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , 
     n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , 
     n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , 
     n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , 
     n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , 
     n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , 
     n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , 
     n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , 
     n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , 
     n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , 
     n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , 
     n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , 
     n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , 
     n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , 
     n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , 
     n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , 
     n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , 
     n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , 
     n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , 
     n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , 
     n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , 
     n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , 
     n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , 
     n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , 
     n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , 
     n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , 
     n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , 
     n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , 
     n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , 
     n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , 
     n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , 
     n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , 
     n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , 
     n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , 
     n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , 
     n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , 
     n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , 
     n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , 
     n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , 
     n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , 
     n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , 
     n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , 
     n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , 
     n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , 
     n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , 
     n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , 
     n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , 
     n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , 
     n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , 
     n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , 
     n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , 
     n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , 
     n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , 
     n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , 
     n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , 
     n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , 
     n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , 
     n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , 
     n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , 
     n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , 
     n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , 
     n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , 
     n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , 
     n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , 
     n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , 
     n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , 
     n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , 
     n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , 
     n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , 
     n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , 
     n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , 
     n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , 
     n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , 
     n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , 
     n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , 
     n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , 
     n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , 
     n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , 
     n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , 
     n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , 
     n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , 
     n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , 
     n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , 
     n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , 
     n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , 
     n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , 
     n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , 
     n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , 
     n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , 
     n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , 
     n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , 
     n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , 
     n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , 
     n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , 
     n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , 
     n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , 
     n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , 
     n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , 
     n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , 
     n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , 
     n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , 
     n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , 
     n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , 
     n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , 
     n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , 
     n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , 
     n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , 
     n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , 
     n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , 
     n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , 
     n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , 
     n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , 
     n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , 
     n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , 
     n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , 
     n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , 
     n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , 
     n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , 
     n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , 
     n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , 
     n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , 
     n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , 
     n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , 
     n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , 
     n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , 
     n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , 
     n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , 
     n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , 
     n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , 
     n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , 
     n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , 
     n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , 
     n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , 
     n32694 , n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , 
     n32704 , n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , 
     n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , 
     n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , 
     n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , 
     n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , 
     n32754 , n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , 
     n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , 
     n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , 
     n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , 
     n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , 
     n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , 
     n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , 
     n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , 
     n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , 
     n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , 
     n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , 
     n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , 
     n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , 
     n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , 
     n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , 
     n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , 
     n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , 
     n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , 
     n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , 
     n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , 
     n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , 
     n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , 
     n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , 
     n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , 
     n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , 
     n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , 
     n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , 
     n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , 
     n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , 
     n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , 
     n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , 
     n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , 
     n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , 
     n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , 
     n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , 
     n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , 
     n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , 
     n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , 
     n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , 
     n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , 
     n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , 
     n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , 
     n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , 
     n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , 
     n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , 
     n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , 
     n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , 
     n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , 
     n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , 
     n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , 
     n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , 
     n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , 
     n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , 
     n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , 
     n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , 
     n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , 
     n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , 
     n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , 
     n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , 
     n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , 
     n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , 
     n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , 
     n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , 
     n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , 
     n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , 
     n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , 
     n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , 
     n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , 
     n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , 
     n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , 
     n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , 
     n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , 
     n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , 
     n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , 
     n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , 
     n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , 
     n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , 
     n33524 , n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , 
     n33534 , n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , 
     n33544 , n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , 
     n33554 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , 
     n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , 
     n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , 
     n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , 
     n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , 
     n33604 , n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , 
     n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , 
     n33624 , n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , 
     n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , 
     n33644 , n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , 
     n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , 
     n33664 , n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , 
     n33674 , n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , 
     n33684 , n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , 
     n33694 , n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , 
     n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , 
     n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , 
     n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , 
     n33734 , n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , 
     n33744 , n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , 
     n33754 , n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , 
     n33764 , n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , 
     n33774 , n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , 
     n33784 , n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , 
     n33794 , n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , 
     n33804 , n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , 
     n33814 , n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , 
     n33824 , n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , 
     n33834 , n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , 
     n33844 , n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , 
     n33854 , n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , 
     n33864 , n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , 
     n33874 , n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , 
     n33884 , n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , 
     n33894 , n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , 
     n33904 , n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , 
     n33914 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , 
     n33924 , n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , 
     n33934 , n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , 
     n33944 , n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , 
     n33954 , n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , 
     n33964 , n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , 
     n33974 , n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , 
     n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , 
     n33994 , n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , 
     n34004 , n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , 
     n34014 , n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , 
     n34024 , n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , 
     n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , 
     n34044 , n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , 
     n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , 
     n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , 
     n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , 
     n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , 
     n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , 
     n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , 
     n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , 
     n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , 
     n34134 , n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , 
     n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , 
     n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , 
     n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , 
     n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , 
     n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , 
     n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , 
     n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , 
     n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , 
     n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , 
     n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , 
     n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , 
     n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , 
     n34264 , n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , 
     n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , 
     n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , 
     n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , 
     n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , 
     n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , 
     n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , 
     n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , 
     n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , 
     n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , 
     n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , 
     n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , 
     n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , 
     n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , 
     n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , 
     n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , 
     n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , 
     n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , 
     n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , 
     n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , 
     n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , 
     n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , 
     n34484 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , 
     n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , 
     n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , 
     n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , 
     n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , 
     n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , 
     n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , 
     n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , 
     n34564 , n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , 
     n34574 , n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , 
     n34584 , n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , 
     n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , 
     n34604 , n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , 
     n34614 , n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , 
     n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , 
     n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , 
     n34644 , n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , 
     n34654 , n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , 
     n34664 , n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , 
     n34674 , n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , 
     n34684 , n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , 
     n34694 , n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , 
     n34704 , n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , 
     n34714 , n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , 
     n34724 , n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , 
     n34734 , n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , 
     n34744 , n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , 
     n34754 , n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , 
     n34764 , n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , 
     n34774 , n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , 
     n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , 
     n34794 , n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , 
     n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , 
     n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , 
     n34824 , n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , 
     n34834 , n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , 
     n34844 , n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , 
     n34854 , n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , 
     n34864 , n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , 
     n34874 , n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , 
     n34884 , n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , 
     n34894 , n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , 
     n34904 , n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , 
     n34914 , n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , 
     n34924 , n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , 
     n34934 , n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , 
     n34944 , n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , 
     n34954 , n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , 
     n34964 , n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , 
     n34974 , n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , 
     n34984 , n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , 
     n34994 , n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , 
     n35004 , n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , 
     n35014 , n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , 
     n35024 , n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , 
     n35034 , n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , 
     n35044 , n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , 
     n35054 , n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , 
     n35064 , n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , 
     n35074 , n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , 
     n35084 , n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , 
     n35094 , n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , 
     n35104 , n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , 
     n35114 , n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , 
     n35124 , n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , 
     n35134 , n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , 
     n35144 , n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , 
     n35154 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , 
     n35164 , n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , 
     n35174 , n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , 
     n35184 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , 
     n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , 
     n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , 
     n35214 , n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , 
     n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , 
     n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , 
     n35244 , n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , 
     n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , 
     n35264 , n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , 
     n35274 , n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , 
     n35284 , n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , 
     n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , 
     n35304 , n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , 
     n35314 , n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , 
     n35324 , n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , 
     n35334 , n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , 
     n35344 , n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , 
     n35354 , n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , 
     n35364 , n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , 
     n35374 , n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , 
     n35384 , n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , 
     n35394 , n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , 
     n35404 , n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , 
     n35414 , n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , 
     n35424 , n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , 
     n35434 , n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , 
     n35444 , n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , 
     n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , 
     n35464 , n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , 
     n35474 , n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , 
     n35484 , n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , 
     n35494 , n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , 
     n35504 , n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , 
     n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , 
     n35524 , n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , 
     n35534 , n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , 
     n35544 , n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , 
     n35554 , n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , 
     n35564 , n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , 
     n35574 , n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , 
     n35584 , n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , 
     n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , 
     n35604 , n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , 
     n35614 , n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , 
     n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , 
     n35634 , n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , 
     n35644 , n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , 
     n35654 , n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , 
     n35664 , n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , 
     n35674 , n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , 
     n35684 , n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , 
     n35694 , n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , 
     n35704 , n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , 
     n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , 
     n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , 
     n35734 , n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , 
     n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , 
     n35754 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , 
     n35764 , n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , 
     n35774 , n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , 
     n35784 , n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , 
     n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , 
     n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , 
     n35814 , n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , 
     n35824 , n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , 
     n35834 , n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , 
     n35844 , n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , 
     n35854 , n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , 
     n35864 , n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , 
     n35874 , n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , 
     n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , 
     n35894 , n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , 
     n35904 , n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , 
     n35914 , n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , 
     n35924 , n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , 
     n35934 , n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , 
     n35944 , n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , 
     n35954 , n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , 
     n35964 , n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , 
     n35974 , n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , 
     n35984 , n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , 
     n35994 , n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , 
     n36004 , n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , 
     n36014 , n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , 
     n36024 , n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , 
     n36034 , n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , 
     n36044 , n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , 
     n36054 , n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , 
     n36064 , n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , 
     n36074 , n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , 
     n36084 , n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , 
     n36094 , n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , 
     n36104 , n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , 
     n36114 , n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , 
     n36124 , n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , 
     n36134 , n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , 
     n36144 , n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , 
     n36154 , n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , 
     n36164 , n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , 
     n36174 , n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , 
     n36184 , n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , 
     n36194 , n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , 
     n36204 , n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , 
     n36214 , n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , 
     n36224 , n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , 
     n36234 , n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , 
     n36244 , n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , 
     n36254 , n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , 
     n36264 , n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , 
     n36274 , n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , 
     n36284 , n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , 
     n36294 , n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , 
     n36304 , n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , 
     n36314 , n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , 
     n36324 , n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , 
     n36334 , n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , 
     n36344 , n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , 
     n36354 , n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , 
     n36364 , n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , 
     n36374 , n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , 
     n36384 , n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , 
     n36394 , n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , 
     n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , 
     n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , 
     n36424 , n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , 
     n36434 , n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , 
     n36444 , n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , 
     n36454 , n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , 
     n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , 
     n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , 
     n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , 
     n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , 
     n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , 
     n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , 
     n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , 
     n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , 
     n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , 
     n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , 
     n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , 
     n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , 
     n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , 
     n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , 
     n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , 
     n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , 
     n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , 
     n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , 
     n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , 
     n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , 
     n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , 
     n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , 
     n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , 
     n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , 
     n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , 
     n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , 
     n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , 
     n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , 
     n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , 
     n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , 
     n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , 
     n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , 
     n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , 
     n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , 
     n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , 
     n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , 
     n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , 
     n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , 
     n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , 
     n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , 
     n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , 
     n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , 
     n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , 
     n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , 
     n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , 
     n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , 
     n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , 
     n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , 
     n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , 
     n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , 
     n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , 
     n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , 
     n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , 
     n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , 
     n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , 
     n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , 
     n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , 
     n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , 
     n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , 
     n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , 
     n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , 
     n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , 
     n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , 
     n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , 
     n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , 
     n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , 
     n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , 
     n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , 
     n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , 
     n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , 
     n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , 
     n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , 
     n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , 
     n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , 
     n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , 
     n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , 
     n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , 
     n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , 
     n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , 
     n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , 
     n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , 
     n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , 
     n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , 
     n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , 
     n37304 , n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , 
     n37314 , n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , 
     n37324 , n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , 
     n37334 , n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , 
     n37344 , n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , 
     n37354 , n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , 
     n37364 , n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , n37373 , 
     n37374 , n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , n37383 , 
     n37384 , n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , n37393 , 
     n37394 , n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , n37403 , 
     n37404 , n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , 
     n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , 
     n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , n37433 , 
     n37434 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , 
     n37444 , n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , 
     n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , 
     n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , 
     n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , 
     n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , 
     n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , 
     n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , 
     n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , 
     n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , 
     n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , 
     n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , 
     n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , 
     n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , 
     n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , 
     n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , 
     n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , 
     n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , 
     n37614 , n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , n37623 , 
     n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , 
     n37634 , n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , 
     n37644 , n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , 
     n37654 , n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , n37663 , 
     n37664 , n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , 
     n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , 
     n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , 
     n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , 
     n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , 
     n37714 , n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , 
     n37724 , n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , n37733 , 
     n37734 , n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , n37743 , 
     n37744 , n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , n37753 , 
     n37754 , n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , 
     n37764 , n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , n37773 , 
     n37774 , n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , n37783 , 
     n37784 , n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , n37793 , 
     n37794 , n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , n37803 , 
     n37804 , n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , n37813 , 
     n37814 , n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , n37823 , 
     n37824 , n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , n37833 , 
     n37834 , n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , n37843 , 
     n37844 , n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , n37853 , 
     n37854 , n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , n37863 , 
     n37864 , n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , n37873 , 
     n37874 , n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , n37883 , 
     n37884 , n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , n37893 , 
     n37894 , n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , 
     n37904 , n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , 
     n37914 , n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , 
     n37924 , n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , n37933 , 
     n37934 , n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , n37943 , 
     n37944 , n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , n37953 , 
     n37954 , n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , n37963 , 
     n37964 , n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , n37973 , 
     n37974 , n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , n37983 , 
     n37984 , n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , n37993 , 
     n37994 , n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , n38003 , 
     n38004 , n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , n38013 , 
     n38014 , n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , n38023 , 
     n38024 , n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , n38033 , 
     n38034 , n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , n38043 , 
     n38044 , n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , n38053 , 
     n38054 , n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , n38063 , 
     n38064 , n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , n38073 , 
     n38074 , n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , n38083 , 
     n38084 , n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , n38093 , 
     n38094 , n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , n38103 , 
     n38104 , n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , n38113 , 
     n38114 , n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , n38123 , 
     n38124 , n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , n38133 , 
     n38134 , n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , n38143 , 
     n38144 , n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , n38153 , 
     n38154 , n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , n38163 , 
     n38164 , n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , n38173 , 
     n38174 , n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , n38183 , 
     n38184 , n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , n38193 , 
     n38194 , n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , n38203 , 
     n38204 , n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , n38213 , 
     n38214 , n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , n38223 , 
     n38224 , n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , n38233 , 
     n38234 , n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , 
     n38244 , n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , n38253 , 
     n38254 , n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , n38263 , 
     n38264 , n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , n38273 , 
     n38274 , n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , n38283 , 
     n38284 , n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , n38291 , n38292 , n38293 , 
     n38294 , n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , n38303 , 
     n38304 , n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , n38313 , 
     n38314 , n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , n38323 , 
     n38324 , n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , n38333 , 
     n38334 , n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , n38343 , 
     n38344 , n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , n38353 , 
     n38354 , n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , n38363 , 
     n38364 , n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , n38371 , n38372 , n38373 , 
     n38374 , n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , n38381 , n38382 , n38383 , 
     n38384 , n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , n38393 , 
     n38394 , n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , n38403 , 
     n38404 , n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , n38413 , 
     n38414 , n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , n38423 , 
     n38424 , n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , n38433 , 
     n38434 , n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , n38443 , 
     n38444 , n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , n38451 , n38452 , n38453 , 
     n38454 , n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , n38463 , 
     n38464 , n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , n38473 , 
     n38474 , n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , n38483 , 
     n38484 , n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , n38493 , 
     n38494 , n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , n38501 , n38502 , n38503 , 
     n38504 , n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , n38513 , 
     n38514 , n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , n38523 , 
     n38524 , n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , n38533 , 
     n38534 , n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , n38543 , 
     n38544 , n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , n38553 , 
     n38554 , n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , n38563 , 
     n38564 , n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , n38573 , 
     n38574 , n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , n38583 , 
     n38584 , n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , n38591 , n38592 , n38593 , 
     n38594 , n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , n38601 , n38602 , n38603 , 
     n38604 , n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , n38611 , n38612 , n38613 , 
     n38614 , n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , n38621 , n38622 , n38623 , 
     n38624 , n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , n38631 , n38632 , n38633 , 
     n38634 , n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , n38641 , n38642 , n38643 , 
     n38644 , n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , n38651 , n38652 , n38653 , 
     n38654 , n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , n38661 , n38662 , n38663 , 
     n38664 , n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , n38671 , n38672 , n38673 , 
     n38674 , n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , n38681 , n38682 , n38683 , 
     n38684 , n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , n38691 , n38692 , n38693 , 
     n38694 , n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , n38701 , n38702 , n38703 , 
     n38704 , n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , n38711 , n38712 , n38713 , 
     n38714 , n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , n38721 , n38722 , n38723 , 
     n38724 , n38725 , n38726 , n38727 , n38728 , n38729 , n38730 , n38731 , n38732 , n38733 , 
     n38734 , n38735 , n38736 , n38737 , n38738 , n38739 , n38740 , n38741 , n38742 , n38743 , 
     n38744 , n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , n38751 , n38752 , n38753 , 
     n38754 , n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , n38761 , n38762 , n38763 , 
     n38764 , n38765 , n38766 , n38767 , n38768 , n38769 , n38770 , n38771 , n38772 , n38773 , 
     n38774 , n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , n38781 , n38782 , n38783 , 
     n38784 , n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , n38791 , n38792 , n38793 , 
     n38794 , n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , n38801 , n38802 , n38803 , 
     n38804 , n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , n38811 , n38812 , n38813 , 
     n38814 , n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , n38821 , n38822 , n38823 , 
     n38824 , n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , n38831 , n38832 , n38833 , 
     n38834 , n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , n38841 , n38842 , n38843 , 
     n38844 , n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , n38851 , n38852 , n38853 , 
     n38854 , n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , n38861 , n38862 , n38863 , 
     n38864 , n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , n38871 , n38872 , n38873 , 
     n38874 , n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , n38881 , n38882 , n38883 , 
     n38884 , n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , n38891 , n38892 , n38893 , 
     n38894 , n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , n38903 , 
     n38904 , n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , n38911 , n38912 , n38913 , 
     n38914 , n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , n38921 , n38922 , n38923 , 
     n38924 , n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , n38931 , n38932 , n38933 , 
     n38934 , n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , n38941 , n38942 , n38943 , 
     n38944 , n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , n38951 , n38952 , n38953 , 
     n38954 , n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , n38961 , n38962 , n38963 , 
     n38964 , n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , n38971 , n38972 , n38973 , 
     n38974 , n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , n38981 , n38982 , n38983 , 
     n38984 , n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , n38991 , n38992 , n38993 , 
     n38994 , n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , n39001 , n39002 , n39003 , 
     n39004 , n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , n39011 , n39012 , n39013 , 
     n39014 , n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , n39021 , n39022 , n39023 , 
     n39024 , n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , n39031 , n39032 , n39033 , 
     n39034 , n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , n39041 , n39042 , n39043 , 
     n39044 , n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , n39051 , n39052 , n39053 , 
     n39054 , n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , n39061 , n39062 , n39063 , 
     n39064 , n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , n39071 , n39072 , n39073 , 
     n39074 , n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , n39081 , n39082 , n39083 , 
     n39084 , n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , n39091 , n39092 , n39093 , 
     n39094 , n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , n39101 , n39102 , n39103 , 
     n39104 , n39105 , n39106 , n39107 , n39108 , n39109 , n39110 , n39111 , n39112 , n39113 , 
     n39114 , n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , n39121 , n39122 , n39123 , 
     n39124 , n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , n39131 , n39132 , n39133 , 
     n39134 , n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , n39141 , n39142 , n39143 , 
     n39144 , n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , n39153 , 
     n39154 , n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , n39161 , n39162 , n39163 , 
     n39164 , n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , n39171 , n39172 , n39173 , 
     n39174 , n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , n39181 , n39182 , n39183 , 
     n39184 , n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , n39191 , n39192 , n39193 , 
     n39194 , n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , n39201 , n39202 , n39203 , 
     n39204 , n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , n39211 , n39212 , n39213 , 
     n39214 , n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , n39221 , n39222 , n39223 , 
     n39224 , n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , n39233 , 
     n39234 , n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , n39241 , n39242 , n39243 , 
     n39244 , n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , n39251 , n39252 , n39253 , 
     n39254 , n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , n39261 , n39262 , n39263 , 
     n39264 , n39265 , n39266 , n39267 , n39268 , n39269 , n39270 , n39271 , n39272 , n39273 , 
     n39274 , n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , n39281 , n39282 , n39283 , 
     n39284 , n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , n39291 , n39292 , n39293 , 
     n39294 , n39295 , n39296 , n39297 , n39298 , n39299 , n39300 , n39301 , n39302 , n39303 , 
     n39304 , n39305 , n39306 , n39307 , n39308 , n39309 , n39310 , n39311 , n39312 , n39313 , 
     n39314 , n39315 , n39316 , n39317 , n39318 , n39319 , n39320 , n39321 , n39322 , n39323 , 
     n39324 , n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , n39331 , n39332 , n39333 , 
     n39334 , n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , n39341 , n39342 , n39343 , 
     n39344 , n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , n39351 , n39352 , n39353 , 
     n39354 , n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , n39361 , n39362 , n39363 , 
     n39364 , n39365 , n39366 , n39367 , n39368 , n39369 , n39370 , n39371 , n39372 , n39373 , 
     n39374 , n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , n39381 , n39382 , n39383 , 
     n39384 , n39385 , n39386 , n39387 , n39388 , n39389 , n39390 , n39391 , n39392 , n39393 , 
     n39394 , n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , n39401 , n39402 , n39403 , 
     n39404 , n39405 , n39406 , n39407 , n39408 , n39409 , n39410 , n39411 , n39412 , n39413 , 
     n39414 , n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , n39421 , n39422 , n39423 , 
     n39424 , n39425 , n39426 , n39427 , n39428 , n39429 , n39430 , n39431 , n39432 , n39433 , 
     n39434 , n39435 , n39436 , n39437 , n39438 , n39439 , n39440 , n39441 , n39442 , n39443 , 
     n39444 , n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , n39451 , n39452 , n39453 , 
     n39454 , n39455 , n39456 , n39457 , n39458 , n39459 , n39460 , n39461 , n39462 , n39463 , 
     n39464 , n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , n39471 , n39472 , n39473 , 
     n39474 , n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , n39481 , n39482 , n39483 , 
     n39484 , n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , n39491 , n39492 , n39493 , 
     n39494 , n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , n39501 , n39502 , n39503 , 
     n39504 , n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , n39511 , n39512 , n39513 , 
     n39514 , n39515 , n39516 , n39517 , n39518 , n39519 , n39520 , n39521 , n39522 , n39523 , 
     n39524 , n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , n39531 , n39532 , n39533 , 
     n39534 , n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , n39541 , n39542 , n39543 , 
     n39544 , n39545 , n39546 , n39547 , n39548 , n39549 , n39550 , n39551 , n39552 , n39553 , 
     n39554 , n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , n39561 , n39562 , n39563 , 
     n39564 , n39565 , n39566 , n39567 , n39568 , n39569 , n39570 , n39571 , n39572 , n39573 , 
     n39574 , n39575 , n39576 , n39577 , n39578 , n39579 , n39580 , n39581 , n39582 , n39583 , 
     n39584 , n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , n39591 , n39592 , n39593 , 
     n39594 , n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , n39601 , n39602 , n39603 , 
     n39604 , n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , n39611 , n39612 , n39613 , 
     n39614 , n39615 , n39616 , n39617 , n39618 , n39619 , n39620 , n39621 , n39622 , n39623 , 
     n39624 , n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , n39631 , n39632 , n39633 , 
     n39634 , n39635 , n39636 , n39637 , n39638 , n39639 , n39640 , n39641 , n39642 , n39643 , 
     n39644 , n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , n39651 , n39652 , n39653 , 
     n39654 , n39655 , n39656 , n39657 , n39658 , n39659 , n39660 , n39661 , n39662 , n39663 , 
     n39664 , n39665 , n39666 , n39667 , n39668 , n39669 , n39670 , n39671 , n39672 , n39673 , 
     n39674 , n39675 , n39676 , n39677 , n39678 , n39679 , n39680 , n39681 , n39682 , n39683 , 
     n39684 , n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , n39691 , n39692 , n39693 , 
     n39694 , n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , n39701 , n39702 , n39703 , 
     n39704 , n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , n39711 , n39712 , n39713 , 
     n39714 , n39715 , n39716 , n39717 , n39718 , n39719 , n39720 , n39721 , n39722 , n39723 , 
     n39724 , n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , n39731 , n39732 , n39733 , 
     n39734 , n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , n39741 , n39742 , n39743 , 
     n39744 , n39745 , n39746 , n39747 , n39748 , n39749 , n39750 , n39751 , n39752 , n39753 , 
     n39754 , n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , n39761 , n39762 , n39763 , 
     n39764 , n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , n39771 , n39772 , n39773 , 
     n39774 , n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , n39781 , n39782 , n39783 , 
     n39784 , n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , n39791 , n39792 , n39793 , 
     n39794 , n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , n39801 , n39802 , n39803 , 
     n39804 , n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , n39811 , n39812 , n39813 , 
     n39814 , n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , n39821 , n39822 , n39823 , 
     n39824 , n39825 , n39826 , n39827 , n39828 , n39829 , n39830 , n39831 , n39832 , n39833 , 
     n39834 , n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , n39841 , n39842 , n39843 , 
     n39844 , n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , n39851 , n39852 , n39853 , 
     n39854 , n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , n39861 , n39862 , n39863 , 
     n39864 , n39865 , n39866 , n39867 , n39868 , n39869 , n39870 , n39871 , n39872 , n39873 , 
     n39874 , n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , n39881 , n39882 , n39883 , 
     n39884 , n39885 , n39886 , n39887 , n39888 , n39889 , n39890 , n39891 , n39892 , n39893 , 
     n39894 , n39895 , n39896 , n39897 , n39898 , n39899 , n39900 , n39901 , n39902 , n39903 , 
     n39904 , n39905 , n39906 , n39907 , n39908 , n39909 , n39910 , n39911 , n39912 , n39913 , 
     n39914 , n39915 , n39916 , n39917 , n39918 , n39919 , n39920 , n39921 , n39922 , n39923 , 
     n39924 , n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , n39931 , n39932 , n39933 , 
     n39934 , n39935 , n39936 , n39937 , n39938 , n39939 , n39940 , n39941 , n39942 , n39943 , 
     n39944 , n39945 , n39946 , n39947 , n39948 , n39949 , n39950 , n39951 , n39952 , n39953 , 
     n39954 , n39955 , n39956 , n39957 , n39958 , n39959 , n39960 , n39961 , n39962 , n39963 , 
     n39964 , n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , n39971 , n39972 , n39973 , 
     n39974 , n39975 , n39976 , n39977 , n39978 , n39979 , n39980 , n39981 , n39982 , n39983 , 
     n39984 , n39985 , n39986 , n39987 , n39988 , n39989 , n39990 , n39991 , n39992 , n39993 , 
     n39994 , n39995 , n39996 , n39997 , n39998 , n39999 , n40000 , n40001 , n40002 , n40003 , 
     n40004 , n40005 , n40006 , n40007 , n40008 , n40009 , n40010 , n40011 , n40012 , n40013 , 
     n40014 , n40015 , n40016 , n40017 , n40018 , n40019 , n40020 , n40021 , n40022 , n40023 , 
     n40024 , n40025 , n40026 , n40027 , n40028 , n40029 , n40030 , n40031 , n40032 , n40033 , 
     n40034 , n40035 , n40036 , n40037 , n40038 , n40039 , n40040 , n40041 , n40042 , n40043 , 
     n40044 , n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , n40051 , n40052 , n40053 , 
     n40054 , n40055 , n40056 , n40057 , n40058 , n40059 , n40060 , n40061 , n40062 , n40063 , 
     n40064 , n40065 , n40066 , n40067 , n40068 , n40069 , n40070 , n40071 , n40072 , n40073 , 
     n40074 , n40075 , n40076 , n40077 , n40078 , n40079 , n40080 , n40081 , n40082 , n40083 , 
     n40084 , n40085 , n40086 , n40087 , n40088 , n40089 , n40090 , n40091 , n40092 , n40093 , 
     n40094 , n40095 , n40096 , n40097 , n40098 , n40099 , n40100 , n40101 , n40102 , n40103 , 
     n40104 , n40105 , n40106 , n40107 , n40108 , n40109 , n40110 , n40111 , n40112 , n40113 , 
     n40114 , n40115 , n40116 , n40117 , n40118 , n40119 , n40120 , n40121 , n40122 , n40123 , 
     n40124 , n40125 , n40126 , n40127 , n40128 , n40129 , n40130 , n40131 , n40132 , n40133 , 
     n40134 , n40135 , n40136 , n40137 , n40138 , n40139 , n40140 , n40141 , n40142 , n40143 , 
     n40144 , n40145 , n40146 , n40147 , n40148 , n40149 , n40150 , n40151 , n40152 , n40153 , 
     n40154 , n40155 , n40156 , n40157 , n40158 , n40159 , n40160 , n40161 , n40162 , n40163 , 
     n40164 , n40165 , n40166 , n40167 , n40168 , n40169 , n40170 , n40171 , n40172 , n40173 , 
     n40174 , n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , n40181 , n40182 , n40183 , 
     n40184 , n40185 , n40186 , n40187 , n40188 , n40189 , n40190 , n40191 , n40192 , n40193 , 
     n40194 , n40195 , n40196 , n40197 , n40198 , n40199 , n40200 , n40201 , n40202 , n40203 , 
     n40204 , n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , n40211 , n40212 , n40213 , 
     n40214 , n40215 , n40216 , n40217 , n40218 , n40219 , n40220 , n40221 , n40222 , n40223 , 
     n40224 , n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , n40231 , n40232 , n40233 , 
     n40234 , n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , n40241 , n40242 , n40243 , 
     n40244 , n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , n40251 , n40252 , n40253 , 
     n40254 , n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , n40261 , n40262 , n40263 , 
     n40264 , n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , n40271 , n40272 , n40273 , 
     n40274 , n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , n40281 , n40282 , n40283 , 
     n40284 , n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , n40291 , n40292 , n40293 , 
     n40294 , n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , n40301 , n40302 , n40303 , 
     n40304 , n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , n40311 , n40312 , n40313 , 
     n40314 , n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , n40321 , n40322 , n40323 , 
     n40324 , n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , n40331 , n40332 , n40333 , 
     n40334 , n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , n40341 , n40342 , n40343 , 
     n40344 , n40345 , n40346 , n40347 , n40348 , n40349 , n40350 , n40351 , n40352 , n40353 , 
     n40354 , n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , n40361 , n40362 , n40363 , 
     n40364 , n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , n40371 , n40372 , n40373 , 
     n40374 , n40375 , n40376 , n40377 , n40378 , n40379 , n40380 , n40381 , n40382 , n40383 , 
     n40384 , n40385 , n40386 , n40387 , n40388 , n40389 , n40390 , n40391 , n40392 , n40393 , 
     n40394 , n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , n40401 , n40402 , n40403 , 
     n40404 , n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , n40411 , n40412 , n40413 , 
     n40414 , n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , n40421 , n40422 , n40423 , 
     n40424 , n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , n40431 , n40432 , n40433 , 
     n40434 , n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , n40441 , n40442 , n40443 , 
     n40444 , n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , n40451 , n40452 , n40453 , 
     n40454 , n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , n40461 , n40462 , n40463 , 
     n40464 , n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , n40471 , n40472 , n40473 , 
     n40474 , n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , n40481 , n40482 , n40483 , 
     n40484 , n40485 , n40486 , n40487 , n40488 , n40489 , n40490 , n40491 , n40492 , n40493 , 
     n40494 , n40495 , n40496 , n40497 , n40498 , n40499 , n40500 , n40501 , n40502 , n40503 , 
     n40504 , n40505 , n40506 , n40507 , n40508 , n40509 , n40510 , n40511 , n40512 , n40513 , 
     n40514 , n40515 , n40516 , n40517 , n40518 , n40519 , n40520 , n40521 , n40522 , n40523 , 
     n40524 , n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , n40531 , n40532 , n40533 , 
     n40534 , n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , n40541 , n40542 , n40543 , 
     n40544 , n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , n40551 , n40552 , n40553 , 
     n40554 , n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , n40561 , n40562 , n40563 , 
     n40564 , n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , n40571 , n40572 , n40573 , 
     n40574 , n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , n40581 , n40582 , n40583 , 
     n40584 , n40585 , n40586 , n40587 , n40588 , n40589 , n40590 , n40591 , n40592 , n40593 , 
     n40594 , n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , n40601 , n40602 , n40603 , 
     n40604 , n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , n40611 , n40612 , n40613 , 
     n40614 , n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , n40621 , n40622 , n40623 , 
     n40624 , n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , n40631 , n40632 , n40633 , 
     n40634 , n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , n40641 , n40642 , n40643 , 
     n40644 , n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , n40651 , n40652 , n40653 , 
     n40654 , n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , n40661 , n40662 , n40663 , 
     n40664 , n40665 , n40666 , n40667 , n40668 , n40669 , n40670 , n40671 , n40672 , n40673 , 
     n40674 , n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , n40681 , n40682 , n40683 , 
     n40684 , n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , n40691 , n40692 , n40693 , 
     n40694 , n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , n40701 , n40702 , n40703 , 
     n40704 , n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , n40711 , n40712 , n40713 , 
     n40714 , n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , n40721 , n40722 , n40723 , 
     n40724 , n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , n40731 , n40732 , n40733 , 
     n40734 , n40735 , n40736 , n40737 , n40738 , n40739 , n40740 , n40741 , n40742 , n40743 , 
     n40744 , n40745 , n40746 , n40747 , n40748 , n40749 , n40750 , n40751 , n40752 , n40753 , 
     n40754 , n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , n40761 , n40762 , n40763 , 
     n40764 , n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , n40771 , n40772 , n40773 , 
     n40774 , n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , n40781 , n40782 , n40783 , 
     n40784 , n40785 , n40786 , n40787 , n40788 , n40789 , n40790 , n40791 , n40792 , n40793 , 
     n40794 , n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , n40801 , n40802 , n40803 , 
     n40804 , n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , n40811 , n40812 , n40813 , 
     n40814 , n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , n40821 , n40822 , n40823 , 
     n40824 , n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , n40831 , n40832 , n40833 , 
     n40834 , n40835 , n40836 , n40837 , n40838 , n40839 , n40840 , n40841 , n40842 , n40843 , 
     n40844 , n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , n40851 , n40852 , n40853 , 
     n40854 , n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , n40861 , n40862 , n40863 , 
     n40864 , n40865 , n40866 , n40867 , n40868 , n40869 , n40870 , n40871 , n40872 , n40873 , 
     n40874 , n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , n40881 , n40882 , n40883 , 
     n40884 , n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , n40891 , n40892 , n40893 , 
     n40894 , n40895 , n40896 , n40897 , n40898 , n40899 , n40900 , n40901 , n40902 , n40903 , 
     n40904 , n40905 , n40906 , n40907 , n40908 , n40909 , n40910 , n40911 , n40912 , n40913 , 
     n40914 , n40915 , n40916 , n40917 , n40918 , n40919 , n40920 , n40921 , n40922 , n40923 , 
     n40924 , n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , n40931 , n40932 , n40933 , 
     n40934 , n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , n40941 , n40942 , n40943 , 
     n40944 , n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , n40951 , n40952 , n40953 , 
     n40954 , n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , n40961 , n40962 , n40963 , 
     n40964 , n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , n40971 , n40972 , n40973 , 
     n40974 , n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , n40981 , n40982 , n40983 , 
     n40984 , n40985 , n40986 , n40987 , n40988 , n40989 , n40990 , n40991 , n40992 , n40993 , 
     n40994 , n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , n41001 , n41002 , n41003 , 
     n41004 , n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , n41011 , n41012 , n41013 , 
     n41014 , n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , n41021 , n41022 , n41023 , 
     n41024 , n41025 , n41026 , n41027 , n41028 , n41029 , n41030 , n41031 , n41032 , n41033 , 
     n41034 , n41035 , n41036 , n41037 , n41038 , n41039 , n41040 , n41041 , n41042 , n41043 , 
     n41044 , n41045 , n41046 , n41047 , n41048 , n41049 , n41050 , n41051 , n41052 , n41053 , 
     n41054 , n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , n41061 , n41062 , n41063 , 
     n41064 , n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , n41071 , n41072 , n41073 , 
     n41074 , n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , n41081 , n41082 , n41083 , 
     n41084 , n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , n41091 , n41092 , n41093 , 
     n41094 , n41095 , n41096 , n41097 , n41098 , n41099 , n41100 , n41101 , n41102 , n41103 , 
     n41104 , n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , n41111 , n41112 , n41113 , 
     n41114 , n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , n41121 , n41122 , n41123 , 
     n41124 , n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , n41131 , n41132 , n41133 , 
     n41134 , n41135 , n41136 , n41137 , n41138 , n41139 , n41140 , n41141 , n41142 , n41143 , 
     n41144 , n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , n41151 , n41152 , n41153 , 
     n41154 , n41155 , n41156 , n41157 , n41158 , n41159 , n41160 , n41161 , n41162 , n41163 , 
     n41164 , n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , n41171 , n41172 , n41173 , 
     n41174 , n41175 , n41176 , n41177 , n41178 , n41179 , n41180 , n41181 , n41182 , n41183 , 
     n41184 , n41185 , n41186 , n41187 , n41188 , n41189 , n41190 , n41191 , n41192 , n41193 , 
     n41194 , n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , n41201 , n41202 , n41203 , 
     n41204 , n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , n41211 , n41212 , n41213 , 
     n41214 , n41215 , n41216 , n41217 , n41218 , n41219 , n41220 , n41221 , n41222 , n41223 , 
     n41224 , n41225 , n41226 , n41227 , n41228 , n41229 , n41230 , n41231 , n41232 , n41233 , 
     n41234 , n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , n41241 , n41242 , n41243 , 
     n41244 , n41245 , n41246 , n41247 , n41248 , n41249 , n41250 , n41251 , n41252 , n41253 , 
     n41254 , n41255 , n41256 , n41257 , n41258 , n41259 , n41260 , n41261 , n41262 , n41263 , 
     n41264 , n41265 , n41266 , n41267 , n41268 , n41269 , n41270 , n41271 , n41272 , n41273 , 
     n41274 , n41275 , n41276 , n41277 , n41278 , n41279 , n41280 , n41281 , n41282 , n41283 , 
     n41284 , n41285 , n41286 , n41287 , n41288 , n41289 , n41290 , n41291 , n41292 , n41293 , 
     n41294 , n41295 , n41296 , n41297 , n41298 , n41299 , n41300 , n41301 , n41302 , n41303 , 
     n41304 , n41305 , n41306 , n41307 , n41308 , n41309 , n41310 , n41311 , n41312 , n41313 , 
     n41314 , n41315 , n41316 , n41317 , n41318 , n41319 , n41320 , n41321 , n41322 , n41323 , 
     n41324 , n41325 , n41326 , n41327 , n41328 , n41329 , n41330 , n41331 , n41332 , n41333 , 
     n41334 , n41335 , n41336 , n41337 , n41338 , n41339 , n41340 , n41341 , n41342 , n41343 , 
     n41344 , n41345 , n41346 , n41347 , n41348 , n41349 , n41350 , n41351 , n41352 , n41353 , 
     n41354 , n41355 , n41356 , n41357 , n41358 , n41359 , n41360 , n41361 , n41362 , n41363 , 
     n41364 , n41365 , n41366 , n41367 , n41368 , n41369 , n41370 , n41371 , n41372 , n41373 , 
     n41374 , n41375 , n41376 , n41377 , n41378 , n41379 , n41380 , n41381 , n41382 , n41383 , 
     n41384 , n41385 , n41386 , n41387 , n41388 , n41389 , n41390 , n41391 , n41392 , n41393 , 
     n41394 , n41395 , n41396 , n41397 , n41398 , n41399 , n41400 , n41401 , n41402 , n41403 , 
     n41404 , n41405 , n41406 , n41407 , n41408 , n41409 , n41410 , n41411 , n41412 , n41413 , 
     n41414 , n41415 , n41416 , n41417 , n41418 , n41419 , n41420 , n41421 , n41422 , n41423 , 
     n41424 , n41425 , n41426 , n41427 , n41428 , n41429 , n41430 , n41431 , n41432 , n41433 , 
     n41434 , n41435 , n41436 , n41437 , n41438 , n41439 , n41440 , n41441 , n41442 , n41443 , 
     n41444 , n41445 , n41446 , n41447 , n41448 , n41449 , n41450 , n41451 , n41452 , n41453 , 
     n41454 , n41455 , n41456 , n41457 , n41458 , n41459 , n41460 , n41461 , n41462 , n41463 , 
     n41464 , n41465 , n41466 , n41467 , n41468 , n41469 , n41470 , n41471 , n41472 , n41473 , 
     n41474 , n41475 , n41476 , n41477 , n41478 , n41479 , n41480 , n41481 , n41482 , n41483 , 
     n41484 , n41485 , n41486 , n41487 , n41488 , n41489 , n41490 , n41491 , n41492 , n41493 , 
     n41494 , n41495 , n41496 , n41497 , n41498 , n41499 , n41500 , n41501 , n41502 , n41503 , 
     n41504 , n41505 , n41506 , n41507 , n41508 , n41509 , n41510 , n41511 , n41512 , n41513 , 
     n41514 , n41515 , n41516 , n41517 , n41518 , n41519 , n41520 , n41521 , n41522 , n41523 , 
     n41524 , n41525 , n41526 , n41527 , n41528 , n41529 , n41530 , n41531 , n41532 , n41533 , 
     n41534 , n41535 , n41536 , n41537 , n41538 , n41539 , n41540 , n41541 , n41542 , n41543 , 
     n41544 , n41545 , n41546 , n41547 , n41548 , n41549 , n41550 , n41551 , n41552 , n41553 , 
     n41554 , n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , n41561 , n41562 , n41563 , 
     n41564 , n41565 , n41566 , n41567 , n41568 , n41569 , n41570 , n41571 , n41572 , n41573 , 
     n41574 , n41575 , n41576 , n41577 , n41578 , n41579 , n41580 , n41581 , n41582 , n41583 , 
     n41584 , n41585 , n41586 , n41587 , n41588 , n41589 , n41590 , n41591 , n41592 , n41593 , 
     n41594 , n41595 , n41596 , n41597 , n41598 , n41599 , n41600 , n41601 , n41602 , n41603 , 
     n41604 , n41605 , n41606 , n41607 , n41608 , n41609 , n41610 , n41611 , n41612 , n41613 , 
     n41614 , n41615 , n41616 , n41617 , n41618 , n41619 , n41620 , n41621 , n41622 , n41623 , 
     n41624 , n41625 , n41626 , n41627 , n41628 , n41629 , n41630 , n41631 , n41632 , n41633 , 
     n41634 , n41635 , n41636 , n41637 , n41638 , n41639 , n41640 , n41641 , n41642 , n41643 , 
     n41644 , n41645 , n41646 , n41647 , n41648 , n41649 , n41650 , n41651 , n41652 , n41653 , 
     n41654 , n41655 , n41656 , n41657 , n41658 , n41659 , n41660 , n41661 , n41662 , n41663 , 
     n41664 , n41665 , n41666 , n41667 , n41668 , n41669 , n41670 , n41671 , n41672 , n41673 , 
     n41674 , n41675 , n41676 , n41677 , n41678 , n41679 , n41680 , n41681 , n41682 , n41683 , 
     n41684 , n41685 , n41686 , n41687 , n41688 , n41689 , n41690 , n41691 , n41692 , n41693 , 
     n41694 , n41695 , n41696 , n41697 , n41698 , n41699 , n41700 , n41701 , n41702 , n41703 , 
     n41704 , n41705 , n41706 , n41707 , n41708 , n41709 , n41710 , n41711 , n41712 , n41713 , 
     n41714 , n41715 , n41716 , n41717 , n41718 , n41719 , n41720 , n41721 , n41722 , n41723 , 
     n41724 , n41725 , n41726 , n41727 , n41728 , n41729 , n41730 , n41731 , n41732 , n41733 , 
     n41734 , n41735 , n41736 , n41737 , n41738 , n41739 , n41740 , n41741 , n41742 , n41743 , 
     n41744 , n41745 , n41746 , n41747 , n41748 , n41749 , n41750 , n41751 , n41752 , n41753 , 
     n41754 , n41755 , n41756 , n41757 , n41758 , n41759 , n41760 , n41761 , n41762 , n41763 , 
     n41764 , n41765 , n41766 , n41767 , n41768 , n41769 , n41770 , n41771 , n41772 , n41773 , 
     n41774 , n41775 , n41776 , n41777 , n41778 , n41779 , n41780 , n41781 , n41782 , n41783 , 
     n41784 , n41785 , n41786 , n41787 , n41788 , n41789 , n41790 , n41791 , n41792 , n41793 , 
     n41794 , n41795 , n41796 , n41797 , n41798 , n41799 , n41800 , n41801 , n41802 , n41803 , 
     n41804 , n41805 , n41806 , n41807 , n41808 , n41809 , n41810 , n41811 , n41812 , n41813 , 
     n41814 , n41815 , n41816 , n41817 , n41818 , n41819 , n41820 , n41821 , n41822 , n41823 , 
     n41824 , n41825 , n41826 , n41827 , n41828 , n41829 , n41830 , n41831 , n41832 , n41833 , 
     n41834 , n41835 , n41836 , n41837 , n41838 , n41839 , n41840 , n41841 , n41842 , n41843 , 
     n41844 , n41845 , n41846 , n41847 , n41848 , n41849 , n41850 , n41851 , n41852 , n41853 , 
     n41854 , n41855 , n41856 , n41857 , n41858 , n41859 , n41860 , n41861 , n41862 , n41863 , 
     n41864 , n41865 , n41866 , n41867 , n41868 , n41869 , n41870 , n41871 , n41872 , n41873 , 
     n41874 , n41875 , n41876 , n41877 , n41878 , n41879 , n41880 , n41881 , n41882 , n41883 , 
     n41884 , n41885 , n41886 , n41887 , n41888 , n41889 , n41890 , n41891 , n41892 , n41893 , 
     n41894 , n41895 , n41896 , n41897 , n41898 , n41899 , n41900 , n41901 , n41902 , n41903 , 
     n41904 , n41905 , n41906 , n41907 , n41908 , n41909 , n41910 , n41911 , n41912 , n41913 , 
     n41914 , n41915 , n41916 , n41917 , n41918 , n41919 , n41920 , n41921 , n41922 , n41923 , 
     n41924 , n41925 , n41926 , n41927 , n41928 , n41929 , n41930 , n41931 , n41932 , n41933 , 
     n41934 , n41935 , n41936 , n41937 , n41938 , n41939 , n41940 , n41941 , n41942 , n41943 , 
     n41944 , n41945 , n41946 , n41947 , n41948 , n41949 , n41950 , n41951 , n41952 , n41953 , 
     n41954 , n41955 , n41956 , n41957 , n41958 , n41959 , n41960 , n41961 , n41962 , n41963 , 
     n41964 , n41965 , n41966 , n41967 , n41968 , n41969 , n41970 , n41971 , n41972 , n41973 , 
     n41974 , n41975 , n41976 , n41977 , n41978 , n41979 , n41980 , n41981 , n41982 , n41983 , 
     n41984 , n41985 , n41986 , n41987 , n41988 , n41989 , n41990 , n41991 , n41992 , n41993 , 
     n41994 , n41995 , n41996 , n41997 , n41998 , n41999 , n42000 , n42001 , n42002 , n42003 , 
     n42004 , n42005 , n42006 , n42007 , n42008 , n42009 , n42010 , n42011 , n42012 , n42013 , 
     n42014 , n42015 , n42016 , n42017 , n42018 , n42019 , n42020 , n42021 , n42022 , n42023 , 
     n42024 , n42025 , n42026 , n42027 , n42028 , n42029 , n42030 , n42031 , n42032 , n42033 , 
     n42034 , n42035 , n42036 , n42037 , n42038 , n42039 , n42040 , n42041 , n42042 , n42043 , 
     n42044 , n42045 , n42046 , n42047 , n42048 , n42049 , n42050 , n42051 , n42052 , n42053 , 
     n42054 , n42055 , n42056 , n42057 , n42058 , n42059 , n42060 , n42061 , n42062 , n42063 , 
     n42064 , n42065 , n42066 , n42067 , n42068 , n42069 , n42070 , n42071 , n42072 , n42073 , 
     n42074 , n42075 , n42076 , n42077 , n42078 , n42079 , n42080 , n42081 , n42082 , n42083 , 
     n42084 , n42085 , n42086 , n42087 , n42088 , n42089 , n42090 , n42091 , n42092 , n42093 , 
     n42094 , n42095 , n42096 , n42097 , n42098 , n42099 , n42100 , n42101 , n42102 , n42103 , 
     n42104 , n42105 , n42106 , n42107 , n42108 , n42109 , n42110 , n42111 , n42112 , n42113 , 
     n42114 , n42115 , n42116 , n42117 , n42118 , n42119 , n42120 , n42121 , n42122 , n42123 , 
     n42124 , n42125 , n42126 , n42127 , n42128 , n42129 , n42130 , n42131 , n42132 , n42133 , 
     n42134 , n42135 , n42136 , n42137 , n42138 , n42139 , n42140 , n42141 , n42142 , n42143 , 
     n42144 , n42145 , n42146 , n42147 , n42148 , n42149 , n42150 , n42151 , n42152 , n42153 , 
     n42154 , n42155 , n42156 , n42157 , n42158 , n42159 , n42160 , n42161 , n42162 , n42163 , 
     n42164 , n42165 , n42166 , n42167 , n42168 , n42169 , n42170 , n42171 , n42172 , n42173 , 
     n42174 , n42175 , n42176 , n42177 , n42178 , n42179 , n42180 , n42181 , n42182 , n42183 , 
     n42184 , n42185 , n42186 , n42187 , n42188 , n42189 , n42190 , n42191 , n42192 , n42193 , 
     n42194 , n42195 , n42196 , n42197 , n42198 , n42199 , n42200 , n42201 , n42202 , n42203 , 
     n42204 , n42205 , n42206 , n42207 , n42208 , n42209 , n42210 , n42211 , n42212 , n42213 , 
     n42214 , n42215 , n42216 , n42217 , n42218 , n42219 , n42220 , n42221 , n42222 , n42223 , 
     n42224 , n42225 , n42226 , n42227 , n42228 , n42229 , n42230 , n42231 , n42232 , n42233 , 
     n42234 , n42235 , n42236 , n42237 , n42238 , n42239 , n42240 , n42241 , n42242 , n42243 , 
     n42244 , n42245 , n42246 , n42247 , n42248 , n42249 , n42250 , n42251 , n42252 , n42253 , 
     n42254 , n42255 , n42256 , n42257 , n42258 , n42259 , n42260 , n42261 , n42262 , n42263 , 
     n42264 , n42265 , n42266 , n42267 , n42268 , n42269 , n42270 , n42271 , n42272 , n42273 , 
     n42274 , n42275 , n42276 , n42277 , n42278 , n42279 , n42280 , n42281 , n42282 , n42283 , 
     n42284 , n42285 , n42286 , n42287 , n42288 , n42289 , n42290 , n42291 , n42292 , n42293 , 
     n42294 , n42295 , n42296 , n42297 , n42298 , n42299 , n42300 , n42301 , n42302 , n42303 , 
     n42304 , n42305 , n42306 , n42307 , n42308 , n42309 , n42310 , n42311 , n42312 , n42313 , 
     n42314 , n42315 , n42316 , n42317 , n42318 , n42319 , n42320 , n42321 , n42322 , n42323 , 
     n42324 , n42325 , n42326 , n42327 , n42328 , n42329 , n42330 , n42331 , n42332 , n42333 , 
     n42334 , n42335 , n42336 , n42337 , n42338 , n42339 , n42340 , n42341 , n42342 , n42343 , 
     n42344 , n42345 , n42346 , n42347 , n42348 , n42349 , n42350 , n42351 , n42352 , n42353 , 
     n42354 , n42355 , n42356 , n42357 , n42358 , n42359 , n42360 , n42361 , n42362 , n42363 , 
     n42364 , n42365 , n42366 , n42367 , n42368 , n42369 , n42370 , n42371 , n42372 , n42373 , 
     n42374 , n42375 , n42376 , n42377 , n42378 , n42379 , n42380 , n42381 , n42382 , n42383 , 
     n42384 , n42385 , n42386 , n42387 , n42388 , n42389 , n42390 , n42391 , n42392 , n42393 , 
     n42394 , n42395 , n42396 , n42397 , n42398 , n42399 , n42400 , n42401 , n42402 , n42403 , 
     n42404 , n42405 , n42406 , n42407 , n42408 , n42409 , n42410 , n42411 , n42412 , n42413 , 
     n42414 , n42415 , n42416 , n42417 , n42418 , n42419 , n42420 , n42421 , n42422 , n42423 , 
     n42424 , n42425 , n42426 , n42427 , n42428 , n42429 , n42430 , n42431 , n42432 , n42433 , 
     n42434 , n42435 , n42436 , n42437 , n42438 , n42439 , n42440 , n42441 , n42442 , n42443 , 
     n42444 , n42445 , n42446 , n42447 , n42448 , n42449 , n42450 , n42451 , n42452 , n42453 , 
     n42454 , n42455 , n42456 , n42457 , n42458 , n42459 , n42460 , n42461 , n42462 , n42463 , 
     n42464 , n42465 , n42466 , n42467 , n42468 , n42469 , n42470 , n42471 , n42472 , n42473 , 
     n42474 , n42475 , n42476 , n42477 , n42478 , n42479 , n42480 , n42481 , n42482 , n42483 , 
     n42484 , n42485 , n42486 , n42487 , n42488 , n42489 , n42490 , n42491 , n42492 , n42493 , 
     n42494 , n42495 , n42496 , n42497 , n42498 , n42499 , n42500 , n42501 , n42502 , n42503 , 
     n42504 , n42505 , n42506 , n42507 , n42508 , n42509 , n42510 , n42511 , n42512 , n42513 , 
     n42514 , n42515 , n42516 , n42517 , n42518 , n42519 , n42520 , n42521 , n42522 , n42523 , 
     n42524 , n42525 , n42526 , n42527 , n42528 , n42529 , n42530 , n42531 , n42532 , n42533 , 
     n42534 , n42535 , n42536 , n42537 , n42538 , n42539 , n42540 , n42541 , n42542 , n42543 , 
     n42544 , n42545 , n42546 , n42547 , n42548 , n42549 , n42550 , n42551 , n42552 , n42553 , 
     n42554 , n42555 , n42556 , n42557 , n42558 , n42559 , n42560 , n42561 , n42562 , n42563 , 
     n42564 , n42565 , n42566 , n42567 , n42568 , n42569 , n42570 , n42571 , n42572 , n42573 , 
     n42574 , n42575 , n42576 , n42577 , n42578 , n42579 , n42580 , n42581 , n42582 , n42583 , 
     n42584 , n42585 , n42586 , n42587 , n42588 , n42589 , n42590 , n42591 , n42592 , n42593 , 
     n42594 , n42595 , n42596 , n42597 , n42598 , n42599 , n42600 , n42601 , n42602 , n42603 , 
     n42604 , n42605 , n42606 , n42607 , n42608 , n42609 , n42610 , n42611 , n42612 , n42613 , 
     n42614 , n42615 , n42616 , n42617 , n42618 , n42619 , n42620 , n42621 , n42622 , n42623 , 
     n42624 , n42625 , n42626 , n42627 , n42628 , n42629 , n42630 , n42631 , n42632 , n42633 , 
     n42634 , n42635 , n42636 , n42637 , n42638 , n42639 , n42640 , n42641 , n42642 , n42643 , 
     n42644 , n42645 , n42646 , n42647 , n42648 , n42649 , n42650 , n42651 , n42652 , n42653 , 
     n42654 , n42655 , n42656 , n42657 , n42658 , n42659 , n42660 , n42661 , n42662 , n42663 , 
     n42664 , n42665 , n42666 , n42667 , n42668 , n42669 , n42670 , n42671 , n42672 , n42673 , 
     n42674 , n42675 , n42676 , n42677 , n42678 , n42679 , n42680 , n42681 , n42682 , n42683 , 
     n42684 , n42685 , n42686 , n42687 , n42688 , n42689 , n42690 , n42691 , n42692 , n42693 , 
     n42694 , n42695 , n42696 , n42697 , n42698 , n42699 , n42700 , n42701 , n42702 , n42703 , 
     n42704 , n42705 , n42706 , n42707 , n42708 , n42709 , n42710 , n42711 , n42712 , n42713 , 
     n42714 , n42715 , n42716 , n42717 , n42718 , n42719 , n42720 , n42721 , n42722 , n42723 , 
     n42724 , n42725 , n42726 , n42727 , n42728 , n42729 , n42730 , n42731 , n42732 , n42733 , 
     n42734 , n42735 , n42736 , n42737 , n42738 , n42739 , n42740 , n42741 , n42742 , n42743 , 
     n42744 , n42745 , n42746 , n42747 , n42748 , n42749 , n42750 , n42751 , n42752 , n42753 , 
     n42754 , n42755 , n42756 , n42757 , n42758 , n42759 , n42760 , n42761 , n42762 , n42763 , 
     n42764 , n42765 , n42766 , n42767 , n42768 , n42769 , n42770 , n42771 , n42772 , n42773 , 
     n42774 , n42775 , n42776 , n42777 , n42778 , n42779 , n42780 , n42781 , n42782 , n42783 , 
     n42784 , n42785 , n42786 , n42787 , n42788 , n42789 , n42790 , n42791 , n42792 , n42793 , 
     n42794 , n42795 , n42796 , n42797 , n42798 , n42799 , n42800 , n42801 , n42802 , n42803 , 
     n42804 , n42805 , n42806 , n42807 , n42808 , n42809 , n42810 , n42811 , n42812 , n42813 , 
     n42814 , n42815 , n42816 , n42817 , n42818 , n42819 , n42820 , n42821 , n42822 , n42823 , 
     n42824 , n42825 , n42826 , n42827 , n42828 , n42829 , n42830 , n42831 , n42832 , n42833 , 
     n42834 , n42835 , n42836 , n42837 , n42838 , n42839 , n42840 , n42841 , n42842 , n42843 , 
     n42844 , n42845 , n42846 , n42847 , n42848 , n42849 , n42850 , n42851 , n42852 , n42853 , 
     n42854 , n42855 , n42856 , n42857 , n42858 , n42859 , n42860 , n42861 , n42862 , n42863 , 
     n42864 , n42865 , n42866 , n42867 , n42868 , n42869 , n42870 , n42871 , n42872 , n42873 , 
     n42874 , n42875 , n42876 , n42877 , n42878 , n42879 , n42880 , n42881 , n42882 , n42883 , 
     n42884 , n42885 , n42886 , n42887 , n42888 , n42889 , n42890 , n42891 , n42892 , n42893 , 
     n42894 , n42895 , n42896 , n42897 , n42898 , n42899 , n42900 , n42901 , n42902 , n42903 , 
     n42904 , n42905 , n42906 , n42907 , n42908 , n42909 , n42910 , n42911 , n42912 , n42913 , 
     n42914 , n42915 , n42916 , n42917 , n42918 , n42919 , n42920 , n42921 , n42922 , n42923 , 
     n42924 , n42925 , n42926 , n42927 , n42928 , n42929 , n42930 , n42931 , n42932 , n42933 , 
     n42934 , n42935 , n42936 , n42937 , n42938 , n42939 , n42940 , n42941 , n42942 , n42943 , 
     n42944 , n42945 , n42946 , n42947 , n42948 , n42949 , n42950 , n42951 , n42952 , n42953 , 
     n42954 , n42955 , n42956 , n42957 , n42958 , n42959 , n42960 , n42961 , n42962 , n42963 , 
     n42964 , n42965 , n42966 , n42967 , n42968 , n42969 , n42970 , n42971 , n42972 , n42973 , 
     n42974 , n42975 , n42976 , n42977 , n42978 , n42979 , n42980 , n42981 , n42982 , n42983 , 
     n42984 , n42985 , n42986 , n42987 , n42988 , n42989 , n42990 , n42991 , n42992 , n42993 , 
     n42994 , n42995 , n42996 , n42997 , n42998 , n42999 , n43000 , n43001 , n43002 , n43003 , 
     n43004 , n43005 , n43006 , n43007 , n43008 , n43009 , n43010 , n43011 , n43012 , n43013 , 
     n43014 , n43015 , n43016 , n43017 , n43018 , n43019 , n43020 , n43021 , n43022 , n43023 , 
     n43024 , n43025 , n43026 , n43027 , n43028 , n43029 , n43030 , n43031 , n43032 , n43033 , 
     n43034 , n43035 , n43036 , n43037 , n43038 , n43039 , n43040 , n43041 , n43042 , n43043 , 
     n43044 , n43045 , n43046 , n43047 , n43048 , n43049 , n43050 , n43051 , n43052 , n43053 , 
     n43054 , n43055 , n43056 , n43057 , n43058 , n43059 , n43060 , n43061 , n43062 , n43063 , 
     n43064 , n43065 , n43066 , n43067 , n43068 , n43069 , n43070 , n43071 , n43072 , n43073 , 
     n43074 , n43075 , n43076 , n43077 , n43078 , n43079 , n43080 , n43081 , n43082 , n43083 , 
     n43084 , n43085 , n43086 , n43087 , n43088 , n43089 , n43090 , n43091 , n43092 , n43093 , 
     n43094 , n43095 , n43096 , n43097 , n43098 , n43099 , n43100 , n43101 , n43102 , n43103 , 
     n43104 , n43105 , n43106 , n43107 , n43108 , n43109 , n43110 , n43111 , n43112 , n43113 , 
     n43114 , n43115 , n43116 , n43117 , n43118 , n43119 , n43120 , n43121 , n43122 , n43123 , 
     n43124 , n43125 , n43126 , n43127 , n43128 , n43129 , n43130 , n43131 , n43132 , n43133 , 
     n43134 , n43135 , n43136 , n43137 , n43138 , n43139 , n43140 , n43141 , n43142 , n43143 , 
     n43144 , n43145 , n43146 , n43147 , n43148 , n43149 , n43150 , n43151 , n43152 , n43153 , 
     n43154 , n43155 , n43156 , n43157 , n43158 , n43159 , n43160 , n43161 , n43162 , n43163 , 
     n43164 , n43165 , n43166 , n43167 , n43168 , n43169 , n43170 , n43171 , n43172 , n43173 , 
     n43174 , n43175 , n43176 , n43177 , n43178 , n43179 , n43180 , n43181 , n43182 , n43183 , 
     n43184 , n43185 , n43186 , n43187 , n43188 , n43189 , n43190 , n43191 , n43192 , n43193 , 
     n43194 , n43195 , n43196 , n43197 , n43198 , n43199 , n43200 , n43201 , n43202 , n43203 , 
     n43204 , n43205 , n43206 , n43207 , n43208 , n43209 , n43210 , n43211 , n43212 , n43213 , 
     n43214 , n43215 , n43216 , n43217 , n43218 , n43219 , n43220 , n43221 , n43222 , n43223 , 
     n43224 , n43225 , n43226 , n43227 , n43228 , n43229 , n43230 , n43231 , n43232 , n43233 , 
     n43234 , n43235 , n43236 , n43237 , n43238 , n43239 , n43240 , n43241 , n43242 , n43243 , 
     n43244 , n43245 , n43246 , n43247 , n43248 , n43249 , n43250 , n43251 , n43252 , n43253 , 
     n43254 , n43255 , n43256 , n43257 , n43258 , n43259 , n43260 , n43261 , n43262 , n43263 , 
     n43264 , n43265 , n43266 , n43267 , n43268 , n43269 , n43270 , n43271 , n43272 , n43273 , 
     n43274 , n43275 , n43276 , n43277 , n43278 , n43279 , n43280 , n43281 , n43282 , n43283 , 
     n43284 , n43285 , n43286 , n43287 , n43288 , n43289 , n43290 , n43291 , n43292 , n43293 , 
     n43294 , n43295 , n43296 , n43297 , n43298 , n43299 , n43300 , n43301 , n43302 , n43303 , 
     n43304 , n43305 , n43306 , n43307 , n43308 , n43309 , n43310 , n43311 , n43312 , n43313 , 
     n43314 , n43315 , n43316 , n43317 , n43318 , n43319 , n43320 , n43321 , n43322 , n43323 , 
     n43324 , n43325 , n43326 , n43327 , n43328 , n43329 , n43330 , n43331 , n43332 , n43333 , 
     n43334 , n43335 , n43336 , n43337 , n43338 , n43339 , n43340 , n43341 , n43342 , n43343 , 
     n43344 , n43345 , n43346 , n43347 , n43348 , n43349 , n43350 , n43351 , n43352 , n43353 , 
     n43354 , n43355 , n43356 , n43357 , n43358 , n43359 , n43360 , n43361 , n43362 , n43363 , 
     n43364 , n43365 , n43366 , n43367 , n43368 , n43369 , n43370 , n43371 , n43372 , n43373 , 
     n43374 , n43375 , n43376 , n43377 , n43378 , n43379 , n43380 , n43381 , n43382 , n43383 , 
     n43384 , n43385 , n43386 , n43387 , n43388 , n43389 , n43390 , n43391 , n43392 , n43393 , 
     n43394 , n43395 , n43396 , n43397 , n43398 , n43399 , n43400 , n43401 , n43402 , n43403 , 
     n43404 , n43405 , n43406 , n43407 , n43408 , n43409 , n43410 , n43411 , n43412 , n43413 , 
     n43414 , n43415 , n43416 , n43417 , n43418 , n43419 , n43420 , n43421 , n43422 , n43423 , 
     n43424 , n43425 , n43426 , n43427 , n43428 , n43429 , n43430 , n43431 , n43432 , n43433 , 
     n43434 , n43435 , n43436 , n43437 , n43438 , n43439 , n43440 , n43441 , n43442 , n43443 , 
     n43444 , n43445 , n43446 , n43447 , n43448 , n43449 , n43450 , n43451 , n43452 , n43453 , 
     n43454 , n43455 , n43456 , n43457 , n43458 , n43459 , n43460 , n43461 , n43462 , n43463 , 
     n43464 , n43465 , n43466 , n43467 , n43468 , n43469 , n43470 , n43471 , n43472 , n43473 , 
     n43474 , n43475 , n43476 , n43477 , n43478 , n43479 , n43480 , n43481 , n43482 , n43483 , 
     n43484 , n43485 , n43486 , n43487 , n43488 , n43489 , n43490 , n43491 , n43492 , n43493 , 
     n43494 , n43495 , n43496 , n43497 , n43498 , n43499 , n43500 , n43501 , n43502 , n43503 , 
     n43504 , n43505 , n43506 , n43507 , n43508 , n43509 , n43510 , n43511 , n43512 , n43513 , 
     n43514 , n43515 , n43516 , n43517 , n43518 , n43519 , n43520 , n43521 , n43522 , n43523 , 
     n43524 , n43525 , n43526 , n43527 , n43528 , n43529 , n43530 , n43531 , n43532 , n43533 , 
     n43534 , n43535 , n43536 , n43537 , n43538 , n43539 , n43540 , n43541 , n43542 , n43543 , 
     n43544 , n43545 , n43546 , n43547 , n43548 , n43549 , n43550 , n43551 , n43552 , n43553 , 
     n43554 , n43555 , n43556 , n43557 , n43558 , n43559 , n43560 , n43561 , n43562 , n43563 , 
     n43564 , n43565 , n43566 , n43567 , n43568 , n43569 , n43570 , n43571 , n43572 , n43573 , 
     n43574 , n43575 , n43576 , n43577 , n43578 , n43579 , n43580 , n43581 , n43582 , n43583 , 
     n43584 , n43585 , n43586 , n43587 , n43588 , n43589 , n43590 , n43591 , n43592 , n43593 , 
     n43594 , n43595 , n43596 , n43597 , n43598 , n43599 , n43600 , n43601 , n43602 , n43603 , 
     n43604 , n43605 , n43606 , n43607 , n43608 , n43609 , n43610 , n43611 , n43612 , n43613 , 
     n43614 , n43615 , n43616 , n43617 , n43618 , n43619 , n43620 , n43621 , n43622 , n43623 , 
     n43624 , n43625 , n43626 , n43627 , n43628 , n43629 , n43630 , n43631 , n43632 , n43633 , 
     n43634 , n43635 , n43636 , n43637 , n43638 , n43639 , n43640 , n43641 , n43642 , n43643 , 
     n43644 , n43645 , n43646 , n43647 , n43648 , n43649 , n43650 , n43651 , n43652 , n43653 , 
     n43654 , n43655 , n43656 , n43657 , n43658 , n43659 , n43660 , n43661 , n43662 , n43663 , 
     n43664 , n43665 , n43666 , n43667 , n43668 , n43669 , n43670 , n43671 , n43672 , n43673 , 
     n43674 , n43675 , n43676 , n43677 , n43678 , n43679 , n43680 , n43681 , n43682 , n43683 , 
     n43684 , n43685 , n43686 , n43687 , n43688 , n43689 , n43690 , n43691 , n43692 , n43693 , 
     n43694 , n43695 , n43696 , n43697 , n43698 , n43699 , n43700 , n43701 , n43702 , n43703 , 
     n43704 , n43705 , n43706 , n43707 , n43708 , n43709 , n43710 , n43711 , n43712 , n43713 , 
     n43714 , n43715 , n43716 , n43717 , n43718 , n43719 , n43720 , n43721 , n43722 , n43723 , 
     n43724 , n43725 , n43726 , n43727 , n43728 , n43729 , n43730 , n43731 , n43732 , n43733 , 
     n43734 , n43735 , n43736 , n43737 , n43738 , n43739 , n43740 , n43741 , n43742 , n43743 , 
     n43744 , n43745 , n43746 , n43747 , n43748 , n43749 , n43750 , n43751 , n43752 , n43753 , 
     n43754 , n43755 , n43756 , n43757 , n43758 , n43759 , n43760 , n43761 , n43762 , n43763 , 
     n43764 , n43765 , n43766 , n43767 , n43768 , n43769 , n43770 , n43771 , n43772 , n43773 , 
     n43774 , n43775 , n43776 , n43777 , n43778 , n43779 , n43780 , n43781 , n43782 , n43783 , 
     n43784 , n43785 , n43786 , n43787 , n43788 , n43789 , n43790 , n43791 , n43792 , n43793 , 
     n43794 , n43795 , n43796 , n43797 , n43798 , n43799 , n43800 , n43801 , n43802 , n43803 , 
     n43804 , n43805 , n43806 , n43807 , n43808 , n43809 , n43810 , n43811 , n43812 , n43813 , 
     n43814 , n43815 , n43816 , n43817 , n43818 , n43819 , n43820 , n43821 , n43822 , n43823 , 
     n43824 , n43825 , n43826 , n43827 , n43828 , n43829 , n43830 , n43831 , n43832 , n43833 , 
     n43834 , n43835 , n43836 , n43837 , n43838 , n43839 , n43840 , n43841 , n43842 , n43843 , 
     n43844 , n43845 , n43846 , n43847 , n43848 , n43849 , n43850 , n43851 , n43852 , n43853 , 
     n43854 , n43855 , n43856 , n43857 , n43858 , n43859 , n43860 , n43861 , n43862 , n43863 , 
     n43864 , n43865 , n43866 , n43867 , n43868 , n43869 , n43870 , n43871 , n43872 , n43873 , 
     n43874 , n43875 , n43876 , n43877 , n43878 , n43879 , n43880 , n43881 , n43882 , n43883 , 
     n43884 , n43885 , n43886 , n43887 , n43888 , n43889 , n43890 , n43891 , n43892 , n43893 , 
     n43894 , n43895 , n43896 , n43897 , n43898 , n43899 , n43900 , n43901 , n43902 , n43903 , 
     n43904 , n43905 , n43906 , n43907 , n43908 , n43909 , n43910 , n43911 , n43912 , n43913 , 
     n43914 , n43915 , n43916 , n43917 , n43918 , n43919 , n43920 , n43921 , n43922 , n43923 , 
     n43924 , n43925 , n43926 , n43927 , n43928 , n43929 , n43930 , n43931 , n43932 , n43933 , 
     n43934 , n43935 , n43936 , n43937 , n43938 , n43939 , n43940 , n43941 , n43942 , n43943 , 
     n43944 , n43945 , n43946 , n43947 , n43948 , n43949 , n43950 , n43951 , n43952 , n43953 , 
     n43954 , n43955 , n43956 , n43957 , n43958 , n43959 , n43960 , n43961 , n43962 , n43963 , 
     n43964 , n43965 , n43966 , n43967 , n43968 , n43969 , n43970 , n43971 , n43972 , n43973 , 
     n43974 , n43975 , n43976 , n43977 , n43978 , n43979 , n43980 , n43981 , n43982 , n43983 , 
     n43984 , n43985 , n43986 , n43987 , n43988 , n43989 , n43990 , n43991 , n43992 , n43993 , 
     n43994 , n43995 , n43996 , n43997 , n43998 , n43999 , n44000 , n44001 , n44002 , n44003 , 
     n44004 , n44005 , n44006 , n44007 , n44008 , n44009 , n44010 , n44011 , n44012 , n44013 , 
     n44014 , n44015 , n44016 , n44017 , n44018 , n44019 , n44020 , n44021 , n44022 , n44023 , 
     n44024 , n44025 , n44026 , n44027 , n44028 , n44029 , n44030 , n44031 , n44032 , n44033 , 
     n44034 , n44035 , n44036 , n44037 , n44038 , n44039 , n44040 , n44041 , n44042 , n44043 , 
     n44044 , n44045 , n44046 , n44047 , n44048 , n44049 , n44050 , n44051 , n44052 , n44053 , 
     n44054 , n44055 , n44056 , n44057 , n44058 , n44059 , n44060 , n44061 , n44062 , n44063 , 
     n44064 , n44065 , n44066 , n44067 , n44068 , n44069 , n44070 , n44071 , n44072 , n44073 , 
     n44074 , n44075 , n44076 , n44077 , n44078 , n44079 , n44080 , n44081 , n44082 , n44083 , 
     n44084 , n44085 , n44086 , n44087 , n44088 , n44089 , n44090 , n44091 , n44092 , n44093 , 
     n44094 , n44095 , n44096 , n44097 , n44098 , n44099 , n44100 , n44101 , n44102 , n44103 , 
     n44104 , n44105 , n44106 , n44107 , n44108 , n44109 , n44110 , n44111 , n44112 , n44113 , 
     n44114 , n44115 , n44116 , n44117 , n44118 , n44119 , n44120 , n44121 , n44122 , n44123 , 
     n44124 , n44125 , n44126 , n44127 , n44128 , n44129 , n44130 , n44131 , n44132 , n44133 , 
     n44134 , n44135 , n44136 , n44137 , n44138 , n44139 , n44140 , n44141 , n44142 , n44143 , 
     n44144 , n44145 , n44146 , n44147 , n44148 , n44149 , n44150 , n44151 , n44152 , n44153 , 
     n44154 , n44155 , n44156 , n44157 , n44158 , n44159 , n44160 , n44161 , n44162 , n44163 , 
     n44164 , n44165 , n44166 , n44167 , n44168 , n44169 , n44170 , n44171 , n44172 , n44173 , 
     n44174 , n44175 , n44176 , n44177 , n44178 , n44179 , n44180 , n44181 , n44182 , n44183 , 
     n44184 , n44185 , n44186 , n44187 , n44188 , n44189 , n44190 , n44191 , n44192 , n44193 , 
     n44194 , n44195 , n44196 , n44197 , n44198 , n44199 , n44200 , n44201 , n44202 , n44203 , 
     n44204 , n44205 , n44206 , n44207 , n44208 , n44209 , n44210 , n44211 , n44212 , n44213 , 
     n44214 , n44215 , n44216 , n44217 , n44218 , n44219 , n44220 , n44221 , n44222 , n44223 , 
     n44224 , n44225 , n44226 , n44227 , n44228 , n44229 , n44230 , n44231 , n44232 , n44233 , 
     n44234 , n44235 , n44236 , n44237 , n44238 , n44239 , n44240 , n44241 , n44242 , n44243 , 
     n44244 , n44245 , n44246 , n44247 , n44248 , n44249 , n44250 , n44251 , n44252 , n44253 , 
     n44254 , n44255 , n44256 , n44257 , n44258 , n44259 , n44260 , n44261 , n44262 , n44263 , 
     n44264 , n44265 , n44266 , n44267 , n44268 , n44269 , n44270 , n44271 , n44272 , n44273 , 
     n44274 , n44275 , n44276 , n44277 , n44278 , n44279 , n44280 , n44281 , n44282 , n44283 , 
     n44284 , n44285 , n44286 , n44287 , n44288 , n44289 , n44290 , n44291 , n44292 , n44293 , 
     n44294 , n44295 , n44296 , n44297 , n44298 , n44299 , n44300 , n44301 , n44302 , n44303 , 
     n44304 , n44305 , n44306 , n44307 , n44308 , n44309 , n44310 , n44311 , n44312 , n44313 , 
     n44314 , n44315 , n44316 , n44317 , n44318 , n44319 , n44320 , n44321 , n44322 , n44323 , 
     n44324 , n44325 , n44326 , n44327 , n44328 , n44329 , n44330 , n44331 , n44332 , n44333 , 
     n44334 , n44335 , n44336 , n44337 , n44338 , n44339 , n44340 , n44341 , n44342 , n44343 , 
     n44344 , n44345 , n44346 , n44347 , n44348 , n44349 , n44350 , n44351 , n44352 , n44353 , 
     n44354 , n44355 , n44356 , n44357 , n44358 , n44359 , n44360 , n44361 , n44362 , n44363 , 
     n44364 , n44365 , n44366 , n44367 , n44368 , n44369 , n44370 , n44371 , n44372 , n44373 , 
     n44374 , n44375 , n44376 , n44377 , n44378 , n44379 , n44380 , n44381 , n44382 , n44383 , 
     n44384 , n44385 , n44386 , n44387 , n44388 , n44389 , n44390 , n44391 , n44392 , n44393 , 
     n44394 , n44395 , n44396 , n44397 , n44398 , n44399 , n44400 , n44401 , n44402 , n44403 , 
     n44404 , n44405 , n44406 , n44407 , n44408 , n44409 , n44410 , n44411 , n44412 , n44413 , 
     n44414 , n44415 , n44416 , n44417 , n44418 , n44419 , n44420 , n44421 , n44422 , n44423 , 
     n44424 , n44425 , n44426 , n44427 , n44428 , n44429 , n44430 , n44431 , n44432 , n44433 , 
     n44434 , n44435 , n44436 , n44437 , n44438 , n44439 , n44440 , n44441 , n44442 , n44443 , 
     n44444 , n44445 , n44446 , n44447 , n44448 , n44449 , n44450 , n44451 , n44452 , n44453 , 
     n44454 , n44455 , n44456 , n44457 , n44458 , n44459 , n44460 , n44461 , n44462 , n44463 , 
     n44464 , n44465 , n44466 , n44467 , n44468 , n44469 , n44470 , n44471 , n44472 , n44473 , 
     n44474 , n44475 , n44476 , n44477 , n44478 , n44479 , n44480 , n44481 , n44482 , n44483 , 
     n44484 , n44485 , n44486 , n44487 , n44488 , n44489 , n44490 , n44491 , n44492 , n44493 , 
     n44494 , n44495 , n44496 , n44497 , n44498 , n44499 , n44500 , n44501 , n44502 , n44503 , 
     n44504 , n44505 , n44506 , n44507 , n44508 , n44509 , n44510 , n44511 , n44512 , n44513 , 
     n44514 , n44515 , n44516 , n44517 , n44518 , n44519 , n44520 , n44521 , n44522 , n44523 , 
     n44524 , n44525 , n44526 , n44527 , n44528 , n44529 , n44530 , n44531 , n44532 , n44533 , 
     n44534 , n44535 , n44536 , n44537 , n44538 , n44539 , n44540 , n44541 , n44542 , n44543 , 
     n44544 , n44545 , n44546 , n44547 , n44548 , n44549 , n44550 , n44551 , n44552 , n44553 , 
     n44554 , n44555 , n44556 , n44557 , n44558 , n44559 , n44560 , n44561 , n44562 , n44563 , 
     n44564 , n44565 , n44566 , n44567 , n44568 , n44569 , n44570 , n44571 , n44572 , n44573 , 
     n44574 , n44575 , n44576 , n44577 , n44578 , n44579 , n44580 , n44581 , n44582 , n44583 , 
     n44584 , n44585 , n44586 , n44587 , n44588 , n44589 , n44590 , n44591 , n44592 , n44593 , 
     n44594 , n44595 , n44596 , n44597 , n44598 , n44599 , n44600 , n44601 , n44602 , n44603 , 
     n44604 , n44605 , n44606 , n44607 , n44608 , n44609 , n44610 , n44611 , n44612 , n44613 , 
     n44614 , n44615 , n44616 , n44617 , n44618 , n44619 , n44620 , n44621 , n44622 , n44623 , 
     n44624 , n44625 , n44626 , n44627 , n44628 , n44629 , n44630 , n44631 , n44632 , n44633 , 
     n44634 , n44635 , n44636 , n44637 , n44638 , n44639 , n44640 , n44641 , n44642 , n44643 , 
     n44644 , n44645 , n44646 , n44647 , n44648 , n44649 , n44650 , n44651 , n44652 , n44653 , 
     n44654 , n44655 , n44656 , n44657 , n44658 , n44659 , n44660 , n44661 , n44662 , n44663 , 
     n44664 , n44665 , n44666 , n44667 , n44668 , n44669 , n44670 , n44671 , n44672 , n44673 , 
     n44674 , n44675 , n44676 , n44677 , n44678 , n44679 , n44680 , n44681 , n44682 , n44683 , 
     n44684 , n44685 , n44686 , n44687 , n44688 , n44689 , n44690 , n44691 , n44692 , n44693 , 
     n44694 , n44695 , n44696 , n44697 , n44698 , n44699 , n44700 , n44701 , n44702 , n44703 , 
     n44704 , n44705 , n44706 , n44707 , n44708 , n44709 , n44710 , n44711 , n44712 , n44713 , 
     n44714 , n44715 , n44716 , n44717 , n44718 , n44719 , n44720 , n44721 , n44722 , n44723 , 
     n44724 , n44725 , n44726 , n44727 , n44728 , n44729 , n44730 , n44731 , n44732 , n44733 , 
     n44734 , n44735 , n44736 , n44737 , n44738 , n44739 , n44740 , n44741 , n44742 , n44743 , 
     n44744 , n44745 , n44746 , n44747 , n44748 , n44749 , n44750 , n44751 , n44752 , n44753 , 
     n44754 , n44755 , n44756 , n44757 , n44758 , n44759 , n44760 , n44761 , n44762 , n44763 , 
     n44764 , n44765 , n44766 , n44767 , n44768 , n44769 , n44770 , n44771 , n44772 , n44773 , 
     n44774 , n44775 , n44776 , n44777 , n44778 , n44779 , n44780 , n44781 , n44782 , n44783 , 
     n44784 , n44785 , n44786 , n44787 , n44788 , n44789 , n44790 , n44791 , n44792 , n44793 , 
     n44794 , n44795 , n44796 , n44797 , n44798 , n44799 , n44800 , n44801 , n44802 , n44803 , 
     n44804 , n44805 , n44806 , n44807 , n44808 , n44809 , n44810 , n44811 , n44812 , n44813 , 
     n44814 , n44815 , n44816 , n44817 , n44818 , n44819 , n44820 , n44821 , n44822 , n44823 , 
     n44824 , n44825 , n44826 , n44827 , n44828 , n44829 , n44830 , n44831 , n44832 , n44833 , 
     n44834 , n44835 , n44836 , n44837 , n44838 , n44839 , n44840 , n44841 , n44842 , n44843 , 
     n44844 , n44845 , n44846 , n44847 , n44848 , n44849 , n44850 , n44851 , n44852 , n44853 , 
     n44854 , n44855 , n44856 , n44857 , n44858 , n44859 , n44860 , n44861 , n44862 , n44863 , 
     n44864 , n44865 , n44866 , n44867 , n44868 , n44869 , n44870 , n44871 , n44872 , n44873 , 
     n44874 , n44875 , n44876 , n44877 , n44878 , n44879 , n44880 , n44881 , n44882 , n44883 , 
     n44884 , n44885 , n44886 , n44887 , n44888 , n44889 , n44890 , n44891 , n44892 , n44893 , 
     n44894 , n44895 , n44896 , n44897 , n44898 , n44899 , n44900 , n44901 , n44902 , n44903 , 
     n44904 , n44905 , n44906 , n44907 , n44908 , n44909 , n44910 , n44911 , n44912 , n44913 , 
     n44914 , n44915 , n44916 , n44917 , n44918 , n44919 , n44920 , n44921 , n44922 , n44923 , 
     n44924 , n44925 , n44926 , n44927 , n44928 , n44929 , n44930 , n44931 , n44932 , n44933 , 
     n44934 , n44935 , n44936 , n44937 , n44938 , n44939 , n44940 , n44941 , n44942 , n44943 , 
     n44944 , n44945 , n44946 , n44947 , n44948 , n44949 , n44950 , n44951 , n44952 , n44953 , 
     n44954 , n44955 , n44956 , n44957 , n44958 , n44959 , n44960 , n44961 , n44962 , n44963 , 
     n44964 , n44965 , n44966 , n44967 , n44968 , n44969 , n44970 , n44971 , n44972 , n44973 , 
     n44974 , n44975 , n44976 , n44977 , n44978 , n44979 , n44980 , n44981 , n44982 , n44983 , 
     n44984 , n44985 , n44986 , n44987 , n44988 , n44989 , n44990 , n44991 , n44992 , n44993 , 
     n44994 , n44995 , n44996 , n44997 , n44998 , n44999 , n45000 , n45001 , n45002 , n45003 , 
     n45004 , n45005 , n45006 , n45007 , n45008 , n45009 , n45010 , n45011 , n45012 , n45013 , 
     n45014 , n45015 , n45016 , n45017 , n45018 , n45019 , n45020 , n45021 , n45022 , n45023 , 
     n45024 , n45025 , n45026 , n45027 , n45028 , n45029 , n45030 , n45031 , n45032 , n45033 , 
     n45034 , n45035 , n45036 , n45037 , n45038 , n45039 , n45040 , n45041 , n45042 , n45043 , 
     n45044 , n45045 , n45046 , n45047 , n45048 , n45049 , n45050 , n45051 , n45052 , n45053 , 
     n45054 , n45055 , n45056 , n45057 , n45058 , n45059 , n45060 , n45061 , n45062 , n45063 , 
     n45064 , n45065 , n45066 , n45067 , n45068 , n45069 , n45070 , n45071 , n45072 , n45073 , 
     n45074 , n45075 , n45076 , n45077 , n45078 , n45079 , n45080 , n45081 , n45082 , n45083 , 
     n45084 , n45085 , n45086 , n45087 , n45088 , n45089 , n45090 , n45091 , n45092 , n45093 , 
     n45094 , n45095 , n45096 , n45097 , n45098 , n45099 , n45100 , n45101 , n45102 , n45103 , 
     n45104 , n45105 , n45106 , n45107 , n45108 , n45109 , n45110 , n45111 , n45112 , n45113 , 
     n45114 , n45115 , n45116 , n45117 , n45118 , n45119 , n45120 , n45121 , n45122 , n45123 , 
     n45124 , n45125 , n45126 , n45127 , n45128 , n45129 , n45130 , n45131 , n45132 , n45133 , 
     n45134 , n45135 , n45136 , n45137 , n45138 , n45139 , n45140 , n45141 , n45142 , n45143 , 
     n45144 , n45145 , n45146 , n45147 , n45148 , n45149 , n45150 , n45151 , n45152 , n45153 , 
     n45154 , n45155 , n45156 , n45157 , n45158 , n45159 , n45160 , n45161 , n45162 , n45163 , 
     n45164 , n45165 , n45166 , n45167 , n45168 , n45169 , n45170 , n45171 , n45172 , n45173 , 
     n45174 , n45175 , n45176 , n45177 , n45178 , n45179 , n45180 , n45181 , n45182 , n45183 , 
     n45184 , n45185 , n45186 , n45187 , n45188 , n45189 , n45190 , n45191 , n45192 , n45193 , 
     n45194 , n45195 , n45196 , n45197 , n45198 , n45199 , n45200 , n45201 , n45202 , n45203 , 
     n45204 , n45205 , n45206 , n45207 , n45208 , n45209 , n45210 , n45211 , n45212 , n45213 , 
     n45214 , n45215 , n45216 , n45217 , n45218 , n45219 , n45220 , n45221 , n45222 , n45223 , 
     n45224 , n45225 , n45226 , n45227 , n45228 , n45229 , n45230 , n45231 , n45232 , n45233 , 
     n45234 , n45235 , n45236 , n45237 , n45238 , n45239 , n45240 , n45241 , n45242 , n45243 , 
     n45244 , n45245 , n45246 , n45247 , n45248 , n45249 , n45250 , n45251 , n45252 , n45253 , 
     n45254 , n45255 , n45256 , n45257 , n45258 , n45259 , n45260 , n45261 , n45262 , n45263 , 
     n45264 , n45265 , n45266 , n45267 , n45268 , n45269 , n45270 , n45271 , n45272 , n45273 , 
     n45274 , n45275 , n45276 , n45277 , n45278 , n45279 , n45280 , n45281 , n45282 , n45283 , 
     n45284 , n45285 , n45286 , n45287 , n45288 , n45289 , n45290 , n45291 , n45292 , n45293 , 
     n45294 , n45295 , n45296 , n45297 , n45298 , n45299 , n45300 , n45301 , n45302 , n45303 , 
     n45304 , n45305 , n45306 , n45307 , n45308 , n45309 , n45310 , n45311 , n45312 , n45313 , 
     n45314 , n45315 , n45316 , n45317 , n45318 , n45319 , n45320 , n45321 , n45322 , n45323 , 
     n45324 , n45325 , n45326 , n45327 , n45328 , n45329 , n45330 , n45331 , n45332 , n45333 , 
     n45334 , n45335 , n45336 , n45337 , n45338 , n45339 , n45340 , n45341 , n45342 , n45343 , 
     n45344 , n45345 , n45346 , n45347 , n45348 , n45349 , n45350 , n45351 , n45352 , n45353 , 
     n45354 , n45355 , n45356 , n45357 , n45358 , n45359 , n45360 , n45361 , n45362 , n45363 , 
     n45364 , n45365 , n45366 , n45367 , n45368 , n45369 , n45370 , n45371 , n45372 , n45373 , 
     n45374 , n45375 , n45376 , n45377 , n45378 , n45379 , n45380 , n45381 , n45382 , n45383 , 
     n45384 , n45385 , n45386 , n45387 , n45388 , n45389 , n45390 , n45391 , n45392 , n45393 , 
     n45394 , n45395 , n45396 , n45397 , n45398 , n45399 , n45400 , n45401 , n45402 , n45403 , 
     n45404 , n45405 , n45406 , n45407 , n45408 , n45409 , n45410 , n45411 , n45412 , n45413 , 
     n45414 , n45415 , n45416 , n45417 , n45418 , n45419 , n45420 , n45421 , n45422 , n45423 , 
     n45424 , n45425 , n45426 , n45427 , n45428 , n45429 , n45430 , n45431 , n45432 , n45433 , 
     n45434 , n45435 , n45436 , n45437 , n45438 , n45439 , n45440 , n45441 , n45442 , n45443 , 
     n45444 , n45445 , n45446 , n45447 , n45448 , n45449 , n45450 , n45451 , n45452 , n45453 , 
     n45454 , n45455 , n45456 , n45457 , n45458 , n45459 , n45460 , n45461 , n45462 , n45463 , 
     n45464 , n45465 , n45466 , n45467 , n45468 , n45469 , n45470 , n45471 , n45472 , n45473 , 
     n45474 , n45475 , n45476 , n45477 , n45478 , n45479 , n45480 , n45481 , n45482 , n45483 , 
     n45484 , n45485 , n45486 , n45487 , n45488 , n45489 , n45490 , n45491 , n45492 , n45493 , 
     n45494 , n45495 , n45496 , n45497 , n45498 , n45499 , n45500 , n45501 , n45502 , n45503 , 
     n45504 , n45505 , n45506 , n45507 , n45508 , n45509 , n45510 , n45511 , n45512 , n45513 , 
     n45514 , n45515 , n45516 , n45517 , n45518 , n45519 , n45520 , n45521 , n45522 , n45523 , 
     n45524 , n45525 , n45526 , n45527 , n45528 , n45529 , n45530 , n45531 , n45532 , n45533 , 
     n45534 , n45535 , n45536 , n45537 , n45538 , n45539 , n45540 , n45541 , n45542 , n45543 , 
     n45544 , n45545 , n45546 , n45547 , n45548 , n45549 , n45550 , n45551 , n45552 , n45553 , 
     n45554 , n45555 , n45556 , n45557 , n45558 , n45559 , n45560 , n45561 , n45562 , n45563 , 
     n45564 , n45565 , n45566 , n45567 , n45568 , n45569 , n45570 , n45571 , n45572 , n45573 , 
     n45574 , n45575 , n45576 , n45577 , n45578 , n45579 , n45580 , n45581 , n45582 , n45583 , 
     n45584 , n45585 , n45586 , n45587 , n45588 , n45589 , n45590 , n45591 , n45592 , n45593 , 
     n45594 , n45595 , n45596 , n45597 , n45598 , n45599 , n45600 , n45601 , n45602 , n45603 , 
     n45604 , n45605 , n45606 , n45607 , n45608 , n45609 , n45610 , n45611 , n45612 , n45613 , 
     n45614 , n45615 , n45616 , n45617 , n45618 , n45619 , n45620 , n45621 , n45622 , n45623 , 
     n45624 , n45625 , n45626 , n45627 , n45628 , n45629 , n45630 , n45631 , n45632 , n45633 , 
     n45634 , n45635 , n45636 , n45637 , n45638 , n45639 , n45640 , n45641 , n45642 , n45643 , 
     n45644 , n45645 , n45646 , n45647 , n45648 , n45649 , n45650 , n45651 , n45652 , n45653 , 
     n45654 , n45655 , n45656 , n45657 , n45658 , n45659 , n45660 , n45661 , n45662 , n45663 , 
     n45664 , n45665 , n45666 , n45667 , n45668 , n45669 , n45670 , n45671 , n45672 , n45673 , 
     n45674 , n45675 , n45676 , n45677 , n45678 , n45679 , n45680 , n45681 , n45682 , n45683 , 
     n45684 , n45685 , n45686 , n45687 , n45688 , n45689 , n45690 , n45691 , n45692 , n45693 , 
     n45694 , n45695 , n45696 , n45697 , n45698 , n45699 , n45700 , n45701 , n45702 , n45703 , 
     n45704 , n45705 , n45706 , n45707 , n45708 , n45709 , n45710 , n45711 , n45712 , n45713 , 
     n45714 , n45715 , n45716 , n45717 , n45718 , n45719 , n45720 , n45721 , n45722 , n45723 , 
     n45724 , n45725 , n45726 , n45727 , n45728 , n45729 , n45730 , n45731 , n45732 , n45733 , 
     n45734 , n45735 , n45736 , n45737 , n45738 , n45739 , n45740 , n45741 , n45742 , n45743 , 
     n45744 , n45745 , n45746 , n45747 , n45748 , n45749 , n45750 , n45751 , n45752 , n45753 , 
     n45754 , n45755 , n45756 , n45757 , n45758 , n45759 , n45760 , n45761 , n45762 , n45763 , 
     n45764 , n45765 , n45766 , n45767 , n45768 , n45769 , n45770 , n45771 , n45772 , n45773 , 
     n45774 , n45775 , n45776 , n45777 , n45778 , n45779 , n45780 , n45781 , n45782 , n45783 , 
     n45784 , n45785 , n45786 , n45787 , n45788 , n45789 , n45790 , n45791 , n45792 , n45793 , 
     n45794 , n45795 , n45796 , n45797 , n45798 , n45799 , n45800 , n45801 , n45802 , n45803 , 
     n45804 , n45805 , n45806 , n45807 , n45808 , n45809 , n45810 , n45811 , n45812 , n45813 , 
     n45814 , n45815 , n45816 , n45817 , n45818 , n45819 , n45820 , n45821 , n45822 , n45823 , 
     n45824 , n45825 , n45826 , n45827 , n45828 , n45829 , n45830 , n45831 , n45832 , n45833 , 
     n45834 , n45835 , n45836 , n45837 , n45838 , n45839 , n45840 , n45841 , n45842 , n45843 , 
     n45844 , n45845 , n45846 , n45847 , n45848 , n45849 , n45850 , n45851 , n45852 , n45853 , 
     n45854 , n45855 , n45856 , n45857 , n45858 , n45859 , n45860 , n45861 , n45862 , n45863 , 
     n45864 , n45865 , n45866 , n45867 , n45868 , n45869 , n45870 , n45871 , n45872 , n45873 , 
     n45874 , n45875 , n45876 , n45877 , n45878 , n45879 , n45880 , n45881 , n45882 , n45883 , 
     n45884 , n45885 , n45886 , n45887 , n45888 , n45889 , n45890 , n45891 , n45892 , n45893 , 
     n45894 , n45895 , n45896 , n45897 , n45898 , n45899 , n45900 , n45901 , n45902 , n45903 , 
     n45904 , n45905 , n45906 , n45907 , n45908 , n45909 , n45910 , n45911 , n45912 , n45913 , 
     n45914 , n45915 , n45916 , n45917 , n45918 , n45919 , n45920 , n45921 , n45922 , n45923 , 
     n45924 , n45925 , n45926 , n45927 , n45928 , n45929 , n45930 , n45931 , n45932 , n45933 , 
     n45934 , n45935 , n45936 , n45937 , n45938 , n45939 , n45940 , n45941 , n45942 , n45943 , 
     n45944 , n45945 , n45946 , n45947 , n45948 , n45949 , n45950 , n45951 , n45952 , n45953 , 
     n45954 , n45955 , n45956 , n45957 , n45958 , n45959 , n45960 , n45961 , n45962 , n45963 , 
     n45964 , n45965 , n45966 , n45967 , n45968 , n45969 , n45970 , n45971 , n45972 , n45973 , 
     n45974 , n45975 , n45976 , n45977 , n45978 , n45979 , n45980 , n45981 , n45982 , n45983 , 
     n45984 , n45985 , n45986 , n45987 , n45988 , n45989 , n45990 , n45991 , n45992 , n45993 , 
     n45994 , n45995 , n45996 , n45997 , n45998 , n45999 , n46000 , n46001 , n46002 , n46003 , 
     n46004 , n46005 , n46006 , n46007 , n46008 , n46009 , n46010 , n46011 , n46012 , n46013 , 
     n46014 , n46015 , n46016 , n46017 , n46018 , n46019 , n46020 , n46021 , n46022 , n46023 , 
     n46024 , n46025 , n46026 , n46027 , n46028 , n46029 , n46030 , n46031 , n46032 , n46033 , 
     n46034 , n46035 , n46036 , n46037 , n46038 , n46039 , n46040 , n46041 , n46042 , n46043 , 
     n46044 , n46045 , n46046 , n46047 , n46048 , n46049 , n46050 , n46051 , n46052 , n46053 , 
     n46054 , n46055 , n46056 , n46057 , n46058 , n46059 , n46060 , n46061 , n46062 , n46063 , 
     n46064 , n46065 , n46066 , n46067 , n46068 , n46069 , n46070 , n46071 , n46072 , n46073 , 
     n46074 , n46075 , n46076 , n46077 , n46078 , n46079 , n46080 , n46081 , n46082 , n46083 , 
     n46084 , n46085 , n46086 , n46087 , n46088 , n46089 , n46090 , n46091 , n46092 , n46093 , 
     n46094 , n46095 , n46096 , n46097 , n46098 , n46099 , n46100 , n46101 , n46102 , n46103 , 
     n46104 , n46105 , n46106 , n46107 , n46108 , n46109 , n46110 , n46111 , n46112 , n46113 , 
     n46114 , n46115 , n46116 , n46117 , n46118 , n46119 , n46120 , n46121 , n46122 , n46123 , 
     n46124 , n46125 , n46126 , n46127 , n46128 , n46129 , n46130 , n46131 , n46132 , n46133 , 
     n46134 , n46135 , n46136 , n46137 , n46138 , n46139 , n46140 , n46141 , n46142 , n46143 , 
     n46144 , n46145 , n46146 , n46147 , n46148 , n46149 , n46150 , n46151 , n46152 , n46153 , 
     n46154 , n46155 , n46156 , n46157 , n46158 , n46159 , n46160 , n46161 , n46162 , n46163 , 
     n46164 , n46165 , n46166 , n46167 , n46168 , n46169 , n46170 , n46171 , n46172 , n46173 , 
     n46174 , n46175 , n46176 , n46177 , n46178 , n46179 , n46180 , n46181 , n46182 , n46183 , 
     n46184 , n46185 , n46186 , n46187 , n46188 , n46189 , n46190 , n46191 , n46192 , n46193 , 
     n46194 , n46195 , n46196 , n46197 , n46198 , n46199 , n46200 , n46201 , n46202 , n46203 , 
     n46204 , n46205 , n46206 , n46207 , n46208 , n46209 , n46210 , n46211 , n46212 , n46213 , 
     n46214 , n46215 , n46216 , n46217 , n46218 , n46219 , n46220 , n46221 , n46222 , n46223 , 
     n46224 , n46225 , n46226 , n46227 , n46228 , n46229 , n46230 , n46231 , n46232 , n46233 , 
     n46234 , n46235 , n46236 , n46237 , n46238 , n46239 , n46240 , n46241 , n46242 , n46243 , 
     n46244 , n46245 , n46246 , n46247 , n46248 , n46249 , n46250 , n46251 , n46252 , n46253 , 
     n46254 , n46255 , n46256 , n46257 , n46258 , n46259 , n46260 , n46261 , n46262 , n46263 , 
     n46264 , n46265 , n46266 , n46267 , n46268 , n46269 , n46270 , n46271 , n46272 , n46273 , 
     n46274 , n46275 , n46276 , n46277 , n46278 , n46279 , n46280 , n46281 , n46282 , n46283 , 
     n46284 , n46285 , n46286 , n46287 , n46288 , n46289 , n46290 , n46291 , n46292 , n46293 , 
     n46294 , n46295 , n46296 , n46297 , n46298 , n46299 , n46300 , n46301 , n46302 , n46303 , 
     n46304 , n46305 , n46306 , n46307 , n46308 , n46309 , n46310 , n46311 , n46312 , n46313 , 
     n46314 , n46315 , n46316 , n46317 , n46318 , n46319 , n46320 , n46321 , n46322 , n46323 , 
     n46324 , n46325 , n46326 , n46327 , n46328 , n46329 , n46330 , n46331 , n46332 , n46333 , 
     n46334 , n46335 , n46336 , n46337 , n46338 , n46339 , n46340 , n46341 , n46342 , n46343 , 
     n46344 , n46345 , n46346 , n46347 , n46348 , n46349 , n46350 , n46351 , n46352 , n46353 , 
     n46354 , n46355 , n46356 , n46357 , n46358 , n46359 , n46360 , n46361 , n46362 , n46363 , 
     n46364 , n46365 , n46366 , n46367 , n46368 , n46369 , n46370 , n46371 , n46372 , n46373 , 
     n46374 , n46375 , n46376 , n46377 , n46378 , n46379 , n46380 , n46381 , n46382 , n46383 , 
     n46384 , n46385 , n46386 , n46387 , n46388 , n46389 , n46390 , n46391 , n46392 , n46393 , 
     n46394 , n46395 , n46396 , n46397 , n46398 , n46399 , n46400 , n46401 , n46402 , n46403 , 
     n46404 , n46405 , n46406 , n46407 , n46408 , n46409 , n46410 , n46411 , n46412 , n46413 , 
     n46414 , n46415 , n46416 , n46417 , n46418 , n46419 , n46420 , n46421 , n46422 , n46423 , 
     n46424 , n46425 , n46426 , n46427 , n46428 , n46429 , n46430 , n46431 , n46432 , n46433 , 
     n46434 , n46435 , n46436 , n46437 , n46438 , n46439 , n46440 , n46441 , n46442 , n46443 , 
     n46444 , n46445 , n46446 , n46447 , n46448 , n46449 , n46450 , n46451 , n46452 , n46453 , 
     n46454 , n46455 , n46456 , n46457 , n46458 , n46459 , n46460 , n46461 , n46462 , n46463 , 
     n46464 , n46465 , n46466 , n46467 , n46468 , n46469 , n46470 , n46471 , n46472 , n46473 , 
     n46474 , n46475 , n46476 , n46477 , n46478 , n46479 , n46480 , n46481 , n46482 , n46483 , 
     n46484 , n46485 , n46486 , n46487 , n46488 , n46489 , n46490 , n46491 , n46492 , n46493 , 
     n46494 , n46495 , n46496 , n46497 , n46498 , n46499 , n46500 , n46501 , n46502 , n46503 , 
     n46504 , n46505 , n46506 , n46507 , n46508 , n46509 , n46510 , n46511 , n46512 , n46513 , 
     n46514 , n46515 , n46516 , n46517 , n46518 , n46519 , n46520 , n46521 , n46522 , n46523 , 
     n46524 , n46525 , n46526 , n46527 , n46528 , n46529 , n46530 , n46531 , n46532 , n46533 , 
     n46534 , n46535 , n46536 , n46537 , n46538 , n46539 , n46540 , n46541 , n46542 , n46543 , 
     n46544 , n46545 , n46546 , n46547 , n46548 , n46549 , n46550 , n46551 , n46552 , n46553 , 
     n46554 , n46555 , n46556 , n46557 , n46558 , n46559 , n46560 , n46561 , n46562 , n46563 , 
     n46564 , n46565 , n46566 , n46567 , n46568 , n46569 , n46570 , n46571 , n46572 , n46573 , 
     n46574 , n46575 , n46576 , n46577 , n46578 , n46579 , n46580 , n46581 , n46582 , n46583 , 
     n46584 , n46585 , n46586 , n46587 , n46588 , n46589 , n46590 , n46591 , n46592 , n46593 , 
     n46594 , n46595 , n46596 , n46597 , n46598 , n46599 , n46600 , n46601 , n46602 , n46603 , 
     n46604 , n46605 , n46606 , n46607 , n46608 , n46609 , n46610 , n46611 , n46612 , n46613 , 
     n46614 , n46615 , n46616 , n46617 , n46618 , n46619 , n46620 , n46621 , n46622 , n46623 , 
     n46624 , n46625 , n46626 , n46627 , n46628 , n46629 , n46630 , n46631 , n46632 , n46633 , 
     n46634 , n46635 , n46636 , n46637 , n46638 , n46639 , n46640 , n46641 , n46642 , n46643 , 
     n46644 , n46645 , n46646 , n46647 , n46648 , n46649 , n46650 , n46651 , n46652 , n46653 , 
     n46654 , n46655 , n46656 , n46657 , n46658 , n46659 , n46660 , n46661 , n46662 , n46663 , 
     n46664 , n46665 , n46666 , n46667 , n46668 , n46669 , n46670 , n46671 , n46672 , n46673 , 
     n46674 , n46675 , n46676 , n46677 , n46678 , n46679 , n46680 , n46681 , n46682 , n46683 , 
     n46684 , n46685 , n46686 , n46687 , n46688 , n46689 , n46690 , n46691 , n46692 , n46693 , 
     n46694 , n46695 , n46696 , n46697 , n46698 , n46699 , n46700 , n46701 , n46702 , n46703 , 
     n46704 , n46705 , n46706 , n46707 , n46708 , n46709 , n46710 , n46711 , n46712 , n46713 , 
     n46714 , n46715 , n46716 , n46717 , n46718 , n46719 , n46720 , n46721 , n46722 , n46723 , 
     n46724 , n46725 , n46726 , n46727 , n46728 , n46729 , n46730 , n46731 , n46732 , n46733 , 
     n46734 , n46735 , n46736 , n46737 , n46738 , n46739 , n46740 , n46741 , n46742 , n46743 , 
     n46744 , n46745 , n46746 , n46747 , n46748 , n46749 , n46750 , n46751 , n46752 , n46753 , 
     n46754 , n46755 , n46756 , n46757 , n46758 , n46759 , n46760 , n46761 , n46762 , n46763 , 
     n46764 , n46765 , n46766 , n46767 , n46768 , n46769 , n46770 , n46771 , n46772 , n46773 , 
     n46774 , n46775 , n46776 , n46777 , n46778 , n46779 , n46780 , n46781 , n46782 , n46783 , 
     n46784 , n46785 , n46786 , n46787 , n46788 , n46789 , n46790 , n46791 , n46792 , n46793 , 
     n46794 , n46795 , n46796 , n46797 , n46798 , n46799 , n46800 , n46801 , n46802 , n46803 , 
     n46804 , n46805 , n46806 , n46807 , n46808 , n46809 , n46810 , n46811 , n46812 , n46813 , 
     n46814 , n46815 , n46816 , n46817 , n46818 , n46819 , n46820 , n46821 , n46822 , n46823 , 
     n46824 , n46825 , n46826 , n46827 , n46828 , n46829 , n46830 , n46831 , n46832 , n46833 , 
     n46834 , n46835 , n46836 , n46837 , n46838 , n46839 , n46840 , n46841 , n46842 , n46843 , 
     n46844 , n46845 , n46846 , n46847 , n46848 , n46849 , n46850 , n46851 , n46852 , n46853 , 
     n46854 , n46855 , n46856 , n46857 , n46858 , n46859 , n46860 , n46861 , n46862 , n46863 , 
     n46864 , n46865 , n46866 , n46867 , n46868 , n46869 , n46870 , n46871 , n46872 , n46873 , 
     n46874 , n46875 , n46876 , n46877 , n46878 , n46879 , n46880 , n46881 , n46882 , n46883 , 
     n46884 , n46885 , n46886 , n46887 , n46888 , n46889 , n46890 , n46891 , n46892 , n46893 , 
     n46894 , n46895 , n46896 , n46897 , n46898 , n46899 , n46900 , n46901 , n46902 , n46903 , 
     n46904 , n46905 , n46906 , n46907 , n46908 , n46909 , n46910 , n46911 , n46912 , n46913 , 
     n46914 , n46915 , n46916 , n46917 , n46918 , n46919 , n46920 , n46921 , n46922 , n46923 , 
     n46924 , n46925 , n46926 , n46927 , n46928 , n46929 , n46930 , n46931 , n46932 , n46933 , 
     n46934 , n46935 , n46936 , n46937 , n46938 , n46939 , n46940 , n46941 , n46942 , n46943 , 
     n46944 , n46945 , n46946 , n46947 , n46948 , n46949 , n46950 , n46951 , n46952 , n46953 , 
     n46954 , n46955 , n46956 , n46957 , n46958 , n46959 , n46960 , n46961 , n46962 , n46963 , 
     n46964 , n46965 , n46966 , n46967 , n46968 , n46969 , n46970 , n46971 , n46972 , n46973 , 
     n46974 , n46975 , n46976 , n46977 , n46978 , n46979 , n46980 , n46981 , n46982 , n46983 , 
     n46984 , n46985 , n46986 , n46987 , n46988 , n46989 , n46990 , n46991 , n46992 , n46993 , 
     n46994 , n46995 , n46996 , n46997 , n46998 , n46999 , n47000 , n47001 , n47002 , n47003 , 
     n47004 , n47005 , n47006 , n47007 , n47008 , n47009 , n47010 , n47011 , n47012 , n47013 , 
     n47014 , n47015 , n47016 , n47017 , n47018 , n47019 , n47020 , n47021 , n47022 , n47023 , 
     n47024 , n47025 , n47026 , n47027 , n47028 , n47029 , n47030 , n47031 , n47032 , n47033 , 
     n47034 , n47035 , n47036 , n47037 , n47038 , n47039 , n47040 , n47041 , n47042 , n47043 , 
     n47044 , n47045 , n47046 , n47047 , n47048 , n47049 , n47050 , n47051 , n47052 , n47053 , 
     n47054 , n47055 , n47056 , n47057 , n47058 , n47059 , n47060 , n47061 , n47062 , n47063 , 
     n47064 , n47065 , n47066 , n47067 , n47068 , n47069 , n47070 , n47071 , n47072 , n47073 , 
     n47074 , n47075 , n47076 , n47077 , n47078 , n47079 , n47080 , n47081 , n47082 , n47083 , 
     n47084 , n47085 , n47086 , n47087 , n47088 , n47089 , n47090 , n47091 , n47092 , n47093 , 
     n47094 , n47095 , n47096 , n47097 , n47098 , n47099 , n47100 , n47101 , n47102 , n47103 , 
     n47104 , n47105 , n47106 , n47107 , n47108 , n47109 , n47110 , n47111 , n47112 , n47113 , 
     n47114 , n47115 , n47116 , n47117 , n47118 , n47119 , n47120 , n47121 , n47122 , n47123 , 
     n47124 , n47125 , n47126 , n47127 , n47128 , n47129 , n47130 , n47131 , n47132 , n47133 , 
     n47134 , n47135 , n47136 , n47137 , n47138 , n47139 , n47140 , n47141 , n47142 , n47143 , 
     n47144 , n47145 , n47146 , n47147 , n47148 , n47149 , n47150 , n47151 , n47152 , n47153 , 
     n47154 , n47155 , n47156 , n47157 , n47158 , n47159 , n47160 , n47161 , n47162 , n47163 , 
     n47164 , n47165 , n47166 , n47167 , n47168 , n47169 , n47170 , n47171 , n47172 , n47173 , 
     n47174 , n47175 , n47176 , n47177 , n47178 , n47179 , n47180 , n47181 , n47182 , n47183 , 
     n47184 , n47185 , n47186 , n47187 , n47188 , n47189 , n47190 , n47191 , n47192 , n47193 , 
     n47194 , n47195 , n47196 , n47197 , n47198 , n47199 , n47200 , n47201 , n47202 , n47203 , 
     n47204 , n47205 , n47206 , n47207 , n47208 , n47209 , n47210 , n47211 , n47212 , n47213 , 
     n47214 , n47215 , n47216 , n47217 , n47218 , n47219 , n47220 , n47221 , n47222 , n47223 , 
     n47224 , n47225 , n47226 , n47227 , n47228 , n47229 , n47230 , n47231 , n47232 , n47233 , 
     n47234 , n47235 , n47236 , n47237 , n47238 , n47239 , n47240 , n47241 , n47242 , n47243 , 
     n47244 , n47245 , n47246 , n47247 , n47248 , n47249 , n47250 , n47251 , n47252 , n47253 , 
     n47254 , n47255 , n47256 , n47257 , n47258 , n47259 , n47260 , n47261 , n47262 , n47263 , 
     n47264 , n47265 , n47266 , n47267 , n47268 , n47269 , n47270 , n47271 , n47272 , n47273 , 
     n47274 , n47275 , n47276 , n47277 , n47278 , n47279 , n47280 , n47281 , n47282 , n47283 , 
     n47284 , n47285 , n47286 , n47287 , n47288 , n47289 , n47290 , n47291 , n47292 , n47293 , 
     n47294 , n47295 , n47296 , n47297 , n47298 , n47299 , n47300 , n47301 , n47302 , n47303 , 
     n47304 , n47305 , n47306 , n47307 , n47308 , n47309 , n47310 , n47311 , n47312 , n47313 , 
     n47314 , n47315 , n47316 , n47317 , n47318 , n47319 , n47320 , n47321 , n47322 , n47323 , 
     n47324 , n47325 , n47326 , n47327 , n47328 , n47329 , n47330 , n47331 , n47332 , n47333 , 
     n47334 , n47335 , n47336 , n47337 , n47338 , n47339 , n47340 , n47341 , n47342 , n47343 , 
     n47344 , n47345 , n47346 , n47347 , n47348 , n47349 , n47350 , n47351 , n47352 , n47353 , 
     n47354 , n47355 , n47356 , n47357 , n47358 , n47359 , n47360 , n47361 , n47362 , n47363 , 
     n47364 , n47365 , n47366 , n47367 , n47368 , n47369 , n47370 , n47371 , n47372 , n47373 , 
     n47374 , n47375 , n47376 , n47377 , n47378 , n47379 , n47380 , n47381 , n47382 , n47383 , 
     n47384 , n47385 , n47386 , n47387 , n47388 , n47389 , n47390 , n47391 , n47392 , n47393 , 
     n47394 , n47395 , n47396 , n47397 , n47398 , n47399 , n47400 , n47401 , n47402 , n47403 , 
     n47404 , n47405 , n47406 , n47407 , n47408 , n47409 , n47410 , n47411 , n47412 , n47413 , 
     n47414 , n47415 , n47416 , n47417 , n47418 , n47419 , n47420 , n47421 , n47422 , n47423 , 
     n47424 , n47425 , n47426 , n47427 , n47428 , n47429 , n47430 , n47431 , n47432 , n47433 , 
     n47434 , n47435 , n47436 , n47437 , n47438 , n47439 , n47440 , n47441 , n47442 , n47443 , 
     n47444 , n47445 , n47446 , n47447 , n47448 , n47449 , n47450 , n47451 , n47452 , n47453 , 
     n47454 , n47455 , n47456 , n47457 , n47458 , n47459 , n47460 , n47461 , n47462 , n47463 , 
     n47464 , n47465 , n47466 , n47467 , n47468 , n47469 , n47470 , n47471 , n47472 , n47473 , 
     n47474 , n47475 , n47476 , n47477 , n47478 , n47479 , n47480 , n47481 , n47482 , n47483 , 
     n47484 , n47485 , n47486 , n47487 , n47488 , n47489 , n47490 , n47491 , n47492 , n47493 , 
     n47494 , n47495 , n47496 , n47497 , n47498 , n47499 , n47500 , n47501 , n47502 , n47503 , 
     n47504 , n47505 , n47506 , n47507 , n47508 , n47509 , n47510 , n47511 , n47512 , n47513 , 
     n47514 , n47515 , n47516 , n47517 , n47518 , n47519 , n47520 , n47521 , n47522 , n47523 , 
     n47524 , n47525 , n47526 , n47527 , n47528 , n47529 , n47530 , n47531 , n47532 , n47533 , 
     n47534 , n47535 , n47536 , n47537 , n47538 , n47539 , n47540 , n47541 , n47542 , n47543 , 
     n47544 , n47545 , n47546 , n47547 , n47548 , n47549 , n47550 , n47551 , n47552 , n47553 , 
     n47554 , n47555 , n47556 , n47557 , n47558 , n47559 , n47560 , n47561 , n47562 , n47563 , 
     n47564 , n47565 , n47566 , n47567 , n47568 , n47569 , n47570 , n47571 , n47572 , n47573 , 
     n47574 , n47575 , n47576 , n47577 , n47578 , n47579 , n47580 , n47581 , n47582 , n47583 , 
     n47584 , n47585 , n47586 , n47587 , n47588 , n47589 , n47590 , n47591 , n47592 , n47593 , 
     n47594 , n47595 , n47596 , n47597 , n47598 , n47599 , n47600 , n47601 , n47602 , n47603 , 
     n47604 , n47605 , n47606 , n47607 , n47608 , n47609 , n47610 , n47611 , n47612 , n47613 , 
     n47614 , n47615 , n47616 , n47617 , n47618 , n47619 , n47620 , n47621 , n47622 , n47623 , 
     n47624 , n47625 , n47626 , n47627 , n47628 , n47629 , n47630 , n47631 , n47632 , n47633 , 
     n47634 , n47635 , n47636 , n47637 , n47638 , n47639 , n47640 , n47641 , n47642 , n47643 , 
     n47644 , n47645 , n47646 , n47647 , n47648 , n47649 , n47650 , n47651 , n47652 , n47653 , 
     n47654 , n47655 , n47656 , n47657 , n47658 , n47659 , n47660 , n47661 , n47662 , n47663 , 
     n47664 , n47665 , n47666 , n47667 , n47668 , n47669 , n47670 , n47671 , n47672 , n47673 , 
     n47674 , n47675 , n47676 , n47677 , n47678 , n47679 , n47680 , n47681 , n47682 , n47683 , 
     n47684 , n47685 , n47686 , n47687 , n47688 , n47689 , n47690 , n47691 , n47692 , n47693 , 
     n47694 , n47695 , n47696 , n47697 , n47698 , n47699 , n47700 , n47701 , n47702 , n47703 , 
     n47704 , n47705 , n47706 , n47707 , n47708 , n47709 , n47710 , n47711 , n47712 , n47713 , 
     n47714 , n47715 , n47716 , n47717 , n47718 , n47719 , n47720 , n47721 , n47722 , n47723 , 
     n47724 , n47725 , n47726 , n47727 , n47728 , n47729 , n47730 , n47731 , n47732 , n47733 , 
     n47734 , n47735 , n47736 , n47737 , n47738 , n47739 , n47740 , n47741 , n47742 , n47743 , 
     n47744 , n47745 , n47746 , n47747 , n47748 , n47749 , n47750 , n47751 , n47752 , n47753 , 
     n47754 , n47755 , n47756 , n47757 , n47758 , n47759 , n47760 , n47761 , n47762 , n47763 , 
     n47764 , n47765 , n47766 , n47767 , n47768 , n47769 , n47770 , n47771 , n47772 , n47773 , 
     n47774 , n47775 , n47776 , n47777 , n47778 , n47779 , n47780 , n47781 , n47782 , n47783 , 
     n47784 , n47785 , n47786 , n47787 , n47788 , n47789 , n47790 , n47791 , n47792 , n47793 , 
     n47794 , n47795 , n47796 , n47797 , n47798 , n47799 , n47800 , n47801 , n47802 , n47803 , 
     n47804 , n47805 , n47806 , n47807 , n47808 , n47809 , n47810 , n47811 , n47812 , n47813 , 
     n47814 , n47815 , n47816 , n47817 , n47818 , n47819 , n47820 , n47821 , n47822 , n47823 , 
     n47824 , n47825 , n47826 , n47827 , n47828 , n47829 , n47830 , n47831 , n47832 , n47833 , 
     n47834 , n47835 , n47836 , n47837 , n47838 , n47839 , n47840 , n47841 , n47842 , n47843 , 
     n47844 , n47845 , n47846 , n47847 , n47848 , n47849 , n47850 , n47851 , n47852 , n47853 , 
     n47854 , n47855 , n47856 , n47857 , n47858 , n47859 , n47860 , n47861 , n47862 , n47863 , 
     n47864 , n47865 , n47866 , n47867 , n47868 , n47869 , n47870 , n47871 , n47872 , n47873 , 
     n47874 , n47875 , n47876 , n47877 , n47878 , n47879 , n47880 , n47881 , n47882 , n47883 , 
     n47884 , n47885 , n47886 , n47887 , n47888 , n47889 , n47890 , n47891 , n47892 , n47893 , 
     n47894 , n47895 , n47896 , n47897 , n47898 , n47899 , n47900 , n47901 , n47902 , n47903 , 
     n47904 , n47905 , n47906 , n47907 , n47908 , n47909 , n47910 , n47911 , n47912 , n47913 , 
     n47914 , n47915 , n47916 , n47917 , n47918 , n47919 , n47920 , n47921 , n47922 , n47923 , 
     n47924 , n47925 , n47926 , n47927 , n47928 , n47929 , n47930 , n47931 , n47932 , n47933 , 
     n47934 , n47935 , n47936 , n47937 , n47938 , n47939 , n47940 , n47941 , n47942 , n47943 , 
     n47944 , n47945 , n47946 , n47947 , n47948 , n47949 , n47950 , n47951 , n47952 , n47953 , 
     n47954 , n47955 , n47956 , n47957 , n47958 , n47959 , n47960 , n47961 , n47962 , n47963 , 
     n47964 , n47965 , n47966 , n47967 , n47968 , n47969 , n47970 , n47971 , n47972 , n47973 , 
     n47974 , n47975 , n47976 , n47977 , n47978 , n47979 , n47980 , n47981 , n47982 , n47983 , 
     n47984 , n47985 , n47986 , n47987 , n47988 , n47989 , n47990 , n47991 , n47992 , n47993 , 
     n47994 , n47995 , n47996 , n47997 , n47998 , n47999 , n48000 , n48001 , n48002 , n48003 , 
     n48004 , n48005 , n48006 , n48007 , n48008 , n48009 , n48010 , n48011 , n48012 , n48013 , 
     n48014 , n48015 , n48016 , n48017 , n48018 , n48019 , n48020 , n48021 , n48022 , n48023 , 
     n48024 , n48025 , n48026 , n48027 , n48028 , n48029 , n48030 , n48031 , n48032 , n48033 , 
     n48034 , n48035 , n48036 , n48037 , n48038 , n48039 , n48040 , n48041 , n48042 , n48043 , 
     n48044 , n48045 , n48046 , n48047 , n48048 , n48049 , n48050 , n48051 , n48052 , n48053 , 
     n48054 , n48055 , n48056 , n48057 , n48058 , n48059 , n48060 , n48061 , n48062 , n48063 , 
     n48064 , n48065 , n48066 , n48067 , n48068 , n48069 , n48070 , n48071 , n48072 , n48073 , 
     n48074 , n48075 , n48076 , n48077 , n48078 , n48079 , n48080 , n48081 , n48082 , n48083 , 
     n48084 , n48085 , n48086 , n48087 , n48088 , n48089 , n48090 , n48091 , n48092 , n48093 , 
     n48094 , n48095 , n48096 , n48097 , n48098 , n48099 , n48100 , n48101 , n48102 , n48103 , 
     n48104 , n48105 , n48106 , n48107 , n48108 , n48109 , n48110 , n48111 , n48112 , n48113 , 
     n48114 , n48115 , n48116 , n48117 , n48118 , n48119 , n48120 , n48121 , n48122 , n48123 , 
     n48124 , n48125 , n48126 , n48127 , n48128 , n48129 , n48130 , n48131 , n48132 , n48133 , 
     n48134 , n48135 , n48136 , n48137 , n48138 , n48139 , n48140 , n48141 , n48142 , n48143 , 
     n48144 , n48145 , n48146 , n48147 , n48148 , n48149 , n48150 , n48151 , n48152 , n48153 , 
     n48154 , n48155 , n48156 , n48157 , n48158 , n48159 , n48160 , n48161 , n48162 , n48163 , 
     n48164 , n48165 , n48166 , n48167 , n48168 , n48169 , n48170 , n48171 , n48172 , n48173 , 
     n48174 , n48175 , n48176 , n48177 , n48178 , n48179 , n48180 , n48181 , n48182 , n48183 , 
     n48184 , n48185 , n48186 , n48187 , n48188 , n48189 , n48190 , n48191 , n48192 , n48193 , 
     n48194 , n48195 , n48196 , n48197 , n48198 , n48199 , n48200 , n48201 , n48202 , n48203 , 
     n48204 , n48205 , n48206 , n48207 , n48208 , n48209 , n48210 , n48211 , n48212 , n48213 , 
     n48214 , n48215 , n48216 , n48217 , n48218 , n48219 , n48220 , n48221 , n48222 , n48223 , 
     n48224 , n48225 , n48226 , n48227 , n48228 , n48229 , n48230 , n48231 , n48232 , n48233 , 
     n48234 , n48235 , n48236 , n48237 , n48238 , n48239 , n48240 , n48241 , n48242 , n48243 , 
     n48244 , n48245 , n48246 , n48247 , n48248 , n48249 , n48250 , n48251 , n48252 , n48253 , 
     n48254 , n48255 , n48256 , n48257 , n48258 , n48259 , n48260 , n48261 , n48262 , n48263 , 
     n48264 , n48265 , n48266 , n48267 , n48268 , n48269 , n48270 , n48271 , n48272 , n48273 , 
     n48274 , n48275 , n48276 , n48277 , n48278 , n48279 , n48280 , n48281 , n48282 , n48283 , 
     n48284 , n48285 , n48286 , n48287 , n48288 , n48289 , n48290 , n48291 , n48292 , n48293 , 
     n48294 , n48295 , n48296 , n48297 , n48298 , n48299 , n48300 , n48301 , n48302 , n48303 , 
     n48304 , n48305 , n48306 , n48307 , n48308 , n48309 , n48310 , n48311 , n48312 , n48313 , 
     n48314 , n48315 , n48316 , n48317 , n48318 , n48319 , n48320 , n48321 , n48322 , n48323 , 
     n48324 , n48325 , n48326 , n48327 , n48328 , n48329 , n48330 , n48331 , n48332 , n48333 , 
     n48334 , n48335 , n48336 , n48337 , n48338 , n48339 , n48340 , n48341 , n48342 , n48343 , 
     n48344 , n48345 , n48346 , n48347 , n48348 , n48349 , n48350 , n48351 , n48352 , n48353 , 
     n48354 , n48355 , n48356 , n48357 , n48358 , n48359 , n48360 , n48361 , n48362 , n48363 , 
     n48364 , n48365 , n48366 , n48367 , n48368 , n48369 , n48370 , n48371 , n48372 , n48373 , 
     n48374 , n48375 , n48376 , n48377 , n48378 , n48379 , n48380 , n48381 , n48382 , n48383 , 
     n48384 , n48385 , n48386 , n48387 , n48388 , n48389 , n48390 , n48391 , n48392 , n48393 , 
     n48394 , n48395 , n48396 , n48397 , n48398 , n48399 , n48400 , n48401 , n48402 , n48403 , 
     n48404 , n48405 , n48406 , n48407 , n48408 , n48409 , n48410 , n48411 , n48412 , n48413 , 
     n48414 , n48415 , n48416 , n48417 , n48418 , n48419 , n48420 , n48421 , n48422 , n48423 , 
     n48424 , n48425 , n48426 , n48427 , n48428 , n48429 , n48430 , n48431 , n48432 , n48433 , 
     n48434 , n48435 , n48436 , n48437 , n48438 , n48439 , n48440 , n48441 , n48442 , n48443 , 
     n48444 , n48445 , n48446 , n48447 , n48448 , n48449 , n48450 , n48451 , n48452 , n48453 , 
     n48454 , n48455 , n48456 , n48457 , n48458 , n48459 , n48460 , n48461 , n48462 , n48463 , 
     n48464 , n48465 , n48466 , n48467 , n48468 , n48469 , n48470 , n48471 , n48472 , n48473 , 
     n48474 , n48475 , n48476 , n48477 , n48478 , n48479 , n48480 , n48481 , n48482 , n48483 , 
     n48484 , n48485 , n48486 , n48487 , n48488 , n48489 , n48490 , n48491 , n48492 , n48493 , 
     n48494 , n48495 , n48496 , n48497 , n48498 , n48499 , n48500 , n48501 , n48502 , n48503 , 
     n48504 , n48505 , n48506 , n48507 , n48508 , n48509 , n48510 , n48511 , n48512 , n48513 , 
     n48514 , n48515 , n48516 , n48517 , n48518 , n48519 , n48520 , n48521 , n48522 , n48523 , 
     n48524 , n48525 , n48526 , n48527 , n48528 , n48529 , n48530 , n48531 , n48532 , n48533 , 
     n48534 , n48535 , n48536 , n48537 , n48538 , n48539 , n48540 , n48541 , n48542 , n48543 , 
     n48544 , n48545 , n48546 , n48547 , n48548 , n48549 , n48550 , n48551 , n48552 , n48553 , 
     n48554 , n48555 , n48556 , n48557 , n48558 , n48559 , n48560 , n48561 , n48562 , n48563 , 
     n48564 , n48565 , n48566 , n48567 , n48568 , n48569 , n48570 , n48571 , n48572 , n48573 , 
     n48574 , n48575 , n48576 , n48577 , n48578 , n48579 , n48580 , n48581 , n48582 , n48583 , 
     n48584 , n48585 , n48586 , n48587 , n48588 , n48589 , n48590 , n48591 , n48592 , n48593 , 
     n48594 , n48595 , n48596 , n48597 , n48598 , n48599 , n48600 , n48601 , n48602 , n48603 , 
     n48604 , n48605 , n48606 , n48607 , n48608 , n48609 , n48610 , n48611 , n48612 , n48613 , 
     n48614 , n48615 , n48616 , n48617 , n48618 , n48619 , n48620 , n48621 , n48622 , n48623 , 
     n48624 , n48625 , n48626 , n48627 , n48628 , n48629 , n48630 , n48631 , n48632 , n48633 , 
     n48634 , n48635 , n48636 , n48637 , n48638 , n48639 , n48640 , n48641 , n48642 , n48643 , 
     n48644 , n48645 , n48646 , n48647 , n48648 , n48649 , n48650 , n48651 , n48652 , n48653 , 
     n48654 , n48655 , n48656 , n48657 , n48658 , n48659 , n48660 , n48661 , n48662 , n48663 , 
     n48664 , n48665 , n48666 , n48667 , n48668 , n48669 , n48670 , n48671 , n48672 , n48673 , 
     n48674 , n48675 , n48676 , n48677 , n48678 , n48679 , n48680 , n48681 , n48682 , n48683 , 
     n48684 , n48685 , n48686 , n48687 , n48688 , n48689 , n48690 , n48691 , n48692 , n48693 , 
     n48694 , n48695 , n48696 , n48697 , n48698 , n48699 , n48700 , n48701 , n48702 , n48703 , 
     n48704 , n48705 , n48706 , n48707 , n48708 , n48709 , n48710 , n48711 , n48712 , n48713 , 
     n48714 , n48715 , n48716 , n48717 , n48718 , n48719 , n48720 , n48721 , n48722 , n48723 , 
     n48724 , n48725 , n48726 , n48727 , n48728 , n48729 , n48730 , n48731 , n48732 , n48733 , 
     n48734 , n48735 , n48736 , n48737 , n48738 , n48739 , n48740 , n48741 , n48742 , n48743 , 
     n48744 , n48745 , n48746 , n48747 , n48748 , n48749 , n48750 , n48751 , n48752 , n48753 , 
     n48754 , n48755 , n48756 , n48757 , n48758 , n48759 , n48760 , n48761 , n48762 , n48763 , 
     n48764 , n48765 , n48766 , n48767 , n48768 , n48769 , n48770 , n48771 , n48772 , n48773 , 
     n48774 , n48775 , n48776 , n48777 , n48778 , n48779 , n48780 , n48781 , n48782 , n48783 , 
     n48784 , n48785 , n48786 , n48787 , n48788 , n48789 , n48790 , n48791 , n48792 , n48793 , 
     n48794 , n48795 , n48796 , n48797 , n48798 , n48799 , n48800 , n48801 , n48802 , n48803 , 
     n48804 , n48805 , n48806 , n48807 , n48808 , n48809 , n48810 , n48811 , n48812 , n48813 , 
     n48814 , n48815 , n48816 , n48817 , n48818 , n48819 , n48820 , n48821 , n48822 , n48823 , 
     n48824 , n48825 , n48826 , n48827 , n48828 , n48829 , n48830 , n48831 , n48832 , n48833 , 
     n48834 , n48835 , n48836 , n48837 , n48838 , n48839 , n48840 , n48841 , n48842 , n48843 , 
     n48844 , n48845 , n48846 , n48847 , n48848 , n48849 , n48850 , n48851 , n48852 , n48853 , 
     n48854 , n48855 , n48856 , n48857 , n48858 , n48859 , n48860 , n48861 , n48862 , n48863 , 
     n48864 , n48865 , n48866 , n48867 , n48868 , n48869 , n48870 , n48871 , n48872 , n48873 , 
     n48874 , n48875 , n48876 , n48877 , n48878 , n48879 , n48880 , n48881 , n48882 , n48883 , 
     n48884 , n48885 , n48886 , n48887 , n48888 , n48889 , n48890 , n48891 , n48892 , n48893 , 
     n48894 , n48895 , n48896 , n48897 , n48898 , n48899 , n48900 , n48901 , n48902 , n48903 , 
     n48904 , n48905 , n48906 , n48907 , n48908 , n48909 , n48910 , n48911 , n48912 , n48913 , 
     n48914 , n48915 , n48916 , n48917 , n48918 , n48919 , n48920 , n48921 , n48922 , n48923 , 
     n48924 , n48925 , n48926 , n48927 , n48928 , n48929 , n48930 , n48931 , n48932 , n48933 , 
     n48934 , n48935 , n48936 , n48937 , n48938 , n48939 , n48940 , n48941 , n48942 , n48943 , 
     n48944 , n48945 , n48946 , n48947 , n48948 , n48949 , n48950 , n48951 , n48952 , n48953 , 
     n48954 , n48955 , n48956 , n48957 , n48958 , n48959 , n48960 , n48961 , n48962 , n48963 , 
     n48964 , n48965 , n48966 , n48967 , n48968 , n48969 , n48970 , n48971 , n48972 , n48973 , 
     n48974 , n48975 , n48976 , n48977 , n48978 , n48979 , n48980 , n48981 , n48982 , n48983 , 
     n48984 , n48985 , n48986 , n48987 , n48988 , n48989 , n48990 , n48991 , n48992 , n48993 , 
     n48994 , n48995 , n48996 , n48997 , n48998 , n48999 , n49000 , n49001 , n49002 , n49003 , 
     n49004 , n49005 , n49006 , n49007 , n49008 , n49009 , n49010 , n49011 , n49012 , n49013 , 
     n49014 , n49015 , n49016 , n49017 , n49018 , n49019 , n49020 , n49021 , n49022 , n49023 , 
     n49024 , n49025 , n49026 , n49027 , n49028 , n49029 , n49030 , n49031 , n49032 , n49033 , 
     n49034 , n49035 , n49036 , n49037 , n49038 , n49039 , n49040 , n49041 , n49042 , n49043 , 
     n49044 , n49045 , n49046 , n49047 , n49048 , n49049 , n49050 , n49051 , n49052 , n49053 , 
     n49054 , n49055 , n49056 , n49057 , n49058 , n49059 , n49060 , n49061 , n49062 , n49063 , 
     n49064 , n49065 , n49066 , n49067 , n49068 , n49069 , n49070 , n49071 , n49072 , n49073 , 
     n49074 , n49075 , n49076 , n49077 , n49078 , n49079 , n49080 , n49081 , n49082 , n49083 , 
     n49084 , n49085 , n49086 , n49087 , n49088 , n49089 , n49090 , n49091 , n49092 , n49093 , 
     n49094 , n49095 , n49096 , n49097 , n49098 , n49099 , n49100 , n49101 , n49102 , n49103 , 
     n49104 , n49105 , n49106 , n49107 , n49108 , n49109 , n49110 , n49111 , n49112 , n49113 , 
     n49114 , n49115 , n49116 , n49117 , n49118 , n49119 , n49120 , n49121 , n49122 , n49123 , 
     n49124 , n49125 , n49126 , n49127 , n49128 , n49129 , n49130 , n49131 , n49132 , n49133 , 
     n49134 , n49135 , n49136 , n49137 , n49138 , n49139 , n49140 , n49141 , n49142 , n49143 , 
     n49144 , n49145 , n49146 , n49147 , n49148 , n49149 , n49150 , n49151 , n49152 , n49153 , 
     n49154 , n49155 , n49156 , n49157 , n49158 , n49159 , n49160 , n49161 , n49162 , n49163 , 
     n49164 , n49165 , n49166 , n49167 , n49168 , n49169 , n49170 , n49171 , n49172 , n49173 , 
     n49174 , n49175 , n49176 , n49177 , n49178 , n49179 , n49180 , n49181 , n49182 , n49183 , 
     n49184 , n49185 , n49186 , n49187 , n49188 , n49189 , n49190 , n49191 , n49192 , n49193 , 
     n49194 , n49195 , n49196 , n49197 , n49198 , n49199 , n49200 , n49201 , n49202 , n49203 , 
     n49204 , n49205 , n49206 , n49207 , n49208 , n49209 , n49210 , n49211 , n49212 , n49213 , 
     n49214 , n49215 , n49216 , n49217 , n49218 , n49219 , n49220 , n49221 , n49222 , n49223 , 
     n49224 , n49225 , n49226 , n49227 , n49228 , n49229 , n49230 , n49231 , n49232 , n49233 , 
     n49234 , n49235 , n49236 , n49237 , n49238 , n49239 , n49240 , n49241 , n49242 , n49243 , 
     n49244 , n49245 , n49246 , n49247 , n49248 , n49249 , n49250 , n49251 , n49252 , n49253 , 
     n49254 , n49255 , n49256 , n49257 , n49258 , n49259 , n49260 , n49261 , n49262 , n49263 , 
     n49264 , n49265 , n49266 , n49267 , n49268 , n49269 , n49270 , n49271 , n49272 , n49273 , 
     n49274 , n49275 , n49276 , n49277 , n49278 , n49279 , n49280 , n49281 , n49282 , n49283 , 
     n49284 , n49285 , n49286 , n49287 , n49288 , n49289 , n49290 , n49291 , n49292 , n49293 , 
     n49294 , n49295 , n49296 , n49297 , n49298 , n49299 , n49300 , n49301 , n49302 , n49303 , 
     n49304 , n49305 , n49306 , n49307 , n49308 , n49309 , n49310 , n49311 , n49312 , n49313 , 
     n49314 , n49315 , n49316 , n49317 , n49318 , n49319 , n49320 , n49321 , n49322 , n49323 , 
     n49324 , n49325 , n49326 , n49327 , n49328 , n49329 , n49330 , n49331 , n49332 , n49333 , 
     n49334 , n49335 , n49336 , n49337 , n49338 , n49339 , n49340 , n49341 , n49342 , n49343 , 
     n49344 , n49345 , n49346 , n49347 , n49348 , n49349 , n49350 , n49351 , n49352 , n49353 , 
     n49354 , n49355 , n49356 , n49357 , n49358 , n49359 , n49360 , n49361 , n49362 , n49363 , 
     n49364 , n49365 , n49366 , n49367 , n49368 , n49369 , n49370 , n49371 , n49372 , n49373 , 
     n49374 , n49375 , n49376 , n49377 , n49378 , n49379 , n49380 , n49381 , n49382 , n49383 , 
     n49384 , n49385 , n49386 , n49387 , n49388 , n49389 , n49390 , n49391 , n49392 , n49393 , 
     n49394 , n49395 , n49396 , n49397 , n49398 , n49399 , n49400 , n49401 , n49402 , n49403 , 
     n49404 , n49405 , n49406 , n49407 , n49408 , n49409 , n49410 , n49411 , n49412 , n49413 , 
     n49414 , n49415 , n49416 , n49417 , n49418 , n49419 , n49420 , n49421 , n49422 , n49423 , 
     n49424 , n49425 , n49426 , n49427 , n49428 , n49429 , n49430 , n49431 , n49432 , n49433 , 
     n49434 , n49435 , n49436 , n49437 , n49438 , n49439 , n49440 , n49441 , n49442 , n49443 , 
     n49444 , n49445 , n49446 , n49447 , n49448 , n49449 , n49450 , n49451 , n49452 , n49453 , 
     n49454 , n49455 , n49456 , n49457 , n49458 , n49459 , n49460 , n49461 , n49462 , n49463 , 
     n49464 , n49465 , n49466 , n49467 , n49468 , n49469 , n49470 , n49471 , n49472 , n49473 , 
     n49474 , n49475 , n49476 , n49477 , n49478 , n49479 , n49480 , n49481 , n49482 , n49483 , 
     n49484 , n49485 , n49486 , n49487 , n49488 , n49489 , n49490 , n49491 , n49492 , n49493 , 
     n49494 , n49495 , n49496 , n49497 , n49498 , n49499 , n49500 , n49501 , n49502 , n49503 , 
     n49504 , n49505 , n49506 , n49507 , n49508 , n49509 , n49510 , n49511 , n49512 , n49513 , 
     n49514 , n49515 , n49516 , n49517 , n49518 , n49519 , n49520 , n49521 , n49522 , n49523 , 
     n49524 , n49525 , n49526 , n49527 , n49528 , n49529 , n49530 , n49531 , n49532 , n49533 , 
     n49534 , n49535 , n49536 , n49537 , n49538 , n49539 , n49540 , n49541 , n49542 , n49543 , 
     n49544 , n49545 , n49546 , n49547 , n49548 , n49549 , n49550 , n49551 , n49552 , n49553 , 
     n49554 , n49555 , n49556 , n49557 , n49558 , n49559 , n49560 , n49561 , n49562 , n49563 , 
     n49564 , n49565 , n49566 , n49567 , n49568 , n49569 , n49570 , n49571 , n49572 , n49573 , 
     n49574 , n49575 , n49576 , n49577 , n49578 , n49579 , n49580 , n49581 , n49582 , n49583 , 
     n49584 , n49585 , n49586 , n49587 , n49588 , n49589 , n49590 , n49591 , n49592 , n49593 , 
     n49594 , n49595 , n49596 , n49597 , n49598 , n49599 , n49600 , n49601 , n49602 , n49603 , 
     n49604 , n49605 , n49606 , n49607 , n49608 , n49609 , n49610 , n49611 , n49612 , n49613 , 
     n49614 , n49615 , n49616 , n49617 , n49618 , n49619 , n49620 , n49621 , n49622 , n49623 , 
     n49624 , n49625 , n49626 , n49627 , n49628 , n49629 , n49630 , n49631 , n49632 , n49633 , 
     n49634 , n49635 , n49636 , n49637 , n49638 , n49639 , n49640 , n49641 , n49642 , n49643 , 
     n49644 , n49645 , n49646 , n49647 , n49648 , n49649 , n49650 , n49651 , n49652 , n49653 , 
     n49654 , n49655 , n49656 , n49657 , n49658 , n49659 , n49660 , n49661 , n49662 , n49663 , 
     n49664 , n49665 , n49666 , n49667 , n49668 , n49669 , n49670 , n49671 , n49672 , n49673 , 
     n49674 , n49675 , n49676 , n49677 , n49678 , n49679 , n49680 , n49681 , n49682 , n49683 , 
     n49684 , n49685 , n49686 , n49687 , n49688 , n49689 , n49690 , n49691 , n49692 , n49693 , 
     n49694 , n49695 , n49696 , n49697 , n49698 , n49699 , n49700 , n49701 , n49702 , n49703 , 
     n49704 , n49705 , n49706 , n49707 , n49708 , n49709 , n49710 , n49711 , n49712 , n49713 , 
     n49714 , n49715 , n49716 , n49717 , n49718 , n49719 , n49720 , n49721 , n49722 , n49723 , 
     n49724 , n49725 , n49726 , n49727 , n49728 , n49729 , n49730 , n49731 , n49732 , n49733 , 
     n49734 , n49735 , n49736 , n49737 , n49738 , n49739 , n49740 , n49741 , n49742 , n49743 , 
     n49744 , n49745 , n49746 , n49747 , n49748 , n49749 , n49750 , n49751 , n49752 , n49753 , 
     n49754 , n49755 , n49756 , n49757 , n49758 , n49759 , n49760 , n49761 , n49762 , n49763 , 
     n49764 , n49765 , n49766 , n49767 , n49768 , n49769 , n49770 , n49771 , n49772 , n49773 , 
     n49774 , n49775 , n49776 , n49777 , n49778 , n49779 , n49780 , n49781 , n49782 , n49783 , 
     n49784 , n49785 , n49786 , n49787 , n49788 , n49789 , n49790 , n49791 , n49792 , n49793 , 
     n49794 , n49795 , n49796 , n49797 , n49798 , n49799 , n49800 , n49801 , n49802 , n49803 , 
     n49804 , n49805 , n49806 , n49807 , n49808 , n49809 , n49810 , n49811 , n49812 , n49813 , 
     n49814 , n49815 , n49816 , n49817 , n49818 , n49819 , n49820 , n49821 , n49822 , n49823 , 
     n49824 , n49825 , n49826 , n49827 , n49828 , n49829 , n49830 , n49831 , n49832 , n49833 , 
     n49834 , n49835 , n49836 , n49837 , n49838 , n49839 , n49840 , n49841 , n49842 , n49843 , 
     n49844 , n49845 , n49846 , n49847 , n49848 , n49849 , n49850 , n49851 , n49852 , n49853 , 
     n49854 , n49855 , n49856 , n49857 , n49858 , n49859 , n49860 , n49861 , n49862 , n49863 , 
     n49864 , n49865 , n49866 , n49867 , n49868 , n49869 , n49870 , n49871 , n49872 , n49873 , 
     n49874 , n49875 , n49876 , n49877 , n49878 , n49879 , n49880 , n49881 , n49882 , n49883 , 
     n49884 , n49885 , n49886 , n49887 , n49888 , n49889 , n49890 , n49891 , n49892 , n49893 , 
     n49894 , n49895 , n49896 , n49897 , n49898 , n49899 , n49900 , n49901 , n49902 , n49903 , 
     n49904 , n49905 , n49906 , n49907 , n49908 , n49909 , n49910 , n49911 , n49912 , n49913 , 
     n49914 , n49915 , n49916 , n49917 , n49918 , n49919 , n49920 , n49921 , n49922 , n49923 , 
     n49924 , n49925 , n49926 , n49927 , n49928 , n49929 , n49930 , n49931 , n49932 , n49933 , 
     n49934 , n49935 , n49936 , n49937 , n49938 , n49939 , n49940 , n49941 , n49942 , n49943 , 
     n49944 , n49945 , n49946 , n49947 , n49948 , n49949 , n49950 , n49951 , n49952 , n49953 , 
     n49954 , n49955 , n49956 , n49957 , n49958 , n49959 , n49960 , n49961 , n49962 , n49963 , 
     n49964 , n49965 , n49966 , n49967 , n49968 , n49969 , n49970 , n49971 , n49972 , n49973 , 
     n49974 , n49975 , n49976 , n49977 , n49978 , n49979 , n49980 , n49981 , n49982 , n49983 , 
     n49984 , n49985 , n49986 , n49987 , n49988 , n49989 , n49990 , n49991 , n49992 , n49993 , 
     n49994 , n49995 , n49996 , n49997 , n49998 , n49999 , n50000 , n50001 , n50002 , n50003 , 
     n50004 , n50005 , n50006 , n50007 , n50008 , n50009 , n50010 , n50011 , n50012 , n50013 , 
     n50014 , n50015 , n50016 , n50017 , n50018 , n50019 , n50020 , n50021 , n50022 , n50023 , 
     n50024 , n50025 , n50026 , n50027 , n50028 , n50029 , n50030 , n50031 , n50032 , n50033 , 
     n50034 , n50035 , n50036 , n50037 , n50038 , n50039 , n50040 , n50041 , n50042 , n50043 , 
     n50044 , n50045 , n50046 , n50047 , n50048 , n50049 , n50050 , n50051 , n50052 , n50053 , 
     n50054 , n50055 , n50056 , n50057 , n50058 , n50059 , n50060 , n50061 , n50062 , n50063 , 
     n50064 , n50065 , n50066 , n50067 , n50068 , n50069 , n50070 , n50071 , n50072 , n50073 , 
     n50074 , n50075 , n50076 , n50077 , n50078 , n50079 , n50080 , n50081 , n50082 , n50083 , 
     n50084 , n50085 , n50086 , n50087 , n50088 , n50089 , n50090 , n50091 , n50092 , n50093 , 
     n50094 , n50095 , n50096 , n50097 , n50098 , n50099 , n50100 , n50101 , n50102 , n50103 , 
     n50104 , n50105 , n50106 , n50107 , n50108 , n50109 , n50110 , n50111 , n50112 , n50113 , 
     n50114 , n50115 , n50116 , n50117 , n50118 , n50119 , n50120 , n50121 , n50122 , n50123 , 
     n50124 , n50125 , n50126 , n50127 , n50128 , n50129 , n50130 , n50131 , n50132 , n50133 , 
     n50134 , n50135 , n50136 , n50137 , n50138 , n50139 , n50140 , n50141 , n50142 , n50143 , 
     n50144 , n50145 , n50146 , n50147 , n50148 , n50149 , n50150 , n50151 , n50152 , n50153 , 
     n50154 , n50155 , n50156 , n50157 , n50158 , n50159 , n50160 , n50161 , n50162 , n50163 , 
     n50164 , n50165 , n50166 , n50167 , n50168 , n50169 , n50170 , n50171 , n50172 , n50173 , 
     n50174 , n50175 , n50176 , n50177 , n50178 , n50179 , n50180 , n50181 , n50182 , n50183 , 
     n50184 , n50185 , n50186 , n50187 , n50188 , n50189 , n50190 , n50191 , n50192 , n50193 , 
     n50194 , n50195 , n50196 , n50197 , n50198 , n50199 , n50200 , n50201 , n50202 , n50203 , 
     n50204 , n50205 , n50206 , n50207 , n50208 , n50209 , n50210 , n50211 , n50212 , n50213 , 
     n50214 , n50215 , n50216 , n50217 , n50218 , n50219 , n50220 , n50221 , n50222 , n50223 , 
     n50224 , n50225 , n50226 , n50227 , n50228 , n50229 , n50230 , n50231 , n50232 , n50233 , 
     n50234 , n50235 , n50236 , n50237 , n50238 , n50239 , n50240 , n50241 , n50242 , n50243 , 
     n50244 , n50245 , n50246 , n50247 , n50248 , n50249 , n50250 , n50251 , n50252 , n50253 , 
     n50254 , n50255 , n50256 , n50257 , n50258 , n50259 , n50260 , n50261 , n50262 , n50263 , 
     n50264 , n50265 , n50266 , n50267 , n50268 , n50269 , n50270 , n50271 , n50272 , n50273 , 
     n50274 , n50275 , n50276 , n50277 , n50278 , n50279 , n50280 , n50281 , n50282 , n50283 , 
     n50284 , n50285 , n50286 , n50287 , n50288 , n50289 , n50290 , n50291 , n50292 , n50293 , 
     n50294 , n50295 , n50296 , n50297 , n50298 , n50299 , n50300 , n50301 , n50302 , n50303 , 
     n50304 , n50305 , n50306 , n50307 , n50308 , n50309 , n50310 , n50311 , n50312 , n50313 , 
     n50314 , n50315 , n50316 , n50317 , n50318 , n50319 , n50320 , n50321 , n50322 , n50323 , 
     n50324 , n50325 , n50326 , n50327 , n50328 , n50329 , n50330 , n50331 , n50332 , n50333 , 
     n50334 , n50335 , n50336 , n50337 , n50338 , n50339 , n50340 , n50341 , n50342 , n50343 , 
     n50344 , n50345 , n50346 , n50347 , n50348 , n50349 , n50350 , n50351 , n50352 , n50353 , 
     n50354 , n50355 , n50356 , n50357 , n50358 , n50359 , n50360 , n50361 , n50362 , n50363 , 
     n50364 , n50365 , n50366 , n50367 , n50368 , n50369 , n50370 , n50371 , n50372 , n50373 , 
     n50374 , n50375 , n50376 , n50377 , n50378 , n50379 , n50380 , n50381 , n50382 , n50383 , 
     n50384 , n50385 , n50386 , n50387 , n50388 , n50389 , n50390 , n50391 , n50392 , n50393 , 
     n50394 , n50395 , n50396 , n50397 , n50398 , n50399 , n50400 , n50401 , n50402 , n50403 , 
     n50404 , n50405 , n50406 , n50407 , n50408 , n50409 , n50410 , n50411 , n50412 , n50413 , 
     n50414 , n50415 , n50416 , n50417 , n50418 , n50419 , n50420 , n50421 , n50422 , n50423 , 
     n50424 , n50425 , n50426 , n50427 , n50428 , n50429 , n50430 , n50431 , n50432 , n50433 , 
     n50434 , n50435 , n50436 , n50437 , n50438 , n50439 , n50440 , n50441 , n50442 , n50443 , 
     n50444 , n50445 , n50446 , n50447 , n50448 , n50449 , n50450 , n50451 , n50452 , n50453 , 
     n50454 , n50455 , n50456 , n50457 , n50458 , n50459 , n50460 , n50461 , n50462 , n50463 , 
     n50464 , n50465 , n50466 , n50467 , n50468 , n50469 , n50470 , n50471 , n50472 , n50473 , 
     n50474 , n50475 , n50476 , n50477 , n50478 , n50479 , n50480 , n50481 , n50482 , n50483 , 
     n50484 , n50485 , n50486 , n50487 , n50488 , n50489 , n50490 , n50491 , n50492 , n50493 , 
     n50494 , n50495 , n50496 , n50497 , n50498 , n50499 , n50500 , n50501 , n50502 , n50503 , 
     n50504 , n50505 , n50506 , n50507 , n50508 , n50509 , n50510 , n50511 , n50512 , n50513 , 
     n50514 , n50515 , n50516 , n50517 , n50518 , n50519 , n50520 , n50521 , n50522 , n50523 , 
     n50524 , n50525 , n50526 , n50527 , n50528 , n50529 , n50530 , n50531 , n50532 , n50533 , 
     n50534 , n50535 , n50536 , n50537 , n50538 , n50539 , n50540 , n50541 , n50542 , n50543 , 
     n50544 , n50545 , n50546 , n50547 , n50548 , n50549 , n50550 ;
buf ( RI21a19c60_2 , n0 );
buf ( RI21a5daf0_1 , n1 );
buf ( RI2107e620_463 , n2 );
buf ( RI210bf4e0_288 , n15 );
buf ( RI21078b30_503 , n48 );
buf ( RI21a13090_74 , n14 );
buf ( RI210bf558_287 , n17 );
buf ( RI21078ba8_502 , n49 );
buf ( RI21a13108_73 , n16 );
buf ( RI21a116c8_87 , n26 );
buf ( RI210bd6e0_301 , n27 );
buf ( RI21077078_516 , n54 );
buf ( RI21a11dd0_86 , n28 );
buf ( RI210bd758_300 , n29 );
buf ( RI210770f0_515 , n55 );
buf ( RI21a11e48_85 , n30 );
buf ( RI210bd7d0_299 , n31 );
buf ( RI21077168_514 , n56 );
buf ( RI21a132e8_69 , n24 );
buf ( RI210bff30_283 , n25 );
buf ( RI210797d8_498 , n53 );
buf ( RI210bfeb8_284 , n23 );
buf ( RI21079760_499 , n52 );
buf ( RI21a13270_70 , n22 );
buf ( RI210be1a8_295 , n39 );
buf ( RI21077d98_510 , n60 );
buf ( RI21a12028_81 , n38 );
buf ( RI21a12730_80 , n40 );
buf ( RI210bea18_294 , n41 );
buf ( RI21077e10_509 , n61 );
buf ( RI21a127a8_79 , n42 );
buf ( RI210bea90_293 , n43 );
buf ( RI21077e88_508 , n62 );
buf ( RI21079850_497 , n5 );
buf ( RI21a139f0_68 , n3 );
buf ( RI21084368_418 , n4 );
buf ( RI21a11f38_83 , n34 );
buf ( RI210be0b8_297 , n35 );
buf ( RI21077258_512 , n58 );
buf ( RI21a11fb0_82 , n36 );
buf ( RI210be130_296 , n37 );
buf ( RI21077d20_511 , n59 );
buf ( RI210be040_298 , n33 );
buf ( RI210771e0_513 , n57 );
buf ( RI21a11ec0_84 , n32 );
buf ( RI21a13180_72 , n18 );
buf ( RI210bfdc8_286 , n19 );
buf ( RI21078c20_501 , n50 );
buf ( RI21a131f8_71 , n20 );
buf ( RI210bfe40_285 , n21 );
buf ( RI21078c98_500 , n51 );
buf ( RI2107a660_489 , n63 );
buf ( RI2107cd48_472 , n78 );
buf ( RI2106bde0_608 , n94 );
buf ( RI2107c118_476 , n93 );
buf ( RI2107a570_491 , n90 );
buf ( RI21079940_495 , n86 );
buf ( RI2107a5e8_490 , n91 );
buf ( RI2107d900_469 , n81 );
buf ( RI2107b1a0_487 , n92 );
buf ( RI2107d978_468 , n82 );
buf ( RI2107a480_493 , n88 );
buf ( RI2107da68_466 , n84 );
buf ( RI210799b8_494 , n87 );
buf ( RI2107d9f0_467 , n83 );
buf ( RI2107a4f8_492 , n89 );
buf ( RI210798c8_496 , n85 );
buf ( RI2107ce38_470 , n80 );
buf ( RI2107cdc0_471 , n79 );
buf ( RI2107ccd0_473 , n77 );
buf ( RI2107cc58_474 , n76 );
buf ( RI2107c028_478 , n73 );
buf ( RI2107cbe0_475 , n75 );
buf ( RI2107c0a0_477 , n74 );
buf ( RI2107bfb0_479 , n72 );
buf ( RI2107b3f8_482 , n69 );
buf ( RI2107bf38_480 , n71 );
buf ( RI2107bec0_481 , n70 );
buf ( RI2107b380_483 , n68 );
buf ( RI2107b308_484 , n67 );
buf ( RI2107b218_486 , n65 );
buf ( RI2107b290_485 , n66 );
buf ( RI2107a6d8_488 , n64 );
buf ( RI2106be58_607 , n320 );
buf ( RI2107dae0_465 , n215 );
buf ( RI2106ddc0_566 , n217 );
buf ( RI210730b8_542 , n218 );
buf ( RI2106cc68_590 , n216 );
buf ( RI2106a2b0_640 , n102 );
buf ( RI21069ab8_644 , n117 );
buf ( RI2106bfc0_604 , n119 );
buf ( RI2106c038_603 , n120 );
buf ( RI2106a148_643 , n121 );
buf ( RI2106bf48_605 , n118 );
buf ( RI21069a40_645 , n115 );
buf ( RI2106a760_630 , n112 );
buf ( RI2106a5f8_633 , n109 );
buf ( RI2106a670_632 , n110 );
buf ( RI2106bed0_606 , n116 );
buf ( RI2106a7d8_629 , n113 );
buf ( RI2106c308_597 , n108 );
buf ( RI2106ae68_628 , n114 );
buf ( RI2106a6e8_631 , n111 );
buf ( RI2106a580_634 , n107 );
buf ( RI2106a508_635 , n106 );
buf ( RI2106a490_636 , n105 );
buf ( RI2106a3a0_638 , n104 );
buf ( RI2106a328_639 , n103 );
buf ( RI2106a238_641 , n101 );
buf ( RI2106c290_598 , n100 );
buf ( RI2106c218_599 , n99 );
buf ( RI2106c1a0_600 , n98 );
buf ( RI2106c128_601 , n97 );
buf ( RI2106c0b0_602 , n96 );
buf ( RI2106dd48_567 , n126 );
buf ( RI21073040_543 , n127 );
buf ( RI2106cbf0_591 , n125 );
buf ( RI21a12820_78 , n6 );
buf ( RI210beb08_292 , n7 );
buf ( RI21a0e608_121 , n219 );
buf ( RI21077f00_507 , n44 );
buf ( RI210b87a8_334 , n220 );
buf ( RI21a11560_90 , n284 );
buf ( RI210bcd80_304 , n285 );
buf ( RI210cfcc8_237 , n282 );
buf ( RI210842f0_419 , n283 );
buf ( RI21a0efe0_114 , n278 );
buf ( RI210b92e8_327 , n279 );
buf ( RI21a0f148_111 , n280 );
buf ( RI21084278_420 , n281 );
buf ( RI21a0ef68_115 , n276 );
buf ( RI210b9270_328 , n277 );
buf ( RI21a0eef0_116 , n274 );
buf ( RI210b91f8_329 , n275 );
buf ( RI21a0e680_120 , n266 );
buf ( RI210b8820_333 , n267 );
buf ( RI21a0e6f8_119 , n268 );
buf ( RI210b8898_332 , n269 );
buf ( RI21a10c00_96 , n254 );
buf ( RI210bc2b8_310 , n255 );
buf ( RI21a11470_92 , n262 );
buf ( RI210bcc90_306 , n263 );
buf ( RI21a10cf0_94 , n258 );
buf ( RI210bc3a8_308 , n259 );
buf ( RI21a0e770_118 , n270 );
buf ( RI210b8910_331 , n271 );
buf ( RI21a10c78_95 , n256 );
buf ( RI210bc330_309 , n257 );
buf ( RI21a114e8_91 , n264 );
buf ( RI210bcd08_305 , n265 );
buf ( RI21a10d68_93 , n260 );
buf ( RI210bc420_307 , n261 );
buf ( RI21a0e7e8_117 , n272 );
buf ( RI210b9180_330 , n273 );
buf ( RI21a102a0_102 , n242 );
buf ( RI210baff8_316 , n243 );
buf ( RI21a10318_101 , n244 );
buf ( RI210bb070_315 , n245 );
buf ( RI21a101b0_104 , n238 );
buf ( RI210baf08_318 , n239 );
buf ( RI21a10228_103 , n240 );
buf ( RI210baf80_317 , n241 );
buf ( RI21a10390_100 , n246 );
buf ( RI210bb8e0_314 , n247 );
buf ( RI21a10408_99 , n248 );
buf ( RI210bb958_313 , n249 );
buf ( RI21a10b10_98 , n250 );
buf ( RI210bb9d0_312 , n251 );
buf ( RI21a10b88_97 , n252 );
buf ( RI210bba48_311 , n253 );
buf ( RI21a0f940_108 , n230 );
buf ( RI210ba530_322 , n231 );
buf ( RI21a0f9b8_107 , n232 );
buf ( RI210ba5a8_321 , n233 );
buf ( RI21a0fa30_106 , n234 );
buf ( RI210ba620_320 , n235 );
buf ( RI21a0faa8_105 , n236 );
buf ( RI210ba698_319 , n237 );
buf ( RI21a0f850_110 , n226 );
buf ( RI210b9c48_324 , n227 );
buf ( RI21a0f8c8_109 , n228 );
buf ( RI210b9cc0_323 , n229 );
buf ( RI21a0f0d0_112 , n224 );
buf ( RI210b9bd0_325 , n225 );
buf ( RI21a19990_4 , n286 );
buf ( RI2106cd58_588 , n128 );
buf ( RI2106deb0_564 , n129 );
buf ( RI21073c70_539 , n130 );
buf ( RI21a198a0_6 , n291 );
buf ( RI2106de38_565 , n288 );
buf ( RI21073bf8_540 , n289 );
buf ( RI2106cce0_589 , n287 );
buf ( RI21a19918_5 , n290 );
buf ( RI21a0f058_113 , n222 );
buf ( RI210b9b58_326 , n223 );
buf ( RI21a19a08_3 , n221 );
buf ( RI21a197b0_8 , n293 );
buf ( RI2106ce48_586 , n134 );
buf ( RI21073d60_537 , n136 );
buf ( RI2106dfa0_562 , n135 );
buf ( RI2106df28_563 , n132 );
buf ( RI2106cdd0_587 , n131 );
buf ( RI21073ce8_538 , n133 );
buf ( RI21a19828_7 , n292 );
buf ( RI2106cec0_585 , n137 );
buf ( RI21073dd8_536 , n139 );
buf ( RI2106e018_561 , n138 );
buf ( RI21a190a8_9 , n294 );
buf ( RI210748a0_535 , n142 );
buf ( RI2106e090_560 , n141 );
buf ( RI2106cf38_584 , n140 );
buf ( RI21a19030_10 , n295 );
buf ( RI2106cfb0_583 , n143 );
buf ( RI21074918_534 , n145 );
buf ( RI2106e108_559 , n144 );
buf ( RI21a18fb8_11 , n296 );
buf ( RI21074990_533 , n148 );
buf ( RI21070a48_558 , n147 );
buf ( RI2106d028_582 , n146 );
buf ( RI21a18f40_12 , n297 );
buf ( RI21a18e50_14 , n299 );
buf ( RI2106d118_580 , n152 );
buf ( RI21074a80_531 , n154 );
buf ( RI21071588_556 , n153 );
buf ( RI21070ac0_557 , n150 );
buf ( RI2106d0a0_581 , n149 );
buf ( RI21074a08_532 , n151 );
buf ( RI21a18ec8_13 , n298 );
buf ( RI21a186d0_16 , n301 );
buf ( RI2106b1b0_621 , n158 );
buf ( RI21075638_528 , n160 );
buf ( RI2106b570_613 , n159 );
buf ( RI2106b4f8_614 , n156 );
buf ( RI2106b138_622 , n155 );
buf ( RI210755c0_529 , n157 );
buf ( RI21a18748_15 , n300 );
buf ( RI2106bc00_612 , n162 );
buf ( RI210756b0_527 , n163 );
buf ( RI2106b228_620 , n161 );
buf ( RI21a18658_17 , n302 );
buf ( RI2106d190_579 , n164 );
buf ( RI21075728_526 , n166 );
buf ( RI21071600_555 , n165 );
buf ( RI21a185e0_18 , n303 );
buf ( RI21a17410_28 , n313 );
buf ( RI21072e60_547 , n196 );
buf ( RI2106af58_626 , n194 );
buf ( RI2106dcd0_568 , n195 );
buf ( RI2106dc58_569 , n192 );
buf ( RI21072398_548 , n193 );
buf ( RI2106aee0_627 , n191 );
buf ( RI21a17488_27 , n312 );
buf ( RI21a17320_30 , n315 );
buf ( RI21072f50_545 , n202 );
buf ( RI2106afd0_625 , n200 );
buf ( RI2106b318_618 , n201 );
buf ( RI2106cb00_593 , n197 );
buf ( RI2106b2a0_619 , n198 );
buf ( RI21072ed8_546 , n199 );
buf ( RI21a17398_29 , n314 );
buf ( RI21a16b28_33 , n318 );
buf ( RI2106b0c0_623 , n209 );
buf ( RI2106b480_615 , n210 );
buf ( RI21074af8_530 , n211 );
buf ( RI2106a418_637 , n123 );
buf ( RI21072230_551 , n213 );
buf ( RI210764c0_519 , n214 );
buf ( RI2106c380_596 , n124 );
buf ( RI2106daf0_572 , n212 );
buf ( RI21a16ab0_34 , n319 );
buf ( RI2106cb78_592 , n203 );
buf ( RI21072fc8_544 , n205 );
buf ( RI2106b390_617 , n204 );
buf ( RI21a172a8_31 , n316 );
buf ( RI2106b048_624 , n206 );
buf ( RI2106b408_616 , n207 );
buf ( RI21073b80_541 , n208 );
buf ( RI2106a1c0_642 , n122 );
buf ( RI21a17230_32 , n317 );
buf ( RI21a184f0_20 , n305 );
buf ( RI2106d898_577 , n170 );
buf ( RI2106bc78_611 , n171 );
buf ( RI21075818_524 , n172 );
buf ( RI210757a0_525 , n169 );
buf ( RI2106d208_578 , n167 );
buf ( RI21071678_554 , n168 );
buf ( RI21a18568_19 , n304 );
buf ( RI21a17d70_22 , n307 );
buf ( RI210716f0_553 , n177 );
buf ( RI2106d988_575 , n176 );
buf ( RI21076358_522 , n178 );
buf ( RI2106d910_576 , n173 );
buf ( RI2106bcf0_610 , n174 );
buf ( RI210762e0_523 , n175 );
buf ( RI21a17de8_21 , n306 );
buf ( RI210721b8_552 , n180 );
buf ( RI2106da00_574 , n179 );
buf ( RI210763d0_521 , n181 );
buf ( RI21a17cf8_23 , n308 );
buf ( RI2106da78_573 , n182 );
buf ( RI21076448_520 , n184 );
buf ( RI2106bd68_609 , n183 );
buf ( RI21a17c80_24 , n309 );
buf ( RI21a17b90_26 , n311 );
buf ( RI2106ca88_594 , n188 );
buf ( RI21072320_549 , n190 );
buf ( RI2106dbe0_570 , n189 );
buf ( RI2106ca10_595 , n185 );
buf ( RI210722a8_550 , n187 );
buf ( RI2106db68_571 , n186 );
buf ( RI21a17c08_25 , n310 );
buf ( RI21a14440_60 , n321 );
buf ( RI21a15f70_44 , n335 );
buf ( RI21a14350_62 , n348 );
buf ( RI21a13ae0_66 , n344 );
buf ( RI21a13b58_65 , n345 );
buf ( RI21a168d0_38 , n341 );
buf ( RI21a13bd0_64 , n346 );
buf ( RI21a16948_37 , n342 );
buf ( RI21a169c0_36 , n352 );
buf ( RI21a15778_47 , n351 );
buf ( RI21a15fe8_43 , n336 );
buf ( RI21a16150_40 , n339 );
buf ( RI21a143c8_61 , n349 );
buf ( RI21a161c8_39 , n340 );
buf ( RI21a14530_58 , n350 );
buf ( RI21a16060_42 , n337 );
buf ( RI21a160d8_41 , n338 );
buf ( RI21a13a68_67 , n343 );
buf ( RI21a13c48_63 , n347 );
buf ( RI21a15868_45 , n334 );
buf ( RI21a15688_49 , n331 );
buf ( RI21a15700_48 , n332 );
buf ( RI21a157f0_46 , n333 );
buf ( RI21a15610_50 , n330 );
buf ( RI21a14f08_51 , n329 );
buf ( RI21a14e90_52 , n328 );
buf ( RI21a14e18_53 , n327 );
buf ( RI21a14da0_54 , n326 );
buf ( RI21a14d28_55 , n325 );
buf ( RI21a145a8_57 , n323 );
buf ( RI21a14cb0_56 , n324 );
buf ( RI21a144b8_59 , n322 );
buf ( RI210d8710_180 , n420 );
buf ( RI21a0b6b0_152 , n421 );
buf ( RI210d41b0_209 , n366 );
buf ( RI21a0de10_124 , n422 );
buf ( RI210d8788_179 , n417 );
buf ( RI21a0b728_151 , n418 );
buf ( RI210d4228_208 , n365 );
buf ( RI21a0de88_123 , n419 );
buf ( RI210d37d8_213 , n370 );
buf ( RI210d7d38_184 , n432 );
buf ( RI21a0ae40_156 , n433 );
buf ( RI21a0dc30_128 , n434 );
buf ( RI21a0aeb8_155 , n430 );
buf ( RI210d7db0_183 , n429 );
buf ( RI210d3850_212 , n369 );
buf ( RI21a0dca8_127 , n431 );
buf ( RI210d5560_201 , n396 );
buf ( RI210d9b38_171 , n397 );
buf ( RI210d1078_229 , n358 );
buf ( RI21a0c100_144 , n398 );
buf ( RI210d9160_175 , n409 );
buf ( RI210d4b88_205 , n408 );
buf ( RI210d06a0_233 , n362 );
buf ( RI21a0b908_147 , n410 );
buf ( RI210d4c00_204 , n405 );
buf ( RI210d99d0_174 , n406 );
buf ( RI210d0718_232 , n361 );
buf ( RI21a0c010_146 , n407 );
buf ( RI210d42a0_207 , n414 );
buf ( RI210d9070_177 , n415 );
buf ( RI210cfdb8_235 , n364 );
buf ( RI21a0b818_149 , n416 );
buf ( RI210d4b10_206 , n411 );
buf ( RI210d90e8_176 , n412 );
buf ( RI210d0628_234 , n363 );
buf ( RI21a0b890_148 , n413 );
buf ( RI210d54e8_202 , n399 );
buf ( RI210d9ac0_172 , n400 );
buf ( RI210d1000_230 , n359 );
buf ( RI210cf2f0_241 , n401 );
buf ( RI210d4c78_203 , n402 );
buf ( RI210d9a48_173 , n403 );
buf ( RI210d0790_231 , n360 );
buf ( RI21a0c088_145 , n404 );
buf ( RI21a0af30_154 , n427 );
buf ( RI210d8620_182 , n426 );
buf ( RI210d38c8_211 , n368 );
buf ( RI21a0dd20_126 , n428 );
buf ( RI210d4138_210 , n367 );
buf ( RI210d8698_181 , n423 );
buf ( RI21a0dd98_125 , n425 );
buf ( RI21a0afa8_153 , n424 );
buf ( RI210d2ef0_215 , n372 );
buf ( RI210cea08_243 , n439 );
buf ( RI210d7cc0_185 , n438 );
buf ( RI210cfc50_238 , n440 );
buf ( RI210d3760_214 , n371 );
buf ( RI210cf278_242 , n436 );
buf ( RI210ce8a0_246 , n435 );
buf ( RI21a0d528_129 , n437 );
buf ( RI210d23b0_222 , n378 );
buf ( RI21a0a558_161 , n457 );
buf ( RI210d6a00_191 , n456 );
buf ( RI21a0d2d0_134 , n458 );
buf ( RI21a0a648_159 , n451 );
buf ( RI210d72e8_189 , n450 );
buf ( RI210d24a0_220 , n376 );
buf ( RI21a0d3c0_132 , n452 );
buf ( RI210ce030_247 , n441 );
buf ( RI21a0adc8_157 , n442 );
buf ( RI21a0d4b0_130 , n443 );
buf ( RI210d2e78_216 , n373 );
buf ( RI21a0a5d0_160 , n454 );
buf ( RI210d7270_190 , n453 );
buf ( RI21a0d348_133 , n455 );
buf ( RI210d2428_221 , n377 );
buf ( RI210ce990_244 , n445 );
buf ( RI210d7c48_186 , n444 );
buf ( RI210d2e00_217 , n374 );
buf ( RI210cf3e0_239 , n446 );
buf ( RI210d2518_219 , n375 );
buf ( RI210ce918_245 , n448 );
buf ( RI210d7360_188 , n447 );
buf ( RI210cf368_240 , n449 );
buf ( RI21a09e50_162 , n460 );
buf ( RI210d1b40_223 , n379 );
buf ( RI21a0cbc8_135 , n461 );
buf ( RI210d6988_192 , n459 );
buf ( RI21a09dd8_163 , n462 );
buf ( RI210d6910_193 , n353 );
buf ( RI21a0cb50_136 , n463 );
buf ( RI210d1ac8_224 , n380 );
buf ( RI21a09478_164 , n465 );
buf ( RI210d6898_194 , n464 );
buf ( RI210d1a50_225 , n381 );
buf ( RI21a0cad8_137 , n466 );
buf ( RI210d2d88_218 , n356 );
buf ( RI21a0d438_131 , n392 );
buf ( RI21a0a6c0_158 , n391 );
buf ( RI210d73d8_187 , n390 );
buf ( RI210d10f0_228 , n357 );
buf ( RI210d5ec0_198 , n393 );
buf ( RI210da498_168 , n394 );
buf ( RI21a0c268_141 , n395 );
buf ( RI210d5fb0_196 , n470 );
buf ( RI210dad80_166 , n471 );
buf ( RI210d1168_227 , n383 );
buf ( RI21a0c9e8_139 , n472 );
buf ( RI210d5f38_197 , n477 );
buf ( RI210da510_167 , n478 );
buf ( RI21a0c970_140 , n479 );
buf ( RI210da420_169 , n475 );
buf ( RI210d5650_199 , n474 );
buf ( RI21a0c1f0_142 , n476 );
buf ( RI210d6028_195 , n467 );
buf ( RI210dadf8_165 , n468 );
buf ( RI21a0ca60_138 , n469 );
buf ( RI210d19d8_226 , n382 );
buf ( RI210da3a8_170 , n388 );
buf ( RI210d55d8_200 , n387 );
buf ( RI21a0c178_143 , n389 );
buf ( RI210cdfb8_248 , n354 );
buf ( RI21a0e590_122 , n386 );
buf ( RI21a0b7a0_150 , n385 );
buf ( RI210d8ff8_178 , n384 );
buf ( RI210cfd40_236 , n482 );
buf ( RI21a16a38_35 , n473 );
buf ( RI21a115d8_89 , n481 );
buf ( RI21a11650_88 , n480 );
buf ( RI210ccb90_257 , n499 );
buf ( RI210c9b48_275 , n483 );
buf ( RI210cd658_251 , n514 );
buf ( RI210cc140_262 , n513 );
buf ( RI210ca430_273 , n512 );
buf ( RI210c9ad0_276 , n511 );
buf ( RI210c91e8_278 , n509 );
buf ( RI210c9a58_277 , n510 );
buf ( RI210c2078_280 , n507 );
buf ( RI210c9170_279 , n508 );
buf ( RI210c07a0_282 , n505 );
buf ( RI210c0818_281 , n506 );
buf ( RI210cd568_253 , n503 );
buf ( RI210cd5e0_252 , n504 );
buf ( RI210ccc80_255 , n501 );
buf ( RI210cd4f0_254 , n502 );
buf ( RI210ccc08_256 , n500 );
buf ( RI210cc2a8_259 , n497 );
buf ( RI210ccb18_258 , n498 );
buf ( RI210cc230_260 , n496 );
buf ( RI210cb8d0_263 , n494 );
buf ( RI210cb858_264 , n493 );
buf ( RI210cc1b8_261 , n495 );
buf ( RI210cb7e0_265 , n492 );
buf ( RI210cb768_266 , n491 );
buf ( RI210caef8_267 , n490 );
buf ( RI210cae80_268 , n489 );
buf ( RI210cae08_269 , n488 );
buf ( RI210cad90_270 , n487 );
buf ( RI210ca4a8_272 , n485 );
buf ( RI210ca520_271 , n486 );
buf ( RI210ca3b8_274 , n484 );
buf ( RI210aeb90_395 , n516 );
buf ( RI210b43b0_360 , n547 );
buf ( RI210b7f38_335 , n548 );
buf ( RI210b2538_374 , n546 );
buf ( RI210b5670_354 , n556 );
buf ( RI21081aa0_439 , n555 );
buf ( RI2107e878_458 , n519 );
buf ( RI210b07b0_386 , n554 );
buf ( RI210af478_393 , n572 );
buf ( RI21080d80_445 , n573 );
buf ( RI2107e698_462 , n525 );
buf ( RI210834e0_427 , n574 );
buf ( RI2107f3b8_456 , n560 );
buf ( RI21080f60_441 , n561 );
buf ( RI210835d0_425 , n562 );
buf ( RI21084458_416 , n521 );
buf ( RI210afdd8_390 , n563 );
buf ( RI21080ee8_442 , n564 );
buf ( RI2107e800_459 , n522 );
buf ( RI210b4d10_357 , n565 );
buf ( RI210aec08_394 , n575 );
buf ( RI210b25b0_373 , n576 );
buf ( RI210843e0_417 , n526 );
buf ( RI210b4428_359 , n577 );
buf ( RI210b08a0_384 , n632 );
buf ( RI210b2f88_369 , n633 );
buf ( RI210b5760_352 , n634 );
buf ( RI21084f98_414 , n545 );
buf ( RI210b2f10_370 , n640 );
buf ( RI210b0828_385 , n639 );
buf ( RI210b56e8_353 , n641 );
buf ( RI210b3078_367 , n627 );
buf ( RI210b1188_382 , n626 );
buf ( RI210b6048_350 , n628 );
buf ( RI21085088_412 , n543 );
buf ( RI210b3000_368 , n630 );
buf ( RI210b0918_383 , n629 );
buf ( RI21085010_413 , n544 );
buf ( RI210b57d8_351 , n631 );
buf ( RI21085c40_409 , n540 );
buf ( RI210b61b0_347 , n619 );
buf ( RI210b12f0_379 , n617 );
buf ( RI210b39d8_364 , n618 );
buf ( RI21085cb8_408 , n539 );
buf ( RI210b6a20_346 , n616 );
buf ( RI210b1b60_378 , n614 );
buf ( RI210b3a50_363 , n615 );
buf ( RI210b73f8_342 , n607 );
buf ( RI21085e20_405 , n536 );
buf ( RI2107f520_453 , n605 );
buf ( RI21081b90_437 , n606 );
buf ( RI210836c0_423 , n604 );
buf ( RI21085e98_404 , n535 );
buf ( RI21081c08_436 , n603 );
buf ( RI210b1c50_376 , n602 );
buf ( RI210b1200_381 , n623 );
buf ( RI210b38e8_366 , n624 );
buf ( RI210b60c0_349 , n625 );
buf ( RI21085100_411 , n542 );
buf ( RI210b6b10_344 , n610 );
buf ( RI21085da8_406 , n537 );
buf ( RI210b4338_361 , n609 );
buf ( RI2107f430_455 , n608 );
buf ( RI210b7470_341 , n595 );
buf ( RI21086a50_401 , n532 );
buf ( RI210800d8_450 , n593 );
buf ( RI210827c0_433 , n594 );
buf ( RI210b74e8_340 , n592 );
buf ( RI21086ac8_400 , n531 );
buf ( RI21082838_432 , n591 );
buf ( RI21080150_449 , n590 );
buf ( RI210802b8_446 , n581 );
buf ( RI210829a0_429 , n582 );
buf ( RI21086e10_397 , n528 );
buf ( RI210b7e48_337 , n583 );
buf ( RI210b1cc8_375 , n578 );
buf ( RI21082a18_428 , n579 );
buf ( RI210a63a0_396 , n527 );
buf ( RI210b7ec0_336 , n580 );
buf ( RI21085178_410 , n541 );
buf ( RI210b6138_348 , n622 );
buf ( RI210b1278_380 , n620 );
buf ( RI210b3960_365 , n621 );
buf ( RI210b6a98_345 , n613 );
buf ( RI21085d30_407 , n538 );
buf ( RI210b42c0_362 , n612 );
buf ( RI210b1bd8_377 , n611 );
buf ( RI210b26a0_371 , n637 );
buf ( RI210b4e00_355 , n638 );
buf ( RI210aff40_387 , n636 );
buf ( RI21083648_424 , n559 );
buf ( RI21084f20_415 , n520 );
buf ( RI210afe50_389 , n557 );
buf ( RI21080fd8_440 , n558 );
buf ( RI210af4f0_392 , n569 );
buf ( RI21080df8_444 , n570 );
buf ( RI2107e710_461 , n524 );
buf ( RI21083558_426 , n571 );
buf ( RI2107e788_460 , n523 );
buf ( RI210b4c98_358 , n568 );
buf ( RI210af568_391 , n566 );
buf ( RI21080e70_443 , n567 );
buf ( RI21083738_422 , n601 );
buf ( RI21086960_403 , n534 );
buf ( RI21081c80_435 , n600 );
buf ( RI2107f598_452 , n599 );
buf ( RI21084200_421 , n598 );
buf ( RI210869d8_402 , n533 );
buf ( RI21081cf8_434 , n597 );
buf ( RI21080060_451 , n596 );
buf ( RI210828b0_431 , n588 );
buf ( RI210801c8_448 , n587 );
buf ( RI21086b40_399 , n530 );
buf ( RI210b7560_339 , n589 );
buf ( RI21082928_430 , n585 );
buf ( RI21080240_447 , n584 );
buf ( RI210b7dd0_338 , n586 );
buf ( RI21086bb8_398 , n529 );
buf ( RI210b2628_372 , n550 );
buf ( RI210afec8_388 , n549 );
buf ( RI210b4d88_356 , n551 );
buf ( RI210b6b88_343 , n553 );
buf ( RI21081b18_438 , n552 );
buf ( RI2107f4a8_454 , n515 );
buf ( RI2107f340_457 , n518 );
buf ( RI210cdec8_250 , n635 );
buf ( RI210bcdf8_303 , n643 );
buf ( RI210bd668_302 , n642 );
buf ( RI21077000_517 , n644 );
buf ( RI21076538_518 , n645 );
buf ( RI21a12988_75 , n12 );
buf ( RI210bf468_289 , n13 );
buf ( RI21078ab8_504 , n47 );
buf ( RI21a12910_76 , n10 );
buf ( RI210bf3f0_290 , n11 );
buf ( RI21078a40_505 , n46 );
buf ( RI21a12898_77 , n8 );
buf ( RI210beb80_291 , n9 );
buf ( RI21077f78_506 , n45 );
buf ( RI210cdf40_249 , n646 );
buf ( RI2107db58_464 , n647 );
buf ( RI21069950_647 , n648 );
buf ( RI210699c8_646 , n649 );
buf ( n650 , R_61e_1dfaf3c8 );
buf ( n651 , R_8f7_1e09b6c8 );
buf ( n652 , R_714_1dfb8888 );
buf ( n653 , R_951_1e17ef68 );
buf ( n654 , R_28c_1d9fb268 );
buf ( n655 , R_9be_1e183888 );
buf ( n656 , R_9ab_1e1827a8 );
buf ( n657 , R_30f_1d9d04a8 );
buf ( n658 , R_959_1e17f468 );
buf ( n659 , R_b13_1e6b0908 );
buf ( n660 , R_519_1dda4b48 );
buf ( n661 , R_92d_1e09d888 );
buf ( n662 , R_c06_1e6bafe8 );
buf ( n663 , R_8c6_1e099d28 );
buf ( n664 , R_845_1e094788 );
buf ( n665 , R_414_1d9da7c8 );
buf ( n666 , R_313_1d9d0728 );
buf ( n667 , R_518_1dda4aa8 );
buf ( n668 , R_9d9_1e184468 );
buf ( n669 , R_4dd_1dda25c8 );
buf ( n670 , R_59f_1dda9f08 );
buf ( n671 , R_517_1dda4a08 );
buf ( n672 , R_509_1dda4148 );
buf ( n673 , R_508_1dda40a8 );
buf ( n674 , R_401_1d9d9be8 );
buf ( n675 , R_5f9_1ddad748 );
buf ( n676 , R_6ef_1dfb7168 );
buf ( n677 , R_a30_1e187ac8 );
buf ( n678 , R_2b0_1d9fc8e8 );
buf ( n679 , R_77c_1dfbc988 );
buf ( n680 , R_8f1_1e09b308 );
buf ( n681 , R_36a_1d9d4288 );
buf ( n682 , R_507_1dda4008 );
buf ( n683 , R_516_1dda4e68 );
buf ( n684 , R_98e_1e181a88 );
buf ( n685 , R_8d5_1e09a188 );
buf ( n686 , R_498_1dd9faa8 );
buf ( n687 , R_68b_1dfb32e8 );
buf ( n688 , R_773_1dfbc3e8 );
buf ( n689 , R_45b_1d9dd428 );
buf ( n690 , R_48d_1dd9f3c8 );
buf ( n691 , R_5ff_1ddadb08 );
buf ( n692 , R_705_1dfb7f28 );
buf ( n693 , R_644_1dfb0688 );
buf ( n694 , R_63a_1dfb0548 );
buf ( n695 , R_ac7_1e18d928 );
buf ( n696 , R_320_1d9d0f48 );
buf ( n697 , R_737_1dfb9e68 );
buf ( n698 , R_506_1dda4468 );
buf ( n699 , R_647_1dfb0868 );
buf ( n700 , R_b86_1e6bb4e8 );
buf ( n701 , R_883_1e096e48 );
buf ( n702 , R_6a8_1dfb4508 );
buf ( n703 , R_aa5_1e18c3e8 );
buf ( n704 , R_440_1d9dc348 );
buf ( n705 , R_2f9_1d9cf6e8 );
buf ( n706 , R_69c_1dfb3d88 );
buf ( n707 , R_65d_1dfb1628 );
buf ( n708 , R_b0c_1e6b04a8 );
buf ( n709 , R_b20_1e6b1128 );
buf ( n710 , R_a2e_1e189788 );
buf ( n711 , R_905_1e09bf88 );
buf ( n712 , R_a57_1e189328 );
buf ( n713 , R_5f8_1ddad6a8 );
buf ( n714 , R_54c_1dda6b28 );
buf ( n715 , R_bd2_1e6b32e8 );
buf ( n716 , R_aca_1e6ae068 );
buf ( n717 , R_58b_1dda9288 );
buf ( n718 , R_2e3_1d9ce928 );
buf ( n719 , R_3e2_1d9d8d88 );
buf ( n720 , R_8f6_1e09bb28 );
buf ( n721 , R_331_1d9d19e8 );
buf ( n722 , R_97d_1e180ae8 );
buf ( n723 , R_5cd_1ddabbc8 );
buf ( n724 , R_45c_1d9dd4c8 );
buf ( n725 , R_999_1e181c68 );
buf ( n726 , R_b99_1e6b5cc8 );
buf ( n727 , R_948_1e17e9c8 );
buf ( n728 , R_97e_1e181308 );
buf ( n729 , R_ab0_1e18cac8 );
buf ( n730 , R_bb8_1e6b7028 );
buf ( n731 , R_489_1dd9f148 );
buf ( n732 , R_4b6_1dda1268 );
buf ( n733 , R_63f_1dfb0368 );
buf ( n734 , R_3e7_1d9d8ba8 );
buf ( n735 , R_2bd_1d9fd108 );
buf ( n736 , R_81b_1e092d48 );
buf ( n737 , R_b54_1e6b31a8 );
buf ( n738 , R_4df_1dda2708 );
buf ( n739 , R_bab_1e6b6808 );
buf ( n740 , R_431_1d9db9e8 );
buf ( n741 , R_2f2_1d9cf788 );
buf ( n742 , R_601_1ddadc48 );
buf ( n743 , R_6e7_1dfb6c68 );
buf ( n744 , R_bdf_1e6b8888 );
buf ( n745 , R_656_1dfb1bc8 );
buf ( n746 , R_4e0_1dda27a8 );
buf ( n747 , R_4de_1dda2b68 );
buf ( n748 , R_a4e_1e189288 );
buf ( n749 , R_8e1_1e09a908 );
buf ( n750 , R_8f0_1e09b268 );
buf ( n751 , R_299_1d9fba88 );
buf ( n752 , R_292_1d9fb628 );
buf ( n753 , R_4e1_1dda2848 );
buf ( n754 , R_a7f_1e18ac28 );
buf ( n755 , R_c04_1e6b9fa8 );
buf ( n756 , R_3ef_1d9d90a8 );
buf ( n757 , R_5de_1dd9f1e8 );
buf ( n758 , R_878_1e096768 );
buf ( n759 , R_720_1dfb9008 );
buf ( n760 , R_ad6_1e6ae7e8 );
buf ( n761 , R_9a2_1e182708 );
buf ( n762 , R_630_1dfafa08 );
buf ( n763 , R_52f_1dda5908 );
buf ( n764 , R_7a9_1e08e608 );
buf ( n765 , R_976_1e180b88 );
buf ( n766 , R_439_1d9dbee8 );
buf ( n767 , R_604_1ddade28 );
buf ( n768 , R_530_1dda59a8 );
buf ( n769 , R_52e_1dda5d68 );
buf ( n770 , R_7ed_1e091088 );
buf ( n771 , R_3f2_1d9d4c88 );
buf ( n772 , R_3d4_1d9d7fc8 );
buf ( n773 , R_84a_1e094fa8 );
buf ( n774 , R_2de_1d9ceb08 );
buf ( n775 , R_690_1dfb3608 );
buf ( n776 , R_4cd_1dda1bc8 );
buf ( n777 , R_531_1dda5a48 );
buf ( n778 , R_b34_1e6b1da8 );
buf ( n779 , R_5f7_1ddad608 );
buf ( n780 , R_806_1e092528 );
buf ( n781 , R_a5b_1e1895a8 );
buf ( n782 , R_718_1dfb8b08 );
buf ( n783 , R_695_1dfb3928 );
buf ( n784 , R_7af_1e08e9c8 );
buf ( n785 , R_62b_1dfaf6e8 );
buf ( n786 , R_904_1e09bee8 );
buf ( n787 , R_501_1dda3c48 );
buf ( n788 , R_585_1dda8ec8 );
buf ( n789 , R_9cd_1e183ce8 );
buf ( n790 , R_78c_1dfbd388 );
buf ( n791 , R_392_1d9d5b88 );
buf ( n792 , R_4b4_1dda0c28 );
buf ( n793 , R_b44_1e6b27a8 );
buf ( n794 , R_969_1e17fe68 );
buf ( n795 , R_40d_1d9da368 );
buf ( n796 , R_627_1dfaf468 );
buf ( n797 , R_67a_1dfadfc8 );
buf ( n798 , R_45d_1d9dd568 );
buf ( n799 , R_7c1_1e08f508 );
buf ( n800 , R_552_1dda73e8 );
buf ( n801 , R_2bf_1d9fd248 );
buf ( n802 , R_5d4_1ddac028 );
buf ( n803 , R_b77_1e6b4788 );
buf ( n804 , R_3fa_1d9db088 );
buf ( n805 , R_6aa_1dfb4b48 );
buf ( n806 , R_82a_1e093ba8 );
buf ( n807 , R_3aa_1d9d6a88 );
buf ( n808 , R_300_1d9cfb48 );
buf ( n809 , R_405_1d9d9e68 );
buf ( n810 , R_953_1e17f0a8 );
buf ( n811 , R_3cf_1d9d7ca8 );
buf ( n812 , R_ac1_1e18d568 );
buf ( n813 , R_61c_1dfaed88 );
buf ( n814 , R_a99_1e18bc68 );
buf ( n815 , R_4ae_1dda0fe8 );
buf ( n816 , R_aec_1e6af0a8 );
buf ( n817 , R_af8_1e6af828 );
buf ( n818 , R_762_1dfbbe48 );
buf ( n819 , R_3a8_1d9d6448 );
buf ( n820 , R_4ca_1dda1ee8 );
buf ( n821 , R_6b7_1dfb4e68 );
buf ( n822 , R_57c_1dda8928 );
buf ( n823 , R_52b_1dda5688 );
buf ( n824 , R_8ef_1e09b1c8 );
buf ( n825 , R_8c5_1e099788 );
buf ( n826 , R_8ab_1e098748 );
buf ( n827 , R_71c_1dfb8d88 );
buf ( n828 , R_388_1d9d5048 );
buf ( n829 , R_b6e_1e6b46e8 );
buf ( n830 , R_9cc_1e183c48 );
buf ( n831 , R_65b_1dfb14e8 );
buf ( n832 , R_bbd_1e6b7348 );
buf ( n833 , R_3b2_1d9d6f88 );
buf ( n834 , R_862_1e095ea8 );
buf ( n835 , R_4a5_1dda02c8 );
buf ( n836 , R_90f_1e09c5c8 );
buf ( n837 , R_702_1dfb8248 );
buf ( n838 , R_29f_1d9fbe48 );
buf ( n839 , R_72b_1dfb96e8 );
buf ( n840 , R_6f4_1dfb7488 );
buf ( n841 , R_5f2_1dda8a68 );
buf ( n842 , R_a64_1e189b48 );
buf ( n843 , R_2e9_1d9cece8 );
buf ( n844 , R_683_1dfb2de8 );
buf ( n845 , R_2fd_1d9cf968 );
buf ( n846 , R_8b2_1e0990a8 );
buf ( n847 , R_5f0_1ddad1a8 );
buf ( n848 , R_bac_1e6b68a8 );
buf ( n849 , R_642_1dfb0a48 );
buf ( n850 , R_5f6_1d9fbda8 );
buf ( n851 , R_568_1dda7ca8 );
buf ( n852 , R_409_1d9da0e8 );
buf ( n853 , R_5a8_1ddaa4a8 );
buf ( n854 , R_5e3_1ddac988 );
buf ( n855 , R_96b_1e17ffa8 );
buf ( n856 , R_bca_1e6b14e8 );
buf ( n857 , R_3b8_1d9d6e48 );
buf ( n858 , R_789_1dfbd1a8 );
buf ( n859 , R_86a_1e0963a8 );
buf ( n860 , R_416_1ddabc68 );
buf ( n861 , R_903_1e09be48 );
buf ( n862 , R_a2d_1e1878e8 );
buf ( n863 , R_9cb_1e183ba8 );
buf ( n864 , R_59b_1dda9c88 );
buf ( n865 , R_a4c_1e188c48 );
buf ( n866 , R_79c_1dfbdd88 );
buf ( n867 , R_888_1e097168 );
buf ( n868 , R_2a7_1d9fc348 );
buf ( n869 , R_7f3_1e091448 );
buf ( n870 , R_73c_1dfba188 );
buf ( n871 , R_bd1_1e6b7fc8 );
buf ( n872 , R_4a6_1dda0868 );
buf ( n873 , R_3dd_1d9d8568 );
buf ( n874 , R_346_1d9d2c08 );
buf ( n875 , R_4c4_1dda1628 );
buf ( n876 , R_b15_1e6b0a48 );
buf ( n877 , R_5ec_1ddacf28 );
buf ( n878 , R_bb4_1e6b6da8 );
buf ( n879 , R_bed_1e6b9148 );
buf ( n880 , R_7bf_1e08f3c8 );
buf ( n881 , R_344_1d9d25c8 );
buf ( n882 , R_c0b_1e6ba408 );
buf ( n883 , R_6a5_1dfb4328 );
buf ( n884 , R_b8c_1e6b54a8 );
buf ( n885 , R_3a1_1d9d5fe8 );
buf ( n886 , R_7ea_1e09d928 );
buf ( n887 , R_46e_1dd9e568 );
buf ( n888 , R_8ee_1e09b628 );
buf ( n889 , R_697_1dfb3a68 );
buf ( n890 , R_77f_1dfbcb68 );
buf ( n891 , R_391_1d9d55e8 );
buf ( n892 , R_746_1dfb6448 );
buf ( n893 , R_b3b_1e6b2208 );
buf ( n894 , R_7f1_1e091308 );
buf ( n895 , R_410_1d9da548 );
buf ( n896 , R_700_1dfb7c08 );
buf ( n897 , R_58f_1dda9508 );
buf ( n898 , R_582_1dda91e8 );
buf ( n899 , R_793_1dfbd7e8 );
buf ( n900 , R_847_1e0948c8 );
buf ( n901 , R_95e_1e17fc88 );
buf ( n902 , R_560_1dda77a8 );
buf ( n903 , R_9ca_1e184008 );
buf ( n904 , R_397_1d9d59a8 );
buf ( n905 , R_46b_1d9dde28 );
buf ( n906 , R_44e_1d9fc028 );
buf ( n907 , R_6cc_1dfb5b88 );
buf ( n908 , R_62e_1dfafdc8 );
buf ( n909 , R_2b1_1d9fc988 );
buf ( n910 , R_6f9_1dfb77a8 );
buf ( n911 , R_af5_1e6af648 );
buf ( n912 , R_b81_1e6b4dc8 );
buf ( n913 , R_427_1d9db3a8 );
buf ( n914 , R_547_1dda6808 );
buf ( n915 , R_c1d_1e6baf48 );
buf ( n916 , R_a2c_1e187848 );
buf ( n917 , R_355_1d9d3068 );
buf ( n918 , R_857_1e0952c8 );
buf ( n919 , R_413_1d9da728 );
buf ( n920 , R_afa_1e6afe68 );
buf ( n921 , R_adc_1e6ae6a8 );
buf ( n922 , R_5fc_1ddad928 );
buf ( n923 , R_c24_1e6bb3a8 );
buf ( n924 , R_421_1d9dafe8 );
buf ( n925 , R_892_1e17e608 );
buf ( n926 , R_70b_1dfb82e8 );
buf ( n927 , R_aad_1e18c8e8 );
buf ( n928 , R_3ca_1d9d8108 );
buf ( n929 , R_7ac_1e08e7e8 );
buf ( n930 , R_8da_1e09a9a8 );
buf ( n931 , R_400_1d9d9b48 );
buf ( n932 , R_bb0_1e6b6b28 );
buf ( n933 , R_893_1e097848 );
buf ( n934 , R_902_1e09c2a8 );
buf ( n935 , R_a93_1e18b8a8 );
buf ( n936 , R_8cd_1e099c88 );
buf ( n937 , R_861_1e095908 );
buf ( n938 , R_3ea_1d9d9288 );
buf ( n939 , R_915_1e09c988 );
buf ( n940 , R_844_1e0946e8 );
buf ( n941 , R_677_1dfb2668 );
buf ( n942 , R_602_1dfae248 );
buf ( n943 , R_39c_1d9d5cc8 );
buf ( n944 , R_be3_1e6b8b08 );
buf ( n945 , R_bea_1e6b9468 );
buf ( n946 , R_993_1e1818a8 );
buf ( n947 , R_bad_1e6b6948 );
buf ( n948 , R_88d_1e097488 );
buf ( n949 , R_5a2_1ddaa5e8 );
buf ( n950 , R_655_1dfb1128 );
buf ( n951 , R_4ad_1dda07c8 );
buf ( n952 , R_493_1dd9f788 );
buf ( n953 , R_894_1e0978e8 );
buf ( n954 , R_668_1dfb1d08 );
buf ( n955 , R_730_1dfb9a08 );
buf ( n956 , R_7dc_1e0905e8 );
buf ( n957 , R_abd_1e18d2e8 );
buf ( n958 , R_662_1dfb1e48 );
buf ( n959 , R_a7c_1e18aa48 );
buf ( n960 , R_5cf_1ddabd08 );
buf ( n961 , R_328_1d9d1448 );
buf ( n962 , R_741_1dfba4a8 );
buf ( n963 , R_9a6_1e182988 );
buf ( n964 , R_36d_1d9d3f68 );
buf ( n965 , R_308_1d9d0048 );
buf ( n966 , R_95b_1e17f5a8 );
buf ( n967 , R_b63_1e6b3b08 );
buf ( n968 , R_2da_1d9ce888 );
buf ( n969 , R_5dc_1ddac528 );
buf ( n970 , R_49f_1dd9ff08 );
buf ( n971 , R_895_1e097988 );
buf ( n972 , R_761_1dfbb8a8 );
buf ( n973 , R_2e4_1d9ce9c8 );
buf ( n974 , R_ab5_1e18cde8 );
buf ( n975 , R_c28_1e6bb628 );
buf ( n976 , R_8d4_1e09a0e8 );
buf ( n977 , R_a8c_1e18b448 );
buf ( n978 , R_597_1dda9a08 );
buf ( n979 , R_5c4_1ddab628 );
buf ( n980 , R_384_1d9d4dc8 );
buf ( n981 , R_31c_1d9d0cc8 );
buf ( n982 , R_987_1e181128 );
buf ( n983 , R_b2e_1e6b1ee8 );
buf ( n984 , R_2f3_1d9cf328 );
buf ( n985 , R_6cf_1dfb5d68 );
buf ( n986 , R_6e4_1dfb6a88 );
buf ( n987 , R_357_1d9d31a8 );
buf ( n988 , R_3c1_1d9d73e8 );
buf ( n989 , R_5e7_1ddacc08 );
buf ( n990 , R_974_1e180548 );
buf ( n991 , R_61a_1dfaf148 );
buf ( n992 , R_3f8_1d9d9648 );
buf ( n993 , R_802_1e0922a8 );
buf ( n994 , R_593_1dda9788 );
buf ( n995 , R_a69_1e189e68 );
buf ( n996 , R_a87_1e18b128 );
buf ( n997 , R_a5d_1e1896e8 );
buf ( n998 , R_a2b_1e1877a8 );
buf ( n999 , R_671_1dfb22a8 );
buf ( n1000 , R_4cf_1dda1d08 );
buf ( n1001 , R_420_1d9daf48 );
buf ( n1002 , R_6bc_1dfb5188 );
buf ( n1003 , R_43f_1d9dc2a8 );
buf ( n1004 , R_692_1dfb3c48 );
buf ( n1005 , R_80b_1e092348 );
buf ( n1006 , R_882_1e0972a8 );
buf ( n1007 , R_871_1e096308 );
buf ( n1008 , R_2c2_1d9fd928 );
buf ( n1009 , R_2ce_1d9cfa08 );
buf ( n1010 , R_a9c_1e18be48 );
buf ( n1011 , R_768_1dfbbd08 );
buf ( n1012 , R_56d_1dda7fc8 );
buf ( n1013 , R_34c_1d9d2ac8 );
buf ( n1014 , R_b8f_1e6b5688 );
buf ( n1015 , R_b07_1e6b0188 );
buf ( n1016 , R_6b5_1dfb4d28 );
buf ( n1017 , R_5ae_1ddaad68 );
buf ( n1018 , R_2df_1d9ce6a8 );
buf ( n1019 , R_674_1dfb2488 );
buf ( n1020 , R_608_1dfae108 );
buf ( n1021 , R_ad3_1e6ae108 );
buf ( n1022 , R_505_1dda3ec8 );
buf ( n1023 , R_8bf_1e0993c8 );
buf ( n1024 , R_542_1dda69e8 );
buf ( n1025 , R_7f6_1e091b28 );
buf ( n1026 , R_504_1dda3e28 );
buf ( n1027 , R_8a7_1e0984c8 );
buf ( n1028 , R_76a_1dfbc5c8 );
buf ( n1029 , R_937_1e09dec8 );
buf ( n1030 , R_6fb_1dfb78e8 );
buf ( n1031 , R_3b0_1d9d6948 );
buf ( n1032 , R_2c0_1d9fd2e8 );
buf ( n1033 , R_37c_1d9d48c8 );
buf ( n1034 , R_782_1dfbd248 );
buf ( n1035 , R_503_1dda3d88 );
buf ( n1036 , R_82e_1e093e28 );
buf ( n1037 , R_8bb_1e099148 );
buf ( n1038 , R_430_1d9db948 );
buf ( n1039 , R_5cb_1ddaba88 );
buf ( n1040 , R_ae6_1e6af1e8 );
buf ( n1041 , R_7a3_1e08e248 );
buf ( n1042 , R_b78_1e6b4828 );
buf ( n1043 , R_bc9_1e6b7ac8 );
buf ( n1044 , R_380_1d9d4b48 );
buf ( n1045 , R_33d_1d9d2168 );
buf ( n1046 , R_8e0_1e09a868 );
buf ( n1047 , R_3c7_1d9d77a8 );
buf ( n1048 , R_2b2_1d9fcf28 );
buf ( n1049 , R_618_1dfaeb08 );
buf ( n1050 , R_823_1e093248 );
buf ( n1051 , R_89e_1e098428 );
buf ( n1052 , R_502_1dda41e8 );
buf ( n1053 , R_b6f_1e6b4288 );
buf ( n1054 , R_c00_1e6b9d28 );
buf ( n1055 , R_98d_1e1814e8 );
buf ( n1056 , R_28b_1d9fb1c8 );
buf ( n1057 , R_a55_1e1891e8 );
buf ( n1058 , R_3c4_1d9d75c8 );
buf ( n1059 , R_40c_1d9da2c8 );
buf ( n1060 , R_2d2_1d9ce388 );
buf ( n1061 , R_c21_1e6bb1c8 );
buf ( n1062 , R_b3d_1e6b2348 );
buf ( n1063 , R_877_1e0966c8 );
buf ( n1064 , R_855_1e095188 );
buf ( n1065 , R_41d_1d9dad68 );
buf ( n1066 , R_438_1d9dbe48 );
buf ( n1067 , R_2d6_1d9ce608 );
buf ( n1068 , R_7da_1e0909a8 );
buf ( n1069 , R_6f6_1dfb7ac8 );
buf ( n1070 , R_9aa_1e182e88 );
buf ( n1071 , R_b47_1e6b2988 );
buf ( n1072 , R_a2a_1e6b3ce8 );
buf ( n1073 , R_41f_1d9daea8 );
buf ( n1074 , R_ae4_1e6aeba8 );
buf ( n1075 , R_a79_1e18a868 );
buf ( n1076 , R_3a3_1d9d6128 );
buf ( n1077 , R_5bd_1ddab1c8 );
buf ( n1078 , R_301_1d9cfbe8 );
buf ( n1079 , R_298_1d9fb9e8 );
buf ( n1080 , R_bb9_1e6b70c8 );
buf ( n1081 , R_82d_1e093888 );
buf ( n1082 , R_404_1d9d9dc8 );
buf ( n1083 , R_a62_1e189f08 );
buf ( n1084 , R_93c_1e17e248 );
buf ( n1085 , R_62d_1dfaf828 );
buf ( n1086 , R_579_1dda8748 );
buf ( n1087 , R_452_1ddac3e8 );
buf ( n1088 , R_54d_1dda6bc8 );
buf ( n1089 , R_4d9_1dda2348 );
buf ( n1090 , R_4d4_1dda2028 );
buf ( n1091 , R_6c1_1dfb54a8 );
buf ( n1092 , R_379_1d9d46e8 );
buf ( n1093 , R_34e_1d9d3108 );
buf ( n1094 , R_94a_1e097ca8 );
buf ( n1095 , R_74b_1dfbaae8 );
buf ( n1096 , R_ade_1e6aece8 );
buf ( n1097 , R_79f_1e08dfc8 );
buf ( n1098 , R_797_1dfbda68 );
buf ( n1099 , R_943_1e17e6a8 );
buf ( n1100 , R_653_1dfb0fe8 );
buf ( n1101 , R_3d8_1d9d8248 );
buf ( n1102 , R_b61_1e6b39c8 );
buf ( n1103 , R_bc4_1e6b77a8 );
buf ( n1104 , R_a02_1e186308 );
buf ( n1105 , R_368_1d9d3c48 );
buf ( n1106 , R_35e_1d9d3b08 );
buf ( n1107 , R_7fe_1e092028 );
buf ( n1108 , R_499_1dd9fb48 );
buf ( n1109 , R_680_1dfb2c08 );
buf ( n1110 , R_2a8_1d9fc3e8 );
buf ( n1111 , R_6ec_1dfb6f88 );
buf ( n1112 , R_776_1dfbcac8 );
buf ( n1113 , R_b5e_1e6b0368 );
buf ( n1114 , R_635_1dfafd28 );
buf ( n1115 , R_7fa_1e091da8 );
buf ( n1116 , R_af7_1e6af788 );
buf ( n1117 , R_8c4_1e0996e8 );
buf ( n1118 , R_408_1d9da048 );
buf ( n1119 , R_ab9_1e18d068 );
buf ( n1120 , R_6a2_1dfb61c8 );
buf ( n1121 , R_291_1d9fb588 );
buf ( n1122 , R_7b8_1e08ef68 );
buf ( n1123 , R_8b6_1e08e6a8 );
buf ( n1124 , R_48a_1dda0d68 );
buf ( n1125 , R_6c7_1dfb5868 );
buf ( n1126 , R_c10_1e6ba728 );
buf ( n1127 , R_bf1_1e6b93c8 );
buf ( n1128 , R_4d6_1dd9e2e8 );
buf ( n1129 , R_5b3_1ddaab88 );
buf ( n1130 , R_771_1dfbc2a8 );
buf ( n1131 , R_af1_1e6af3c8 );
buf ( n1132 , R_6e1_1dfb68a8 );
buf ( n1133 , R_a9f_1e18c028 );
buf ( n1134 , R_b17_1e6b0b88 );
buf ( n1135 , R_b30_1e6b1b28 );
buf ( n1136 , R_bde_1e6b37e8 );
buf ( n1137 , R_998_1e181bc8 );
buf ( n1138 , R_a4a_1e189008 );
buf ( n1139 , R_48e_1dd9f968 );
buf ( n1140 , R_688_1dfb3108 );
buf ( n1141 , R_810_1e092668 );
buf ( n1142 , R_75c_1dfbb588 );
buf ( n1143 , R_3bb_1d9d7028 );
buf ( n1144 , R_c2e_1e17f008 );
buf ( n1145 , R_5d2_1d9db308 );
buf ( n1146 , R_32e_1d9d1d08 );
buf ( n1147 , R_580_1dda8ba8 );
buf ( n1148 , R_453_1d9dcf28 );
buf ( n1149 , R_83a_1e0913a8 );
buf ( n1150 , R_41e_1d9dc988 );
buf ( n1151 , R_97c_1e180a48 );
buf ( n1152 , R_5b8_1ddaaea8 );
buf ( n1153 , R_363_1d9d3928 );
buf ( n1154 , R_94e_1ddadce8 );
buf ( n1155 , R_7c4_1e08f6e8 );
buf ( n1156 , R_52c_1dda5728 );
buf ( n1157 , R_aa2_1e18c708 );
buf ( n1158 , R_625_1dfaf328 );
buf ( n1159 , R_4b7_1dda0e08 );
buf ( n1160 , R_55d_1dda75c8 );
buf ( n1161 , R_b0e_1e6b0ae8 );
buf ( n1162 , R_425_1d9db268 );
buf ( n1163 , R_30c_1d9d02c8 );
buf ( n1164 , R_3db_1d9d8428 );
buf ( n1165 , R_a48_1e1889c8 );
buf ( n1166 , R_aaf_1e18ca28 );
buf ( n1167 , R_5ad_1ddaa7c8 );
buf ( n1168 , R_589_1dda9148 );
buf ( n1169 , R_338_1d9d1e48 );
buf ( n1170 , R_832_1e0940a8 );
buf ( n1171 , R_790_1dfbd608 );
buf ( n1172 , R_318_1d9d0a48 );
buf ( n1173 , R_869_1e095e08 );
buf ( n1174 , R_6d3_1dfb5fe8 );
buf ( n1175 , R_60c_1dfae388 );
buf ( n1176 , R_56a_1dda82e8 );
buf ( n1177 , R_887_1e0970c8 );
buf ( n1178 , R_815_1e092988 );
buf ( n1179 , R_66b_1dfb1ee8 );
buf ( n1180 , R_a34_1e187d48 );
buf ( n1181 , R_40f_1d9da4a8 );
buf ( n1182 , R_ac3_1e18d6a8 );
buf ( n1183 , R_324_1d9d11c8 );
buf ( n1184 , R_614_1dfae888 );
buf ( n1185 , R_752_1dfbb448 );
buf ( n1186 , R_4c0_1dda13a8 );
buf ( n1187 , R_7d9_1e090408 );
buf ( n1188 , R_ad0_1e18dec8 );
buf ( n1189 , R_bee_1e6b96e8 );
buf ( n1190 , R_736_1dfba2c8 );
buf ( n1191 , R_727_1dfb9468 );
buf ( n1192 , R_a8a_1e18b808 );
buf ( n1193 , R_933_1e09dc48 );
buf ( n1194 , R_8b1_1e098b08 );
buf ( n1195 , R_606_1dfae4c8 );
buf ( n1196 , R_927_1e09d4c8 );
buf ( n1197 , R_a7a_1e18ae08 );
buf ( n1198 , R_333_1d9d1b28 );
buf ( n1199 , R_968_1e17fdc8 );
buf ( n1200 , R_574_1dda8428 );
buf ( n1201 , R_836_1e094328 );
buf ( n1202 , R_757_1dfbb268 );
buf ( n1203 , R_2db_1d9ce428 );
buf ( n1204 , R_af4_1e6af5a8 );
buf ( n1205 , R_454_1d9dcfc8 );
buf ( n1206 , R_412_1d9dab88 );
buf ( n1207 , R_709_1dfb81a8 );
buf ( n1208 , R_8a4_1e0982e8 );
buf ( n1209 , R_c1b_1e6bae08 );
buf ( n1210 , R_846_1e094d28 );
buf ( n1211 , R_3ff_1d9d9aa8 );
buf ( n1212 , R_76e_1dfbdec8 );
buf ( n1213 , R_33f_1d9d22a8 );
buf ( n1214 , R_4af_1dda0908 );
buf ( n1215 , R_a67_1e189d28 );
buf ( n1216 , R_616_1dfaeec8 );
buf ( n1217 , R_b49_1e6b2ac8 );
buf ( n1218 , R_2f4_1d9cf3c8 );
buf ( n1219 , R_426_1d9db808 );
buf ( n1220 , R_2e5_1d9cea68 );
buf ( n1221 , R_bb5_1e6b6e48 );
buf ( n1222 , R_7b6_1e08f328 );
buf ( n1223 , R_751_1dfbaea8 );
buf ( n1224 , R_bd0_1e6b7f28 );
buf ( n1225 , R_610_1dfae608 );
buf ( n1226 , R_918_1e09cb68 );
buf ( n1227 , R_35c_1d9d34c8 );
buf ( n1228 , R_924_1e09d2e8 );
buf ( n1229 , R_912_1e09cca8 );
buf ( n1230 , R_77d_1dfbca28 );
buf ( n1231 , R_774_1dfbc488 );
buf ( n1232 , R_a71_1e18a368 );
buf ( n1233 , R_32d_1d9d1768 );
buf ( n1234 , R_99d_1e181ee8 );
buf ( n1235 , R_87d_1e096a88 );
buf ( n1236 , R_472_1dd9e7e8 );
buf ( n1237 , R_b2a_1e6b1c68 );
buf ( n1238 , R_56f_1dda8108 );
buf ( n1239 , R_b87_1e6b5188 );
buf ( n1240 , R_921_1e09d108 );
buf ( n1241 , R_375_1d9d4468 );
buf ( n1242 , R_576_1dda8ce8 );
buf ( n1243 , R_b82_1e6b5368 );
buf ( n1244 , R_39e_1d9d6308 );
buf ( n1245 , R_856_1e095728 );
buf ( n1246 , R_6c2_1dfb5a48 );
buf ( n1247 , R_2c3_1d9fd4c8 );
buf ( n1248 , R_90b_1e09c348 );
buf ( n1249 , R_92f_1e09d9c8 );
buf ( n1250 , R_38e_1d9d5908 );
buf ( n1251 , R_b9e_1e18d388 );
buf ( n1252 , R_8cc_1e099be8 );
buf ( n1253 , R_860_1e095868 );
buf ( n1254 , R_c09_1e6ba2c8 );
buf ( n1255 , R_b09_1e6b02c8 );
buf ( n1256 , R_521_1dda5048 );
buf ( n1257 , R_b4a_1e6b3068 );
buf ( n1258 , R_88c_1e0973e8 );
buf ( n1259 , R_520_1dda4fa8 );
buf ( n1260 , R_8b5_1e098d88 );
buf ( n1261 , R_b5d_1e6b3748 );
buf ( n1262 , R_843_1e094648 );
buf ( n1263 , R_633_1dfafbe8 );
buf ( n1264 , R_7c2_1e08faa8 );
buf ( n1265 , R_6d8_1dfb6308 );
buf ( n1266 , R_38d_1d9d5368 );
buf ( n1267 , R_7e7_1e090cc8 );
buf ( n1268 , R_bfc_1e6b9aa8 );
buf ( n1269 , R_841_1e094508 );
buf ( n1270 , R_a96_1e18bf88 );
buf ( n1271 , R_7e5_1e090b88 );
buf ( n1272 , R_51f_1dda4f08 );
buf ( n1273 , R_949_1e17ea68 );
buf ( n1274 , R_b5a_1e6b3a68 );
buf ( n1275 , R_2e0_1d9ce748 );
buf ( n1276 , R_acd_1e18dce8 );
buf ( n1277 , R_70f_1dfb8568 );
buf ( n1278 , R_c15_1e6baa48 );
buf ( n1279 , R_310_1d9d0548 );
buf ( n1280 , R_bf5_1e6b9648 );
buf ( n1281 , R_314_1d9d07c8 );
buf ( n1282 , R_6af_1dfb4968 );
buf ( n1283 , R_445_1d9dc668 );
buf ( n1284 , R_658_1dfb1308 );
buf ( n1285 , R_a6c_1e18a048 );
buf ( n1286 , R_2c1_1d9fd388 );
buf ( n1287 , R_2b3_1d9fcac8 );
buf ( n1288 , R_6de_1dfb6bc8 );
buf ( n1289 , R_9b9_1e183068 );
buf ( n1290 , R_6ad_1dfb4828 );
buf ( n1291 , R_548_1dda68a8 );
buf ( n1292 , R_4c9_1dda1948 );
buf ( n1293 , R_51e_1dda5368 );
buf ( n1294 , R_96a_1e180408 );
buf ( n1295 , R_455_1d9dd068 );
buf ( n1296 , R_8d3_1e09a048 );
buf ( n1297 , R_bb1_1e6b6bc8 );
buf ( n1298 , R_7d7_1e0902c8 );
buf ( n1299 , R_6a0_1dfb4008 );
buf ( n1300 , R_b79_1e6b48c8 );
buf ( n1301 , R_565_1dda7ac8 );
buf ( n1302 , R_586_1dda9468 );
buf ( n1303 , R_4a7_1dda0408 );
buf ( n1304 , R_b70_1e6b4328 );
buf ( n1305 , R_661_1dfb18a8 );
buf ( n1306 , R_2d3_1d9fdec8 );
buf ( n1307 , R_ad9_1e6ae4c8 );
buf ( n1308 , R_a85_1e18afe8 );
buf ( n1309 , R_a77_1e18a728 );
buf ( n1310 , R_2d7_1d9ce1a8 );
buf ( n1311 , R_7b3_1e08ec48 );
buf ( n1312 , R_870_1e096268 );
buf ( n1313 , R_43e_1d9dc708 );
buf ( n1314 , R_6db_1dfb64e8 );
buf ( n1315 , R_807_1e0920c8 );
buf ( n1316 , R_a74_1e18a548 );
buf ( n1317 , R_bf9_1e6b98c8 );
buf ( n1318 , R_321_1d9d0fe8 );
buf ( n1319 , R_a53_1e1890a8 );
buf ( n1320 , R_4e3_1dda2988 );
buf ( n1321 , R_831_1e093b08 );
buf ( n1322 , R_66e_1dfb25c8 );
buf ( n1323 , R_ac6_1e18dd88 );
buf ( n1324 , R_55a_1dda78e8 );
buf ( n1325 , R_4c6_1dda1c68 );
buf ( n1326 , R_4e4_1dda2a28 );
buf ( n1327 , R_4e2_1dda2de8 );
buf ( n1328 , R_c22_1e6b55e8 );
buf ( n1329 , R_92c_1e09d7e8 );
buf ( n1330 , R_7c9_1e08fa08 );
buf ( n1331 , R_623_1dfaf1e8 );
buf ( n1332 , R_b58_1e6b3428 );
buf ( n1333 , R_370_1d9d4148 );
buf ( n1334 , R_3be_1d9d7708 );
buf ( n1335 , R_4e5_1dda2ac8 );
buf ( n1336 , R_a03_1e185ea8 );
buf ( n1337 , R_c12_1e6bad68 );
buf ( n1338 , R_456_1d9dd608 );
buf ( n1339 , R_bf2_1e6b9968 );
buf ( n1340 , R_6a7_1dfb4468 );
buf ( n1341 , R_c30_1e6bbb28 );
buf ( n1342 , R_40b_1d9da228 );
buf ( n1343 , R_42f_1d9db8a8 );
buf ( n1344 , R_68d_1dfb3428 );
buf ( n1345 , R_735_1dfb9d28 );
buf ( n1346 , R_78d_1dfbd428 );
buf ( n1347 , R_8df_1e09a7c8 );
buf ( n1348 , R_41c_1d9dacc8 );
buf ( n1349 , R_46f_1dd9e108 );
buf ( n1350 , R_2a9_1d9fc488 );
buf ( n1351 , R_81e_1e093428 );
buf ( n1352 , R_5e0_1ddac7a8 );
buf ( n1353 , R_462_1d9ddd88 );
buf ( n1354 , R_60a_1dfae748 );
buf ( n1355 , R_5a7_1ddaa408 );
buf ( n1356 , R_403_1d9d9d28 );
buf ( n1357 , R_2c6_1d9fdba8 );
buf ( n1358 , R_7e3_1e090a48 );
buf ( n1359 , R_7ee_1e09c528 );
buf ( n1360 , R_706_1dfb84c8 );
buf ( n1361 , R_c17_1e6bab88 );
buf ( n1362 , R_c1f_1e6bb088 );
buf ( n1363 , R_b93_1e6b5908 );
buf ( n1364 , R_854_1e0950e8 );
buf ( n1365 , R_b9f_1e6b6088 );
buf ( n1366 , R_8e5_1e09ab88 );
buf ( n1367 , R_437_1d9dbda8 );
buf ( n1368 , R_612_1dfaec48 );
buf ( n1369 , R_816_1e0931a8 );
buf ( n1370 , R_b19_1e6b0cc8 );
buf ( n1371 , R_73b_1dfba0e8 );
buf ( n1372 , R_a44_1e188748 );
buf ( n1373 , R_93e_1e17e888 );
buf ( n1374 , R_67c_1dfb2988 );
buf ( n1375 , R_992_1e181d08 );
buf ( n1376 , R_494_1dd9f828 );
buf ( n1377 , R_3e0_1d9d8748 );
buf ( n1378 , R_7a7_1e08e4c8 );
buf ( n1379 , R_876_1e096b28 );
buf ( n1380 , R_543_1dda6588 );
buf ( n1381 , R_8ae_1dfbc0c8 );
buf ( n1382 , R_351_1d9d2de8 );
buf ( n1383 , R_457_1d9dd1a8 );
buf ( n1384 , R_bf6_1e6b3f68 );
buf ( n1385 , R_a38_1e187fc8 );
buf ( n1386 , R_6f1_1dfb72a8 );
buf ( n1387 , R_b3e_1e6b28e8 );
buf ( n1388 , R_53e_1dda6768 );
buf ( n1389 , R_ac0_1e18d4c8 );
buf ( n1390 , R_763_1dfbb9e8 );
buf ( n1391 , R_c26_1e6b8ce8 );
buf ( n1392 , R_650_1dfb0e08 );
buf ( n1393 , R_361_1d9d37e8 );
buf ( n1394 , R_aaa_1e187e88 );
buf ( n1395 , R_b10_1e6b0728 );
buf ( n1396 , R_b2c_1e6b18a8 );
buf ( n1397 , R_5a1_1ddaa048 );
buf ( n1398 , R_be7_1e6b8d88 );
buf ( n1399 , R_b26_1e6b19e8 );
buf ( n1400 , R_4a0_1dd9ffa8 );
buf ( n1401 , R_95a_1e17fa08 );
buf ( n1402 , R_909_1e09c208 );
buf ( n1403 , R_463_1d9dd928 );
buf ( n1404 , R_407_1d9d9fa8 );
buf ( n1405 , R_5c5_1ddab6c8 );
buf ( n1406 , R_986_1e181588 );
buf ( n1407 , R_515_1dda48c8 );
buf ( n1408 , R_5c1_1ddab448 );
buf ( n1409 , R_297_1d9fb948 );
buf ( n1410 , R_514_1dda4828 );
buf ( n1411 , R_b4c_1e6b2ca8 );
buf ( n1412 , R_973_1e1804a8 );
buf ( n1413 , R_60e_1dfae9c8 );
buf ( n1414 , R_7d4_1e0900e8 );
buf ( n1415 , R_7c7_1e08f8c8 );
buf ( n1416 , R_513_1dda4788 );
buf ( n1417 , R_65f_1dfb1768 );
buf ( n1418 , R_9b5_1e182de8 );
buf ( n1419 , R_2ee_1d9cf508 );
buf ( n1420 , R_91b_1e09cd48 );
buf ( n1421 , R_af6_1e6afbe8 );
buf ( n1422 , R_83d_1e094288 );
buf ( n1423 , R_8c3_1e099648 );
buf ( n1424 , R_458_1d9dd248 );
buf ( n1425 , R_512_1dda4be8 );
buf ( n1426 , R_ba6_1e6b69e8 );
buf ( n1427 , R_5e5_1ddacac8 );
buf ( n1428 , R_57b_1dda8888 );
buf ( n1429 , R_aeb_1e6af008 );
buf ( n1430 , R_7f4_1e0914e8 );
buf ( n1431 , R_a46_1e188d88 );
buf ( n1432 , R_b8d_1e6b5548 );
buf ( n1433 , R_562_1dda7de8 );
buf ( n1434 , R_745_1dfba728 );
buf ( n1435 , R_557_1dda7208 );
buf ( n1436 , R_464_1d9dd9c8 );
buf ( n1437 , R_835_1e093d88 );
buf ( n1438 , R_49a_1dda00e8 );
buf ( n1439 , R_7d1_1e08ff08 );
buf ( n1440 , R_911_1e09c708 );
buf ( n1441 , R_6e9_1dfb6da8 );
buf ( n1442 , R_723_1dfb91e8 );
buf ( n1443 , R_a95_1e18b9e8 );
buf ( n1444 , R_58d_1dda93c8 );
buf ( n1445 , R_a89_1e18b268 );
buf ( n1446 , R_780_1dfbcc08 );
buf ( n1447 , R_740_1dfba408 );
buf ( n1448 , R_72f_1dfb9968 );
buf ( n1449 , R_828_1e093568 );
buf ( n1450 , R_89c_1e097de8 );
buf ( n1451 , R_a32_1e188108 );
buf ( n1452 , R_840_1e094468 );
buf ( n1453 , R_b37_1e6b1f88 );
buf ( n1454 , R_9db_1e1845a8 );
buf ( n1455 , R_b22_1e6b1768 );
buf ( n1456 , R_9dc_1e184648 );
buf ( n1457 , R_9da_1e184a08 );
buf ( n1458 , R_794_1dfbd888 );
buf ( n1459 , R_33a_1d9d2488 );
buf ( n1460 , R_424_1d9db1c8 );
buf ( n1461 , R_2dc_1d9ce4c8 );
buf ( n1462 , R_a6f_1e18a228 );
buf ( n1463 , R_98c_1e181448 );
buf ( n1464 , R_6b6_1dfb52c8 );
buf ( n1465 , R_908_1e09c168 );
buf ( n1466 , R_9dd_1e1846e8 );
buf ( n1467 , R_965_1e17fbe8 );
buf ( n1468 , R_28a_1d9fb128 );
buf ( n1469 , R_529_1dda5548 );
buf ( n1470 , R_40e_1d9da908 );
buf ( n1471 , R_bcd_1e6b7d48 );
buf ( n1472 , R_476_1dd9ea68 );
buf ( n1473 , R_393_1d9d5728 );
buf ( n1474 , R_a40_1e1884c8 );
buf ( n1475 , R_528_1dda54a8 );
buf ( n1476 , R_2fa_1d9d0188 );
buf ( n1477 , R_a3c_1e188248 );
buf ( n1478 , R_868_1e095d68 );
buf ( n1479 , R_2cf_1d9fdc48 );
buf ( n1480 , R_2c4_1d9fd568 );
buf ( n1481 , R_7cc_1e08fbe8 );
buf ( n1482 , R_8fd_1e09ba88 );
buf ( n1483 , R_3d5_1d9d8068 );
buf ( n1484 , R_b64_1e6b3ba8 );
buf ( n1485 , R_527_1dda5408 );
buf ( n1486 , R_9d1_1e183f68 );
buf ( n1487 , R_46c_1d9ddec8 );
buf ( n1488 , R_2f5_1d9cf468 );
buf ( n1489 , R_839_1e094008 );
buf ( n1490 , R_554_1dda7028 );
buf ( n1491 , R_3ab_1d9d6628 );
buf ( n1492 , R_459_1d9dd2e8 );
buf ( n1493 , R_b4f_1e6b2e88 );
buf ( n1494 , R_886_1e097528 );
buf ( n1495 , R_3e5_1d9d8a68 );
buf ( n1496 , R_52d_1dda57c8 );
buf ( n1497 , R_290_1d9fb4e8 );
buf ( n1498 , R_b7a_1e18cc08 );
buf ( n1499 , R_526_1dda5ae8 );
buf ( n1500 , R_79a_1e098e28 );
buf ( n1501 , R_ba0_1e6b6128 );
buf ( n1502 , R_6d1_1dfb5ea8 );
buf ( n1503 , R_713_1dfb87e8 );
buf ( n1504 , R_685_1dfb2f28 );
buf ( n1505 , R_3fe_1d9d9f08 );
buf ( n1506 , R_638_1dfaff08 );
buf ( n1507 , R_465_1d9dda68 );
buf ( n1508 , R_b91_1e6b57c8 );
buf ( n1509 , R_b53_1e6b3108 );
buf ( n1510 , R_8ad_1e098888 );
buf ( n1511 , R_59e_1dd9e068 );
buf ( n1512 , R_9c5_1e1837e8 );
buf ( n1513 , R_3a9_1d9d64e8 );
buf ( n1514 , R_3b3_1d9d6b28 );
buf ( n1515 , R_2b4_1d9fcb68 );
buf ( n1516 , R_af3_1e6af508 );
buf ( n1517 , R_4f9_1dda3748 );
buf ( n1518 , R_a90_1e18b6c8 );
buf ( n1519 , R_389_1d9d50e8 );
buf ( n1520 , R_a6a_1e18a408 );
buf ( n1521 , R_b1b_1e6b0e08 );
buf ( n1522 , R_4f8_1dda36a8 );
buf ( n1523 , R_b66_1e6b9be8 );
buf ( n1524 , R_9d0_1e183ec8 );
buf ( n1525 , R_2e1_1d9ce7e8 );
buf ( n1526 , R_7d2_1e0904a8 );
buf ( n1527 , R_803_1e091e48 );
buf ( n1528 , R_91e_1e09d428 );
buf ( n1529 , R_4f7_1dda3608 );
buf ( n1530 , R_ab4_1e18cd48 );
buf ( n1531 , R_6ee_1dfb75c8 );
buf ( n1532 , R_c05_1e6ba048 );
buf ( n1533 , R_704_1dfb7e88 );
buf ( n1534 , R_353_1d9d2f28 );
buf ( n1535 , R_ba7_1e6b6588 );
buf ( n1536 , R_87c_1e0969e8 );
buf ( n1537 , R_3f5_1d9d9468 );
buf ( n1538 , R_abc_1e18d248 );
buf ( n1539 , R_a83_1e18aea8 );
buf ( n1540 , R_b40_1e6b2528 );
buf ( n1541 , R_a06_1e186588 );
buf ( n1542 , R_907_1e09c0c8 );
buf ( n1543 , R_664_1dfb1a88 );
buf ( n1544 , R_b71_1e6b43c8 );
buf ( n1545 , R_4f6_1ddad2e8 );
buf ( n1546 , R_8b9_1e099008 );
buf ( n1547 , R_971_1e180368 );
buf ( n1548 , R_64e_1dfb11c8 );
buf ( n1549 , R_679_1dfb27a8 );
buf ( n1550 , R_80c_1e0923e8 );
buf ( n1551 , R_347_1d9d27a8 );
buf ( n1552 , R_b28_1e6b1628 );
buf ( n1553 , R_7cf_1e08fdc8 );
buf ( n1554 , R_8fc_1e09b9e8 );
buf ( n1555 , R_72d_1dfb9828 );
buf ( n1556 , R_9c4_1e183748 );
buf ( n1557 , R_997_1e181b28 );
buf ( n1558 , R_85f_1e0957c8 );
buf ( n1559 , R_2d4_1d9cdfc8 );
buf ( n1560 , R_48f_1dd9f508 );
buf ( n1561 , R_adb_1e6ae608 );
buf ( n1562 , R_3b9_1d9d6ee8 );
buf ( n1563 , R_a51_1e188f68 );
buf ( n1564 , R_8cb_1e099b48 );
buf ( n1565 , R_2d8_1d9ce248 );
buf ( n1566 , R_a72_1e18a908 );
buf ( n1567 , R_7f7_1e0916c8 );
buf ( n1568 , R_4b5_1dda0cc8 );
buf ( n1569 , R_88b_1e097348 );
buf ( n1570 , R_aa7_1e18c528 );
buf ( n1571 , R_699_1dfb3ba8 );
buf ( n1572 , R_68a_1dfb3748 );
buf ( n1573 , R_9cf_1e183e28 );
buf ( n1574 , R_345_1d9d2668 );
buf ( n1575 , R_76b_1dfbbee8 );
buf ( n1576 , R_7aa_1e099328 );
buf ( n1577 , R_5e9_1ddacd48 );
buf ( n1578 , R_a04_1e185f48 );
buf ( n1579 , R_36b_1d9d3e28 );
buf ( n1580 , R_444_1d9dc5c8 );
buf ( n1581 , R_842_1e094aa8 );
buf ( n1582 , R_58a_1dda96e8 );
buf ( n1583 , R_97b_1e1809a8 );
buf ( n1584 , R_5bc_1ddab128 );
buf ( n1585 , R_ae9_1e6aeec8 );
buf ( n1586 , R_74e_1dfbc348 );
buf ( n1587 , R_69b_1dfb3ce8 );
buf ( n1588 , R_783_1dfbcde8 );
buf ( n1589 , R_64d_1dfb0c28 );
buf ( n1590 , R_938_1e17dfc8 );
buf ( n1591 , R_7bd_1e08f288 );
buf ( n1592 , R_7ca_1e08ffa8 );
buf ( n1593 , R_482_1ddac668 );
buf ( n1594 , R_2c7_1d9fd748 );
buf ( n1595 , R_621_1dfaf0a8 );
buf ( n1596 , R_9c3_1e1836a8 );
buf ( n1597 , R_309_1d9d00e8 );
buf ( n1598 , R_5f1_1ddad248 );
buf ( n1599 , R_4b8_1dda0ea8 );
buf ( n1600 , R_bcf_1e6b7e88 );
buf ( n1601 , R_824_1e0932e8 );
buf ( n1602 , R_6e6_1dfb70c8 );
buf ( n1603 , R_7a4_1e08e2e8 );
buf ( n1604 , R_59d_1dda9dc8 );
buf ( n1605 , R_769_1dfbbda8 );
buf ( n1606 , R_38a_1d9d5688 );
buf ( n1607 , R_4cb_1dda1a88 );
buf ( n1608 , R_8d9_1e09a408 );
buf ( n1609 , R_8d2_1e09a4a8 );
buf ( n1610 , R_b24_1e6b13a8 );
buf ( n1611 , R_4ba_1d9d9a08 );
buf ( n1612 , R_bdd_1e6b8748 );
buf ( n1613 , R_398_1d9d5a48 );
buf ( n1614 , R_31d_1d9d0d68 );
buf ( n1615 , R_47a_1dd9ece8 );
buf ( n1616 , R_2ca_1d9ce108 );
buf ( n1617 , R_b03_1e6aff08 );
buf ( n1618 , R_2a0_1d9fbee8 );
buf ( n1619 , R_71f_1dfb8f68 );
buf ( n1620 , R_950_1e17eec8 );
buf ( n1621 , R_9ce_1e184288 );
buf ( n1622 , R_aae_1e6b6c68 );
buf ( n1623 , R_b39_1e6b20c8 );
buf ( n1624 , R_906_1e090ea8 );
buf ( n1625 , R_786_1dfbd4c8 );
buf ( n1626 , R_81c_1e092de8 );
buf ( n1627 , R_94b_1e17eba8 );
buf ( n1628 , R_8fb_1e09b948 );
buf ( n1629 , R_3cb_1d9d7a28 );
buf ( n1630 , R_86f_1e0961c8 );
buf ( n1631 , R_584_1dda8e28 );
buf ( n1632 , R_40a_1d9da688 );
buf ( n1633 , R_954_1e17f148 );
buf ( n1634 , R_944_1e17e748 );
buf ( n1635 , R_bc8_1e6b7a28 );
buf ( n1636 , R_9a1_1e182168 );
buf ( n1637 , R_c02_1e6ba5e8 );
buf ( n1638 , R_967_1e17fd28 );
buf ( n1639 , R_7ff_1e091bc8 );
buf ( n1640 , R_329_1d9d14e8 );
buf ( n1641 , R_ba1_1e6b61c8 );
buf ( n1642 , R_717_1dfb8a68 );
buf ( n1643 , R_aa1_1e18c168 );
buf ( n1644 , R_591_1dda9648 );
buf ( n1645 , R_99c_1e181e48 );
buf ( n1646 , R_a42_1e188b08 );
buf ( n1647 , R_ba8_1e6b6628 );
buf ( n1648 , R_ae1_1e6ae9c8 );
buf ( n1649 , R_9c2_1e183b08 );
buf ( n1650 , R_6bb_1dfb50e8 );
buf ( n1651 , R_41b_1d9dac28 );
buf ( n1652 , R_93d_1e17e2e8 );
buf ( n1653 , R_5b2_1ddaafe8 );
buf ( n1654 , R_5d6_1d9dd388 );
buf ( n1655 , R_402_1d9da188 );
buf ( n1656 , R_4b0_1dda09a8 );
buf ( n1657 , R_549_1dda6948 );
buf ( n1658 , R_53a_1dda64e8 );
buf ( n1659 , R_70d_1dfb8428 );
buf ( n1660 , R_aa4_1e18c348 );
buf ( n1661 , R_798_1dfbdb08 );
buf ( n1662 , R_7fb_1e091948 );
buf ( n1663 , R_32a_1d9d1a88 );
buf ( n1664 , R_a36_1e188388 );
buf ( n1665 , R_5ed_1ddacfc8 );
buf ( n1666 , R_b9a_1e6b6268 );
buf ( n1667 , R_c07_1e6ba188 );
buf ( n1668 , R_47e_1dd9ef68 );
buf ( n1669 , R_ad2_1e6ae568 );
buf ( n1670 , R_39d_1d9d5d68 );
buf ( n1671 , R_83f_1e0943c8 );
buf ( n1672 , R_7eb_1e090f48 );
buf ( n1673 , R_42e_1d9dbd08 );
buf ( n1674 , R_b51_1e6b2fc8 );
buf ( n1675 , R_6b4_1dfb4c88 );
buf ( n1676 , R_694_1dfb3888 );
buf ( n1677 , R_68f_1dfb3568 );
buf ( n1678 , R_777_1dfbc668 );
buf ( n1679 , R_7b0_1e08ea68 );
buf ( n1680 , R_7a0_1e08e068 );
buf ( n1681 , R_75e_1dfbbbc8 );
buf ( n1682 , R_5b7_1ddaae08 );
buf ( n1683 , R_63d_1dfb0228 );
buf ( n1684 , R_636_1dfb02c8 );
buf ( n1685 , R_8de_1e09ac28 );
buf ( n1686 , R_2ef_1d9cf0a8 );
buf ( n1687 , R_302_1d9d4508 );
buf ( n1688 , R_9b8_1e182fc8 );
buf ( n1689 , R_4b2_1dda14e8 );
buf ( n1690 , R_8e4_1e09aae8 );
buf ( n1691 , R_3de_1d9d8b08 );
buf ( n1692 , R_ab8_1e18cfc8 );
buf ( n1693 , R_71b_1dfb8ce8 );
buf ( n1694 , R_c0c_1e6ba4a8 );
buf ( n1695 , R_c2b_1e6bb808 );
buf ( n1696 , R_5ac_1ddaa728 );
buf ( n1697 , R_853_1e095048 );
buf ( n1698 , R_2aa_1d9fca28 );
buf ( n1699 , R_385_1d9d4e68 );
buf ( n1700 , R_436_1d9dc208 );
buf ( n1701 , R_a60_1e1898c8 );
buf ( n1702 , R_7bb_1e08f148 );
buf ( n1703 , R_811_1e092708 );
buf ( n1704 , R_4c5_1dda16c8 );
buf ( n1705 , R_406_1d9da408 );
buf ( n1706 , R_473_1dd9e388 );
buf ( n1707 , R_8aa_1e098ba8 );
buf ( n1708 , R_b7e_1e6b50e8 );
buf ( n1709 , R_7b5_1e08ed88 );
buf ( n1710 , R_5fb_1ddad888 );
buf ( n1711 , R_34d_1d9d2b68 );
buf ( n1712 , R_ae3_1e6aeb08 );
buf ( n1713 , R_6f3_1dfb73e8 );
buf ( n1714 , R_82b_1e093748 );
buf ( n1715 , R_72a_1dfbacc8 );
buf ( n1716 , R_bc3_1e6b7708 );
buf ( n1717 , R_8fa_1e09bda8 );
buf ( n1718 , R_567_1dda7c08 );
buf ( n1719 , R_89f_1e097fc8 );
buf ( n1720 , R_3ed_1d9d8f68 );
buf ( n1721 , R_599_1dda9b48 );
buf ( n1722 , R_851_1e094f08 );
buf ( n1723 , R_2dd_1d9ce568 );
buf ( n1724 , R_4a8_1dda04a8 );
buf ( n1725 , R_8a9_1e098608 );
buf ( n1726 , R_366_1d9d4008 );
buf ( n1727 , R_376_1ddad568 );
buf ( n1728 , R_75d_1dfbb628 );
buf ( n1729 , R_59a_1ddaa0e8 );
buf ( n1730 , R_4c2_1dda19e8 );
buf ( n1731 , R_8be_1e08eba8 );
buf ( n1732 , R_2c5_1d9fd608 );
buf ( n1733 , R_595_1dda98c8 );
buf ( n1734 , R_446_1d9dd108 );
buf ( n1735 , R_6c5_1dfb5728 );
buf ( n1736 , R_5d8_1ddac2a8 );
buf ( n1737 , R_682_1dfb3248 );
buf ( n1738 , R_64b_1dfb0ae8 );
buf ( n1739 , R_791_1dfbd6a8 );
buf ( n1740 , R_b7b_1e6b4a08 );
buf ( n1741 , R_3b1_1d9d69e8 );
buf ( n1742 , R_7e9_1e090e08 );
buf ( n1743 , R_beb_1e6b9008 );
buf ( n1744 , R_6c0_1dfb5408 );
buf ( n1745 , R_8ba_1e0995a8 );
buf ( n1746 , R_a8e_1e17f508 );
buf ( n1747 , R_3c8_1d9d7848 );
buf ( n1748 , R_be4_1e6b8ba8 );
buf ( n1749 , R_544_1dda6628 );
buf ( n1750 , R_53f_1dda6308 );
buf ( n1751 , R_90e_1e09ca28 );
buf ( n1752 , R_381_1d9d4be8 );
buf ( n1753 , R_a3e_1e188888 );
buf ( n1754 , R_6fd_1dfb7a28 );
buf ( n1755 , R_a3a_1e188608 );
buf ( n1756 , R_8c2_1e099aa8 );
buf ( n1757 , R_af0_1e6af328 );
buf ( n1758 , R_296_1d9fb8a8 );
buf ( n1759 , R_b12_1e6b0d68 );
buf ( n1760 , R_ba9_1e6b66c8 );
buf ( n1761 , R_b1d_1e6b0f48 );
buf ( n1762 , R_2b5_1d9fcc08 );
buf ( n1763 , R_6ff_1dfb7b68 );
buf ( n1764 , R_a98_1e18bbc8 );
buf ( n1765 , R_58e_1dda9968 );
buf ( n1766 , R_753_1dfbafe8 );
buf ( n1767 , R_3c5_1d9d7668 );
buf ( n1768 , R_447_1d9dc7a8 );
buf ( n1769 , R_61f_1dfaef68 );
buf ( n1770 , R_54e_1dda28e8 );
buf ( n1771 , R_6f8_1dfb7708 );
buf ( n1772 , R_3a4_1d9d61c8 );
buf ( n1773 , R_423_1d9db128 );
buf ( n1774 , R_6a4_1dfb4288 );
buf ( n1775 , R_b9b_1e6b5e08 );
buf ( n1776 , R_a07_1e186128 );
buf ( n1777 , R_55f_1dda7708 );
buf ( n1778 , R_79d_1dfbde28 );
buf ( n1779 , R_66d_1dfb2028 );
buf ( n1780 , R_5e2_1ddacde8 );
buf ( n1781 , R_48b_1dd9f288 );
buf ( n1782 , R_5ee_1dda3a68 );
buf ( n1783 , R_6c6_1dfb2d48 );
buf ( n1784 , R_3e3_1d9d8928 );
buf ( n1785 , R_b83_1e6b4f08 );
buf ( n1786 , R_533_1dda5b88 );
buf ( n1787 , R_42d_1d9db768 );
buf ( n1788 , R_7e0_1e090868 );
buf ( n1789 , R_696_1dfb3ec8 );
buf ( n1790 , R_3f9_1d9d96e8 );
buf ( n1791 , R_b88_1e6b5228 );
buf ( n1792 , R_758_1dfbb308 );
buf ( n1793 , R_3d2_1d9d8388 );
buf ( n1794 , R_534_1dda5c28 );
buf ( n1795 , R_532_1d9d1308 );
buf ( n1796 , R_867_1e095cc8 );
buf ( n1797 , R_2b6_1d9fd1a8 );
buf ( n1798 , R_775_1dfbc528 );
buf ( n1799 , R_3e8_1d9d8c48 );
buf ( n1800 , R_4d0_1dda1da8 );
buf ( n1801 , R_30d_1d9d0368 );
buf ( n1802 , R_4e7_1dda2c08 );
buf ( n1803 , R_70a_1dfb8748 );
buf ( n1804 , R_a58_1e1893c8 );
buf ( n1805 , R_4e8_1dda2ca8 );
buf ( n1806 , R_4e6_1dda3068 );
buf ( n1807 , R_535_1dda5cc8 );
buf ( n1808 , R_5ea_1dda37e8 );
buf ( n1809 , R_929_1e09d608 );
buf ( n1810 , R_448_1d9dc848 );
buf ( n1811 , R_b0b_1e6b0408 );
buf ( n1812 , R_319_1d9d0ae8 );
buf ( n1813 , R_985_1e180fe8 );
buf ( n1814 , R_32f_1d9d18a8 );
buf ( n1815 , R_4e9_1dda2d48 );
buf ( n1816 , R_b1f_1e6b1088 );
buf ( n1817 , R_495_1dd9f8c8 );
buf ( n1818 , R_63b_1dfb00e8 );
buf ( n1819 , R_536_1dda6268 );
buf ( n1820 , R_3d9_1d9d82e8 );
buf ( n1821 , R_a4f_1e188e28 );
buf ( n1822 , R_470_1dd9e1a8 );
buf ( n1823 , R_2d5_1d9ce068 );
buf ( n1824 , R_3f0_1d9d9148 );
buf ( n1825 , R_acf_1e18de28 );
buf ( n1826 , R_ac2_1e18db08 );
buf ( n1827 , R_9b4_1e182d48 );
buf ( n1828 , R_a05_1e185fe8 );
buf ( n1829 , R_2d9_1d9ce2e8 );
buf ( n1830 , R_8ed_1e09b088 );
buf ( n1831 , R_3f3_1d9d9328 );
buf ( n1832 , R_af2_1e6af968 );
buf ( n1833 , R_44d_1d9dcb68 );
buf ( n1834 , R_645_1dfb0728 );
buf ( n1835 , R_648_1dfb0908 );
buf ( n1836 , R_4a1_1dda0048 );
buf ( n1837 , R_749_1dfba9a8 );
buf ( n1838 , R_2c8_1d9fd7e8 );
buf ( n1839 , R_3bc_1d9d70c8 );
buf ( n1840 , R_3f6_1ddad7e8 );
buf ( n1841 , R_596_1dda9e68 );
buf ( n1842 , R_c01_1e6b9dc8 );
buf ( n1843 , R_734_1dfb9c88 );
buf ( n1844 , R_5a5_1ddaa2c8 );
buf ( n1845 , R_6e3_1dfb69e8 );
buf ( n1846 , R_914_1e09c8e8 );
buf ( n1847 , R_43d_1d9dc168 );
buf ( n1848 , R_2cb_1d9fd9c8 );
buf ( n1849 , R_3d0_1d9d7d48 );
buf ( n1850 , R_b67_1e6b3d88 );
buf ( n1851 , R_b01_1e6afdc8 );
buf ( n1852 , R_37d_1d9d4968 );
buf ( n1853 , R_a80_1e18acc8 );
buf ( n1854 , R_9bd_1e1832e8 );
buf ( n1855 , R_339_1d9d1ee8 );
buf ( n1856 , R_7ad_1e08e888 );
buf ( n1857 , R_972_1e180908 );
buf ( n1858 , R_a22_1e184788 );
buf ( n1859 , R_486_1ddacb68 );
buf ( n1860 , R_5d5_1ddac0c8 );
buf ( n1861 , R_592_1dda9be8 );
buf ( n1862 , R_449_1d9dc8e8 );
buf ( n1863 , R_87b_1e096948 );
buf ( n1864 , R_8f5_1e09b588 );
buf ( n1865 , R_35a_1d9d3888 );
buf ( n1866 , R_37a_1ddab9e8 );
buf ( n1867 , R_991_1e181768 );
buf ( n1868 , R_62a_1dfb1448 );
buf ( n1869 , R_808_1e092168 );
buf ( n1870 , R_3a6_1d9d6808 );
buf ( n1871 , R_b95_1e6b5a48 );
buf ( n1872 , R_83e_1e17e108 );
buf ( n1873 , R_386_1d9d5408 );
buf ( n1874 , R_90d_1e09c488 );
buf ( n1875 , R_931_1e09db08 );
buf ( n1876 , R_ac9_1e18da68 );
buf ( n1877 , R_a31_1e187b68 );
buf ( n1878 , R_640_1dfb0408 );
buf ( n1879 , R_667_1dfb1c68 );
buf ( n1880 , R_6cb_1dfb5ae8 );
buf ( n1881 , R_74a_1e17f288 );
buf ( n1882 , R_676_1dfb2ac8 );
buf ( n1883 , R_372_1d9d4788 );
buf ( n1884 , R_56c_1dda7f28 );
buf ( n1885 , R_334_1d9d1bc8 );
buf ( n1886 , R_31e_1d9fc528 );
buf ( n1887 , R_981_1e180d68 );
buf ( n1888 , R_8ca_1e099fa8 );
buf ( n1889 , R_85e_1e095c28 );
buf ( n1890 , R_bbe_1e6af6e8 );
buf ( n1891 , R_49b_1dd9fc88 );
buf ( n1892 , R_73a_1dfba548 );
buf ( n1893 , R_5fe_1dfaf8c8 );
buf ( n1894 , R_98b_1e1813a8 );
buf ( n1895 , R_88e_1e097a28 );
buf ( n1896 , R_28f_1d9fb448 );
buf ( n1897 , R_9bc_1e183248 );
buf ( n1898 , R_5db_1ddac488 );
buf ( n1899 , R_88a_1e08ee28 );
buf ( n1900 , R_5a6_1ddaa868 );
buf ( n1901 , R_443_1d9dc528 );
buf ( n1902 , R_a0a_1e186808 );
buf ( n1903 , R_358_1d9d3248 );
buf ( n1904 , R_88f_1e0975c8 );
buf ( n1905 , R_acc_1e18dc48 );
buf ( n1906 , R_aac_1e18c848 );
buf ( n1907 , R_2a2_1d9fde28 );
buf ( n1908 , R_8a5_1e098388 );
buf ( n1909 , R_8ec_1e09afe8 );
buf ( n1910 , R_289_1d9fb088 );
buf ( n1911 , R_340_1d9d2348 );
buf ( n1912 , R_c2d_1e6bb948 );
buf ( n1913 , R_964_1e17fb48 );
buf ( n1914 , R_85d_1e095688 );
buf ( n1915 , R_6fa_1dfb7d48 );
buf ( n1916 , R_4d5_1dda20c8 );
buf ( n1917 , R_a5a_1e18b308 );
buf ( n1918 , R_7de_1e090c28 );
buf ( n1919 , R_605_1ddadec8 );
buf ( n1920 , R_311_1d9d05e8 );
buf ( n1921 , R_8a6_1e098928 );
buf ( n1922 , R_a2f_1e187a28 );
buf ( n1923 , R_81f_1e092fc8 );
buf ( n1924 , R_3b6_1d9d7208 );
buf ( n1925 , R_315_1d9d0868 );
buf ( n1926 , R_93f_1e17e428 );
buf ( n1927 , R_5b1_1ddaaa48 );
buf ( n1928 , R_631_1dfafaa8 );
buf ( n1929 , R_890_1e097668 );
buf ( n1930 , R_670_1dfb2208 );
buf ( n1931 , R_b9c_1e6b5ea8 );
buf ( n1932 , R_8e9_1e09ae08 );
buf ( n1933 , R_932_1e093928 );
buf ( n1934 , R_817_1e092ac8 );
buf ( n1935 , R_b60_1e6b3928 );
buf ( n1936 , R_979_1e180868 );
buf ( n1937 , R_8d8_1e09a368 );
buf ( n1938 , R_628_1dfaf508 );
buf ( n1939 , R_729_1dfb95a8 );
buf ( n1940 , R_a92_1e18bd08 );
buf ( n1941 , R_b33_1e6b1d08 );
buf ( n1942 , R_2ab_1d9fc5c8 );
buf ( n1943 , R_5e6_1dd9f6e8 );
buf ( n1944 , R_5c0_1ddab3a8 );
buf ( n1945 , R_600_1ddadba8 );
buf ( n1946 , R_8f4_1e09b4e8 );
buf ( n1947 , R_29d_1d9fbd08 );
buf ( n1948 , R_c11_1e6ba7c8 );
buf ( n1949 , R_4d7_1dda2208 );
buf ( n1950 , R_b43_1e6b2708 );
buf ( n1951 , R_881_1e096d08 );
buf ( n1952 , R_891_1e097708 );
buf ( n1953 , R_8b4_1e098ce8 );
buf ( n1954 , R_6ac_1dfb4788 );
buf ( n1955 , R_2f0_1d9cf148 );
buf ( n1956 , R_ad8_1e6ae428 );
buf ( n1957 , R_9bb_1e1831a8 );
buf ( n1958 , R_bd9_1e6b84c8 );
buf ( n1959 , R_39f_1d9d5ea8 );
buf ( n1960 , R_a5e_1e189c88 );
buf ( n1961 , R_303_1d9cfd28 );
buf ( n1962 , R_6ae_1dfb4dc8 );
buf ( n1963 , R_477_1dd9e608 );
buf ( n1964 , R_6d2_1e0981a8 );
buf ( n1965 , R_38f_1d9d54a8 );
buf ( n1966 , R_4d2_1dda23e8 );
buf ( n1967 , R_82f_1e0939c8 );
buf ( n1968 , R_61d_1dfaee28 );
buf ( n1969 , R_673_1dfb23e8 );
buf ( n1970 , R_578_1dda86a8 );
buf ( n1971 , R_a65_1e189be8 );
buf ( n1972 , R_9a5_1e1823e8 );
buf ( n1973 , R_744_1dfba688 );
buf ( n1974 , R_bfe_1e6ba0e8 );
buf ( n1975 , R_86e_1e096628 );
buf ( n1976 , R_6ce_1e0945a8 );
buf ( n1977 , R_9df_1e184828 );
buf ( n1978 , R_571_1dda8248 );
buf ( n1979 , R_9e0_1e1848c8 );
buf ( n1980 , R_9de_1e184c88 );
buf ( n1981 , R_41a_1ddabee8 );
buf ( n1982 , R_36e_1d9d1588 );
buf ( n1983 , R_6b9_1dfb4fa8 );
buf ( n1984 , R_b72_1e6b4968 );
buf ( n1985 , R_73f_1dfba368 );
buf ( n1986 , R_a4d_1e188ce8 );
buf ( n1987 , R_9e1_1e184968 );
buf ( n1988 , R_2d0_1d9fdce8 );
buf ( n1989 , R_72e_1dfb9dc8 );
buf ( n1990 , R_c25_1e6bb448 );
buf ( n1991 , R_8eb_1e09af48 );
buf ( n1992 , R_6eb_1dfb6ee8 );
buf ( n1993 , R_764_1dfbba88 );
buf ( n1994 , R_9b1_1e182b68 );
buf ( n1995 , R_970_1e1802c8 );
buf ( n1996 , R_bce_1e6b82e8 );
buf ( n1997 , R_325_1d9d1268 );
buf ( n1998 , R_65c_1dfb1588 );
buf ( n1999 , R_643_1dfb05e8 );
buf ( n2000 , R_abf_1e18d428 );
buf ( n2001 , R_a9b_1e18bda8 );
buf ( n2002 , R_b7c_1e6b4aa8 );
buf ( n2003 , R_9ba_1e183608 );
buf ( n2004 , R_bef_1e6b9288 );
buf ( n2005 , R_b14_1e6b09a8 );
buf ( n2006 , R_996_1e181f88 );
buf ( n2007 , R_812_1e092ca8 );
buf ( n2008 , R_4a2_1dda05e8 );
buf ( n2009 , R_6e0_1dfb6808 );
buf ( n2010 , R_490_1dd9f5a8 );
buf ( n2011 , R_711_1dfb86a8 );
buf ( n2012 , R_a86_1e18ba88 );
buf ( n2013 , R_342_1d9d2988 );
buf ( n2014 , R_c0e_1e6baae8 );
buf ( n2015 , R_8e3_1e09aa48 );
buf ( n2016 , R_646_1dfb0cc8 );
buf ( n2017 , R_74d_1dfbac28 );
buf ( n2018 , R_67f_1dfb2b68 );
buf ( n2019 , R_34f_1d9d2ca8 );
buf ( n2020 , R_8f3_1e09b448 );
buf ( n2021 , R_bdc_1e6b86a8 );
buf ( n2022 , R_57f_1dda8b08 );
buf ( n2023 , R_77a_1dfbcd48 );
buf ( n2024 , R_4c1_1dda1448 );
buf ( n2025 , R_b8e_1e6b5ae8 );
buf ( n2026 , R_c29_1e6bb6c8 );
buf ( n2027 , R_875_1e096588 );
buf ( n2028 , R_852_1e0954a8 );
buf ( n2029 , R_6a6_1dfb48c8 );
buf ( n2030 , R_76f_1dfbc168 );
buf ( n2031 , R_984_1e180f48 );
buf ( n2032 , R_39a_1d9d6088 );
buf ( n2033 , R_35f_1d9d36a8 );
buf ( n2034 , R_5d0_1ddabda8 );
buf ( n2035 , R_b65_1e6b3c48 );
buf ( n2036 , R_92b_1e09d748 );
buf ( n2037 , R_3eb_1d9d8e28 );
buf ( n2038 , R_53b_1dda6088 );
buf ( n2039 , R_97a_1e180e08 );
buf ( n2040 , R_369_1d9d3ce8 );
buf ( n2041 , R_7f5_1e091588 );
buf ( n2042 , R_588_1dda90a8 );
buf ( n2043 , R_b6a_1e6b4468 );
buf ( n2044 , R_435_1d9dbc68 );
buf ( n2045 , R_a08_1e1861c8 );
buf ( n2046 , R_7ef_1e0911c8 );
buf ( n2047 , R_781_1dfbcca8 );
buf ( n2048 , R_55c_1dda7528 );
buf ( n2049 , R_3bf_1d9d72a8 );
buf ( n2050 , R_850_1e094e68 );
buf ( n2051 , R_2ea_1d9cf288 );
buf ( n2052 , R_687_1dfb3068 );
buf ( n2053 , R_795_1dfbd928 );
buf ( n2054 , R_382_1d9d5188 );
buf ( n2055 , R_63e_1dfb07c8 );
buf ( n2056 , R_2b7_1d9fcd48 );
buf ( n2057 , R_9b0_1e182ac8 );
buf ( n2058 , R_6dd_1dfb6628 );
buf ( n2059 , R_4be_1dda1768 );
buf ( n2060 , R_bfd_1e6b9b48 );
buf ( n2061 , R_b0d_1e6b0548 );
buf ( n2062 , R_b9d_1e6b5f48 );
buf ( n2063 , R_b3a_1e6b2668 );
buf ( n2064 , R_4b9_1dda0f48 );
buf ( n2065 , R_4bb_1dda1088 );
buf ( n2066 , R_9a0_1e1820c8 );
buf ( n2067 , R_83b_1e094148 );
buf ( n2068 , R_8ea_1e09b3a8 );
buf ( n2069 , R_b21_1e6b11c8 );
buf ( n2070 , R_62f_1dfaf968 );
buf ( n2071 , R_91d_1e09ce88 );
buf ( n2072 , R_483_1dd9ed88 );
buf ( n2073 , R_7c0_1e08f468 );
buf ( n2074 , R_bd5_1e6b8248 );
buf ( n2075 , R_364_1d9d39c8 );
buf ( n2076 , R_322_1d9d2e88 );
buf ( n2077 , R_326_1d9d1808 );
buf ( n2078 , R_99b_1e181da8 );
buf ( n2079 , R_961_1e17f968 );
buf ( n2080 , R_726_1dfb98c8 );
buf ( n2081 , R_a7d_1e18aae8 );
buf ( n2082 , R_826_1e09de28 );
buf ( n2083 , R_89a_1dfb4648 );
buf ( n2084 , R_511_1dda4648 );
buf ( n2085 , R_2fb_1d9cf828 );
buf ( n2086 , R_b5c_1e6b36a8 );
buf ( n2087 , R_8b0_1e098a68 );
buf ( n2088 , R_708_1dfb8108 );
buf ( n2089 , R_603_1ddadd88 );
buf ( n2090 , R_804_1e091ee8 );
buf ( n2091 , R_573_1dda8388 );
buf ( n2092 , R_a56_1e189a08 );
buf ( n2093 , R_510_1dda45a8 );
buf ( n2094 , R_833_1e093c48 );
buf ( n2095 , R_8c1_1e099508 );
buf ( n2096 , R_966_1e180188 );
buf ( n2097 , R_46d_1dd9dfc8 );
buf ( n2098 , R_bcc_1e6b7ca8 );
buf ( n2099 , R_47b_1dd9e888 );
buf ( n2100 , R_aea_1e6af468 );
buf ( n2101 , R_8d1_1e099f08 );
buf ( n2102 , R_57a_1ddaa368 );
buf ( n2103 , R_8f2_1e09b8a8 );
buf ( n2104 , R_b35_1e6b1e48 );
buf ( n2105 , R_b05_1e6b0048 );
buf ( n2106 , R_aa9_1e18c668 );
buf ( n2107 , R_9b7_1e182f28 );
buf ( n2108 , R_3ae_1d9d6d08 );
buf ( n2109 , R_50f_1dda4508 );
buf ( n2110 , R_a23_1e1872a8 );
buf ( n2111 , R_2c9_1d9fd888 );
buf ( n2112 , R_5c6_1d9d7e88 );
buf ( n2113 , R_8bd_1e099288 );
buf ( n2114 , R_4b1_1dda0a48 );
buf ( n2115 , R_b45_1e6b2848 );
buf ( n2116 , R_422_1d9db588 );
buf ( n2117 , R_2cc_1d9fda68 );
buf ( n2118 , R_9d5_1e1841e8 );
buf ( n2119 , R_37e_1d9d4f08 );
buf ( n2120 , R_42c_1d9db6c8 );
buf ( n2121 , R_a7e_1e18b088 );
buf ( n2122 , R_a8d_1e18b4e8 );
buf ( n2123 , R_50e_1dda4968 );
buf ( n2124 , R_626_1dfafb48 );
buf ( n2125 , R_5cc_1ddabb28 );
buf ( n2126 , R_295_1d9fb808 );
buf ( n2127 , R_a9e_1e18c488 );
buf ( n2128 , R_80d_1e092488 );
buf ( n2129 , R_9af_1e182a28 );
buf ( n2130 , R_946_1e17ed88 );
buf ( n2131 , R_a5c_1e189648 );
buf ( n2132 , R_5bb_1ddab088 );
buf ( n2133 , R_3e6_1d9d9008 );
buf ( n2134 , R_ab3_1e18cca8 );
buf ( n2135 , R_a1e_1e187488 );
buf ( n2136 , R_66a_1dfb2348 );
buf ( n2137 , R_7f8_1e091768 );
buf ( n2138 , R_56e_1dda8568 );
buf ( n2139 , R_3c2_1d9d7988 );
buf ( n2140 , R_837_1e093ec8 );
buf ( n2141 , R_866_1e096128 );
buf ( n2142 , R_65a_1dfb1948 );
buf ( n2143 , R_4aa_1dda0ae8 );
buf ( n2144 , R_540_1dda63a8 );
buf ( n2145 , R_61b_1dfaece8 );
buf ( n2146 , R_78a_1dfbd748 );
buf ( n2147 , R_76c_1dfbbf88 );
buf ( n2148 , R_4c7_1dda1808 );
buf ( n2149 , R_47f_1dd9eb08 );
buf ( n2150 , R_34a_1d9d4a08 );
buf ( n2151 , R_b57_1e6b3388 );
buf ( n2152 , R_545_1dda66c8 );
buf ( n2153 , R_c13_1e6ba908 );
buf ( n2154 , R_44c_1d9dcac8 );
buf ( n2155 , R_a0b_1e1863a8 );
buf ( n2156 , R_6d5_1dfb6128 );
buf ( n2157 , R_bf3_1e6b9508 );
buf ( n2158 , R_3ee_1d9d9508 );
buf ( n2159 , R_6d7_1dfb6268 );
buf ( n2160 , R_3d6_1d9d9788 );
buf ( n2161 , R_b06_1e6b05e8 );
buf ( n2162 , R_9d4_1e184148 );
buf ( n2163 , R_33b_1d9d2028 );
buf ( n2164 , R_739_1dfb9fa8 );
buf ( n2165 , R_a0e_1e186a88 );
buf ( n2166 , R_7dd_1e090688 );
buf ( n2167 , R_54f_1dda6d08 );
buf ( n2168 , R_926_1e09dba8 );
buf ( n2169 , R_abb_1e18d1a8 );
buf ( n2170 , R_70e_1dfb89c8 );
buf ( n2171 , R_ba2_1e6b6768 );
buf ( n2172 , R_917_1e09cac8 );
buf ( n2173 , R_923_1e09d248 );
buf ( n2174 , R_784_1dfbce88 );
buf ( n2175 , R_920_1e09d068 );
buf ( n2176 , R_564_1dda7a28 );
buf ( n2177 , R_9a9_1e182668 );
buf ( n2178 , R_bfa_1e6b9e68 );
buf ( n2179 , R_62c_1dfaf788 );
buf ( n2180 , R_8c9_1e099a08 );
buf ( n2181 , R_43c_1d9dc0c8 );
buf ( n2182 , R_b00_1e6afd28 );
buf ( n2183 , R_35d_1d9d3568 );
buf ( n2184 , R_c18_1e6bac28 );
buf ( n2185 , R_306_1d9d0408 );
buf ( n2186 , R_939_1e17e068 );
buf ( n2187 , R_474_1dd9e428 );
buf ( n2188 , R_4a9_1dda0548 );
buf ( n2189 , R_2ac_1d9fc668 );
buf ( n2190 , R_609_1dfae1a8 );
buf ( n2191 , R_94c_1e17ec48 );
buf ( n2192 , R_90a_1e09c7a8 );
buf ( n2193 , R_92e_1e0918a8 );
buf ( n2194 , R_7be_1e08f828 );
buf ( n2195 , R_825_1e093388 );
buf ( n2196 , R_559_1dda7348 );
buf ( n2197 , R_bf7_1e6b9788 );
buf ( n2198 , R_87a_1e096da8 );
buf ( n2199 , R_9d3_1e1840a8 );
buf ( n2200 , R_394_1d9d57c8 );
buf ( n2201 , R_31a_1d9d1088 );
buf ( n2202 , R_69f_1dfb3f68 );
buf ( n2203 , R_787_1dfbd068 );
buf ( n2204 , R_a63_1e189aa8 );
buf ( n2205 , R_9ae_1e183388 );
buf ( n2206 , R_945_1e17e7e8 );
buf ( n2207 , R_537_1dda5e08 );
buf ( n2208 , R_725_1dfb9328 );
buf ( n2209 , R_b68_1e6b3e28 );
buf ( n2210 , R_7a5_1e08e388 );
buf ( n2211 , R_4eb_1dda2e88 );
buf ( n2212 , R_619_1dfaeba8 );
buf ( n2213 , R_800_1e091c68 );
buf ( n2214 , R_be8_1e6b8e28 );
buf ( n2215 , R_4ec_1dda2f28 );
buf ( n2216 , R_4ea_1dda32e8 );
buf ( n2217 , R_2f1_1d9cf1e8 );
buf ( n2218 , R_5d3_1ddabf88 );
buf ( n2219 , R_6da_1dfb6948 );
buf ( n2220 , R_5b6_1ddab268 );
buf ( n2221 , R_3ac_1d9d66c8 );
buf ( n2222 , R_983_1e180ea8 );
buf ( n2223 , R_b73_1e6b4508 );
buf ( n2224 , R_4ed_1dda2fc8 );
buf ( n2225 , R_ada_1e6aea68 );
buf ( n2226 , R_7fc_1e0919e8 );
buf ( n2227 , R_b3c_1e6b22a8 );
buf ( n2228 , R_304_1d9cfdc8 );
buf ( n2229 , R_5ab_1ddaa688 );
buf ( n2230 , R_85c_1e0955e8 );
buf ( n2231 , R_442_1d9dcc08 );
buf ( n2232 , R_3ce_1d9d8608 );
buf ( n2233 , R_ad5_1e6ae248 );
buf ( n2234 , R_ae8_1e6aee28 );
buf ( n2235 , R_3b4_1d9d6bc8 );
buf ( n2236 , R_8b8_1e098f68 );
buf ( n2237 , R_b46_1e6b2de8 );
buf ( n2238 , R_8e8_1e09ad68 );
buf ( n2239 , R_bbf_1e6b7488 );
buf ( n2240 , R_799_1dfbdba8 );
buf ( n2241 , R_778_1dfbc708 );
buf ( n2242 , R_a4b_1e188ba8 );
buf ( n2243 , R_51d_1dda4dc8 );
buf ( n2244 , R_657_1dfb1268 );
buf ( n2245 , R_9d2_1e17f788 );
buf ( n2246 , R_348_1d9d2848 );
buf ( n2247 , R_51c_1dda4d28 );
buf ( n2248 , R_8d7_1e09a2c8 );
buf ( n2249 , R_9b3_1e182ca8 );
buf ( n2250 , R_7db_1e090548 );
buf ( n2251 , R_715_1dfb8928 );
buf ( n2252 , R_68c_1dfb3388 );
buf ( n2253 , R_880_1e096c68 );
buf ( n2254 , R_29c_1d9fbc68 );
buf ( n2255 , R_b7d_1e6b4b48 );
buf ( n2256 , R_51b_1dda4c88 );
buf ( n2257 , R_bba_1e6b7668 );
buf ( n2258 , R_3dc_1d9d84c8 );
buf ( n2259 , R_5a0_1dda9fa8 );
buf ( n2260 , R_75f_1dfbb768 );
buf ( n2261 , R_b7f_1e6b4c88 );
buf ( n2262 , R_b16_1e6b0fe8 );
buf ( n2263 , R_ba3_1e6b6308 );
buf ( n2264 , R_654_1dfb1088 );
buf ( n2265 , R_bc7_1e6b7988 );
buf ( n2266 , R_2a3_1d9fc0c8 );
buf ( n2267 , R_6f0_1dfb7208 );
buf ( n2268 , R_7a1_1e08e108 );
buf ( n2269 , R_371_1d9d41e8 );
buf ( n2270 , R_51a_1dda50e8 );
buf ( n2271 , R_ab7_1e18cf28 );
buf ( n2272 , R_7e6_1e099828 );
buf ( n2273 , R_b6b_1e6b4008 );
buf ( n2274 , R_9ad_1e1828e8 );
buf ( n2275 , R_935_1e09dd88 );
buf ( n2276 , R_b8a_1e6bb768 );
buf ( n2277 , R_69d_1dfb3e28 );
buf ( n2278 , R_45e_1d9ddb08 );
buf ( n2279 , R_a1a_1e187208 );
buf ( n2280 , R_a49_1e188a68 );
buf ( n2281 , R_a09_1e186268 );
buf ( n2282 , R_496_1dd9fe68 );
buf ( n2283 , R_336_1d9d2208 );
buf ( n2284 , R_5df_1ddac708 );
buf ( n2285 , R_5c7_1ddab808 );
buf ( n2286 , R_990_1e1816c8 );
buf ( n2287 , R_6c9_1dfb59a8 );
buf ( n2288 , R_2eb_1d9cee28 );
buf ( n2289 , R_2b8_1d9fcde8 );
buf ( n2290 , R_ae0_1e6ae928 );
buf ( n2291 , R_b2f_1e6b1a88 );
buf ( n2292 , R_84d_1e094c88 );
buf ( n2293 , R_a12_1e186d08 );
buf ( n2294 , R_74f_1dfbad68 );
buf ( n2295 , R_a35_1e187de8 );
buf ( n2296 , R_28e_1d9fb3a8 );
buf ( n2297 , R_81a_1e0936a8 );
buf ( n2298 , R_487_1dd9f008 );
buf ( n2299 , R_c1c_1e6baea8 );
buf ( n2300 , R_7a8_1e08e568 );
buf ( n2301 , R_471_1dd9e248 );
buf ( n2302 , R_766_1e0986a8 );
buf ( n2303 , R_38b_1d9d5228 );
buf ( n2304 , R_a7b_1e18a9a8 );
buf ( n2305 , R_b52_1e6b8568 );
buf ( n2306 , R_9ff_1e185c28 );
buf ( n2307 , R_7b9_1e08f008 );
buf ( n2308 , R_67b_1dfb28e8 );
buf ( n2309 , R_a00_1e185cc8 );
buf ( n2310 , R_9fe_1e6bb9e8 );
buf ( n2311 , R_980_1e180cc8 );
buf ( n2312 , R_874_1e0964e8 );
buf ( n2313 , R_49c_1dd9fd28 );
buf ( n2314 , R_58c_1dda9328 );
buf ( n2315 , R_45f_1d9dd6a8 );
buf ( n2316 , R_98a_1e181808 );
buf ( n2317 , R_8e2_1e09aea8 );
buf ( n2318 , R_6ba_1dfb5548 );
buf ( n2319 , R_bd8_1e6b8428 );
buf ( n2320 , R_a8b_1e18b3a8 );
buf ( n2321 , R_a01_1e185d68 );
buf ( n2322 , R_6b3_1dfb4be8 );
buf ( n2323 , R_60d_1dfae428 );
buf ( n2324 , R_6e8_1dfb6d08 );
buf ( n2325 , R_399_1d9d5ae8 );
buf ( n2326 , R_a16_1e186f88 );
buf ( n2327 , R_bc2_1e6b7b68 );
buf ( n2328 , R_32b_1d9d1628 );
buf ( n2329 , R_434_1d9dbbc8 );
buf ( n2330 , R_a24_1e187348 );
buf ( n2331 , R_377_1d9d45a8 );
buf ( n2332 , R_3cc_1d9d7ac8 );
buf ( n2333 , R_a68_1e189dc8 );
buf ( n2334 , R_963_1e17faa8 );
buf ( n2335 , R_7c5_1e08f788 );
buf ( n2336 , R_615_1dfae928 );
buf ( n2337 , R_8a2_1dfb9b48 );
buf ( n2338 , R_722_1dfb9648 );
buf ( n2339 , R_288_1d9f96e8 );
buf ( n2340 , R_556_1dda7668 );
buf ( n2341 , R_748_1dfba908 );
buf ( n2342 , R_865_1e095b88 );
buf ( n2343 , R_607_1dfae068 );
buf ( n2344 , R_691_1dfb36a8 );
buf ( n2345 , R_978_1e1807c8 );
buf ( n2346 , R_84f_1e094dc8 );
buf ( n2347 , R_2cd_1d9fdb08 );
buf ( n2348 , R_ae2_1e6aef68 );
buf ( n2349 , R_a1f_1e187028 );
buf ( n2350 , R_721_1dfb90a8 );
buf ( n2351 , R_733_1dfb9be8 );
buf ( n2352 , R_9e3_1e184aa8 );
buf ( n2353 , R_9e4_1e184b48 );
buf ( n2354 , R_c23_1e6bb308 );
buf ( n2355 , R_9e2_1e184f08 );
buf ( n2356 , R_7ae_1dfbb1c8 );
buf ( n2357 , R_91a_1e09d1a8 );
buf ( n2358 , R_b84_1e6b4fa8 );
buf ( n2359 , R_b92_1e181088 );
buf ( n2360 , R_ba4_1e6b63a8 );
buf ( n2361 , R_754_1dfbb088 );
buf ( n2362 , R_5a4_1ddaa228 );
buf ( n2363 , R_9a4_1e182348 );
buf ( n2364 , R_b08_1e6b0228 );
buf ( n2365 , R_9e5_1e184be8 );
buf ( n2366 , R_617_1dfaea68 );
buf ( n2367 , R_5ce_1ddac168 );
buf ( n2368 , R_b89_1e6b52c8 );
buf ( n2369 , R_7b2_1e09b128 );
buf ( n2370 , R_460_1d9dd748 );
buf ( n2371 , R_5e4_1ddaca28 );
buf ( n2372 , R_30a_1d9d0688 );
buf ( n2373 , R_a0c_1e186448 );
buf ( n2374 , R_910_1e09c668 );
buf ( n2375 , R_553_1dda6f88 );
buf ( n2376 , R_86d_1e096088 );
buf ( n2377 , R_a0f_1e186628 );
buf ( n2378 , R_719_1dfb8ba8 );
buf ( n2379 , R_b48_1e6b2a28 );
buf ( n2380 , R_316_1d9d0e08 );
buf ( n2381 , R_901_1e09bd08 );
buf ( n2382 , R_611_1dfae6a8 );
buf ( n2383 , R_ac5_1e18d7e8 );
buf ( n2384 , R_6c4_1dfb5688 );
buf ( n2385 , R_53c_1dda6128 );
buf ( n2386 , R_712_1dfb8c48 );
buf ( n2387 , R_2f6_1d9cfc88 );
buf ( n2388 , R_829_1e093608 );
buf ( n2389 , R_89d_1e097e88 );
buf ( n2390 , R_8d0_1e099e68 );
buf ( n2391 , R_8ac_1e0987e8 );
buf ( n2392 , R_8a0_1e098068 );
buf ( n2393 , R_aef_1e6af288 );
buf ( n2394 , R_759_1dfbb3a8 );
buf ( n2395 , R_a6d_1e18a0e8 );
buf ( n2396 , R_6bf_1dfb5368 );
buf ( n2397 , R_982_1e182c08 );
buf ( n2398 , R_bdb_1e6b8608 );
buf ( n2399 , R_684_1dfb2e88 );
buf ( n2400 , R_7b7_1e08eec8 );
buf ( n2401 , R_478_1dd9e6a8 );
buf ( n2402 , R_be1_1e6b89c8 );
buf ( n2403 , R_b55_1e6b3248 );
buf ( n2404 , R_79b_1dfbdce8 );
buf ( n2405 , R_c27_1e6bb588 );
buf ( n2406 , R_96f_1e180228 );
buf ( n2407 , R_42b_1d9db628 );
buf ( n2408 , R_6cd_1dfb5c28 );
buf ( n2409 , R_652_1dfb16c8 );
buf ( n2410 , R_71d_1dfb8e28 );
buf ( n2411 , R_703_1dfb7de8 );
buf ( n2412 , R_a54_1e189148 );
buf ( n2413 , R_4a3_1dda0188 );
buf ( n2414 , R_634_1dfafc88 );
buf ( n2415 , R_2ad_1d9fc708 );
buf ( n2416 , R_4cc_1dda1b28 );
buf ( n2417 , R_2a1_1d9fbf88 );
buf ( n2418 , R_93a_1e0977a8 );
buf ( n2419 , R_a78_1e18a7c8 );
buf ( n2420 , R_c03_1e6b9f08 );
buf ( n2421 , R_72c_1dfb9788 );
buf ( n2422 , R_809_1e092208 );
buf ( n2423 , R_5b0_1ddaa9a8 );
buf ( n2424 , R_44b_1d9dca28 );
buf ( n2425 , R_952_1ddab768 );
buf ( n2426 , R_899_1e097c08 );
buf ( n2427 , R_bd4_1e6b81a8 );
buf ( n2428 , R_a94_1e18b948 );
buf ( n2429 , R_6b1_1dfb4aa8 );
buf ( n2430 , R_491_1dd9f648 );
buf ( n2431 , R_5ca_1d9dae08 );
buf ( n2432 , R_6f5_1dfb7528 );
buf ( n2433 , R_9c9_1e183a68 );
buf ( n2434 , R_75a_1dfbb948 );
buf ( n2435 , R_461_1d9dd7e8 );
buf ( n2436 , R_7c3_1e08f648 );
buf ( n2437 , R_569_1dda7d48 );
buf ( n2438 , R_a75_1e18a5e8 );
buf ( n2439 , R_7ec_1e090fe8 );
buf ( n2440 , R_c20_1e6bb128 );
buf ( n2441 , R_96d_1e1800e8 );
buf ( n2442 , R_54a_1dda6ee8 );
buf ( n2443 , R_b31_1e6b1bc8 );
buf ( n2444 , R_5bf_1ddab308 );
buf ( n2445 , R_900_1e09bc68 );
buf ( n2446 , R_b74_1e6b45a8 );
buf ( n2447 , R_940_1e17e4c8 );
buf ( n2448 , R_8dd_1e09a688 );
buf ( n2449 , R_a88_1e18b1c8 );
buf ( n2450 , R_743_1dfba5e8 );
buf ( n2451 , R_2d1_1d9fdd88 );
buf ( n2452 , R_4b3_1dda0b88 );
buf ( n2453 , R_48c_1dd9f328 );
buf ( n2454 , R_419_1d9daae8 );
buf ( n2455 , R_2ba_1d9fd428 );
buf ( n2456 , R_898_1e097b68 );
buf ( n2457 , R_354_1d9d2fc8 );
buf ( n2458 , R_3c9_1d9d78e8 );
buf ( n2459 , R_afd_1e6afb48 );
buf ( n2460 , R_698_1dfb3b08 );
buf ( n2461 , R_8c8_1e099968 );
buf ( n2462 , R_aff_1e6afc88 );
buf ( n2463 , R_59c_1dda9d28 );
buf ( n2464 , R_43b_1d9dc028 );
buf ( n2465 , R_3e1_1d9d87e8 );
buf ( n2466 , R_7d8_1e090368 );
buf ( n2467 , R_624_1dfaf288 );
buf ( n2468 , R_ace_1e6ae2e8 );
buf ( n2469 , R_294_1d9fb768 );
buf ( n2470 , R_818_1e092b68 );
buf ( n2471 , R_9c8_1e1839c8 );
buf ( n2472 , R_5c8_1ddab8a8 );
buf ( n2473 , R_c2f_1e6bba88 );
buf ( n2474 , R_ba5_1e6b6448 );
buf ( n2475 , R_6d0_1dfb5e08 );
buf ( n2476 , R_820_1e093068 );
buf ( n2477 , R_30e_1d9d0908 );
buf ( n2478 , R_99f_1e182028 );
buf ( n2479 , R_73e_1dfba7c8 );
buf ( n2480 , R_4ef_1dda3108 );
buf ( n2481 , R_451_1d9dcde8 );
buf ( n2482 , R_678_1dfb2708 );
buf ( n2483 , R_663_1dfb19e8 );
buf ( n2484 , R_5fa_1e091128 );
buf ( n2485 , R_312_1d9d0b88 );
buf ( n2486 , R_a45_1e1887e8 );
buf ( n2487 , R_b18_1e6b0c28 );
buf ( n2488 , R_4f0_1dda31a8 );
buf ( n2489 , R_4ee_1dda3568 );
buf ( n2490 , R_7ab_1e08e748 );
buf ( n2491 , R_305_1d9cfe68 );
buf ( n2492 , R_955_1e17f1e8 );
buf ( n2493 , R_373_1d9d4328 );
buf ( n2494 , R_a39_1e188068 );
buf ( n2495 , R_669_1dfb1da8 );
buf ( n2496 , R_3a5_1d9d6268 );
buf ( n2497 , R_c0d_1e6ba548 );
buf ( n2498 , R_4f1_1dda3248 );
buf ( n2499 , R_541_1dda6448 );
buf ( n2500 , R_69a_1dfb4148 );
buf ( n2501 , R_b90_1e6b5728 );
buf ( n2502 , R_99a_1e182208 );
buf ( n2503 , R_960_1e17f8c8 );
buf ( n2504 , R_6a9_1dfb45a8 );
buf ( n2505 , R_4bc_1dda1128 );
buf ( n2506 , R_897_1e097ac8 );
buf ( n2507 , R_701_1dfb7ca8 );
buf ( n2508 , R_36c_1d9d3ec8 );
buf ( n2509 , R_60b_1dfae2e8 );
buf ( n2510 , R_583_1dda8d88 );
buf ( n2511 , R_330_1d9d1948 );
buf ( n2512 , R_bb6_1e6b73e8 );
buf ( n2513 , R_71e_1dfb93c8 );
buf ( n2514 , R_590_1dda95a8 );
buf ( n2515 , R_29e_1dda2668 );
buf ( n2516 , R_b0f_1e6b0688 );
buf ( n2517 , R_a1b_1e186da8 );
buf ( n2518 , R_550_1dda6da8 );
buf ( n2519 , R_ac8_1e18d9c8 );
buf ( n2520 , R_a9d_1e18bee8 );
buf ( n2521 , R_561_1dda7848 );
buf ( n2522 , R_80e_1e092a28 );
buf ( n2523 , R_9b6_1e187708 );
buf ( n2524 , R_5e8_1ddacca8 );
buf ( n2525 , R_613_1dfae7e8 );
buf ( n2526 , R_b6c_1e6b40a8 );
buf ( n2527 , R_3d3_1d9d7f28 );
buf ( n2528 , R_31f_1d9d0ea8 );
buf ( n2529 , R_9c7_1e183928 );
buf ( n2530 , R_5dd_1ddac5c8 );
buf ( n2531 , R_78e_1dfbd9c8 );
buf ( n2532 , R_a13_1e1868a8 );
buf ( n2533 , R_70c_1dfb8388 );
buf ( n2534 , R_885_1e096f88 );
buf ( n2535 , R_85b_1e095548 );
buf ( n2536 , R_8ff_1e09bbc8 );
buf ( n2537 , R_716_1dfb8ec8 );
buf ( n2538 , R_2b9_1d9fce88 );
buf ( n2539 , R_b69_1e6b3ec8 );
buf ( n2540 , R_356_1d9d3608 );
buf ( n2541 , R_2e6_1d9cf008 );
buf ( n2542 , R_484_1dd9ee28 );
buf ( n2543 , R_2ec_1d9ceec8 );
buf ( n2544 , R_acb_1e18dba8 );
buf ( n2545 , R_813_1e092848 );
buf ( n2546 , R_4c3_1dda1588 );
buf ( n2547 , R_a47_1e188928 );
buf ( n2548 , R_81d_1e092e88 );
buf ( n2549 , R_8e7_1e09acc8 );
buf ( n2550 , R_5ef_1ddad108 );
buf ( n2551 , R_896_1e094828 );
buf ( n2552 , R_bec_1e6b90a8 );
buf ( n2553 , R_b2b_1e6b1808 );
buf ( n2554 , R_4ab_1dda0688 );
buf ( n2555 , R_7e4_1e090ae8 );
buf ( n2556 , R_a33_1e187ca8 );
buf ( n2557 , R_47c_1dd9e928 );
buf ( n2558 , R_8d6_1e09a728 );
buf ( n2559 , R_87f_1e096bc8 );
buf ( n2560 , R_5b5_1ddaacc8 );
buf ( n2561 , R_651_1dfb0ea8 );
buf ( n2562 , R_3da_1d9d8888 );
buf ( n2563 , R_538_1dda5ea8 );
buf ( n2564 , R_675_1dfb2528 );
buf ( n2565 , R_60f_1dfae568 );
buf ( n2566 , R_29b_1d9fbbc8 );
buf ( n2567 , R_aa6_1e18c988 );
buf ( n2568 , R_3bd_1d9d7168 );
buf ( n2569 , R_be5_1e6b8c48 );
buf ( n2570 , R_c0a_1e6ba868 );
buf ( n2571 , R_5f5_1ddad4c8 );
buf ( n2572 , R_b4b_1e6b2c08 );
buf ( n2573 , R_7b1_1e08eb08 );
buf ( n2574 , R_95d_1e17f6e8 );
buf ( n2575 , R_a17_1e186b28 );
buf ( n2576 , R_a29_1e187668 );
buf ( n2577 , R_71a_1dfb9148 );
buf ( n2578 , R_693_1dfb37e8 );
buf ( n2579 , R_77b_1dfbc8e8 );
buf ( n2580 , R_9c6_1e183d88 );
buf ( n2581 , R_3a7_1d9d63a8 );
buf ( n2582 , R_bc0_1e6b7528 );
buf ( n2583 , R_68e_1dfb39c8 );
buf ( n2584 , R_335_1d9d1c68 );
buf ( n2585 , R_5eb_1ddace88 );
buf ( n2586 , R_ad7_1e6ae388 );
buf ( n2587 , R_765_1dfbbb28 );
buf ( n2588 , R_387_1d9d4fa8 );
buf ( n2589 , R_9a8_1e1825c8 );
buf ( n2590 , R_632_1dfb0048 );
buf ( n2591 , R_6e5_1dfb6b28 );
buf ( n2592 , R_772_1dfbc848 );
buf ( n2593 , R_995_1e1819e8 );
buf ( n2594 , R_7d6_1e090728 );
buf ( n2595 , R_598_1dda9aa8 );
buf ( n2596 , R_a70_1e18a2c8 );
buf ( n2597 , R_a25_1e1873e8 );
buf ( n2598 , R_bbb_1e6b7208 );
buf ( n2599 , R_6f2_1dfb7848 );
buf ( n2600 , R_a41_1e188568 );
buf ( n2601 , R_a66_1e18a188 );
buf ( n2602 , R_a3d_1e1882e8 );
buf ( n2603 , R_341_1d9d23e8 );
buf ( n2604 , R_594_1dda9828 );
buf ( n2605 , R_4fe_1dda5868 );
buf ( n2606 , R_480_1dd9eba8 );
buf ( n2607 , R_6ab_1dfb46e8 );
buf ( n2608 , R_84c_1e094be8 );
buf ( n2609 , R_660_1dfb1808 );
buf ( n2610 , R_a20_1e1870c8 );
buf ( n2611 , R_abe_1e6b64e8 );
buf ( n2612 , R_566_1dda8068 );
buf ( n2613 , R_7c8_1e08f968 );
buf ( n2614 , R_5c2_1d9fc2a8 );
buf ( n2615 , R_989_1e181268 );
buf ( n2616 , R_8a8_1e098568 );
buf ( n2617 , R_2a4_1d9fc168 );
buf ( n2618 , R_7d5_1e090188 );
buf ( n2619 , R_8fe_1e09c028 );
buf ( n2620 , R_3b7_1d9d6da8 );
buf ( n2621 , R_6b8_1dfb4f08 );
buf ( n2622 , R_8b3_1e098c48 );
buf ( n2623 , R_94f_1e17ee28 );
buf ( n2624 , R_9fb_1e1859a8 );
buf ( n2625 , R_a10_1e1866c8 );
buf ( n2626 , R_b36_1e6b23e8 );
buf ( n2627 , R_aa0_1e18c0c8 );
buf ( n2628 , R_c1a_1e6bb268 );
buf ( n2629 , R_82c_1e0937e8 );
buf ( n2630 , R_4d1_1dda1e48 );
buf ( n2631 , R_6fc_1dfb7988 );
buf ( n2632 , R_9fa_1e185e08 );
buf ( n2633 , R_9fc_1e185a48 );
buf ( n2634 , R_a0d_1e1864e8 );
buf ( n2635 , R_be2_1e6b8f68 );
buf ( n2636 , R_b02_1e6b8068 );
buf ( n2637 , R_a28_1e1875c8 );
buf ( n2638 , R_4fd_1dda39c8 );
buf ( n2639 , R_5fd_1ddad9c8 );
buf ( n2640 , R_873_1e096448 );
buf ( n2641 , R_9fd_1e185ae8 );
buf ( n2642 , R_a6b_1e189fa8 );
buf ( n2643 , R_aa3_1e18c2a8 );
buf ( n2644 , R_738_1dfb9f08 );
buf ( n2645 , R_805_1e091f88 );
buf ( n2646 , R_2f7_1d9cf5a8 );
buf ( n2647 , R_5ba_1ddab4e8 );
buf ( n2648 , R_57d_1dda89c8 );
buf ( n2649 , R_475_1dd9e4c8 );
buf ( n2650 , R_433_1d9dbb28 );
buf ( n2651 , R_aed_1e6af148 );
buf ( n2652 , R_4fc_1dda3928 );
buf ( n2653 , R_3a0_1d9d5f48 );
buf ( n2654 , R_3f7_1d9d95a8 );
buf ( n2655 , R_367_1d9d3ba8 );
buf ( n2656 , R_947_1e17e928 );
buf ( n2657 , R_b1a_1e6b1268 );
buf ( n2658 , R_525_1dda52c8 );
buf ( n2659 , R_50d_1dda43c8 );
buf ( n2660 , R_390_1d9d5548 );
buf ( n2661 , R_6fe_1dfb7fc8 );
buf ( n2662 , R_6f7_1dfb7668 );
buf ( n2663 , R_2ae_1d9fcca8 );
buf ( n2664 , R_864_1e095ae8 );
buf ( n2665 , R_9e7_1e184d28 );
buf ( n2666 , R_524_1dda5228 );
buf ( n2667 , R_50c_1dda4328 );
buf ( n2668 , R_9e6_1e185188 );
buf ( n2669 , R_9e8_1e184dc8 );
buf ( n2670 , R_9b2_1e183108 );
buf ( n2671 , R_7e2_1dfbaf48 );
buf ( n2672 , R_622_1dfaf648 );
buf ( n2673 , R_b4e_1e184508 );
buf ( n2674 , R_a91_1e18b768 );
buf ( n2675 , R_a84_1e18af48 );
buf ( n2676 , R_4ce_1dda2168 );
buf ( n2677 , R_bb2_1e6b7168 );
buf ( n2678 , R_523_1dda5188 );
buf ( n2679 , R_50b_1dda4288 );
buf ( n2680 , R_9e9_1e184e68 );
buf ( n2681 , R_4f3_1dda3388 );
buf ( n2682 , R_4fb_1dda3888 );
buf ( n2683 , R_4f2_1ddad068 );
buf ( n2684 , R_4f4_1dda3428 );
buf ( n2685 , R_55e_1dda7b68 );
buf ( n2686 , R_84e_1e095228 );
buf ( n2687 , R_a76_1e18ab88 );
buf ( n2688 , R_5c9_1ddab948 );
buf ( n2689 , R_343_1d9d2528 );
buf ( n2690 , R_a73_1e18a4a8 );
buf ( n2691 , R_7cd_1e08fc88 );
buf ( n2692 , R_522_1dda55e8 );
buf ( n2693 , R_50a_1dda46e8 );
buf ( n2694 , R_4f5_1dda34c8 );
buf ( n2695 , R_396_1d9d5e08 );
buf ( n2696 , R_7f9_1e091808 );
buf ( n2697 , R_681_1dfb2ca8 );
buf ( n2698 , R_37b_1d9d4828 );
buf ( n2699 , R_639_1dfaffa8 );
buf ( n2700 , R_76d_1dfbc028 );
buf ( n2701 , R_78b_1dfbd2e8 );
buf ( n2702 , R_6a3_1dfb41e8 );
buf ( n2703 , R_9ac_1e182848 );
buf ( n2704 , R_86c_1e095fe8 );
buf ( n2705 , R_c08_1e6ba228 );
buf ( n2706 , R_2fc_1d9cf8c8 );
buf ( n2707 , R_7f0_1e091268 );
buf ( n2708 , R_c31_1e6bbbc8 );
buf ( n2709 , R_a52_1e189508 );
buf ( n2710 , R_ab2_1e18d108 );
buf ( n2711 , R_28d_1d9fb308 );
buf ( n2712 , R_bcb_1e6b7c08 );
buf ( n2713 , R_4fa_1dda3f68 );
buf ( n2714 , R_2bb_1d9fcfc8 );
buf ( n2715 , R_b3f_1e6b2488 );
buf ( n2716 , R_a27_1e187528 );
buf ( n2717 , R_362_1d9d3d88 );
buf ( n2718 , R_497_1dd9fa08 );
buf ( n2719 , R_64f_1dfb0d68 );
buf ( n2720 , R_bd7_1e6b8388 );
buf ( n2721 , R_b75_1e6b4648 );
buf ( n2722 , R_98f_1e181628 );
buf ( n2723 , R_6ed_1dfb7028 );
buf ( n2724 , R_7d3_1e090048 );
buf ( n2725 , R_b27_1e6b1588 );
buf ( n2726 , R_39b_1d9d5c28 );
buf ( n2727 , R_8cf_1e099dc8 );
buf ( n2728 , R_689_1dfb31a8 );
buf ( n2729 , R_7c6_1e08fd28 );
buf ( n2730 , R_b2d_1e6b1948 );
buf ( n2731 , R_92a_1e092f28 );
buf ( n2732 , R_66c_1dfb1f88 );
buf ( n2733 , R_956_1e6b00e8 );
buf ( n2734 , R_b96_1e18ce88 );
buf ( n2735 , R_bae_1e6b6ee8 );
buf ( n2736 , R_94d_1e17ece8 );
buf ( n2737 , R_785_1dfbcf28 );
buf ( n2738 , R_6e2_1dfb6e48 );
buf ( n2739 , R_65e_1dfb5cc8 );
buf ( n2740 , R_42a_1d9dba88 );
buf ( n2741 , R_7e8_1e090d68 );
buf ( n2742 , R_b4d_1e6b2d48 );
buf ( n2743 , R_bff_1e6b9c88 );
buf ( n2744 , R_3c0_1d9d7348 );
buf ( n2745 , R_44a_1d9dce88 );
buf ( n2746 , R_2fe_1d9cff08 );
buf ( n2747 , R_383_1d9d4d28 );
buf ( n2748 , R_928_1e09d568 );
buf ( n2749 , R_488_1dd9f0a8 );
buf ( n2750 , R_5aa_1ddaaae8 );
buf ( n2751 , R_3fd_1d9d9968 );
buf ( n2752 , R_7d0_1e08fe68 );
buf ( n2753 , R_7b4_1e08ece8 );
buf ( n2754 , R_4d8_1dda22a8 );
buf ( n2755 , R_418_1d9daa48 );
buf ( n2756 , R_a43_1e1886a8 );
buf ( n2757 , R_327_1d9d13a8 );
buf ( n2758 , R_849_1e094a08 );
buf ( n2759 , R_b5f_1e6b3888 );
buf ( n2760 , R_4d3_1dda1f88 );
buf ( n2761 , R_a97_1e18bb28 );
buf ( n2762 , R_aba_1e18d608 );
buf ( n2763 , R_ab1_1e18cb68 );
buf ( n2764 , R_97f_1e180c28 );
buf ( n2765 , R_788_1dfbd108 );
buf ( n2766 , R_a1c_1e186e48 );
buf ( n2767 , R_b11_1e6b07c8 );
buf ( n2768 , R_a37_1e187f28 );
buf ( n2769 , R_801_1e091d08 );
buf ( n2770 , R_581_1dda8c48 );
buf ( n2771 , R_49d_1dd9fdc8 );
buf ( n2772 , R_56b_1dda7e88 );
buf ( n2773 , R_4da_1dda3ce8 );
buf ( n2774 , R_7f2_1e09d6a8 );
buf ( n2775 , R_53d_1dda61c8 );
buf ( n2776 , R_3df_1d9d86a8 );
buf ( n2777 , R_429_1d9db4e8 );
buf ( n2778 , R_8dc_1e09a5e8 );
buf ( n2779 , R_a14_1e186948 );
buf ( n2780 , R_9d6_1e186088 );
buf ( n2781 , R_add_1e6ae748 );
buf ( n2782 , R_b6d_1e6b4148 );
buf ( n2783 , R_c1e_1e6b4e68 );
buf ( n2784 , R_7fd_1e091a88 );
buf ( n2785 , R_859_1e095408 );
buf ( n2786 , R_b23_1e6b1308 );
buf ( n2787 , R_afc_1e6afaa8 );
buf ( n2788 , R_913_1e09c848 );
buf ( n2789 , R_450_1d9dcd48 );
buf ( n2790 , R_7cb_1e08fb48 );
buf ( n2791 , R_b38_1e6b2028 );
buf ( n2792 , R_a26_1e187988 );
buf ( n2793 , R_74c_1dfbab88 );
buf ( n2794 , R_35b_1d9d3428 );
buf ( n2795 , R_962_1e17ff08 );
buf ( n2796 , R_2e7_1d9ceba8 );
buf ( n2797 , R_8c0_1e099468 );
buf ( n2798 , R_8c7_1e0998c8 );
buf ( n2799 , R_afe_1e6b5d68 );
buf ( n2800 , R_977_1e180728 );
buf ( n2801 , R_925_1e09d388 );
buf ( n2802 , R_919_1e09cc08 );
buf ( n2803 , R_728_1dfb9508 );
buf ( n2804 , R_43a_1d9dc488 );
buf ( n2805 , R_bf0_1e6b9328 );
buf ( n2806 , R_9a3_1e1822a8 );
buf ( n2807 , R_3af_1d9d68a8 );
buf ( n2808 , R_930_1e09da68 );
buf ( n2809 , R_90c_1e09c3e8 );
buf ( n2810 , R_5a9_1ddaa548 );
buf ( n2811 , R_659_1dfb13a8 );
buf ( n2812 , R_c0f_1e6ba688 );
buf ( n2813 , R_307_1d9cffa8 );
buf ( n2814 , R_8bc_1e0991e8 );
buf ( n2815 , R_2ed_1d9cef68 );
buf ( n2816 , R_770_1dfbc208 );
buf ( n2817 , R_34b_1d9d2a28 );
buf ( n2818 , R_37f_1d9d4aa8 );
buf ( n2819 , R_5f4_1ddad428 );
buf ( n2820 , R_779_1dfbc7a8 );
buf ( n2821 , R_46a_1dd9f468 );
buf ( n2822 , R_be0_1e6b8928 );
buf ( n2823 , R_bd3_1e6b8108 );
buf ( n2824 , R_466_1d9d9c88 );
buf ( n2825 , R_77e_1dfbcfc8 );
buf ( n2826 , R_575_1dda84c8 );
buf ( n2827 , R_4ff_1dda3b08 );
buf ( n2828 , R_a18_1e186bc8 );
buf ( n2829 , R_bda_1e6b8a68 );
buf ( n2830 , R_31b_1d9d0c28 );
buf ( n2831 , R_3c6_1d9d7c08 );
buf ( n2832 , R_792_1dfbdc48 );
buf ( n2833 , R_54b_1dda6a88 );
buf ( n2834 , R_6bd_1dfb5228 );
buf ( n2835 , R_b50_1e6b2f28 );
buf ( n2836 , R_a61_1e189968 );
buf ( n2837 , R_b8b_1e6b5408 );
buf ( n2838 , R_b80_1e6b4d28 );
buf ( n2839 , R_33c_1d9d20c8 );
buf ( n2840 , R_3c3_1d9d7528 );
buf ( n2841 , R_666_1dfb20c8 );
buf ( n2842 , R_c2a_1e6bbc68 );
buf ( n2843 , R_359_1d9d32e8 );
buf ( n2844 , R_415_1d9da868 );
buf ( n2845 , R_5da_1ddac8e8 );
buf ( n2846 , R_577_1dda8608 );
buf ( n2847 , R_637_1dfafe68 );
buf ( n2848 , R_9f7_1e185728 );
buf ( n2849 , R_570_1dda81a8 );
buf ( n2850 , R_9f6_1e185b88 );
buf ( n2851 , R_9f8_1e1857c8 );
buf ( n2852 , R_a6e_1e18a688 );
buf ( n2853 , R_73d_1dfba228 );
buf ( n2854 , R_293_1d9fb6c8 );
buf ( n2855 , R_884_1e096ee8 );
buf ( n2856 , R_3a2_1d9d6588 );
buf ( n2857 , R_9f9_1e185868 );
buf ( n2858 , R_957_1e17f328 );
buf ( n2859 , R_ab6_1e6b5fe8 );
buf ( n2860 , R_760_1dfbb808 );
buf ( n2861 , R_a21_1e187168 );
buf ( n2862 , R_bb7_1e6b6f88 );
buf ( n2863 , R_9eb_1e184fa8 );
buf ( n2864 , R_a3f_1e188428 );
buf ( n2865 , R_747_1dfba868 );
buf ( n2866 , R_4bf_1dda1308 );
buf ( n2867 , R_3d7_1d9d81a8 );
buf ( n2868 , R_4a4_1dda0228 );
buf ( n2869 , R_441_1d9dc3e8 );
buf ( n2870 , R_7ce_1e090228 );
buf ( n2871 , R_85a_1e0959a8 );
buf ( n2872 , R_66f_1dfb2168 );
buf ( n2873 , R_9ea_1e185408 );
buf ( n2874 , R_9ec_1e185048 );
buf ( n2875 , R_a3b_1e1881a8 );
buf ( n2876 , R_ad4_1e6ae1a8 );
buf ( n2877 , R_b94_1e6b59a8 );
buf ( n2878 , R_467_1d9ddba8 );
buf ( n2879 , R_96e_1e180688 );
buf ( n2880 , R_323_1d9d1128 );
buf ( n2881 , R_6ea_1dfb7348 );
buf ( n2882 , R_6ca_1dfb5f48 );
buf ( n2883 , R_9ed_1e1850e8 );
buf ( n2884 , R_ae7_1e6aed88 );
buf ( n2885 , R_830_1e093a68 );
buf ( n2886 , R_6d9_1dfb63a8 );
buf ( n2887 , R_8e6_1e08f0a8 );
buf ( n2888 , R_6a1_1dfb40a8 );
buf ( n2889 , R_710_1dfb8608 );
buf ( n2890 , R_b41_1e6b25c8 );
buf ( n2891 , R_732_1dfba048 );
buf ( n2892 , R_6df_1dfb6768 );
buf ( n2893 , R_a11_1e186768 );
buf ( n2894 , R_a8f_1e18b628 );
buf ( n2895 , R_b97_1e6b5b88 );
buf ( n2896 , R_bc6_1e6b7de8 );
buf ( n2897 , R_4db_1dda2488 );
buf ( n2898 , R_9d7_1e184328 );
buf ( n2899 , R_b29_1e6b16c8 );
buf ( n2900 , R_57e_1dda8f68 );
buf ( n2901 , R_29a_1d9fbb28 );
buf ( n2902 , R_36f_1d9d40a8 );
buf ( n2903 , R_3e4_1d9d89c8 );
buf ( n2904 , R_7bc_1e08f1e8 );
buf ( n2905 , R_87e_1e097028 );
buf ( n2906 , R_b1c_1e6b0ea8 );
buf ( n2907 , R_aab_1e18c7a8 );
buf ( n2908 , R_96c_1e180048 );
buf ( n2909 , R_551_1dda6e48 );
buf ( n2910 , R_6d4_1dfb6088 );
buf ( n2911 , R_2af_1d9fc848 );
buf ( n2912 , R_479_1dd9e748 );
buf ( n2913 , R_5a3_1ddaa188 );
buf ( n2914 , R_672_1dfb2848 );
buf ( n2915 , R_587_1dda9008 );
buf ( n2916 , R_767_1dfbbc68 );
buf ( n2917 , R_395_1d9d5868 );
buf ( n2918 , R_3e9_1d9d8ce8 );
buf ( n2919 , R_2f8_1d9cf648 );
buf ( n2920 , R_64c_1dfb0b88 );
buf ( n2921 , R_5e1_1ddac848 );
buf ( n2922 , R_3fc_1d9d98c8 );
buf ( n2923 , R_468_1d9ddc48 );
buf ( n2924 , R_3ba_1d9d7488 );
buf ( n2925 , R_55b_1dda7488 );
buf ( n2926 , R_67e_1dfb2fc8 );
buf ( n2927 , R_8b7_1e098ec8 );
buf ( n2928 , R_879_1e096808 );
buf ( n2929 , R_b5b_1e6b3608 );
buf ( n2930 , R_a82_1e18b588 );
buf ( n2931 , R_ae5_1e6aec48 );
buf ( n2932 , R_84b_1e094b48 );
buf ( n2933 , R_99e_1e182488 );
buf ( n2934 , R_6dc_1dfb6588 );
buf ( n2935 , R_3ad_1d9d6768 );
buf ( n2936 , R_a59_1e189468 );
buf ( n2937 , R_b62_1e6ba368 );
buf ( n2938 , R_731_1dfb9aa8 );
buf ( n2939 , R_3f1_1d9d91e8 );
buf ( n2940 , R_620_1dfaf008 );
buf ( n2941 , R_67d_1dfb2a28 );
buf ( n2942 , R_adf_1e6ae888 );
buf ( n2943 , R_349_1d9d28e8 );
buf ( n2944 , R_3d1_1d9d7de8 );
buf ( n2945 , R_3f4_1d9d93c8 );
buf ( n2946 , R_80a_1e0927a8 );
buf ( n2947 , R_350_1d9d2d48 );
buf ( n2948 , R_a50_1e188ec8 );
buf ( n2949 , R_bc1_1e6b75c8 );
buf ( n2950 , R_b85_1e6b5048 );
buf ( n2951 , R_5d7_1ddac208 );
buf ( n2952 , R_7a2_1ddada68 );
buf ( n2953 , R_539_1dda5f48 );
buf ( n2954 , R_bbc_1e6b72a8 );
buf ( n2955 , R_c14_1e6ba9a8 );
buf ( n2956 , R_6c8_1dfb5908 );
buf ( n2957 , R_4c8_1dda18a8 );
buf ( n2958 , R_360_1d9d3748 );
buf ( n2959 , R_2e2_1d9ced88 );
buf ( n2960 , R_936_1e17e388 );
buf ( n2961 , R_9f3_1e1854a8 );
buf ( n2962 , R_b25_1e6b1448 );
buf ( n2963 , R_b0a_1e6b0868 );
buf ( n2964 , R_b56_1e6b87e8 );
buf ( n2965 , R_bf4_1e6b95a8 );
buf ( n2966 , R_95f_1e17f828 );
buf ( n2967 , R_3b5_1d9d6c68 );
buf ( n2968 , R_52a_1dda5fe8 );
buf ( n2969 , R_9f2_1e185908 );
buf ( n2970 , R_9f4_1e185548 );
buf ( n2971 , R_686_1dfb34c8 );
buf ( n2972 , R_2bc_1d9fd068 );
buf ( n2973 , R_7a6_1e08e928 );
buf ( n2974 , R_9ef_1e185228 );
buf ( n2975 , R_b1e_1e6b78e8 );
buf ( n2976 , R_bfb_1e6b9a08 );
buf ( n2977 , R_378_1d9d4648 );
buf ( n2978 , R_9ee_1e185688 );
buf ( n2979 , R_9f0_1e1852c8 );
buf ( n2980 , R_9f5_1e1855e8 );
buf ( n2981 , R_4bd_1dda11c8 );
buf ( n2982 , R_5af_1ddaa908 );
buf ( n2983 , R_822_1e097f28 );
buf ( n2984 , R_872_1e0968a8 );
buf ( n2985 , R_9f1_1e185368 );
buf ( n2986 , R_337_1d9d1da8 );
buf ( n2987 , R_707_1dfb8068 );
buf ( n2988 , R_755_1dfbb128 );
buf ( n2989 , R_8f9_1e09b808 );
buf ( n2990 , R_432_1d9dbf88 );
buf ( n2991 , R_8af_1e0989c8 );
buf ( n2992 , R_bc5_1e6b7848 );
buf ( n2993 , R_934_1e09dce8 );
buf ( n2994 , R_469_1d9ddce8 );
buf ( n2995 , R_572_1dda87e8 );
buf ( n2996 , R_863_1e095a48 );
buf ( n2997 , R_958_1e17f3c8 );
buf ( n2998 , R_742_1dfbaa48 );
buf ( n2999 , R_2a5_1d9fc208 );
buf ( n3000 , R_a9a_1e18c208 );
buf ( n3001 , R_af9_1e6af8c8 );
buf ( n3002 , R_9c1_1e183568 );
buf ( n3003 , R_83c_1e0941e8 );
buf ( n3004 , R_a81_1e18ad68 );
buf ( n3005 , R_c19_1e6bacc8 );
buf ( n3006 , R_91c_1e09cde8 );
buf ( n3007 , R_4ac_1dda0728 );
buf ( n3008 , R_bf8_1e6b9828 );
buf ( n3009 , R_5be_1dda7168 );
buf ( n3010 , R_93b_1e17e1a8 );
buf ( n3011 , R_63c_1dfb0188 );
buf ( n3012 , R_7e1_1e090908 );
buf ( n3013 , R_7ba_1e08f5a8 );
buf ( n3014 , R_6b2_1dfb5048 );
buf ( n3015 , R_4dc_1dda2528 );
buf ( n3016 , R_79e_1e08e428 );
buf ( n3017 , R_492_1dd9fbe8 );
buf ( n3018 , R_750_1dfbae08 );
buf ( n3019 , R_9d8_1e1843c8 );
buf ( n3020 , R_365_1d9d3a68 );
buf ( n3021 , R_994_1e181948 );
buf ( n3022 , R_95c_1e17f648 );
buf ( n3023 , R_2ff_1d9cfaa8 );
buf ( n3024 , R_89b_1e097d48 );
buf ( n3025 , R_827_1e0934c8 );
buf ( n3026 , R_332_1d9d1f88 );
buf ( n3027 , R_9a7_1e182528 );
buf ( n3028 , R_834_1e093ce8 );
buf ( n3029 , R_30b_1d9d0228 );
buf ( n3030 , R_86b_1e095f48 );
buf ( n3031 , R_649_1dfb09a8 );
buf ( n3032 , R_a1d_1e186ee8 );
buf ( n3033 , R_b59_1e6b34c8 );
buf ( n3034 , R_bb3_1e6b6d08 );
buf ( n3035 , R_796_1e08e1a8 );
buf ( n3036 , R_941_1e17e568 );
buf ( n3037 , R_be9_1e6b8ec8 );
buf ( n3038 , R_485_1dd9eec8 );
buf ( n3039 , R_317_1d9d09a8 );
buf ( n3040 , R_8a3_1e098248 );
buf ( n3041 , R_49e_1dda0368 );
buf ( n3042 , R_9c0_1e1834c8 );
buf ( n3043 , R_32c_1d9d16c8 );
buf ( n3044 , R_6d6_1dfb66c8 );
buf ( n3045 , R_a15_1e1869e8 );
buf ( n3046 , R_33e_1d9d2708 );
buf ( n3047 , R_38c_1d9d52c8 );
buf ( n3048 , R_75b_1dfbb4e8 );
buf ( n3049 , R_ac4_1e18d748 );
buf ( n3050 , R_5d9_1ddac348 );
buf ( n3051 , R_546_1dda6c68 );
buf ( n3052 , R_2be_1d9fd6a8 );
buf ( n3053 , R_b76_1e6b4be8 );
buf ( n3054 , R_975_1e1805e8 );
buf ( n3055 , R_5c3_1ddab588 );
buf ( n3056 , R_500_1dda3ba8 );
buf ( n3057 , R_889_1e097208 );
buf ( n3058 , R_988_1e1811c8 );
buf ( n3059 , R_c2c_1e6bb8a8 );
buf ( n3060 , R_b98_1e6b5c28 );
buf ( n3061 , R_47d_1dd9e9c8 );
buf ( n3062 , R_417_1d9da9a8 );
buf ( n3063 , R_819_1e092c08 );
buf ( n3064 , R_8f8_1e09b768 );
buf ( n3065 , R_942_1e17eb08 );
buf ( n3066 , R_ad1_1e6adfc8 );
buf ( n3067 , R_8ce_1e09a228 );
buf ( n3068 , R_563_1dda7988 );
buf ( n3069 , R_2e8_1d9cec48 );
buf ( n3070 , R_838_1e093f68 );
buf ( n3071 , R_aee_1e187c08 );
buf ( n3072 , R_641_1dfb04a8 );
buf ( n3073 , R_c16_1e6b41e8 );
buf ( n3074 , R_6c3_1dfb55e8 );
buf ( n3075 , R_5f3_1ddad388 );
buf ( n3076 , R_558_1dda72a8 );
buf ( n3077 , R_821_1e093108 );
buf ( n3078 , R_a5f_1e189828 );
buf ( n3079 , R_3cd_1d9d7b68 );
buf ( n3080 , R_80f_1e0925c8 );
buf ( n3081 , R_724_1dfb9288 );
buf ( n3082 , R_848_1e094968 );
buf ( n3083 , R_9bf_1e183428 );
buf ( n3084 , R_a19_1e186c68 );
buf ( n3085 , R_baf_1e6b6a88 );
buf ( n3086 , R_64a_1dfb0f48 );
buf ( n3087 , R_aa8_1e18c5c8 );
buf ( n3088 , R_6be_1dfb57c8 );
buf ( n3089 , R_481_1dd9ec48 );
buf ( n3090 , R_428_1d9db448 );
buf ( n3091 , R_be6_1e6b91e8 );
buf ( n3092 , R_44f_1d9dcca8 );
buf ( n3093 , R_5b4_1ddaac28 );
buf ( n3094 , R_629_1dfaf5a8 );
buf ( n3095 , R_78f_1dfbd568 );
buf ( n3096 , R_91f_1e09cfc8 );
buf ( n3097 , R_858_1e095368 );
buf ( n3098 , R_afb_1e6afa08 );
buf ( n3099 , R_3fb_1d9d9828 );
buf ( n3100 , R_922_1e091628 );
buf ( n3101 , R_916_1e09cf28 );
buf ( n3102 , R_8a1_1e098108 );
buf ( n3103 , R_8db_1e09a548 );
buf ( n3104 , R_b32_1e6b2168 );
buf ( n3105 , R_411_1d9da5e8 );
buf ( n3106 , R_6b0_1dfb4a08 );
buf ( n3107 , R_5d1_1ddabe48 );
buf ( n3108 , R_7df_1e0907c8 );
buf ( n3109 , R_b04_1e6affa8 );
buf ( n3110 , R_45a_1d9dd888 );
buf ( n3111 , R_814_1e0928e8 );
buf ( n3112 , R_665_1dfb1b28 );
buf ( n3113 , R_69e_1dfb43c8 );
buf ( n3114 , R_b42_1e6b2b68 );
buf ( n3115 , R_555_1dda70c8 );
buf ( n3116 , R_374_1d9d43c8 );
buf ( n3117 , R_352_1d9d3388 );
buf ( n3118 , R_2a6_1d9fc7a8 );
buf ( n3119 , R_756_1dfbb6c8 );
buf ( n3120 , R_bd6_1e6b3568 );
buf ( n3121 , R_baa_1e18d888 );
buf ( n3122 , R_5b9_1ddaaf48 );
buf ( n3123 , R_3ec_1d9d8ec8 );
buf ( R_61e_1dfaf3c8 , C0 );
buf ( R_8f7_1e09b6c8 , n275553 );
buf ( R_714_1dfb8888 , n275555 );
buf ( R_951_1e17ef68 , n275559 );
buf ( R_28c_1d9fb268 , n275924 );
buf ( R_9be_1e183888 , C0 );
buf ( R_9ab_1e1827a8 , n275928 );
buf ( R_30f_1d9d04a8 , n275932 );
buf ( R_959_1e17f468 , n12699 );
buf ( R_b13_1e6b0908 , n12702 );
buf ( R_519_1dda4b48 , n17569 );
buf ( R_92d_1e09d888 , n19393 );
buf ( R_c06_1e6bafe8 , C0 );
buf ( R_8c6_1e099d28 , C0 );
buf ( R_845_1e094788 , n20573 );
buf ( R_414_1d9da7c8 , n20574 );
buf ( R_313_1d9d0728 , n20577 );
buf ( R_518_1dda4aa8 , n20578 );
buf ( R_9d9_1e184468 , n20662 );
buf ( R_4dd_1dda25c8 , n20704 );
buf ( R_59f_1dda9f08 , n20707 );
buf ( R_517_1dda4a08 , n20710 );
buf ( R_509_1dda4148 , n20818 );
buf ( R_508_1dda40a8 , n20819 );
buf ( R_401_1d9d9be8 , n20957 );
buf ( R_5f9_1ddad748 , n20964 );
buf ( R_6ef_1dfb7168 , n20967 );
buf ( R_a30_1e187ac8 , n20968 );
buf ( R_2b0_1d9fc8e8 , n20969 );
buf ( R_77c_1dfbc988 , n20970 );
buf ( R_8f1_1e09b308 , n21035 );
buf ( R_36a_1d9d4288 , C0 );
buf ( R_507_1dda4008 , n21038 );
buf ( R_516_1dda4e68 , C0 );
buf ( R_98e_1e181a88 , C0 );
buf ( R_8d5_1e09a188 , n21634 );
buf ( R_498_1dd9faa8 , n21635 );
buf ( R_68b_1dfb32e8 , n21638 );
buf ( R_773_1dfbc3e8 , n21641 );
buf ( R_45b_1d9dd428 , n21644 );
buf ( R_48d_1dd9f3c8 , n21702 );
buf ( R_5ff_1ddadb08 , n21705 );
buf ( R_705_1dfb7f28 , n21778 );
buf ( R_644_1dfb0688 , n21779 );
buf ( R_63a_1dfb0548 , C0 );
buf ( R_ac7_1e18d928 , n21782 );
buf ( R_320_1d9d0f48 , n21783 );
buf ( R_737_1dfb9e68 , n21786 );
buf ( R_506_1dda4468 , C0 );
buf ( R_647_1dfb0868 , n21789 );
buf ( R_b86_1e6bb4e8 , C0 );
buf ( R_883_1e096e48 , n21792 );
buf ( R_6a8_1dfb4508 , n21793 );
buf ( R_aa5_1e18c3e8 , n22199 );
buf ( R_440_1d9dc348 , n22200 );
buf ( R_2f9_1d9cf6e8 , n22333 );
buf ( R_69c_1dfb3d88 , n22334 );
buf ( R_65d_1dfb1628 , n22795 );
buf ( R_b0c_1e6b04a8 , n22796 );
buf ( R_b20_1e6b1128 , n22797 );
buf ( R_a2e_1e189788 , C0 );
buf ( R_905_1e09bf88 , n22882 );
buf ( R_a57_1e189328 , n22885 );
buf ( R_5f8_1ddad6a8 , n22886 );
buf ( R_54c_1dda6b28 , n22887 );
buf ( R_bd2_1e6b32e8 , C0 );
buf ( R_aca_1e6ae068 , C0 );
buf ( R_58b_1dda9288 , n22890 );
buf ( R_2e3_1d9ce928 , n22893 );
buf ( R_3e2_1d9d8d88 , C0 );
buf ( R_8f6_1e09bb28 , C0 );
buf ( R_331_1d9d19e8 , n23378 );
buf ( R_97d_1e180ae8 , n23385 );
buf ( R_5cd_1ddabbc8 , n23457 );
buf ( R_45c_1d9dd4c8 , n23458 );
buf ( R_999_1e181c68 , n23464 );
buf ( R_b99_1e6b5cc8 , n23712 );
buf ( R_948_1e17e9c8 , n23713 );
buf ( R_97e_1e181308 , C0 );
buf ( R_ab0_1e18cac8 , n23714 );
buf ( R_bb8_1e6b7028 , n23715 );
buf ( R_489_1dd9f148 , n23796 );
buf ( R_4b6_1dda1268 , C0 );
buf ( R_63f_1dfb0368 , n23799 );
buf ( R_3e7_1d9d8ba8 , n23802 );
buf ( R_2bd_1d9fd108 , n23811 );
buf ( R_81b_1e092d48 , n23814 );
buf ( R_b54_1e6b31a8 , n23815 );
buf ( R_4df_1dda2708 , n23818 );
buf ( R_bab_1e6b6808 , n23821 );
buf ( R_431_1d9db9e8 , n23892 );
buf ( R_2f2_1d9cf788 , C0 );
buf ( R_601_1ddadc48 , n23898 );
buf ( R_6e7_1dfb6c68 , n23901 );
buf ( R_bdf_1e6b8888 , n23904 );
buf ( R_656_1dfb1bc8 , C0 );
buf ( R_4e0_1dda27a8 , n23905 );
buf ( R_4de_1dda2b68 , C0 );
buf ( R_a4e_1e189288 , C0 );
buf ( R_8e1_1e09a908 , n24335 );
buf ( R_8f0_1e09b268 , n24336 );
buf ( R_299_1d9fba88 , n24344 );
buf ( R_292_1d9fb628 , n24356 );
buf ( R_4e1_1dda2848 , n24372 );
buf ( R_a7f_1e18ac28 , n24375 );
buf ( R_c04_1e6b9fa8 , n24376 );
buf ( R_3ef_1d9d90a8 , n24379 );
buf ( R_5de_1dd9f1e8 , C0 );
buf ( R_878_1e096768 , n24380 );
buf ( R_720_1dfb9008 , n24381 );
buf ( R_ad6_1e6ae7e8 , C0 );
buf ( R_9a2_1e182708 , C0 );
buf ( R_630_1dfafa08 , n24382 );
buf ( R_52f_1dda5908 , n24385 );
buf ( R_7a9_1e08e608 , n24456 );
buf ( R_976_1e180b88 , C0 );
buf ( R_439_1d9dbee8 , n24628 );
buf ( R_604_1ddade28 , n24629 );
buf ( R_530_1dda59a8 , n24630 );
buf ( R_52e_1dda5d68 , C0 );
buf ( R_7ed_1e091088 , n24669 );
buf ( R_3f2_1d9d4c88 , C0 );
buf ( R_3d4_1d9d7fc8 , n24670 );
buf ( R_84a_1e094fa8 , C0 );
buf ( R_2de_1d9ceb08 , C0 );
buf ( R_690_1dfb3608 , n24671 );
buf ( R_4cd_1dda1bc8 , n24733 );
buf ( R_531_1dda5a48 , n25035 );
buf ( R_b34_1e6b1da8 , n25036 );
buf ( R_5f7_1ddad608 , n25040 );
buf ( R_806_1e092528 , C0 );
buf ( R_a5b_1e1895a8 , n25043 );
buf ( R_718_1dfb8b08 , n25044 );
buf ( R_695_1dfb3928 , n26330 );
buf ( R_7af_1e08e9c8 , n26333 );
buf ( R_62b_1dfaf6e8 , n26336 );
buf ( R_904_1e09bee8 , n26337 );
buf ( R_501_1dda3c48 , n26356 );
buf ( R_585_1dda8ec8 , n26403 );
buf ( R_9cd_1e183ce8 , n26412 );
buf ( R_78c_1dfbd388 , n26413 );
buf ( R_392_1d9d5b88 , C0 );
buf ( R_4b4_1dda0c28 , n26414 );
buf ( R_b44_1e6b27a8 , n26415 );
buf ( R_969_1e17fe68 , n26422 );
buf ( R_40d_1d9da368 , n26507 );
buf ( R_627_1dfaf468 , n26510 );
buf ( R_67a_1dfadfc8 , C0 );
buf ( R_45d_1d9dd568 , n26515 );
buf ( R_7c1_1e08f508 , n27089 );
buf ( R_552_1dda73e8 , C0 );
buf ( R_2bf_1d9fd248 , n27092 );
buf ( R_5d4_1ddac028 , n27093 );
buf ( R_b77_1e6b4788 , n27096 );
buf ( R_3fa_1d9db088 , C0 );
buf ( R_6aa_1dfb4b48 , C0 );
buf ( R_82a_1e093ba8 , C0 );
buf ( R_3aa_1d9d6a88 , C0 );
buf ( R_300_1d9cfb48 , n27097 );
buf ( R_405_1d9d9e68 , n27170 );
buf ( R_953_1e17f0a8 , n27174 );
buf ( R_3cf_1d9d7ca8 , n27177 );
buf ( R_ac1_1e18d568 , n27530 );
buf ( R_61c_1dfaed88 , n27531 );
buf ( R_a99_1e18bc68 , n27596 );
buf ( R_4ae_1dda0fe8 , C0 );
buf ( R_aec_1e6af0a8 , n27597 );
buf ( R_af8_1e6af828 , n27598 );
buf ( R_762_1dfbbe48 , C0 );
buf ( R_3a8_1d9d6448 , n27599 );
buf ( R_4ca_1dda1ee8 , C0 );
buf ( R_6b7_1dfb4e68 , n27602 );
buf ( R_57c_1dda8928 , n27603 );
buf ( R_52b_1dda5688 , n27606 );
buf ( R_8ef_1e09b1c8 , n27609 );
buf ( R_8c5_1e099788 , n27629 );
buf ( R_8ab_1e098748 , n27632 );
buf ( R_71c_1dfb8d88 , n27633 );
buf ( R_388_1d9d5048 , n27634 );
buf ( R_b6e_1e6b46e8 , C0 );
buf ( R_9cc_1e183c48 , n27635 );
buf ( R_65b_1dfb14e8 , n27638 );
buf ( R_bbd_1e6b7348 , n27645 );
buf ( R_3b2_1d9d6f88 , C0 );
buf ( R_862_1e095ea8 , C0 );
buf ( R_4a5_1dda02c8 , n27651 );
buf ( R_90f_1e09c5c8 , n27654 );
buf ( R_702_1dfb8248 , C0 );
buf ( R_29f_1d9fbe48 , n27657 );
buf ( R_72b_1dfb96e8 , n27660 );
buf ( R_6f4_1dfb7488 , n27661 );
buf ( R_5f2_1dda8a68 , C0 );
buf ( R_a64_1e189b48 , n27662 );
buf ( R_2e9_1d9cece8 , n27672 );
buf ( R_683_1dfb2de8 , n27675 );
buf ( R_2fd_1d9cf968 , n27681 );
buf ( R_8b2_1e0990a8 , C0 );
buf ( R_5f0_1ddad1a8 , n27682 );
buf ( R_bac_1e6b68a8 , n27683 );
buf ( R_642_1dfb0a48 , C0 );
buf ( R_5f6_1d9fbda8 , C0 );
buf ( R_568_1dda7ca8 , n27684 );
buf ( R_409_1d9da0e8 , n27747 );
buf ( R_5a8_1ddaa4a8 , n27748 );
buf ( R_5e3_1ddac988 , n27751 );
buf ( R_96b_1e17ffa8 , n27754 );
buf ( R_bca_1e6b14e8 , C0 );
buf ( R_3b8_1d9d6e48 , n27755 );
buf ( R_789_1dfbd1a8 , n28152 );
buf ( R_86a_1e0963a8 , C0 );
buf ( R_416_1ddabc68 , C0 );
buf ( R_903_1e09be48 , n28155 );
buf ( R_a2d_1e1878e8 , n28162 );
buf ( R_9cb_1e183ba8 , n28165 );
buf ( R_59b_1dda9c88 , n28168 );
buf ( R_a4c_1e188c48 , n28169 );
buf ( R_79c_1dfbdd88 , n28170 );
buf ( R_888_1e097168 , n28171 );
buf ( R_2a7_1d9fc348 , n28174 );
buf ( R_7f3_1e091448 , n28177 );
buf ( R_73c_1dfba188 , n28178 );
buf ( R_bd1_1e6b7fc8 , n28246 );
buf ( R_4a6_1dda0868 , C0 );
buf ( R_3dd_1d9d8568 , n28256 );
buf ( R_346_1d9d2c08 , C0 );
buf ( R_4c4_1dda1628 , n28257 );
buf ( R_b15_1e6b0a48 , n28363 );
buf ( R_5ec_1ddacf28 , n28364 );
buf ( R_bb4_1e6b6da8 , n28365 );
buf ( R_bed_1e6b9148 , n28467 );
buf ( R_7bf_1e08f3c8 , n28470 );
buf ( R_344_1d9d25c8 , n28471 );
buf ( R_c0b_1e6ba408 , n28474 );
buf ( R_6a5_1dfb4328 , n29040 );
buf ( R_b8c_1e6b54a8 , n29041 );
buf ( R_3a1_1d9d5fe8 , n29050 );
buf ( R_7ea_1e09d928 , C0 );
buf ( R_46e_1dd9e568 , C0 );
buf ( R_8ee_1e09b628 , C0 );
buf ( R_697_1dfb3a68 , n29053 );
buf ( R_77f_1dfbcb68 , n29056 );
buf ( R_391_1d9d55e8 , n29063 );
buf ( R_746_1dfb6448 , C0 );
buf ( R_b3b_1e6b2208 , n29066 );
buf ( R_7f1_1e091308 , n29084 );
buf ( R_410_1d9da548 , n29085 );
buf ( R_700_1dfb7c08 , n29086 );
buf ( R_58f_1dda9508 , n29089 );
buf ( R_582_1dda91e8 , C0 );
buf ( R_793_1dfbd7e8 , n29092 );
buf ( R_847_1e0948c8 , n29095 );
buf ( R_95e_1e17fc88 , C0 );
buf ( R_560_1dda77a8 , n29096 );
buf ( R_9ca_1e184008 , C0 );
buf ( R_397_1d9d59a8 , n29099 );
buf ( R_46b_1d9dde28 , n29102 );
buf ( R_44e_1d9fc028 , C0 );
buf ( R_6cc_1dfb5b88 , n29103 );
buf ( R_62e_1dfafdc8 , C0 );
buf ( R_2b1_1d9fc988 , n29109 );
buf ( R_6f9_1dfb77a8 , n29116 );
buf ( R_af5_1e6af648 , n29161 );
buf ( R_b81_1e6b4dc8 , n29182 );
buf ( R_427_1d9db3a8 , n29185 );
buf ( R_547_1dda6808 , n29188 );
buf ( R_c1d_1e6baf48 , n29238 );
buf ( R_a2c_1e187848 , n29239 );
buf ( R_355_1d9d3068 , n29301 );
buf ( R_857_1e0952c8 , n29304 );
buf ( R_413_1d9da728 , n29307 );
buf ( R_afa_1e6afe68 , C0 );
buf ( R_adc_1e6ae6a8 , n29308 );
buf ( R_5fc_1ddad928 , n29309 );
buf ( R_c24_1e6bb3a8 , n29310 );
buf ( R_421_1d9dafe8 , n29317 );
buf ( R_892_1e17e608 , C0 );
buf ( R_70b_1dfb82e8 , n29320 );
buf ( R_aad_1e18c8e8 , n29384 );
buf ( R_3ca_1d9d8108 , C0 );
buf ( R_7ac_1e08e7e8 , n29385 );
buf ( R_8da_1e09a9a8 , C0 );
buf ( R_400_1d9d9b48 , n29386 );
buf ( R_bb0_1e6b6b28 , n29387 );
buf ( R_893_1e097848 , n29390 );
buf ( R_902_1e09c2a8 , C0 );
buf ( R_a93_1e18b8a8 , n29393 );
buf ( R_8cd_1e099c88 , n29469 );
buf ( R_861_1e095908 , n29505 );
buf ( R_3ea_1d9d9288 , C0 );
buf ( R_915_1e09c988 , n29584 );
buf ( R_844_1e0946e8 , n29585 );
buf ( R_677_1dfb2668 , n29588 );
buf ( R_602_1dfae248 , C0 );
buf ( R_39c_1d9d5cc8 , n29589 );
buf ( R_be3_1e6b8b08 , n29592 );
buf ( R_bea_1e6b9468 , C0 );
buf ( R_993_1e1818a8 , n29595 );
buf ( R_bad_1e6b6948 , n29777 );
buf ( R_88d_1e097488 , n30186 );
buf ( R_5a2_1ddaa5e8 , C0 );
buf ( R_655_1dfb1128 , n30243 );
buf ( R_4ad_1dda07c8 , n30384 );
buf ( R_493_1dd9f788 , n30387 );
buf ( R_894_1e0978e8 , n30388 );
buf ( R_668_1dfb1d08 , n30389 );
buf ( R_730_1dfb9a08 , n30390 );
buf ( R_7dc_1e0905e8 , n30391 );
buf ( R_abd_1e18d2e8 , n30500 );
buf ( R_662_1dfb1e48 , C0 );
buf ( R_a7c_1e18aa48 , n30501 );
buf ( R_5cf_1ddabd08 , n30504 );
buf ( R_328_1d9d1448 , n30505 );
buf ( R_741_1dfba4a8 , n30512 );
buf ( R_9a6_1e182988 , C0 );
buf ( R_36d_1d9d3f68 , n30587 );
buf ( R_308_1d9d0048 , n30588 );
buf ( R_95b_1e17f5a8 , n30591 );
buf ( R_b63_1e6b3b08 , n30594 );
buf ( R_2da_1d9ce888 , C0 );
buf ( R_5dc_1ddac528 , n30595 );
buf ( R_49f_1dd9ff08 , n30598 );
buf ( R_895_1e097988 , n30654 );
buf ( R_761_1dfbb8a8 , n30673 );
buf ( R_2e4_1d9ce9c8 , n30674 );
buf ( R_ab5_1e18cde8 , n30753 );
buf ( R_c28_1e6bb628 , n30754 );
buf ( R_8d4_1e09a0e8 , n30755 );
buf ( R_a8c_1e18b448 , n30756 );
buf ( R_597_1dda9a08 , n30759 );
buf ( R_5c4_1ddab628 , n30760 );
buf ( R_384_1d9d4dc8 , n30761 );
buf ( R_31c_1d9d0cc8 , n30762 );
buf ( R_987_1e181128 , n30765 );
buf ( R_b2e_1e6b1ee8 , C0 );
buf ( R_2f3_1d9cf328 , n30768 );
buf ( R_6cf_1dfb5d68 , n30771 );
buf ( R_6e4_1dfb6a88 , n30772 );
buf ( R_357_1d9d31a8 , n30775 );
buf ( R_3c1_1d9d73e8 , n30781 );
buf ( R_5e7_1ddacc08 , n30784 );
buf ( R_974_1e180548 , n30785 );
buf ( R_61a_1dfaf148 , C0 );
buf ( R_3f8_1d9d9648 , n30786 );
buf ( R_802_1e0922a8 , C0 );
buf ( R_593_1dda9788 , n30789 );
buf ( R_a69_1e189e68 , n31000 );
buf ( R_a87_1e18b128 , n31003 );
buf ( R_a5d_1e1896e8 , n31018 );
buf ( R_a2b_1e1877a8 , n31021 );
buf ( R_671_1dfb22a8 , n31028 );
buf ( R_4cf_1dda1d08 , n31031 );
buf ( R_420_1d9daf48 , n31032 );
buf ( R_6bc_1dfb5188 , n31033 );
buf ( R_43f_1d9dc2a8 , n31036 );
buf ( R_692_1dfb3c48 , C0 );
buf ( R_80b_1e092348 , n31039 );
buf ( R_882_1e0972a8 , C0 );
buf ( R_871_1e096308 , n31127 );
buf ( R_2c2_1d9fd928 , C0 );
buf ( R_2ce_1d9cfa08 , C0 );
buf ( R_a9c_1e18be48 , n31128 );
buf ( R_768_1dfbbd08 , n31129 );
buf ( R_56d_1dda7fc8 , n31189 );
buf ( R_34c_1d9d2ac8 , n31190 );
buf ( R_b8f_1e6b5688 , n31193 );
buf ( R_b07_1e6b0188 , n31196 );
buf ( R_6b5_1dfb4d28 , n31282 );
buf ( R_5ae_1ddaad68 , C0 );
buf ( R_2df_1d9ce6a8 , n31285 );
buf ( R_674_1dfb2488 , n31286 );
buf ( R_608_1dfae108 , n31287 );
buf ( R_ad3_1e6ae108 , n31290 );
buf ( R_505_1dda3ec8 , n31361 );
buf ( R_8bf_1e0993c8 , n31364 );
buf ( R_542_1dda69e8 , C0 );
buf ( R_7f6_1e091b28 , C0 );
buf ( R_504_1dda3e28 , n31365 );
buf ( R_8a7_1e0984c8 , n31368 );
buf ( R_76a_1dfbc5c8 , C0 );
buf ( R_937_1e09dec8 , n31371 );
buf ( R_6fb_1dfb78e8 , n31374 );
buf ( R_3b0_1d9d6948 , n31375 );
buf ( R_2c0_1d9fd2e8 , n31376 );
buf ( R_37c_1d9d48c8 , n31377 );
buf ( R_782_1dfbd248 , C0 );
buf ( R_503_1dda3d88 , n31380 );
buf ( R_82e_1e093e28 , C0 );
buf ( R_8bb_1e099148 , n31383 );
buf ( R_430_1d9db948 , n31384 );
buf ( R_5cb_1ddaba88 , n31387 );
buf ( R_ae6_1e6af1e8 , C0 );
buf ( R_7a3_1e08e248 , n31390 );
buf ( R_b78_1e6b4828 , n31391 );
buf ( R_bc9_1e6b7ac8 , n31465 );
buf ( R_380_1d9d4b48 , n31466 );
buf ( R_33d_1d9d2168 , n31661 );
buf ( R_8e0_1e09a868 , n31662 );
buf ( R_3c7_1d9d77a8 , n31665 );
buf ( R_2b2_1d9fcf28 , C0 );
buf ( R_618_1dfaeb08 , n31666 );
buf ( R_823_1e093248 , n31669 );
buf ( R_89e_1e098428 , C0 );
buf ( R_502_1dda41e8 , C0 );
buf ( R_b6f_1e6b4288 , n31672 );
buf ( R_c00_1e6b9d28 , n31673 );
buf ( R_98d_1e1814e8 , n31679 );
buf ( R_28b_1d9fb1c8 , n31718 );
buf ( R_a55_1e1891e8 , n31738 );
buf ( R_3c4_1d9d75c8 , n31739 );
buf ( R_40c_1d9da2c8 , n31740 );
buf ( R_2d2_1d9ce388 , C0 );
buf ( R_c21_1e6bb1c8 , n31792 );
buf ( R_b3d_1e6b2348 , n32069 );
buf ( R_877_1e0966c8 , n32072 );
buf ( R_855_1e095188 , n32095 );
buf ( R_41d_1d9dad68 , n32100 );
buf ( R_438_1d9dbe48 , n32101 );
buf ( R_2d6_1d9ce608 , C0 );
buf ( R_7da_1e0909a8 , C0 );
buf ( R_6f6_1dfb7ac8 , C0 );
buf ( R_9aa_1e182e88 , C0 );
buf ( R_b47_1e6b2988 , n32104 );
buf ( R_a2a_1e6b3ce8 , C0 );
buf ( R_41f_1d9daea8 , n32107 );
buf ( R_ae4_1e6aeba8 , n32108 );
buf ( R_a79_1e18a868 , n32127 );
buf ( R_3a3_1d9d6128 , n32130 );
buf ( R_5bd_1ddab1c8 , n32199 );
buf ( R_301_1d9cfbe8 , n32205 );
buf ( R_298_1d9fb9e8 , n32213 );
buf ( R_bb9_1e6b70c8 , n32233 );
buf ( R_82d_1e093888 , n32256 );
buf ( R_404_1d9d9dc8 , n32257 );
buf ( R_a62_1e189f08 , C0 );
buf ( R_93c_1e17e248 , n32258 );
buf ( R_62d_1dfaf828 , n32264 );
buf ( R_579_1dda8748 , n32334 );
buf ( R_452_1ddac3e8 , C0 );
buf ( R_54d_1dda6bc8 , n32352 );
buf ( R_4d9_1dda2348 , n32414 );
buf ( R_4d4_1dda2028 , n32415 );
buf ( R_6c1_1dfb54a8 , n32578 );
buf ( R_379_1d9d46e8 , n32583 );
buf ( R_34e_1d9d3108 , C0 );
buf ( R_94a_1e097ca8 , C0 );
buf ( R_74b_1dfbaae8 , n32586 );
buf ( R_ade_1e6aece8 , C0 );
buf ( R_79f_1e08dfc8 , n32589 );
buf ( R_797_1dfbda68 , n32592 );
buf ( R_943_1e17e6a8 , n32595 );
buf ( R_653_1dfb0fe8 , n32598 );
buf ( R_3d8_1d9d8248 , n32599 );
buf ( R_b61_1e6b39c8 , n32614 );
buf ( R_bc4_1e6b77a8 , n32615 );
buf ( R_a02_1e186308 , C0 );
buf ( R_368_1d9d3c48 , n32616 );
buf ( R_35e_1d9d3b08 , C0 );
buf ( R_7fe_1e092028 , C0 );
buf ( R_499_1dd9fb48 , n32704 );
buf ( R_680_1dfb2c08 , n32705 );
buf ( R_2a8_1d9fc3e8 , n32706 );
buf ( R_6ec_1dfb6f88 , n32707 );
buf ( R_776_1dfbcac8 , C0 );
buf ( R_b5e_1e6b0368 , C0 );
buf ( R_635_1dfafd28 , n32713 );
buf ( R_7fa_1e091da8 , C0 );
buf ( R_af7_1e6af788 , n32716 );
buf ( R_8c4_1e0996e8 , n32717 );
buf ( R_408_1d9da048 , n32718 );
buf ( R_ab9_1e18d068 , n32733 );
buf ( R_6a2_1dfb61c8 , C0 );
buf ( R_291_1d9fb588 , n32744 );
buf ( R_7b8_1e08ef68 , n32745 );
buf ( R_8b6_1e08e6a8 , C0 );
buf ( R_48a_1dda0d68 , C0 );
buf ( R_6c7_1dfb5868 , n32748 );
buf ( R_c10_1e6ba728 , n32749 );
buf ( R_bf1_1e6b93c8 , n32765 );
buf ( R_4d6_1dd9e2e8 , C0 );
buf ( R_5b3_1ddaab88 , n32768 );
buf ( R_771_1dfbc2a8 , n32789 );
buf ( R_af1_1e6af3c8 , n32840 );
buf ( R_6e1_1dfb68a8 , n32846 );
buf ( R_a9f_1e18c028 , n32849 );
buf ( R_b17_1e6b0b88 , n32852 );
buf ( R_b30_1e6b1b28 , n32853 );
buf ( R_bde_1e6b37e8 , C0 );
buf ( R_998_1e181bc8 , n32854 );
buf ( R_a4a_1e189008 , C0 );
buf ( R_48e_1dd9f968 , C0 );
buf ( R_688_1dfb3108 , n32855 );
buf ( R_810_1e092668 , n32856 );
buf ( R_75c_1dfbb588 , n32857 );
buf ( R_3bb_1d9d7028 , n32860 );
buf ( R_c2e_1e17f008 , C0 );
buf ( R_5d2_1d9db308 , C0 );
buf ( R_32e_1d9d1d08 , C0 );
buf ( R_580_1dda8ba8 , n32861 );
buf ( R_453_1d9dcf28 , n32864 );
buf ( R_83a_1e0913a8 , C0 );
buf ( R_41e_1d9dc988 , C0 );
buf ( R_97c_1e180a48 , n32865 );
buf ( R_5b8_1ddaaea8 , n32866 );
buf ( R_363_1d9d3928 , n32869 );
buf ( R_94e_1ddadce8 , C0 );
buf ( R_7c4_1e08f6e8 , n32870 );
buf ( R_52c_1dda5728 , n32871 );
buf ( R_aa2_1e18c708 , C0 );
buf ( R_625_1dfaf328 , n32880 );
buf ( R_4b7_1dda0e08 , n32883 );
buf ( R_55d_1dda75c8 , n32899 );
buf ( R_b0e_1e6b0ae8 , C0 );
buf ( R_425_1d9db268 , n32919 );
buf ( R_30c_1d9d02c8 , n32920 );
buf ( R_3db_1d9d8428 , n32923 );
buf ( R_a48_1e1889c8 , n32924 );
buf ( R_aaf_1e18ca28 , n32927 );
buf ( R_5ad_1ddaa7c8 , n32979 );
buf ( R_589_1dda9148 , n33052 );
buf ( R_338_1d9d1e48 , n33053 );
buf ( R_832_1e0940a8 , C0 );
buf ( R_790_1dfbd608 , n33054 );
buf ( R_318_1d9d0a48 , n33055 );
buf ( R_869_1e095e08 , n33148 );
buf ( R_6d3_1dfb5fe8 , n33151 );
buf ( R_60c_1dfae388 , n33152 );
buf ( R_56a_1dda82e8 , C0 );
buf ( R_887_1e0970c8 , n33155 );
buf ( R_815_1e092988 , n33169 );
buf ( R_66b_1dfb1ee8 , n33172 );
buf ( R_a34_1e187d48 , n33173 );
buf ( R_40f_1d9da4a8 , n33176 );
buf ( R_ac3_1e18d6a8 , n33179 );
buf ( R_324_1d9d11c8 , n33180 );
buf ( R_614_1dfae888 , n33181 );
buf ( R_752_1dfbb448 , C0 );
buf ( R_4c0_1dda13a8 , n33182 );
buf ( R_7d9_1e090408 , n33201 );
buf ( R_ad0_1e18dec8 , n33202 );
buf ( R_bee_1e6b96e8 , C0 );
buf ( R_736_1dfba2c8 , C0 );
buf ( R_727_1dfb9468 , n33205 );
buf ( R_a8a_1e18b808 , C0 );
buf ( R_933_1e09dc48 , n33208 );
buf ( R_8b1_1e098b08 , n33279 );
buf ( R_606_1dfae4c8 , C0 );
buf ( R_927_1e09d4c8 , n33282 );
buf ( R_a7a_1e18ae08 , C0 );
buf ( R_333_1d9d1b28 , n33285 );
buf ( R_968_1e17fdc8 , n33286 );
buf ( R_574_1dda8428 , n33287 );
buf ( R_836_1e094328 , C0 );
buf ( R_757_1dfbb268 , n33290 );
buf ( R_2db_1d9ce428 , n33293 );
buf ( R_af4_1e6af5a8 , n33294 );
buf ( R_454_1d9dcfc8 , n33295 );
buf ( R_412_1d9dab88 , C0 );
buf ( R_709_1dfb81a8 , n33303 );
buf ( R_8a4_1e0982e8 , n33304 );
buf ( R_c1b_1e6bae08 , n33307 );
buf ( R_846_1e094d28 , C0 );
buf ( R_3ff_1d9d9aa8 , n33310 );
buf ( R_76e_1dfbdec8 , C0 );
buf ( R_33f_1d9d22a8 , n33313 );
buf ( R_4af_1dda0908 , n33316 );
buf ( R_a67_1e189d28 , n33319 );
buf ( R_616_1dfaeec8 , C0 );
buf ( R_b49_1e6b2ac8 , n33507 );
buf ( R_2f4_1d9cf3c8 , n33508 );
buf ( R_426_1d9db808 , C0 );
buf ( R_2e5_1d9cea68 , n33516 );
buf ( R_bb5_1e6b6e48 , n33532 );
buf ( R_7b6_1e08f328 , C0 );
buf ( R_751_1dfbaea8 , n33550 );
buf ( R_bd0_1e6b7f28 , n33551 );
buf ( R_610_1dfae608 , n33552 );
buf ( R_918_1e09cb68 , n33553 );
buf ( R_35c_1d9d34c8 , n33554 );
buf ( R_924_1e09d2e8 , n33555 );
buf ( R_912_1e09cca8 , C0 );
buf ( R_77d_1dfbca28 , n33560 );
buf ( R_774_1dfbc488 , n33561 );
buf ( R_a71_1e18a368 , n33633 );
buf ( R_32d_1d9d1768 , n33705 );
buf ( R_99d_1e181ee8 , n33711 );
buf ( R_87d_1e096a88 , n33778 );
buf ( R_472_1dd9e7e8 , C0 );
buf ( R_b2a_1e6b1c68 , C0 );
buf ( R_56f_1dda8108 , n33781 );
buf ( R_b87_1e6b5188 , n33784 );
buf ( R_921_1e09d108 , n33847 );
buf ( R_375_1d9d4468 , n33852 );
buf ( R_576_1dda8ce8 , C0 );
buf ( R_b82_1e6b5368 , C0 );
buf ( R_39e_1d9d6308 , C0 );
buf ( R_856_1e095728 , C0 );
buf ( R_6c2_1dfb5a48 , C0 );
buf ( R_2c3_1d9fd4c8 , n33855 );
buf ( R_90b_1e09c348 , n33858 );
buf ( R_92f_1e09d9c8 , n33861 );
buf ( R_38e_1d9d5908 , C0 );
buf ( R_b9e_1e18d388 , C0 );
buf ( R_8cc_1e099be8 , n33862 );
buf ( R_860_1e095868 , n33863 );
buf ( R_c09_1e6ba2c8 , n33873 );
buf ( R_b09_1e6b02c8 , n33888 );
buf ( R_521_1dda5048 , n33977 );
buf ( R_b4a_1e6b3068 , C0 );
buf ( R_88c_1e0973e8 , n33978 );
buf ( R_520_1dda4fa8 , n33979 );
buf ( R_8b5_1e098d88 , n34040 );
buf ( R_b5d_1e6b3748 , n34084 );
buf ( R_843_1e094648 , n34087 );
buf ( R_633_1dfafbe8 , n34090 );
buf ( R_7c2_1e08faa8 , C0 );
buf ( R_6d8_1dfb6308 , n34091 );
buf ( R_38d_1d9d5368 , n34098 );
buf ( R_7e7_1e090cc8 , n34101 );
buf ( R_bfc_1e6b9aa8 , n34102 );
buf ( R_841_1e094508 , n34116 );
buf ( R_a96_1e18bf88 , C0 );
buf ( R_7e5_1e090b88 , n34267 );
buf ( R_51f_1dda4f08 , n34270 );
buf ( R_949_1e17ea68 , n34289 );
buf ( R_b5a_1e6b3a68 , C0 );
buf ( R_2e0_1d9ce748 , n34290 );
buf ( R_acd_1e18dce8 , n34296 );
buf ( R_70f_1dfb8568 , n34299 );
buf ( R_c15_1e6baa48 , n34321 );
buf ( R_310_1d9d0548 , n34322 );
buf ( R_bf5_1e6b9648 , n34395 );
buf ( R_314_1d9d07c8 , n34396 );
buf ( R_6af_1dfb4968 , n34399 );
buf ( R_445_1d9dc668 , n34522 );
buf ( R_658_1dfb1308 , n34523 );
buf ( R_a6c_1e18a048 , n34524 );
buf ( R_2c1_1d9fd388 , n34533 );
buf ( R_2b3_1d9fcac8 , n34536 );
buf ( R_6de_1dfb6bc8 , C0 );
buf ( R_9b9_1e183068 , n34542 );
buf ( R_6ad_1dfb4828 , n34621 );
buf ( R_548_1dda68a8 , n34622 );
buf ( R_4c9_1dda1948 , n34679 );
buf ( R_51e_1dda5368 , C0 );
buf ( R_96a_1e180408 , C0 );
buf ( R_455_1d9dd068 , n34743 );
buf ( R_8d3_1e09a048 , n34746 );
buf ( R_bb1_1e6b6bc8 , n34751 );
buf ( R_7d7_1e0902c8 , n34754 );
buf ( R_6a0_1dfb4008 , n34755 );
buf ( R_b79_1e6b48c8 , n34856 );
buf ( R_565_1dda7ac8 , n34936 );
buf ( R_586_1dda9468 , C0 );
buf ( R_4a7_1dda0408 , n34939 );
buf ( R_b70_1e6b4328 , n34940 );
buf ( R_661_1dfb18a8 , n34946 );
buf ( R_2d3_1d9fdec8 , n34949 );
buf ( R_ad9_1e6ae4c8 , n35056 );
buf ( R_a85_1e18afe8 , n35077 );
buf ( R_a77_1e18a728 , n35080 );
buf ( R_2d7_1d9ce1a8 , n35083 );
buf ( R_7b3_1e08ec48 , n35086 );
buf ( R_870_1e096268 , n35087 );
buf ( R_43e_1d9dc708 , C0 );
buf ( R_6db_1dfb64e8 , n35090 );
buf ( R_807_1e0920c8 , n35093 );
buf ( R_a74_1e18a548 , n35094 );
buf ( R_bf9_1e6b98c8 , n35107 );
buf ( R_321_1d9d0fe8 , n35114 );
buf ( R_a53_1e1890a8 , n35117 );
buf ( R_4e3_1dda2988 , n35120 );
buf ( R_831_1e093b08 , n35196 );
buf ( R_66e_1dfb25c8 , C0 );
buf ( R_ac6_1e18dd88 , C0 );
buf ( R_55a_1dda78e8 , C0 );
buf ( R_4c6_1dda1c68 , C0 );
buf ( R_4e4_1dda2a28 , n35197 );
buf ( R_4e2_1dda2de8 , C0 );
buf ( R_c22_1e6b55e8 , C0 );
buf ( R_92c_1e09d7e8 , n35198 );
buf ( R_7c9_1e08fa08 , n35217 );
buf ( R_623_1dfaf1e8 , n35220 );
buf ( R_b58_1e6b3428 , n35221 );
buf ( R_370_1d9d4148 , n35222 );
buf ( R_3be_1d9d7708 , C0 );
buf ( R_4e5_1dda2ac8 , n35238 );
buf ( R_a03_1e185ea8 , n35241 );
buf ( R_c12_1e6bad68 , C0 );
buf ( R_456_1d9dd608 , C0 );
buf ( R_bf2_1e6b9968 , C0 );
buf ( R_6a7_1dfb4468 , n35244 );
buf ( R_c30_1e6bbb28 , n35245 );
buf ( R_40b_1d9da228 , n35248 );
buf ( R_42f_1d9db8a8 , n35251 );
buf ( R_68d_1dfb3428 , n35393 );
buf ( R_735_1dfb9d28 , n35399 );
buf ( R_78d_1dfbd428 , n35478 );
buf ( R_8df_1e09a7c8 , n35481 );
buf ( R_41c_1d9dacc8 , n35482 );
buf ( R_46f_1dd9e108 , n35485 );
buf ( R_2a9_1d9fc488 , n35492 );
buf ( R_81e_1e093428 , C0 );
buf ( R_5e0_1ddac7a8 , n35493 );
buf ( R_462_1d9ddd88 , C0 );
buf ( R_60a_1dfae748 , C0 );
buf ( R_5a7_1ddaa408 , n35496 );
buf ( R_403_1d9d9d28 , n35499 );
buf ( R_2c6_1d9fdba8 , C0 );
buf ( R_7e3_1e090a48 , n35502 );
buf ( R_7ee_1e09c528 , C0 );
buf ( R_706_1dfb84c8 , C0 );
buf ( R_c17_1e6bab88 , n35505 );
buf ( R_c1f_1e6bb088 , n35508 );
buf ( R_b93_1e6b5908 , n35511 );
buf ( R_854_1e0950e8 , n35512 );
buf ( R_b9f_1e6b6088 , n35515 );
buf ( R_8e5_1e09ab88 , n35520 );
buf ( R_437_1d9dbda8 , n35523 );
buf ( R_612_1dfaec48 , C0 );
buf ( R_816_1e0931a8 , C0 );
buf ( R_b19_1e6b0cc8 , n35536 );
buf ( R_73b_1dfba0e8 , n35539 );
buf ( R_a44_1e188748 , n35540 );
buf ( R_93e_1e17e888 , C0 );
buf ( R_67c_1dfb2988 , n35541 );
buf ( R_992_1e181d08 , C0 );
buf ( R_494_1dd9f828 , n35542 );
buf ( R_3e0_1d9d8748 , n35543 );
buf ( R_7a7_1e08e4c8 , n35546 );
buf ( R_876_1e096b28 , C0 );
buf ( R_543_1dda6588 , n35549 );
buf ( R_8ae_1dfbc0c8 , C0 );
buf ( R_351_1d9d2de8 , n35572 );
buf ( R_457_1d9dd1a8 , n35575 );
buf ( R_bf6_1e6b3f68 , C0 );
buf ( R_a38_1e187fc8 , n35576 );
buf ( R_6f1_1dfb72a8 , n35581 );
buf ( R_b3e_1e6b28e8 , C0 );
buf ( R_53e_1dda6768 , C0 );
buf ( R_ac0_1e18d4c8 , n35582 );
buf ( R_763_1dfbb9e8 , n35585 );
buf ( R_c26_1e6b8ce8 , C0 );
buf ( R_650_1dfb0e08 , n35586 );
buf ( R_361_1d9d37e8 , n35646 );
buf ( R_aaa_1e187e88 , C0 );
buf ( R_b10_1e6b0728 , n35647 );
buf ( R_b2c_1e6b18a8 , n35648 );
buf ( R_5a1_1ddaa048 , n35668 );
buf ( R_be7_1e6b8d88 , n35671 );
buf ( R_b26_1e6b19e8 , C0 );
buf ( R_4a0_1dd9ffa8 , n35672 );
buf ( R_95a_1e17fa08 , C0 );
buf ( R_909_1e09c208 , n35723 );
buf ( R_463_1d9dd928 , n35726 );
buf ( R_407_1d9d9fa8 , n35729 );
buf ( R_5c5_1ddab6c8 , n35731 );
buf ( R_986_1e181588 , C0 );
buf ( R_515_1dda48c8 , n35748 );
buf ( R_5c1_1ddab448 , n35766 );
buf ( R_297_1d9fb948 , n35775 );
buf ( R_514_1dda4828 , n35776 );
buf ( R_b4c_1e6b2ca8 , n35777 );
buf ( R_973_1e1804a8 , n35780 );
buf ( R_60e_1dfae9c8 , C0 );
buf ( R_7d4_1e0900e8 , n35781 );
buf ( R_7c7_1e08f8c8 , n35784 );
buf ( R_513_1dda4788 , n35787 );
buf ( R_65f_1dfb1768 , n35790 );
buf ( R_9b5_1e182de8 , n35796 );
buf ( R_2ee_1d9cf508 , C0 );
buf ( R_91b_1e09cd48 , n35799 );
buf ( R_af6_1e6afbe8 , C0 );
buf ( R_83d_1e094288 , n35868 );
buf ( R_8c3_1e099648 , n35871 );
buf ( R_458_1d9dd248 , n35872 );
buf ( R_512_1dda4be8 , C0 );
buf ( R_ba6_1e6b69e8 , C0 );
buf ( R_5e5_1ddacac8 , n35891 );
buf ( R_57b_1dda8888 , n35894 );
buf ( R_aeb_1e6af008 , n35897 );
buf ( R_7f4_1e0914e8 , n35898 );
buf ( R_a46_1e188d88 , C0 );
buf ( R_b8d_1e6b5548 , n35913 );
buf ( R_562_1dda7de8 , C0 );
buf ( R_745_1dfba728 , n35918 );
buf ( R_557_1dda7208 , n35921 );
buf ( R_464_1d9dd9c8 , n35922 );
buf ( R_835_1e093d88 , n35938 );
buf ( R_49a_1dda00e8 , C0 );
buf ( R_7d1_1e08ff08 , n35943 );
buf ( R_911_1e09c708 , n35963 );
buf ( R_6e9_1dfb6da8 , n35970 );
buf ( R_723_1dfb91e8 , n35973 );
buf ( R_a95_1e18b9e8 , n35979 );
buf ( R_58d_1dda93c8 , n35997 );
buf ( R_a89_1e18b268 , n36003 );
buf ( R_780_1dfbcc08 , n36004 );
buf ( R_740_1dfba408 , n36005 );
buf ( R_72f_1dfb9968 , n36008 );
buf ( R_828_1e093568 , n36009 );
buf ( R_89c_1e097de8 , n36010 );
buf ( R_a32_1e188108 , C0 );
buf ( R_840_1e094468 , n36011 );
buf ( R_b37_1e6b1f88 , n36014 );
buf ( R_9db_1e1845a8 , n36017 );
buf ( R_b22_1e6b1768 , C0 );
buf ( R_9dc_1e184648 , n36018 );
buf ( R_9da_1e184a08 , C0 );
buf ( R_794_1dfbd888 , n36019 );
buf ( R_33a_1d9d2488 , C0 );
buf ( R_424_1d9db1c8 , n36020 );
buf ( R_2dc_1d9ce4c8 , n36021 );
buf ( R_a6f_1e18a228 , n36024 );
buf ( R_98c_1e181448 , n36025 );
buf ( R_6b6_1dfb52c8 , C0 );
buf ( R_908_1e09c168 , n36026 );
buf ( R_9dd_1e1846e8 , n36482 );
buf ( R_965_1e17fbe8 , n36489 );
buf ( R_28a_1d9fb128 , n36514 );
buf ( R_529_1dda5548 , n36526 );
buf ( R_40e_1d9da908 , C0 );
buf ( R_bcd_1e6b7d48 , n36541 );
buf ( R_476_1dd9ea68 , C0 );
buf ( R_393_1d9d5728 , n36544 );
buf ( R_a40_1e1884c8 , n36545 );
buf ( R_528_1dda54a8 , n36546 );
buf ( R_2fa_1d9d0188 , C0 );
buf ( R_a3c_1e188248 , n36547 );
buf ( R_868_1e095d68 , n36548 );
buf ( R_2cf_1d9fdc48 , n36551 );
buf ( R_2c4_1d9fd568 , n36552 );
buf ( R_7cc_1e08fbe8 , n36553 );
buf ( R_8fd_1e09ba88 , n36558 );
buf ( R_3d5_1d9d8068 , n36564 );
buf ( R_b64_1e6b3ba8 , n36565 );
buf ( R_527_1dda5408 , n36568 );
buf ( R_9d1_1e183f68 , n36575 );
buf ( R_46c_1d9ddec8 , n36576 );
buf ( R_2f5_1d9cf468 , n36582 );
buf ( R_839_1e094008 , n36602 );
buf ( R_554_1dda7028 , n36603 );
buf ( R_3ab_1d9d6628 , n36606 );
buf ( R_459_1d9dd2e8 , n36611 );
buf ( R_b4f_1e6b2e88 , n36614 );
buf ( R_886_1e097528 , C0 );
buf ( R_3e5_1d9d8a68 , n36620 );
buf ( R_52d_1dda57c8 , n36670 );
buf ( R_290_1d9fb4e8 , n36680 );
buf ( R_b7a_1e18cc08 , C0 );
buf ( R_526_1dda5ae8 , C0 );
buf ( R_79a_1e098e28 , C0 );
buf ( R_ba0_1e6b6128 , n36681 );
buf ( R_6d1_1dfb5ea8 , n36686 );
buf ( R_713_1dfb87e8 , n36689 );
buf ( R_685_1dfb2f28 , n36832 );
buf ( R_3fe_1d9d9f08 , C0 );
buf ( R_638_1dfaff08 , n36833 );
buf ( R_465_1d9dda68 , n36847 );
buf ( R_b91_1e6b57c8 , n36849 );
buf ( R_b53_1e6b3108 , n36852 );
buf ( R_8ad_1e098888 , n36857 );
buf ( R_59e_1dd9e068 , C0 );
buf ( R_9c5_1e1837e8 , n36865 );
buf ( R_3a9_1d9d64e8 , n36871 );
buf ( R_3b3_1d9d6b28 , n36874 );
buf ( R_2b4_1d9fcb68 , n36875 );
buf ( R_af3_1e6af508 , n36878 );
buf ( R_4f9_1dda3748 , n36896 );
buf ( R_a90_1e18b6c8 , n36897 );
buf ( R_389_1d9d50e8 , n36903 );
buf ( R_a6a_1e18a408 , C0 );
buf ( R_b1b_1e6b0e08 , n36906 );
buf ( R_4f8_1dda36a8 , n36907 );
buf ( R_b66_1e6b9be8 , C0 );
buf ( R_9d0_1e183ec8 , n36908 );
buf ( R_2e1_1d9ce7e8 , n36914 );
buf ( R_7d2_1e0904a8 , C0 );
buf ( R_803_1e091e48 , n36917 );
buf ( R_91e_1e09d428 , C0 );
buf ( R_4f7_1dda3608 , n36920 );
buf ( R_ab4_1e18cd48 , n36921 );
buf ( R_6ee_1dfb75c8 , C0 );
buf ( R_c05_1e6ba048 , n36936 );
buf ( R_704_1dfb7e88 , n36937 );
buf ( R_353_1d9d2f28 , n36940 );
buf ( R_ba7_1e6b6588 , n36943 );
buf ( R_87c_1e0969e8 , n36944 );
buf ( R_3f5_1d9d9468 , n36950 );
buf ( R_abc_1e18d248 , n36951 );
buf ( R_a83_1e18aea8 , n36954 );
buf ( R_b40_1e6b2528 , n36955 );
buf ( R_a06_1e186588 , C0 );
buf ( R_907_1e09c0c8 , n36958 );
buf ( R_664_1dfb1a88 , n36959 );
buf ( R_b71_1e6b43c8 , n36974 );
buf ( R_4f6_1ddad2e8 , C0 );
buf ( R_8b9_1e099008 , n36991 );
buf ( R_971_1e180368 , n36998 );
buf ( R_64e_1dfb11c8 , C0 );
buf ( R_679_1dfb27a8 , n37005 );
buf ( R_80c_1e0923e8 , n37006 );
buf ( R_347_1d9d27a8 , n37009 );
buf ( R_b28_1e6b1628 , n37010 );
buf ( R_7cf_1e08fdc8 , n37013 );
buf ( R_8fc_1e09b9e8 , n37014 );
buf ( R_72d_1dfb9828 , n37020 );
buf ( R_9c4_1e183748 , n37021 );
buf ( R_997_1e181b28 , n37024 );
buf ( R_85f_1e0957c8 , n37027 );
buf ( R_2d4_1d9cdfc8 , n37028 );
buf ( R_48f_1dd9f508 , n37031 );
buf ( R_adb_1e6ae608 , n37034 );
buf ( R_3b9_1d9d6ee8 , n37040 );
buf ( R_a51_1e188f68 , n37095 );
buf ( R_8cb_1e099b48 , n37098 );
buf ( R_2d8_1d9ce248 , n37099 );
buf ( R_a72_1e18a908 , C0 );
buf ( R_7f7_1e0916c8 , n37102 );
buf ( R_4b5_1dda0cc8 , n37121 );
buf ( R_88b_1e097348 , n37124 );
buf ( R_aa7_1e18c528 , n37127 );
buf ( R_699_1dfb3ba8 , n37267 );
buf ( R_68a_1dfb3748 , C0 );
buf ( R_9cf_1e183e28 , n37270 );
buf ( R_345_1d9d2668 , n37431 );
buf ( R_76b_1dfbbee8 , n37434 );
buf ( R_7aa_1e099328 , C0 );
buf ( R_5e9_1ddacd48 , n37452 );
buf ( R_a04_1e185f48 , n37453 );
buf ( R_36b_1d9d3e28 , n37456 );
buf ( R_444_1d9dc5c8 , n37457 );
buf ( R_842_1e094aa8 , C0 );
buf ( R_58a_1dda96e8 , C0 );
buf ( R_97b_1e1809a8 , n37460 );
buf ( R_5bc_1ddab128 , n37461 );
buf ( R_ae9_1e6aeec8 , n37468 );
buf ( R_74e_1dfbc348 , C0 );
buf ( R_69b_1dfb3ce8 , n37471 );
buf ( R_783_1dfbcde8 , n37474 );
buf ( R_64d_1dfb0c28 , n37482 );
buf ( R_938_1e17dfc8 , n37483 );
buf ( R_7bd_1e08f288 , n37502 );
buf ( R_7ca_1e08ffa8 , C0 );
buf ( R_482_1ddac668 , C0 );
buf ( R_2c7_1d9fd748 , n37505 );
buf ( R_621_1dfaf0a8 , n37511 );
buf ( R_9c3_1e1836a8 , n37514 );
buf ( R_309_1d9d00e8 , n37522 );
buf ( R_5f1_1ddad248 , n37539 );
buf ( R_4b8_1dda0ea8 , n37540 );
buf ( R_bcf_1e6b7e88 , n37543 );
buf ( R_824_1e0932e8 , n37544 );
buf ( R_6e6_1dfb70c8 , C0 );
buf ( R_7a4_1e08e2e8 , n37545 );
buf ( R_59d_1dda9dc8 , n37561 );
buf ( R_769_1dfbbda8 , n37651 );
buf ( R_38a_1d9d5688 , C0 );
buf ( R_4cb_1dda1a88 , n37654 );
buf ( R_8d9_1e09a408 , n37659 );
buf ( R_8d2_1e09a4a8 , C0 );
buf ( R_b24_1e6b13a8 , n37660 );
buf ( R_4ba_1d9d9a08 , C0 );
buf ( R_bdd_1e6b8748 , n37679 );
buf ( R_398_1d9d5a48 , n37680 );
buf ( R_31d_1d9d0d68 , n37687 );
buf ( R_47a_1dd9ece8 , C0 );
buf ( R_2ca_1d9ce108 , C0 );
buf ( R_b03_1e6aff08 , n37690 );
buf ( R_2a0_1d9fbee8 , n37691 );
buf ( R_71f_1dfb8f68 , n37694 );
buf ( R_950_1e17eec8 , n37695 );
buf ( R_9ce_1e184288 , C0 );
buf ( R_aae_1e6b6c68 , C0 );
buf ( R_b39_1e6b20c8 , n37710 );
buf ( R_906_1e090ea8 , C0 );
buf ( R_786_1dfbd4c8 , C0 );
buf ( R_81c_1e092de8 , n37711 );
buf ( R_94b_1e17eba8 , n37714 );
buf ( R_8fb_1e09b948 , n37717 );
buf ( R_3cb_1d9d7a28 , n37720 );
buf ( R_86f_1e0961c8 , n37723 );
buf ( R_584_1dda8e28 , n37724 );
buf ( R_40a_1d9da688 , C0 );
buf ( R_954_1e17f148 , n37725 );
buf ( R_944_1e17e748 , n37726 );
buf ( R_bc8_1e6b7a28 , n37727 );
buf ( R_9a1_1e182168 , n37733 );
buf ( R_c02_1e6ba5e8 , C0 );
buf ( R_967_1e17fd28 , n37736 );
buf ( R_7ff_1e091bc8 , n37739 );
buf ( R_329_1d9d14e8 , n37790 );
buf ( R_ba1_1e6b61c8 , n37803 );
buf ( R_717_1dfb8a68 , n37806 );
buf ( R_aa1_1e18c168 , n37812 );
buf ( R_591_1dda9648 , n37826 );
buf ( R_99c_1e181e48 , n37827 );
buf ( R_a42_1e188b08 , C0 );
buf ( R_ba8_1e6b6628 , n37828 );
buf ( R_ae1_1e6ae9c8 , n37841 );
buf ( R_9c2_1e183b08 , C0 );
buf ( R_6bb_1dfb50e8 , n37844 );
buf ( R_41b_1d9dac28 , n37847 );
buf ( R_93d_1e17e2e8 , n37858 );
buf ( R_5b2_1ddaafe8 , C0 );
buf ( R_5d6_1d9dd388 , C0 );
buf ( R_402_1d9da188 , C0 );
buf ( R_4b0_1dda09a8 , n37859 );
buf ( R_549_1dda6948 , n37941 );
buf ( R_53a_1dda64e8 , C0 );
buf ( R_70d_1dfb8428 , n37947 );
buf ( R_aa4_1e18c348 , n37948 );
buf ( R_798_1dfbdb08 , n37949 );
buf ( R_7fb_1e091948 , n37952 );
buf ( R_32a_1d9d1a88 , C0 );
buf ( R_a36_1e188388 , C0 );
buf ( R_5ed_1ddacfc8 , n37969 );
buf ( R_b9a_1e6b6268 , C0 );
buf ( R_c07_1e6ba188 , n37972 );
buf ( R_47e_1dd9ef68 , C0 );
buf ( R_ad2_1e6ae568 , C0 );
buf ( R_39d_1d9d5d68 , n37978 );
buf ( R_83f_1e0943c8 , n37981 );
buf ( R_7eb_1e090f48 , n37984 );
buf ( R_42e_1d9dbd08 , C0 );
buf ( R_b51_1e6b2fc8 , n37993 );
buf ( R_6b4_1dfb4c88 , n37994 );
buf ( R_694_1dfb3888 , n37995 );
buf ( R_68f_1dfb3568 , n37998 );
buf ( R_777_1dfbc668 , n38001 );
buf ( R_7b0_1e08ea68 , n38002 );
buf ( R_7a0_1e08e068 , n38003 );
buf ( R_75e_1dfbbbc8 , C0 );
buf ( R_5b7_1ddaae08 , n38006 );
buf ( R_63d_1dfb0228 , n38014 );
buf ( R_636_1dfb02c8 , C0 );
buf ( R_8de_1e09ac28 , C0 );
buf ( R_2ef_1d9cf0a8 , n38017 );
buf ( R_302_1d9d4508 , C0 );
buf ( R_9b8_1e182fc8 , n38018 );
buf ( R_4b2_1dda14e8 , C0 );
buf ( R_8e4_1e09aae8 , n38019 );
buf ( R_3de_1d9d8b08 , C0 );
buf ( R_ab8_1e18cfc8 , n38020 );
buf ( R_71b_1dfb8ce8 , n38023 );
buf ( R_c0c_1e6ba4a8 , n38024 );
buf ( R_c2b_1e6bb808 , n38028 );
buf ( R_5ac_1ddaa728 , n38029 );
buf ( R_853_1e095048 , n38032 );
buf ( R_2aa_1d9fca28 , C0 );
buf ( R_385_1d9d4e68 , n38038 );
buf ( R_436_1d9dc208 , C0 );
buf ( R_a60_1e1898c8 , n38039 );
buf ( R_7bb_1e08f148 , n38042 );
buf ( R_811_1e092708 , n38132 );
buf ( R_4c5_1dda16c8 , n38151 );
buf ( R_406_1d9da408 , C0 );
buf ( R_473_1dd9e388 , n38154 );
buf ( R_8aa_1e098ba8 , C0 );
buf ( R_b7e_1e6b50e8 , C0 );
buf ( R_7b5_1e08ed88 , n38159 );
buf ( R_5fb_1ddad888 , n38162 );
buf ( R_34d_1d9d2b68 , n38309 );
buf ( R_ae3_1e6aeb08 , n38312 );
buf ( R_6f3_1dfb73e8 , n38315 );
buf ( R_82b_1e093748 , n38318 );
buf ( R_72a_1dfbacc8 , C0 );
buf ( R_bc3_1e6b7708 , n38321 );
buf ( R_8fa_1e09bda8 , C0 );
buf ( R_567_1dda7c08 , n38324 );
buf ( R_89f_1e097fc8 , n38327 );
buf ( R_3ed_1d9d8f68 , n38333 );
buf ( R_599_1dda9b48 , n38351 );
buf ( R_851_1e094f08 , n38368 );
buf ( R_2dd_1d9ce568 , n38374 );
buf ( R_4a8_1dda04a8 , n38375 );
buf ( R_8a9_1e098608 , n38393 );
buf ( R_366_1d9d4008 , C0 );
buf ( R_376_1ddad568 , C0 );
buf ( R_75d_1dfbb628 , n38398 );
buf ( R_59a_1ddaa0e8 , C0 );
buf ( R_4c2_1dda19e8 , C0 );
buf ( R_8be_1e08eba8 , C0 );
buf ( R_2c5_1d9fd608 , n38404 );
buf ( R_595_1dda98c8 , n38418 );
buf ( R_446_1d9dd108 , C0 );
buf ( R_6c5_1dfb5728 , n38497 );
buf ( R_5d8_1ddac2a8 , n38498 );
buf ( R_682_1dfb3248 , C0 );
buf ( R_64b_1dfb0ae8 , n38501 );
buf ( R_791_1dfbd6a8 , n38520 );
buf ( R_b7b_1e6b4a08 , n38523 );
buf ( R_3b1_1d9d69e8 , n38529 );
buf ( R_7e9_1e090e08 , n38548 );
buf ( R_beb_1e6b9008 , n38551 );
buf ( R_6c0_1dfb5408 , n38552 );
buf ( R_8ba_1e0995a8 , C0 );
buf ( R_a8e_1e17f508 , C0 );
buf ( R_3c8_1d9d7848 , n38553 );
buf ( R_be4_1e6b8ba8 , n38554 );
buf ( R_544_1dda6628 , n38555 );
buf ( R_53f_1dda6308 , n38558 );
buf ( R_90e_1e09ca28 , C0 );
buf ( R_381_1d9d4be8 , n38564 );
buf ( R_a3e_1e188888 , C0 );
buf ( R_6fd_1dfb7a28 , n38572 );
buf ( R_a3a_1e188608 , C0 );
buf ( R_8c2_1e099aa8 , C0 );
buf ( R_af0_1e6af328 , n38573 );
buf ( R_296_1d9fb8a8 , n38586 );
buf ( R_b12_1e6b0d68 , C0 );
buf ( R_ba9_1e6b66c8 , n38594 );
buf ( R_b1d_1e6b0f48 , n38607 );
buf ( R_2b5_1d9fcc08 , n38613 );
buf ( R_6ff_1dfb7b68 , n38616 );
buf ( R_a98_1e18bbc8 , n38617 );
buf ( R_58e_1dda9968 , C0 );
buf ( R_753_1dfbafe8 , n38620 );
buf ( R_3c5_1d9d7668 , n38626 );
buf ( R_447_1d9dc7a8 , n38629 );
buf ( R_61f_1dfaef68 , n38632 );
buf ( R_54e_1dda28e8 , C0 );
buf ( R_6f8_1dfb7708 , n38633 );
buf ( R_3a4_1d9d61c8 , n38634 );
buf ( R_423_1d9db128 , n38637 );
buf ( R_6a4_1dfb4288 , n38638 );
buf ( R_b9b_1e6b5e08 , n38641 );
buf ( R_a07_1e186128 , n38644 );
buf ( R_55f_1dda7708 , n38647 );
buf ( R_79d_1dfbde28 , n38654 );
buf ( R_66d_1dfb2028 , n38661 );
buf ( R_5e2_1ddacde8 , C0 );
buf ( R_48b_1dd9f288 , n38664 );
buf ( R_5ee_1dda3a68 , C0 );
buf ( R_6c6_1dfb2d48 , C0 );
buf ( R_3e3_1d9d8928 , n38667 );
buf ( R_b83_1e6b4f08 , n38670 );
buf ( R_533_1dda5b88 , n38673 );
buf ( R_42d_1d9db768 , n38678 );
buf ( R_7e0_1e090868 , n38679 );
buf ( R_696_1dfb3ec8 , C0 );
buf ( R_3f9_1d9d96e8 , n38688 );
buf ( R_b88_1e6b5228 , n38689 );
buf ( R_758_1dfbb308 , n38690 );
buf ( R_3d2_1d9d8388 , C0 );
buf ( R_534_1dda5c28 , n38691 );
buf ( R_532_1d9d1308 , C0 );
buf ( R_867_1e095cc8 , n38694 );
buf ( R_2b6_1d9fd1a8 , C0 );
buf ( R_775_1dfbc528 , n38760 );
buf ( R_3e8_1d9d8c48 , n38761 );
buf ( R_4d0_1dda1da8 , n38762 );
buf ( R_30d_1d9d0368 , n38769 );
buf ( R_4e7_1dda2c08 , n38772 );
buf ( R_70a_1dfb8748 , C0 );
buf ( R_a58_1e1893c8 , n38773 );
buf ( R_4e8_1dda2ca8 , n38774 );
buf ( R_4e6_1dda3068 , C0 );
buf ( R_535_1dda5cc8 , n38860 );
buf ( R_5ea_1dda37e8 , C0 );
buf ( R_929_1e09d608 , n38876 );
buf ( R_448_1d9dc848 , n38877 );
buf ( R_b0b_1e6b0408 , n38880 );
buf ( R_319_1d9d0ae8 , n38887 );
buf ( R_985_1e180fe8 , n38895 );
buf ( R_32f_1d9d18a8 , n38898 );
buf ( R_4e9_1dda2d48 , n38910 );
buf ( R_b1f_1e6b1088 , n38913 );
buf ( R_495_1dd9f8c8 , n38933 );
buf ( R_63b_1dfb00e8 , n38936 );
buf ( R_536_1dda6268 , C0 );
buf ( R_3d9_1d9d82e8 , n38942 );
buf ( R_a4f_1e188e28 , n38945 );
buf ( R_470_1dd9e1a8 , n38946 );
buf ( R_2d5_1d9ce068 , n38952 );
buf ( R_3f0_1d9d9148 , n38953 );
buf ( R_acf_1e18de28 , n38956 );
buf ( R_ac2_1e18db08 , C0 );
buf ( R_9b4_1e182d48 , n38957 );
buf ( R_a05_1e185fe8 , n38991 );
buf ( R_2d9_1d9ce2e8 , n38997 );
buf ( R_8ed_1e09b088 , n39002 );
buf ( R_3f3_1d9d9328 , n39005 );
buf ( R_af2_1e6af968 , C0 );
buf ( R_44d_1d9dcb68 , n39011 );
buf ( R_645_1dfb0728 , n39019 );
buf ( R_648_1dfb0908 , n39020 );
buf ( R_4a1_1dda0048 , n39039 );
buf ( R_749_1dfba9a8 , n39045 );
buf ( R_2c8_1d9fd7e8 , n39046 );
buf ( R_3bc_1d9d70c8 , n39047 );
buf ( R_3f6_1ddad7e8 , C0 );
buf ( R_596_1dda9e68 , C0 );
buf ( R_c01_1e6b9dc8 , n39062 );
buf ( R_734_1dfb9c88 , n39063 );
buf ( R_5a5_1ddaa2c8 , n39075 );
buf ( R_6e3_1dfb69e8 , n39078 );
buf ( R_914_1e09c8e8 , n39079 );
buf ( R_43d_1d9dc168 , n39096 );
buf ( R_2cb_1d9fd9c8 , n39099 );
buf ( R_3d0_1d9d7d48 , n39100 );
buf ( R_b67_1e6b3d88 , n39103 );
buf ( R_b01_1e6afdc8 , n39108 );
buf ( R_37d_1d9d4968 , n39115 );
buf ( R_a80_1e18acc8 , n39116 );
buf ( R_9bd_1e1832e8 , n39123 );
buf ( R_339_1d9d1ee8 , n39185 );
buf ( R_7ad_1e08e888 , n39202 );
buf ( R_972_1e180908 , C0 );
buf ( R_a22_1e184788 , C0 );
buf ( R_486_1ddacb68 , C0 );
buf ( R_5d5_1ddac0c8 , n39207 );
buf ( R_592_1dda9be8 , C0 );
buf ( R_449_1d9dc8e8 , n39214 );
buf ( R_87b_1e096948 , n39217 );
buf ( R_8f5_1e09b588 , n39222 );
buf ( R_35a_1d9d3888 , C0 );
buf ( R_37a_1ddab9e8 , C0 );
buf ( R_991_1e181768 , n39228 );
buf ( R_62a_1dfb1448 , C0 );
buf ( R_808_1e092168 , n39229 );
buf ( R_3a6_1d9d6808 , C0 );
buf ( R_b95_1e6b5a48 , n39235 );
buf ( R_83e_1e17e108 , C0 );
buf ( R_386_1d9d5408 , C0 );
buf ( R_90d_1e09c488 , n39311 );
buf ( R_931_1e09db08 , n39334 );
buf ( R_ac9_1e18da68 , n39424 );
buf ( R_a31_1e187b68 , n39497 );
buf ( R_640_1dfb0408 , n39498 );
buf ( R_667_1dfb1c68 , n39501 );
buf ( R_6cb_1dfb5ae8 , n39504 );
buf ( R_74a_1e17f288 , C0 );
buf ( R_676_1dfb2ac8 , C0 );
buf ( R_372_1d9d4788 , C0 );
buf ( R_56c_1dda7f28 , n39505 );
buf ( R_334_1d9d1bc8 , n39506 );
buf ( R_31e_1d9fc528 , C0 );
buf ( R_981_1e180d68 , n39512 );
buf ( R_8ca_1e099fa8 , C0 );
buf ( R_85e_1e095c28 , C0 );
buf ( R_bbe_1e6af6e8 , C0 );
buf ( R_49b_1dd9fc88 , n39515 );
buf ( R_73a_1dfba548 , C0 );
buf ( R_5fe_1dfaf8c8 , C0 );
buf ( R_98b_1e1813a8 , n39518 );
buf ( R_88e_1e097a28 , C0 );
buf ( R_28f_1d9fb448 , n39528 );
buf ( R_9bc_1e183248 , n39529 );
buf ( R_5db_1ddac488 , n39532 );
buf ( R_88a_1e08ee28 , C0 );
buf ( R_5a6_1ddaa868 , C0 );
buf ( R_443_1d9dc528 , n39535 );
buf ( R_a0a_1e186808 , C0 );
buf ( R_358_1d9d3248 , n39536 );
buf ( R_88f_1e0975c8 , n39539 );
buf ( R_acc_1e18dc48 , n39540 );
buf ( R_aac_1e18c848 , n39541 );
buf ( R_2a2_1d9fde28 , C0 );
buf ( R_8a5_1e098388 , n39549 );
buf ( R_8ec_1e09afe8 , n39550 );
buf ( R_289_1d9fb088 , n39584 );
buf ( R_340_1d9d2348 , n39585 );
buf ( R_c2d_1e6bb948 , n39593 );
buf ( R_964_1e17fb48 , n39594 );
buf ( R_85d_1e095688 , n39608 );
buf ( R_6fa_1dfb7d48 , C0 );
buf ( R_4d5_1dda20c8 , n39613 );
buf ( R_a5a_1e18b308 , C0 );
buf ( R_7de_1e090c28 , C0 );
buf ( R_605_1ddadec8 , n39621 );
buf ( R_311_1d9d05e8 , n39628 );
buf ( R_8a6_1e098928 , C0 );
buf ( R_a2f_1e187a28 , n39631 );
buf ( R_81f_1e092fc8 , n39634 );
buf ( R_3b6_1d9d7208 , C0 );
buf ( R_315_1d9d0868 , n39641 );
buf ( R_93f_1e17e428 , n39644 );
buf ( R_5b1_1ddaaa48 , n39663 );
buf ( R_631_1dfafaa8 , n39669 );
buf ( R_890_1e097668 , n39670 );
buf ( R_670_1dfb2208 , n39671 );
buf ( R_b9c_1e6b5ea8 , n39672 );
buf ( R_8e9_1e09ae08 , n39691 );
buf ( R_932_1e093928 , C0 );
buf ( R_817_1e092ac8 , n39694 );
buf ( R_b60_1e6b3928 , n39695 );
buf ( R_979_1e180868 , n39703 );
buf ( R_8d8_1e09a368 , n39704 );
buf ( R_628_1dfaf508 , n39705 );
buf ( R_729_1dfb95a8 , n39711 );
buf ( R_a92_1e18bd08 , C0 );
buf ( R_b33_1e6b1d08 , n39714 );
buf ( R_2ab_1d9fc5c8 , n39717 );
buf ( R_5e6_1dd9f6e8 , C0 );
buf ( R_5c0_1ddab3a8 , n39718 );
buf ( R_600_1ddadba8 , n39719 );
buf ( R_8f4_1e09b4e8 , n39720 );
buf ( R_29d_1d9fbd08 , n39736 );
buf ( R_c11_1e6ba7c8 , n39752 );
buf ( R_4d7_1dda2208 , n39755 );
buf ( R_b43_1e6b2708 , n39758 );
buf ( R_881_1e096d08 , n39778 );
buf ( R_891_1e097708 , n39793 );
buf ( R_8b4_1e098ce8 , n39794 );
buf ( R_6ac_1dfb4788 , n39795 );
buf ( R_2f0_1d9cf148 , n39796 );
buf ( R_ad8_1e6ae428 , n39797 );
buf ( R_9bb_1e1831a8 , n39800 );
buf ( R_bd9_1e6b84c8 , n39814 );
buf ( R_39f_1d9d5ea8 , n39817 );
buf ( R_a5e_1e189c88 , C0 );
buf ( R_303_1d9cfd28 , n39820 );
buf ( R_6ae_1dfb4dc8 , C0 );
buf ( R_477_1dd9e608 , n39823 );
buf ( R_6d2_1e0981a8 , C0 );
buf ( R_38f_1d9d54a8 , n39826 );
buf ( R_4d2_1dda23e8 , C0 );
buf ( R_82f_1e0939c8 , n39829 );
buf ( R_61d_1dfaee28 , n39835 );
buf ( R_673_1dfb23e8 , n39838 );
buf ( R_578_1dda86a8 , n39839 );
buf ( R_a65_1e189be8 , n39845 );
buf ( R_9a5_1e1823e8 , n39851 );
buf ( R_744_1dfba688 , n39852 );
buf ( R_bfe_1e6ba0e8 , C0 );
buf ( R_86e_1e096628 , C0 );
buf ( R_6ce_1e0945a8 , C0 );
buf ( R_9df_1e184828 , n39855 );
buf ( R_571_1dda8248 , n39869 );
buf ( R_9e0_1e1848c8 , n39870 );
buf ( R_9de_1e184c88 , C0 );
buf ( R_41a_1ddabee8 , C0 );
buf ( R_36e_1d9d1588 , C0 );
buf ( R_6b9_1dfb4fa8 , n39976 );
buf ( R_b72_1e6b4968 , C0 );
buf ( R_73f_1dfba368 , n39979 );
buf ( R_a4d_1e188ce8 , n39985 );
buf ( R_9e1_1e184968 , n40078 );
buf ( R_2d0_1d9fdce8 , n40079 );
buf ( R_72e_1dfb9dc8 , C0 );
buf ( R_c25_1e6bb448 , n40093 );
buf ( R_8eb_1e09af48 , n40096 );
buf ( R_6eb_1dfb6ee8 , n40099 );
buf ( R_764_1dfbba88 , n40100 );
buf ( R_9b1_1e182b68 , n40107 );
buf ( R_970_1e1802c8 , n40108 );
buf ( R_bce_1e6b82e8 , C0 );
buf ( R_325_1d9d1268 , n40126 );
buf ( R_65c_1dfb1588 , n40127 );
buf ( R_643_1dfb05e8 , n40130 );
buf ( R_abf_1e18d428 , n40133 );
buf ( R_a9b_1e18bda8 , n40136 );
buf ( R_b7c_1e6b4aa8 , n40137 );
buf ( R_9ba_1e183608 , C0 );
buf ( R_bef_1e6b9288 , n40140 );
buf ( R_b14_1e6b09a8 , n40141 );
buf ( R_996_1e181f88 , C0 );
buf ( R_812_1e092ca8 , C0 );
buf ( R_4a2_1dda05e8 , C0 );
buf ( R_6e0_1dfb6808 , n40142 );
buf ( R_490_1dd9f5a8 , n40143 );
buf ( R_711_1dfb86a8 , n40149 );
buf ( R_a86_1e18ba88 , C0 );
buf ( R_342_1d9d2988 , C0 );
buf ( R_c0e_1e6baae8 , C0 );
buf ( R_8e3_1e09aa48 , n40152 );
buf ( R_646_1dfb0cc8 , C0 );
buf ( R_74d_1dfbac28 , n40158 );
buf ( R_67f_1dfb2b68 , n40161 );
buf ( R_34f_1d9d2ca8 , n40164 );
buf ( R_8f3_1e09b448 , n40167 );
buf ( R_bdc_1e6b86a8 , n40168 );
buf ( R_57f_1dda8b08 , n40171 );
buf ( R_77a_1dfbcd48 , C0 );
buf ( R_4c1_1dda1448 , n40176 );
buf ( R_b8e_1e6b5ae8 , C0 );
buf ( R_c29_1e6bb6c8 , n40189 );
buf ( R_875_1e096588 , n40210 );
buf ( R_852_1e0954a8 , C0 );
buf ( R_6a6_1dfb48c8 , C0 );
buf ( R_76f_1dfbc168 , n40213 );
buf ( R_984_1e180f48 , n40214 );
buf ( R_39a_1d9d6088 , C0 );
buf ( R_35f_1d9d36a8 , n40217 );
buf ( R_5d0_1ddabda8 , n40218 );
buf ( R_b65_1e6b3c48 , n40229 );
buf ( R_92b_1e09d748 , n40232 );
buf ( R_3eb_1d9d8e28 , n40235 );
buf ( R_53b_1dda6088 , n40238 );
buf ( R_97a_1e180e08 , C0 );
buf ( R_369_1d9d3ce8 , n40315 );
buf ( R_7f5_1e091588 , n40334 );
buf ( R_588_1dda90a8 , n40335 );
buf ( R_b6a_1e6b4468 , C0 );
buf ( R_435_1d9dbc68 , n40340 );
buf ( R_a08_1e1861c8 , n40341 );
buf ( R_7ef_1e0911c8 , n40344 );
buf ( R_781_1dfbcca8 , n40431 );
buf ( R_55c_1dda7528 , n40432 );
buf ( R_3bf_1d9d72a8 , n40435 );
buf ( R_850_1e094e68 , n40436 );
buf ( R_2ea_1d9cf288 , C0 );
buf ( R_687_1dfb3068 , n40439 );
buf ( R_795_1dfbd928 , n40444 );
buf ( R_382_1d9d5188 , C0 );
buf ( R_63e_1dfb07c8 , C0 );
buf ( R_2b7_1d9fcd48 , n40447 );
buf ( R_9b0_1e182ac8 , n40448 );
buf ( R_6dd_1dfb6628 , n40454 );
buf ( R_4be_1dda1768 , C0 );
buf ( R_bfd_1e6b9b48 , n40470 );
buf ( R_b0d_1e6b0548 , n40484 );
buf ( R_b9d_1e6b5f48 , n40497 );
buf ( R_b3a_1e6b2668 , C0 );
buf ( R_4b9_1dda0f48 , n40503 );
buf ( R_4bb_1dda1088 , n40506 );
buf ( R_9a0_1e1820c8 , n40507 );
buf ( R_83b_1e094148 , n40510 );
buf ( R_8ea_1e09b3a8 , C0 );
buf ( R_b21_1e6b11c8 , n40524 );
buf ( R_62f_1dfaf968 , n40527 );
buf ( R_91d_1e09ce88 , n40547 );
buf ( R_483_1dd9ed88 , n40550 );
buf ( R_7c0_1e08f468 , n40551 );
buf ( R_bd5_1e6b8248 , n40565 );
buf ( R_364_1d9d39c8 , n40566 );
buf ( R_322_1d9d2e88 , C0 );
buf ( R_326_1d9d1808 , C0 );
buf ( R_99b_1e181da8 , n40569 );
buf ( R_961_1e17f968 , n40575 );
buf ( R_726_1dfb98c8 , C0 );
buf ( R_a7d_1e18aae8 , n40581 );
buf ( R_826_1e09de28 , C0 );
buf ( R_89a_1dfb4648 , C0 );
buf ( R_511_1dda4648 , n40597 );
buf ( R_2fb_1d9cf828 , n40600 );
buf ( R_b5c_1e6b36a8 , n40601 );
buf ( R_8b0_1e098a68 , n40602 );
buf ( R_708_1dfb8108 , n40603 );
buf ( R_603_1ddadd88 , n40606 );
buf ( R_804_1e091ee8 , n40607 );
buf ( R_573_1dda8388 , n40610 );
buf ( R_a56_1e189a08 , C0 );
buf ( R_510_1dda45a8 , n40611 );
buf ( R_833_1e093c48 , n40614 );
buf ( R_8c1_1e099508 , n40619 );
buf ( R_966_1e180188 , C0 );
buf ( R_46d_1dd9dfc8 , n40636 );
buf ( R_bcc_1e6b7ca8 , n40637 );
buf ( R_47b_1dd9e888 , n40640 );
buf ( R_aea_1e6af468 , C0 );
buf ( R_8d1_1e099f08 , n40645 );
buf ( R_57a_1ddaa368 , C0 );
buf ( R_8f2_1e09b8a8 , C0 );
buf ( R_b35_1e6b1e48 , n40660 );
buf ( R_b05_1e6b0048 , n40673 );
buf ( R_aa9_1e18c668 , n40688 );
buf ( R_9b7_1e182f28 , n40691 );
buf ( R_3ae_1d9d6d08 , C0 );
buf ( R_50f_1dda4508 , n40694 );
buf ( R_a23_1e1872a8 , n40697 );
buf ( R_2c9_1d9fd888 , n40703 );
buf ( R_5c6_1d9d7e88 , C0 );
buf ( R_8bd_1e099288 , n40708 );
buf ( R_4b1_1dda0a48 , n40713 );
buf ( R_b45_1e6b2848 , n40799 );
buf ( R_422_1d9db588 , C0 );
buf ( R_2cc_1d9fda68 , n40800 );
buf ( R_9d5_1e1841e8 , n40807 );
buf ( R_37e_1d9d4f08 , C0 );
buf ( R_42c_1d9db6c8 , n40808 );
buf ( R_a7e_1e18b088 , C0 );
buf ( R_a8d_1e18b4e8 , n40820 );
buf ( R_50e_1dda4968 , C0 );
buf ( R_626_1dfafb48 , C0 );
buf ( R_5cc_1ddabb28 , n40821 );
buf ( R_295_1d9fb808 , n40832 );
buf ( R_a9e_1e18c488 , C0 );
buf ( R_80d_1e092488 , n40848 );
buf ( R_9af_1e182a28 , n40851 );
buf ( R_946_1e17ed88 , C0 );
buf ( R_a5c_1e189648 , n40852 );
buf ( R_5bb_1ddab088 , n40855 );
buf ( R_3e6_1d9d9008 , C0 );
buf ( R_ab3_1e18cca8 , n40858 );
buf ( R_a1e_1e187488 , C0 );
buf ( R_66a_1dfb2348 , C0 );
buf ( R_7f8_1e091768 , n40859 );
buf ( R_56e_1dda8568 , C0 );
buf ( R_3c2_1d9d7988 , C0 );
buf ( R_837_1e093ec8 , n40862 );
buf ( R_866_1e096128 , C0 );
buf ( R_65a_1dfb1948 , C0 );
buf ( R_4aa_1dda0ae8 , C0 );
buf ( R_540_1dda63a8 , n40863 );
buf ( R_61b_1dfaece8 , n40866 );
buf ( R_78a_1dfbd748 , C0 );
buf ( R_76c_1dfbbf88 , n40867 );
buf ( R_4c7_1dda1808 , n40870 );
buf ( R_47f_1dd9eb08 , n40873 );
buf ( R_34a_1d9d4a08 , C0 );
buf ( R_b57_1e6b3388 , n40876 );
buf ( R_545_1dda66c8 , n40899 );
buf ( R_c13_1e6ba908 , n40902 );
buf ( R_44c_1d9dcac8 , n40903 );
buf ( R_a0b_1e1863a8 , n40906 );
buf ( R_6d5_1dfb6128 , n40913 );
buf ( R_bf3_1e6b9508 , n40916 );
buf ( R_3ee_1d9d9508 , C0 );
buf ( R_6d7_1dfb6268 , n40919 );
buf ( R_3d6_1d9d9788 , C0 );
buf ( R_b06_1e6b05e8 , C0 );
buf ( R_9d4_1e184148 , n40920 );
buf ( R_33b_1d9d2028 , n40923 );
buf ( R_739_1dfb9fa8 , n40929 );
buf ( R_a0e_1e186a88 , C0 );
buf ( R_7dd_1e090688 , n41044 );
buf ( R_54f_1dda6d08 , n41047 );
buf ( R_926_1e09dba8 , C0 );
buf ( R_abb_1e18d1a8 , n41050 );
buf ( R_70e_1dfb89c8 , C0 );
buf ( R_ba2_1e6b6768 , C0 );
buf ( R_917_1e09cac8 , n41053 );
buf ( R_923_1e09d248 , n41056 );
buf ( R_784_1dfbce88 , n41057 );
buf ( R_920_1e09d068 , n41058 );
buf ( R_564_1dda7a28 , n41059 );
buf ( R_9a9_1e182668 , n41067 );
buf ( R_bfa_1e6b9e68 , C0 );
buf ( R_62c_1dfaf788 , n41068 );
buf ( R_8c9_1e099a08 , n41087 );
buf ( R_43c_1d9dc0c8 , n41088 );
buf ( R_b00_1e6afd28 , n41089 );
buf ( R_35d_1d9d3568 , n41131 );
buf ( R_c18_1e6bac28 , n41132 );
buf ( R_306_1d9d0408 , C0 );
buf ( R_939_1e17e068 , n41144 );
buf ( R_474_1dd9e428 , n41145 );
buf ( R_4a9_1dda0548 , n41150 );
buf ( R_2ac_1d9fc668 , n41151 );
buf ( R_609_1dfae1a8 , n41159 );
buf ( R_94c_1e17ec48 , n41160 );
buf ( R_90a_1e09c7a8 , C0 );
buf ( R_92e_1e0918a8 , C0 );
buf ( R_7be_1e08f828 , C0 );
buf ( R_825_1e093388 , n41166 );
buf ( R_559_1dda7348 , n41178 );
buf ( R_bf7_1e6b9788 , n41181 );
buf ( R_87a_1e096da8 , C0 );
buf ( R_9d3_1e1840a8 , n41184 );
buf ( R_394_1d9d57c8 , n41185 );
buf ( R_31a_1d9d1088 , C0 );
buf ( R_69f_1dfb3f68 , n41188 );
buf ( R_787_1dfbd068 , n41191 );
buf ( R_a63_1e189aa8 , n41194 );
buf ( R_9ae_1e183388 , C0 );
buf ( R_945_1e17e7e8 , n41208 );
buf ( R_537_1dda5e08 , n41211 );
buf ( R_725_1dfb9328 , n41217 );
buf ( R_b68_1e6b3e28 , n41218 );
buf ( R_7a5_1e08e388 , n41224 );
buf ( R_4eb_1dda2e88 , n41227 );
buf ( R_619_1dfaeba8 , n41233 );
buf ( R_800_1e091c68 , n41234 );
buf ( R_be8_1e6b8e28 , n41235 );
buf ( R_4ec_1dda2f28 , n41236 );
buf ( R_4ea_1dda32e8 , C0 );
buf ( R_2f1_1d9cf1e8 , n41244 );
buf ( R_5d3_1ddabf88 , n41247 );
buf ( R_6da_1dfb6948 , C0 );
buf ( R_5b6_1ddab268 , C0 );
buf ( R_3ac_1d9d66c8 , n41248 );
buf ( R_983_1e180ea8 , n41251 );
buf ( R_b73_1e6b4508 , n41254 );
buf ( R_4ed_1dda2fc8 , n41271 );
buf ( R_ada_1e6aea68 , C0 );
buf ( R_7fc_1e0919e8 , n41272 );
buf ( R_b3c_1e6b22a8 , n41273 );
buf ( R_304_1d9cfdc8 , n41274 );
buf ( R_5ab_1ddaa688 , n41277 );
buf ( R_85c_1e0955e8 , n41278 );
buf ( R_442_1d9dcc08 , C0 );
buf ( R_3ce_1d9d8608 , C0 );
buf ( R_ad5_1e6ae248 , n41284 );
buf ( R_ae8_1e6aee28 , n41285 );
buf ( R_3b4_1d9d6bc8 , n41286 );
buf ( R_8b8_1e098f68 , n41287 );
buf ( R_b46_1e6b2de8 , C0 );
buf ( R_8e8_1e09ad68 , n41288 );
buf ( R_bbf_1e6b7488 , n41291 );
buf ( R_799_1dfbdba8 , n41296 );
buf ( R_778_1dfbc708 , n41297 );
buf ( R_a4b_1e188ba8 , n41300 );
buf ( R_51d_1dda4dc8 , n41313 );
buf ( R_657_1dfb1268 , n41316 );
buf ( R_9d2_1e17f788 , C0 );
buf ( R_348_1d9d2848 , n41317 );
buf ( R_51c_1dda4d28 , n41318 );
buf ( R_8d7_1e09a2c8 , n41321 );
buf ( R_9b3_1e182ca8 , n41324 );
buf ( R_7db_1e090548 , n41327 );
buf ( R_715_1dfb8928 , n41333 );
buf ( R_68c_1dfb3388 , n41334 );
buf ( R_880_1e096c68 , n41335 );
buf ( R_29c_1d9fbc68 , n41347 );
buf ( R_b7d_1e6b4b48 , n41362 );
buf ( R_51b_1dda4c88 , n41365 );
buf ( R_bba_1e6b7668 , C0 );
buf ( R_3dc_1d9d84c8 , n41366 );
buf ( R_5a0_1dda9fa8 , n41367 );
buf ( R_75f_1dfbb768 , n41370 );
buf ( R_b7f_1e6b4c88 , n41373 );
buf ( R_b16_1e6b0fe8 , C0 );
buf ( R_ba3_1e6b6308 , n41376 );
buf ( R_654_1dfb1088 , n41377 );
buf ( R_bc7_1e6b7988 , n41380 );
buf ( R_2a3_1d9fc0c8 , n41383 );
buf ( R_6f0_1dfb7208 , n41384 );
buf ( R_7a1_1e08e108 , n41401 );
buf ( R_371_1d9d41e8 , n41459 );
buf ( R_51a_1dda50e8 , C0 );
buf ( R_ab7_1e18cf28 , n41462 );
buf ( R_7e6_1e099828 , C0 );
buf ( R_b6b_1e6b4008 , n41465 );
buf ( R_9ad_1e1828e8 , n41471 );
buf ( R_935_1e09dd88 , n41489 );
buf ( R_b8a_1e6bb768 , C0 );
buf ( R_69d_1dfb3e28 , n41616 );
buf ( R_45e_1d9ddb08 , C0 );
buf ( R_a1a_1e187208 , C0 );
buf ( R_a49_1e188a68 , n41621 );
buf ( R_a09_1e186268 , n41674 );
buf ( R_496_1dd9fe68 , C0 );
buf ( R_336_1d9d2208 , C0 );
buf ( R_5df_1ddac708 , n41677 );
buf ( R_5c7_1ddab808 , n41680 );
buf ( R_990_1e1816c8 , n41681 );
buf ( R_6c9_1dfb59a8 , n41793 );
buf ( R_2eb_1d9cee28 , n41796 );
buf ( R_2b8_1d9fcde8 , n41797 );
buf ( R_ae0_1e6ae928 , n41798 );
buf ( R_b2f_1e6b1a88 , n41801 );
buf ( R_84d_1e094c88 , n41818 );
buf ( R_a12_1e186d08 , C0 );
buf ( R_74f_1dfbad68 , n41821 );
buf ( R_a35_1e187de8 , n41826 );
buf ( R_28e_1d9fb3a8 , n41837 );
buf ( R_81a_1e0936a8 , C0 );
buf ( R_487_1dd9f008 , n41840 );
buf ( R_c1c_1e6baea8 , n41841 );
buf ( R_7a8_1e08e568 , n41842 );
buf ( R_471_1dd9e248 , n41847 );
buf ( R_766_1e0986a8 , C0 );
buf ( R_38b_1d9d5228 , n41850 );
buf ( R_a7b_1e18a9a8 , n41853 );
buf ( R_b52_1e6b8568 , C0 );
buf ( R_9ff_1e185c28 , n41856 );
buf ( R_7b9_1e08f008 , n41861 );
buf ( R_67b_1dfb28e8 , n41864 );
buf ( R_a00_1e185cc8 , n41865 );
buf ( R_9fe_1e6bb9e8 , C0 );
buf ( R_980_1e180cc8 , n41866 );
buf ( R_874_1e0964e8 , n41867 );
buf ( R_49c_1dd9fd28 , n41868 );
buf ( R_58c_1dda9328 , n41869 );
buf ( R_45f_1d9dd6a8 , n41872 );
buf ( R_98a_1e181808 , C0 );
buf ( R_8e2_1e09aea8 , C0 );
buf ( R_6ba_1dfb5548 , C0 );
buf ( R_bd8_1e6b8428 , n41873 );
buf ( R_a8b_1e18b3a8 , n41876 );
buf ( R_a01_1e185d68 , n42258 );
buf ( R_6b3_1dfb4be8 , n42261 );
buf ( R_60d_1dfae428 , n42269 );
buf ( R_6e8_1dfb6d08 , n42270 );
buf ( R_399_1d9d5ae8 , n42276 );
buf ( R_a16_1e186f88 , C0 );
buf ( R_bc2_1e6b7b68 , C0 );
buf ( R_32b_1d9d1628 , n42279 );
buf ( R_434_1d9dbbc8 , n42280 );
buf ( R_a24_1e187348 , n42281 );
buf ( R_377_1d9d45a8 , n42284 );
buf ( R_3cc_1d9d7ac8 , n42285 );
buf ( R_a68_1e189dc8 , n42286 );
buf ( R_963_1e17faa8 , n42289 );
buf ( R_7c5_1e08f788 , n42294 );
buf ( R_615_1dfae928 , n42301 );
buf ( R_8a2_1dfb9b48 , C0 );
buf ( R_722_1dfb9648 , C0 );
buf ( R_288_1d9f96e8 , n42328 );
buf ( R_556_1dda7668 , C0 );
buf ( R_748_1dfba908 , n42329 );
buf ( R_865_1e095b88 , n42341 );
buf ( R_607_1dfae068 , n42344 );
buf ( R_691_1dfb36a8 , n42473 );
buf ( R_978_1e1807c8 , n42474 );
buf ( R_84f_1e094dc8 , n42477 );
buf ( R_2cd_1d9fdb08 , n42483 );
buf ( R_ae2_1e6aef68 , C0 );
buf ( R_a1f_1e187028 , n42486 );
buf ( R_721_1dfb90a8 , n42492 );
buf ( R_733_1dfb9be8 , n42495 );
buf ( R_9e3_1e184aa8 , n42498 );
buf ( R_9e4_1e184b48 , n42499 );
buf ( R_c23_1e6bb308 , n42502 );
buf ( R_9e2_1e184f08 , C0 );
buf ( R_7ae_1dfbb1c8 , C0 );
buf ( R_91a_1e09d1a8 , C0 );
buf ( R_b84_1e6b4fa8 , n42503 );
buf ( R_b92_1e181088 , C0 );
buf ( R_ba4_1e6b63a8 , n42504 );
buf ( R_754_1dfbb088 , n42505 );
buf ( R_5a4_1ddaa228 , n42506 );
buf ( R_9a4_1e182348 , n42507 );
buf ( R_b08_1e6b0228 , n42508 );
buf ( R_9e5_1e184be8 , n42558 );
buf ( R_617_1dfaea68 , n42561 );
buf ( R_5ce_1ddac168 , C0 );
buf ( R_b89_1e6b52c8 , n42578 );
buf ( R_7b2_1e09b128 , C0 );
buf ( R_460_1d9dd748 , n42579 );
buf ( R_5e4_1ddaca28 , n42580 );
buf ( R_30a_1d9d0688 , C0 );
buf ( R_a0c_1e186448 , n42581 );
buf ( R_910_1e09c668 , n42582 );
buf ( R_553_1dda6f88 , n42585 );
buf ( R_86d_1e096088 , n42601 );
buf ( R_a0f_1e186628 , n42604 );
buf ( R_719_1dfb8ba8 , n42610 );
buf ( R_b48_1e6b2a28 , n42611 );
buf ( R_316_1d9d0e08 , C0 );
buf ( R_901_1e09bd08 , n42616 );
buf ( R_611_1dfae6a8 , n42624 );
buf ( R_ac5_1e18d7e8 , n42688 );
buf ( R_6c4_1dfb5688 , n42689 );
buf ( R_53c_1dda6128 , n42690 );
buf ( R_712_1dfb8c48 , C0 );
buf ( R_2f6_1d9cfc88 , C0 );
buf ( R_829_1e093608 , n42705 );
buf ( R_89d_1e097e88 , n42735 );
buf ( R_8d0_1e099e68 , n42736 );
buf ( R_8ac_1e0987e8 , n42737 );
buf ( R_8a0_1e098068 , n42738 );
buf ( R_aef_1e6af288 , n42741 );
buf ( R_759_1dfbb3a8 , n42746 );
buf ( R_a6d_1e18a0e8 , n42841 );
buf ( R_6bf_1dfb5368 , n42844 );
buf ( R_982_1e182c08 , C0 );
buf ( R_bdb_1e6b8608 , n42847 );
buf ( R_684_1dfb2e88 , n42848 );
buf ( R_7b7_1e08eec8 , n42851 );
buf ( R_478_1dd9e6a8 , n42852 );
buf ( R_be1_1e6b89c8 , n42871 );
buf ( R_b55_1e6b3248 , n42885 );
buf ( R_79b_1dfbdce8 , n42888 );
buf ( R_c27_1e6bb588 , n42891 );
buf ( R_96f_1e180228 , n42894 );
buf ( R_42b_1d9db628 , n42897 );
buf ( R_6cd_1dfb5c28 , n42901 );
buf ( R_652_1dfb16c8 , C0 );
buf ( R_71d_1dfb8e28 , n42907 );
buf ( R_703_1dfb7de8 , n42910 );
buf ( R_a54_1e189148 , n42911 );
buf ( R_4a3_1dda0188 , n42914 );
buf ( R_634_1dfafc88 , n42915 );
buf ( R_2ad_1d9fc708 , n42921 );
buf ( R_4cc_1dda1b28 , n42922 );
buf ( R_2a1_1d9fbf88 , n44733 );
buf ( R_93a_1e0977a8 , C0 );
buf ( R_a78_1e18a7c8 , n44734 );
buf ( R_c03_1e6b9f08 , n44737 );
buf ( R_72c_1dfb9788 , n44738 );
buf ( R_809_1e092208 , n44754 );
buf ( R_5b0_1ddaa9a8 , n44755 );
buf ( R_44b_1d9dca28 , n44758 );
buf ( R_952_1ddab768 , C0 );
buf ( R_899_1e097c08 , n44774 );
buf ( R_bd4_1e6b81a8 , n44775 );
buf ( R_a94_1e18b948 , n44776 );
buf ( R_6b1_1dfb4aa8 , n44869 );
buf ( R_491_1dd9f648 , n44874 );
buf ( R_5ca_1d9dae08 , C0 );
buf ( R_6f5_1dfb7528 , n44880 );
buf ( R_9c9_1e183a68 , n44888 );
buf ( R_75a_1dfbb948 , C0 );
buf ( R_461_1d9dd7e8 , n44903 );
buf ( R_7c3_1e08f648 , n44906 );
buf ( R_569_1dda7d48 , n44985 );
buf ( R_a75_1e18a5e8 , n44991 );
buf ( R_7ec_1e090fe8 , n44992 );
buf ( R_c20_1e6bb128 , n44993 );
buf ( R_96d_1e1800e8 , n45000 );
buf ( R_54a_1dda6ee8 , C0 );
buf ( R_b31_1e6b1bc8 , n45015 );
buf ( R_5bf_1ddab308 , n45018 );
buf ( R_900_1e09bc68 , n45019 );
buf ( R_b74_1e6b45a8 , n45020 );
buf ( R_940_1e17e4c8 , n45021 );
buf ( R_8dd_1e09a688 , n45026 );
buf ( R_a88_1e18b1c8 , n45027 );
buf ( R_743_1dfba5e8 , n45030 );
buf ( R_2d1_1d9fdd88 , n45036 );
buf ( R_4b3_1dda0b88 , n45039 );
buf ( R_48c_1dd9f328 , n45040 );
buf ( R_419_1d9daae8 , n45053 );
buf ( R_2ba_1d9fd428 , C0 );
buf ( R_898_1e097b68 , n45054 );
buf ( R_354_1d9d2fc8 , n45055 );
buf ( R_3c9_1d9d78e8 , n45061 );
buf ( R_afd_1e6afb48 , n45066 );
buf ( R_698_1dfb3b08 , n45067 );
buf ( R_8c8_1e099968 , n45068 );
buf ( R_aff_1e6afc88 , n45071 );
buf ( R_59c_1dda9d28 , n45072 );
buf ( R_43b_1d9dc028 , n45075 );
buf ( R_3e1_1d9d87e8 , n45081 );
buf ( R_7d8_1e090368 , n45082 );
buf ( R_624_1dfaf288 , n45083 );
buf ( R_ace_1e6ae2e8 , C0 );
buf ( R_294_1d9fb768 , n45094 );
buf ( R_818_1e092b68 , n45095 );
buf ( R_9c8_1e1839c8 , n45096 );
buf ( R_5c8_1ddab8a8 , n45097 );
buf ( R_c2f_1e6bba88 , n45100 );
buf ( R_ba5_1e6b6448 , n45108 );
buf ( R_6d0_1dfb5e08 , n45109 );
buf ( R_820_1e093068 , n45110 );
buf ( R_30e_1d9d0908 , C0 );
buf ( R_99f_1e182028 , n45113 );
buf ( R_73e_1dfba7c8 , C0 );
buf ( R_4ef_1dda3108 , n45116 );
buf ( R_451_1d9dcde8 , n45122 );
buf ( R_678_1dfb2708 , n45123 );
buf ( R_663_1dfb19e8 , n45126 );
buf ( R_5fa_1e091128 , C0 );
buf ( R_312_1d9d0b88 , C0 );
buf ( R_a45_1e1887e8 , n45131 );
buf ( R_b18_1e6b0c28 , n45132 );
buf ( R_4f0_1dda31a8 , n45133 );
buf ( R_4ee_1dda3568 , C0 );
buf ( R_7ab_1e08e748 , n45136 );
buf ( R_305_1d9cfe68 , n45142 );
buf ( R_955_1e17f1e8 , n45145 );
buf ( R_373_1d9d4328 , n45148 );
buf ( R_a39_1e188068 , n45153 );
buf ( R_669_1dfb1da8 , n45160 );
buf ( R_3a5_1d9d6268 , n45166 );
buf ( R_c0d_1e6ba548 , n45182 );
buf ( R_4f1_1dda3248 , n45194 );
buf ( R_541_1dda6448 , n45217 );
buf ( R_69a_1dfb4148 , C0 );
buf ( R_b90_1e6b5728 , n45218 );
buf ( R_99a_1e182208 , C0 );
buf ( R_960_1e17f8c8 , n45219 );
buf ( R_6a9_1dfb45a8 , n45253 );
buf ( R_4bc_1dda1128 , n45254 );
buf ( R_897_1e097ac8 , n45257 );
buf ( R_701_1dfb7ca8 , n45263 );
buf ( R_36c_1d9d3ec8 , n45264 );
buf ( R_60b_1dfae2e8 , n45267 );
buf ( R_583_1dda8d88 , n45270 );
buf ( R_330_1d9d1948 , n45271 );
buf ( R_bb6_1e6b73e8 , C0 );
buf ( R_71e_1dfb93c8 , C0 );
buf ( R_590_1dda95a8 , n45272 );
buf ( R_29e_1dda2668 , C0 );
buf ( R_b0f_1e6b0688 , n45275 );
buf ( R_a1b_1e186da8 , n45278 );
buf ( R_550_1dda6da8 , n45279 );
buf ( R_ac8_1e18d9c8 , n45280 );
buf ( R_a9d_1e18bee8 , n45341 );
buf ( R_561_1dda7848 , n45354 );
buf ( R_80e_1e092a28 , C0 );
buf ( R_9b6_1e187708 , C0 );
buf ( R_5e8_1ddacca8 , n45355 );
buf ( R_613_1dfae7e8 , n45358 );
buf ( R_b6c_1e6b40a8 , n45359 );
buf ( R_3d3_1d9d7f28 , n45362 );
buf ( R_31f_1d9d0ea8 , n45365 );
buf ( R_9c7_1e183928 , n45368 );
buf ( R_5dd_1ddac5c8 , n45373 );
buf ( R_78e_1dfbd9c8 , C0 );
buf ( R_a13_1e1868a8 , n45376 );
buf ( R_70c_1dfb8388 , n45377 );
buf ( R_885_1e096f88 , n45393 );
buf ( R_85b_1e095548 , n45396 );
buf ( R_8ff_1e09bbc8 , n45399 );
buf ( R_716_1dfb8ec8 , C0 );
buf ( R_2b9_1d9fce88 , n45405 );
buf ( R_b69_1e6b3ec8 , n45419 );
buf ( R_356_1d9d3608 , C0 );
buf ( R_2e6_1d9cf008 , C0 );
buf ( R_484_1dd9ee28 , n45420 );
buf ( R_2ec_1d9ceec8 , n45421 );
buf ( R_acb_1e18dba8 , n45424 );
buf ( R_813_1e092848 , n45427 );
buf ( R_4c3_1dda1588 , n45430 );
buf ( R_a47_1e188928 , n45433 );
buf ( R_81d_1e092e88 , n45450 );
buf ( R_8e7_1e09acc8 , n45453 );
buf ( R_5ef_1ddad108 , n45456 );
buf ( R_896_1e094828 , C0 );
buf ( R_bec_1e6b90a8 , n45457 );
buf ( R_b2b_1e6b1808 , n45460 );
buf ( R_4ab_1dda0688 , n45463 );
buf ( R_7e4_1e090ae8 , n45464 );
buf ( R_a33_1e187ca8 , n45467 );
buf ( R_47c_1dd9e928 , n45468 );
buf ( R_8d6_1e09a728 , C0 );
buf ( R_87f_1e096bc8 , n45471 );
buf ( R_5b5_1ddaacc8 , n45488 );
buf ( R_651_1dfb0ea8 , n45494 );
buf ( R_3da_1d9d8888 , C0 );
buf ( R_538_1dda5ea8 , n45495 );
buf ( R_675_1dfb2528 , n45502 );
buf ( R_60f_1dfae568 , n45505 );
buf ( R_29b_1d9fbbc8 , n45512 );
buf ( R_aa6_1e18c988 , C0 );
buf ( R_3bd_1d9d7168 , n45518 );
buf ( R_be5_1e6b8c48 , n45530 );
buf ( R_c0a_1e6ba868 , C0 );
buf ( R_5f5_1ddad4c8 , n45540 );
buf ( R_b4b_1e6b2c08 , n45543 );
buf ( R_7b1_1e08eb08 , n45548 );
buf ( R_95d_1e17f6e8 , n45554 );
buf ( R_a17_1e186b28 , n45557 );
buf ( R_a29_1e187668 , n45561 );
buf ( R_71a_1dfb9148 , C0 );
buf ( R_693_1dfb37e8 , n45564 );
buf ( R_77b_1dfbc8e8 , n45567 );
buf ( R_9c6_1e183d88 , C0 );
buf ( R_3a7_1d9d63a8 , n45570 );
buf ( R_bc0_1e6b7528 , n45571 );
buf ( R_68e_1dfb39c8 , C0 );
buf ( R_335_1d9d1c68 , n45643 );
buf ( R_5eb_1ddace88 , n45646 );
buf ( R_ad7_1e6ae388 , n45649 );
buf ( R_765_1dfbbb28 , n45656 );
buf ( R_387_1d9d4fa8 , n45659 );
buf ( R_9a8_1e1825c8 , n45660 );
buf ( R_632_1dfb0048 , C0 );
buf ( R_6e5_1dfb6b28 , n45666 );
buf ( R_772_1dfbc848 , C0 );
buf ( R_995_1e1819e8 , n45672 );
buf ( R_7d6_1e090728 , C0 );
buf ( R_598_1dda9aa8 , n45673 );
buf ( R_a70_1e18a2c8 , n45674 );
buf ( R_a25_1e1873e8 , n45739 );
buf ( R_bbb_1e6b7208 , n45742 );
buf ( R_6f2_1dfb7848 , C0 );
buf ( R_a41_1e188568 , n45747 );
buf ( R_a66_1e18a188 , C0 );
buf ( R_a3d_1e1882e8 , n45752 );
buf ( R_341_1d9d23e8 , n45816 );
buf ( R_594_1dda9828 , n45817 );
buf ( R_4fe_1dda5868 , C0 );
buf ( R_480_1dd9eba8 , n45818 );
buf ( R_6ab_1dfb46e8 , n45821 );
buf ( R_84c_1e094be8 , n45822 );
buf ( R_660_1dfb1808 , n45823 );
buf ( R_a20_1e1870c8 , n45824 );
buf ( R_abe_1e6b64e8 , C0 );
buf ( R_566_1dda8068 , C0 );
buf ( R_7c8_1e08f968 , n45825 );
buf ( R_5c2_1d9fc2a8 , C0 );
buf ( R_989_1e181268 , n45831 );
buf ( R_8a8_1e098568 , n45832 );
buf ( R_2a4_1d9fc168 , n45833 );
buf ( R_7d5_1e090188 , n45838 );
buf ( R_8fe_1e09c028 , C0 );
buf ( R_3b7_1d9d6da8 , n45841 );
buf ( R_6b8_1dfb4f08 , n45842 );
buf ( R_8b3_1e098c48 , n45845 );
buf ( R_94f_1e17ee28 , n45848 );
buf ( R_9fb_1e1859a8 , n45851 );
buf ( R_a10_1e1866c8 , n45852 );
buf ( R_b36_1e6b23e8 , C0 );
buf ( R_aa0_1e18c0c8 , n45853 );
buf ( R_c1a_1e6bb268 , C0 );
buf ( R_82c_1e0937e8 , n45854 );
buf ( R_4d1_1dda1e48 , n45859 );
buf ( R_6fc_1dfb7988 , n45860 );
buf ( R_9fa_1e185e08 , C0 );
buf ( R_9fc_1e185a48 , n45861 );
buf ( R_a0d_1e1864e8 , n45918 );
buf ( R_be2_1e6b8f68 , C0 );
buf ( R_b02_1e6b8068 , C0 );
buf ( R_a28_1e1875c8 , n45919 );
buf ( R_4fd_1dda39c8 , n45935 );
buf ( R_5fd_1ddad9c8 , n47765 );
buf ( R_873_1e096448 , n47768 );
buf ( R_9fd_1e185ae8 , n47847 );
buf ( R_a6b_1e189fa8 , n47850 );
buf ( R_aa3_1e18c2a8 , n47853 );
buf ( R_738_1dfb9f08 , n47854 );
buf ( R_805_1e091f88 , n47868 );
buf ( R_2f7_1d9cf5a8 , n47871 );
buf ( R_5ba_1ddab4e8 , C0 );
buf ( R_57d_1dda89c8 , n47883 );
buf ( R_475_1dd9e4c8 , n47888 );
buf ( R_433_1d9dbb28 , n47891 );
buf ( R_aed_1e6af148 , n47899 );
buf ( R_4fc_1dda3928 , n47900 );
buf ( R_3a0_1d9d5f48 , n47901 );
buf ( R_3f7_1d9d95a8 , n47904 );
buf ( R_367_1d9d3ba8 , n47907 );
buf ( R_947_1e17e928 , n47910 );
buf ( R_b1a_1e6b1268 , C0 );
buf ( R_525_1dda52c8 , n47923 );
buf ( R_50d_1dda43c8 , n47939 );
buf ( R_390_1d9d5548 , n47940 );
buf ( R_6fe_1dfb7fc8 , C0 );
buf ( R_6f7_1dfb7668 , n47943 );
buf ( R_2ae_1d9fcca8 , C0 );
buf ( R_864_1e095ae8 , n47944 );
buf ( R_9e7_1e184d28 , n47947 );
buf ( R_524_1dda5228 , n47948 );
buf ( R_50c_1dda4328 , n47949 );
buf ( R_9e6_1e185188 , C0 );
buf ( R_9e8_1e184dc8 , n47950 );
buf ( R_9b2_1e183108 , C0 );
buf ( R_7e2_1dfbaf48 , C0 );
buf ( R_622_1dfaf648 , C0 );
buf ( R_b4e_1e184508 , C0 );
buf ( R_a91_1e18b768 , n47956 );
buf ( R_a84_1e18af48 , n47957 );
buf ( R_4ce_1dda2168 , C0 );
buf ( R_bb2_1e6b7168 , C0 );
buf ( R_523_1dda5188 , n47960 );
buf ( R_50b_1dda4288 , n47963 );
buf ( R_9e9_1e184e68 , n48035 );
buf ( R_4f3_1dda3388 , n48038 );
buf ( R_4fb_1dda3888 , n48041 );
buf ( R_4f2_1ddad068 , C0 );
buf ( R_4f4_1dda3428 , n48042 );
buf ( R_55e_1dda7b68 , C0 );
buf ( R_84e_1e095228 , C0 );
buf ( R_a76_1e18ab88 , C0 );
buf ( R_5c9_1ddab948 , n48049 );
buf ( R_343_1d9d2528 , n48052 );
buf ( R_a73_1e18a4a8 , n48055 );
buf ( R_7cd_1e08fc88 , n48061 );
buf ( R_522_1dda55e8 , C0 );
buf ( R_50a_1dda46e8 , C0 );
buf ( R_4f5_1dda34c8 , n48073 );
buf ( R_396_1d9d5e08 , C0 );
buf ( R_7f9_1e091808 , n48088 );
buf ( R_681_1dfb2ca8 , n48185 );
buf ( R_37b_1d9d4828 , n48188 );
buf ( R_639_1dfaffa8 , n48194 );
buf ( R_76d_1dfbc028 , n48199 );
buf ( R_78b_1dfbd2e8 , n48202 );
buf ( R_6a3_1dfb41e8 , n48205 );
buf ( R_9ac_1e182848 , n48206 );
buf ( R_86c_1e095fe8 , n48207 );
buf ( R_c08_1e6ba228 , n48208 );
buf ( R_2fc_1d9cf8c8 , n48209 );
buf ( R_7f0_1e091268 , n48210 );
buf ( R_c31_1e6bbbc8 , n48214 );
buf ( R_a52_1e189508 , C0 );
buf ( R_ab2_1e18d108 , C0 );
buf ( R_28d_1d9fb308 , n48222 );
buf ( R_bcb_1e6b7c08 , n48225 );
buf ( R_4fa_1dda3f68 , C0 );
buf ( R_2bb_1d9fcfc8 , n48228 );
buf ( R_b3f_1e6b2488 , n48231 );
buf ( R_a27_1e187528 , n48234 );
buf ( R_362_1d9d3d88 , C0 );
buf ( R_497_1dd9fa08 , n48237 );
buf ( R_64f_1dfb0d68 , n48240 );
buf ( R_bd7_1e6b8388 , n48243 );
buf ( R_b75_1e6b4648 , n48258 );
buf ( R_98f_1e181628 , n48261 );
buf ( R_6ed_1dfb7028 , n48267 );
buf ( R_7d3_1e090048 , n48270 );
buf ( R_b27_1e6b1588 , n48273 );
buf ( R_39b_1d9d5c28 , n48276 );
buf ( R_8cf_1e099dc8 , n48279 );
buf ( R_689_1dfb31a8 , n48356 );
buf ( R_7c6_1e08fd28 , C0 );
buf ( R_b2d_1e6b1948 , n48371 );
buf ( R_92a_1e092f28 , C0 );
buf ( R_66c_1dfb1f88 , n48372 );
buf ( R_956_1e6b00e8 , C0 );
buf ( R_b96_1e18ce88 , C0 );
buf ( R_bae_1e6b6ee8 , C0 );
buf ( R_94d_1e17ece8 , n48384 );
buf ( R_785_1dfbcf28 , n48389 );
buf ( R_6e2_1dfb6e48 , C0 );
buf ( R_65e_1dfb5cc8 , C0 );
buf ( R_42a_1d9dba88 , C0 );
buf ( R_7e8_1e090d68 , n48390 );
buf ( R_b4d_1e6b2d48 , n48418 );
buf ( R_bff_1e6b9c88 , n48421 );
buf ( R_3c0_1d9d7348 , n48422 );
buf ( R_44a_1d9dce88 , C0 );
buf ( R_2fe_1d9cff08 , C0 );
buf ( R_383_1d9d4d28 , n48425 );
buf ( R_928_1e09d568 , n48426 );
buf ( R_488_1dd9f0a8 , n48427 );
buf ( R_5aa_1ddaaae8 , C0 );
buf ( R_3fd_1d9d9968 , n48433 );
buf ( R_7d0_1e08fe68 , n48434 );
buf ( R_7b4_1e08ece8 , n48435 );
buf ( R_4d8_1dda22a8 , n48436 );
buf ( R_418_1d9daa48 , n48437 );
buf ( R_a43_1e1886a8 , n48440 );
buf ( R_327_1d9d13a8 , n48443 );
buf ( R_849_1e094a08 , n48459 );
buf ( R_b5f_1e6b3888 , n48462 );
buf ( R_4d3_1dda1f88 , n48465 );
buf ( R_a97_1e18bb28 , n48468 );
buf ( R_aba_1e18d608 , C0 );
buf ( R_ab1_1e18cb68 , n48473 );
buf ( R_97f_1e180c28 , n48476 );
buf ( R_788_1dfbd108 , n48477 );
buf ( R_a1c_1e186e48 , n48478 );
buf ( R_b11_1e6b07c8 , n48491 );
buf ( R_a37_1e187f28 , n48494 );
buf ( R_801_1e091d08 , n48512 );
buf ( R_581_1dda8c48 , n48526 );
buf ( R_49d_1dd9fdc8 , n48531 );
buf ( R_56b_1dda7e88 , n48534 );
buf ( R_4da_1dda3ce8 , C0 );
buf ( R_7f2_1e09d6a8 , C0 );
buf ( R_53d_1dda61c8 , n48553 );
buf ( R_3df_1d9d86a8 , n48556 );
buf ( R_429_1d9db4e8 , n48561 );
buf ( R_8dc_1e09a5e8 , n48562 );
buf ( R_a14_1e186948 , n48563 );
buf ( R_9d6_1e186088 , C0 );
buf ( R_add_1e6ae748 , n48569 );
buf ( R_b6d_1e6b4148 , n48584 );
buf ( R_c1e_1e6b4e68 , C0 );
buf ( R_7fd_1e091a88 , n48598 );
buf ( R_859_1e095408 , n48614 );
buf ( R_b23_1e6b1308 , n48617 );
buf ( R_afc_1e6afaa8 , n48618 );
buf ( R_913_1e09c848 , n48621 );
buf ( R_450_1d9dcd48 , n48622 );
buf ( R_7cb_1e08fb48 , n48625 );
buf ( R_b38_1e6b2028 , n48626 );
buf ( R_a26_1e187988 , C0 );
buf ( R_74c_1dfbab88 , n48627 );
buf ( R_35b_1d9d3428 , n48630 );
buf ( R_962_1e17ff08 , C0 );
buf ( R_2e7_1d9ceba8 , n48633 );
buf ( R_8c0_1e099468 , n48634 );
buf ( R_8c7_1e0998c8 , n48637 );
buf ( R_afe_1e6b5d68 , C0 );
buf ( R_977_1e180728 , n48640 );
buf ( R_925_1e09d388 , n48655 );
buf ( R_919_1e09cc08 , n48671 );
buf ( R_728_1dfb9508 , n48672 );
buf ( R_43a_1d9dc488 , C0 );
buf ( R_bf0_1e6b9328 , n48673 );
buf ( R_9a3_1e1822a8 , n48676 );
buf ( R_3af_1d9d68a8 , n48679 );
buf ( R_930_1e09da68 , n48680 );
buf ( R_90c_1e09c3e8 , n48681 );
buf ( R_5a9_1ddaa548 , n48696 );
buf ( R_659_1dfb13a8 , n48704 );
buf ( R_c0f_1e6ba688 , n48707 );
buf ( R_307_1d9cffa8 , n48710 );
buf ( R_8bc_1e0991e8 , n48711 );
buf ( R_2ed_1d9cef68 , n48719 );
buf ( R_770_1dfbc208 , n48720 );
buf ( R_34b_1d9d2a28 , n48723 );
buf ( R_37f_1d9d4aa8 , n48726 );
buf ( R_5f4_1ddad428 , n48727 );
buf ( R_779_1dfbc7a8 , n48732 );
buf ( R_46a_1dd9f468 , C0 );
buf ( R_be0_1e6b8928 , n48733 );
buf ( R_bd3_1e6b8108 , n48736 );
buf ( R_466_1d9d9c88 , C0 );
buf ( R_77e_1dfbcfc8 , C0 );
buf ( R_575_1dda84c8 , n48754 );
buf ( R_4ff_1dda3b08 , n48757 );
buf ( R_a18_1e186bc8 , n48758 );
buf ( R_bda_1e6b8a68 , C0 );
buf ( R_31b_1d9d0c28 , n48761 );
buf ( R_3c6_1d9d7c08 , C0 );
buf ( R_792_1dfbdc48 , C0 );
buf ( R_54b_1dda6a88 , n48764 );
buf ( R_6bd_1dfb5228 , n48856 );
buf ( R_b50_1e6b2f28 , n48857 );
buf ( R_a61_1e189968 , n48863 );
buf ( R_b8b_1e6b5408 , n48866 );
buf ( R_b80_1e6b4d28 , n48867 );
buf ( R_33c_1d9d20c8 , n48868 );
buf ( R_3c3_1d9d7528 , n48871 );
buf ( R_666_1dfb20c8 , C0 );
buf ( R_c2a_1e6bbc68 , C0 );
buf ( R_359_1d9d32e8 , n48919 );
buf ( R_415_1d9da868 , n48933 );
buf ( R_5da_1ddac8e8 , C0 );
buf ( R_577_1dda8608 , n48936 );
buf ( R_637_1dfafe68 , n48939 );
buf ( R_9f7_1e185728 , n48942 );
buf ( R_570_1dda81a8 , n48943 );
buf ( R_9f6_1e185b88 , C0 );
buf ( R_9f8_1e1857c8 , n48944 );
buf ( R_a6e_1e18a688 , C0 );
buf ( R_73d_1dfba228 , n48950 );
buf ( R_293_1d9fb6c8 , n48960 );
buf ( R_884_1e096ee8 , n48961 );
buf ( R_3a2_1d9d6588 , C0 );
buf ( R_9f9_1e185868 , n49036 );
buf ( R_957_1e17f328 , n49039 );
buf ( R_ab6_1e6b5fe8 , C0 );
buf ( R_760_1dfbb808 , n49040 );
buf ( R_a21_1e187168 , n49091 );
buf ( R_bb7_1e6b6f88 , n49094 );
buf ( R_9eb_1e184fa8 , n49097 );
buf ( R_a3f_1e188428 , n49100 );
buf ( R_747_1dfba868 , n49103 );
buf ( R_4bf_1dda1308 , n49106 );
buf ( R_3d7_1d9d81a8 , n49109 );
buf ( R_4a4_1dda0228 , n49110 );
buf ( R_441_1d9dc3e8 , n49115 );
buf ( R_7ce_1e090228 , C0 );
buf ( R_85a_1e0959a8 , C0 );
buf ( R_66f_1dfb2168 , n49118 );
buf ( R_9ea_1e185408 , C0 );
buf ( R_9ec_1e185048 , n49119 );
buf ( R_a3b_1e1881a8 , n49122 );
buf ( R_ad4_1e6ae1a8 , n49123 );
buf ( R_b94_1e6b59a8 , n49124 );
buf ( R_467_1d9ddba8 , n49127 );
buf ( R_96e_1e180688 , C0 );
buf ( R_323_1d9d1128 , n49130 );
buf ( R_6ea_1dfb7348 , C0 );
buf ( R_6ca_1dfb5f48 , C0 );
buf ( R_9ed_1e1850e8 , n49201 );
buf ( R_ae7_1e6aed88 , n49204 );
buf ( R_830_1e093a68 , n49205 );
buf ( R_6d9_1dfb63a8 , n49211 );
buf ( R_8e6_1e08f0a8 , C0 );
buf ( R_6a1_1dfb40a8 , n49358 );
buf ( R_710_1dfb8608 , n49359 );
buf ( R_b41_1e6b25c8 , n49374 );
buf ( R_732_1dfba048 , C0 );
buf ( R_6df_1dfb6768 , n49377 );
buf ( R_a11_1e186768 , n49431 );
buf ( R_a8f_1e18b628 , n49434 );
buf ( R_b97_1e6b5b88 , n49437 );
buf ( R_bc6_1e6b7de8 , C0 );
buf ( R_4db_1dda2488 , n49440 );
buf ( R_9d7_1e184328 , n49443 );
buf ( R_b29_1e6b16c8 , n49458 );
buf ( R_57e_1dda8f68 , C0 );
buf ( R_29a_1d9fbb28 , n49462 );
buf ( R_36f_1d9d40a8 , n49465 );
buf ( R_3e4_1d9d89c8 , n49466 );
buf ( R_7bc_1e08f1e8 , n49467 );
buf ( R_87e_1e097028 , C0 );
buf ( R_b1c_1e6b0ea8 , n49468 );
buf ( R_aab_1e18c7a8 , n49471 );
buf ( R_96c_1e180048 , n49472 );
buf ( R_551_1dda6e48 , n49484 );
buf ( R_6d4_1dfb6088 , n49485 );
buf ( R_2af_1d9fc848 , n49488 );
buf ( R_479_1dd9e748 , n49493 );
buf ( R_5a3_1ddaa188 , n49496 );
buf ( R_672_1dfb2848 , C0 );
buf ( R_587_1dda9008 , n49499 );
buf ( R_767_1dfbbc68 , n49502 );
buf ( R_395_1d9d5868 , n49508 );
buf ( R_3e9_1d9d8ce8 , n49514 );
buf ( R_2f8_1d9cf648 , n49515 );
buf ( R_64c_1dfb0b88 , n49516 );
buf ( R_5e1_1ddac848 , n49521 );
buf ( R_3fc_1d9d98c8 , n49522 );
buf ( R_468_1d9ddc48 , n49523 );
buf ( R_3ba_1d9d7488 , C0 );
buf ( R_55b_1dda7488 , n49526 );
buf ( R_67e_1dfb2fc8 , C0 );
buf ( R_8b7_1e098ec8 , n49529 );
buf ( R_879_1e096808 , n49546 );
buf ( R_b5b_1e6b3608 , n49549 );
buf ( R_a82_1e18b588 , C0 );
buf ( R_ae5_1e6aec48 , n49564 );
buf ( R_84b_1e094b48 , n49567 );
buf ( R_99e_1e182488 , C0 );
buf ( R_6dc_1dfb6588 , n49568 );
buf ( R_3ad_1d9d6768 , n49574 );
buf ( R_a59_1e189468 , n49580 );
buf ( R_b62_1e6ba368 , C0 );
buf ( R_731_1dfb9aa8 , n49587 );
buf ( R_3f1_1d9d91e8 , n49592 );
buf ( R_620_1dfaf008 , n49593 );
buf ( R_67d_1dfb2a28 , n49601 );
buf ( R_adf_1e6ae888 , n49604 );
buf ( R_349_1d9d28e8 , n49676 );
buf ( R_3d1_1d9d7de8 , n49682 );
buf ( R_3f4_1d9d93c8 , n49683 );
buf ( R_80a_1e0927a8 , C0 );
buf ( R_350_1d9d2d48 , n49684 );
buf ( R_a50_1e188ec8 , n49685 );
buf ( R_bc1_1e6b75c8 , n49692 );
buf ( R_b85_1e6b5048 , n49705 );
buf ( R_5d7_1ddac208 , n49708 );
buf ( R_7a2_1ddada68 , C0 );
buf ( R_539_1dda5f48 , n49724 );
buf ( R_bbc_1e6b72a8 , n49725 );
buf ( R_c14_1e6ba9a8 , n49726 );
buf ( R_6c8_1dfb5908 , n49727 );
buf ( R_4c8_1dda18a8 , n49728 );
buf ( R_360_1d9d3748 , n49729 );
buf ( R_2e2_1d9ced88 , C0 );
buf ( R_936_1e17e388 , C0 );
buf ( R_9f3_1e1854a8 , n49732 );
buf ( R_b25_1e6b1448 , n49747 );
buf ( R_b0a_1e6b0868 , C0 );
buf ( R_b56_1e6b87e8 , C0 );
buf ( R_bf4_1e6b95a8 , n49748 );
buf ( R_95f_1e17f828 , n49751 );
buf ( R_3b5_1d9d6c68 , n49757 );
buf ( R_52a_1dda5fe8 , C0 );
buf ( R_9f2_1e185908 , C0 );
buf ( R_9f4_1e185548 , n49758 );
buf ( R_686_1dfb34c8 , C0 );
buf ( R_2bc_1d9fd068 , n49759 );
buf ( R_7a6_1e08e928 , C0 );
buf ( R_9ef_1e185228 , n49762 );
buf ( R_b1e_1e6b78e8 , C0 );
buf ( R_bfb_1e6b9a08 , n49765 );
buf ( R_378_1d9d4648 , n49766 );
buf ( R_9ee_1e185688 , C0 );
buf ( R_9f0_1e1852c8 , n49767 );
buf ( R_9f5_1e1855e8 , n49837 );
buf ( R_4bd_1dda11c8 , n49843 );
buf ( R_5af_1ddaa908 , n49846 );
buf ( R_822_1e097f28 , C0 );
buf ( R_872_1e0968a8 , C0 );
buf ( R_9f1_1e185368 , n49925 );
buf ( R_337_1d9d1da8 , n49928 );
buf ( R_707_1dfb8068 , n49931 );
buf ( R_755_1dfbb128 , n49936 );
buf ( R_8f9_1e09b808 , n49941 );
buf ( R_432_1d9dbf88 , C0 );
buf ( R_8af_1e0989c8 , n49944 );
buf ( R_bc5_1e6b7848 , n49958 );
buf ( R_934_1e09dce8 , n49959 );
buf ( R_469_1d9ddce8 , n49964 );
buf ( R_572_1dda87e8 , C0 );
buf ( R_863_1e095a48 , n49967 );
buf ( R_958_1e17f3c8 , n49968 );
buf ( R_742_1dfbaa48 , C0 );
buf ( R_2a5_1d9fc208 , n49974 );
buf ( R_a9a_1e18c208 , C0 );
buf ( R_af9_1e6af8c8 , n49979 );
buf ( R_9c1_1e183568 , n49985 );
buf ( R_83c_1e0941e8 , n49986 );
buf ( R_a81_1e18ad68 , n49992 );
buf ( R_c19_1e6bacc8 , n50008 );
buf ( R_91c_1e09cde8 , n50009 );
buf ( R_4ac_1dda0728 , n50010 );
buf ( R_bf8_1e6b9828 , n50011 );
buf ( R_5be_1dda7168 , C0 );
buf ( R_93b_1e17e1a8 , n50014 );
buf ( R_63c_1dfb0188 , n50015 );
buf ( R_7e1_1e090908 , n50020 );
buf ( R_7ba_1e08f5a8 , C0 );
buf ( R_6b2_1dfb5048 , C0 );
buf ( R_4dc_1dda2528 , n50021 );
buf ( R_79e_1e08e428 , C0 );
buf ( R_492_1dd9fbe8 , C0 );
buf ( R_750_1dfbae08 , n50022 );
buf ( R_9d8_1e1843c8 , n50023 );
buf ( R_365_1d9d3a68 , n50071 );
buf ( R_994_1e181948 , n50072 );
buf ( R_95c_1e17f648 , n50073 );
buf ( R_2ff_1d9cfaa8 , n50076 );
buf ( R_89b_1e097d48 , n50079 );
buf ( R_827_1e0934c8 , n50082 );
buf ( R_332_1d9d1f88 , C0 );
buf ( R_9a7_1e182528 , n50085 );
buf ( R_834_1e093ce8 , n50086 );
buf ( R_30b_1d9d0228 , n50089 );
buf ( R_86b_1e095f48 , n50092 );
buf ( R_649_1dfb09a8 , n50098 );
buf ( R_a1d_1e186ee8 , n50172 );
buf ( R_b59_1e6b34c8 , n50192 );
buf ( R_bb3_1e6b6d08 , n50195 );
buf ( R_796_1e08e1a8 , C0 );
buf ( R_941_1e17e568 , n50208 );
buf ( R_be9_1e6b8ec8 , n50220 );
buf ( R_485_1dd9eec8 , n50225 );
buf ( R_317_1d9d09a8 , n50228 );
buf ( R_8a3_1e098248 , n50231 );
buf ( R_49e_1dda0368 , C0 );
buf ( R_9c0_1e1834c8 , n50232 );
buf ( R_32c_1d9d16c8 , n50233 );
buf ( R_6d6_1dfb66c8 , C0 );
buf ( R_a15_1e1869e8 , n50288 );
buf ( R_33e_1d9d2708 , C0 );
buf ( R_38c_1d9d52c8 , n50289 );
buf ( R_75b_1dfbb4e8 , n50292 );
buf ( R_ac4_1e18d748 , n50293 );
buf ( R_5d9_1ddac348 , n50298 );
buf ( R_546_1dda6c68 , C0 );
buf ( R_2be_1d9fd6a8 , C0 );
buf ( R_b76_1e6b4be8 , C0 );
buf ( R_975_1e1805e8 , n50304 );
buf ( R_5c3_1ddab588 , n50307 );
buf ( R_500_1dda3ba8 , n50308 );
buf ( R_889_1e097208 , n50323 );
buf ( R_988_1e1811c8 , n50324 );
buf ( R_c2c_1e6bb8a8 , n50325 );
buf ( R_b98_1e6b5c28 , n50326 );
buf ( R_47d_1dd9e9c8 , n50331 );
buf ( R_417_1d9da9a8 , n50334 );
buf ( R_819_1e092c08 , n50346 );
buf ( R_8f8_1e09b768 , n50347 );
buf ( R_942_1e17eb08 , C0 );
buf ( R_ad1_1e6adfc8 , n50353 );
buf ( R_8ce_1e09a228 , C0 );
buf ( R_563_1dda7988 , n50356 );
buf ( R_2e8_1d9cec48 , n50357 );
buf ( R_838_1e093f68 , n50358 );
buf ( R_aee_1e187c08 , C0 );
buf ( R_641_1dfb04a8 , n50366 );
buf ( R_c16_1e6b41e8 , C0 );
buf ( R_6c3_1dfb55e8 , n50369 );
buf ( R_5f3_1ddad388 , n50372 );
buf ( R_558_1dda72a8 , n50373 );
buf ( R_821_1e093108 , n50378 );
buf ( R_a5f_1e189828 , n50381 );
buf ( R_3cd_1d9d7b68 , n50387 );
buf ( R_80f_1e0925c8 , n50390 );
buf ( R_724_1dfb9288 , n50391 );
buf ( R_848_1e094968 , n50392 );
buf ( R_9bf_1e183428 , n50395 );
buf ( R_a19_1e186c68 , n50446 );
buf ( R_baf_1e6b6a88 , n50449 );
buf ( R_64a_1dfb0f48 , C0 );
buf ( R_aa8_1e18c5c8 , n50450 );
buf ( R_6be_1dfb57c8 , C0 );
buf ( R_481_1dd9ec48 , n50464 );
buf ( R_428_1d9db448 , n50465 );
buf ( R_be6_1e6b91e8 , C0 );
buf ( R_44f_1d9dcca8 , n50468 );
buf ( R_5b4_1ddaac28 , n50469 );
buf ( R_629_1dfaf5a8 , n50475 );
buf ( R_78f_1dfbd568 , n50478 );
buf ( R_91f_1e09cfc8 , n50481 );
buf ( R_858_1e095368 , n50482 );
buf ( R_afb_1e6afa08 , n50485 );
buf ( R_3fb_1d9d9828 , n50488 );
buf ( R_922_1e091628 , C0 );
buf ( R_916_1e09cf28 , C0 );
buf ( R_8a1_1e098108 , n50495 );
buf ( R_8db_1e09a548 , n50498 );
buf ( R_b32_1e6b2168 , C0 );
buf ( R_411_1d9da5e8 , n50503 );
buf ( R_6b0_1dfb4a08 , n50504 );
buf ( R_5d1_1ddabe48 , n50509 );
buf ( R_7df_1e0907c8 , n50512 );
buf ( R_b04_1e6affa8 , n50513 );
buf ( R_45a_1d9dd888 , C0 );
buf ( R_814_1e0928e8 , n50514 );
buf ( R_665_1dfb1b28 , n50521 );
buf ( R_69e_1dfb43c8 , C0 );
buf ( R_b42_1e6b2b68 , C0 );
buf ( R_555_1dda70c8 , n50533 );
buf ( R_374_1d9d43c8 , n50534 );
buf ( R_352_1d9d3388 , C0 );
buf ( R_2a6_1d9fc7a8 , C0 );
buf ( R_756_1dfbb6c8 , C0 );
buf ( R_bd6_1e6b3568 , C0 );
buf ( R_baa_1e18d888 , C0 );
buf ( R_5b9_1ddaaf48 , n50549 );
buf ( R_3ec_1d9d8ec8 , n50550 );
buf ( n275549 , RI21a19c60_2);
not ( n275550 , n275549 );
not ( n275551 , n275550 );
buf ( n275552 , n275551 );
buf ( n275553 , n275552 );
buf ( n275554 , RI21a5daf0_1);
buf ( n275555 , n275554 );
buf ( n275556 , RI2107e620_463);
not ( n275557 , n275556 );
buf ( n275558 , n275557 );
buf ( n275559 , n275558 );
buf ( n275560 , RI210bf4e0_288);
not ( n275561 , n275560 );
not ( n275562 , n275561 );
buf ( n275563 , n275562 );
buf ( n275564 , RI21078b30_503);
not ( n275565 , n275564 );
not ( n275566 , n275565 );
buf ( n275567 , n275566 );
not ( n275568 , n275567 );
xor ( n275569 , n275563 , n275568 );
buf ( n275570 , RI21a13090_74);
buf ( n275571 , n275570 );
buf ( n275572 , n275571 );
xor ( n275573 , n275569 , n275572 );
buf ( n275574 , RI210bf558_287);
not ( n275575 , n275574 );
not ( n275576 , n275575 );
buf ( n275577 , n275576 );
buf ( n275578 , RI21078ba8_502);
not ( n275579 , n275578 );
not ( n275580 , n275579 );
buf ( n275581 , n275580 );
not ( n275582 , n275581 );
xor ( n275583 , n275577 , n275582 );
buf ( n275584 , RI21a13108_73);
buf ( n275585 , n275584 );
buf ( n275586 , n275585 );
and ( n275587 , n275583 , n275586 );
and ( n275588 , n275577 , n275582 );
or ( n275589 , n275587 , n275588 );
nor ( n275590 , n275573 , n275589 );
not ( n275591 , n275590 );
nand ( n275592 , n275573 , n275589 );
nand ( n275593 , n275591 , n275592 );
not ( n275594 , n275593 );
buf ( n275595 , RI21a116c8_87);
buf ( n275596 , n275595 );
buf ( n275597 , n275596 );
buf ( n275598 , RI210bd6e0_301);
not ( n275599 , n275598 );
not ( n275600 , n275599 );
buf ( n275601 , n275600 );
xor ( n275602 , n275597 , n275601 );
buf ( n275603 , RI21077078_516);
not ( n275604 , n275603 );
not ( n275605 , n275604 );
buf ( n275606 , n275605 );
not ( n275607 , n275606 );
xor ( n275608 , n275602 , n275607 );
buf ( n275609 , RI21a11dd0_86);
buf ( n275610 , n275609 );
buf ( n275611 , n275610 );
buf ( n275612 , RI210bd758_300);
not ( n275613 , n275612 );
not ( n275614 , n275613 );
buf ( n275615 , n275614 );
xor ( n275616 , n275611 , n275615 );
buf ( n275617 , RI210770f0_515);
not ( n275618 , n275617 );
not ( n275619 , n275618 );
buf ( n275620 , n275619 );
not ( n275621 , n275620 );
and ( n275622 , n275616 , n275621 );
and ( n275623 , n275611 , n275615 );
or ( n275624 , n275622 , n275623 );
nor ( n275625 , n275608 , n275624 );
xor ( n275626 , n275611 , n275615 );
xor ( n275627 , n275626 , n275621 );
buf ( n275628 , RI21a11e48_85);
buf ( n275629 , n275628 );
buf ( n275630 , n275629 );
buf ( n275631 , RI210bd7d0_299);
not ( n275632 , n275631 );
not ( n275633 , n275632 );
buf ( n275634 , n275633 );
xor ( n275635 , n275630 , n275634 );
buf ( n275636 , RI21077168_514);
not ( n275637 , n275636 );
not ( n275638 , n275637 );
buf ( n275639 , n275638 );
not ( n275640 , n275639 );
and ( n275641 , n275635 , n275640 );
and ( n275642 , n275630 , n275634 );
or ( n275643 , n275641 , n275642 );
nor ( n275644 , n275627 , n275643 );
nor ( n275645 , n275625 , n275644 );
not ( n275646 , n275645 );
buf ( n275647 , RI21a132e8_69);
buf ( n275648 , n275647 );
buf ( n275649 , n275648 );
buf ( n275650 , RI210bff30_283);
not ( n275651 , n275650 );
not ( n275652 , n275651 );
buf ( n275653 , n275652 );
xor ( n275654 , n275649 , n275653 );
buf ( n275655 , RI210797d8_498);
not ( n275656 , n275655 );
not ( n275657 , n275656 );
buf ( n275658 , n275657 );
not ( n275659 , n275658 );
xor ( n275660 , n275654 , n275659 );
xor ( n275661 , n275597 , n275601 );
and ( n275662 , n275661 , n275607 );
and ( n275663 , n275597 , n275601 );
or ( n275664 , n275662 , n275663 );
nor ( n275665 , n275660 , n275664 );
buf ( n275666 , RI210bfeb8_284);
not ( n275667 , n275666 );
not ( n275668 , n275667 );
buf ( n275669 , n275668 );
buf ( n275670 , RI21079760_499);
not ( n275671 , n275670 );
not ( n275672 , n275671 );
buf ( n275673 , n275672 );
not ( n275674 , n275673 );
xor ( n275675 , n275669 , n275674 );
buf ( n275676 , RI21a13270_70);
buf ( n275677 , n275676 );
buf ( n275678 , n275677 );
xor ( n275679 , n275675 , n275678 );
xor ( n275680 , n275649 , n275653 );
and ( n275681 , n275680 , n275659 );
and ( n275682 , n275649 , n275653 );
or ( n275683 , n275681 , n275682 );
nor ( n275684 , n275679 , n275683 );
nor ( n275685 , n275646 , n275665 , n275684 );
not ( n275686 , n275685 );
buf ( n275687 , RI210be1a8_295);
not ( n275688 , n275687 );
not ( n275689 , n275688 );
buf ( n275690 , n275689 );
buf ( n275691 , RI21077d98_510);
not ( n275692 , n275691 );
not ( n275693 , n275692 );
buf ( n275694 , n275693 );
not ( n275695 , n275694 );
xor ( n275696 , n275690 , n275695 );
buf ( n275697 , RI21a12028_81);
buf ( n275698 , n275697 );
buf ( n275699 , n275698 );
xor ( n275700 , n275696 , n275699 );
buf ( n275701 , RI21a12730_80);
buf ( n275702 , n275701 );
buf ( n275703 , n275702 );
buf ( n275704 , RI210bea18_294);
not ( n275705 , n275704 );
not ( n275706 , n275705 );
buf ( n275707 , n275706 );
xor ( n275708 , n275703 , n275707 );
buf ( n275709 , RI21077e10_509);
not ( n275710 , n275709 );
not ( n275711 , n275710 );
buf ( n275712 , n275711 );
not ( n275713 , n275712 );
and ( n275714 , n275708 , n275713 );
and ( n275715 , n275703 , n275707 );
or ( n275716 , n275714 , n275715 );
or ( n275717 , n275700 , n275716 );
not ( n275718 , n275717 );
xor ( n275719 , n275703 , n275707 );
xor ( n275720 , n275719 , n275713 );
buf ( n275721 , RI21a127a8_79);
buf ( n275722 , n275721 );
buf ( n275723 , RI210bea90_293);
not ( n275724 , n275723 );
not ( n275725 , n275724 );
buf ( n275726 , n275725 );
xor ( n275727 , n275722 , n275726 );
buf ( n275728 , RI21077e88_508);
not ( n275729 , n275728 );
not ( n275730 , n275729 );
buf ( n275731 , n275730 );
not ( n275732 , n275731 );
and ( n275733 , n275727 , n275732 );
and ( n275734 , n275722 , n275726 );
or ( n275735 , n275733 , n275734 );
or ( n275736 , n275720 , n275735 );
not ( n275737 , n275736 );
buf ( n275738 , RI21079850_497);
not ( n275739 , n275738 );
not ( n275740 , n275739 );
buf ( n275741 , n275740 );
not ( n275742 , n275741 );
not ( n275743 , n275741 );
buf ( n275744 , RI21a139f0_68);
buf ( n275745 , n275744 );
not ( n275746 , n275745 );
or ( n275747 , n275743 , n275746 );
or ( n275748 , n275741 , n275745 );
buf ( n275749 , RI21084368_418);
buf ( n275750 , n275749 );
buf ( n275751 , n275750 );
nand ( n275752 , n275748 , n275751 );
nand ( n275753 , n275747 , n275752 );
xor ( n275754 , n275742 , n275753 );
xor ( n275755 , n275722 , n275726 );
xor ( n275756 , n275755 , n275732 );
and ( n275757 , n275754 , n275756 );
and ( n275758 , n275742 , n275753 );
or ( n275759 , n275757 , n275758 );
not ( n275760 , n275759 );
or ( n275761 , n275737 , n275760 );
nand ( n275762 , n275720 , n275735 );
nand ( n275763 , n275761 , n275762 );
not ( n275764 , n275763 );
or ( n275765 , n275718 , n275764 );
nand ( n275766 , n275700 , n275716 );
nand ( n275767 , n275765 , n275766 );
buf ( n275768 , RI21a11f38_83);
buf ( n275769 , n275768 );
buf ( n275770 , n275769 );
buf ( n275771 , RI210be0b8_297);
not ( n275772 , n275771 );
not ( n275773 , n275772 );
buf ( n275774 , n275773 );
xor ( n275775 , n275770 , n275774 );
buf ( n275776 , RI21077258_512);
not ( n275777 , n275776 );
not ( n275778 , n275777 );
buf ( n275779 , n275778 );
not ( n275780 , n275779 );
xor ( n275781 , n275775 , n275780 );
buf ( n275782 , RI21a11fb0_82);
buf ( n275783 , n275782 );
buf ( n275784 , n275783 );
buf ( n275785 , RI210be130_296);
not ( n275786 , n275785 );
not ( n275787 , n275786 );
buf ( n275788 , n275787 );
xor ( n275789 , n275784 , n275788 );
buf ( n275790 , RI21077d20_511);
not ( n275791 , n275790 );
not ( n275792 , n275791 );
buf ( n275793 , n275792 );
not ( n275794 , n275793 );
and ( n275795 , n275789 , n275794 );
and ( n275796 , n275784 , n275788 );
or ( n275797 , n275795 , n275796 );
nor ( n275798 , n275781 , n275797 );
xor ( n275799 , n275784 , n275788 );
xor ( n275800 , n275799 , n275794 );
xor ( n275801 , n275690 , n275695 );
and ( n275802 , n275801 , n275699 );
and ( n275803 , n275690 , n275695 );
or ( n275804 , n275802 , n275803 );
nor ( n275805 , n275800 , n275804 );
nor ( n275806 , n275798 , n275805 );
nand ( n275807 , n275767 , n275806 );
xor ( n275808 , n275630 , n275634 );
xor ( n275809 , n275808 , n275640 );
buf ( n275810 , RI210be040_298);
not ( n275811 , n275810 );
not ( n275812 , n275811 );
buf ( n275813 , n275812 );
buf ( n275814 , RI210771e0_513);
not ( n275815 , n275814 );
not ( n275816 , n275815 );
buf ( n275817 , n275816 );
not ( n275818 , n275817 );
xor ( n275819 , n275813 , n275818 );
buf ( n275820 , RI21a11ec0_84);
buf ( n275821 , n275820 );
buf ( n275822 , n275821 );
and ( n275823 , n275819 , n275822 );
and ( n275824 , n275813 , n275818 );
or ( n275825 , n275823 , n275824 );
nor ( n275826 , n275809 , n275825 );
xor ( n275827 , n275813 , n275818 );
xor ( n275828 , n275827 , n275822 );
xor ( n275829 , n275770 , n275774 );
and ( n275830 , n275829 , n275780 );
and ( n275831 , n275770 , n275774 );
or ( n275832 , n275830 , n275831 );
nor ( n275833 , n275828 , n275832 );
nor ( n275834 , n275826 , n275833 );
not ( n275835 , n275834 );
or ( n275836 , n275807 , n275835 );
nand ( n275837 , n275800 , n275804 );
or ( n275838 , n275798 , n275837 );
nand ( n275839 , n275781 , n275797 );
nand ( n275840 , n275838 , n275839 );
and ( n275841 , n275834 , n275840 );
nand ( n275842 , n275828 , n275832 );
or ( n275843 , n275826 , n275842 );
nand ( n275844 , n275809 , n275825 );
nand ( n275845 , n275843 , n275844 );
nor ( n275846 , n275841 , n275845 );
nand ( n275847 , n275836 , n275846 );
not ( n275848 , n275847 );
or ( n275849 , n275686 , n275848 );
nand ( n275850 , n275627 , n275643 );
or ( n275851 , n275625 , n275850 );
nand ( n275852 , n275608 , n275624 );
nand ( n275853 , n275851 , n275852 );
not ( n275854 , n275853 );
or ( n275855 , n275854 , n275665 );
nand ( n275856 , n275660 , n275664 );
nand ( n275857 , n275855 , n275856 );
not ( n275858 , n275684 );
and ( n275859 , n275857 , n275858 );
and ( n275860 , n275679 , n275683 );
nor ( n275861 , n275859 , n275860 );
nand ( n275862 , n275849 , n275861 );
buf ( n275863 , RI21a13180_72);
buf ( n275864 , n275863 );
buf ( n275865 , n275864 );
buf ( n275866 , RI210bfdc8_286);
not ( n275867 , n275866 );
not ( n275868 , n275867 );
buf ( n275869 , n275868 );
xor ( n275870 , n275865 , n275869 );
buf ( n275871 , RI21078c20_501);
not ( n275872 , n275871 );
not ( n275873 , n275872 );
buf ( n275874 , n275873 );
not ( n275875 , n275874 );
xor ( n275876 , n275870 , n275875 );
buf ( n275877 , RI21a131f8_71);
buf ( n275878 , n275877 );
buf ( n275879 , n275878 );
buf ( n275880 , RI210bfe40_285);
not ( n275881 , n275880 );
not ( n275882 , n275881 );
buf ( n275883 , n275882 );
xor ( n275884 , n275879 , n275883 );
buf ( n275885 , RI21078c98_500);
not ( n275886 , n275885 );
not ( n275887 , n275886 );
buf ( n275888 , n275887 );
not ( n275889 , n275888 );
and ( n275890 , n275884 , n275889 );
and ( n275891 , n275879 , n275883 );
or ( n275892 , n275890 , n275891 );
nor ( n275893 , n275876 , n275892 );
xor ( n275894 , n275879 , n275883 );
xor ( n275895 , n275894 , n275889 );
xor ( n275896 , n275669 , n275674 );
and ( n275897 , n275896 , n275678 );
and ( n275898 , n275669 , n275674 );
or ( n275899 , n275897 , n275898 );
nor ( n275900 , n275895 , n275899 );
nor ( n275901 , n275893 , n275900 );
and ( n275902 , n275862 , n275901 );
nand ( n275903 , n275895 , n275899 );
or ( n275904 , n275893 , n275903 );
nand ( n275905 , n275876 , n275892 );
nand ( n275906 , n275904 , n275905 );
nor ( n275907 , n275902 , n275906 );
xor ( n275908 , n275577 , n275582 );
xor ( n275909 , n275908 , n275586 );
xor ( n275910 , n275865 , n275869 );
and ( n275911 , n275910 , n275875 );
and ( n275912 , n275865 , n275869 );
or ( n275913 , n275911 , n275912 );
nor ( n275914 , n275909 , n275913 );
or ( n275915 , n275907 , n275914 );
and ( n275916 , n275909 , n275913 );
not ( n275917 , n275916 );
nand ( n275918 , n275915 , n275917 );
not ( n275919 , n275918 );
or ( n275920 , n275594 , n275919 );
or ( n275921 , n275918 , n275593 );
nand ( n275922 , n275920 , n275921 );
buf ( n275923 , n275922 );
buf ( n275924 , n275923 );
not ( n275925 , n275549 );
not ( n275926 , n275925 );
buf ( n275927 , n275926 );
buf ( n275928 , n275927 );
not ( n275929 , n275549 );
not ( n275930 , n275929 );
buf ( n275931 , n275930 );
buf ( n275932 , n275931 );
buf ( n275933 , RI2107a660_489);
not ( n275934 , n275933 );
not ( n275935 , n275934 );
not ( n275936 , n275935 );
not ( n275937 , n275936 );
buf ( n275938 , n275937 );
buf ( n275939 , RI2107cd48_472);
buf ( n275940 , n275939 );
buf ( n275941 , n275940 );
buf ( n275942 , n275941 );
not ( n275943 , n275942 );
not ( n275944 , n275943 );
buf ( n275945 , RI2106bde0_608);
buf ( n275946 , n275945 );
buf ( n275947 , n275946 );
not ( n275948 , n275947 );
buf ( n275949 , RI2107c118_476);
buf ( n275950 , n275949 );
buf ( n275951 , n275950 );
not ( n275952 , n275951 );
nand ( n275953 , n275948 , n275952 );
buf ( n275954 , RI2107a570_491);
buf ( n275955 , n275954 );
buf ( n275956 , n275955 );
not ( n275957 , n275956 );
buf ( n275958 , RI21079940_495);
buf ( n275959 , n275958 );
buf ( n275960 , n275959 );
not ( n275961 , n275960 );
nand ( n275962 , n275957 , n275961 );
nor ( n275963 , n275953 , n275962 );
buf ( n275964 , RI2107a5e8_490);
buf ( n275965 , n275964 );
buf ( n275966 , n275965 );
buf ( n275967 , RI2107d900_469);
buf ( n275968 , n275967 );
buf ( n275969 , n275968 );
nor ( n275970 , n275966 , n275969 );
buf ( n275971 , RI2107b1a0_487);
buf ( n275972 , n275971 );
buf ( n275973 , n275972 );
buf ( n275974 , RI2107d978_468);
buf ( n275975 , n275974 );
buf ( n275976 , n275975 );
nor ( n275977 , n275973 , n275976 );
nand ( n275978 , n275970 , n275977 );
not ( n275979 , n275978 );
buf ( n275980 , RI2107a480_493);
buf ( n275981 , n275980 );
buf ( n275982 , n275981 );
not ( n275983 , n275982 );
buf ( n275984 , RI2107da68_466);
buf ( n275985 , n275984 );
buf ( n275986 , n275985 );
not ( n275987 , n275986 );
nand ( n275988 , n275983 , n275987 );
buf ( n275989 , RI210799b8_494);
buf ( n275990 , n275989 );
buf ( n275991 , n275990 );
not ( n275992 , n275991 );
buf ( n275993 , RI2107d9f0_467);
buf ( n275994 , n275993 );
buf ( n275995 , n275994 );
not ( n275996 , n275995 );
nand ( n275997 , n275992 , n275996 );
nor ( n275998 , n275988 , n275997 );
buf ( n275999 , RI2107a4f8_492);
buf ( n276000 , n275999 );
buf ( n276001 , n276000 );
not ( n276002 , n276001 );
buf ( n276003 , RI210798c8_496);
buf ( n276004 , n276003 );
buf ( n276005 , n276004 );
not ( n276006 , n276005 );
nand ( n276007 , n276002 , n276006 );
buf ( n276008 , RI2107ce38_470);
buf ( n276009 , n276008 );
buf ( n276010 , n276009 );
not ( n276011 , n276010 );
buf ( n276012 , RI2107cdc0_471);
buf ( n276013 , n276012 );
buf ( n276014 , n276013 );
not ( n276015 , n276014 );
nand ( n276016 , n276011 , n276015 );
nor ( n276017 , n276007 , n276016 );
and ( n276018 , n275963 , n275979 , n275998 , n276017 );
buf ( n276019 , n276018 );
not ( n276020 , n276019 );
not ( n276021 , n276020 );
or ( n276022 , n275944 , n276021 );
not ( n276023 , n276019 );
or ( n276024 , n276023 , n275943 );
nand ( n276025 , n276022 , n276024 );
buf ( n276026 , n276025 );
and ( n276027 , n275938 , n276026 );
not ( n276028 , n275938 );
buf ( n276029 , n275940 );
and ( n276030 , n276028 , n276029 );
nor ( n276031 , n276027 , n276030 );
buf ( n276032 , n276010 );
not ( n276033 , n276032 );
not ( n276034 , n276033 );
not ( n276035 , n275947 );
not ( n276036 , n275973 );
nand ( n276037 , n276035 , n276036 );
not ( n276038 , n275966 );
not ( n276039 , n275951 );
nand ( n276040 , n276038 , n276039 );
nor ( n276041 , n276037 , n276040 );
not ( n276042 , n276001 );
not ( n276043 , n275956 );
nand ( n276044 , n276042 , n276043 );
not ( n276045 , n275982 );
not ( n276046 , n275991 );
nand ( n276047 , n276045 , n276046 );
nor ( n276048 , n276044 , n276047 );
and ( n276049 , n276041 , n276048 );
buf ( n276050 , n276049 );
buf ( n276051 , n276006 );
nand ( n276052 , n276051 , n275961 );
buf ( n276053 , n275996 );
buf ( n276054 , n275987 );
nand ( n276055 , n276053 , n276054 );
nor ( n276056 , n276052 , n276055 );
buf ( n276057 , n275969 );
buf ( n276058 , n275976 );
nor ( n276059 , n276057 , n276058 );
and ( n276060 , n276056 , n276059 );
nand ( n276061 , n276050 , n276060 );
not ( n276062 , n276061 );
or ( n276063 , n276034 , n276062 );
nand ( n276064 , n276050 , n276060 );
or ( n276065 , n276064 , n276033 );
nand ( n276066 , n276063 , n276065 );
buf ( n276067 , n276066 );
buf ( n276068 , n276067 );
not ( n276069 , n276057 );
not ( n276070 , n276069 );
not ( n276071 , n276058 );
and ( n276072 , n276056 , n276071 );
nand ( n276073 , n276050 , n276072 );
not ( n276074 , n276073 );
or ( n276075 , n276070 , n276074 );
nand ( n276076 , n276050 , n276072 );
or ( n276077 , n276076 , n276069 );
nand ( n276078 , n276075 , n276077 );
buf ( n276079 , n276078 );
buf ( n276080 , n276079 );
nor ( n276081 , n276068 , n276080 );
not ( n276082 , n276071 );
buf ( n276083 , n276056 );
nand ( n276084 , n276050 , n276083 );
not ( n276085 , n276084 );
or ( n276086 , n276082 , n276085 );
nand ( n276087 , n276050 , n276083 );
or ( n276088 , n276087 , n276071 );
nand ( n276089 , n276086 , n276088 );
buf ( n276090 , n276089 );
buf ( n276091 , RI2107ccd0_473);
buf ( n276092 , n276091 );
buf ( n276093 , n276092 );
not ( n276094 , n276093 );
not ( n276095 , n276094 );
nand ( n276096 , n276019 , n275943 );
not ( n276097 , n276096 );
or ( n276098 , n276095 , n276097 );
nand ( n276099 , n276019 , n275943 );
or ( n276100 , n276099 , n276094 );
nand ( n276101 , n276098 , n276100 );
buf ( n276102 , n276101 );
nor ( n276103 , n276090 , n276102 );
nand ( n276104 , n276031 , n276081 , n276103 );
not ( n276105 , n276104 );
nor ( n276106 , n275941 , n276093 );
buf ( n276107 , n276106 );
nand ( n276108 , n276019 , n276107 );
buf ( n276109 , RI2107cc58_474);
buf ( n276110 , n276109 );
buf ( n276111 , n276110 );
buf ( n276112 , n276111 );
not ( n276113 , n276112 );
xnor ( n276114 , n276108 , n276113 );
buf ( n276115 , n276114 );
not ( n276116 , n276053 );
not ( n276117 , n276054 );
buf ( n276118 , n276052 );
nor ( n276119 , n276117 , n276118 );
nand ( n276120 , n276050 , n276119 );
not ( n276121 , n276120 );
or ( n276122 , n276116 , n276121 );
or ( n276123 , n276120 , n276053 );
nand ( n276124 , n276122 , n276123 );
buf ( n276125 , n276124 );
nor ( n276126 , n276115 , n276125 );
not ( n276127 , n276126 );
buf ( n276128 , n276015 );
not ( n276129 , n276128 );
not ( n276130 , n276059 );
nor ( n276131 , n276130 , n276032 );
and ( n276132 , n276056 , n276131 );
nand ( n276133 , n276050 , n276132 );
not ( n276134 , n276133 );
or ( n276135 , n276129 , n276134 );
nand ( n276136 , n276050 , n276132 );
or ( n276137 , n276136 , n276128 );
nand ( n276138 , n276135 , n276137 );
buf ( n276139 , n276138 );
buf ( n276140 , n276139 );
nor ( n276141 , n276127 , n276140 );
nand ( n276142 , n276105 , n276141 );
buf ( n276143 , n275935 );
not ( n276144 , n276143 );
buf ( n276145 , RI2107c028_478);
buf ( n276146 , n276145 );
buf ( n276147 , n276146 );
and ( n276148 , n276144 , n276147 );
not ( n276149 , n276144 );
buf ( n276150 , n276146 );
not ( n276151 , n276150 );
not ( n276152 , n276151 );
not ( n276153 , n275998 );
nor ( n276154 , n276153 , n275978 );
not ( n276155 , n276017 );
not ( n276156 , n275962 );
buf ( n276157 , RI2107cbe0_475);
buf ( n276158 , n276157 );
buf ( n276159 , n276158 );
nor ( n276160 , n276111 , n276159 );
nand ( n276161 , n276156 , n276160 );
nor ( n276162 , n276155 , n276161 );
buf ( n276163 , n276035 );
buf ( n276164 , n276039 );
buf ( n276165 , RI2107c0a0_477);
buf ( n276166 , n276165 );
buf ( n276167 , n276166 );
not ( n276168 , n276167 );
buf ( n276169 , n276168 );
nand ( n276170 , n276163 , n276164 , n276169 );
not ( n276171 , n276107 );
nor ( n276172 , n276170 , n276171 );
nand ( n276173 , n276154 , n276162 , n276172 );
not ( n276174 , n276173 );
or ( n276175 , n276152 , n276174 );
or ( n276176 , n276173 , n276151 );
nand ( n276177 , n276175 , n276176 );
buf ( n276178 , n276177 );
and ( n276179 , n276149 , n276178 );
nor ( n276180 , n276148 , n276179 );
buf ( n276181 , n276166 );
and ( n276182 , n276144 , n276181 );
not ( n276183 , n276144 );
not ( n276184 , n276169 );
nand ( n276185 , n276160 , n276106 );
buf ( n276186 , n276185 );
not ( n276187 , n276186 );
nand ( n276188 , n276019 , n276187 );
not ( n276189 , n276188 );
or ( n276190 , n276184 , n276189 );
nand ( n276191 , n276019 , n276187 );
or ( n276192 , n276191 , n276169 );
nand ( n276193 , n276190 , n276192 );
buf ( n276194 , n276193 );
and ( n276195 , n276183 , n276194 );
nor ( n276196 , n276182 , n276195 );
nand ( n276197 , n276180 , n276196 );
not ( n276198 , n276197 );
not ( n276199 , n275938 );
buf ( n276200 , RI2107bfb0_479);
buf ( n276201 , n276200 );
buf ( n276202 , n276201 );
and ( n276203 , n276199 , n276202 );
not ( n276204 , n276199 );
nand ( n276205 , n276151 , n276168 );
buf ( n276206 , n276205 );
nor ( n276207 , n276186 , n276206 );
nand ( n276208 , n276019 , n276207 );
buf ( n276209 , n276201 );
not ( n276210 , n276209 );
buf ( n276211 , n276210 );
not ( n276212 , n276211 );
and ( n276213 , n276208 , n276212 );
not ( n276214 , n276208 );
and ( n276215 , n276214 , n276211 );
nor ( n276216 , n276213 , n276215 );
buf ( n276217 , n276216 );
not ( n276218 , n276217 );
not ( n276219 , n276218 );
and ( n276220 , n276204 , n276219 );
nor ( n276221 , n276203 , n276220 );
nor ( n276222 , n276171 , n276112 );
nand ( n276223 , n276019 , n276222 );
buf ( n276224 , n276159 );
and ( n276225 , n276223 , n276224 );
not ( n276226 , n276223 );
not ( n276227 , n276224 );
and ( n276228 , n276226 , n276227 );
nor ( n276229 , n276225 , n276228 );
buf ( n276230 , n276229 );
not ( n276231 , n276230 );
nand ( n276232 , n276198 , n276221 , n276231 );
nor ( n276233 , n276142 , n276232 );
buf ( n276234 , n276046 );
not ( n276235 , n276234 );
buf ( n276236 , n276041 );
buf ( n276237 , n276044 );
buf ( n276238 , n276045 );
not ( n276239 , n276238 );
nor ( n276240 , n276237 , n276239 );
nand ( n276241 , n276236 , n276240 );
not ( n276242 , n276241 );
or ( n276243 , n276235 , n276242 );
or ( n276244 , n276241 , n276234 );
nand ( n276245 , n276243 , n276244 );
buf ( n276246 , n276245 );
buf ( n276247 , n276246 );
and ( n276248 , n276247 , n275938 );
and ( n276249 , n276144 , n275990 );
nor ( n276250 , n276248 , n276249 );
buf ( n276251 , n276042 );
not ( n276252 , n276251 );
buf ( n276253 , n276043 );
nand ( n276254 , n276236 , n276253 );
not ( n276255 , n276254 );
or ( n276256 , n276252 , n276255 );
or ( n276257 , n276254 , n276251 );
nand ( n276258 , n276256 , n276257 );
buf ( n276259 , n276258 );
buf ( n276260 , n276259 );
and ( n276261 , n276260 , n275938 );
and ( n276262 , n276144 , n276000 );
nor ( n276263 , n276261 , n276262 );
not ( n276264 , n276253 );
not ( n276265 , n276264 );
not ( n276266 , n276236 );
or ( n276267 , n276265 , n276266 );
or ( n276268 , n276236 , n276264 );
nand ( n276269 , n276267 , n276268 );
buf ( n276270 , n276269 );
and ( n276271 , n275935 , n276270 );
not ( n276272 , n275935 );
buf ( n276273 , n275955 );
and ( n276274 , n276272 , n276273 );
nor ( n276275 , n276271 , n276274 );
not ( n276276 , n275935 );
buf ( n276277 , n276036 );
not ( n276278 , n276277 );
buf ( n276279 , n275953 );
not ( n276280 , n276279 );
or ( n276281 , n276278 , n276280 );
not ( n276282 , n276277 );
not ( n276283 , n276282 );
or ( n276284 , n276279 , n276283 );
nand ( n276285 , n276281 , n276284 );
buf ( n276286 , n276285 );
not ( n276287 , n276286 );
or ( n276288 , n276276 , n276287 );
not ( n276289 , n275935 );
buf ( n276290 , n275972 );
nand ( n276291 , n276289 , n276290 );
nand ( n276292 , n276288 , n276291 );
not ( n276293 , n275935 );
not ( n276294 , n276164 );
not ( n276295 , n276163 );
and ( n276296 , n276294 , n276295 );
not ( n276297 , n276294 );
and ( n276298 , n276297 , n276163 );
nor ( n276299 , n276296 , n276298 );
buf ( n276300 , n276299 );
not ( n276301 , n276300 );
or ( n276302 , n276293 , n276301 );
not ( n276303 , n275935 );
buf ( n276304 , n275950 );
nand ( n276305 , n276303 , n276304 );
nand ( n276306 , n276302 , n276305 );
nor ( n276307 , n276292 , n276306 );
nand ( n276308 , n276275 , n276307 );
not ( n276309 , n276308 );
not ( n276310 , n276143 );
not ( n276311 , n276038 );
not ( n276312 , n276311 );
nor ( n276313 , n276279 , n276282 );
not ( n276314 , n276313 );
or ( n276315 , n276312 , n276314 );
or ( n276316 , n276311 , n276313 );
nand ( n276317 , n276315 , n276316 );
buf ( n276318 , n276317 );
not ( n276319 , n276318 );
or ( n276320 , n276310 , n276319 );
buf ( n276321 , n275965 );
nand ( n276322 , n275936 , n276321 );
nand ( n276323 , n276320 , n276322 );
buf ( n276324 , n275946 );
buf ( n276325 , n276324 );
nor ( n276326 , n276323 , n276325 );
and ( n276327 , n276250 , n276263 , n276309 , n276326 );
not ( n276328 , n276054 );
not ( n276329 , n276118 );
nand ( n276330 , n276050 , n276329 );
not ( n276331 , n276330 );
or ( n276332 , n276328 , n276331 );
nand ( n276333 , n276050 , n276329 );
or ( n276334 , n276333 , n276054 );
nand ( n276335 , n276332 , n276334 );
buf ( n276336 , n276335 );
buf ( n276337 , n276336 );
not ( n276338 , n276051 );
not ( n276339 , n276049 );
not ( n276340 , n276339 );
buf ( n276341 , n275961 );
nand ( n276342 , n276340 , n276341 );
not ( n276343 , n276342 );
or ( n276344 , n276338 , n276343 );
or ( n276345 , n276051 , n276342 );
nand ( n276346 , n276344 , n276345 );
buf ( n276347 , n276346 );
buf ( n276348 , n276347 );
nor ( n276349 , n276337 , n276348 );
not ( n276350 , n276341 );
not ( n276351 , n276339 );
or ( n276352 , n276350 , n276351 );
not ( n276353 , n276050 );
or ( n276354 , n276353 , n276341 );
nand ( n276355 , n276352 , n276354 );
buf ( n276356 , n276355 );
and ( n276357 , n276356 , n275937 );
not ( n276358 , n275959 );
nor ( n276359 , n276358 , n275937 );
nor ( n276360 , n276357 , n276359 );
buf ( n276361 , n276360 );
buf ( n276362 , n275981 );
and ( n276363 , n275936 , n276362 );
not ( n276364 , n275936 );
not ( n276365 , n276238 );
not ( n276366 , n276237 );
nand ( n276367 , n276236 , n276366 );
not ( n276368 , n276367 );
or ( n276369 , n276365 , n276368 );
or ( n276370 , n276238 , n276367 );
nand ( n276371 , n276369 , n276370 );
buf ( n276372 , n276371 );
and ( n276373 , n276364 , n276372 );
nor ( n276374 , n276363 , n276373 );
buf ( n276375 , n276374 );
nand ( n276376 , n276327 , n276349 , n276361 , n276375 );
buf ( n276377 , RI2107b3f8_482);
buf ( n276378 , n276377 );
buf ( n276379 , n276378 );
not ( n276380 , n276379 );
not ( n276381 , n276380 );
not ( n276382 , n276185 );
buf ( n276383 , RI2107bf38_480);
buf ( n276384 , n276383 );
buf ( n276385 , n276384 );
not ( n276386 , n276385 );
nand ( n276387 , n276210 , n276386 );
nor ( n276388 , n276205 , n276387 );
nand ( n276389 , n276382 , n276388 );
buf ( n276390 , RI2107bec0_481);
buf ( n276391 , n276390 );
buf ( n276392 , n276391 );
buf ( n276393 , n276392 );
nor ( n276394 , n276389 , n276393 );
nand ( n276395 , n276394 , n276019 );
not ( n276396 , n276395 );
or ( n276397 , n276381 , n276396 );
not ( n276398 , n276389 );
not ( n276399 , n276393 );
nand ( n276400 , n276019 , n276398 , n276399 );
or ( n276401 , n276400 , n276380 );
nand ( n276402 , n276397 , n276401 );
buf ( n276403 , n276402 );
buf ( n276404 , n276403 );
not ( n276405 , n276399 );
nand ( n276406 , n276019 , n276398 );
not ( n276407 , n276406 );
or ( n276408 , n276405 , n276407 );
or ( n276409 , n276406 , n276399 );
nand ( n276410 , n276408 , n276409 );
buf ( n276411 , n276410 );
buf ( n276412 , n276411 );
nor ( n276413 , n276404 , n276412 );
not ( n276414 , n276392 );
nand ( n276415 , n276414 , n276380 );
nor ( n276416 , n276389 , n276415 );
nand ( n276417 , n276019 , n276416 );
buf ( n276418 , RI2107b380_483);
buf ( n276419 , n276418 );
buf ( n276420 , n276419 );
buf ( n276421 , n276420 );
and ( n276422 , n276417 , n276421 );
not ( n276423 , n276417 );
not ( n276424 , n276421 );
and ( n276425 , n276423 , n276424 );
nor ( n276426 , n276422 , n276425 );
buf ( n276427 , n276426 );
not ( n276428 , n276427 );
not ( n276429 , n276428 );
buf ( n276430 , n276143 );
nand ( n276431 , n276429 , n276430 );
not ( n276432 , n276206 );
nand ( n276433 , n276432 , n276210 );
nor ( n276434 , n276186 , n276433 );
nand ( n276435 , n276019 , n276434 );
buf ( n276436 , n276386 );
not ( n276437 , n276436 );
and ( n276438 , n276435 , n276437 );
not ( n276439 , n276435 );
and ( n276440 , n276439 , n276436 );
nor ( n276441 , n276438 , n276440 );
buf ( n276442 , n276441 );
not ( n276443 , n276442 );
not ( n276444 , n276443 );
buf ( n276445 , n276143 );
nand ( n276446 , n276444 , n276445 );
nand ( n276447 , n276413 , n276431 , n276446 );
nor ( n276448 , n276376 , n276447 );
and ( n276449 , n276233 , n276448 );
buf ( n276450 , n276019 );
not ( n276451 , n276398 );
nor ( n276452 , n276379 , n276392 );
buf ( n276453 , RI2107b308_484);
buf ( n276454 , n276453 );
buf ( n276455 , n276454 );
nor ( n276456 , n276455 , n276420 );
nand ( n276457 , n276452 , n276456 );
not ( n276458 , n276457 );
buf ( n276459 , RI2107b218_486);
buf ( n276460 , n276459 );
buf ( n276461 , n276460 );
not ( n276462 , n276461 );
buf ( n276463 , RI2107b290_485);
buf ( n276464 , n276463 );
buf ( n276465 , n276464 );
not ( n276466 , n276465 );
nand ( n276467 , n276462 , n276466 );
buf ( n276468 , RI2107a6d8_488);
buf ( n276469 , n276468 );
buf ( n276470 , n276469 );
nor ( n9008 , n276467 , n276470 );
nand ( n9009 , n276458 , n9008 );
nor ( n9010 , n276451 , n9009 );
nand ( n9011 , n276450 , n9010 );
buf ( n9012 , n275935 );
buf ( n9013 , n9012 );
and ( n9014 , n9011 , n9013 );
not ( n9015 , n9011 );
not ( n9016 , n9013 );
and ( n9017 , n9015 , n9016 );
nor ( n9018 , n9014 , n9017 );
buf ( n9019 , n9018 );
nand ( n9020 , n9019 , n276445 );
not ( n9021 , n9020 );
not ( n9022 , n9021 );
nor ( n9023 , n276449 , n9022 );
buf ( n9024 , n9023 );
not ( n9025 , n276445 );
not ( n9026 , n276455 );
not ( n9027 , n9026 );
nor ( n9028 , n276415 , n276420 );
not ( n9029 , n9028 );
nor ( n9030 , n9029 , n276389 );
nand ( n9031 , n276019 , n9030 );
not ( n9032 , n9031 );
or ( n9033 , n9027 , n9032 );
or ( n9034 , n9031 , n9026 );
nand ( n9035 , n9033 , n9034 );
buf ( n9036 , n9035 );
not ( n9037 , n9036 );
or ( n9038 , n9025 , n9037 );
not ( n9039 , n276445 );
nand ( n9040 , n9039 , n276454 );
nand ( n9041 , n9038 , n9040 );
buf ( n9042 , n9041 );
buf ( n9043 , n9042 );
nand ( n9044 , n9024 , n9043 );
nor ( n9045 , n276389 , n276457 );
nand ( n9046 , n276019 , n9045 );
and ( n9047 , n9046 , n276465 );
not ( n9048 , n9046 );
and ( n9049 , n9048 , n276466 );
nor ( n9050 , n9047 , n9049 );
buf ( n9051 , n9050 );
buf ( n9052 , n9051 );
not ( n9053 , n275938 );
not ( n9054 , n9053 );
and ( n9055 , n9052 , n9054 );
not ( n9056 , n276430 );
and ( n9057 , n9056 , n276464 );
nor ( n9058 , n9055 , n9057 );
and ( n9059 , n9044 , n9058 );
not ( n9060 , n9044 );
not ( n9061 , n9058 );
and ( n9062 , n9060 , n9061 );
nor ( n9063 , n9059 , n9062 );
not ( n9064 , n276445 );
not ( n9065 , n276412 );
or ( n9066 , n9064 , n9065 );
nand ( n9067 , n9039 , n276391 );
nand ( n9068 , n9066 , n9067 );
not ( n9069 , n276384 );
not ( n9070 , n9056 );
or ( n9071 , n9069 , n9070 );
nand ( n9072 , n9071 , n276446 );
and ( n9073 , n9068 , n9072 );
not ( n9074 , n276430 );
not ( n9075 , n276404 );
or ( n9076 , n9074 , n9075 );
nand ( n9077 , n9039 , n276378 );
nand ( n9078 , n9076 , n9077 );
nand ( n9079 , n9073 , n9078 );
not ( n9080 , n276419 );
not ( n9081 , n9053 );
or ( n9082 , n9080 , n9081 );
nand ( n9083 , n9082 , n276431 );
not ( n9084 , n9083 );
and ( n9085 , n9079 , n9084 );
not ( n9086 , n9079 );
and ( n9087 , n9086 , n9083 );
nor ( n9088 , n9085 , n9087 );
not ( n9089 , n9073 );
not ( n9090 , n9078 );
and ( n9091 , n9089 , n9090 );
not ( n9092 , n9089 );
and ( n9093 , n9092 , n9078 );
nor ( n9094 , n9091 , n9093 );
not ( n9095 , n9068 );
and ( n9096 , n9072 , n9095 );
not ( n9097 , n9072 );
and ( n9098 , n9097 , n9068 );
or ( n9099 , n9096 , n9098 );
and ( n9100 , n9088 , n9094 , n9099 );
not ( n9101 , n9100 );
nand ( n9102 , n9063 , n9101 );
not ( n9103 , n9102 );
not ( n9104 , n276376 );
not ( n9105 , n9104 );
not ( n9106 , n276142 );
not ( n9107 , n9106 );
or ( n9108 , n9105 , n9107 );
not ( n9109 , n9022 );
nand ( n9110 , n9108 , n9109 );
not ( n9111 , n276231 );
nand ( n9112 , n9111 , n276445 );
nand ( n9113 , n9056 , n276158 );
and ( n9114 , n9112 , n9113 );
nor ( n9115 , n9110 , n9114 );
buf ( n9116 , n276196 );
not ( n9117 , n9116 );
nand ( n9118 , n9115 , n9117 );
not ( n9119 , n9118 );
not ( n9120 , n276180 );
buf ( n9121 , n9120 );
nand ( n9122 , n9119 , n9121 );
not ( n9123 , n276221 );
buf ( n9124 , n9123 );
and ( n9125 , n9122 , n9124 );
not ( n9126 , n9122 );
not ( n9127 , n9124 );
and ( n9128 , n9126 , n9127 );
nor ( n9129 , n9125 , n9128 );
not ( n9130 , n9129 );
not ( n9131 , n9121 );
and ( n9132 , n9118 , n9131 );
not ( n9133 , n9118 );
and ( n9134 , n9133 , n9121 );
nor ( n9135 , n9132 , n9134 );
not ( n9136 , n9135 );
not ( n9137 , n9114 );
not ( n9138 , n9137 );
buf ( n9139 , n9110 );
not ( n9140 , n9139 );
not ( n9141 , n9140 );
not ( n9142 , n9141 );
or ( n9143 , n9138 , n9142 );
not ( n9144 , n9137 );
nand ( n9145 , n9140 , n9144 );
nand ( n9146 , n9143 , n9145 );
nor ( n9147 , n9136 , n9146 );
nand ( n9148 , n9130 , n9147 );
not ( n9149 , n9148 );
not ( n9150 , n9115 );
xor ( n9151 , n9117 , n9150 );
buf ( n9152 , n9151 );
nand ( n9153 , n9149 , n9152 );
buf ( n9154 , n9153 );
not ( n9155 , n9154 );
buf ( n9156 , RI2106be58_607);
not ( n9157 , n9156 );
not ( n9158 , n9157 );
buf ( n9159 , n9158 );
nand ( n9160 , n9103 , n9155 , n9159 );
buf ( n9161 , RI2107dae0_465);
not ( n9162 , n9161 );
not ( n9163 , n9162 );
nand ( n9164 , n9160 , n9163 );
nand ( n9165 , n276233 , n276448 );
nand ( n9166 , n9165 , n9021 );
nor ( n9167 , n9166 , n9043 );
not ( n9168 , n9167 );
nand ( n9169 , n9166 , n9042 );
buf ( n9170 , n9169 );
nand ( n9171 , n9168 , n9170 );
nand ( n9172 , n9171 , n9163 );
and ( n9173 , n9164 , n9172 );
not ( n9174 , n9021 );
not ( n9175 , n276232 );
or ( n9176 , n9174 , n9175 );
nand ( n9177 , n9176 , n9139 );
buf ( n9178 , n9072 );
and ( n9179 , n9177 , n9178 );
not ( n9180 , n9177 );
not ( n9181 , n9178 );
and ( n9182 , n9180 , n9181 );
nor ( n9183 , n9179 , n9182 );
and ( n9184 , n9183 , n9159 );
nor ( n9185 , n9173 , n9184 );
not ( n9186 , n9185 );
not ( n9187 , n9183 );
not ( n9188 , n9149 );
or ( n9189 , n9187 , n9188 );
nor ( n9190 , n276102 , n9036 );
not ( n9191 , n276139 );
and ( n9192 , n276126 , n9190 , n9191 );
nor ( n9193 , n276090 , n276336 );
not ( n9194 , n276325 );
and ( n9195 , n276360 , n9194 );
nor ( n9196 , n276411 , n276308 );
and ( n9197 , n276026 , n276143 );
nor ( n9198 , n9197 , n276323 );
nand ( n9199 , n9193 , n9195 , n9196 , n9198 );
not ( n9200 , n9199 );
not ( n9201 , n9051 );
nor ( n9202 , n276246 , n276259 );
and ( n9203 , n276374 , n9202 );
nand ( n9204 , n9201 , n9203 , n276231 );
nor ( n9205 , n276197 , n9204 );
nor ( n9206 , n276403 , n276079 );
nor ( n9207 , n276067 , n276347 );
nand ( n9208 , n9206 , n9207 );
nand ( n9209 , n276218 , n276428 , n276443 );
nor ( n9210 , n9208 , n9209 );
nand ( n9211 , n9192 , n9200 , n9205 , n9210 );
nand ( n9212 , n9211 , n9021 );
nand ( n9213 , n276458 , n276466 );
nor ( n9214 , n276451 , n9213 );
nand ( n9215 , n276450 , n9214 );
not ( n9216 , n276462 );
and ( n9217 , n9215 , n9216 );
not ( n9218 , n9215 );
and ( n9219 , n9218 , n276462 );
nor ( n9220 , n9217 , n9219 );
buf ( n9221 , n9220 );
and ( n9222 , n9221 , n276445 );
and ( n9223 , n276144 , n276460 );
nor ( n9224 , n9222 , n9223 );
buf ( n9225 , n9224 );
and ( n9226 , n9212 , n9225 );
not ( n9227 , n9212 );
not ( n9228 , n9225 );
and ( n9229 , n9227 , n9228 );
nor ( n9230 , n9226 , n9229 );
buf ( n9231 , n9230 );
nor ( n9232 , n9224 , n9020 );
nand ( n9233 , n9211 , n9232 );
not ( n9234 , n9233 );
not ( n9235 , n276467 );
nand ( n9236 , n9235 , n276458 );
nor ( n9237 , n276451 , n9236 );
nand ( n9238 , n276450 , n9237 );
xor ( n9239 , n9238 , n276470 );
buf ( n9240 , n9239 );
not ( n9241 , n9053 );
nand ( n9242 , n9240 , n9241 );
nand ( n9243 , n9053 , n276469 );
nand ( n9244 , n9242 , n9243 );
not ( n9245 , n9244 );
and ( n9246 , n9234 , n9245 );
and ( n9247 , n9233 , n9244 );
nor ( n9248 , n9246 , n9247 );
buf ( n9249 , n9248 );
and ( n9250 , n9231 , n9249 );
buf ( n9251 , n9250 );
buf ( n9252 , RI2106ddc0_566);
not ( n9253 , n9252 );
not ( n9254 , n9253 );
nand ( n9255 , n9251 , n9254 );
not ( n9256 , n9231 );
and ( n9257 , n9256 , n9249 );
buf ( n9258 , n9257 );
buf ( n9259 , n9258 );
buf ( n9260 , RI210730b8_542);
not ( n9261 , n9260 );
not ( n9262 , n9261 );
nand ( n9263 , n9259 , n9262 );
not ( n9264 , n9248 );
not ( n9265 , n9264 );
not ( n9266 , n9265 );
nand ( n9267 , n9266 , n9256 );
not ( n9268 , n9267 );
buf ( n9269 , RI2106cc68_590);
not ( n9270 , n9269 );
not ( n9271 , n9270 );
nand ( n9272 , n9268 , n9271 );
buf ( n9273 , RI2106a2b0_640);
buf ( n9274 , n9273 );
not ( n9275 , n9274 );
buf ( n9276 , RI21069ab8_644);
buf ( n9277 , n9276 );
not ( n9278 , n9277 );
buf ( n9279 , RI2106bfc0_604);
not ( n9280 , n9279 );
not ( n9281 , n9280 );
not ( n9282 , n9281 );
buf ( n9283 , RI2106c038_603);
not ( n9284 , n9283 );
not ( n9285 , n9284 );
buf ( n9286 , RI2106a148_643);
buf ( n9287 , n9286 );
nor ( n9288 , n9285 , n9287 );
nand ( n9289 , n9282 , n9288 );
buf ( n9290 , RI2106bf48_605);
buf ( n9291 , n9290 );
nor ( n9292 , n9289 , n9291 );
nand ( n9293 , n9278 , n9292 );
buf ( n9294 , RI21069a40_645);
buf ( n9295 , n9294 );
not ( n9296 , n9295 );
buf ( n9297 , RI2106a760_630);
buf ( n9298 , n9297 );
buf ( n9299 , RI2106a5f8_633);
buf ( n9300 , n9299 );
nor ( n9301 , n9298 , n9300 );
buf ( n9302 , RI2106a670_632);
buf ( n9303 , n9302 );
buf ( n9304 , RI2106bed0_606);
not ( n9305 , n9304 );
not ( n9306 , n9305 );
nor ( n9307 , n9303 , n9306 );
and ( n9308 , n9301 , n9307 );
buf ( n9309 , RI2106a7d8_629);
buf ( n9310 , n9309 );
buf ( n9311 , RI2106c308_597);
buf ( n9312 , n9311 );
nor ( n9313 , n9310 , n9312 );
buf ( n9314 , RI2106ae68_628);
buf ( n9315 , n9314 );
buf ( n9316 , RI2106a6e8_631);
buf ( n9317 , n9316 );
nor ( n9318 , n9315 , n9317 );
and ( n9319 , n9313 , n9318 );
nand ( n9320 , n9296 , n9308 , n9319 );
nor ( n9321 , n9293 , n9320 );
buf ( n9322 , RI2106a580_634);
buf ( n9323 , n9322 );
not ( n9324 , n9323 );
and ( n9325 , n9321 , n9324 );
buf ( n9326 , RI2106a508_635);
buf ( n9327 , n9326 );
buf ( n9328 , RI2106a490_636);
buf ( n9329 , n9328 );
nor ( n9330 , n9327 , n9329 );
nand ( n9331 , n9325 , n9330 );
buf ( n9332 , RI2106a3a0_638);
buf ( n9333 , n9332 );
nor ( n9334 , n9331 , n9333 );
buf ( n9335 , RI2106a328_639);
buf ( n9336 , n9335 );
not ( n9337 , n9336 );
and ( n9338 , n9334 , n9337 );
nand ( n9339 , n9275 , n9338 );
buf ( n9340 , RI2106a238_641);
buf ( n9341 , n9340 );
nor ( n9342 , n9339 , n9341 );
buf ( n9343 , RI2106c290_598);
not ( n9344 , n9343 );
not ( n9345 , n9344 );
not ( n9346 , n9345 );
and ( n9347 , n9342 , n9346 );
buf ( n9348 , RI2106c218_599);
not ( n9349 , n9348 );
not ( n9350 , n9349 );
not ( n9351 , n9350 );
nand ( n9352 , n9347 , n9351 );
buf ( n9353 , RI2106c1a0_600);
not ( n9354 , n9353 );
not ( n9355 , n9354 );
nor ( n9356 , n9352 , n9355 );
not ( n9357 , n9356 );
buf ( n9358 , RI2106c128_601);
not ( n9359 , n9358 );
not ( n9360 , n9359 );
nor ( n9361 , n9357 , n9360 );
buf ( n9362 , RI2106c0b0_602);
not ( n9363 , n9362 );
not ( n9364 , n9363 );
not ( n9365 , n9364 );
nand ( n9366 , n9361 , n9365 );
not ( n9367 , n9366 );
not ( n9368 , n9231 );
buf ( n9369 , n9244 );
not ( n9370 , n9369 );
nor ( n9371 , n9368 , n9370 );
buf ( n9372 , n9371 );
nand ( n9373 , n9367 , n9372 );
nand ( n9374 , n9255 , n9263 , n9272 , n9373 );
buf ( n9375 , RI2106dd48_567);
not ( n9376 , n9375 );
not ( n9377 , n9376 );
not ( n9378 , n9377 );
not ( n9379 , n9231 );
not ( n9380 , n9379 );
not ( n9381 , n9380 );
or ( n9382 , n9378 , n9381 );
not ( n9383 , n9231 );
not ( n9384 , n9383 );
buf ( n9385 , RI21073040_543);
not ( n9386 , n9385 );
not ( n9387 , n9386 );
not ( n9388 , n9387 );
or ( n9389 , n9384 , n9388 );
nand ( n9390 , n9382 , n9389 );
not ( n9391 , n9249 );
not ( n9392 , n9391 );
and ( n9393 , n9390 , n9392 );
not ( n9394 , n9267 );
buf ( n9395 , RI2106cbf0_591);
not ( n9396 , n9395 );
not ( n9397 , n9396 );
and ( n9398 , n9394 , n9397 );
nor ( n9399 , n9393 , n9398 );
nand ( n9400 , n9399 , n9373 );
nand ( n9401 , n9374 , n9400 );
not ( n9402 , n9401 );
buf ( n9403 , n9402 );
not ( n9404 , n9058 );
not ( n9405 , n9041 );
and ( n9406 , n9404 , n9405 );
and ( n9407 , n9023 , n9058 );
nor ( n9408 , n9406 , n9407 );
nand ( n9409 , n9408 , n9169 );
buf ( n9410 , n9409 );
buf ( n9411 , n9410 );
buf ( n9412 , RI21a12820_78);
buf ( n9413 , n9412 );
not ( n9414 , n9413 );
buf ( n9415 , RI210beb08_292);
buf ( n9416 , n9415 );
not ( n9417 , n9416 );
buf ( n9418 , RI21a0e608_121);
buf ( n9419 , n9418 );
not ( n9420 , n9419 );
buf ( n9421 , RI21077f00_507);
not ( n9422 , n9421 );
not ( n9423 , n9422 );
nand ( n9424 , n9414 , n9417 , n9420 , n9423 );
buf ( n9425 , RI210b87a8_334);
buf ( n9426 , n9425 );
nor ( n9427 , n9423 , n9426 );
nand ( n9428 , n9427 , n9416 , n9413 );
nand ( n9429 , n9424 , n9428 );
not ( n9430 , n9429 );
not ( n9431 , n9430 );
not ( n9432 , n9431 );
not ( n9433 , n9432 );
not ( n9434 , n9433 );
buf ( n9435 , RI21a11560_90);
buf ( n9436 , n9435 );
buf ( n9437 , n9436 );
not ( n9438 , n9437 );
buf ( n9439 , RI210bcd80_304);
buf ( n9440 , n9439 );
buf ( n9441 , n9440 );
nand ( n9442 , n9438 , n9441 );
not ( n9443 , n9442 );
buf ( n9444 , RI210cfcc8_237);
buf ( n9445 , n9444 );
buf ( n9446 , n9445 );
not ( n9447 , n9446 );
buf ( n9448 , RI210842f0_419);
buf ( n9449 , n9448 );
buf ( n9450 , n9449 );
nand ( n9451 , n9447 , n9450 );
not ( n9452 , n9451 );
or ( n9453 , n9443 , n9452 );
or ( n9454 , n9450 , n9447 );
nand ( n9455 , n9453 , n9454 );
not ( n9456 , n9455 );
buf ( n9457 , RI21a0efe0_114);
buf ( n9458 , n9457 );
buf ( n9459 , n9458 );
not ( n9460 , n9459 );
buf ( n9461 , RI210b92e8_327);
buf ( n9462 , n9461 );
buf ( n9463 , n9462 );
nand ( n9464 , n9460 , n9463 );
buf ( n9465 , RI21a0f148_111);
buf ( n9466 , n9465 );
buf ( n9467 , n9466 );
not ( n9468 , n9467 );
buf ( n9469 , RI21084278_420);
buf ( n9470 , n9469 );
buf ( n9471 , n9470 );
nand ( n9472 , n9468 , n9471 );
and ( n9473 , n9464 , n9472 );
not ( n9474 , n9473 );
or ( n9475 , n9456 , n9474 );
not ( n9476 , n9467 );
nor ( n9477 , n9476 , n9471 );
not ( n9478 , n9477 );
not ( n9479 , n9464 );
or ( n9480 , n9478 , n9479 );
not ( n9481 , n9463 );
buf ( n9482 , n9459 );
nand ( n9483 , n9481 , n9482 );
nand ( n9484 , n9480 , n9483 );
not ( n9485 , n9484 );
nand ( n9486 , n9475 , n9485 );
buf ( n9487 , RI21a0ef68_115);
buf ( n9488 , n9487 );
buf ( n9489 , n9488 );
not ( n9490 , n9489 );
buf ( n9491 , RI210b9270_328);
buf ( n9492 , n9491 );
buf ( n9493 , n9492 );
nand ( n9494 , n9490 , n9493 );
buf ( n9495 , RI21a0eef0_116);
buf ( n9496 , n9495 );
buf ( n9497 , n9496 );
not ( n9498 , n9497 );
buf ( n9499 , RI210b91f8_329);
buf ( n9500 , n9499 );
buf ( n9501 , n9500 );
nand ( n9502 , n9498 , n9501 );
and ( n9503 , n9494 , n9502 );
buf ( n9504 , RI21a0e680_120);
buf ( n9505 , n9504 );
buf ( n9506 , n9505 );
not ( n9507 , n9506 );
buf ( n9508 , RI210b8820_333);
buf ( n9509 , n9508 );
buf ( n9510 , n9509 );
nand ( n9511 , n9507 , n9510 );
buf ( n9512 , RI21a0e6f8_119);
buf ( n9513 , n9512 );
buf ( n9514 , n9513 );
not ( n9515 , n9514 );
buf ( n9516 , RI210b8898_332);
buf ( n9517 , n9516 );
buf ( n9518 , n9517 );
nand ( n9519 , n9515 , n9518 );
and ( n9520 , n9511 , n9519 );
nand ( n9521 , n9503 , n9520 );
buf ( n9522 , RI21a10c00_96);
buf ( n9523 , n9522 );
buf ( n9524 , n9523 );
not ( n9525 , n9524 );
buf ( n9526 , RI210bc2b8_310);
buf ( n9527 , n9526 );
buf ( n9528 , n9527 );
nand ( n9529 , n9525 , n9528 );
buf ( n9530 , RI21a11470_92);
buf ( n9531 , n9530 );
buf ( n9532 , n9531 );
not ( n9533 , n9532 );
buf ( n9534 , RI210bcc90_306);
buf ( n9535 , n9534 );
buf ( n9536 , n9535 );
nand ( n9537 , n9533 , n9536 );
nand ( n9538 , n9529 , n9537 );
buf ( n9539 , RI21a10cf0_94);
buf ( n9540 , n9539 );
buf ( n9541 , n9540 );
not ( n9542 , n9541 );
buf ( n9543 , RI210bc3a8_308);
buf ( n9544 , n9543 );
buf ( n9545 , n9544 );
nand ( n9546 , n9542 , n9545 );
buf ( n9547 , RI21a0e770_118);
buf ( n9548 , n9547 );
buf ( n9549 , n9548 );
not ( n9550 , n9549 );
buf ( n9551 , RI210b8910_331);
buf ( n9552 , n9551 );
buf ( n9553 , n9552 );
nand ( n9554 , n9550 , n9553 );
nand ( n9555 , n9546 , n9554 );
nor ( n9556 , n9538 , n9555 );
buf ( n9557 , RI21a10c78_95);
buf ( n9558 , n9557 );
buf ( n9559 , n9558 );
not ( n9560 , n9559 );
buf ( n9561 , RI210bc330_309);
buf ( n9562 , n9561 );
buf ( n9563 , n9562 );
nand ( n9564 , n9560 , n9563 );
buf ( n9565 , RI21a114e8_91);
buf ( n9566 , n9565 );
buf ( n9567 , n9566 );
not ( n9568 , n9567 );
buf ( n9569 , RI210bcd08_305);
buf ( n9570 , n9569 );
buf ( n9571 , n9570 );
nand ( n9572 , n9568 , n9571 );
nand ( n9573 , n9564 , n9572 );
buf ( n9574 , RI21a10d68_93);
buf ( n9575 , n9574 );
buf ( n9576 , n9575 );
not ( n9577 , n9576 );
buf ( n9578 , RI210bc420_307);
buf ( n9579 , n9578 );
buf ( n9580 , n9579 );
nand ( n9581 , n9577 , n9580 );
buf ( n9582 , RI21a0e7e8_117);
buf ( n9583 , n9582 );
buf ( n9584 , n9583 );
not ( n9585 , n9584 );
buf ( n9586 , RI210b9180_330);
buf ( n9587 , n9586 );
buf ( n9588 , n9587 );
nand ( n9589 , n9585 , n9588 );
nand ( n9590 , n9581 , n9589 );
nor ( n9591 , n9573 , n9590 );
nand ( n9592 , n9556 , n9591 );
nor ( n9593 , n9521 , n9592 );
nand ( n9594 , n9486 , n9593 );
and ( n9595 , n9537 , n9572 );
and ( n9596 , n9529 , n9564 );
and ( n9597 , n9546 , n9581 );
nand ( n9598 , n9595 , n9520 , n9596 , n9597 );
not ( n9599 , n9598 );
not ( n9600 , n9554 );
not ( n9601 , n9584 );
nor ( n9602 , n9601 , n9588 );
not ( n9603 , n9602 );
or ( n9604 , n9600 , n9603 );
not ( n9605 , n9553 );
nand ( n9606 , n9605 , n9549 );
nand ( n9607 , n9604 , n9606 );
not ( n9608 , n9607 );
nand ( n9609 , n9554 , n9589 );
nand ( n9610 , n9608 , n9609 );
not ( n9611 , n9502 );
not ( n9612 , n9489 );
nor ( n9613 , n9612 , n9493 );
not ( n9614 , n9613 );
or ( n9615 , n9611 , n9614 );
not ( n9616 , n9501 );
nand ( n9617 , n9616 , n9497 );
nand ( n9618 , n9615 , n9617 );
not ( n9619 , n9618 );
nand ( n9620 , n9608 , n9619 );
nand ( n9621 , n9599 , n9610 , n9620 );
not ( n9622 , n9511 );
not ( n9623 , n9514 );
nor ( n9624 , n9623 , n9518 );
not ( n9625 , n9624 );
or ( n9626 , n9622 , n9625 );
or ( n9627 , n9510 , n9507 );
nand ( n9628 , n9626 , n9627 );
not ( n9629 , n9628 );
not ( n9630 , n9595 );
or ( n9631 , n9629 , n9630 );
not ( n9632 , n9567 );
buf ( n9633 , n9571 );
nor ( n9634 , n9632 , n9633 );
and ( n9635 , n9634 , n9537 );
not ( n9636 , n9532 );
nor ( n9637 , n9636 , n9536 );
nor ( n9638 , n9635 , n9637 );
nand ( n9639 , n9631 , n9638 );
not ( n9640 , n9596 );
not ( n9641 , n9597 );
nor ( n9642 , n9640 , n9641 );
nand ( n9643 , n9639 , n9642 );
not ( n9644 , n9596 );
not ( n9645 , n9546 );
not ( n9646 , n9576 );
nor ( n9647 , n9646 , n9580 );
not ( n9648 , n9647 );
or ( n9649 , n9645 , n9648 );
not ( n9650 , n9545 );
nand ( n9651 , n9650 , n9541 );
nand ( n9652 , n9649 , n9651 );
not ( n9653 , n9652 );
or ( n9654 , n9644 , n9653 );
buf ( n9655 , n9563 );
nor ( n9656 , n9560 , n9655 );
and ( n9657 , n9656 , n9529 );
not ( n9658 , n9524 );
nor ( n9659 , n9658 , n9528 );
nor ( n9660 , n9657 , n9659 );
nand ( n9661 , n9654 , n9660 );
not ( n9662 , n9661 );
nand ( n9663 , n9594 , n9621 , n9643 , n9662 );
buf ( n9664 , n9663 );
not ( n9665 , n9664 );
buf ( n9666 , RI21a102a0_102);
buf ( n9667 , n9666 );
buf ( n9668 , n9667 );
not ( n9669 , n9668 );
buf ( n9670 , RI210baff8_316);
buf ( n9671 , n9670 );
buf ( n9672 , n9671 );
nand ( n9673 , n9669 , n9672 );
buf ( n9674 , RI21a10318_101);
buf ( n9675 , n9674 );
buf ( n9676 , n9675 );
not ( n9677 , n9676 );
buf ( n9678 , RI210bb070_315);
buf ( n9679 , n9678 );
buf ( n9680 , n9679 );
nand ( n9681 , n9677 , n9680 );
nand ( n9682 , n9673 , n9681 );
buf ( n9683 , RI21a101b0_104);
buf ( n9684 , n9683 );
buf ( n9685 , n9684 );
not ( n9686 , n9685 );
buf ( n9687 , RI210baf08_318);
buf ( n9688 , n9687 );
buf ( n9689 , n9688 );
nand ( n9690 , n9686 , n9689 );
buf ( n9691 , RI21a10228_103);
buf ( n9692 , n9691 );
buf ( n9693 , n9692 );
not ( n9694 , n9693 );
buf ( n9695 , RI210baf80_317);
buf ( n9696 , n9695 );
buf ( n9697 , n9696 );
nand ( n9698 , n9694 , n9697 );
nand ( n9699 , n9690 , n9698 );
nor ( n9700 , n9682 , n9699 );
buf ( n9701 , RI21a10390_100);
buf ( n9702 , n9701 );
buf ( n9703 , n9702 );
not ( n9704 , n9703 );
buf ( n9705 , RI210bb8e0_314);
buf ( n9706 , n9705 );
buf ( n9707 , n9706 );
nand ( n9708 , n9704 , n9707 );
buf ( n9709 , RI21a10408_99);
buf ( n9710 , n9709 );
buf ( n9711 , n9710 );
not ( n9712 , n9711 );
buf ( n9713 , RI210bb958_313);
buf ( n9714 , n9713 );
buf ( n9715 , n9714 );
nand ( n9716 , n9712 , n9715 );
and ( n9717 , n9708 , n9716 );
not ( n9718 , n9717 );
buf ( n9719 , RI21a10b10_98);
buf ( n9720 , n9719 );
buf ( n9721 , n9720 );
not ( n9722 , n9721 );
buf ( n9723 , RI210bb9d0_312);
buf ( n9724 , n9723 );
buf ( n9725 , n9724 );
nand ( n9726 , n9722 , n9725 );
buf ( n9727 , RI21a10b88_97);
buf ( n9728 , n9727 );
buf ( n9729 , n9728 );
not ( n9730 , n9729 );
buf ( n9731 , RI210bba48_311);
buf ( n9732 , n9731 );
buf ( n9733 , n9732 );
nand ( n9734 , n9730 , n9733 );
nand ( n9735 , n9726 , n9734 );
nor ( n9736 , n9718 , n9735 );
nand ( n9737 , n9700 , n9736 );
not ( n9738 , n9737 );
buf ( n9739 , RI21a0f940_108);
buf ( n9740 , n9739 );
buf ( n9741 , n9740 );
not ( n9742 , n9741 );
buf ( n9743 , RI210ba530_322);
buf ( n9744 , n9743 );
buf ( n9745 , n9744 );
nand ( n9746 , n9742 , n9745 );
buf ( n9747 , RI21a0f9b8_107);
buf ( n9748 , n9747 );
buf ( n9749 , n9748 );
not ( n9750 , n9749 );
buf ( n9751 , RI210ba5a8_321);
buf ( n9752 , n9751 );
buf ( n9753 , n9752 );
nand ( n9754 , n9750 , n9753 );
and ( n9755 , n9746 , n9754 );
buf ( n9756 , RI21a0fa30_106);
buf ( n9757 , n9756 );
buf ( n9758 , n9757 );
not ( n9759 , n9758 );
buf ( n9760 , RI210ba620_320);
buf ( n9761 , n9760 );
buf ( n9762 , n9761 );
nand ( n9763 , n9759 , n9762 );
buf ( n9764 , RI21a0faa8_105);
buf ( n9765 , n9764 );
buf ( n9766 , n9765 );
not ( n9767 , n9766 );
buf ( n9768 , RI210ba698_319);
buf ( n9769 , n9768 );
buf ( n9770 , n9769 );
nand ( n9771 , n9767 , n9770 );
and ( n9772 , n9763 , n9771 );
nand ( n9773 , n9755 , n9772 );
buf ( n9774 , RI21a0f850_110);
buf ( n9775 , n9774 );
buf ( n9776 , n9775 );
not ( n9777 , n9776 );
buf ( n9778 , RI210b9c48_324);
buf ( n9779 , n9778 );
buf ( n9780 , n9779 );
nand ( n9781 , n9777 , n9780 );
buf ( n9782 , RI21a0f8c8_109);
buf ( n9783 , n9782 );
buf ( n9784 , n9783 );
not ( n9785 , n9784 );
buf ( n9786 , RI210b9cc0_323);
buf ( n9787 , n9786 );
buf ( n9788 , n9787 );
nand ( n9789 , n9785 , n9788 );
nand ( n9790 , n9781 , n9789 );
nor ( n9791 , n9773 , n9790 );
nand ( n9792 , n9738 , n9791 );
or ( n9793 , n9665 , n9792 );
not ( n9794 , n9700 );
not ( n9795 , n9726 );
not ( n9796 , n9729 );
nor ( n9797 , n9796 , n9733 );
not ( n9798 , n9797 );
or ( n9799 , n9795 , n9798 );
not ( n9800 , n9725 );
nand ( n9801 , n9800 , n9721 );
nand ( n9802 , n9799 , n9801 );
not ( n9803 , n9802 );
not ( n9804 , n9717 );
or ( n9805 , n9803 , n9804 );
not ( n9806 , n9711 );
nor ( n9807 , n9806 , n9715 );
not ( n9808 , n9807 );
not ( n9809 , n9708 );
or ( n277273 , n9808 , n9809 );
not ( n277274 , n9707 );
nand ( n277275 , n277274 , n9703 );
nand ( n277276 , n277273 , n277275 );
not ( n277277 , n277276 );
nand ( n277278 , n9805 , n277277 );
not ( n277279 , n277278 );
or ( n277280 , n9794 , n277279 );
not ( n277281 , n9676 );
nor ( n277282 , n277281 , n9680 );
not ( n277283 , n277282 );
not ( n277284 , n9673 );
or ( n277285 , n277283 , n277284 );
not ( n277286 , n9672 );
nand ( n277287 , n277286 , n9668 );
nand ( n277288 , n277285 , n277287 );
not ( n277289 , n9699 );
and ( n277290 , n277288 , n277289 );
not ( n277291 , n9693 );
nor ( n277292 , n277291 , n9697 );
nand ( n277293 , n277292 , n9690 );
not ( n277294 , n9689 );
nand ( n277295 , n277294 , n9685 );
nand ( n277296 , n277293 , n277295 );
nor ( n277297 , n277290 , n277296 );
nand ( n277298 , n277280 , n277297 );
and ( n277299 , n277298 , n9791 );
not ( n277300 , n9763 );
not ( n277301 , n9766 );
nor ( n277302 , n277301 , n9770 );
not ( n277303 , n277302 );
or ( n277304 , n277300 , n277303 );
not ( n277305 , n9762 );
nand ( n277306 , n277305 , n9758 );
nand ( n277307 , n277304 , n277306 );
not ( n277308 , n277307 );
not ( n277309 , n9755 );
or ( n277310 , n277308 , n277309 );
not ( n277311 , n9749 );
nor ( n277312 , n277311 , n9753 );
not ( n277313 , n277312 );
not ( n277314 , n9746 );
or ( n277315 , n277313 , n277314 );
not ( n277316 , n9745 );
nand ( n277317 , n277316 , n9741 );
nand ( n277318 , n277315 , n277317 );
not ( n277319 , n277318 );
nand ( n277320 , n277310 , n277319 );
not ( n277321 , n277320 );
or ( n277322 , n277321 , n9790 );
not ( n277323 , n9784 );
nor ( n277324 , n277323 , n9788 );
not ( n277325 , n277324 );
not ( n277326 , n9781 );
or ( n277327 , n277325 , n277326 );
not ( n277328 , n9780 );
nand ( n277329 , n277328 , n9776 );
nand ( n277330 , n277327 , n277329 );
not ( n277331 , n277330 );
nand ( n277332 , n277322 , n277331 );
nor ( n277333 , n277299 , n277332 );
nand ( n277334 , n9793 , n277333 );
buf ( n277335 , RI21a0f0d0_112);
buf ( n277336 , n277335 );
buf ( n277337 , n277336 );
not ( n277338 , n277337 );
buf ( n277339 , RI210b9bd0_325);
buf ( n277340 , n277339 );
buf ( n277341 , n277340 );
nand ( n277342 , n277338 , n277341 );
not ( n277343 , n277341 );
nand ( n277344 , n277343 , n277337 );
nand ( n277345 , n277342 , n277344 );
xnor ( n277346 , n277334 , n277345 );
buf ( n277347 , n277346 );
not ( n277348 , n277347 );
or ( n277349 , n9434 , n277348 );
not ( n277350 , n9429 );
not ( n277351 , n277350 );
not ( n277352 , n277351 );
buf ( n277353 , RI21a19990_4);
nand ( n277354 , n277352 , n277353 );
nand ( n277355 , n277349 , n277354 );
and ( n277356 , n9411 , n277355 );
buf ( n277357 , n277356 );
not ( n277358 , n277357 );
nor ( n277359 , n9403 , n277358 );
nor ( n277360 , n9361 , n9365 );
not ( n277361 , n277360 );
nand ( n277362 , n277361 , n9366 );
and ( n277363 , n277362 , n9372 );
not ( n277364 , n9249 );
and ( n277365 , n9379 , n277364 );
not ( n277366 , n277365 );
buf ( n277367 , RI2106cd58_588);
not ( n277368 , n277367 );
not ( n277369 , n277368 );
not ( n277370 , n277369 );
nor ( n277371 , n277366 , n277370 );
nor ( n277372 , n277363 , n277371 );
buf ( n277373 , n9251 );
buf ( n277374 , RI2106deb0_564);
not ( n277375 , n277374 );
not ( n277376 , n277375 );
and ( n277377 , n277373 , n277376 );
not ( n277378 , n9258 );
buf ( n277379 , RI21073c70_539);
not ( n277380 , n277379 );
not ( n277381 , n277380 );
not ( n277382 , n277381 );
nor ( n277383 , n277378 , n277382 );
nor ( n277384 , n277377 , n277383 );
nand ( n277385 , n277372 , n277384 );
buf ( n277386 , n277385 );
buf ( n277387 , n277386 );
not ( n277388 , n277387 );
buf ( n277389 , n9410 );
not ( n277390 , n9430 );
not ( n277391 , n277390 );
not ( n277392 , n9789 );
or ( n277393 , n277324 , n277392 );
not ( n277394 , n277393 );
not ( n277395 , n9773 );
nand ( n277396 , n9738 , n277395 );
or ( n277397 , n9665 , n277396 );
nand ( n277398 , n277298 , n277395 );
and ( n277399 , n277398 , n277321 );
nand ( n277400 , n277397 , n277399 );
not ( n277401 , n277400 );
or ( n277402 , n277394 , n277401 );
or ( n277403 , n277400 , n277393 );
nand ( n277404 , n277402 , n277403 );
buf ( n277405 , n277404 );
not ( n277406 , n277405 );
or ( n277407 , n277391 , n277406 );
buf ( n277408 , RI21a198a0_6);
nand ( n277409 , n9432 , n277408 );
nand ( n277410 , n277407 , n277409 );
and ( n277411 , n277389 , n277410 );
buf ( n277412 , n277411 );
nand ( n277413 , n277388 , n277412 );
buf ( n277414 , RI2106de38_565);
not ( n277415 , n277414 );
not ( n277416 , n277415 );
nand ( n277417 , n277373 , n277416 );
buf ( n277418 , RI21073bf8_540);
not ( n277419 , n277418 );
not ( n277420 , n277419 );
nand ( n277421 , n9259 , n277420 );
buf ( n277422 , RI2106cce0_589);
not ( n277423 , n277422 );
not ( n277424 , n277423 );
nand ( n277425 , n9268 , n277424 );
nand ( n277426 , n9373 , n277417 , n277421 , n277425 );
buf ( n277427 , n277426 );
not ( n277428 , n277427 );
not ( n277429 , n9433 );
nor ( n277430 , n9773 , n277392 );
and ( n277431 , n9738 , n277430 );
not ( n277432 , n277431 );
not ( n277433 , n9664 );
or ( n277434 , n277432 , n277433 );
and ( n277435 , n277298 , n277430 );
or ( n277436 , n277321 , n277392 );
not ( n277437 , n277324 );
nand ( n277438 , n277436 , n277437 );
nor ( n277439 , n277435 , n277438 );
nand ( n277440 , n277434 , n277439 );
nand ( n277441 , n9781 , n277329 );
not ( n277442 , n277441 );
and ( n277443 , n277440 , n277442 );
not ( n277444 , n277440 );
and ( n277445 , n277444 , n277441 );
nor ( n277446 , n277443 , n277445 );
buf ( n277447 , n277446 );
not ( n277448 , n277447 );
or ( n277449 , n277429 , n277448 );
buf ( n277450 , RI21a19918_5);
nand ( n277451 , n9432 , n277450 );
nand ( n277452 , n277449 , n277451 );
and ( n277453 , n277389 , n277452 );
buf ( n277454 , n277453 );
nand ( n277455 , n277428 , n277454 );
buf ( n277456 , RI21a0f058_113);
buf ( n277457 , n277456 );
buf ( n277458 , n277457 );
buf ( n277459 , RI210b9b58_326);
buf ( n277460 , n277459 );
buf ( n277461 , n277460 );
xnor ( n277462 , n277458 , n277461 );
not ( n277463 , n277462 );
not ( n277464 , n9594 );
nand ( n277465 , n9621 , n9643 , n9662 );
nor ( n277466 , n277464 , n277465 );
nor ( n277467 , n277466 , n9737 );
not ( n277468 , n277298 );
not ( n277469 , n277342 );
nor ( n277470 , n277469 , n9790 );
not ( n277471 , n277470 );
not ( n277472 , n277320 );
or ( n277473 , n277471 , n277472 );
not ( n277474 , n277342 );
not ( n277475 , n277330 );
or ( n277476 , n277474 , n277475 );
nand ( n277477 , n277476 , n277344 );
not ( n277478 , n277477 );
nand ( n277479 , n277473 , n277478 );
not ( n277480 , n277479 );
nand ( n277481 , n277468 , n277480 );
or ( n277482 , n277467 , n277481 );
not ( n277483 , n277395 );
not ( n277484 , n277470 );
or ( n277485 , n277483 , n277484 );
nand ( n277486 , n277485 , n277480 );
nand ( n277487 , n277482 , n277486 );
not ( n277488 , n277487 );
or ( n277489 , n277463 , n277488 );
or ( n277490 , n277487 , n277462 );
nand ( n277491 , n277489 , n277490 );
buf ( n277492 , n277491 );
not ( n277493 , n277492 );
or ( n277494 , n277493 , n9432 );
buf ( n277495 , RI21a19a08_3);
nand ( n277496 , n9432 , n277495 );
nand ( n277497 , n277494 , n277496 );
and ( n277498 , n277389 , n277497 );
buf ( n277499 , n277498 );
not ( n277500 , n277499 );
buf ( n277501 , n9400 );
buf ( n277502 , n277501 );
nand ( n277503 , n277500 , n277502 );
nand ( n277504 , n277413 , n277455 , n277503 );
nor ( n277505 , n277359 , n277504 );
not ( n277506 , n9754 );
or ( n277507 , n277312 , n277506 );
not ( n277508 , n277507 );
not ( n277509 , n9772 );
nor ( n277510 , n277509 , n9737 );
not ( n277511 , n277510 );
not ( n277512 , n9664 );
or ( n277513 , n277511 , n277512 );
not ( n277514 , n9772 );
not ( n277515 , n277298 );
or ( n277516 , n277514 , n277515 );
not ( n277517 , n277307 );
nand ( n277518 , n277516 , n277517 );
not ( n277519 , n277518 );
nand ( n277520 , n277513 , n277519 );
not ( n277521 , n277520 );
or ( n277522 , n277508 , n277521 );
or ( n277523 , n277520 , n277507 );
nand ( n277524 , n277522 , n277523 );
buf ( n277525 , n277524 );
not ( n277526 , n277525 );
not ( n277527 , n277390 );
or ( n277528 , n277526 , n277527 );
buf ( n277529 , RI21a197b0_8);
nand ( n277530 , n277527 , n277529 );
nand ( n277531 , n277528 , n277530 );
nand ( n277532 , n9411 , n277531 );
not ( n277533 , n277532 );
buf ( n277534 , n277533 );
not ( n277535 , n277534 );
not ( n277536 , n9267 );
buf ( n277537 , RI2106ce48_586);
not ( n277538 , n277537 );
not ( n277539 , n277538 );
and ( n277540 , n277536 , n277539 );
not ( n277541 , n9372 );
nand ( n277542 , n9352 , n9355 );
not ( n277543 , n277542 );
nor ( n277544 , n277543 , n9356 );
nor ( n277545 , n277541 , n277544 );
nor ( n277546 , n277540 , n277545 );
buf ( n277547 , RI21073d60_537);
buf ( n277548 , n277547 );
nand ( n277549 , n9258 , n277548 );
buf ( n277550 , RI2106dfa0_562);
buf ( n277551 , n277550 );
nand ( n277552 , n9251 , n277551 );
nand ( n277553 , n277546 , n277549 , n277552 );
buf ( n277554 , n277553 );
buf ( n277555 , n277554 );
not ( n277556 , n277555 );
not ( n277557 , n277556 );
or ( n277558 , n277535 , n277557 );
buf ( n277559 , RI2106df28_563);
not ( n277560 , n277559 );
not ( n277561 , n277560 );
nand ( n277562 , n9251 , n277561 );
buf ( n277563 , RI2106cdd0_587);
not ( n277564 , n277563 );
not ( n277565 , n277564 );
nand ( n277566 , n277536 , n277565 );
buf ( n277567 , RI21073ce8_538);
not ( n277568 , n277567 );
not ( n277569 , n277568 );
nand ( n277570 , n9258 , n277569 );
not ( n277571 , n9360 );
nor ( n277572 , n277571 , n9356 );
or ( n277573 , n277572 , n9361 );
nand ( n277574 , n9372 , n277573 );
nand ( n277575 , n277562 , n277566 , n277570 , n277574 );
buf ( n277576 , n277575 );
not ( n277577 , n277576 );
nand ( n277578 , n9746 , n277317 );
not ( n277579 , n277578 );
not ( n277580 , n9772 );
nor ( n277581 , n277580 , n277506 );
not ( n277582 , n277581 );
nor ( n277583 , n277582 , n9737 );
not ( n277584 , n277583 );
not ( n277585 , n9664 );
or ( n277586 , n277584 , n277585 );
not ( n277587 , n277581 );
not ( n277588 , n277298 );
or ( n277589 , n277587 , n277588 );
not ( n277590 , n277517 );
not ( n277591 , n277506 );
and ( n277592 , n277590 , n277591 );
nor ( n277593 , n277592 , n277312 );
nand ( n277594 , n277589 , n277593 );
not ( n277595 , n277594 );
nand ( n277596 , n277586 , n277595 );
not ( n277597 , n277596 );
or ( n277598 , n277579 , n277597 );
or ( n277599 , n277596 , n277578 );
nand ( n277600 , n277598 , n277599 );
buf ( n277601 , n277600 );
not ( n277602 , n277601 );
buf ( n277603 , n277350 );
or ( n277604 , n277602 , n277603 );
buf ( n277605 , RI21a19828_7);
nand ( n277606 , n277527 , n277605 );
nand ( n277607 , n277604 , n277606 );
nand ( n277608 , n277389 , n277607 );
not ( n277609 , n277608 );
buf ( n277610 , n277609 );
nand ( n277611 , n277577 , n277610 );
nand ( n277612 , n277558 , n277611 );
buf ( n277613 , RI2106cec0_585);
not ( n277614 , n277613 );
not ( n277615 , n277614 );
nand ( n277616 , n277365 , n277615 );
buf ( n277617 , RI21073dd8_536);
buf ( n277618 , n277617 );
nand ( n277619 , n9258 , n277618 );
buf ( n277620 , RI2106e018_561);
buf ( n277621 , n277620 );
nand ( n277622 , n9251 , n277621 );
nor ( n277623 , n9347 , n9351 );
not ( n277624 , n277623 );
nand ( n277625 , n277624 , n9352 );
nand ( n277626 , n9372 , n277625 );
nand ( n277627 , n277616 , n277619 , n277622 , n277626 );
buf ( n277628 , n277627 );
buf ( n277629 , n277628 );
not ( n277630 , n277629 );
not ( n277631 , n277390 );
nand ( n277632 , n9738 , n9771 );
or ( n277633 , n9665 , n277632 );
not ( n277634 , n9771 );
not ( n277635 , n277298 );
or ( n277636 , n277634 , n277635 );
not ( n277637 , n277302 );
nand ( n277638 , n277636 , n277637 );
not ( n277639 , n277638 );
nand ( n277640 , n277633 , n277639 );
nand ( n277641 , n9763 , n277306 );
xnor ( n277642 , n277640 , n277641 );
buf ( n277643 , n277642 );
not ( n277644 , n277643 );
or ( n277645 , n277631 , n277644 );
buf ( n277646 , RI21a190a8_9);
nand ( n277647 , n277603 , n277646 );
nand ( n277648 , n277645 , n277647 );
and ( n277649 , n277389 , n277648 );
buf ( n277650 , n277649 );
nand ( n277651 , n277630 , n277650 );
buf ( n277652 , RI210748a0_535);
buf ( n277653 , n277652 );
not ( n277654 , n277653 );
not ( n277655 , n9258 );
or ( n277656 , n277654 , n277655 );
buf ( n277657 , RI2106e090_560);
buf ( n277658 , n277657 );
nand ( n277659 , n9251 , n277658 );
nand ( n277660 , n277656 , n277659 );
buf ( n277661 , RI2106cf38_584);
not ( n277662 , n277661 );
not ( n277663 , n277662 );
not ( n277664 , n277663 );
not ( n277665 , n9268 );
or ( n277666 , n277664 , n277665 );
not ( n277667 , n9345 );
not ( n277668 , n9342 );
not ( n277669 , n277668 );
or ( n277670 , n277667 , n277669 );
not ( n277671 , n9347 );
nand ( n277672 , n277670 , n277671 );
nand ( n277673 , n9372 , n277672 );
nand ( n277674 , n277666 , n277673 );
nor ( n277675 , n277660 , n277674 );
not ( n277676 , n277675 );
buf ( n277677 , n277676 );
not ( n277678 , n277677 );
nand ( n277679 , n9771 , n277637 );
not ( n277680 , n277679 );
not ( n277681 , n9738 );
not ( n277682 , n9664 );
or ( n277683 , n277681 , n277682 );
nand ( n277684 , n277683 , n277468 );
not ( n277685 , n277684 );
or ( n277686 , n277680 , n277685 );
or ( n277687 , n277684 , n277679 );
nand ( n277688 , n277686 , n277687 );
buf ( n277689 , n277688 );
not ( n277690 , n277689 );
or ( n277691 , n277690 , n277603 );
buf ( n277692 , RI21a19030_10);
nand ( n277693 , n9432 , n277692 );
nand ( n277694 , n277691 , n277693 );
nand ( n277695 , n9411 , n277694 );
not ( n277696 , n277695 );
buf ( n277697 , n277696 );
nand ( n277698 , n277678 , n277697 );
nand ( n277699 , n277651 , n277698 );
nor ( n277700 , n277612 , n277699 );
and ( n277701 , n277505 , n277700 );
buf ( n277702 , RI2106cfb0_583);
not ( n277703 , n277702 );
not ( n277704 , n277703 );
nand ( n277705 , n277536 , n277704 );
buf ( n277706 , RI21074918_534);
buf ( n277707 , n277706 );
nand ( n277708 , n9258 , n277707 );
buf ( n277709 , RI2106e108_559);
buf ( n277710 , n277709 );
nand ( n277711 , n9251 , n277710 );
not ( n277712 , n9341 );
not ( n277713 , n9339 );
or ( n277714 , n277712 , n277713 );
nand ( n277715 , n277714 , n277668 );
nand ( n277716 , n9372 , n277715 );
nand ( n277717 , n277705 , n277708 , n277711 , n277716 );
not ( n277718 , n277717 );
not ( n277719 , n277718 );
buf ( n277720 , n277719 );
not ( n277721 , n277720 );
nand ( n277722 , n9690 , n277295 );
not ( n277723 , n277722 );
not ( n277724 , n9682 );
and ( n277725 , n277724 , n9698 );
and ( n277726 , n277725 , n9736 );
not ( n277727 , n277726 );
not ( n277728 , n9664 );
or ( n277729 , n277727 , n277728 );
and ( n277730 , n277278 , n277725 );
not ( n277731 , n9698 );
not ( n277732 , n277288 );
or ( n277733 , n277731 , n277732 );
not ( n277734 , n277292 );
nand ( n277735 , n277733 , n277734 );
nor ( n277736 , n277730 , n277735 );
nand ( n277737 , n277729 , n277736 );
not ( n277738 , n277737 );
or ( n277739 , n277723 , n277738 );
or ( n277740 , n277737 , n277722 );
nand ( n277741 , n277739 , n277740 );
buf ( n277742 , n277741 );
not ( n277743 , n277742 );
or ( n277744 , n277743 , n277603 );
buf ( n277745 , RI21a18fb8_11);
nand ( n277746 , n9432 , n277745 );
nand ( n277747 , n277744 , n277746 );
nand ( n277748 , n277389 , n277747 );
not ( n277749 , n277748 );
buf ( n277750 , n277749 );
nand ( n277751 , n277721 , n277750 );
buf ( n277752 , RI21074990_533);
buf ( n277753 , n277752 );
not ( n277754 , n277753 );
not ( n277755 , n9258 );
or ( n277756 , n277754 , n277755 );
buf ( n277757 , RI21070a48_558);
buf ( n277758 , n277757 );
nand ( n277759 , n9251 , n277758 );
nand ( n277760 , n277756 , n277759 );
buf ( n277761 , RI2106d028_582);
not ( n277762 , n277761 );
not ( n277763 , n277762 );
not ( n277764 , n277763 );
not ( n277765 , n277365 );
or ( n277766 , n277764 , n277765 );
not ( n277767 , n9274 );
not ( n277768 , n9338 );
not ( n277769 , n277768 );
or ( n277770 , n277767 , n277769 );
nand ( n277771 , n277770 , n9339 );
nand ( n277772 , n9372 , n277771 );
nand ( n277773 , n277766 , n277772 );
nor ( n277774 , n277760 , n277773 );
not ( n277775 , n277774 );
buf ( n277776 , n277775 );
not ( n277777 , n277776 );
nand ( n277778 , n9698 , n277734 );
not ( n277779 , n277778 );
and ( n277780 , n9736 , n277724 );
not ( n277781 , n277780 );
not ( n277782 , n9664 );
or ( n277783 , n277781 , n277782 );
and ( n277784 , n277278 , n277724 );
nor ( n277785 , n277784 , n277288 );
nand ( n277786 , n277783 , n277785 );
not ( n277787 , n277786 );
or ( n277788 , n277779 , n277787 );
or ( n277789 , n277786 , n277778 );
nand ( n277790 , n277788 , n277789 );
buf ( n277791 , n277790 );
not ( n277792 , n277791 );
or ( n277793 , n277792 , n277352 );
buf ( n277794 , RI21a18f40_12);
nand ( n277795 , n9432 , n277794 );
nand ( n277796 , n277793 , n277795 );
nand ( n277797 , n9411 , n277796 );
not ( n277798 , n277797 );
buf ( n277799 , n277798 );
nand ( n277800 , n277777 , n277799 );
nand ( n277801 , n277751 , n277800 );
not ( n277802 , n277282 );
nand ( n277803 , n277802 , n9681 );
not ( n277804 , n277803 );
not ( n277805 , n9736 );
not ( n277806 , n9664 );
or ( n277807 , n277805 , n277806 );
not ( n277808 , n277278 );
nand ( n277809 , n277807 , n277808 );
not ( n277810 , n277809 );
or ( n277811 , n277804 , n277810 );
or ( n277812 , n277809 , n277803 );
nand ( n277813 , n277811 , n277812 );
buf ( n277814 , n277813 );
not ( n277815 , n277814 );
or ( n277816 , n277815 , n277352 );
not ( n277817 , n9431 );
buf ( n277818 , RI21a18e50_14);
nand ( n277819 , n277817 , n277818 );
nand ( n277820 , n277816 , n277819 );
nand ( n277821 , n277389 , n277820 );
not ( n277822 , n277821 );
buf ( n277823 , n277822 );
not ( n277824 , n277823 );
buf ( n277825 , RI2106d118_580);
not ( n277826 , n277825 );
not ( n277827 , n277826 );
nand ( n277828 , n277536 , n277827 );
buf ( n277829 , RI21074a80_531);
buf ( n277830 , n277829 );
nand ( n277831 , n9258 , n277830 );
buf ( n277832 , RI21071588_556);
buf ( n277833 , n277832 );
nand ( n277834 , n9251 , n277833 );
not ( n277835 , n9333 );
not ( n277836 , n9331 );
or ( n277837 , n277835 , n277836 );
not ( n277838 , n9334 );
nand ( n277839 , n277837 , n277838 );
nand ( n277840 , n9372 , n277839 );
nand ( n277841 , n277828 , n277831 , n277834 , n277840 );
buf ( n277842 , n277841 );
buf ( n277843 , n277842 );
not ( n277844 , n277843 );
not ( n277845 , n277844 );
or ( n277846 , n277824 , n277845 );
buf ( n277847 , RI21070ac0_557);
buf ( n277848 , n277847 );
not ( n277849 , n277848 );
not ( n277850 , n9251 );
or ( n277851 , n277849 , n277850 );
buf ( n277852 , RI2106d0a0_581);
not ( n277853 , n277852 );
not ( n277854 , n277853 );
not ( n277855 , n277854 );
or ( n277856 , n9392 , n277855 );
not ( n277857 , n9249 );
not ( n277858 , n277857 );
buf ( n277859 , RI21074a08_532);
buf ( n277860 , n277859 );
nand ( n277861 , n277858 , n277860 );
nand ( n277862 , n277856 , n277861 );
buf ( n277863 , n9379 );
and ( n277864 , n277862 , n277863 );
not ( n277865 , n9336 );
not ( n277866 , n277838 );
or ( n277867 , n277865 , n277866 );
nand ( n277868 , n277867 , n277768 );
and ( n277869 , n9372 , n277868 );
nor ( n277870 , n277864 , n277869 );
nand ( n277871 , n277851 , n277870 );
buf ( n277872 , n277871 );
buf ( n277873 , n277872 );
not ( n277874 , n277873 );
nand ( n277875 , n9673 , n277287 );
not ( n277876 , n277875 );
and ( n277877 , n9736 , n9681 );
not ( n277878 , n277877 );
not ( n277879 , n9664 );
or ( n277880 , n277878 , n277879 );
and ( n277881 , n277278 , n9681 );
nor ( n277882 , n277881 , n277282 );
nand ( n277883 , n277880 , n277882 );
not ( n277884 , n277883 );
or ( n277885 , n277876 , n277884 );
or ( n277886 , n277883 , n277875 );
nand ( n277887 , n277885 , n277886 );
buf ( n277888 , n277887 );
not ( n277889 , n277888 );
or ( n277890 , n277889 , n277603 );
buf ( n277891 , RI21a18ec8_13);
nand ( n277892 , n9432 , n277891 );
nand ( n277893 , n277890 , n277892 );
not ( n277894 , n277893 );
not ( n277895 , n9410 );
nor ( n277896 , n277894 , n277895 );
buf ( n277897 , n277896 );
nand ( n277898 , n277874 , n277897 );
nand ( n277899 , n277846 , n277898 );
nor ( n277900 , n277801 , n277899 );
not ( n277901 , n277900 );
not ( n277902 , n276110 );
not ( n277903 , n9056 );
or ( n277904 , n277902 , n277903 );
nand ( n277905 , n276115 , n276445 );
nand ( n277906 , n277904 , n277905 );
not ( n277907 , n277906 );
not ( n277908 , n277895 );
or ( n277909 , n277907 , n277908 );
not ( n277910 , n277603 );
not ( n277911 , n277910 );
not ( n277912 , n9716 );
or ( n277913 , n9807 , n277912 );
not ( n277914 , n277913 );
not ( n277915 , n9664 );
or ( n277916 , n277915 , n9735 );
not ( n277917 , n9802 );
nand ( n277918 , n277916 , n277917 );
not ( n277919 , n277918 );
or ( n277920 , n277914 , n277919 );
or ( n277921 , n277918 , n277913 );
nand ( n277922 , n277920 , n277921 );
buf ( n277923 , n277922 );
not ( n277924 , n277923 );
or ( n277925 , n277911 , n277924 );
buf ( n277926 , RI21a186d0_16);
nand ( n277927 , n277603 , n277926 );
nand ( n277928 , n277925 , n277927 );
nand ( n277929 , n9410 , n277928 );
nand ( n277930 , n277909 , n277929 );
buf ( n277931 , n277930 );
not ( n277932 , n277931 );
buf ( n277933 , RI2106b1b0_621);
buf ( n277934 , n277933 );
and ( n277935 , n9394 , n277934 );
not ( n277936 , n9327 );
not ( n277937 , n9325 );
not ( n277938 , n277937 );
or ( n277939 , n277936 , n277938 );
or ( n277940 , n277937 , n9327 );
nand ( n277941 , n277939 , n277940 );
and ( n277942 , n9372 , n277941 );
nor ( n277943 , n277935 , n277942 );
buf ( n277944 , RI21075638_528);
buf ( n277945 , n277944 );
nand ( n277946 , n9258 , n277945 );
buf ( n277947 , RI2106b570_613);
buf ( n277948 , n277947 );
nand ( n277949 , n9251 , n277948 );
nand ( n277950 , n277943 , n277946 , n277949 );
buf ( n277951 , n277950 );
buf ( n277952 , n277951 );
not ( n277953 , n277952 );
not ( n277954 , n277953 );
or ( n277955 , n277932 , n277954 );
buf ( n277956 , RI2106b4f8_614);
buf ( n277957 , n277956 );
not ( n277958 , n277957 );
not ( n277959 , n9251 );
or ( n277960 , n277958 , n277959 );
buf ( n277961 , RI2106b138_622);
buf ( n277962 , n277961 );
nand ( n277963 , n277365 , n277962 );
nand ( n277964 , n277960 , n277963 );
buf ( n277965 , RI210755c0_529);
buf ( n277966 , n277965 );
not ( n277967 , n277966 );
not ( n277968 , n9258 );
or ( n277969 , n277967 , n277968 );
not ( n277970 , n9329 );
not ( n277971 , n277940 );
or ( n277972 , n277970 , n277971 );
nand ( n277973 , n277972 , n9331 );
nand ( n277974 , n9372 , n277973 );
nand ( n277975 , n277969 , n277974 );
nor ( n277976 , n277964 , n277975 );
not ( n277977 , n277976 );
buf ( n277978 , n277977 );
not ( n277979 , n277978 );
not ( n277980 , n9137 );
not ( n277981 , n277895 );
or ( n277982 , n277980 , n277981 );
not ( n277983 , n277603 );
not ( n277984 , n277983 );
nand ( n277985 , n9708 , n277275 );
not ( n277986 , n277985 );
or ( n277987 , n9735 , n277912 );
or ( n277988 , n277915 , n277987 );
not ( n277989 , n277917 );
not ( n277990 , n277912 );
and ( n277991 , n277989 , n277990 );
nor ( n277992 , n277991 , n9807 );
nand ( n277993 , n277988 , n277992 );
not ( n277994 , n277993 );
or ( n277995 , n277986 , n277994 );
or ( n277996 , n277993 , n277985 );
nand ( n277997 , n277995 , n277996 );
buf ( n277998 , n277997 );
not ( n277999 , n277998 );
or ( n278000 , n277984 , n277999 );
buf ( n278001 , RI21a18748_15);
nand ( n278002 , n277603 , n278001 );
nand ( n278003 , n278000 , n278002 );
nand ( n278004 , n277389 , n278003 );
nand ( n278005 , n277982 , n278004 );
buf ( n278006 , n278005 );
nand ( n278007 , n277979 , n278006 );
nand ( n278008 , n277955 , n278007 );
buf ( n278009 , RI2106bc00_612);
buf ( n278010 , n278009 );
nand ( n278011 , n9251 , n278010 );
buf ( n278012 , RI210756b0_527);
buf ( n278013 , n278012 );
nand ( n278014 , n9258 , n278013 );
buf ( n278015 , RI2106b228_620);
buf ( n278016 , n278015 );
nand ( n278017 , n277365 , n278016 );
not ( n278018 , n9323 );
not ( n278019 , n9321 );
not ( n278020 , n278019 );
or ( n278021 , n278018 , n278020 );
nand ( n278022 , n278021 , n277937 );
nand ( n278023 , n9372 , n278022 );
nand ( n278024 , n278011 , n278014 , n278017 , n278023 );
buf ( n278025 , n278024 );
buf ( n278026 , n278025 );
not ( n278027 , n278026 );
not ( n278028 , n9241 );
not ( n278029 , n276102 );
or ( n278030 , n278028 , n278029 );
nand ( n278031 , n9039 , n276092 );
nand ( n278032 , n278030 , n278031 );
not ( n278033 , n278032 );
or ( n278034 , n277389 , n278033 );
not ( n278035 , n277910 );
nand ( n278036 , n9726 , n9801 );
not ( n278037 , n278036 );
not ( n278038 , n9734 );
or ( n278039 , n277915 , n278038 );
not ( n278040 , n9797 );
nand ( n278041 , n278039 , n278040 );
not ( n278042 , n278041 );
or ( n278043 , n278037 , n278042 );
or ( n278044 , n278041 , n278036 );
nand ( n278045 , n278043 , n278044 );
buf ( n278046 , n278045 );
not ( n278047 , n278046 );
or ( n278048 , n278035 , n278047 );
buf ( n278049 , RI21a18658_17);
nand ( n278050 , n277603 , n278049 );
nand ( n278051 , n278048 , n278050 );
nand ( n278052 , n9410 , n278051 );
nand ( n278053 , n278034 , n278052 );
buf ( n278054 , n278053 );
buf ( n278055 , n278054 );
nand ( n278056 , n278027 , n278055 );
buf ( n278057 , RI2106d190_579);
not ( n278058 , n278057 );
not ( n278059 , n278058 );
nand ( n278060 , n277365 , n278059 );
buf ( n278061 , RI21075728_526);
not ( n278062 , n278061 );
not ( n278063 , n278062 );
nand ( n278064 , n9258 , n278063 );
buf ( n278065 , RI21071600_555);
buf ( n278066 , n278065 );
nand ( n278067 , n9251 , n278066 );
not ( n278068 , n9312 );
not ( n278069 , n9300 );
not ( n278070 , n9317 );
not ( n278071 , n9315 );
not ( n278072 , n9306 );
not ( n278073 , n9293 );
nand ( n278074 , n278072 , n278073 );
nor ( n278075 , n278074 , n9295 );
nand ( n10613 , n278071 , n278075 );
buf ( n10614 , n9310 );
nor ( n10615 , n10613 , n10614 );
not ( n10616 , n10615 );
nor ( n10617 , n10616 , n9298 );
nand ( n10618 , n278070 , n10617 );
buf ( n10619 , n9303 );
nor ( n10620 , n10618 , n10619 );
nand ( n10621 , n278069 , n10620 );
not ( n10622 , n10621 );
or ( n10623 , n278068 , n10622 );
nand ( n10624 , n10623 , n278019 );
nand ( n10625 , n9372 , n10624 );
nand ( n10626 , n278060 , n278064 , n278067 , n10625 );
buf ( n10627 , n10626 );
buf ( n10628 , n10627 );
not ( n10629 , n10628 );
buf ( n10630 , n276031 );
or ( n10631 , n277389 , n10630 );
not ( n10632 , n277910 );
nor ( n10633 , n278038 , n9797 );
not ( n10634 , n10633 );
not ( n10635 , n277915 );
or ( n10636 , n10634 , n10635 );
or ( n10637 , n9665 , n10633 );
nand ( n10638 , n10636 , n10637 );
buf ( n10639 , n10638 );
not ( n10640 , n10639 );
or ( n10641 , n10632 , n10640 );
buf ( n10642 , RI21a185e0_18);
nand ( n10643 , n277352 , n10642 );
nand ( n10644 , n10641 , n10643 );
nand ( n10645 , n9410 , n10644 );
nand ( n10646 , n10631 , n10645 );
buf ( n10647 , n10646 );
buf ( n10648 , n10647 );
nor ( n10649 , n10629 , n10648 );
and ( n10650 , n278056 , n10649 );
nor ( n10651 , n278027 , n278055 );
nor ( n10652 , n10650 , n10651 );
or ( n10653 , n278008 , n10652 );
nor ( n10654 , n277953 , n277931 );
and ( n10655 , n278007 , n10654 );
not ( n10656 , n277978 );
nor ( n10657 , n10656 , n278006 );
nor ( n10658 , n10655 , n10657 );
nand ( n10659 , n10653 , n10658 );
not ( n10660 , n10659 );
or ( n10661 , n277901 , n10660 );
not ( n10662 , n277801 );
nor ( n10663 , n277844 , n277823 );
not ( n10664 , n10663 );
not ( n10665 , n277898 );
or ( n10666 , n10664 , n10665 );
not ( n10667 , n277897 );
nand ( n10668 , n10667 , n277873 );
nand ( n10669 , n10666 , n10668 );
and ( n10670 , n10662 , n10669 );
nor ( n10671 , n277777 , n277799 );
not ( n10672 , n10671 );
not ( n10673 , n277751 );
or ( n10674 , n10672 , n10673 );
not ( n10675 , n277750 );
nand ( n10676 , n10675 , n277720 );
nand ( n10677 , n10674 , n10676 );
nor ( n10678 , n10670 , n10677 );
nand ( n10679 , n10661 , n10678 );
and ( n10680 , n277701 , n10679 );
nor ( n10681 , n277678 , n277697 );
and ( n10682 , n277651 , n10681 );
nor ( n10683 , n277630 , n277650 );
nor ( n10684 , n10682 , n10683 );
or ( n10685 , n277612 , n10684 );
not ( n10686 , n277534 );
and ( n10687 , n277611 , n277555 , n10686 );
nor ( n10688 , n277577 , n277610 );
nor ( n10689 , n10687 , n10688 );
nand ( n10690 , n10685 , n10689 );
not ( n10691 , n10690 );
not ( n10692 , n277505 );
or ( n10693 , n10691 , n10692 );
not ( n10694 , n277359 );
nor ( n10695 , n277388 , n277412 );
not ( n10696 , n10695 );
not ( n10697 , n277455 );
or ( n10698 , n10696 , n10697 );
or ( n10699 , n277428 , n277454 );
nand ( n10700 , n10698 , n10699 );
and ( n10701 , n10694 , n10700 , n277503 );
not ( n10702 , n277499 );
not ( n10703 , n277502 );
not ( n10704 , n10703 );
or ( n10705 , n10702 , n10704 );
nand ( n10706 , n277503 , n9403 , n277358 );
nand ( n10707 , n10705 , n10706 );
nor ( n10708 , n10701 , n10707 );
nand ( n10709 , n10693 , n10708 );
nor ( n10710 , n10680 , n10709 );
not ( n10711 , n9022 );
nand ( n10712 , n10711 , n9165 );
not ( n10713 , n10712 );
not ( n10714 , n9042 );
or ( n10715 , n10713 , n10714 );
nand ( n10716 , n10715 , n9408 );
buf ( n10717 , n10716 );
not ( n10718 , n276375 );
not ( n10719 , n10718 );
or ( n10720 , n10717 , n10719 );
not ( n10721 , n9602 );
nand ( n10722 , n9589 , n10721 );
not ( n10723 , n10722 );
not ( n10724 , n9503 );
not ( n10725 , n9486 );
or ( n10726 , n10724 , n10725 );
nand ( n10727 , n10726 , n9619 );
not ( n10728 , n10727 );
or ( n10729 , n10723 , n10728 );
or ( n10730 , n10727 , n10722 );
nand ( n10731 , n10729 , n10730 );
buf ( n10732 , n10731 );
not ( n10733 , n10732 );
or ( n10734 , n10733 , n277603 );
buf ( n10735 , RI21a17410_28);
nand ( n10736 , n9432 , n10735 );
nand ( n10737 , n10734 , n10736 );
nand ( n10738 , n10717 , n10737 );
nand ( n10739 , n10720 , n10738 );
buf ( n10740 , n10739 );
buf ( n10741 , n10740 );
not ( n10742 , n10741 );
buf ( n10743 , n9383 );
not ( n10744 , n10743 );
buf ( n10745 , RI21072e60_547);
buf ( n10746 , n10745 );
not ( n10747 , n10746 );
not ( n10748 , n9264 );
not ( n10749 , n10748 );
or ( n10750 , n10747 , n10749 );
not ( n10751 , n277857 );
buf ( n10752 , RI2106af58_626);
buf ( n10753 , n10752 );
not ( n10754 , n10753 );
or ( n10755 , n10751 , n10754 );
nand ( n10756 , n10750 , n10755 );
not ( n10757 , n10756 );
or ( n10758 , n10744 , n10757 );
not ( n10759 , n10748 );
and ( n10760 , n9289 , n9291 );
nor ( n10761 , n10760 , n9292 );
and ( n10762 , n10759 , n10761 );
not ( n10763 , n10759 );
buf ( n10764 , RI2106dcd0_568);
buf ( n10765 , n10764 );
not ( n10766 , n10765 );
and ( n10767 , n10763 , n10766 );
nor ( n10768 , n10762 , n10767 );
buf ( n10769 , n9231 );
buf ( n10770 , n10769 );
nand ( n10771 , n10768 , n10770 );
nand ( n10772 , n10758 , n10771 );
buf ( n10773 , n10772 );
buf ( n10774 , n10773 );
not ( n10775 , n10774 );
not ( n10776 , n10775 );
or ( n10777 , n10742 , n10776 );
not ( n10778 , n10770 );
buf ( n10779 , RI2106dc58_569);
buf ( n10780 , n10779 );
not ( n10781 , n10780 );
not ( n10782 , n10748 );
or ( n10783 , n10781 , n10782 );
not ( n10784 , n9265 );
not ( n10785 , n10784 );
not ( n10786 , n9292 );
and ( n10787 , n10786 , n9277 );
nor ( n10788 , n10787 , n278073 );
or ( n10789 , n10785 , n10788 );
nand ( n10790 , n10783 , n10789 );
not ( n10791 , n10790 );
or ( n10792 , n10778 , n10791 );
buf ( n10793 , RI21072398_548);
not ( n10794 , n10793 );
not ( n10795 , n10794 );
not ( n10796 , n10795 );
not ( n10797 , n10748 );
or ( n10798 , n10796 , n10797 );
buf ( n10799 , RI2106aee0_627);
buf ( n10800 , n10799 );
nand ( n10801 , n10759 , n10800 );
nand ( n10802 , n10798 , n10801 );
not ( n10803 , n10770 );
nand ( n10804 , n10802 , n10803 );
nand ( n10805 , n10792 , n10804 );
buf ( n10806 , n10805 );
buf ( n10807 , n10806 );
not ( n10808 , n10807 );
buf ( n10809 , n276250 );
or ( n10810 , n10717 , n10809 );
not ( n10811 , n277983 );
nand ( n10812 , n9554 , n9606 );
not ( n10813 , n10812 );
not ( n10814 , n9589 );
not ( n10815 , n9503 );
nor ( n10816 , n10814 , n10815 );
not ( n10817 , n10816 );
not ( n10818 , n9486 );
or ( n10819 , n10817 , n10818 );
nand ( n10820 , n9618 , n9589 );
and ( n10821 , n10820 , n10721 );
nand ( n10822 , n10819 , n10821 );
not ( n10823 , n10822 );
or ( n10824 , n10813 , n10823 );
or ( n10825 , n10822 , n10812 );
nand ( n10826 , n10824 , n10825 );
buf ( n10827 , n10826 );
not ( n10828 , n10827 );
or ( n10829 , n10811 , n10828 );
buf ( n10830 , RI21a17488_27);
nand ( n10831 , n277350 , n10830 );
nand ( n10832 , n10829 , n10831 );
nand ( n10833 , n10717 , n10832 );
nand ( n10834 , n10810 , n10833 );
not ( n10835 , n10834 );
not ( n10836 , n10835 );
buf ( n10837 , n10836 );
nand ( n10838 , n10808 , n10837 );
nand ( n10839 , n10777 , n10838 );
buf ( n10840 , n276275 );
not ( n10841 , n10840 );
not ( n10842 , n10841 );
not ( n10843 , n9410 );
not ( n10844 , n10843 );
or ( n10845 , n10842 , n10844 );
buf ( n10846 , RI21a17320_30);
and ( n10847 , n9430 , n10846 );
not ( n10848 , n9430 );
not ( n10849 , n9613 );
nand ( n10850 , n9494 , n10849 );
not ( n10851 , n10850 );
not ( n10852 , n9486 );
or ( n10853 , n10851 , n10852 );
or ( n10854 , n9486 , n10850 );
nand ( n10855 , n10853 , n10854 );
buf ( n10856 , n10855 );
and ( n10857 , n10848 , n10856 );
or ( n10858 , n10847 , n10857 );
nand ( n10859 , n9410 , n10858 );
nand ( n10860 , n10845 , n10859 );
not ( n10861 , n10860 );
not ( n10862 , n10861 );
buf ( n10863 , n10862 );
not ( n10864 , n10863 );
not ( n10865 , n10769 );
buf ( n10866 , RI21072f50_545);
not ( n10867 , n10866 );
not ( n10868 , n10867 );
not ( n10869 , n10868 );
not ( n10870 , n277364 );
not ( n10871 , n10870 );
or ( n10872 , n10869 , n10871 );
buf ( n10873 , RI2106afd0_625);
buf ( n10874 , n10873 );
not ( n10875 , n10874 );
or ( n10876 , n10785 , n10875 );
nand ( n10877 , n10872 , n10876 );
and ( n10878 , n10865 , n10877 );
not ( n10879 , n10865 );
buf ( n10880 , RI2106b318_618);
buf ( n10881 , n10880 );
not ( n10882 , n10881 );
not ( n10883 , n10870 );
or ( n10884 , n10882 , n10883 );
buf ( n10885 , n9287 );
and ( n10886 , n9285 , n10885 );
buf ( n10887 , n9288 );
nor ( n10888 , n10886 , n10887 );
or ( n10889 , n10870 , n10888 );
nand ( n10890 , n10884 , n10889 );
and ( n10891 , n10879 , n10890 );
nor ( n10892 , n10878 , n10891 );
not ( n10893 , n10892 );
buf ( n10894 , n10893 );
not ( n10895 , n10894 );
not ( n10896 , n10895 );
or ( n10897 , n10864 , n10896 );
not ( n10898 , n10784 );
not ( n10899 , n10898 );
not ( n10900 , n10769 );
buf ( n10901 , RI2106cb00_593);
buf ( n10902 , n10901 );
nand ( n10903 , n10899 , n10900 , n10902 );
not ( n10904 , n9249 );
not ( n10905 , n10904 );
buf ( n10906 , RI2106b2a0_619);
buf ( n10907 , n10906 );
nand ( n10908 , n10905 , n9380 , n10907 );
buf ( n10909 , RI21072ed8_546);
not ( n10910 , n10909 );
not ( n10911 , n10910 );
nand ( n10912 , n10898 , n9383 , n10911 );
not ( n10913 , n9281 );
not ( n10914 , n10887 );
not ( n10915 , n10914 );
or ( n10916 , n10913 , n10915 );
nand ( n10917 , n10916 , n9289 );
and ( n10918 , n9369 , n10917 );
nand ( n10919 , n9384 , n10918 );
nand ( n10920 , n10903 , n10908 , n10912 , n10919 );
buf ( n10921 , n10920 );
buf ( n10922 , n10921 );
not ( n10923 , n10922 );
buf ( n10924 , n276263 );
or ( n10925 , n9410 , n10924 );
nand ( n10926 , n9502 , n9617 );
not ( n10927 , n10926 );
nand ( n10928 , n9494 , n9472 );
not ( n10929 , n10928 );
not ( n10930 , n9438 );
nand ( n10931 , n9464 , n9451 , n10930 );
not ( n10932 , n10931 );
and ( n10933 , n10929 , n10932 );
not ( n10934 , n9494 );
or ( n10935 , n10934 , n9483 );
nand ( n10936 , n10935 , n10849 );
nor ( n10937 , n10933 , n10936 );
not ( n10938 , n9464 );
nor ( n10939 , n10934 , n10938 );
not ( n10940 , n9472 );
nor ( n10941 , n10940 , n9454 );
nand ( n10942 , n10939 , n10941 );
not ( n10943 , n10928 );
not ( n10944 , n9441 );
and ( n10945 , n9464 , n9451 , n10944 );
nand ( n10946 , n10943 , n10945 );
nand ( n10947 , n10939 , n9477 );
nand ( n10948 , n10937 , n10942 , n10946 , n10947 );
not ( n10949 , n10948 );
or ( n10950 , n10927 , n10949 );
or ( n10951 , n10948 , n10926 );
nand ( n10952 , n10950 , n10951 );
buf ( n10953 , n10952 );
not ( n10954 , n10953 );
or ( n10955 , n10954 , n277603 );
buf ( n10956 , RI21a17398_29);
nand ( n10957 , n9432 , n10956 );
nand ( n10958 , n10955 , n10957 );
nand ( n10959 , n10717 , n10958 );
nand ( n10960 , n10925 , n10959 );
buf ( n10961 , n10960 );
buf ( n10962 , n10961 );
nand ( n10963 , n10923 , n10962 );
nand ( n10964 , n10897 , n10963 );
nor ( n10965 , n10839 , n10964 );
buf ( n10966 , n276306 );
not ( n10967 , n10966 );
not ( n10968 , n10717 );
not ( n10969 , n10968 );
or ( n10970 , n10967 , n10969 );
buf ( n10971 , RI21a16b28_33);
and ( n10972 , n277350 , n10971 );
not ( n10973 , n277350 );
not ( n10974 , n9442 );
nand ( n10975 , n9451 , n9454 );
not ( n10976 , n10975 );
or ( n10977 , n10974 , n10976 );
or ( n10978 , n10975 , n9442 );
nand ( n10979 , n10977 , n10978 );
buf ( n10980 , n10979 );
and ( n10981 , n10973 , n10980 );
or ( n10982 , n10972 , n10981 );
nand ( n10983 , n10717 , n10982 );
nand ( n10984 , n10970 , n10983 );
not ( n10985 , n10984 );
not ( n10986 , n10985 );
buf ( n10987 , n10986 );
not ( n10988 , n10987 );
not ( n10989 , n9231 );
buf ( n10990 , RI2106b0c0_623);
buf ( n10991 , n10990 );
nand ( n10992 , n10989 , n10991 );
nor ( n10993 , n10748 , n10992 );
not ( n10994 , n10993 );
buf ( n10995 , RI2106b480_615);
buf ( n10996 , n10995 );
not ( n10997 , n10996 );
nor ( n10998 , n9379 , n10997 );
nand ( n10999 , n10998 , n10870 );
not ( n11000 , n9231 );
buf ( n11001 , RI21074af8_530);
not ( n11002 , n11001 );
not ( n11003 , n11002 );
nand ( n11004 , n10748 , n11000 , n11003 );
buf ( n11005 , RI2106a418_637);
buf ( n11006 , n11005 );
and ( n11007 , n9369 , n11006 );
nand ( n11008 , n9380 , n11007 );
nand ( n11009 , n10994 , n10999 , n11004 , n11008 );
buf ( n11010 , n11009 );
buf ( n11011 , n11010 );
not ( n11012 , n11011 );
not ( n11013 , n11012 );
or ( n11014 , n10988 , n11013 );
not ( n11015 , n9392 );
buf ( n11016 , RI21072230_551);
not ( n11017 , n11016 );
not ( n11018 , n11017 );
not ( n11019 , n11018 );
not ( n11020 , n9231 );
or ( n11021 , n11019 , n11020 );
buf ( n11022 , RI210764c0_519);
not ( n11023 , n11022 );
not ( n11024 , n11023 );
not ( n11025 , n11024 );
or ( n11026 , n9231 , n11025 );
nand ( n11027 , n11021 , n11026 );
not ( n11028 , n11027 );
or ( n11029 , n11015 , n11028 );
buf ( n11030 , n9265 );
not ( n11031 , n11030 );
buf ( n11032 , RI2106c380_596);
not ( n11033 , n11032 );
not ( n11034 , n11033 );
not ( n11035 , n11034 );
not ( n11036 , n9231 );
or ( n11037 , n11035 , n11036 );
buf ( n11038 , RI2106daf0_572);
not ( n11039 , n11038 );
not ( n11040 , n11039 );
not ( n11041 , n11040 );
or ( n11042 , n9231 , n11041 );
nand ( n11043 , n11037 , n11042 );
nand ( n11044 , n11031 , n11043 );
nand ( n11045 , n11029 , n11044 );
buf ( n11046 , n11045 );
buf ( n11047 , n11046 );
not ( n11048 , n11047 );
or ( n11049 , n10717 , n9194 );
buf ( n11050 , RI21a16ab0_34);
not ( n11051 , n11050 );
not ( n11052 , n9430 );
or ( n11053 , n11051 , n11052 );
not ( n11054 , n10930 );
not ( n11055 , n10944 );
or ( n11056 , n11054 , n11055 );
nand ( n11057 , n11056 , n9442 );
buf ( n11058 , n11057 );
nand ( n11059 , n9431 , n11058 );
nand ( n11060 , n11053 , n11059 );
nand ( n11061 , n10717 , n11060 );
nand ( n11062 , n11049 , n11061 );
buf ( n11063 , n11062 );
buf ( n11064 , n11063 );
nand ( n11065 , n11048 , n11064 );
nand ( n11066 , n11014 , n11065 );
not ( n11067 , n10987 );
nand ( n11068 , n11067 , n11011 );
nand ( n11069 , n11066 , n11068 );
not ( n11070 , n9231 );
buf ( n11071 , RI2106cb78_592);
not ( n11072 , n11071 );
not ( n11073 , n11072 );
not ( n11074 , n11073 );
not ( n11075 , n277857 );
or ( n11076 , n11074 , n11075 );
not ( n11077 , n9249 );
buf ( n11078 , RI21072fc8_544);
not ( n11079 , n11078 );
not ( n11080 , n11079 );
not ( n11081 , n11080 );
or ( n11082 , n11077 , n11081 );
nand ( n11083 , n11076 , n11082 );
and ( n11084 , n11070 , n11083 );
not ( n11085 , n11070 );
not ( n11086 , n10784 );
or ( n11087 , n11086 , n10885 );
not ( n11088 , n10904 );
buf ( n11089 , RI2106b390_617);
buf ( n11090 , n11089 );
not ( n11091 , n11090 );
not ( n11092 , n11091 );
nand ( n11093 , n11088 , n11092 );
nand ( n11094 , n11087 , n11093 );
and ( n11095 , n11085 , n11094 );
or ( n11096 , n11084 , n11095 );
buf ( n11097 , n11096 );
buf ( n11098 , n11097 );
not ( n11099 , n11098 );
not ( n11100 , n276323 );
not ( n11101 , n10968 );
or ( n11102 , n11100 , n11101 );
buf ( n11103 , RI21a172a8_31);
and ( n11104 , n277817 , n11103 );
not ( n11105 , n277817 );
not ( n11106 , n10938 );
nand ( n11107 , n11106 , n9483 );
not ( n11108 , n11107 );
not ( n11109 , n9472 );
not ( n11110 , n9455 );
or ( n11111 , n11109 , n11110 );
not ( n11112 , n9477 );
nand ( n11113 , n11111 , n11112 );
not ( n11114 , n11113 );
or ( n11115 , n11108 , n11114 );
or ( n11116 , n11113 , n11107 );
nand ( n11117 , n11115 , n11116 );
buf ( n11118 , n11117 );
and ( n11119 , n11105 , n11118 );
or ( n11120 , n11104 , n11119 );
nand ( n11121 , n10717 , n11120 );
nand ( n11122 , n11102 , n11121 );
buf ( n11123 , n11122 );
nand ( n11124 , n11099 , n11123 );
not ( n11125 , n10748 );
buf ( n11126 , RI2106b048_624);
buf ( n11127 , n11126 );
nand ( n11128 , n11125 , n11070 , n11127 );
buf ( n11129 , RI2106b408_616);
buf ( n11130 , n11129 );
nand ( n11131 , n10905 , n10769 , n11130 );
buf ( n11132 , RI21073b80_541);
not ( n11133 , n11132 );
not ( n11134 , n11133 );
nand ( n11135 , n11030 , n9383 , n11134 );
buf ( n11136 , RI2106a1c0_642);
buf ( n11137 , n11136 );
and ( n11138 , n9369 , n11137 );
nand ( n11139 , n10769 , n11138 );
nand ( n11140 , n11128 , n11131 , n11135 , n11139 );
buf ( n11141 , n11140 );
buf ( n11142 , n11141 );
not ( n11143 , n11142 );
buf ( n11144 , n276292 );
not ( n11145 , n11144 );
or ( n11146 , n10717 , n11145 );
buf ( n11147 , RI21a17230_32);
not ( n11148 , n11147 );
not ( n11149 , n277350 );
or ( n11150 , n11148 , n11149 );
nand ( n11151 , n9472 , n11112 );
not ( n11152 , n11151 );
not ( n11153 , n9455 );
or ( n11154 , n11152 , n11153 );
or ( n11155 , n9455 , n11151 );
nand ( n11156 , n11154 , n11155 );
buf ( n11157 , n11156 );
nand ( n11158 , n11157 , n9431 );
nand ( n11159 , n11150 , n11158 );
nand ( n11160 , n10717 , n11159 );
nand ( n11161 , n11146 , n11160 );
buf ( n11162 , n11161 );
nand ( n11163 , n11143 , n11162 );
nand ( n11164 , n11069 , n11124 , n11163 );
not ( n11165 , n11123 );
nand ( n11166 , n11165 , n11098 );
not ( n11167 , n11166 );
not ( n11168 , n11162 );
nand ( n11169 , n11168 , n11142 );
not ( n11170 , n11169 );
or ( n11171 , n11167 , n11170 );
nand ( n11172 , n11171 , n11124 );
nand ( n11173 , n11164 , n11172 );
nand ( n11174 , n10965 , n11173 );
not ( n11175 , n11174 );
not ( n11176 , n10839 );
nor ( n11177 , n10895 , n10863 );
not ( n11178 , n11177 );
not ( n11179 , n10963 );
or ( n11180 , n11178 , n11179 );
not ( n11181 , n10962 );
nand ( n11182 , n11181 , n10922 );
nand ( n11183 , n11180 , n11182 );
and ( n11184 , n11176 , n11183 );
nor ( n11185 , n10775 , n10741 );
not ( n11186 , n11185 );
not ( n11187 , n10838 );
or ( n11188 , n11186 , n11187 );
not ( n11189 , n10837 );
nand ( n11190 , n11189 , n10807 );
nand ( n11191 , n11188 , n11190 );
nor ( n11192 , n11184 , n11191 );
not ( n11193 , n11192 );
or ( n11194 , n11175 , n11193 );
not ( n11195 , n276445 );
buf ( n11196 , n276009 );
and ( n11197 , n11195 , n11196 );
not ( n11198 , n11195 );
buf ( n11199 , n276068 );
and ( n11200 , n11198 , n11199 );
nor ( n11201 , n11197 , n11200 );
not ( n11202 , n11201 );
not ( n11203 , n11202 );
not ( n11204 , n277895 );
or ( n11205 , n11203 , n11204 );
not ( n11206 , n9433 );
not ( n11207 , n9656 );
nand ( n11208 , n9564 , n11207 );
not ( n11209 , n11208 );
and ( n11210 , n9595 , n9520 );
and ( n11211 , n11210 , n9597 );
not ( n11212 , n11211 );
nor ( n11213 , n10815 , n9609 );
not ( n11214 , n11213 );
not ( n11215 , n9486 );
or ( n11216 , n11214 , n11215 );
not ( n11217 , n9609 );
not ( n11218 , n11217 );
not ( n11219 , n9618 );
or ( n11220 , n11218 , n11219 );
nand ( n11221 , n11220 , n9608 );
not ( n11222 , n11221 );
nand ( n11223 , n11216 , n11222 );
not ( n11224 , n11223 );
or ( n11225 , n11212 , n11224 );
and ( n11226 , n9639 , n9597 );
nor ( n11227 , n11226 , n9652 );
nand ( n11228 , n11225 , n11227 );
not ( n11229 , n11228 );
or ( n11230 , n11209 , n11229 );
or ( n11231 , n11228 , n11208 );
nand ( n11232 , n11230 , n11231 );
buf ( n11233 , n11232 );
not ( n11234 , n11233 );
or ( n11235 , n11206 , n11234 );
buf ( n11236 , RI21a184f0_20);
nand ( n11237 , n277527 , n11236 );
nand ( n11238 , n11235 , n11237 );
nand ( n11239 , n9410 , n11238 );
nand ( n11240 , n11205 , n11239 );
buf ( n11241 , n11240 );
buf ( n11242 , n11241 );
not ( n11243 , n11242 );
not ( n11244 , n10620 );
nand ( n11245 , n10618 , n10619 );
nand ( n11246 , n11244 , n11245 );
nand ( n11247 , n11246 , n9369 );
nor ( n11248 , n9379 , n11247 );
not ( n11249 , n11248 );
buf ( n11250 , RI2106d898_577);
not ( n11251 , n11250 );
not ( n11252 , n11251 );
nand ( n11253 , n11031 , n9383 , n11252 );
not ( n11254 , n11077 );
buf ( n11255 , RI2106bc78_611);
buf ( n11256 , n11255 );
nand ( n11257 , n11254 , n10769 , n11256 );
buf ( n11258 , RI21075818_524);
not ( n11259 , n11258 );
not ( n11260 , n11259 );
nand ( n11261 , n11030 , n9383 , n11260 );
nand ( n11262 , n11249 , n11253 , n11257 , n11261 );
buf ( n11263 , n11262 );
not ( n11264 , n11263 );
not ( n11265 , n11264 );
or ( n11266 , n11243 , n11265 );
buf ( n11267 , RI210757a0_525);
not ( n11268 , n11267 );
not ( n11269 , n11268 );
not ( n11270 , n11269 );
not ( n11271 , n10748 );
or ( n11272 , n11270 , n11271 );
buf ( n11273 , RI2106d208_578);
not ( n11274 , n11273 );
not ( n11275 , n11274 );
nand ( n11276 , n11125 , n11275 );
nand ( n11277 , n11272 , n11276 );
and ( n11278 , n10743 , n11277 );
not ( n11279 , n10743 );
not ( n11280 , n9300 );
nor ( n11281 , n11280 , n10620 );
not ( n11282 , n11281 );
nand ( n11283 , n11282 , n10621 );
not ( n11284 , n11283 );
buf ( n11285 , n277364 );
not ( n11286 , n11285 );
or ( n11287 , n11284 , n11286 );
buf ( n11288 , n9249 );
buf ( n11289 , RI21071678_554);
buf ( n11290 , n11289 );
nand ( n11291 , n11288 , n11290 );
nand ( n11292 , n11287 , n11291 );
and ( n11293 , n11279 , n11292 );
nor ( n11294 , n11278 , n11293 );
not ( n11295 , n11294 );
buf ( n11296 , n11295 );
not ( n11297 , n11296 );
buf ( n11298 , n276013 );
and ( n11299 , n9053 , n11298 );
not ( n11300 , n9053 );
and ( n11301 , n11300 , n276140 );
or ( n11302 , n11299 , n11301 );
not ( n11303 , n11302 );
not ( n11304 , n10843 );
or ( n11305 , n11303 , n11304 );
not ( n11306 , n9433 );
not ( n11307 , n9659 );
nand ( n11308 , n11307 , n9529 );
not ( n11309 , n11308 );
and ( n11310 , n9597 , n9564 );
and ( n11311 , n11210 , n11310 );
not ( n11312 , n11311 );
not ( n11313 , n11223 );
or ( n11314 , n11312 , n11313 );
and ( n11315 , n9639 , n11310 );
not ( n11316 , n9564 );
not ( n11317 , n9652 );
or ( n11318 , n11316 , n11317 );
nand ( n11319 , n11318 , n11207 );
nor ( n11320 , n11315 , n11319 );
nand ( n11321 , n11314 , n11320 );
not ( n11322 , n11321 );
or ( n11323 , n11309 , n11322 );
or ( n11324 , n11321 , n11308 );
nand ( n11325 , n11323 , n11324 );
buf ( n11326 , n11325 );
not ( n11327 , n11326 );
or ( n11328 , n11306 , n11327 );
buf ( n11329 , RI21a18568_19);
nand ( n11330 , n277527 , n11329 );
nand ( n11331 , n11328 , n11330 );
nand ( n11332 , n10717 , n11331 );
nand ( n11333 , n11305 , n11332 );
buf ( n11334 , n11333 );
nand ( n11335 , n11297 , n11334 );
nand ( n11336 , n11266 , n11335 );
buf ( n11337 , n276090 );
and ( n11338 , n276445 , n11337 );
not ( n11339 , n276445 );
buf ( n11340 , n275975 );
and ( n11341 , n11339 , n11340 );
nor ( n11342 , n11338 , n11341 );
not ( n11343 , n11342 );
not ( n11344 , n11343 );
not ( n11345 , n9410 );
not ( n11346 , n11345 );
or ( n11347 , n11344 , n11346 );
not ( n11348 , n9433 );
not ( n11349 , n9647 );
nand ( n11350 , n11349 , n9581 );
not ( n11351 , n11350 );
not ( n11352 , n11210 );
not ( n11353 , n11223 );
or ( n11354 , n11352 , n11353 );
not ( n11355 , n9639 );
nand ( n11356 , n11354 , n11355 );
not ( n11357 , n11356 );
or ( n11358 , n11351 , n11357 );
or ( n11359 , n11356 , n11350 );
nand ( n11360 , n11358 , n11359 );
buf ( n11361 , n11360 );
not ( n11362 , n11361 );
or ( n11363 , n11348 , n11362 );
buf ( n11364 , RI21a17d70_22);
nand ( n11365 , n277527 , n11364 );
nand ( n11366 , n11363 , n11365 );
nand ( n11367 , n9410 , n11366 );
nand ( n11368 , n11347 , n11367 );
buf ( n11369 , n11368 );
not ( n11370 , n11369 );
buf ( n11371 , RI210716f0_553);
buf ( n11372 , n11371 );
not ( n11373 , n11372 );
not ( n11374 , n9251 );
or ( n11375 , n11373 , n11374 );
buf ( n11376 , RI2106d988_575);
not ( n11377 , n11376 );
not ( n11378 , n11377 );
not ( n11379 , n11378 );
or ( n11380 , n11086 , n11379 );
buf ( n11381 , RI21076358_522);
not ( n11382 , n11381 );
not ( n11383 , n11382 );
nand ( n11384 , n11086 , n11383 );
nand ( n11385 , n11380 , n11384 );
and ( n11386 , n11385 , n10743 );
not ( n11387 , n9298 );
not ( n11388 , n10615 );
not ( n11389 , n11388 );
or ( n11390 , n11387 , n11389 );
not ( n11391 , n10617 );
nand ( n11392 , n11390 , n11391 );
and ( n11393 , n9372 , n11392 );
nor ( n11394 , n11386 , n11393 );
nand ( n11395 , n11375 , n11394 );
buf ( n11396 , n11395 );
buf ( n11397 , n11396 );
not ( n11398 , n11397 );
not ( n11399 , n11398 );
or ( n11400 , n11370 , n11399 );
not ( n11401 , n9317 );
not ( n11402 , n11391 );
or ( n11403 , n11401 , n11402 );
nand ( n11404 , n11403 , n10618 );
nand ( n11405 , n11404 , n9369 );
nor ( n11406 , n9383 , n11405 );
not ( n11407 , n11406 );
not ( n11408 , n10905 );
buf ( n11409 , RI2106d910_576);
not ( n11410 , n11409 );
not ( n11411 , n11410 );
nand ( n11412 , n11408 , n9383 , n11411 );
not ( n11413 , n11070 );
buf ( n11414 , RI2106bcf0_610);
buf ( n11415 , n11414 );
nand ( n11416 , n11288 , n11413 , n11415 );
buf ( n11417 , RI210762e0_523);
not ( n11418 , n11417 );
not ( n11419 , n11418 );
nand ( n11420 , n11254 , n9379 , n11419 );
nand ( n11421 , n11407 , n11412 , n11416 , n11420 );
buf ( n11422 , n11421 );
buf ( n11423 , n11422 );
not ( n11424 , n11423 );
not ( n11425 , n276430 );
buf ( n11426 , n275968 );
and ( n11427 , n11425 , n11426 );
not ( n11428 , n11425 );
buf ( n11429 , n276080 );
and ( n11430 , n11428 , n11429 );
nor ( n11431 , n11427 , n11430 );
not ( n11432 , n11431 );
not ( n11433 , n11432 );
or ( n11434 , n9410 , n11433 );
not ( n11435 , n9431 );
nand ( n11436 , n9546 , n9651 );
not ( n11437 , n11436 );
and ( n11438 , n11210 , n9581 );
not ( n11439 , n11438 );
not ( n11440 , n11223 );
or ( n11441 , n11439 , n11440 );
and ( n11442 , n9639 , n9581 );
nor ( n11443 , n11442 , n9647 );
nand ( n11444 , n11441 , n11443 );
not ( n11445 , n11444 );
or ( n11446 , n11437 , n11445 );
or ( n11447 , n11444 , n11436 );
nand ( n11448 , n11446 , n11447 );
buf ( n11449 , n11448 );
not ( n11450 , n11449 );
or ( n11451 , n11435 , n11450 );
buf ( n11452 , RI21a17de8_21);
nand ( n11453 , n277352 , n11452 );
nand ( n11454 , n11451 , n11453 );
nand ( n11455 , n9410 , n11454 );
nand ( n11456 , n11434 , n11455 );
buf ( n11457 , n11456 );
buf ( n11458 , n11457 );
nand ( n11459 , n11424 , n11458 );
nand ( n11460 , n11400 , n11459 );
nor ( n11461 , n11336 , n11460 );
not ( n11462 , n11285 );
and ( n11463 , n10613 , n10614 );
nor ( n11464 , n11463 , n10615 );
or ( n11465 , n11462 , n11464 );
buf ( n11466 , RI210721b8_552);
buf ( n11467 , n11466 );
nand ( n11468 , n10748 , n11467 );
nand ( n11469 , n11465 , n11468 );
not ( n11470 , n10743 );
and ( n11471 , n11469 , n11470 );
buf ( n11472 , RI2106da00_574);
not ( n11473 , n11472 );
not ( n11474 , n11473 );
nand ( n11475 , n9391 , n11474 );
buf ( n11476 , RI210763d0_521);
not ( n11477 , n11476 );
not ( n11478 , n11477 );
nand ( n11479 , n10905 , n11478 );
and ( n11480 , n11475 , n11479 );
nor ( n11481 , n11480 , n10770 );
nor ( n11482 , n11471 , n11481 );
not ( n11483 , n11482 );
buf ( n11484 , n11483 );
not ( n11485 , n11484 );
buf ( n11486 , n276125 );
and ( n11487 , n11486 , n276445 );
and ( n11488 , n9039 , n275994 );
nor ( n11489 , n11487 , n11488 );
not ( n11490 , n11489 );
not ( n11491 , n11490 );
not ( n11492 , n11345 );
or ( n11493 , n11491 , n11492 );
not ( n11494 , n277910 );
not ( n11495 , n9637 );
nand ( n11496 , n11495 , n9537 );
not ( n11497 , n11496 );
and ( n11498 , n9520 , n9572 );
not ( n11499 , n11498 );
not ( n11500 , n11223 );
or ( n11501 , n11499 , n11500 );
and ( n11502 , n9628 , n9572 );
nor ( n11503 , n11502 , n9634 );
nand ( n11504 , n11501 , n11503 );
not ( n11505 , n11504 );
or ( n11506 , n11497 , n11505 );
or ( n11507 , n11504 , n11496 );
nand ( n11508 , n11506 , n11507 );
buf ( n11509 , n11508 );
not ( n11510 , n11509 );
or ( n11511 , n11494 , n11510 );
buf ( n11512 , RI21a17cf8_23);
nand ( n11513 , n9432 , n11512 );
nand ( n11514 , n11511 , n11513 );
nand ( n11515 , n9410 , n11514 );
nand ( n11516 , n11493 , n11515 );
buf ( n11517 , n11516 );
buf ( n11518 , n11517 );
nand ( n11519 , n11485 , n11518 );
buf ( n11520 , RI2106da78_573);
not ( n11521 , n11520 );
not ( n11522 , n11521 );
not ( n11523 , n11522 );
or ( n11524 , n11288 , n11523 );
buf ( n11525 , RI21076448_520);
not ( n11526 , n11525 );
not ( n11527 , n11526 );
nand ( n11528 , n11288 , n11527 );
nand ( n11529 , n11524 , n11528 );
and ( n11530 , n10865 , n11529 );
not ( n11531 , n10865 );
not ( n11532 , n278075 );
and ( n11533 , n11532 , n9315 );
not ( n11534 , n10613 );
nor ( n11535 , n11533 , n11534 );
or ( n11536 , n11086 , n11535 );
buf ( n11537 , RI2106bd68_609);
buf ( n11538 , n11537 );
nand ( n11539 , n10870 , n11538 );
nand ( n11540 , n11536 , n11539 );
and ( n11541 , n11531 , n11540 );
or ( n11542 , n11530 , n11541 );
buf ( n11543 , n11542 );
buf ( n11544 , n11543 );
not ( n11545 , n11544 );
buf ( n11546 , n275985 );
and ( n11547 , n11425 , n11546 );
not ( n11548 , n11425 );
and ( n11549 , n11548 , n276337 );
nor ( n11550 , n11547 , n11549 );
or ( n11551 , n9410 , n11550 );
not ( n11552 , n9433 );
not ( n11553 , n9634 );
nand ( n11554 , n11553 , n9572 );
not ( n11555 , n11554 );
not ( n11556 , n9520 );
not ( n11557 , n11223 );
or ( n11558 , n11556 , n11557 );
not ( n11559 , n9628 );
nand ( n11560 , n11558 , n11559 );
not ( n11561 , n11560 );
or ( n11562 , n11555 , n11561 );
or ( n11563 , n11560 , n11554 );
nand ( n11564 , n11562 , n11563 );
buf ( n11565 , n11564 );
not ( n11566 , n11565 );
or ( n11567 , n11552 , n11566 );
buf ( n11568 , RI21a17c80_24);
nand ( n11569 , n277527 , n11568 );
nand ( n11570 , n11567 , n11569 );
nand ( n11571 , n9410 , n11570 );
nand ( n11572 , n11551 , n11571 );
buf ( n11573 , n11572 );
buf ( n11574 , n11573 );
nand ( n11575 , n11545 , n11574 );
nand ( n11576 , n11519 , n11575 );
not ( n11577 , n276361 );
not ( n11578 , n11577 );
not ( n11579 , n10843 );
or ( n11580 , n11578 , n11579 );
not ( n11581 , n9433 );
not ( n11582 , n9624 );
nand ( n11583 , n9519 , n11582 );
not ( n11584 , n11583 );
not ( n11585 , n11223 );
or ( n11586 , n11584 , n11585 );
or ( n11587 , n11223 , n11583 );
nand ( n11588 , n11586 , n11587 );
buf ( n11589 , n11588 );
not ( n11590 , n11589 );
or ( n11591 , n11581 , n11590 );
buf ( n11592 , RI21a17b90_26);
nand ( n11593 , n277352 , n11592 );
nand ( n11594 , n11591 , n11593 );
nand ( n11595 , n9410 , n11594 );
nand ( n11596 , n11580 , n11595 );
buf ( n11597 , n11596 );
not ( n11598 , n11597 );
not ( n11599 , n11288 );
buf ( n11600 , RI2106ca88_594);
not ( n11601 , n11600 );
not ( n11602 , n11601 );
nand ( n11603 , n11599 , n11070 , n11602 );
not ( n11604 , n9306 );
not ( n11605 , n9293 );
or ( n11606 , n11604 , n11605 );
nand ( n11607 , n11606 , n278074 );
not ( n11608 , n11607 );
nor ( n11609 , n11608 , n9370 );
nand ( n11610 , n11413 , n11609 );
buf ( n11611 , RI21072320_549);
not ( n11612 , n11611 );
not ( n11613 , n11612 );
nand ( n11614 , n10905 , n11070 , n11613 );
buf ( n11615 , RI2106dbe0_570);
buf ( n11616 , n11615 );
nand ( n11617 , n11254 , n10769 , n11616 );
nand ( n11618 , n11603 , n11610 , n11614 , n11617 );
buf ( n11619 , n11618 );
buf ( n11620 , n11619 );
not ( n11621 , n11620 );
not ( n11622 , n11621 );
or ( n11623 , n11598 , n11622 );
buf ( n11624 , RI2106ca10_595);
not ( n11625 , n11624 );
not ( n11626 , n11625 );
not ( n11627 , n11626 );
not ( n11628 , n277857 );
or ( n11629 , n11627 , n11628 );
buf ( n11630 , RI210722a8_550);
not ( n11631 , n11630 );
not ( n11632 , n11631 );
not ( n11633 , n11632 );
or ( n11634 , n11077 , n11633 );
nand ( n11635 , n11629 , n11634 );
and ( n11636 , n277863 , n11635 );
not ( n11637 , n277863 );
buf ( n11638 , RI2106db68_571);
buf ( n11639 , n11638 );
not ( n11640 , n11639 );
not ( n11641 , n11030 );
or ( n11642 , n11640 , n11641 );
and ( n11643 , n278074 , n9295 );
nor ( n11644 , n11643 , n278075 );
or ( n11645 , n11088 , n11644 );
nand ( n11646 , n11642 , n11645 );
and ( n11647 , n11637 , n11646 );
or ( n11648 , n11636 , n11647 );
buf ( n11649 , n11648 );
buf ( n11650 , n11649 );
not ( n11651 , n11650 );
buf ( n11652 , n276348 );
and ( n11653 , n11652 , n276430 );
and ( n11654 , n9053 , n276004 );
nor ( n11655 , n11653 , n11654 );
buf ( n11656 , n11655 );
or ( n11657 , n9410 , n11656 );
not ( n11658 , n9431 );
nand ( n11659 , n9511 , n9627 );
not ( n11660 , n11659 );
not ( n11661 , n9519 );
not ( n11662 , n11223 );
or ( n11663 , n11661 , n11662 );
nand ( n11664 , n11663 , n11582 );
not ( n11665 , n11664 );
or ( n11666 , n11660 , n11665 );
or ( n11667 , n11664 , n11659 );
nand ( n11668 , n11666 , n11667 );
buf ( n11669 , n11668 );
not ( n11670 , n11669 );
or ( n11671 , n11658 , n11670 );
buf ( n11672 , RI21a17c08_25);
nand ( n11673 , n277352 , n11672 );
nand ( n11674 , n11671 , n11673 );
nand ( n11675 , n10717 , n11674 );
nand ( n11676 , n11657 , n11675 );
buf ( n11677 , n11676 );
buf ( n11678 , n11677 );
nand ( n11679 , n11651 , n11678 );
nand ( n11680 , n11623 , n11679 );
nor ( n11681 , n11576 , n11680 );
and ( n11682 , n11461 , n11681 );
nand ( n11683 , n11194 , n11682 );
nor ( n11684 , n11621 , n11597 );
not ( n11685 , n11684 );
not ( n11686 , n11679 );
or ( n11687 , n11685 , n11686 );
not ( n11688 , n11678 );
nand ( n11689 , n11688 , n11650 );
nand ( n11690 , n11687 , n11689 );
not ( n11691 , n11690 );
not ( n11692 , n11576 );
not ( n11693 , n11692 );
or ( n11694 , n11691 , n11693 );
not ( n11695 , n11544 );
nor ( n11696 , n11695 , n11574 );
and ( n11697 , n11519 , n11696 );
nor ( n11698 , n11485 , n11518 );
nor ( n11699 , n11697 , n11698 );
nand ( n11700 , n11694 , n11699 );
and ( n11701 , n11700 , n11461 );
nor ( n11702 , n11398 , n11369 );
and ( n11703 , n11459 , n11702 );
not ( n11704 , n11423 );
nor ( n11705 , n11704 , n11458 );
nor ( n11706 , n11703 , n11705 );
or ( n11707 , n11706 , n11336 );
nor ( n11708 , n11264 , n11242 );
and ( n11709 , n11335 , n11708 );
not ( n11710 , n11296 );
nor ( n11711 , n11710 , n11334 );
nor ( n11712 , n11709 , n11711 );
nand ( n11713 , n11707 , n11712 );
nor ( n11714 , n11701 , n11713 );
nand ( n11715 , n11683 , n11714 );
not ( n11716 , n10628 );
nand ( n11717 , n11716 , n10648 );
nand ( n11718 , n278056 , n11717 );
nor ( n11719 , n278008 , n11718 );
and ( n11720 , n277900 , n11719 );
nand ( n11721 , n11715 , n277701 , n11720 );
nand ( n11722 , n10710 , n11721 );
not ( n11723 , n11722 );
buf ( n11724 , n11723 );
not ( n11725 , n11724 );
nand ( n11726 , n9189 , n11725 );
not ( n11727 , n9130 );
not ( n11728 , n11727 );
not ( n11729 , n9136 );
nand ( n11730 , n11728 , n11729 );
buf ( n11731 , n11730 );
not ( n11732 , n11731 );
and ( n11733 , n11732 , n9146 );
not ( n11734 , n11733 );
nand ( n11735 , n11734 , n11724 );
nand ( n11736 , n11726 , n11735 , n9163 );
not ( n11737 , n11736 );
nand ( n11738 , n11725 , n11733 );
nand ( n11739 , n11724 , n9149 );
and ( n11740 , n11738 , n11739 );
not ( n11741 , n9152 );
nand ( n11742 , n11741 , n9184 );
nor ( n11743 , n11740 , n11742 );
nor ( n11744 , n11737 , n11743 );
buf ( n11745 , n277356 );
not ( n11746 , n11745 );
not ( n11747 , n11746 );
buf ( n11748 , n9374 );
buf ( n11749 , n11748 );
not ( n11750 , n11749 );
or ( n11751 , n11747 , n11750 );
buf ( n11752 , n277501 );
not ( n11753 , n11752 );
buf ( n11754 , n277498 );
nand ( n11755 , n11753 , n11754 );
nand ( n11756 , n11751 , n11755 );
buf ( n11757 , n277411 );
not ( n11758 , n11757 );
not ( n11759 , n11758 );
buf ( n11760 , n277386 );
not ( n11761 , n11760 );
or ( n11762 , n11759 , n11761 );
buf ( n11763 , n277453 );
not ( n11764 , n11763 );
not ( n11765 , n277426 );
not ( n11766 , n11765 );
buf ( n11767 , n11766 );
nand ( n11768 , n11764 , n11767 );
nand ( n11769 , n11762 , n11768 );
nor ( n11770 , n11756 , n11769 );
not ( n11771 , n11770 );
buf ( n11772 , n277609 );
not ( n11773 , n11772 );
buf ( n11774 , n277575 );
buf ( n11775 , n11774 );
nand ( n11776 , n11773 , n11775 );
buf ( n11777 , n277533 );
not ( n11778 , n11777 );
buf ( n11779 , n277554 );
nand ( n11780 , n11778 , n11779 );
nand ( n11781 , n11776 , n11780 );
not ( n11782 , n11781 );
buf ( n11783 , n277649 );
not ( n11784 , n11783 );
buf ( n11785 , n277628 );
nand ( n11786 , n11784 , n11785 );
buf ( n11787 , n277696 );
not ( n11788 , n11787 );
buf ( n11789 , n277676 );
buf ( n11790 , n11789 );
nand ( n11791 , n11788 , n11790 );
and ( n11792 , n11786 , n11791 );
nand ( n11793 , n11782 , n11792 );
nor ( n11794 , n11771 , n11793 );
buf ( n11795 , n277749 );
not ( n11796 , n11795 );
not ( n11797 , n277718 );
buf ( n11798 , n11797 );
nand ( n11799 , n11796 , n11798 );
buf ( n11800 , n277798 );
not ( n11801 , n11800 );
buf ( n11802 , n277775 );
buf ( n11803 , n11802 );
nand ( n11804 , n11801 , n11803 );
and ( n11805 , n11799 , n11804 );
buf ( n11806 , n277896 );
not ( n11807 , n11806 );
buf ( n11808 , n277872 );
nand ( n11809 , n11807 , n11808 );
buf ( n11810 , n277822 );
not ( n11811 , n11810 );
buf ( n11812 , n277842 );
nand ( n11813 , n11811 , n11812 );
and ( n11814 , n11809 , n11813 );
nand ( n11815 , n11805 , n11814 );
buf ( n11816 , n277930 );
not ( n11817 , n11816 );
not ( n11818 , n11817 );
not ( n11819 , n277951 );
not ( n11820 , n11819 );
buf ( n11821 , n11820 );
not ( n11822 , n11821 );
or ( n11823 , n11818 , n11822 );
buf ( n11824 , n278005 );
not ( n11825 , n11824 );
buf ( n11826 , n277977 );
buf ( n11827 , n11826 );
nand ( n11828 , n11825 , n11827 );
nand ( n11829 , n11823 , n11828 );
not ( n11830 , n11829 );
buf ( n11831 , n278054 );
not ( n11832 , n11831 );
buf ( n11833 , n278025 );
buf ( n11834 , n11833 );
nand ( n11835 , n11832 , n11834 );
not ( n11836 , n11835 );
buf ( n11837 , n10627 );
not ( n11838 , n11837 );
buf ( n11839 , n10647 );
nor ( n11840 , n11838 , n11839 );
nor ( n11841 , n11836 , n11840 );
nand ( n11842 , n11830 , n11841 );
nor ( n11843 , n11815 , n11842 );
nand ( n11844 , n11794 , n11843 );
not ( n11845 , n11844 );
buf ( n11846 , n10921 );
buf ( n11847 , n11846 );
buf ( n11848 , n10961 );
buf ( n11849 , n11848 );
not ( n11850 , n11849 );
nand ( n11851 , n11847 , n11850 );
not ( n11852 , n10893 );
not ( n11853 , n11852 );
buf ( n11854 , n11853 );
not ( n11855 , n10861 );
buf ( n11856 , n11855 );
not ( n11857 , n11856 );
nor ( n11858 , n11854 , n11857 );
and ( n11859 , n11851 , n11858 );
nor ( n11860 , n11847 , n11850 );
nor ( n11861 , n11859 , n11860 );
buf ( n11862 , n10740 );
not ( n11863 , n11862 );
not ( n11864 , n11863 );
not ( n11865 , n10773 );
not ( n11866 , n11865 );
buf ( n11867 , n11866 );
not ( n11868 , n11867 );
or ( n11869 , n11864 , n11868 );
buf ( n11870 , n10836 );
not ( n11871 , n11870 );
buf ( n11872 , n10806 );
nand ( n11873 , n11871 , n11872 );
nand ( n11874 , n11869 , n11873 );
nor ( n11875 , n11861 , n11874 );
nor ( n11876 , n11867 , n11863 );
not ( n11877 , n11876 );
not ( n11878 , n11873 );
or ( n11879 , n11877 , n11878 );
not ( n11880 , n11872 );
nand ( n11881 , n11880 , n11870 );
nand ( n11882 , n11879 , n11881 );
nor ( n11883 , n11875 , n11882 );
not ( n11884 , n11857 );
not ( n11885 , n11854 );
or ( n11886 , n11884 , n11885 );
nand ( n11887 , n11886 , n11851 );
nor ( n11888 , n11874 , n11887 );
not ( n11889 , n10985 );
buf ( n11890 , n11889 );
not ( n11891 , n11890 );
not ( n11892 , n11891 );
buf ( n11893 , n11010 );
not ( n11894 , n11893 );
or ( n11895 , n11892 , n11894 );
buf ( n11896 , n11063 );
not ( n11897 , n11896 );
buf ( n11898 , n11046 );
nand ( n11899 , n11897 , n11898 );
nand ( n11900 , n11895 , n11899 );
not ( n11901 , n11893 );
nand ( n11902 , n11901 , n11890 );
nand ( n11903 , n11900 , n11902 );
not ( n11904 , n11097 );
not ( n11905 , n11904 );
buf ( n11906 , n11905 );
buf ( n11907 , n11122 );
buf ( n11908 , n11907 );
not ( n11909 , n11908 );
nand ( n11910 , n11906 , n11909 );
not ( n11911 , n11141 );
not ( n11912 , n11911 );
buf ( n11913 , n11912 );
buf ( n11914 , n11161 );
buf ( n11915 , n11914 );
not ( n11916 , n11915 );
nand ( n11917 , n11913 , n11916 );
nand ( n11918 , n11903 , n11910 , n11917 );
nor ( n11919 , n11913 , n11916 );
nor ( n11920 , n11906 , n11909 );
or ( n11921 , n11919 , n11920 );
nand ( n11922 , n11921 , n11910 );
nand ( n11923 , n11918 , n11922 );
nand ( n11924 , n11888 , n11923 );
and ( n11925 , n11883 , n11924 );
buf ( n11926 , n11241 );
not ( n11927 , n11926 );
not ( n11928 , n11927 );
not ( n11929 , n11262 );
not ( n11930 , n11929 );
buf ( n11931 , n11930 );
not ( n11932 , n11931 );
or ( n11933 , n11928 , n11932 );
buf ( n11934 , n11333 );
not ( n11935 , n11934 );
not ( n11936 , n11295 );
not ( n11937 , n11936 );
buf ( n11938 , n11937 );
nand ( n11939 , n11935 , n11938 );
nand ( n11940 , n11933 , n11939 );
buf ( n11941 , n11368 );
not ( n11942 , n11941 );
not ( n11943 , n11942 );
buf ( n11944 , n11396 );
not ( n11945 , n11944 );
or ( n11946 , n11943 , n11945 );
buf ( n11947 , n11457 );
not ( n11948 , n11947 );
buf ( n11949 , n11422 );
nand ( n11950 , n11948 , n11949 );
nand ( n11951 , n11946 , n11950 );
nor ( n11952 , n11940 , n11951 );
buf ( n11953 , n11516 );
buf ( n11954 , n11953 );
not ( n11955 , n11954 );
not ( n11956 , n11483 );
not ( n11957 , n11956 );
buf ( n11958 , n11957 );
nand ( n11959 , n11955 , n11958 );
buf ( n11960 , n11573 );
not ( n11961 , n11960 );
buf ( n11962 , n11543 );
nand ( n11963 , n11961 , n11962 );
nand ( n11964 , n11959 , n11963 );
buf ( n11965 , n11596 );
not ( n11966 , n11965 );
not ( n11967 , n11966 );
not ( n11968 , n11619 );
not ( n11969 , n11968 );
buf ( n11970 , n11969 );
not ( n11971 , n11970 );
or ( n11972 , n11967 , n11971 );
buf ( n11973 , n11677 );
not ( n11974 , n11973 );
buf ( n11975 , n11649 );
nand ( n11976 , n11974 , n11975 );
nand ( n11977 , n11972 , n11976 );
nor ( n11978 , n11964 , n11977 );
nand ( n11979 , n11952 , n11978 );
nor ( n11980 , n11925 , n11979 );
not ( n11981 , n11964 );
nor ( n11982 , n11970 , n11966 );
not ( n11983 , n11982 );
not ( n11984 , n11976 );
or ( n11985 , n11983 , n11984 );
not ( n11986 , n11975 );
nand ( n11987 , n11986 , n11973 );
nand ( n11988 , n11985 , n11987 );
and ( n11989 , n11981 , n11988 );
not ( n11990 , n11960 );
nor ( n11991 , n11990 , n11962 );
not ( n11992 , n11991 );
not ( n11993 , n11959 );
or ( n11994 , n11992 , n11993 );
not ( n11995 , n11958 );
nand ( n11996 , n11995 , n11954 );
nand ( n11997 , n11994 , n11996 );
nor ( n11998 , n11989 , n11997 );
not ( n11999 , n11952 );
or ( n12000 , n11998 , n11999 );
not ( n12001 , n11940 );
nor ( n12002 , n11944 , n11942 );
not ( n12003 , n12002 );
not ( n12004 , n11950 );
or ( n12005 , n12003 , n12004 );
not ( n12006 , n11949 );
nand ( n12007 , n12006 , n11947 );
nand ( n12008 , n12005 , n12007 );
and ( n12009 , n12001 , n12008 );
nor ( n12010 , n11931 , n11927 );
not ( n12011 , n12010 );
not ( n12012 , n11939 );
or ( n12013 , n12011 , n12012 );
not ( n12014 , n11938 );
nand ( n12015 , n12014 , n11934 );
nand ( n12016 , n12013 , n12015 );
nor ( n12017 , n12009 , n12016 );
nand ( n12018 , n12000 , n12017 );
nor ( n12019 , n11980 , n12018 );
not ( n12020 , n12019 );
and ( n12021 , n11845 , n12020 );
not ( n12022 , n11839 );
nor ( n12023 , n12022 , n11837 );
nand ( n12024 , n11835 , n12023 );
not ( n12025 , n11834 );
nand ( n12026 , n12025 , n11831 );
and ( n12027 , n12024 , n12026 );
nor ( n12028 , n12027 , n11829 );
nor ( n12029 , n11821 , n11817 );
not ( n12030 , n12029 );
not ( n12031 , n11828 );
or ( n12032 , n12030 , n12031 );
not ( n12033 , n11827 );
nand ( n12034 , n12033 , n11824 );
nand ( n12035 , n12032 , n12034 );
nor ( n12036 , n12028 , n12035 );
or ( n12037 , n12036 , n11815 );
not ( n12038 , n11810 );
nor ( n12039 , n12038 , n11812 );
not ( n12040 , n12039 );
not ( n12041 , n11809 );
or ( n12042 , n12040 , n12041 );
not ( n12043 , n11808 );
nand ( n12044 , n12043 , n11806 );
nand ( n12045 , n12042 , n12044 );
and ( n12046 , n11805 , n12045 );
not ( n12047 , n11800 );
nor ( n12048 , n12047 , n11803 );
not ( n12049 , n12048 );
not ( n12050 , n11799 );
or ( n12051 , n12049 , n12050 );
not ( n12052 , n11798 );
nand ( n12053 , n12052 , n11795 );
nand ( n12054 , n12051 , n12053 );
nor ( n12055 , n12046 , n12054 );
nand ( n12056 , n12037 , n12055 );
not ( n12057 , n12056 );
not ( n12058 , n11794 );
or ( n12059 , n12057 , n12058 );
not ( n12060 , n11787 );
nor ( n12061 , n12060 , n11790 );
and ( n12062 , n11786 , n12061 );
not ( n12063 , n11783 );
nor ( n12064 , n12063 , n11785 );
nor ( n12065 , n12062 , n12064 );
or ( n12066 , n12065 , n11781 );
not ( n12067 , n11777 );
nor ( n12068 , n12067 , n11779 );
and ( n12069 , n11776 , n12068 );
not ( n12070 , n11772 );
nor ( n12071 , n12070 , n11775 );
nor ( n12072 , n12069 , n12071 );
nand ( n12073 , n12066 , n12072 );
nand ( n12074 , n11770 , n12073 );
not ( n12075 , n11756 );
not ( n12076 , n11757 );
nor ( n12077 , n12076 , n11760 );
and ( n12078 , n11768 , n12077 );
not ( n12079 , n11763 );
nor ( n12080 , n12079 , n11767 );
nor ( n12081 , n12078 , n12080 );
not ( n12082 , n12081 );
and ( n12083 , n12075 , n12082 );
nor ( n12084 , n11749 , n11746 );
not ( n12085 , n12084 );
not ( n12086 , n11755 );
or ( n12087 , n12085 , n12086 );
or ( n12088 , n11753 , n11754 );
nand ( n12089 , n12087 , n12088 );
nor ( n12090 , n12083 , n12089 );
and ( n12091 , n12074 , n12090 );
nand ( n12092 , n12059 , n12091 );
nor ( n12093 , n12021 , n12092 );
buf ( n12094 , n12093 );
not ( n12095 , n12094 );
not ( n12096 , n9146 );
and ( n12097 , n9152 , n12096 );
nand ( n12098 , n12095 , n12097 );
not ( n12099 , n9152 );
not ( n12100 , n12099 );
nor ( n12101 , n12100 , n12096 );
not ( n12102 , n12101 );
not ( n12103 , n12102 );
nand ( n12104 , n12103 , n11725 );
and ( n12105 , n9151 , n9146 );
nand ( n12106 , n12094 , n12105 );
nand ( n12107 , n12099 , n12096 );
not ( n12108 , n12107 );
nand ( n12109 , n11724 , n12108 );
nand ( n12110 , n12098 , n12104 , n12106 , n12109 );
nor ( n12111 , n9130 , n9136 );
and ( n12112 , n12111 , n9184 );
nand ( n12113 , n12110 , n12112 );
and ( n12114 , n11744 , n12113 );
not ( n12115 , n9162 );
not ( n12116 , n12095 );
or ( n12117 , n12115 , n12116 );
not ( n12118 , n11741 );
nand ( n12119 , n11733 , n12118 );
not ( n12120 , n12119 );
nand ( n12121 , n12117 , n12120 );
not ( n12122 , n9155 );
and ( n12123 , n12121 , n12122 );
and ( n12124 , n12094 , n12119 );
nor ( n12125 , n12123 , n12124 );
buf ( n12126 , n10806 );
buf ( n12127 , n10836 );
not ( n12128 , n12127 );
and ( n12129 , n12126 , n12128 );
buf ( n12130 , n11677 );
not ( n12131 , n12130 );
and ( n12132 , n11649 , n12131 );
nor ( n12133 , n12129 , n12132 );
not ( n12134 , n11649 );
and ( n12135 , n12134 , n12130 );
not ( n12136 , n12126 );
and ( n12137 , n12136 , n12127 );
nor ( n12138 , n12135 , n12137 );
not ( n12139 , n11748 );
nand ( n12140 , n12139 , n277356 );
buf ( n12141 , n11889 );
buf ( n12142 , n11010 );
not ( n12143 , n12142 );
and ( n12144 , n12141 , n12143 );
not ( n12145 , n12141 );
and ( n12146 , n12145 , n12142 );
nor ( n12147 , n12144 , n12146 );
and ( n12148 , n12133 , n12138 , n12140 , n12147 );
not ( n12149 , n11936 );
not ( n12150 , n12149 );
not ( n12151 , n12150 );
not ( n12152 , n11333 );
not ( n12153 , n12152 );
not ( n12154 , n12153 );
and ( n12155 , n12151 , n12154 );
buf ( n12156 , n278005 );
not ( n12157 , n12156 );
and ( n12158 , n11826 , n12157 );
nor ( n12159 , n12155 , n12158 );
not ( n12160 , n277386 );
and ( n12161 , n277411 , n12160 );
not ( n12162 , n277411 );
and ( n12163 , n12162 , n277386 );
nor ( n12164 , n12161 , n12163 );
nand ( n12165 , n12159 , n12164 );
not ( n12166 , n277609 );
not ( n12167 , n12166 );
buf ( n12168 , n11774 );
not ( n12169 , n12168 );
or ( n12170 , n12167 , n12169 );
or ( n12171 , n12168 , n12166 );
nand ( n12172 , n12170 , n12171 );
not ( n12173 , n12153 );
not ( n12174 , n12149 );
not ( n12175 , n12174 );
or ( n12176 , n12173 , n12175 );
not ( n12177 , n11826 );
nand ( n12178 , n12177 , n12156 );
nand ( n12179 , n12176 , n12178 );
nor ( n12180 , n12165 , n12172 , n12179 );
nand ( n12181 , n12148 , n12180 );
buf ( n12182 , n277896 );
not ( n12183 , n12182 );
not ( n12184 , n277872 );
not ( n12185 , n12184 );
not ( n12186 , n12185 );
not ( n12187 , n12186 );
or ( n12188 , n12183 , n12187 );
not ( n12189 , n11904 );
not ( n12190 , n12189 );
not ( n12191 , n11907 );
not ( n12192 , n12191 );
nand ( n12193 , n12190 , n12192 );
nand ( n12194 , n12188 , n12193 );
not ( n12195 , n277696 );
not ( n12196 , n12195 );
not ( n12197 , n277676 );
not ( n12198 , n12197 );
not ( n12199 , n12198 );
or ( n12200 , n12196 , n12199 );
not ( n12201 , n277533 );
nand ( n12202 , n12201 , n277554 );
nand ( n12203 , n12200 , n12202 );
nor ( n12204 , n12194 , n12203 );
buf ( n12205 , n11241 );
not ( n12206 , n12205 );
not ( n12207 , n11929 );
not ( n12208 , n12207 );
not ( n12209 , n12208 );
or ( n12210 , n12206 , n12209 );
not ( n12211 , n12198 );
nand ( n12212 , n12211 , n277696 );
nand ( n12213 , n12210 , n12212 );
not ( n12214 , n277533 );
not ( n12215 , n277554 );
not ( n12216 , n12215 );
or ( n12217 , n12214 , n12216 );
not ( n12218 , n11396 );
not ( n12219 , n12218 );
buf ( n12220 , n11368 );
not ( n12221 , n12220 );
nand ( n12222 , n12219 , n12221 );
nand ( n12223 , n12217 , n12222 );
nor ( n12224 , n12213 , n12223 );
not ( n12225 , n277453 );
not ( n12226 , n11765 );
not ( n12227 , n12226 );
not ( n12228 , n12227 );
or ( n12229 , n12225 , n12228 );
not ( n12230 , n12182 );
nand ( n12231 , n12230 , n12185 );
nand ( n12232 , n12229 , n12231 );
buf ( n12233 , n11855 );
not ( n12234 , n12233 );
not ( n12235 , n12234 );
not ( n12236 , n11852 );
not ( n12237 , n12236 );
or ( n12238 , n12235 , n12237 );
not ( n12239 , n11956 );
not ( n12240 , n11953 );
nand ( n12241 , n12239 , n12240 );
nand ( n12242 , n12238 , n12241 );
nor ( n12243 , n12232 , n12242 );
not ( n12244 , n12219 );
and ( n12245 , n12244 , n12220 );
not ( n12246 , n277842 );
not ( n12247 , n12246 );
buf ( n12248 , n277822 );
not ( n12249 , n12248 );
and ( n12250 , n12247 , n12249 );
nor ( n12251 , n12245 , n12250 );
nand ( n12252 , n12204 , n12224 , n12243 , n12251 );
nor ( n12253 , n12181 , n12252 );
not ( n12254 , n11543 );
not ( n12255 , n12254 );
not ( n12256 , n12255 );
buf ( n12257 , n11573 );
not ( n12258 , n12257 );
not ( n12259 , n12258 );
and ( n12260 , n12256 , n12259 );
not ( n12261 , n12236 );
and ( n12262 , n12261 , n12233 );
nor ( n12263 , n12260 , n12262 );
buf ( n12264 , n11846 );
not ( n12265 , n12264 );
not ( n12266 , n11848 );
not ( n12267 , n12266 );
and ( n12268 , n12265 , n12267 );
not ( n12269 , n11968 );
not ( n12270 , n12269 );
buf ( n12271 , n11596 );
and ( n12272 , n12270 , n12271 );
nor ( n12273 , n12268 , n12272 );
not ( n12274 , n12269 );
not ( n12275 , n12274 );
not ( n12276 , n12271 );
and ( n12277 , n12275 , n12276 );
and ( n12278 , n12264 , n12266 );
nor ( n12279 , n12277 , n12278 );
buf ( n12280 , n11914 );
not ( n12281 , n11911 );
not ( n12282 , n12281 );
and ( n12283 , n12280 , n12282 );
not ( n12284 , n12280 );
and ( n12285 , n12284 , n12281 );
nor ( n12286 , n12283 , n12285 );
nand ( n12287 , n12263 , n12273 , n12279 , n12286 );
buf ( n12288 , n10627 );
not ( n12289 , n12288 );
buf ( n12290 , n10647 );
not ( n12291 , n12290 );
not ( n12292 , n12291 );
and ( n12293 , n12289 , n12292 );
buf ( n12294 , n11833 );
buf ( n12295 , n278054 );
not ( n12296 , n12295 );
and ( n12297 , n12294 , n12296 );
nor ( n12298 , n12293 , n12297 );
not ( n12299 , n12227 );
not ( n12300 , n277453 );
and ( n12301 , n12299 , n12300 );
buf ( n12302 , n11797 );
not ( n12303 , n277749 );
not ( n12304 , n12303 );
not ( n12305 , n12304 );
and ( n12306 , n12302 , n12305 );
nor ( n12307 , n12301 , n12306 );
not ( n12308 , n12239 );
not ( n12309 , n12240 );
and ( n12310 , n12308 , n12309 );
and ( n12311 , n12255 , n12258 );
nor ( n12312 , n12310 , n12311 );
not ( n12313 , n12302 );
nand ( n12314 , n12313 , n12304 );
nand ( n12315 , n12298 , n12307 , n12312 , n12314 );
buf ( n12316 , n11063 );
buf ( n12317 , n11046 );
buf ( n12318 , n12317 );
xor ( n12319 , n12316 , n12318 );
nor ( n12320 , n12287 , n12315 , n12319 );
not ( n12321 , n277501 );
not ( n12322 , n12321 );
xnor ( n12323 , n277498 , n12322 );
not ( n12324 , n12208 );
not ( n12325 , n12205 );
and ( n12326 , n12324 , n12325 );
not ( n12327 , n277356 );
and ( n12328 , n11748 , n12327 );
nor ( n12329 , n12326 , n12328 );
not ( n12330 , n12190 );
not ( n12331 , n12192 );
and ( n12332 , n12330 , n12331 );
not ( n12333 , n12247 );
and ( n12334 , n12333 , n12248 );
nor ( n12335 , n12332 , n12334 );
not ( n12336 , n10740 );
not ( n12337 , n11865 );
and ( n12338 , n12336 , n12337 );
not ( n12339 , n12336 );
not ( n12340 , n12337 );
and ( n12341 , n12339 , n12340 );
nor ( n12342 , n12338 , n12341 );
nand ( n12343 , n12323 , n12329 , n12335 , n12342 );
not ( n12344 , n12288 );
not ( n12345 , n12344 );
not ( n12346 , n12290 );
and ( n12347 , n12345 , n12346 );
not ( n12348 , n12294 );
and ( n12349 , n12348 , n12295 );
nor ( n12350 , n12347 , n12349 );
buf ( n12351 , n11422 );
not ( n12352 , n12351 );
buf ( n12353 , n11457 );
and ( n12354 , n12352 , n12353 );
not ( n12355 , n11819 );
not ( n12356 , n12355 );
buf ( n12357 , n277930 );
and ( n12358 , n12356 , n12357 );
nor ( n12359 , n12354 , n12358 );
not ( n12360 , n12353 );
and ( n12361 , n12351 , n12360 );
not ( n12362 , n12357 );
and ( n12363 , n12355 , n12362 );
nor ( n12364 , n12361 , n12363 );
buf ( n12365 , n277649 );
xnor ( n12366 , n12365 , n277628 );
nand ( n12367 , n12350 , n12359 , n12364 , n12366 );
nor ( n12368 , n12343 , n12367 );
buf ( n12369 , n277798 );
buf ( n12370 , n12369 );
buf ( n12371 , n11802 );
xnor ( n12372 , n12370 , n12371 );
nand ( n12373 , n12253 , n12320 , n12368 , n12372 );
buf ( n12374 , n12373 );
not ( n12375 , n12374 );
nand ( n12376 , n9130 , n9136 );
not ( n12377 , n12376 );
nand ( n12378 , n12377 , n12101 );
or ( n12379 , n12375 , n12378 );
nand ( n12380 , n12378 , n9153 );
nand ( n12381 , n12380 , n9163 );
nand ( n12382 , n12379 , n12381 );
or ( n12383 , n12125 , n12382 );
nand ( n12384 , n12383 , n9184 );
buf ( n12385 , n277356 );
not ( n12386 , n12385 );
buf ( n12387 , n11748 );
not ( n12388 , n12387 );
not ( n12389 , n12388 );
or ( n12390 , n12386 , n12389 );
not ( n12391 , n12321 );
buf ( n12392 , n12391 );
buf ( n12393 , n277498 );
not ( n12394 , n12393 );
nand ( n12395 , n12392 , n12394 );
nand ( n12396 , n12390 , n12395 );
buf ( n12397 , n277411 );
not ( n12398 , n12397 );
buf ( n12399 , n277386 );
not ( n12400 , n12399 );
not ( n12401 , n12400 );
or ( n12402 , n12398 , n12401 );
buf ( n12403 , n12226 );
not ( n12404 , n12403 );
buf ( n12405 , n277453 );
nand ( n12406 , n12404 , n12405 );
nand ( n12407 , n12402 , n12406 );
nor ( n12408 , n12396 , n12407 );
buf ( n12409 , n277533 );
not ( n12410 , n12409 );
buf ( n12411 , n277554 );
not ( n12412 , n12411 );
not ( n12413 , n12412 );
or ( n12414 , n12410 , n12413 );
buf ( n12415 , n277575 );
buf ( n12416 , n12415 );
not ( n12417 , n12416 );
buf ( n12418 , n277609 );
nand ( n12419 , n12417 , n12418 );
nand ( n12420 , n12414 , n12419 );
buf ( n12421 , n277628 );
not ( n12422 , n12421 );
buf ( n12423 , n12365 );
nand ( n12424 , n12422 , n12423 );
not ( n12425 , n12197 );
buf ( n12426 , n12425 );
not ( n12427 , n12426 );
buf ( n12428 , n277696 );
nand ( n12429 , n12427 , n12428 );
nand ( n12430 , n12424 , n12429 );
nor ( n12431 , n12420 , n12430 );
nand ( n12432 , n12408 , n12431 );
buf ( n12433 , n12369 );
not ( n12434 , n12433 );
buf ( n12435 , n11802 );
not ( n12436 , n12435 );
not ( n12437 , n12436 );
or ( n12438 , n12434 , n12437 );
buf ( n12439 , n11797 );
not ( n12440 , n12439 );
not ( n12441 , n12303 );
buf ( n12442 , n12441 );
nand ( n12443 , n12440 , n12442 );
nand ( n12444 , n12438 , n12443 );
not ( n12445 , n12184 );
buf ( n12446 , n12445 );
not ( n12447 , n12446 );
buf ( n12448 , n277896 );
buf ( n12449 , n12448 );
nand ( n12450 , n12447 , n12449 );
not ( n12451 , n12246 );
buf ( n12452 , n12451 );
not ( n12453 , n12452 );
buf ( n12454 , n12248 );
nand ( n12455 , n12453 , n12454 );
nand ( n12456 , n12450 , n12455 );
nor ( n12457 , n12444 , n12456 );
buf ( n12458 , n12357 );
not ( n12459 , n12458 );
not ( n12460 , n11819 );
buf ( n12461 , n12460 );
not ( n12462 , n12461 );
not ( n12463 , n12462 );
or ( n12464 , n12459 , n12463 );
buf ( n12465 , n11826 );
not ( n12466 , n12465 );
buf ( n12467 , n12156 );
nand ( n12468 , n12466 , n12467 );
nand ( n12469 , n12464 , n12468 );
buf ( n12470 , n12290 );
not ( n12471 , n12470 );
buf ( n12472 , n10627 );
not ( n12473 , n12472 );
not ( n12474 , n12473 );
or ( n12475 , n12471 , n12474 );
buf ( n12476 , n11833 );
not ( n12477 , n12476 );
buf ( n12478 , n12295 );
nand ( n12479 , n12477 , n12478 );
nand ( n12480 , n12475 , n12479 );
nor ( n12481 , n12469 , n12480 );
nand ( n12482 , n12457 , n12481 );
nor ( n12483 , n12432 , n12482 );
buf ( n12484 , n10740 );
not ( n12485 , n12484 );
buf ( n12486 , n12337 );
not ( n12487 , n12486 );
not ( n12488 , n12487 );
or ( n12489 , n12485 , n12488 );
buf ( n12490 , n12126 );
not ( n12491 , n12490 );
buf ( n12492 , n12127 );
nand ( n12493 , n12491 , n12492 );
nand ( n12494 , n12489 , n12493 );
buf ( n12495 , n11846 );
not ( n12496 , n12495 );
buf ( n12497 , n11848 );
nand ( n12498 , n12496 , n12497 );
buf ( n12499 , n12236 );
not ( n12500 , n12499 );
buf ( n12501 , n12233 );
nand ( n12502 , n12500 , n12501 );
nand ( n12503 , n12498 , n12502 );
nor ( n12504 , n12494 , n12503 );
buf ( n12505 , n12189 );
not ( n12506 , n12505 );
not ( n12507 , n12191 );
buf ( n12508 , n12507 );
nand ( n12509 , n12506 , n12508 );
not ( n12510 , n12509 );
buf ( n12511 , n11914 );
not ( n12512 , n12511 );
not ( n12513 , n12512 );
buf ( n12514 , n12281 );
not ( n12515 , n12514 );
or ( n12516 , n12513 , n12515 );
not ( n12517 , n12508 );
nand ( n12518 , n12517 , n12505 );
nand ( n12519 , n12516 , n12518 );
not ( n12520 , n12519 );
or ( n12521 , n12510 , n12520 );
buf ( n12522 , n12141 );
not ( n12523 , n12522 );
not ( n12524 , n12523 );
buf ( n12525 , n12142 );
not ( n12526 , n12525 );
or ( n12527 , n12524 , n12526 );
not ( n12528 , n12522 );
not ( n12529 , n12525 );
not ( n12530 , n12529 );
or ( n12531 , n12528 , n12530 );
buf ( n12532 , n12317 );
not ( n12533 , n12532 );
buf ( n12534 , n12316 );
nand ( n12535 , n12533 , n12534 );
nand ( n12536 , n12531 , n12535 );
nand ( n12537 , n12527 , n12536 );
not ( n12538 , n12514 );
nand ( n12539 , n12538 , n12511 );
nand ( n12540 , n12537 , n12509 , n12539 );
nand ( n12541 , n12521 , n12540 );
and ( n12542 , n12504 , n12541 );
nor ( n12543 , n12500 , n12501 );
and ( n12544 , n12498 , n12543 );
nor ( n12545 , n12496 , n12497 );
nor ( n12546 , n12544 , n12545 );
or ( n12547 , n12546 , n12494 );
nor ( n12548 , n12487 , n12484 );
and ( n12549 , n12493 , n12548 );
nor ( n12550 , n12491 , n12492 );
nor ( n12551 , n12549 , n12550 );
nand ( n12552 , n12547 , n12551 );
nor ( n12553 , n12542 , n12552 );
buf ( n12554 , n12205 );
not ( n12555 , n12554 );
buf ( n12556 , n12207 );
not ( n12557 , n12556 );
not ( n12558 , n12557 );
or ( n12559 , n12555 , n12558 );
buf ( n12560 , n12149 );
not ( n12561 , n12560 );
not ( n12562 , n12152 );
buf ( n12563 , n12562 );
nand ( n12564 , n12561 , n12563 );
nand ( n12565 , n12559 , n12564 );
buf ( n12566 , n12351 );
not ( n12567 , n12566 );
buf ( n12568 , n12353 );
nand ( n12569 , n12567 , n12568 );
not ( n12570 , n12218 );
buf ( n12571 , n12570 );
not ( n12572 , n12571 );
buf ( n12573 , n12220 );
nand ( n12574 , n12572 , n12573 );
nand ( n12575 , n12569 , n12574 );
nor ( n12576 , n12565 , n12575 );
buf ( n12577 , n12257 );
not ( n12578 , n12577 );
not ( n12579 , n12254 );
buf ( n12580 , n12579 );
not ( n12581 , n12580 );
not ( n12582 , n12581 );
or ( n12583 , n12578 , n12582 );
buf ( n12584 , n12239 );
not ( n12585 , n12584 );
buf ( n12586 , n11953 );
nand ( n12587 , n12585 , n12586 );
nand ( n12588 , n12583 , n12587 );
buf ( n12589 , n12271 );
not ( n12590 , n12589 );
buf ( n12591 , n12269 );
not ( n12592 , n12591 );
not ( n12593 , n12592 );
or ( n12594 , n12590 , n12593 );
buf ( n12595 , n11649 );
not ( n12596 , n12595 );
buf ( n12597 , n12130 );
nand ( n12598 , n12596 , n12597 );
nand ( n12599 , n12594 , n12598 );
nor ( n12600 , n12588 , n12599 );
nand ( n12601 , n12576 , n12600 );
or ( n12602 , n12553 , n12601 );
nor ( n12603 , n12592 , n12589 );
and ( n12604 , n12598 , n12603 );
nor ( n12605 , n12596 , n12597 );
nor ( n12606 , n12604 , n12605 );
or ( n12607 , n12606 , n12588 );
nor ( n12608 , n12581 , n12577 );
and ( n12609 , n12587 , n12608 );
nor ( n12610 , n12585 , n12586 );
nor ( n12611 , n12609 , n12610 );
nand ( n12612 , n12607 , n12611 );
and ( n12613 , n12612 , n12576 );
nor ( n12614 , n12572 , n12573 );
and ( n12615 , n12569 , n12614 );
nor ( n12616 , n12567 , n12568 );
nor ( n12617 , n12615 , n12616 );
or ( n12618 , n12617 , n12565 );
nor ( n12619 , n12557 , n12554 );
and ( n12620 , n12564 , n12619 );
nor ( n12621 , n12561 , n12563 );
nor ( n12622 , n12620 , n12621 );
nand ( n12623 , n12618 , n12622 );
nor ( n12624 , n12613 , n12623 );
nand ( n12625 , n12602 , n12624 );
and ( n12626 , n12483 , n12625 );
nor ( n12627 , n12473 , n12470 );
and ( n12628 , n12479 , n12627 );
nor ( n12629 , n12477 , n12478 );
nor ( n12630 , n12628 , n12629 );
or ( n12631 , n12630 , n12469 );
nor ( n12632 , n12462 , n12458 );
and ( n12633 , n12468 , n12632 );
nor ( n12634 , n12466 , n12467 );
nor ( n12635 , n12633 , n12634 );
nand ( n12636 , n12631 , n12635 );
and ( n12637 , n12636 , n12457 );
nor ( n12638 , n12453 , n12454 );
and ( n12639 , n12450 , n12638 );
nor ( n12640 , n12447 , n12449 );
nor ( n12641 , n12639 , n12640 );
or ( n12642 , n12641 , n12444 );
nor ( n12643 , n12436 , n12433 );
and ( n12644 , n12443 , n12643 );
nor ( n12645 , n12440 , n12442 );
nor ( n12646 , n12644 , n12645 );
nand ( n12647 , n12642 , n12646 );
nor ( n12648 , n12637 , n12647 );
or ( n12649 , n12432 , n12648 );
not ( n12650 , n12426 );
nor ( n12651 , n12650 , n12428 );
and ( n12652 , n12424 , n12651 );
nor ( n12653 , n12422 , n12423 );
nor ( n12654 , n12652 , n12653 );
or ( n12655 , n12654 , n12420 );
not ( n12656 , n12409 );
nand ( n12657 , n12656 , n12419 , n12411 );
not ( n12658 , n12418 );
nand ( n12659 , n12658 , n12416 );
and ( n12660 , n12657 , n12659 );
nand ( n12661 , n12655 , n12660 );
and ( n12662 , n12408 , n12661 );
nor ( n12663 , n12400 , n12397 );
and ( n12664 , n12406 , n12663 );
nor ( n12665 , n12404 , n12405 );
nor ( n12666 , n12664 , n12665 );
or ( n12667 , n12396 , n12666 );
nor ( n12668 , n12388 , n12385 );
and ( n12669 , n12395 , n12668 );
nor ( n12670 , n12392 , n12394 );
nor ( n12671 , n12669 , n12670 );
nand ( n12672 , n12667 , n12671 );
nor ( n12673 , n12662 , n12672 );
nand ( n12674 , n12649 , n12673 );
nor ( n12675 , n12626 , n12674 );
buf ( n12676 , n12675 );
nand ( n12677 , n12676 , n12097 );
not ( n12678 , n12677 );
not ( n12679 , n12105 );
or ( n12680 , n12676 , n12679 );
not ( n12681 , n12373 );
nand ( n12682 , n12681 , n12108 );
nand ( n12683 , n12680 , n12682 );
nor ( n12684 , n12678 , n12683 );
not ( n12685 , n9135 );
nand ( n12686 , n12685 , n9129 );
buf ( n12687 , n12686 );
not ( n12688 , n12687 );
nor ( n12689 , n12377 , n12688 );
or ( n12690 , n12684 , n12689 );
nor ( n12691 , n12687 , n12102 );
and ( n12692 , n12374 , n12691 );
nor ( n12693 , n12376 , n9162 );
nor ( n12694 , n12692 , n12693 );
nand ( n12695 , n12690 , n12694 );
nand ( n12696 , n12695 , n9184 );
nand ( n12697 , n9186 , n12114 , n12384 , n12696 );
buf ( n12698 , n12697 );
buf ( n12699 , n12698 );
not ( n12700 , n275925 );
buf ( n12701 , n12700 );
buf ( n12702 , n12701 );
buf ( n12703 , RI21a14440_60);
not ( n12704 , n12703 );
not ( n12705 , n12704 );
buf ( n12706 , n12705 );
not ( n12707 , n12706 );
buf ( n12708 , RI21a15f70_44);
buf ( n12709 , n12708 );
buf ( n12710 , n12709 );
and ( n12711 , n12707 , n12710 );
not ( n12712 , n12707 );
buf ( n12713 , RI21a14350_62);
buf ( n12714 , n12713 );
buf ( n12715 , n12714 );
not ( n12716 , n12715 );
not ( n12717 , n12716 );
buf ( n12718 , RI21a13ae0_66);
buf ( n12719 , n12718 );
buf ( n12720 , n12719 );
buf ( n12721 , n12720 );
nor ( n12722 , n12717 , n12721 );
buf ( n12723 , RI21a13b58_65);
buf ( n12724 , n12723 );
buf ( n12725 , n12724 );
buf ( n12726 , RI21a168d0_38);
buf ( n12727 , n12726 );
buf ( n12728 , n12727 );
buf ( n12729 , n12728 );
nor ( n12730 , n12725 , n12729 );
nand ( n12731 , n12722 , n12730 );
buf ( n12732 , RI21a13bd0_64);
buf ( n12733 , n12732 );
buf ( n12734 , n12733 );
buf ( n12735 , RI21a16948_37);
buf ( n12736 , n12735 );
buf ( n12737 , n12736 );
buf ( n12738 , n12737 );
nor ( n12739 , n12734 , n12738 );
buf ( n12740 , RI21a169c0_36);
not ( n12741 , n12740 );
not ( n12742 , n12741 );
buf ( n12743 , n12742 );
buf ( n12744 , n12743 );
not ( n12745 , n12744 );
buf ( n12746 , RI21a15778_47);
buf ( n12747 , n12746 );
buf ( n12748 , n12747 );
buf ( n12749 , n12748 );
buf ( n12750 , RI21a15fe8_43);
buf ( n12751 , n12750 );
buf ( n12752 , n12751 );
nor ( n12753 , n12749 , n12752 );
nand ( n12754 , n12739 , n12745 , n12753 );
nor ( n12755 , n12731 , n12754 );
buf ( n12756 , RI21a16150_40);
buf ( n12757 , n12756 );
buf ( n12758 , n12757 );
buf ( n12759 , RI21a143c8_61);
buf ( n12760 , n12759 );
buf ( n12761 , n12760 );
nor ( n12762 , n12758 , n12761 );
buf ( n12763 , RI21a161c8_39);
buf ( n12764 , n12763 );
buf ( n12765 , n12764 );
buf ( n12766 , RI21a14530_58);
buf ( n12767 , n12766 );
buf ( n12768 , n12767 );
nor ( n12769 , n12765 , n12768 );
nand ( n12770 , n12762 , n12769 );
buf ( n12771 , RI21a16060_42);
buf ( n12772 , n12771 );
buf ( n12773 , n12772 );
buf ( n12774 , RI21a160d8_41);
buf ( n12775 , n12774 );
buf ( n12776 , n12775 );
nor ( n12777 , n12773 , n12776 );
buf ( n12778 , RI21a13a68_67);
buf ( n12779 , n12778 );
buf ( n12780 , n12779 );
buf ( n12781 , RI21a13c48_63);
buf ( n12782 , n12781 );
buf ( n12783 , n12782 );
nor ( n12784 , n12780 , n12783 );
nand ( n12785 , n12777 , n12784 );
nor ( n12786 , n12770 , n12785 );
buf ( n12787 , n12786 );
nand ( n12788 , n12755 , n12787 );
buf ( n12789 , n12709 );
buf ( n12790 , n12789 );
and ( n12791 , n12788 , n12790 );
not ( n12792 , n12788 );
not ( n12793 , n12790 );
and ( n12794 , n12792 , n12793 );
nor ( n12795 , n12791 , n12794 );
buf ( n12796 , n12795 );
and ( n12797 , n12712 , n12796 );
nor ( n12798 , n12711 , n12797 );
not ( n12799 , n12798 );
buf ( n12800 , n12707 );
not ( n12801 , n12800 );
not ( n12802 , n12801 );
buf ( n12803 , n12752 );
nor ( n12804 , n12743 , n12748 );
not ( n12805 , n12804 );
nor ( n12806 , n12734 , n12715 );
nor ( n12807 , n12728 , n12737 );
nor ( n12808 , n12725 , n12720 );
nand ( n12809 , n12806 , n12807 , n12808 );
nor ( n12810 , n12805 , n12809 );
nand ( n12811 , n12786 , n12810 );
buf ( n12812 , n12811 );
and ( n12813 , n12803 , n12812 );
not ( n12814 , n12803 );
not ( n12815 , n12811 );
buf ( n12816 , n12815 );
and ( n12817 , n12814 , n12816 );
nor ( n12818 , n12813 , n12817 );
buf ( n12819 , n12818 );
not ( n12820 , n12819 );
or ( n12821 , n12802 , n12820 );
nand ( n12822 , n12800 , n12751 );
nand ( n12823 , n12821 , n12822 );
nor ( n12824 , n12799 , n12823 );
not ( n12825 , n12800 );
not ( n12826 , n12825 );
not ( n12827 , n12773 );
not ( n12828 , n12827 );
nor ( n12829 , n12743 , n12748 );
nor ( n12830 , n12768 , n12761 );
nand ( n12831 , n12829 , n12830 );
not ( n12832 , n12831 );
not ( n12833 , n12783 );
nand ( n12834 , n12833 , n12716 );
not ( n12835 , n12725 );
not ( n12836 , n12734 );
nand ( n12837 , n12835 , n12836 );
nor ( n12838 , n12834 , n12837 );
nand ( n12839 , n12832 , n12838 );
not ( n12840 , n12839 );
buf ( n12841 , n12780 );
not ( n12842 , n12841 );
not ( n12843 , n12721 );
nand ( n12844 , n12842 , n12843 );
not ( n12845 , n12807 );
nor ( n12846 , n12844 , n12845 );
not ( n12847 , n12758 );
not ( n12848 , n12765 );
nand ( n12849 , n12847 , n12848 );
buf ( n12850 , n12776 );
nor ( n12851 , n12849 , n12850 );
and ( n12852 , n12846 , n12851 );
nand ( n12853 , n12840 , n12852 );
not ( n12854 , n12853 );
or ( n12855 , n12828 , n12854 );
nand ( n12856 , n12840 , n12852 );
or ( n12857 , n12856 , n12827 );
nand ( n12858 , n12855 , n12857 );
buf ( n12859 , n12858 );
not ( n12860 , n12859 );
or ( n12861 , n12826 , n12860 );
nand ( n12862 , n12800 , n12772 );
nand ( n12863 , n12861 , n12862 );
not ( n12864 , n12863 );
not ( n12865 , n12801 );
nor ( n12866 , n12789 , n12752 );
buf ( n12867 , n12866 );
not ( n12868 , n12867 );
not ( n12869 , n12868 );
nand ( n12870 , n12810 , n12786 );
not ( n12871 , n12870 );
nand ( n12872 , n12869 , n12871 );
buf ( n12873 , RI21a15868_45);
buf ( n12874 , n12873 );
buf ( n12875 , n12874 );
not ( n12876 , n12875 );
xnor ( n12877 , n12872 , n12876 );
buf ( n12878 , n12877 );
not ( n12879 , n12878 );
or ( n12880 , n12865 , n12879 );
nand ( n12881 , n12800 , n12874 );
nand ( n12882 , n12880 , n12881 );
not ( n12883 , n12882 );
nand ( n12884 , n12824 , n12864 , n12883 );
not ( n12885 , n12706 );
not ( n12886 , n12885 );
not ( n12887 , n12886 );
buf ( n12888 , RI21a15688_49);
buf ( n12889 , n12888 );
buf ( n12890 , n12889 );
buf ( n12891 , RI21a15700_48);
buf ( n12892 , n12891 );
buf ( n12893 , n12892 );
nor ( n12894 , n12890 , n12893 );
not ( n12895 , n12894 );
buf ( n12896 , RI21a157f0_46);
buf ( n12897 , n12896 );
buf ( n12898 , n12897 );
nor ( n12899 , n12898 , n12875 );
nand ( n12900 , n12899 , n12866 );
nor ( n12901 , n12895 , n12900 );
nand ( n12902 , n12871 , n12901 );
buf ( n12903 , RI21a15610_50);
buf ( n12904 , n12903 );
buf ( n12905 , n12904 );
not ( n12906 , n12905 );
xnor ( n12907 , n12902 , n12906 );
buf ( n12908 , n12907 );
not ( n12909 , n12908 );
or ( n12910 , n12887 , n12909 );
nand ( n12911 , n12885 , n12904 );
nand ( n12912 , n12910 , n12911 );
not ( n12913 , n12912 );
not ( n12914 , n12706 );
buf ( n12915 , n12724 );
and ( n12916 , n12914 , n12915 );
not ( n12917 , n12914 );
not ( n12918 , n12725 );
not ( n12919 , n12918 );
not ( n12920 , n12783 );
nand ( n12921 , n12920 , n12716 );
not ( n12922 , n12734 );
not ( n12923 , n12922 );
nor ( n12924 , n12921 , n12923 );
nand ( n12925 , n12832 , n12924 );
not ( n12926 , n12925 );
or ( n12927 , n12919 , n12926 );
buf ( n12928 , n12831 );
not ( n12929 , n12928 );
nand ( n12930 , n12929 , n12924 );
or ( n12931 , n12930 , n12918 );
nand ( n12932 , n12927 , n12931 );
buf ( n12933 , n12932 );
and ( n12934 , n12917 , n12933 );
nor ( n12935 , n12916 , n12934 );
not ( n12936 , n12935 );
not ( n12937 , n12936 );
buf ( n12938 , n12893 );
nor ( n12939 , n12900 , n12938 );
nand ( n12940 , n12871 , n12939 );
not ( n12941 , n12890 );
xnor ( n12942 , n12940 , n12941 );
buf ( n12943 , n12942 );
not ( n12944 , n12943 );
or ( n12945 , n12944 , n12800 );
nand ( n12946 , n12800 , n12889 );
nand ( n12947 , n12945 , n12946 );
buf ( n12948 , n12892 );
and ( n12949 , n12707 , n12948 );
not ( n12950 , n12707 );
not ( n12951 , n12900 );
not ( n12952 , n12951 );
not ( n12953 , n12815 );
or ( n12954 , n12952 , n12953 );
not ( n12955 , n12938 );
nand ( n12956 , n12954 , n12955 );
not ( n12957 , n12749 );
and ( n12958 , n12957 , n12938 );
nand ( n12959 , n12745 , n12769 , n12958 );
buf ( n12960 , n12785 );
nor ( n12961 , n12959 , n12960 );
nor ( n12962 , n12717 , n12721 );
and ( n12963 , n12962 , n12730 , n12739 );
and ( n12964 , n12762 , n12867 , n12899 );
nand ( n12965 , n12961 , n12963 , n12964 );
nand ( n12966 , n12956 , n12965 );
buf ( n12967 , n12966 );
and ( n12968 , n12950 , n12967 );
nor ( n12969 , n12949 , n12968 );
not ( n12970 , n12969 );
nor ( n12971 , n12947 , n12970 );
not ( n12972 , n12825 );
not ( n12973 , n12876 );
nor ( n12974 , n12973 , n12868 );
nand ( n12975 , n12871 , n12974 );
not ( n12976 , n12898 );
xnor ( n12977 , n12975 , n12976 );
buf ( n12978 , n12977 );
not ( n12979 , n12978 );
or ( n12980 , n12972 , n12979 );
nand ( n12981 , n12885 , n12897 );
nand ( n12982 , n12980 , n12981 );
not ( n12983 , n12982 );
nand ( n12984 , n12913 , n12937 , n12971 , n12983 );
nor ( n12985 , n12884 , n12984 );
not ( n12986 , n12825 );
not ( n12987 , n12738 );
not ( n12988 , n12987 );
buf ( n12989 , n12844 );
nor ( n12990 , n12988 , n12989 );
nand ( n12991 , n12840 , n12990 );
and ( n12992 , n12991 , n12729 );
not ( n12993 , n12991 );
not ( n12994 , n12729 );
and ( n12995 , n12993 , n12994 );
nor ( n12996 , n12992 , n12995 );
buf ( n12997 , n12996 );
not ( n12998 , n12997 );
not ( n12999 , n12998 );
not ( n13000 , n12999 );
or ( n13001 , n12986 , n13000 );
nand ( n13002 , n12885 , n12727 );
nand ( n13003 , n13001 , n13002 );
not ( n13004 , n13003 );
not ( n13005 , n12922 );
not ( n13006 , n12921 );
nand ( n13007 , n12929 , n13006 );
not ( n13008 , n13007 );
or ( n13009 , n13005 , n13008 );
not ( n13010 , n12923 );
or ( n13011 , n13007 , n13010 );
nand ( n13012 , n13009 , n13011 );
buf ( n13013 , n13012 );
and ( n13014 , n12706 , n13013 );
not ( n13015 , n12706 );
buf ( n13016 , n12733 );
and ( n13017 , n13015 , n13016 );
nor ( n13018 , n13014 , n13017 );
not ( n13019 , n13018 );
not ( n13020 , n13019 );
buf ( n13021 , n12782 );
and ( n13022 , n12914 , n13021 );
not ( n13023 , n12914 );
nand ( n13024 , n12832 , n12716 );
not ( n13025 , n12920 );
and ( n13026 , n13024 , n13025 );
not ( n13027 , n13024 );
and ( n13028 , n13027 , n12920 );
nor ( n13029 , n13026 , n13028 );
buf ( n13030 , n13029 );
and ( n13031 , n13023 , n13030 );
nor ( n13032 , n13022 , n13031 );
not ( n13033 , n13032 );
not ( n13034 , n13033 );
not ( n13035 , n12705 );
buf ( n13036 , n12714 );
and ( n13037 , n13035 , n13036 );
not ( n13038 , n13035 );
not ( n13039 , n12717 );
not ( n13040 , n12928 );
not ( n13041 , n13040 );
or ( n13042 , n13039 , n13041 );
not ( n13043 , n12928 );
or ( n13044 , n13043 , n12717 );
nand ( n13045 , n13042 , n13044 );
buf ( n13046 , n13045 );
and ( n13047 , n13038 , n13046 );
nor ( n13048 , n13037 , n13047 );
not ( n13049 , n13048 );
buf ( n13050 , n12761 );
not ( n13051 , n13050 );
not ( n13052 , n13051 );
buf ( n13053 , n12804 );
buf ( n13054 , n12768 );
not ( n13055 , n13054 );
nand ( n13056 , n13053 , n13055 );
not ( n13057 , n13056 );
or ( n13058 , n13052 , n13057 );
or ( n13059 , n13056 , n13051 );
nand ( n13060 , n13058 , n13059 );
buf ( n13061 , n13060 );
and ( n13062 , n12705 , n13061 );
not ( n13063 , n12705 );
buf ( n13064 , n12760 );
and ( n13065 , n13063 , n13064 );
nor ( n13066 , n13062 , n13065 );
not ( n13067 , n13066 );
nor ( n13068 , n13049 , n13067 );
and ( n13069 , n13020 , n13034 , n13068 );
not ( n13070 , n12705 );
not ( n13071 , n13055 );
not ( n13072 , n13053 );
not ( n13073 , n13072 );
or ( n13074 , n13071 , n13073 );
or ( n13075 , n13072 , n13055 );
nand ( n13076 , n13074 , n13075 );
buf ( n13077 , n13076 );
not ( n13078 , n13077 );
or ( n13079 , n13070 , n13078 );
not ( n13080 , n12705 );
buf ( n13081 , n12767 );
nand ( n13082 , n13080 , n13081 );
nand ( n13083 , n13079 , n13082 );
buf ( n13084 , n13083 );
not ( n13085 , n12705 );
not ( n13086 , n12749 );
not ( n13087 , n12745 );
or ( n13088 , n13086 , n13087 );
not ( n13089 , n12749 );
nand ( n13090 , n13089 , n12744 );
nand ( n13091 , n13088 , n13090 );
buf ( n13092 , n13091 );
not ( n13093 , n13092 );
or ( n13094 , n13085 , n13093 );
not ( n13095 , n12705 );
buf ( n13096 , n12747 );
nand ( n13097 , n13095 , n13096 );
nand ( n13098 , n13094 , n13097 );
buf ( n13099 , n13098 );
not ( n13100 , n13099 );
buf ( n13101 , n12742 );
buf ( n13102 , n13101 );
not ( n13103 , n13102 );
nand ( n13104 , n13100 , n13103 );
nor ( n13105 , n13084 , n13104 );
nand ( n13106 , n13004 , n13069 , n13105 );
not ( n13107 , n12825 );
not ( n13108 , n12987 );
not ( n13109 , n12989 );
nand ( n13110 , n12840 , n13109 );
not ( n13111 , n13110 );
or ( n13112 , n13108 , n13111 );
nand ( n13113 , n12840 , n13109 );
or ( n13114 , n13113 , n12987 );
nand ( n13115 , n13112 , n13114 );
buf ( n13116 , n13115 );
not ( n13117 , n13116 );
or ( n13118 , n13107 , n13117 );
nand ( n13119 , n12800 , n12736 );
nand ( n13120 , n13118 , n13119 );
not ( n13121 , n13120 );
not ( n13122 , n12801 );
not ( n13123 , n12841 );
not ( n13124 , n12957 );
nor ( n13125 , n13124 , n13054 );
nor ( n13126 , n13025 , n12721 );
nand ( n13127 , n12745 , n13125 , n13126 );
not ( n13128 , n12918 );
nor ( n13129 , n13050 , n13128 );
nand ( n13130 , n12806 , n13129 );
nor ( n13131 , n13127 , n13130 );
not ( n13132 , n13131 );
or ( n13133 , n13123 , n13132 );
or ( n13134 , n13131 , n12841 );
nand ( n13135 , n13133 , n13134 );
buf ( n13136 , n13135 );
not ( n13137 , n13136 );
or ( n13138 , n13122 , n13137 );
nand ( n13139 , n12800 , n12779 );
nand ( n13140 , n13138 , n13139 );
not ( n13141 , n13140 );
buf ( n13142 , n12719 );
not ( n13143 , n13142 );
not ( n13144 , n12800 );
or ( n13145 , n13143 , n13144 );
buf ( n13146 , n12721 );
not ( n13147 , n13146 );
not ( n13148 , n12840 );
or ( n13149 , n13147 , n13148 );
or ( n13150 , n12840 , n13146 );
nand ( n13151 , n13149 , n13150 );
buf ( n13152 , n13151 );
nand ( n13153 , n13152 , n12886 );
nand ( n13154 , n13145 , n13153 );
not ( n13155 , n13154 );
nand ( n13156 , n13121 , n13141 , n13155 );
nor ( n13157 , n13106 , n13156 );
not ( n13158 , n12825 );
not ( n13159 , n12848 );
nand ( n13160 , n12840 , n12846 );
not ( n13161 , n13160 );
or ( n13162 , n13159 , n13161 );
nand ( n13163 , n12840 , n12846 );
or ( n13164 , n13163 , n12848 );
nand ( n13165 , n13162 , n13164 );
buf ( n13166 , n13165 );
not ( n13167 , n13166 );
not ( n13168 , n13167 );
not ( n13169 , n13168 );
or ( n13170 , n13158 , n13169 );
nand ( n13171 , n12800 , n12764 );
nand ( n13172 , n13170 , n13171 );
not ( n13173 , n13172 );
not ( n13174 , n12825 );
not ( n13175 , n12850 );
not ( n13176 , n13175 );
not ( n13177 , n12849 );
and ( n13178 , n12846 , n13177 );
nand ( n13179 , n12840 , n13178 );
not ( n13180 , n13179 );
or ( n13181 , n13176 , n13180 );
nand ( n13182 , n12840 , n13178 );
or ( n13183 , n13182 , n13175 );
nand ( n13184 , n13181 , n13183 );
buf ( n13185 , n13184 );
not ( n13186 , n13185 );
or ( n13187 , n13174 , n13186 );
nand ( n13188 , n12885 , n12775 );
nand ( n13189 , n13187 , n13188 );
not ( n13190 , n13189 );
not ( n13191 , n12800 );
not ( n13192 , n13191 );
not ( n13193 , n12847 );
and ( n13194 , n12846 , n12848 );
nand ( n13195 , n12840 , n13194 );
not ( n13196 , n13195 );
or ( n13197 , n13193 , n13196 );
nand ( n13198 , n12840 , n13194 );
or ( n13199 , n13198 , n12847 );
nand ( n13200 , n13197 , n13199 );
buf ( n13201 , n13200 );
not ( n13202 , n13201 );
or ( n13203 , n13192 , n13202 );
nand ( n13204 , n12800 , n12757 );
nand ( n13205 , n13203 , n13204 );
not ( n13206 , n13205 );
nand ( n13207 , n13173 , n13190 , n13206 );
not ( n13208 , n12825 );
nand ( n13209 , n12894 , n12906 );
nor ( n13210 , n12900 , n13209 );
not ( n13211 , n12962 );
nor ( n13212 , n13211 , n13072 );
nand ( n13213 , n12922 , n12987 );
nand ( n13214 , n12918 , n12994 );
nor ( n13215 , n13213 , n13214 );
nand ( n13216 , n12787 , n13210 , n13212 , n13215 );
buf ( n13217 , RI21a14f08_51);
buf ( n13218 , n13217 );
buf ( n13219 , n13218 );
not ( n13220 , n13219 );
xnor ( n13221 , n13216 , n13220 );
buf ( n13222 , n13221 );
not ( n13223 , n13222 );
or ( n13224 , n13208 , n13223 );
nand ( n13225 , n12800 , n13218 );
nand ( n13226 , n13224 , n13225 );
not ( n13227 , n13226 );
not ( n13228 , n13191 );
nor ( n13229 , n12898 , n12890 );
nor ( n13230 , n12789 , n13219 );
nand ( n13231 , n13229 , n13230 );
not ( n13232 , n13231 );
not ( n13233 , n12752 );
nand ( n13234 , n13233 , n12906 );
not ( n13235 , n12893 );
nand ( n13236 , n13235 , n12876 );
nor ( n13237 , n13234 , n13236 );
nand ( n13238 , n13232 , n13237 );
buf ( n13239 , RI21a14e90_52);
buf ( n13240 , n13239 );
buf ( n13241 , n13240 );
buf ( n13242 , n13241 );
nor ( n13243 , n13238 , n13242 );
nand ( n13244 , n12871 , n13243 );
buf ( n13245 , RI21a14e18_53);
buf ( n13246 , n13245 );
buf ( n13247 , n13246 );
not ( n13248 , n13247 );
xnor ( n13249 , n13244 , n13248 );
buf ( n13250 , n13249 );
not ( n13251 , n13250 );
or ( n13252 , n13228 , n13251 );
nand ( n13253 , n12885 , n13246 );
nand ( n13254 , n13252 , n13253 );
not ( n13255 , n13254 );
not ( n13256 , n12886 );
not ( n13257 , n12811 );
nor ( n13258 , n13247 , n13241 );
not ( n13259 , n13258 );
nand ( n13260 , n13237 , n13232 );
nor ( n13261 , n13259 , n13260 );
nand ( n13262 , n13257 , n13261 );
buf ( n13263 , RI21a14da0_54);
buf ( n13264 , n13263 );
buf ( n13265 , n13264 );
not ( n13266 , n13265 );
not ( n13267 , n13266 );
and ( n13268 , n13262 , n13267 );
not ( n13269 , n13262 );
and ( n13270 , n13269 , n13266 );
nor ( n13271 , n13268 , n13270 );
buf ( n13272 , n13271 );
not ( n13273 , n13272 );
not ( n13274 , n13273 );
not ( n13275 , n13274 );
or ( n13276 , n13256 , n13275 );
nand ( n13277 , n12800 , n13264 );
nand ( n13278 , n13276 , n13277 );
not ( n13279 , n13278 );
not ( n13280 , n12825 );
not ( n13281 , n13260 );
not ( n13282 , n13281 );
not ( n13283 , n12815 );
or ( n13284 , n13282 , n13283 );
not ( n13285 , n13242 );
nand ( n13286 , n13284 , n13285 );
not ( n13287 , n12731 );
not ( n13288 , n13241 );
nor ( n13289 , n13288 , n13124 );
nand ( n13290 , n13289 , n12739 , n12745 );
nor ( n13291 , n13290 , n12960 );
not ( n13292 , n13237 );
nor ( n13293 , n13292 , n12770 );
nand ( n13294 , n13287 , n13291 , n13293 , n13232 );
nand ( n13295 , n13286 , n13294 );
buf ( n13296 , n13295 );
not ( n13297 , n13296 );
or ( n13298 , n13280 , n13297 );
nand ( n13299 , n12800 , n13240 );
nand ( n13300 , n13298 , n13299 );
not ( n13301 , n13300 );
nand ( n13302 , n13227 , n13255 , n13279 , n13301 );
nor ( n13303 , n13207 , n13302 );
nand ( n13304 , n12985 , n13157 , n13303 );
not ( n13305 , n12812 );
not ( n13306 , n13281 );
buf ( n13307 , RI21a14d28_55);
buf ( n13308 , n13307 );
buf ( n13309 , n13308 );
nor ( n13310 , n13265 , n13309 );
nand ( n13311 , n13258 , n13310 );
not ( n13312 , n13311 );
buf ( n13313 , RI21a145a8_57);
buf ( n13314 , n13313 );
buf ( n13315 , n13314 );
not ( n13316 , n13315 );
buf ( n13317 , RI21a14cb0_56);
buf ( n13318 , n13317 );
buf ( n13319 , n13318 );
not ( n13320 , n13319 );
nand ( n13321 , n13316 , n13320 );
buf ( n13322 , RI21a144b8_59);
buf ( n13323 , n13322 );
buf ( n13324 , n13323 );
nor ( n13325 , n13321 , n13324 );
nand ( n13326 , n13312 , n13325 );
nor ( n13327 , n13306 , n13326 );
nand ( n13328 , n13305 , n13327 );
buf ( n13329 , n12705 );
buf ( n13330 , n13329 );
and ( n13331 , n13328 , n13330 );
not ( n13332 , n13328 );
not ( n13333 , n13330 );
and ( n13334 , n13332 , n13333 );
nor ( n13335 , n13331 , n13334 );
buf ( n13336 , n13335 );
nand ( n13337 , n13336 , n12801 );
not ( n13338 , n13337 );
buf ( n13339 , n13338 );
nand ( n13340 , n13304 , n13339 );
not ( n13341 , n13340 );
not ( n13342 , n13191 );
nand ( n13343 , n13258 , n13266 );
nor ( n13344 , n13260 , n13343 );
nand ( n13345 , n13257 , n13344 );
buf ( n13346 , n13309 );
and ( n13347 , n13345 , n13346 );
not ( n13348 , n13345 );
not ( n13349 , n13346 );
and ( n13350 , n13348 , n13349 );
nor ( n13351 , n13347 , n13350 );
buf ( n13352 , n13351 );
not ( n13353 , n13352 );
not ( n13354 , n13353 );
not ( n13355 , n13354 );
or ( n13356 , n13342 , n13355 );
nand ( n13357 , n12800 , n13308 );
nand ( n13358 , n13356 , n13357 );
and ( n13359 , n13341 , n13358 );
not ( n13360 , n13318 );
not ( n13361 , n12800 );
or ( n13362 , n13360 , n13361 );
nor ( n13363 , n13238 , n13311 );
nand ( n13364 , n12871 , n13363 );
xnor ( n13365 , n13364 , n13320 );
buf ( n13366 , n13365 );
buf ( n13367 , n13366 );
nand ( n13368 , n13367 , n13191 );
nand ( n13369 , n13362 , n13368 );
or ( n13370 , n13359 , n13369 );
nand ( n13371 , n13359 , n13369 );
nand ( n13372 , n13370 , n13371 );
not ( n13373 , n13372 );
buf ( n13374 , n13373 );
nand ( n13375 , n13312 , n13320 );
nor ( n13376 , n13306 , n13375 );
nand ( n13377 , n12816 , n13376 );
not ( n13378 , n13316 );
and ( n13379 , n13377 , n13378 );
not ( n13380 , n13377 );
and ( n13381 , n13380 , n13316 );
nor ( n13382 , n13379 , n13381 );
buf ( n13383 , n13382 );
not ( n13384 , n12800 );
and ( n13385 , n13383 , n13384 );
and ( n13386 , n12885 , n13314 );
nor ( n13387 , n13385 , n13386 );
not ( n13388 , n13387 );
not ( n13389 , n13388 );
nand ( n13390 , n12935 , n13032 );
not ( n13391 , n13390 );
nor ( n13392 , n13083 , n13098 );
nand ( n13393 , n13066 , n13048 , n13392 );
not ( n13394 , n13393 );
nand ( n13395 , n13391 , n13153 , n13394 , n13018 );
not ( n13396 , n13366 );
nor ( n13397 , n13222 , n13101 );
nand ( n13398 , n13396 , n13167 , n13353 , n13397 );
nor ( n13399 , n13395 , n13398 );
nor ( n13400 , n12859 , n13136 );
nand ( n13401 , n13400 , n12969 , n12798 );
nor ( n13402 , n13185 , n13201 );
nor ( n13403 , n13116 , n12943 );
nand ( n13404 , n13402 , n13403 );
nor ( n13405 , n13401 , n13404 );
nor ( n13406 , n13250 , n13296 );
nand ( n13407 , n12998 , n13406 , n13273 );
nor ( n13408 , n12978 , n12878 );
nor ( n13409 , n12908 , n12819 );
nand ( n13410 , n13408 , n13409 );
nor ( n13411 , n13407 , n13410 );
nand ( n13412 , n13399 , n13405 , n13411 );
nand ( n13413 , n13412 , n13338 );
not ( n13414 , n13413 );
or ( n13415 , n13389 , n13414 );
or ( n13416 , n13413 , n13388 );
nand ( n13417 , n13415 , n13416 );
not ( n13418 , n13417 );
buf ( n13419 , n13324 );
not ( n13420 , n13419 );
nor ( n13421 , n13311 , n13321 );
nand ( n13422 , n13281 , n13421 );
nor ( n13423 , n12812 , n13422 );
not ( n13424 , n13423 );
or ( n13425 , n13420 , n13424 );
nor ( n13426 , n12812 , n13422 );
or ( n13427 , n13426 , n13419 );
nand ( n13428 , n13425 , n13427 );
buf ( n13429 , n13428 );
and ( n13430 , n13429 , n13384 );
not ( n13431 , n13323 );
nor ( n13432 , n13431 , n13384 );
nor ( n13433 , n13430 , n13432 );
not ( n13434 , n13433 );
not ( n13435 , n13434 );
nor ( n13436 , n13387 , n13337 );
nand ( n13437 , n13412 , n13436 );
not ( n13438 , n13437 );
or ( n13439 , n13435 , n13438 );
nand ( n13440 , n13412 , n13436 , n13433 );
nand ( n13441 , n13439 , n13440 );
nand ( n13442 , n13418 , n13441 );
buf ( n13443 , n13442 );
not ( n13444 , n13443 );
buf ( n13445 , RI210d8710_180);
buf ( n13446 , n13445 );
nand ( n13447 , n13444 , n13446 );
nor ( n13448 , n13441 , n13418 );
not ( n13449 , n13448 );
not ( n13450 , n13449 );
buf ( n13451 , RI21a0b6b0_152);
buf ( n13452 , n13451 );
nand ( n13453 , n13450 , n13452 );
not ( n13454 , n13441 );
nor ( n13455 , n13454 , n13418 );
buf ( n13456 , n13455 );
buf ( n13457 , RI210d41b0_209);
buf ( n13458 , n13457 );
nand ( n13459 , n13456 , n13458 );
nor ( n13460 , n13417 , n13441 );
buf ( n13461 , n13460 );
buf ( n13462 , n13461 );
buf ( n13463 , RI21a0de10_124);
buf ( n13464 , n13463 );
nand ( n13465 , n13462 , n13464 );
nand ( n13466 , n13447 , n13453 , n13459 , n13465 );
buf ( n13467 , n13466 );
buf ( n13468 , n13467 );
not ( n13469 , n13443 );
buf ( n13470 , RI210d8788_179);
buf ( n13471 , n13470 );
nand ( n13472 , n13469 , n13471 );
buf ( n13473 , RI21a0b728_151);
buf ( n13474 , n13473 );
nand ( n13475 , n13450 , n13474 );
buf ( n13476 , RI210d4228_208);
buf ( n13477 , n13476 );
nand ( n13478 , n13456 , n13477 );
buf ( n13479 , RI21a0de88_123);
not ( n13480 , n13479 );
not ( n13481 , n13480 );
nand ( n13482 , n13462 , n13481 );
nand ( n13483 , n13472 , n13475 , n13478 , n13482 );
buf ( n13484 , n13483 );
buf ( n13485 , n13484 );
nand ( n13486 , n13468 , n13485 );
buf ( n13487 , n13486 );
buf ( n13488 , n13487 );
not ( n13489 , n13455 );
buf ( n13490 , RI210d37d8_213);
buf ( n13491 , n13490 );
not ( n13492 , n13491 );
nor ( n13493 , n13489 , n13492 );
buf ( n13494 , RI210d7d38_184);
buf ( n13495 , n13494 );
not ( n13496 , n13495 );
buf ( n13497 , n13443 );
nor ( n13498 , n13496 , n13497 );
nor ( n13499 , n13493 , n13498 );
buf ( n13500 , RI21a0ae40_156);
buf ( n13501 , n13500 );
not ( n13502 , n13501 );
nor ( n13503 , n13502 , n13449 );
not ( n13504 , n13461 );
buf ( n13505 , RI21a0dc30_128);
buf ( n13506 , n13505 );
not ( n13507 , n13506 );
nor ( n13508 , n13504 , n13507 );
nor ( n13509 , n13503 , n13508 );
nand ( n13510 , n13499 , n13509 );
buf ( n13511 , n13510 );
buf ( n13512 , n13511 );
nor ( n13513 , n13441 , n13418 );
not ( n13514 , n13513 );
not ( n13515 , n13514 );
buf ( n13516 , RI21a0aeb8_155);
buf ( n13517 , n13516 );
not ( n13518 , n13517 );
not ( n13519 , n13518 );
and ( n13520 , n13515 , n13519 );
buf ( n13521 , RI210d7db0_183);
buf ( n13522 , n13521 );
and ( n13523 , n13444 , n13522 );
nor ( n13524 , n13520 , n13523 );
buf ( n13525 , RI210d3850_212);
buf ( n13526 , n13525 );
not ( n13527 , n13526 );
nor ( n13528 , n13489 , n13527 );
buf ( n13529 , RI21a0dca8_127);
not ( n13530 , n13529 );
not ( n13531 , n13530 );
not ( n13532 , n13531 );
nor ( n13533 , n13504 , n13532 );
nor ( n13534 , n13528 , n13533 );
nand ( n13535 , n13524 , n13534 );
buf ( n13536 , n13535 );
buf ( n13537 , n13536 );
nand ( n13538 , n13512 , n13537 );
buf ( n13539 , n13538 );
buf ( n13540 , n13539 );
nor ( n13541 , n13488 , n13540 );
buf ( n13542 , n13541 );
buf ( n13543 , n13542 );
not ( n13544 , n13443 );
buf ( n13545 , RI210d5560_201);
buf ( n13546 , n13545 );
nand ( n13547 , n13544 , n13546 );
buf ( n13548 , RI210d9b38_171);
buf ( n13549 , n13548 );
nand ( n13550 , n13513 , n13549 );
nor ( n13551 , n13454 , n13418 );
not ( n13552 , n13551 );
not ( n13553 , n13552 );
buf ( n13554 , RI210d1078_229);
buf ( n13555 , n13554 );
nand ( n13556 , n13553 , n13555 );
nor ( n13557 , n13441 , n13417 );
not ( n13558 , n13557 );
not ( n13559 , n13558 );
buf ( n13560 , RI21a0c100_144);
not ( n13561 , n13560 );
not ( n13562 , n13561 );
nand ( n13563 , n13559 , n13562 );
nand ( n13564 , n13547 , n13550 , n13556 , n13563 );
buf ( n13565 , n13564 );
buf ( n13566 , n13565 );
buf ( n13567 , RI210d9160_175);
buf ( n13568 , n13567 );
nand ( n13569 , n13450 , n13568 );
buf ( n13570 , RI210d4b88_205);
buf ( n13571 , n13570 );
nand ( n13572 , n13469 , n13571 );
buf ( n13573 , RI210d06a0_233);
buf ( n13574 , n13573 );
nand ( n13575 , n13553 , n13574 );
buf ( n13576 , n13557 );
buf ( n13577 , RI21a0b908_147);
buf ( n13578 , n13577 );
nand ( n13579 , n13576 , n13578 );
nand ( n13580 , n13569 , n13572 , n13575 , n13579 );
buf ( n13581 , n13580 );
buf ( n13582 , n13581 );
not ( n13583 , n13443 );
buf ( n13584 , RI210d4c00_204);
buf ( n13585 , n13584 );
nand ( n13586 , n13583 , n13585 );
not ( n13587 , n13514 );
buf ( n13588 , RI210d99d0_174);
buf ( n13589 , n13588 );
nand ( n13590 , n13587 , n13589 );
not ( n13591 , n13552 );
buf ( n13592 , RI210d0718_232);
buf ( n13593 , n13592 );
nand ( n13594 , n13591 , n13593 );
buf ( n13595 , RI21a0c010_146);
buf ( n13596 , n13595 );
nand ( n13597 , n13559 , n13596 );
nand ( n13598 , n13586 , n13590 , n13594 , n13597 );
buf ( n13599 , n13598 );
buf ( n13600 , n13599 );
buf ( n13601 , n13456 );
buf ( n13602 , n13601 );
buf ( n13603 , n13602 );
nand ( n13604 , n13566 , n13582 , n13600 , n13603 );
buf ( n13605 , n13604 );
buf ( n13606 , n13605 );
not ( n13607 , n13606 );
buf ( n13608 , n13607 );
buf ( n13609 , n13608 );
buf ( n13610 , RI210d42a0_207);
buf ( n13611 , n13610 );
nand ( n13612 , n13583 , n13611 );
buf ( n13613 , RI210d9070_177);
buf ( n13614 , n13613 );
nand ( n13615 , n13587 , n13614 );
buf ( n13616 , RI210cfdb8_235);
buf ( n13617 , n13616 );
nand ( n13618 , n13591 , n13617 );
buf ( n13619 , RI21a0b818_149);
buf ( n13620 , n13619 );
nand ( n13621 , n13576 , n13620 );
nand ( n13622 , n13612 , n13615 , n13618 , n13621 );
buf ( n13623 , n13622 );
buf ( n13624 , n13623 );
buf ( n13625 , RI210d4b10_206);
buf ( n13626 , n13625 );
nand ( n13627 , n13544 , n13626 );
buf ( n13628 , RI210d90e8_176);
buf ( n13629 , n13628 );
nand ( n13630 , n13587 , n13629 );
buf ( n13631 , RI210d0628_234);
buf ( n13632 , n13631 );
nand ( n13633 , n13591 , n13632 );
buf ( n13634 , RI21a0b890_148);
buf ( n13635 , n13634 );
nand ( n13636 , n13576 , n13635 );
nand ( n13637 , n13627 , n13630 , n13633 , n13636 );
buf ( n13638 , n13637 );
buf ( n13639 , n13638 );
nand ( n13640 , n13624 , n13639 );
buf ( n13641 , n13640 );
buf ( n13642 , n13641 );
not ( n13643 , n13443 );
buf ( n13644 , RI210d54e8_202);
buf ( n13645 , n13644 );
nand ( n13646 , n13643 , n13645 );
not ( n13647 , n13514 );
buf ( n13648 , RI210d9ac0_172);
buf ( n13649 , n13648 );
nand ( n13650 , n13647 , n13649 );
not ( n13651 , n13552 );
buf ( n13652 , RI210d1000_230);
buf ( n13653 , n13652 );
nand ( n13654 , n13651 , n13653 );
not ( n13655 , n13558 );
buf ( n13656 , RI210cf2f0_241);
buf ( n13657 , n13656 );
nand ( n13658 , n13655 , n13657 );
nand ( n13659 , n13646 , n13650 , n13654 , n13658 );
buf ( n13660 , n13659 );
buf ( n13661 , n13660 );
not ( n13662 , n13661 );
buf ( n13663 , n13662 );
buf ( n13664 , n13663 );
nor ( n13665 , n13642 , n13664 );
buf ( n13666 , n13665 );
buf ( n13667 , n13666 );
not ( n13668 , n13443 );
buf ( n13669 , RI210d4c78_203);
buf ( n13670 , n13669 );
nand ( n13671 , n13668 , n13670 );
not ( n13672 , n13449 );
buf ( n13673 , RI210d9a48_173);
buf ( n13674 , n13673 );
nand ( n13675 , n13672 , n13674 );
buf ( n13676 , RI210d0790_231);
buf ( n13677 , n13676 );
nand ( n13678 , n13591 , n13677 );
not ( n13679 , n13558 );
buf ( n13680 , RI21a0c088_145);
not ( n13681 , n13680 );
not ( n13682 , n13681 );
nand ( n13683 , n13679 , n13682 );
nand ( n13684 , n13671 , n13675 , n13678 , n13683 );
buf ( n13685 , n13684 );
buf ( n13686 , n13685 );
not ( n13687 , n13514 );
buf ( n13688 , RI21a0af30_154);
buf ( n13689 , n13688 );
not ( n13690 , n13689 );
not ( n13691 , n13690 );
and ( n13692 , n13687 , n13691 );
not ( n13693 , n13443 );
buf ( n13694 , RI210d8620_182);
buf ( n13695 , n13694 );
and ( n13696 , n13693 , n13695 );
nor ( n13697 , n13692 , n13696 );
buf ( n13698 , RI210d38c8_211);
buf ( n13699 , n13698 );
not ( n13700 , n13699 );
nor ( n13701 , n13552 , n13700 );
not ( n13702 , n13576 );
buf ( n13703 , RI21a0dd20_126);
buf ( n13704 , n13703 );
not ( n13705 , n13704 );
nor ( n13706 , n13702 , n13705 );
nor ( n13707 , n13701 , n13706 );
nand ( n13708 , n13697 , n13707 );
buf ( n13709 , n13708 );
buf ( n13710 , n13709 );
nand ( n13711 , n13686 , n13710 );
buf ( n13712 , n13711 );
buf ( n13713 , n13712 );
buf ( n13714 , RI210d4138_210);
buf ( n13715 , n13714 );
nand ( n13716 , n13456 , n13715 );
buf ( n13717 , RI210d8698_181);
buf ( n13718 , n13717 );
nand ( n13719 , n13444 , n13718 );
buf ( n13720 , RI21a0dd98_125);
buf ( n13721 , n13720 );
nand ( n13722 , n13462 , n13721 );
buf ( n13723 , RI21a0afa8_153);
buf ( n13724 , n13723 );
nand ( n13725 , n13450 , n13724 );
nand ( n13726 , n13716 , n13719 , n13722 , n13725 );
buf ( n13727 , n13726 );
buf ( n13728 , n13727 );
not ( n13729 , n13728 );
buf ( n13730 , n13729 );
buf ( n13731 , n13730 );
nor ( n13732 , n13713 , n13731 );
buf ( n13733 , n13732 );
buf ( n13734 , n13733 );
and ( n13735 , n13543 , n13609 , n13667 , n13734 );
buf ( n13736 , n13735 );
buf ( n13737 , n13736 );
not ( n13738 , n13737 );
buf ( n13739 , n13738 );
buf ( n13740 , n13739 );
not ( n13741 , n13740 );
buf ( n13742 , n13741 );
buf ( n13743 , n13742 );
buf ( n13744 , n13743 );
buf ( n13745 , RI210d2ef0_215);
buf ( n13746 , n13745 );
not ( n13747 , n13746 );
nor ( n13748 , n13489 , n13747 );
buf ( n13749 , RI210cea08_243);
buf ( n13750 , n13749 );
not ( n13751 , n13750 );
buf ( n13752 , n13448 );
not ( n13753 , n13752 );
nor ( n13754 , n13751 , n13753 );
nor ( n13755 , n13748 , n13754 );
buf ( n13756 , RI210d7cc0_185);
buf ( n13757 , n13756 );
not ( n13758 , n13757 );
not ( n13759 , n13469 );
nor ( n13760 , n13758 , n13759 );
buf ( n13761 , RI210cfc50_238);
buf ( n13762 , n13761 );
not ( n13763 , n13762 );
nor ( n13764 , n13504 , n13763 );
nor ( n13765 , n13760 , n13764 );
nand ( n13766 , n13755 , n13765 );
buf ( n13767 , n13766 );
buf ( n13768 , n13767 );
buf ( n13769 , RI210d3760_214);
buf ( n13770 , n13769 );
not ( n13771 , n13770 );
nor ( n13772 , n13489 , n13771 );
buf ( n13773 , RI210cf278_242);
buf ( n13774 , n13773 );
not ( n13775 , n13774 );
nor ( n13776 , n13775 , n13753 );
nor ( n13777 , n13772 , n13776 );
buf ( n13778 , RI210ce8a0_246);
buf ( n13779 , n13778 );
not ( n13780 , n13779 );
nor ( n13781 , n13780 , n13759 );
buf ( n13782 , RI21a0d528_129);
buf ( n13783 , n13782 );
not ( n13784 , n13783 );
nor ( n13785 , n13504 , n13784 );
nor ( n13786 , n13781 , n13785 );
nand ( n13787 , n13777 , n13786 );
buf ( n13788 , n13787 );
buf ( n13789 , n13788 );
nand ( n13790 , n13768 , n13789 );
buf ( n13791 , n13790 );
buf ( n13792 , n13791 );
not ( n13793 , n13456 );
buf ( n13794 , RI210d23b0_222);
buf ( n13795 , n13794 );
not ( n13796 , n13795 );
nor ( n13797 , n13793 , n13796 );
buf ( n13798 , n13449 );
buf ( n13799 , RI21a0a558_161);
buf ( n13800 , n13799 );
not ( n13801 , n13800 );
nor ( n13802 , n13798 , n13801 );
nor ( n13803 , n13797 , n13802 );
not ( n13804 , n13497 );
buf ( n13805 , RI210d6a00_191);
buf ( n13806 , n13805 );
and ( n13807 , n13804 , n13806 );
buf ( n13808 , RI21a0d2d0_134);
buf ( n13809 , n13808 );
not ( n13810 , n13809 );
nor ( n13811 , n13504 , n13810 );
nor ( n13812 , n13807 , n13811 );
nand ( n13813 , n13803 , n13812 );
buf ( n13814 , n13813 );
buf ( n13815 , n13814 );
not ( n13816 , n13753 );
buf ( n13817 , RI21a0a648_159);
buf ( n13818 , n13817 );
not ( n13819 , n13818 );
not ( n13820 , n13819 );
and ( n13821 , n13816 , n13820 );
buf ( n13822 , RI210d72e8_189);
buf ( n13823 , n13822 );
and ( n13824 , n13804 , n13823 );
nor ( n13825 , n13821 , n13824 );
not ( n13826 , n13456 );
buf ( n13827 , RI210d24a0_220);
buf ( n13828 , n13827 );
not ( n13829 , n13828 );
nor ( n13830 , n13826 , n13829 );
buf ( n13831 , RI21a0d3c0_132);
buf ( n13832 , n13831 );
not ( n13833 , n13832 );
nor ( n13834 , n13504 , n13833 );
nor ( n13835 , n13830 , n13834 );
nand ( n13836 , n13825 , n13835 );
buf ( n13837 , n13836 );
buf ( n13838 , n13837 );
nand ( n13839 , n13815 , n13838 );
buf ( n13840 , n13839 );
buf ( n13841 , n13840 );
nor ( n13842 , n13792 , n13841 );
buf ( n13843 , n13842 );
buf ( n13844 , n13843 );
buf ( n13845 , RI210ce030_247);
buf ( n13846 , n13845 );
nand ( n13847 , n13804 , n13846 );
buf ( n13848 , RI21a0adc8_157);
buf ( n13849 , n13848 );
nand ( n13850 , n13752 , n13849 );
not ( n13851 , n13504 );
buf ( n13852 , RI21a0d4b0_130);
buf ( n13853 , n13852 );
nand ( n13854 , n13851 , n13853 );
buf ( n13855 , RI210d2e78_216);
buf ( n13856 , n13855 );
nand ( n13857 , n13456 , n13856 );
nand ( n13858 , n13847 , n13850 , n13854 , n13857 );
buf ( n13859 , n13858 );
buf ( n13860 , n13859 );
not ( n13861 , n13752 );
not ( n13862 , n13861 );
buf ( n13863 , RI21a0a5d0_160);
buf ( n13864 , n13863 );
not ( n13865 , n13864 );
not ( n13866 , n13865 );
and ( n13867 , n13862 , n13866 );
buf ( n13868 , RI210d7270_190);
not ( n13869 , n13868 );
not ( n13870 , n13869 );
and ( n13871 , n13804 , n13870 );
nor ( n13872 , n13867 , n13871 );
not ( n13873 , n13504 );
buf ( n13874 , RI21a0d348_133);
buf ( n13875 , n13874 );
not ( n13876 , n13875 );
not ( n13877 , n13876 );
and ( n13878 , n13873 , n13877 );
buf ( n13879 , RI210d2428_221);
buf ( n13880 , n13879 );
and ( n13881 , n13456 , n13880 );
nor ( n13882 , n13878 , n13881 );
nand ( n13883 , n13872 , n13882 );
buf ( n13884 , n13883 );
buf ( n13885 , n13884 );
not ( n13886 , n13861 );
buf ( n13887 , RI210ce990_244);
buf ( n13888 , n13887 );
not ( n13889 , n13888 );
not ( n13890 , n13889 );
and ( n13891 , n13886 , n13890 );
buf ( n13892 , RI210d7c48_186);
buf ( n13893 , n13892 );
and ( n13894 , n13804 , n13893 );
nor ( n13895 , n13891 , n13894 );
buf ( n13896 , RI210d2e00_217);
buf ( n13897 , n13896 );
not ( n13898 , n13897 );
nor ( n13899 , n13793 , n13898 );
not ( n13900 , n13462 );
buf ( n13901 , RI210cf3e0_239);
buf ( n13902 , n13901 );
not ( n13903 , n13902 );
nor ( n13904 , n13900 , n13903 );
nor ( n13905 , n13899 , n13904 );
nand ( n13906 , n13895 , n13905 );
buf ( n13907 , n13906 );
buf ( n13908 , n13907 );
buf ( n13909 , RI210d2518_219);
buf ( n13910 , n13909 );
not ( n13911 , n13910 );
nor ( n13912 , n13793 , n13911 );
buf ( n13913 , RI210ce918_245);
buf ( n13914 , n13913 );
not ( n13915 , n13914 );
nor ( n13916 , n13753 , n13915 );
nor ( n13917 , n13912 , n13916 );
not ( n13918 , n13693 );
buf ( n13919 , RI210d7360_188);
buf ( n13920 , n13919 );
not ( n13921 , n13920 );
nor ( n13922 , n13918 , n13921 );
buf ( n13923 , RI210cf368_240);
buf ( n13924 , n13923 );
not ( n13925 , n13924 );
nor ( n13926 , n13504 , n13925 );
nor ( n13927 , n13922 , n13926 );
nand ( n13928 , n13917 , n13927 );
buf ( n13929 , n13928 );
buf ( n13930 , n13929 );
and ( n13931 , n13860 , n13885 , n13908 , n13930 );
buf ( n13932 , n13931 );
buf ( n13933 , n13932 );
nand ( n13934 , n13844 , n13933 );
buf ( n13935 , n13934 );
buf ( n13936 , n13935 );
not ( n13937 , n13936 );
buf ( n13938 , n13937 );
buf ( n13939 , n13938 );
nand ( n13940 , n13744 , n13939 );
buf ( n13941 , n13940 );
buf ( n13942 , n13941 );
buf ( n13943 , RI21a09e50_162);
not ( n13944 , n13943 );
not ( n13945 , n13944 );
not ( n13946 , n13945 );
nor ( n13947 , n13753 , n13946 );
buf ( n13948 , RI210d1b40_223);
buf ( n13949 , n13948 );
not ( n13950 , n13949 );
nor ( n13951 , n13826 , n13950 );
nor ( n13952 , n13947 , n13951 );
buf ( n13953 , RI21a0cbc8_135);
not ( n13954 , n13953 );
not ( n13955 , n13954 );
and ( n13956 , n13462 , n13955 );
buf ( n13957 , RI210d6988_192);
not ( n13958 , n13957 );
not ( n13959 , n13958 );
not ( n13960 , n13959 );
nor ( n13961 , n13918 , n13960 );
nor ( n13962 , n13956 , n13961 );
nand ( n13963 , n13952 , n13962 );
buf ( n13964 , n13963 );
buf ( n13965 , n13964 );
buf ( n13966 , n13965 );
not ( n13967 , n13966 );
buf ( n13968 , n13967 );
buf ( n13969 , n13968 );
and ( n13970 , n13942 , n13969 );
not ( n13971 , n13942 );
buf ( n13972 , n13965 );
and ( n13973 , n13971 , n13972 );
nor ( n13974 , n13970 , n13973 );
buf ( n13975 , n13974 );
buf ( n13976 , n13975 );
and ( n13977 , n13374 , n13976 );
not ( n13978 , n13374 );
buf ( n13979 , n13743 );
buf ( n13980 , n13964 );
not ( n13981 , n13753 );
buf ( n13982 , RI21a09dd8_163);
not ( n13983 , n13982 );
not ( n13984 , n13983 );
not ( n13985 , n13984 );
not ( n13986 , n13985 );
and ( n13987 , n13981 , n13986 );
buf ( n13988 , RI210d6910_193);
not ( n13989 , n13988 );
not ( n13990 , n13989 );
and ( n13991 , n13804 , n13990 );
nor ( n13992 , n13987 , n13991 );
not ( n13993 , n13504 );
buf ( n13994 , RI21a0cb50_136);
not ( n13995 , n13994 );
not ( n13996 , n13995 );
not ( n13997 , n13996 );
not ( n13998 , n13997 );
and ( n13999 , n13993 , n13998 );
not ( n14000 , n13826 );
buf ( n14001 , RI210d1ac8_224);
buf ( n14002 , n14001 );
and ( n14003 , n14000 , n14002 );
nor ( n14004 , n13999 , n14003 );
nand ( n14005 , n13992 , n14004 );
buf ( n14006 , n14005 );
buf ( n14007 , n14006 );
and ( n14008 , n13980 , n14007 );
buf ( n14009 , n14008 );
buf ( n14010 , n14009 );
not ( n14011 , n14010 );
buf ( n14012 , n13938 );
not ( n14013 , n14012 );
buf ( n14014 , n14013 );
buf ( n14015 , n14014 );
nor ( n14016 , n14011 , n14015 );
buf ( n14017 , n14016 );
buf ( n14018 , n14017 );
nand ( n14019 , n13979 , n14018 );
buf ( n14020 , n14019 );
buf ( n14021 , n14020 );
not ( n14022 , n13861 );
buf ( n14023 , RI21a09478_164);
not ( n14024 , n14023 );
not ( n14025 , n14024 );
and ( n14026 , n14022 , n14025 );
buf ( n14027 , RI210d6898_194);
not ( n14028 , n14027 );
not ( n14029 , n14028 );
not ( n14030 , n14029 );
nor ( n14031 , n13918 , n14030 );
nor ( n14032 , n14026 , n14031 );
buf ( n14033 , RI210d1a50_225);
buf ( n14034 , n14033 );
and ( n14035 , n13456 , n14034 );
not ( n14036 , n13462 );
buf ( n14037 , RI21a0cad8_137);
not ( n14038 , n14037 );
not ( n14039 , n14038 );
not ( n14040 , n14039 );
nor ( n14041 , n14036 , n14040 );
nor ( n14042 , n14035 , n14041 );
nand ( n14043 , n14032 , n14042 );
buf ( n14044 , n14043 );
buf ( n14045 , n14044 );
buf ( n14046 , n14045 );
not ( n14047 , n14046 );
buf ( n14048 , n14047 );
buf ( n14049 , n14048 );
and ( n14050 , n14021 , n14049 );
not ( n14051 , n14021 );
buf ( n14052 , n14045 );
and ( n14053 , n14051 , n14052 );
nor ( n14054 , n14050 , n14053 );
buf ( n14055 , n14054 );
buf ( n14056 , n14055 );
buf ( n14057 , n14056 );
buf ( n14058 , n14057 );
not ( n14059 , n14058 );
not ( n14060 , n14059 );
buf ( n14061 , n13736 );
buf ( n14062 , n14061 );
buf ( n14063 , n13788 );
buf ( n14064 , n14063 );
nand ( n14065 , n14062 , n14064 );
buf ( n14066 , n14065 );
buf ( n14067 , n14066 );
buf ( n14068 , n13767 );
buf ( n14069 , n14068 );
not ( n14070 , n14069 );
buf ( n14071 , n14070 );
buf ( n14072 , n14071 );
and ( n14073 , n14067 , n14072 );
not ( n14074 , n14067 );
buf ( n14075 , n14068 );
and ( n14076 , n14074 , n14075 );
nor ( n14077 , n14073 , n14076 );
buf ( n14078 , n14077 );
buf ( n14079 , n14078 );
buf ( n14080 , n14079 );
buf ( n14081 , n13605 );
not ( n14082 , n14081 );
buf ( n14083 , n13685 );
buf ( n14084 , n14083 );
buf ( n14085 , n13660 );
nand ( n14086 , n14084 , n14085 );
buf ( n14087 , n14086 );
buf ( n14088 , n14087 );
not ( n14089 , n14088 );
buf ( n14090 , n14089 );
buf ( n14091 , n14090 );
nand ( n14092 , n14082 , n14091 );
buf ( n14093 , n14092 );
buf ( n14094 , n14093 );
not ( n14095 , n14094 );
buf ( n14096 , n14095 );
buf ( n14097 , n14096 );
buf ( n14098 , n13487 );
buf ( n14099 , n13641 );
nor ( n14100 , n14098 , n14099 );
buf ( n14101 , n14100 );
buf ( n14102 , n14101 );
not ( n14103 , n14102 );
buf ( n14104 , n13727 );
buf ( n14105 , n13709 );
and ( n14106 , n14104 , n14105 );
buf ( n14107 , n14106 );
buf ( n14108 , n14107 );
buf ( n14109 , n13536 );
buf ( n14110 , n14109 );
nand ( n14111 , n14108 , n14110 );
buf ( n14112 , n14111 );
buf ( n14113 , n14112 );
nor ( n14114 , n14103 , n14113 );
buf ( n14115 , n14114 );
buf ( n14116 , n14115 );
nand ( n14117 , n14097 , n14116 );
buf ( n14118 , n14117 );
buf ( n14119 , n14118 );
buf ( n14120 , n13511 );
buf ( n14121 , n14120 );
not ( n14122 , n14121 );
buf ( n14123 , n14122 );
buf ( n14124 , n14123 );
and ( n14125 , n14119 , n14124 );
not ( n14126 , n14119 );
buf ( n14127 , n14120 );
and ( n14128 , n14126 , n14127 );
nor ( n14129 , n14125 , n14128 );
buf ( n14130 , n14129 );
buf ( n14131 , n14130 );
buf ( n14132 , n14131 );
buf ( n14133 , n14096 );
buf ( n14134 , n14101 );
buf ( n14135 , n14107 );
and ( n14136 , n14134 , n14135 );
buf ( n14137 , n14136 );
buf ( n14138 , n14137 );
nand ( n14139 , n14133 , n14138 );
buf ( n14140 , n14139 );
buf ( n14141 , n14140 );
buf ( n14142 , n14109 );
buf ( n14143 , n14142 );
not ( n14144 , n14143 );
buf ( n14145 , n14144 );
buf ( n14146 , n14145 );
and ( n14147 , n14141 , n14146 );
not ( n14148 , n14141 );
buf ( n14149 , n14142 );
and ( n14150 , n14148 , n14149 );
nor ( n14151 , n14147 , n14150 );
buf ( n14152 , n14151 );
buf ( n14153 , n14152 );
buf ( n14154 , n14153 );
and ( n14155 , n14080 , n14132 , n14154 );
buf ( n14156 , n13739 );
not ( n14157 , n14156 );
buf ( n14158 , n14157 );
buf ( n14159 , n14158 );
buf ( n14160 , n13859 );
buf ( n14161 , n14160 );
not ( n14162 , n14161 );
buf ( n14163 , n13791 );
buf ( n14164 , n14163 );
buf ( n14165 , n14164 );
nor ( n14166 , n14162 , n14165 );
buf ( n14167 , n14166 );
buf ( n14168 , n14167 );
nand ( n14169 , n14159 , n14168 );
buf ( n14170 , n14169 );
buf ( n14171 , n14170 );
buf ( n14172 , n13907 );
buf ( n14173 , n14172 );
buf ( n14174 , n14173 );
not ( n14175 , n14174 );
buf ( n14176 , n14175 );
buf ( n14177 , n14176 );
and ( n14178 , n14171 , n14177 );
not ( n14179 , n14171 );
buf ( n14180 , n14173 );
and ( n14181 , n14179 , n14180 );
nor ( n14182 , n14178 , n14181 );
buf ( n14183 , n14182 );
buf ( n14184 , n14183 );
buf ( n14185 , n14184 );
buf ( n14186 , n14096 );
buf ( n14187 , n13641 );
buf ( n14188 , n14187 );
buf ( n14189 , n13484 );
buf ( n14190 , n14189 );
not ( n14191 , n14190 );
buf ( n14192 , n14191 );
buf ( n14193 , n14192 );
nor ( n14194 , n14188 , n14193 );
buf ( n14195 , n14194 );
buf ( n14196 , n14195 );
nand ( n14197 , n14186 , n14196 );
buf ( n14198 , n14197 );
buf ( n14199 , n14198 );
buf ( n14200 , n13467 );
buf ( n14201 , n14200 );
not ( n14202 , n14201 );
buf ( n14203 , n14202 );
buf ( n14204 , n14203 );
and ( n14205 , n14199 , n14204 );
not ( n14206 , n14199 );
buf ( n14207 , n14200 );
and ( n14208 , n14206 , n14207 );
nor ( n14209 , n14205 , n14208 );
buf ( n14210 , n14209 );
buf ( n14211 , n14210 );
buf ( n14212 , n14211 );
buf ( n14213 , n14212 );
nand ( n14214 , n14185 , n14213 );
not ( n14215 , n14214 );
buf ( n14216 , n13739 );
buf ( n14217 , n14063 );
not ( n14218 , n14217 );
buf ( n14219 , n14218 );
buf ( n14220 , n14219 );
and ( n14221 , n14216 , n14220 );
not ( n14222 , n14216 );
buf ( n14223 , n14063 );
and ( n14224 , n14222 , n14223 );
nor ( n14225 , n14221 , n14224 );
buf ( n14226 , n14225 );
buf ( n14227 , n14226 );
buf ( n14228 , n14227 );
buf ( n14229 , n14096 );
buf ( n14230 , n14101 );
buf ( n14231 , n13727 );
buf ( n14232 , n14231 );
and ( n14233 , n14230 , n14232 );
buf ( n14234 , n14233 );
buf ( n14235 , n14234 );
nand ( n14236 , n14229 , n14235 );
buf ( n14237 , n14236 );
buf ( n14238 , n14237 );
buf ( n14239 , n13709 );
buf ( n14240 , n14239 );
not ( n14241 , n14240 );
buf ( n14242 , n14241 );
buf ( n14243 , n14242 );
and ( n14244 , n14238 , n14243 );
not ( n14245 , n14238 );
buf ( n14246 , n14239 );
and ( n14247 , n14245 , n14246 );
nor ( n14248 , n14244 , n14247 );
buf ( n14249 , n14248 );
buf ( n14250 , n14249 );
buf ( n14251 , n14250 );
nand ( n14252 , n14228 , n14251 );
not ( n14253 , n14252 );
and ( n14254 , n14155 , n14215 , n14253 );
buf ( n14255 , n14093 );
not ( n14256 , n14255 );
buf ( n14257 , n14256 );
buf ( n14258 , n14257 );
buf ( n14259 , n13638 );
buf ( n14260 , n14259 );
nand ( n14261 , n14258 , n14260 );
buf ( n14262 , n14261 );
buf ( n14263 , n14262 );
buf ( n14264 , n13623 );
buf ( n14265 , n14264 );
not ( n14266 , n14265 );
buf ( n14267 , n14266 );
buf ( n14268 , n14267 );
and ( n14269 , n14263 , n14268 );
not ( n14270 , n14263 );
buf ( n14271 , n14264 );
and ( n14272 , n14270 , n14271 );
nor ( n14273 , n14269 , n14272 );
buf ( n14274 , n14273 );
buf ( n14275 , n14274 );
buf ( n14276 , n14275 );
buf ( n14277 , n14257 );
buf ( n14278 , n14101 );
nand ( n14279 , n14277 , n14278 );
buf ( n14280 , n14279 );
buf ( n14281 , n14280 );
buf ( n14282 , n14231 );
not ( n14283 , n14282 );
buf ( n14284 , n14283 );
buf ( n14285 , n14284 );
and ( n14286 , n14281 , n14285 );
not ( n14287 , n14281 );
buf ( n14288 , n14231 );
and ( n14289 , n14287 , n14288 );
nor ( n14290 , n14286 , n14289 );
buf ( n14291 , n14290 );
buf ( n14292 , n14291 );
buf ( n14293 , n14292 );
nand ( n14294 , n14276 , n14293 );
not ( n14295 , n14294 );
buf ( n14296 , n14061 );
buf ( n14297 , n14163 );
buf ( n14298 , n14172 );
buf ( n14299 , n14160 );
nand ( n14300 , n14298 , n14299 );
buf ( n14301 , n14300 );
buf ( n14302 , n14301 );
nor ( n14303 , n14297 , n14302 );
buf ( n14304 , n14303 );
buf ( n14305 , n14304 );
buf ( n14306 , n13884 );
buf ( n14307 , n14306 );
not ( n14308 , n14307 );
buf ( n14309 , n13837 );
buf ( n14310 , n14309 );
buf ( n14311 , n13929 );
buf ( n14312 , n14311 );
nand ( n14313 , n14310 , n14312 );
buf ( n14314 , n14313 );
buf ( n14315 , n14314 );
nor ( n14316 , n14308 , n14315 );
buf ( n14317 , n14316 );
buf ( n14318 , n14317 );
and ( n14319 , n14305 , n14318 );
buf ( n14320 , n14319 );
buf ( n14321 , n14320 );
nand ( n14322 , n14296 , n14321 );
buf ( n14323 , n14322 );
buf ( n14324 , n14323 );
buf ( n14325 , n13814 );
buf ( n14326 , n14325 );
not ( n14327 , n14326 );
buf ( n14328 , n14327 );
buf ( n14329 , n14328 );
and ( n14330 , n14324 , n14329 );
not ( n14331 , n14324 );
buf ( n14332 , n14325 );
and ( n14333 , n14331 , n14332 );
nor ( n14334 , n14330 , n14333 );
buf ( n14335 , n14334 );
buf ( n14336 , n14335 );
buf ( n14337 , n14336 );
buf ( n14338 , n14304 );
buf ( n14339 , n14311 );
buf ( n14340 , n14339 );
and ( n14341 , n14338 , n14340 );
buf ( n14342 , n14341 );
buf ( n14343 , n14342 );
buf ( n14344 , n14061 );
nand ( n14345 , n14343 , n14344 );
buf ( n14346 , n14345 );
buf ( n14347 , n14346 );
buf ( n14348 , n14309 );
buf ( n14349 , n14348 );
not ( n14350 , n14349 );
buf ( n14351 , n14350 );
buf ( n14352 , n14351 );
and ( n14353 , n14347 , n14352 );
not ( n14354 , n14347 );
buf ( n14355 , n14348 );
and ( n14356 , n14354 , n14355 );
nor ( n14357 , n14353 , n14356 );
buf ( n14358 , n14357 );
buf ( n14359 , n14358 );
buf ( n14360 , n14359 );
buf ( n14361 , n14061 );
buf ( n14362 , n14304 );
buf ( n14363 , n14314 );
not ( n14364 , n14363 );
buf ( n14365 , n14364 );
buf ( n14366 , n14365 );
and ( n14367 , n14362 , n14366 );
buf ( n14368 , n14367 );
buf ( n14369 , n14368 );
nand ( n14370 , n14361 , n14369 );
buf ( n14371 , n14370 );
buf ( n14372 , n14371 );
buf ( n14373 , n14306 );
not ( n14374 , n14373 );
buf ( n14375 , n14374 );
buf ( n14376 , n14375 );
and ( n14377 , n14372 , n14376 );
not ( n14378 , n14372 );
buf ( n14379 , n14306 );
and ( n14380 , n14378 , n14379 );
nor ( n14381 , n14377 , n14380 );
buf ( n14382 , n14381 );
buf ( n14383 , n14382 );
buf ( n14384 , n14383 );
nand ( n14385 , n14295 , n14337 , n14360 , n14384 );
buf ( n14386 , n13739 );
not ( n14387 , n14386 );
buf ( n14388 , n14387 );
buf ( n14389 , n14388 );
buf ( n14390 , n14304 );
nand ( n14391 , n14389 , n14390 );
buf ( n14392 , n14391 );
buf ( n14393 , n14392 );
buf ( n14394 , n14339 );
not ( n14395 , n14394 );
buf ( n14396 , n14395 );
buf ( n14397 , n14396 );
and ( n14398 , n14393 , n14397 );
not ( n14399 , n14393 );
buf ( n14400 , n14339 );
and ( n14401 , n14399 , n14400 );
nor ( n14402 , n14398 , n14401 );
buf ( n14403 , n14402 );
buf ( n14404 , n14403 );
buf ( n14405 , n14404 );
buf ( n14406 , n14388 );
buf ( n14407 , n14164 );
not ( n14408 , n14407 );
buf ( n14409 , n14408 );
buf ( n14410 , n14409 );
nand ( n14411 , n14406 , n14410 );
buf ( n14412 , n14411 );
buf ( n14413 , n14412 );
buf ( n14414 , n14160 );
buf ( n14415 , n14414 );
not ( n14416 , n14415 );
buf ( n14417 , n14416 );
buf ( n14418 , n14417 );
and ( n14419 , n14413 , n14418 );
not ( n14420 , n14413 );
buf ( n14421 , n14414 );
and ( n14422 , n14420 , n14421 );
nor ( n14423 , n14419 , n14422 );
buf ( n14424 , n14423 );
buf ( n14425 , n14424 );
buf ( n14426 , n14425 );
nand ( n14427 , n14405 , n14426 );
buf ( n14428 , n14083 );
buf ( n14429 , n13660 );
nand ( n14430 , n14428 , n14429 );
buf ( n14431 , n14430 );
buf ( n14432 , n14431 );
buf ( n14433 , n14187 );
nor ( n14434 , n14432 , n14433 );
buf ( n14435 , n14434 );
buf ( n14436 , n14435 );
buf ( n14437 , n13608 );
nand ( n14438 , n14436 , n14437 );
buf ( n14439 , n14438 );
buf ( n14440 , n14439 );
buf ( n14441 , n14192 );
and ( n14442 , n14440 , n14441 );
not ( n14443 , n14440 );
buf ( n14444 , n14189 );
and ( n14445 , n14443 , n14444 );
nor ( n14446 , n14442 , n14445 );
buf ( n14447 , n14446 );
buf ( n14448 , n14447 );
buf ( n14449 , n14448 );
not ( n14450 , n14449 );
buf ( n14451 , n14090 );
buf ( n14452 , n13599 );
buf ( n14453 , n14452 );
not ( n14454 , n14453 );
buf ( n14455 , n13565 );
not ( n14456 , n14455 );
buf ( n14457 , n14456 );
buf ( n14458 , n14457 );
nor ( n14459 , n14454 , n14458 );
buf ( n14460 , n14459 );
buf ( n14461 , n14460 );
buf ( n14462 , n13581 );
not ( n14463 , n14462 );
buf ( n14464 , n14463 );
buf ( n14465 , n14464 );
buf ( n14466 , n13602 );
not ( n14467 , n14466 );
buf ( n14468 , n14467 );
buf ( n14469 , n14468 );
nor ( n14470 , n14465 , n14469 );
buf ( n14471 , n14470 );
buf ( n14472 , n14471 );
nand ( n14473 , n14451 , n14461 , n14472 );
buf ( n14474 , n14473 );
buf ( n14475 , n14474 );
buf ( n14476 , n14259 );
not ( n14477 , n14476 );
buf ( n14478 , n14477 );
buf ( n14479 , n14478 );
and ( n14480 , n14475 , n14479 );
not ( n14481 , n14475 );
buf ( n14482 , n14259 );
and ( n14483 , n14481 , n14482 );
nor ( n14484 , n14480 , n14483 );
buf ( n14485 , n14484 );
buf ( n14486 , n14485 );
buf ( n14487 , n14486 );
buf ( n14488 , n14431 );
not ( n14489 , n14488 );
buf ( n14490 , n13565 );
buf ( n14491 , n13602 );
nand ( n14492 , n14490 , n14491 );
buf ( n14493 , n14492 );
buf ( n14494 , n14493 );
not ( n14495 , n14494 );
buf ( n14496 , n14495 );
buf ( n14497 , n14496 );
buf ( n14498 , n14452 );
buf ( n14499 , n14498 );
nand ( n14500 , n14489 , n14497 , n14499 );
buf ( n14501 , n14500 );
buf ( n14502 , n14501 );
buf ( n14503 , n14464 );
and ( n14504 , n14502 , n14503 );
not ( n14505 , n14502 );
buf ( n14506 , n14464 );
not ( n14507 , n14506 );
buf ( n14508 , n14507 );
buf ( n14509 , n14508 );
and ( n14510 , n14505 , n14509 );
nor ( n14511 , n14504 , n14510 );
buf ( n14512 , n14511 );
buf ( n14513 , n14512 );
buf ( n14514 , n14513 );
nand ( n14515 , n14487 , n14514 );
nor ( n14516 , n14450 , n14515 );
buf ( n14517 , n14493 );
buf ( n14518 , n14457 );
buf ( n14519 , n14468 );
nand ( n14520 , n14518 , n14519 );
buf ( n14521 , n14520 );
buf ( n14522 , n14521 );
and ( n14523 , n14517 , n14522 );
buf ( n14524 , n14523 );
buf ( n14525 , n14524 );
buf ( n14526 , n14525 );
buf ( n14527 , RI210d2d88_218);
buf ( n14528 , n14527 );
nand ( n14529 , n13601 , n14528 );
buf ( n14530 , RI21a0d438_131);
not ( n14531 , n14530 );
not ( n14532 , n14531 );
nand ( n14533 , n13462 , n14532 );
buf ( n14534 , RI21a0a6c0_158);
buf ( n14535 , n14534 );
nand ( n14536 , n14022 , n14535 );
not ( n14537 , n13918 );
buf ( n14538 , RI210d73d8_187);
buf ( n14539 , n14538 );
nand ( n14540 , n14537 , n14539 );
nand ( n14541 , n14529 , n14533 , n14536 , n14540 );
buf ( n14542 , n14541 );
buf ( n14543 , n14542 );
buf ( n14544 , RI210d10f0_228);
buf ( n14545 , n14544 );
not ( n14546 , n14545 );
not ( n14547 , n13601 );
or ( n14548 , n14546 , n14547 );
buf ( n14549 , RI210d5ec0_198);
buf ( n14550 , n14549 );
nand ( n14551 , n14537 , n14550 );
nand ( n14552 , n14548 , n14551 );
buf ( n14553 , RI210da498_168);
buf ( n14554 , n14553 );
not ( n14555 , n14554 );
not ( n14556 , n14022 );
or ( n14557 , n14555 , n14556 );
buf ( n14558 , RI21a0c268_141);
not ( n14559 , n14558 );
not ( n14560 , n14559 );
nand ( n14561 , n13462 , n14560 );
nand ( n14562 , n14557 , n14561 );
nor ( n14563 , n14552 , n14562 );
not ( n14564 , n14563 );
buf ( n14565 , n14564 );
and ( n14566 , n14543 , n14565 );
and ( n14567 , n14526 , n14566 );
buf ( n14568 , n14496 );
buf ( n14569 , n13660 );
buf ( n14570 , n14569 );
nand ( n14571 , n14568 , n14570 );
buf ( n14572 , n14571 );
buf ( n14573 , n14572 );
buf ( n14574 , n14083 );
not ( n14575 , n14574 );
buf ( n14576 , n14575 );
buf ( n14577 , n14576 );
xor ( n14578 , n14573 , n14577 );
buf ( n14579 , n14578 );
buf ( n14580 , n14579 );
buf ( n14581 , n14580 );
buf ( n14582 , n14431 );
not ( n14583 , n14582 );
buf ( n14584 , n14496 );
nand ( n14585 , n14583 , n14584 );
buf ( n14586 , n14585 );
buf ( n14587 , n14586 );
buf ( n14588 , n14498 );
buf ( n14589 , n14588 );
not ( n14590 , n14589 );
buf ( n14591 , n14590 );
buf ( n14592 , n14591 );
and ( n14593 , n14587 , n14592 );
not ( n14594 , n14587 );
buf ( n14595 , n14588 );
and ( n14596 , n14594 , n14595 );
nor ( n14597 , n14593 , n14596 );
buf ( n14598 , n14597 );
buf ( n14599 , n14598 );
buf ( n14600 , n14599 );
buf ( n14601 , n14569 );
not ( n14602 , n14601 );
buf ( n14603 , n14496 );
not ( n14604 , n14603 );
buf ( n14605 , n14604 );
buf ( n14606 , n14605 );
not ( n14607 , n14606 );
or ( n14608 , n14602 , n14607 );
buf ( n14609 , n14605 );
buf ( n14610 , n14569 );
or ( n14611 , n14609 , n14610 );
nand ( n14612 , n14608 , n14611 );
buf ( n14613 , n14612 );
buf ( n14614 , n14613 );
buf ( n14615 , n14614 );
and ( n14616 , n14567 , n14581 , n14600 , n14615 );
nand ( n14617 , n14516 , n14616 );
nor ( n14618 , n14385 , n14427 , n14617 );
buf ( n14619 , n13932 );
buf ( n14620 , n14009 );
buf ( n14621 , n13542 );
buf ( n14622 , n13666 );
nand ( n14623 , n14619 , n14620 , n14621 , n14622 );
buf ( n14624 , n14623 );
buf ( n14625 , n14624 );
not ( n14626 , n14625 );
buf ( n14627 , n13608 );
not ( n14628 , n13759 );
buf ( n14629 , RI210d5fb0_196);
not ( n14630 , n14629 );
not ( n14631 , n14630 );
and ( n14632 , n14628 , n14631 );
buf ( n14633 , RI210dad80_166);
not ( n14634 , n14633 );
not ( n14635 , n14634 );
not ( n14636 , n14635 );
nor ( n14637 , n13798 , n14636 );
nor ( n14638 , n14632 , n14637 );
buf ( n14639 , RI210d1168_227);
not ( n14640 , n14639 );
not ( n14641 , n14640 );
and ( n14642 , n14000 , n14641 );
buf ( n14643 , RI21a0c9e8_139);
not ( n14644 , n14643 );
not ( n14645 , n14644 );
not ( n14646 , n14645 );
nor ( n14647 , n13900 , n14646 );
nor ( n14648 , n14642 , n14647 );
nand ( n14649 , n14638 , n14648 );
buf ( n14650 , n14649 );
buf ( n14651 , n14650 );
buf ( n14652 , RI210d5f38_197);
not ( n14653 , n14652 );
not ( n14654 , n14653 );
nand ( n14655 , n13444 , n14654 );
buf ( n14656 , RI210da510_167);
not ( n14657 , n14656 );
not ( n14658 , n14657 );
nand ( n14659 , n14022 , n14658 );
buf ( n14660 , RI21a0c970_140);
not ( n14661 , n14660 );
not ( n14662 , n14661 );
nand ( n14663 , n13462 , n14662 );
nand ( n14664 , n14655 , n14659 , n14663 );
buf ( n14665 , n14664 );
buf ( n14666 , n14665 );
nand ( n14667 , n14651 , n14666 );
buf ( n14668 , n14667 );
buf ( n14669 , n14668 );
buf ( n14670 , RI210da420_169);
not ( n14671 , n14670 );
not ( n14672 , n14671 );
nand ( n14673 , n14022 , n14672 );
buf ( n14674 , RI210d5650_199);
not ( n14675 , n14674 );
not ( n14676 , n14675 );
nand ( n14677 , n13444 , n14676 );
not ( n14678 , n13504 );
buf ( n14679 , RI21a0c1f0_142);
not ( n14680 , n14679 );
not ( n14681 , n14680 );
nand ( n14682 , n14678 , n14681 );
nand ( n14683 , n14673 , n14677 , n14682 );
buf ( n14684 , n14683 );
buf ( n14685 , n14684 );
not ( n14686 , n14685 );
buf ( n14687 , n14686 );
buf ( n14688 , n14687 );
nor ( n14689 , n14669 , n14688 );
buf ( n14690 , n14689 );
buf ( n14691 , n14690 );
buf ( n14692 , n14107 );
nand ( n14693 , n14627 , n14691 , n14692 );
buf ( n14694 , n14693 );
buf ( n14695 , n14694 );
buf ( n14696 , n14044 );
not ( n14697 , n13444 );
buf ( n14698 , RI210d6028_195);
not ( n14699 , n14698 );
not ( n14700 , n14699 );
not ( n14701 , n14700 );
nor ( n14702 , n14697 , n14701 );
buf ( n14703 , RI210dadf8_165);
not ( n14704 , n14703 );
not ( n14705 , n14704 );
not ( n14706 , n14705 );
nor ( n14707 , n13861 , n14706 );
nor ( n14708 , n14702 , n14707 );
buf ( n14709 , RI21a0ca60_138);
not ( n14710 , n14709 );
not ( n14711 , n14710 );
and ( n14712 , n14678 , n14711 );
buf ( n14713 , RI210d19d8_226);
buf ( n14714 , n14713 );
not ( n14715 , n14714 );
nor ( n14716 , n13793 , n14715 );
nor ( n14717 , n14712 , n14716 );
nand ( n14718 , n14708 , n14717 );
buf ( n14719 , n14718 );
buf ( n14720 , n14719 );
nand ( n14721 , n14696 , n14720 );
buf ( n14722 , n14721 );
buf ( n14723 , n14722 );
buf ( n14724 , n14576 );
nor ( n14725 , n14723 , n14724 );
buf ( n14726 , n14725 );
buf ( n14727 , n14726 );
buf ( n14728 , n13843 );
nand ( n14729 , n14727 , n14728 );
buf ( n14730 , n14729 );
buf ( n14731 , n14730 );
nor ( n14732 , n14695 , n14731 );
buf ( n14733 , n14732 );
buf ( n14734 , n14733 );
nand ( n14735 , n14626 , n14734 );
buf ( n14736 , n14735 );
buf ( n14737 , n14736 );
buf ( n14738 , RI210da3a8_170);
buf ( n14739 , n14738 );
nand ( n14740 , n14022 , n14739 );
buf ( n14741 , RI210d55d8_200);
buf ( n14742 , n14741 );
nand ( n14743 , n14628 , n14742 );
buf ( n14744 , RI21a0c178_143);
buf ( n14745 , n14744 );
nand ( n14746 , n14678 , n14745 );
nand ( n14747 , n14740 , n14743 , n14746 );
buf ( n14748 , n14747 );
buf ( n14749 , n14748 );
not ( n14750 , n14749 );
buf ( n14751 , n14750 );
buf ( n14752 , n14751 );
and ( n14753 , n14737 , n14752 );
not ( n14754 , n14737 );
buf ( n14755 , n14748 );
and ( n14756 , n14754 , n14755 );
nor ( n14757 , n14753 , n14756 );
buf ( n14758 , n14757 );
buf ( n14759 , n14758 );
buf ( n14760 , RI210cdfb8_248);
buf ( n14761 , n14760 );
nand ( n14762 , n13601 , n14761 );
buf ( n14763 , n13462 );
buf ( n14764 , RI21a0e590_122);
not ( n14765 , n14764 );
not ( n14766 , n14765 );
nand ( n14767 , n14763 , n14766 );
buf ( n14768 , n14022 );
buf ( n14769 , RI21a0b7a0_150);
buf ( n14770 , n14769 );
nand ( n14771 , n14768 , n14770 );
buf ( n14772 , RI210d8ff8_178);
buf ( n14773 , n14772 );
nand ( n14774 , n14537 , n14773 );
nand ( n14775 , n14762 , n14767 , n14771 , n14774 );
and ( n14776 , n14759 , n14775 );
buf ( n14777 , n14776 );
buf ( n14778 , n14777 );
nand ( n14779 , n14254 , n14618 , n14778 );
buf ( n14780 , n13976 );
not ( n14781 , n14780 );
nor ( n14782 , n14779 , n14781 );
buf ( n14783 , n13743 );
buf ( n14784 , n14014 );
buf ( n14785 , n13968 );
nor ( n14786 , n14784 , n14785 );
buf ( n14787 , n14786 );
buf ( n14788 , n14787 );
nand ( n14789 , n14783 , n14788 );
buf ( n14790 , n14789 );
buf ( n14791 , n14790 );
buf ( n14792 , n14006 );
xnor ( n14793 , n14791 , n14792 );
buf ( n14794 , n14793 );
buf ( n14795 , n14794 );
buf ( n14796 , n14795 );
buf ( n14797 , n14796 );
nand ( n14798 , n14782 , n14797 );
not ( n14799 , n14798 );
not ( n14800 , n14799 );
or ( n14801 , n14060 , n14800 );
or ( n14802 , n14799 , n14059 );
nand ( n14803 , n14801 , n14802 );
buf ( n14804 , n14803 );
and ( n14805 , n13978 , n14804 );
nor ( n14806 , n13977 , n14805 );
buf ( n14807 , n13254 );
buf ( n14808 , n13226 );
not ( n14809 , n14808 );
not ( n14810 , n13339 );
or ( n14811 , n14809 , n14810 );
not ( n14812 , n13207 );
nand ( n14813 , n12985 , n13157 , n14812 );
nand ( n14814 , n14813 , n13339 );
nand ( n14815 , n14811 , n14814 );
not ( n14816 , n14815 );
nor ( n14817 , n14816 , n13301 );
and ( n14818 , n14807 , n14817 );
not ( n14819 , n13279 );
and ( n14820 , n14818 , n14819 );
not ( n14821 , n14818 );
and ( n14822 , n14821 , n13279 );
nor ( n14823 , n14820 , n14822 );
xor ( n14824 , n14807 , n14817 );
xnor ( n14825 , n14815 , n13301 );
and ( n14826 , n14824 , n14825 );
nand ( n14827 , n14823 , n14826 );
buf ( n14828 , RI210cfd40_236);
buf ( n14829 , n14828 );
buf ( n14830 , n14829 );
and ( n14831 , n14827 , n14830 );
buf ( n14832 , n14814 );
not ( n14833 , n14832 );
not ( n14834 , n14808 );
and ( n14835 , n14833 , n14834 );
and ( n14836 , n14832 , n14808 );
nor ( n14837 , n14835 , n14836 );
not ( n14838 , n14837 );
not ( n14839 , n14838 );
and ( n14840 , n14831 , n14839 );
not ( n14841 , n14840 );
not ( n14842 , n14841 );
buf ( n14843 , n14823 );
not ( n14844 , n14843 );
nand ( n14845 , n14844 , n14824 );
buf ( n14846 , RI21a16a38_35);
buf ( n14847 , n14846 );
not ( n14848 , n14847 );
not ( n14849 , n14825 );
or ( n14850 , n14848 , n14849 );
or ( n14851 , n14825 , n14847 );
nand ( n14852 , n14850 , n14851 );
nor ( n14853 , n14852 , n14824 );
nand ( n14854 , n14843 , n14853 );
buf ( n14855 , RI21a115d8_89);
buf ( n14856 , n14855 );
nand ( n14857 , n14843 , n14856 );
nand ( n14858 , n14845 , n14854 , n14857 );
nand ( n14859 , n14842 , n14858 );
not ( n14860 , n14859 );
buf ( n14861 , RI21a11650_88);
buf ( n14862 , n14861 );
and ( n14863 , n14843 , n14862 );
not ( n14864 , n14825 );
nor ( n14865 , n14843 , n14864 );
nor ( n14866 , n14863 , n14865 );
nand ( n14867 , n14866 , n14854 );
not ( n14868 , n14867 );
nand ( n14869 , n14860 , n14868 );
not ( n14870 , n14869 );
nor ( n14871 , n13156 , n12936 );
not ( n14872 , n12884 );
and ( n14873 , n13069 , n13105 );
and ( n14874 , n14871 , n14872 , n14873 );
not ( n14875 , n14812 );
nor ( n14876 , n14875 , n13003 );
and ( n14877 , n14874 , n14876 );
not ( n14878 , n13339 );
nor ( n14879 , n14877 , n14878 );
buf ( n14880 , n12982 );
nand ( n14881 , n14879 , n14880 );
buf ( n14882 , n12970 );
not ( n14883 , n14882 );
nor ( n14884 , n14881 , n14883 );
buf ( n14885 , n12947 );
xnor ( n14886 , n14884 , n14885 );
not ( n14887 , n14886 );
nand ( n14888 , n14884 , n14885 );
buf ( n14889 , n12912 );
not ( n14890 , n14889 );
and ( n14891 , n14888 , n14890 );
not ( n14892 , n14888 );
and ( n14893 , n14892 , n14889 );
nor ( n14894 , n14891 , n14893 );
nand ( n14895 , n14887 , n14894 );
not ( n14896 , n14895 );
and ( n14897 , n14881 , n14882 );
not ( n14898 , n14881 );
and ( n14899 , n14898 , n14883 );
nor ( n14900 , n14897 , n14899 );
and ( n14901 , n14879 , n14880 );
not ( n14902 , n14879 );
not ( n14903 , n14880 );
and ( n14904 , n14902 , n14903 );
or ( n14905 , n14901 , n14904 );
and ( n14906 , n14900 , n14905 );
and ( n14907 , n14896 , n14906 );
nand ( n14908 , n14870 , n14907 );
buf ( n14909 , n14908 );
or ( n14910 , n14806 , n14909 );
not ( n14911 , n13340 );
not ( n14912 , n13358 );
and ( n14913 , n14911 , n14912 );
and ( n14914 , n13340 , n13358 );
nor ( n14915 , n14913 , n14914 );
xnor ( n14916 , n13358 , n13369 );
nand ( n14917 , n14915 , n14916 );
buf ( n14918 , n14917 );
not ( n14919 , n14918 );
not ( n14920 , n14919 );
not ( n14921 , n277910 );
buf ( n14922 , n9761 );
buf ( n14923 , n14922 );
buf ( n14924 , n277646 );
buf ( n14925 , n14924 );
or ( n14926 , n14923 , n14925 );
buf ( n14927 , n14926 );
buf ( n14928 , n14927 );
buf ( n14929 , n14922 );
buf ( n14930 , n14924 );
nand ( n14931 , n14929 , n14930 );
buf ( n14932 , n14931 );
buf ( n14933 , n14932 );
nand ( n14934 , n14928 , n14933 );
buf ( n14935 , n14934 );
buf ( n14936 , n14935 );
not ( n14937 , n14936 );
buf ( n14938 , n9706 );
buf ( n14939 , n14938 );
buf ( n14940 , n278001 );
buf ( n14941 , n14940 );
nor ( n14942 , n14939 , n14941 );
buf ( n14943 , n14942 );
buf ( n14944 , n14943 );
buf ( n14945 , n9714 );
buf ( n14946 , n14945 );
buf ( n14947 , n277926 );
buf ( n14948 , n14947 );
nor ( n14949 , n14946 , n14948 );
buf ( n14950 , n14949 );
buf ( n14951 , n14950 );
nor ( n14952 , n14944 , n14951 );
buf ( n14953 , n14952 );
buf ( n14954 , n14953 );
buf ( n14955 , n9732 );
buf ( n14956 , n14955 );
buf ( n14957 , n10642 );
buf ( n14958 , n14957 );
nor ( n14959 , n14956 , n14958 );
buf ( n14960 , n14959 );
buf ( n14961 , n14960 );
buf ( n14962 , n9724 );
buf ( n14963 , n14962 );
buf ( n14964 , n278049 );
buf ( n14965 , n14964 );
nor ( n14966 , n14963 , n14965 );
buf ( n14967 , n14966 );
buf ( n14968 , n14967 );
nor ( n14969 , n14961 , n14968 );
buf ( n14970 , n14969 );
buf ( n14971 , n14970 );
and ( n14972 , n14954 , n14971 );
buf ( n14973 , n14972 );
buf ( n14974 , n14973 );
buf ( n14975 , n9671 );
buf ( n14976 , n14975 );
buf ( n14977 , n277891 );
buf ( n14978 , n14977 );
nor ( n14979 , n14976 , n14978 );
buf ( n14980 , n14979 );
buf ( n14981 , n14980 );
buf ( n14982 , n9679 );
buf ( n14983 , n14982 );
buf ( n14984 , n277818 );
buf ( n14985 , n14984 );
nor ( n14986 , n14983 , n14985 );
buf ( n14987 , n14986 );
buf ( n14988 , n14987 );
nor ( n14989 , n14981 , n14988 );
buf ( n14990 , n14989 );
buf ( n14991 , n14990 );
buf ( n14992 , n9696 );
buf ( n14993 , n14992 );
buf ( n14994 , n277794 );
buf ( n14995 , n14994 );
nor ( n14996 , n14993 , n14995 );
buf ( n14997 , n14996 );
buf ( n14998 , n14997 );
buf ( n14999 , n9688 );
buf ( n15000 , n14999 );
buf ( n15001 , n277745 );
buf ( n15002 , n15001 );
nor ( n15003 , n15000 , n15002 );
buf ( n15004 , n15003 );
buf ( n15005 , n15004 );
nor ( n15006 , n14998 , n15005 );
buf ( n15007 , n15006 );
buf ( n15008 , n15007 );
and ( n15009 , n14991 , n15008 );
buf ( n15010 , n15009 );
buf ( n15011 , n15010 );
and ( n15012 , n14974 , n15011 );
buf ( n15013 , n15012 );
buf ( n15014 , n15013 );
buf ( n15015 , n277692 );
buf ( n15016 , n15015 );
buf ( n15017 , n9769 );
buf ( n15018 , n15017 );
or ( n15019 , n15016 , n15018 );
buf ( n15020 , n15019 );
buf ( n15021 , n15020 );
and ( n15022 , n15014 , n15021 );
buf ( n15023 , n15022 );
buf ( n15024 , n15023 );
not ( n15025 , n15024 );
buf ( n15026 , n9552 );
buf ( n15027 , n15026 );
buf ( n15028 , n10830 );
buf ( n15029 , n15028 );
or ( n15030 , n15027 , n15029 );
buf ( n15031 , n15030 );
buf ( n15032 , n15031 );
buf ( n15033 , n10735 );
buf ( n15034 , n15033 );
not ( n15035 , n15034 );
buf ( n15036 , n9587 );
not ( n15037 , n15036 );
buf ( n15038 , n15037 );
buf ( n15039 , n15038 );
nand ( n15040 , n15035 , n15039 );
buf ( n15041 , n15040 );
buf ( n15042 , n15041 );
and ( n15043 , n15032 , n15042 );
buf ( n15044 , n15043 );
buf ( n15045 , n15044 );
not ( n15046 , n15045 );
buf ( n15047 , n9509 );
buf ( n15048 , n15047 );
buf ( n15049 , n11672 );
buf ( n15050 , n15049 );
or ( n15051 , n15048 , n15050 );
buf ( n15052 , n15051 );
buf ( n15053 , n15052 );
buf ( n15054 , n9517 );
buf ( n15055 , n15054 );
buf ( n15056 , n11592 );
buf ( n15057 , n15056 );
or ( n15058 , n15055 , n15057 );
buf ( n15059 , n15058 );
buf ( n15060 , n15059 );
and ( n15061 , n15053 , n15060 );
buf ( n15062 , n15061 );
buf ( n15063 , n15062 );
not ( n15064 , n15063 );
or ( n15065 , n15046 , n15064 );
buf ( n15066 , n15054 );
buf ( n15067 , n15056 );
and ( n15068 , n15066 , n15067 );
buf ( n15069 , n15068 );
buf ( n15070 , n15069 );
not ( n15071 , n15070 );
buf ( n15072 , n15052 );
not ( n15073 , n15072 );
or ( n15074 , n15071 , n15073 );
buf ( n15075 , n15047 );
buf ( n15076 , n15049 );
nand ( n15077 , n15075 , n15076 );
buf ( n15078 , n15077 );
buf ( n15079 , n15078 );
nand ( n15080 , n15074 , n15079 );
buf ( n15081 , n15080 );
buf ( n15082 , n15081 );
not ( n15083 , n15082 );
buf ( n15084 , n15083 );
buf ( n15085 , n15084 );
nand ( n15086 , n15065 , n15085 );
buf ( n15087 , n15086 );
buf ( n15088 , n15087 );
buf ( n15089 , n9527 );
buf ( n15090 , n15089 );
buf ( n15091 , n11329 );
buf ( n15092 , n15091 );
or ( n15093 , n15090 , n15092 );
buf ( n15094 , n15093 );
buf ( n15095 , n15094 );
buf ( n15096 , n9562 );
buf ( n15097 , n15096 );
buf ( n15098 , n11236 );
buf ( n15099 , n15098 );
or ( n15100 , n15097 , n15099 );
buf ( n15101 , n15100 );
buf ( n15102 , n15101 );
nand ( n15103 , n15095 , n15102 );
buf ( n15104 , n15103 );
buf ( n15105 , n15104 );
not ( n15106 , n15105 );
buf ( n15107 , n9535 );
buf ( n15108 , n15107 );
buf ( n15109 , n11512 );
buf ( n15110 , n15109 );
nor ( n15111 , n15108 , n15110 );
buf ( n15112 , n15111 );
buf ( n15113 , n15112 );
buf ( n15114 , n9570 );
buf ( n15115 , n15114 );
buf ( n15116 , n11568 );
buf ( n15117 , n15116 );
nor ( n15118 , n15115 , n15117 );
buf ( n15119 , n15118 );
buf ( n15120 , n15119 );
nor ( n15121 , n15113 , n15120 );
buf ( n15122 , n15121 );
buf ( n15123 , n15122 );
nand ( n15124 , n15106 , n15123 );
buf ( n15125 , n15124 );
buf ( n15126 , n15125 );
buf ( n15127 , n9544 );
buf ( n15128 , n15127 );
buf ( n15129 , n11452 );
buf ( n15130 , n15129 );
or ( n15131 , n15128 , n15130 );
buf ( n15132 , n15131 );
buf ( n15133 , n15132 );
buf ( n15134 , n9579 );
buf ( n15135 , n15134 );
buf ( n15136 , n11364 );
buf ( n15137 , n15136 );
or ( n15138 , n15135 , n15137 );
buf ( n15139 , n15138 );
buf ( n15140 , n15139 );
nand ( n15141 , n15133 , n15140 );
buf ( n15142 , n15141 );
buf ( n15143 , n15142 );
nor ( n15144 , n15126 , n15143 );
buf ( n15145 , n15144 );
buf ( n15146 , n15145 );
buf ( n15147 , n9500 );
buf ( n15148 , n15147 );
buf ( n15149 , n10956 );
buf ( n15150 , n15149 );
or ( n15151 , n15148 , n15150 );
buf ( n15152 , n15151 );
buf ( n15153 , n15152 );
buf ( n15154 , n9492 );
buf ( n15155 , n15154 );
buf ( n15156 , n10846 );
buf ( n15157 , n15156 );
or ( n15158 , n15155 , n15157 );
buf ( n15159 , n15158 );
buf ( n15160 , n15159 );
nand ( n15161 , n15153 , n15160 );
buf ( n15162 , n15161 );
buf ( n15163 , n15162 );
not ( n15164 , n15163 );
buf ( n15165 , n15164 );
buf ( n15166 , n15165 );
not ( n15167 , n15166 );
buf ( n15168 , n9462 );
buf ( n15169 , n15168 );
buf ( n15170 , n11103 );
buf ( n15171 , n15170 );
or ( n15172 , n15169 , n15171 );
buf ( n15173 , n15172 );
buf ( n15174 , n15173 );
not ( n15175 , n15174 );
buf ( n15176 , n9470 );
buf ( n15177 , n15176 );
buf ( n15178 , n11147 );
buf ( n15179 , n15178 );
and ( n15180 , n15177 , n15179 );
buf ( n15181 , n15180 );
buf ( n15182 , n15181 );
not ( n15183 , n15182 );
or ( n15184 , n15175 , n15183 );
buf ( n15185 , n15168 );
buf ( n15186 , n15170 );
nand ( n15187 , n15185 , n15186 );
buf ( n15188 , n15187 );
buf ( n15189 , n15188 );
nand ( n15190 , n15184 , n15189 );
buf ( n15191 , n15190 );
buf ( n15192 , n15191 );
not ( n15193 , n15192 );
or ( n15194 , n15167 , n15193 );
buf ( n15195 , n15084 );
nand ( n15196 , n15194 , n15195 );
buf ( n15197 , n15196 );
buf ( n15198 , n15197 );
nand ( n15199 , n15088 , n15146 , n15198 );
buf ( n15200 , n15199 );
buf ( n15201 , n15200 );
buf ( n15202 , n15125 );
not ( n15203 , n15202 );
buf ( n15204 , n9449 );
buf ( n15205 , n15204 );
buf ( n15206 , n10971 );
buf ( n15207 , n15206 );
or ( n15208 , n15205 , n15207 );
buf ( n15209 , n15208 );
buf ( n15210 , n15209 );
not ( n15211 , n15210 );
buf ( n15212 , n9440 );
buf ( n15213 , n15212 );
buf ( n15214 , n11050 );
buf ( n15215 , n15214 );
and ( n15216 , n15213 , n15215 );
buf ( n15217 , n15216 );
buf ( n15218 , n15217 );
not ( n15219 , n15218 );
or ( n15220 , n15211 , n15219 );
buf ( n15221 , n15204 );
buf ( n15222 , n15206 );
nand ( n15223 , n15221 , n15222 );
buf ( n15224 , n15223 );
buf ( n15225 , n15224 );
nand ( n15226 , n15220 , n15225 );
buf ( n15227 , n15226 );
buf ( n15228 , n15227 );
buf ( n15229 , n15176 );
buf ( n15230 , n15178 );
nor ( n15231 , n15229 , n15230 );
buf ( n15232 , n15231 );
buf ( n15233 , n15232 );
buf ( n15234 , n15168 );
buf ( n15235 , n15170 );
nor ( n15236 , n15234 , n15235 );
buf ( n15237 , n15236 );
buf ( n15238 , n15237 );
nor ( n15239 , n15233 , n15238 );
buf ( n15240 , n15239 );
buf ( n15241 , n15240 );
and ( n15242 , n15228 , n15241 );
buf ( n15243 , n15242 );
buf ( n15244 , n15243 );
buf ( n15245 , n15062 );
buf ( n15246 , n15044 );
and ( n15247 , n15245 , n15246 );
buf ( n15248 , n15247 );
buf ( n15249 , n15248 );
buf ( n15250 , n15142 );
buf ( n15251 , n15162 );
nor ( n15252 , n15250 , n15251 );
buf ( n15253 , n15252 );
buf ( n15254 , n15253 );
nand ( n15255 , n15203 , n15244 , n15249 , n15254 );
buf ( n15256 , n15255 );
buf ( n15257 , n15256 );
buf ( n15258 , n15127 );
buf ( n15259 , n15129 );
nand ( n15260 , n15258 , n15259 );
buf ( n15261 , n15260 );
buf ( n15262 , n15261 );
buf ( n15263 , n15089 );
buf ( n15264 , n15091 );
nand ( n15265 , n15263 , n15264 );
buf ( n15266 , n15265 );
buf ( n15267 , n15266 );
nand ( n15268 , n15262 , n15267 );
buf ( n15269 , n15268 );
buf ( n15270 , n15269 );
buf ( n15271 , n15096 );
buf ( n15272 , n15098 );
and ( n15273 , n15271 , n15272 );
buf ( n15274 , n15273 );
buf ( n15275 , n15274 );
nor ( n15276 , n15270 , n15275 );
buf ( n15277 , n15276 );
buf ( n15278 , n15277 );
not ( n15279 , n15278 );
buf ( n15280 , n15132 );
buf ( n15281 , n15134 );
buf ( n15282 , n15136 );
and ( n15283 , n15281 , n15282 );
buf ( n15284 , n15283 );
buf ( n15285 , n15284 );
nand ( n15286 , n15280 , n15285 );
buf ( n15287 , n15286 );
buf ( n15288 , n15287 );
not ( n15289 , n15288 );
or ( n15290 , n15279 , n15289 );
buf ( n15291 , n15104 );
buf ( n15292 , n15266 );
nand ( n15293 , n15291 , n15292 );
buf ( n15294 , n15293 );
buf ( n15295 , n15294 );
nand ( n15296 , n15290 , n15295 );
buf ( n15297 , n15296 );
buf ( n15298 , n15297 );
buf ( n15299 , n15132 );
buf ( n15300 , n15094 );
buf ( n15301 , n15139 );
buf ( n15302 , n15101 );
and ( n15303 , n15299 , n15300 , n15301 , n15302 );
buf ( n15304 , n15303 );
buf ( n15305 , n15304 );
buf ( n15306 , n15112 );
not ( n15307 , n15306 );
buf ( n15308 , n15307 );
buf ( n15309 , n15308 );
not ( n15310 , n15309 );
buf ( n15311 , n15114 );
buf ( n15312 , n15116 );
and ( n15313 , n15311 , n15312 );
buf ( n15314 , n15313 );
buf ( n15315 , n15314 );
not ( n15316 , n15315 );
or ( n15317 , n15310 , n15316 );
buf ( n15318 , n15107 );
buf ( n15319 , n15109 );
nand ( n15320 , n15318 , n15319 );
buf ( n15321 , n15320 );
buf ( n15322 , n15321 );
nand ( n15323 , n15317 , n15322 );
buf ( n15324 , n15323 );
buf ( n15325 , n15324 );
nand ( n15326 , n15305 , n15325 );
buf ( n15327 , n15326 );
buf ( n15328 , n15327 );
and ( n15329 , n15298 , n15328 );
buf ( n15330 , n15329 );
buf ( n15331 , n15330 );
buf ( n15332 , n15304 );
not ( n15333 , n15332 );
buf ( n15334 , n15333 );
buf ( n15335 , n15334 );
not ( n15336 , n15335 );
buf ( n15337 , n15062 );
buf ( n15338 , n15122 );
and ( n15339 , n15337 , n15338 );
buf ( n15340 , n15339 );
buf ( n15341 , n15340 );
buf ( n15342 , n15044 );
not ( n15343 , n15342 );
buf ( n15344 , n15152 );
not ( n15345 , n15344 );
buf ( n15346 , n15154 );
buf ( n15347 , n15156 );
and ( n15348 , n15346 , n15347 );
buf ( n15349 , n15348 );
buf ( n15350 , n15349 );
not ( n15351 , n15350 );
or ( n15352 , n15345 , n15351 );
buf ( n15353 , n15147 );
buf ( n15354 , n15149 );
nand ( n15355 , n15353 , n15354 );
buf ( n15356 , n15355 );
buf ( n15357 , n15356 );
nand ( n15358 , n15352 , n15357 );
buf ( n15359 , n15358 );
buf ( n15360 , n15359 );
not ( n15361 , n15360 );
or ( n15362 , n15343 , n15361 );
buf ( n15363 , n15031 );
buf ( n15364 , n15033 );
not ( n15365 , n15364 );
buf ( n15366 , n15038 );
nor ( n15367 , n15365 , n15366 );
buf ( n15368 , n15367 );
buf ( n15369 , n15368 );
and ( n15370 , n15363 , n15369 );
buf ( n15371 , n15026 );
buf ( n15372 , n15028 );
and ( n15373 , n15371 , n15372 );
buf ( n15374 , n15373 );
buf ( n15375 , n15374 );
nor ( n15376 , n15370 , n15375 );
buf ( n15377 , n15376 );
buf ( n15378 , n15377 );
nand ( n15379 , n15362 , n15378 );
buf ( n15380 , n15379 );
buf ( n15381 , n15380 );
nand ( n15382 , n15336 , n15341 , n15381 );
buf ( n15383 , n15382 );
buf ( n15384 , n15383 );
nand ( n15385 , n15201 , n15257 , n15331 , n15384 );
buf ( n15386 , n15385 );
buf ( n15387 , n15386 );
buf ( n15388 , n15387 );
not ( n15389 , n15388 );
or ( n15390 , n15025 , n15389 );
buf ( n15391 , n15010 );
not ( n15392 , n15391 );
buf ( n15393 , n14955 );
buf ( n15394 , n14957 );
and ( n15395 , n15393 , n15394 );
buf ( n15396 , n15395 );
buf ( n15397 , n15396 );
buf ( n15398 , n14967 );
not ( n15399 , n15398 );
buf ( n15400 , n15399 );
buf ( n15401 , n15400 );
nand ( n15402 , n15397 , n15401 );
buf ( n15403 , n15402 );
buf ( n15404 , n15403 );
buf ( n15405 , n14962 );
buf ( n15406 , n14964 );
nand ( n15407 , n15405 , n15406 );
buf ( n15408 , n15407 );
buf ( n15409 , n15408 );
nand ( n15410 , n15404 , n15409 );
buf ( n15411 , n15410 );
buf ( n15412 , n15411 );
not ( n15413 , n15412 );
buf ( n15414 , n14953 );
not ( n15415 , n15414 );
or ( n15416 , n15413 , n15415 );
buf ( n15417 , n14943 );
not ( n15418 , n15417 );
buf ( n15419 , n15418 );
buf ( n15420 , n15419 );
buf ( n15421 , n14945 );
buf ( n15422 , n14947 );
and ( n15423 , n15421 , n15422 );
buf ( n15424 , n15423 );
buf ( n15425 , n15424 );
and ( n15426 , n15420 , n15425 );
buf ( n15427 , n14938 );
buf ( n15428 , n14940 );
and ( n15429 , n15427 , n15428 );
buf ( n15430 , n15429 );
buf ( n15431 , n15430 );
nor ( n15432 , n15426 , n15431 );
buf ( n15433 , n15432 );
buf ( n15434 , n15433 );
nand ( n15435 , n15416 , n15434 );
buf ( n15436 , n15435 );
buf ( n15437 , n15436 );
not ( n15438 , n15437 );
or ( n15439 , n15392 , n15438 );
buf ( n15440 , n14982 );
buf ( n15441 , n14984 );
and ( n15442 , n15440 , n15441 );
buf ( n15443 , n15442 );
buf ( n15444 , n15443 );
not ( n15445 , n15444 );
buf ( n15446 , n14980 );
not ( n15447 , n15446 );
buf ( n15448 , n15447 );
buf ( n15449 , n15448 );
not ( n15450 , n15449 );
or ( n15451 , n15445 , n15450 );
buf ( n15452 , n14975 );
buf ( n15453 , n14977 );
nand ( n15454 , n15452 , n15453 );
buf ( n15455 , n15454 );
buf ( n15456 , n15455 );
nand ( n15457 , n15451 , n15456 );
buf ( n15458 , n15457 );
buf ( n15459 , n15458 );
buf ( n15460 , n15007 );
and ( n15461 , n15459 , n15460 );
buf ( n15462 , n14992 );
buf ( n15463 , n14994 );
nand ( n15464 , n15462 , n15463 );
buf ( n15465 , n15464 );
buf ( n15466 , n15465 );
buf ( n15467 , n15004 );
or ( n15468 , n15466 , n15467 );
buf ( n15469 , n14999 );
buf ( n15470 , n15001 );
nand ( n15471 , n15469 , n15470 );
buf ( n15472 , n15471 );
buf ( n15473 , n15472 );
nand ( n15474 , n15468 , n15473 );
buf ( n15475 , n15474 );
buf ( n15476 , n15475 );
nor ( n15477 , n15461 , n15476 );
buf ( n15478 , n15477 );
buf ( n15479 , n15478 );
nand ( n15480 , n15439 , n15479 );
buf ( n15481 , n15480 );
buf ( n15482 , n15481 );
buf ( n15483 , n15020 );
and ( n15484 , n15482 , n15483 );
buf ( n15485 , n15017 );
buf ( n15486 , n15015 );
and ( n15487 , n15485 , n15486 );
buf ( n15488 , n15487 );
buf ( n15489 , n15488 );
nor ( n15490 , n15484 , n15489 );
buf ( n15491 , n15490 );
buf ( n15492 , n15491 );
nand ( n15493 , n15390 , n15492 );
buf ( n15494 , n15493 );
buf ( n15495 , n15494 );
not ( n15496 , n15495 );
or ( n15497 , n14937 , n15496 );
buf ( n15498 , n15494 );
buf ( n15499 , n14935 );
or ( n15500 , n15498 , n15499 );
nand ( n15501 , n15497 , n15500 );
buf ( n15502 , n15501 );
buf ( n15503 , n15502 );
not ( n15504 , n15503 );
or ( n15505 , n14921 , n15504 );
nand ( n15506 , n277603 , n9761 );
nand ( n15507 , n15505 , n15506 );
nand ( n15508 , n14920 , n15507 );
not ( n15509 , n15508 );
buf ( n15510 , n15509 );
not ( n15511 , n15510 );
buf ( n15512 , n14005 );
buf ( n15513 , n15512 );
buf ( n15514 , n15513 );
not ( n15515 , n15514 );
or ( n15516 , n15511 , n15515 );
not ( n15517 , n15514 );
not ( n15518 , n15510 );
nand ( n15519 , n15517 , n15518 );
nand ( n15520 , n15516 , n15519 );
not ( n15521 , n14917 );
not ( n15522 , n15521 );
buf ( n15523 , n15522 );
not ( n15524 , n277910 );
buf ( n15525 , n15488 );
not ( n15526 , n15525 );
buf ( n15527 , n15020 );
nand ( n15528 , n15526 , n15527 );
buf ( n15529 , n15528 );
buf ( n15530 , n15529 );
not ( n15531 , n15530 );
buf ( n15532 , n15013 );
not ( n15533 , n15532 );
buf ( n15534 , n15387 );
not ( n15535 , n15534 );
or ( n15536 , n15533 , n15535 );
buf ( n15537 , n15481 );
not ( n15538 , n15537 );
buf ( n15539 , n15538 );
buf ( n15540 , n15539 );
nand ( n15541 , n15536 , n15540 );
buf ( n15542 , n15541 );
buf ( n15543 , n15542 );
not ( n15544 , n15543 );
or ( n15545 , n15531 , n15544 );
buf ( n15546 , n15542 );
buf ( n15547 , n15529 );
or ( n15548 , n15546 , n15547 );
nand ( n15549 , n15545 , n15548 );
buf ( n15550 , n15549 );
buf ( n15551 , n15550 );
not ( n15552 , n15551 );
or ( n15553 , n15524 , n15552 );
nand ( n15554 , n277527 , n9769 );
nand ( n15555 , n15553 , n15554 );
and ( n15556 , n15523 , n15555 );
buf ( n15557 , n15556 );
buf ( n15558 , n15557 );
not ( n15559 , n15558 );
buf ( n15560 , n13963 );
buf ( n15561 , n15560 );
buf ( n15562 , n15561 );
and ( n15563 , n15559 , n15562 );
nor ( n15564 , n15520 , n15563 );
not ( n15565 , n15564 );
nand ( n15566 , n15520 , n15563 );
nand ( n15567 , n15565 , n15566 );
not ( n15568 , n15567 );
buf ( n15569 , n13858 );
buf ( n15570 , n15569 );
not ( n15571 , n15570 );
buf ( n15572 , n14917 );
not ( n15573 , n15572 );
not ( n15574 , n12883 );
and ( n15575 , n15573 , n15574 );
not ( n15576 , n9431 );
buf ( n15577 , n15424 );
not ( n15578 , n15577 );
buf ( n15579 , n14950 );
not ( n15580 , n15579 );
buf ( n15581 , n15580 );
buf ( n15582 , n15581 );
nand ( n15583 , n15578 , n15582 );
buf ( n15584 , n15583 );
buf ( n15585 , n15584 );
not ( n15586 , n15585 );
buf ( n15587 , n14970 );
not ( n15588 , n15587 );
buf ( n15589 , n15386 );
not ( n15590 , n15589 );
or ( n15591 , n15588 , n15590 );
buf ( n15592 , n15411 );
not ( n15593 , n15592 );
buf ( n15594 , n15593 );
buf ( n15595 , n15594 );
nand ( n15596 , n15591 , n15595 );
buf ( n15597 , n15596 );
buf ( n15598 , n15597 );
not ( n15599 , n15598 );
or ( n15600 , n15586 , n15599 );
buf ( n15601 , n15597 );
buf ( n15602 , n15584 );
or ( n15603 , n15601 , n15602 );
nand ( n15604 , n15600 , n15603 );
buf ( n15605 , n15604 );
buf ( n15606 , n15605 );
not ( n15607 , n15606 );
or ( n15608 , n15576 , n15607 );
nand ( n15609 , n277352 , n9714 );
nand ( n15610 , n15608 , n15609 );
and ( n15611 , n15523 , n15610 );
nor ( n15612 , n15575 , n15611 );
not ( n15613 , n15612 );
buf ( n15614 , n15613 );
not ( n15615 , n15614 );
or ( n15616 , n15571 , n15615 );
not ( n15617 , n15570 );
not ( n15618 , n15614 );
nand ( n15619 , n15617 , n15618 );
nand ( n15620 , n15616 , n15619 );
buf ( n15621 , n13766 );
buf ( n15622 , n15621 );
not ( n15623 , n15622 );
not ( n15624 , n15521 );
not ( n15625 , n15624 );
not ( n15626 , n12799 );
not ( n15627 , n15626 );
and ( n15628 , n15625 , n15627 );
buf ( n15629 , n14918 );
not ( n15630 , n277983 );
buf ( n15631 , n15081 );
buf ( n15632 , n15122 );
and ( n15633 , n15631 , n15632 );
buf ( n15634 , n15324 );
nor ( n15635 , n15633 , n15634 );
buf ( n15636 , n15635 );
buf ( n15637 , n15636 );
buf ( n15638 , n15181 );
not ( n15639 , n15638 );
buf ( n15640 , n15639 );
buf ( n15641 , n15640 );
buf ( n15642 , n15188 );
and ( n15643 , n15641 , n15642 );
buf ( n15644 , n15643 );
buf ( n15645 , n15644 );
not ( n15646 , n15645 );
buf ( n15647 , n15227 );
buf ( n15648 , n15232 );
not ( n15649 , n15648 );
buf ( n15650 , n15649 );
buf ( n15651 , n15650 );
nand ( n15652 , n15647 , n15651 );
buf ( n15653 , n15652 );
buf ( n15654 , n15653 );
not ( n15655 , n15654 );
or ( n15656 , n15646 , n15655 );
buf ( n15657 , n15165 );
buf ( n15658 , n15044 );
buf ( n15659 , n15188 );
buf ( n15660 , n15237 );
nand ( n15661 , n15659 , n15660 );
buf ( n15662 , n15661 );
buf ( n15663 , n15662 );
and ( n15664 , n15657 , n15658 , n15663 );
buf ( n15665 , n15664 );
buf ( n15666 , n15665 );
nand ( n15667 , n15656 , n15666 );
buf ( n15668 , n15667 );
buf ( n15669 , n15668 );
buf ( n15670 , n15297 );
not ( n15671 , n15670 );
buf ( n15672 , n15671 );
buf ( n15673 , n15672 );
buf ( n15674 , n15380 );
nor ( n15675 , n15673 , n15674 );
buf ( n15676 , n15675 );
buf ( n15677 , n15676 );
nand ( n15678 , n15637 , n15669 , n15677 );
buf ( n15679 , n15678 );
buf ( n15680 , n15679 );
buf ( n15681 , n15636 );
buf ( n15682 , n15672 );
buf ( n15683 , n15340 );
nor ( n15684 , n15682 , n15683 );
buf ( n15685 , n15684 );
buf ( n15686 , n15685 );
nand ( n15687 , n15681 , n15686 );
buf ( n15688 , n15687 );
buf ( n15689 , n15688 );
buf ( n15690 , n15297 );
buf ( n15691 , n15334 );
and ( n15692 , n15690 , n15691 );
buf ( n15693 , n14960 );
nor ( n15694 , n15692 , n15693 );
buf ( n15695 , n15694 );
buf ( n15696 , n15695 );
nand ( n15697 , n15680 , n15689 , n15696 );
buf ( n15698 , n15697 );
buf ( n15699 , n15698 );
buf ( n15700 , n15396 );
not ( n15701 , n15700 );
buf ( n15702 , n15701 );
buf ( n15703 , n15702 );
nand ( n15704 , n15699 , n15703 );
buf ( n15705 , n15704 );
buf ( n15706 , n15705 );
buf ( n15707 , n15400 );
buf ( n15708 , n15408 );
nand ( n15709 , n15707 , n15708 );
buf ( n15710 , n15709 );
buf ( n15711 , n15710 );
not ( n15712 , n15711 );
buf ( n15713 , n15712 );
buf ( n15714 , n15713 );
and ( n15715 , n15706 , n15714 );
not ( n15716 , n15706 );
buf ( n15717 , n15710 );
and ( n15718 , n15716 , n15717 );
nor ( n15719 , n15715 , n15718 );
buf ( n15720 , n15719 );
buf ( n15721 , n15720 );
not ( n15722 , n15721 );
or ( n15723 , n15630 , n15722 );
nand ( n15724 , n9432 , n9724 );
nand ( n15725 , n15723 , n15724 );
and ( n15726 , n15629 , n15725 );
nor ( n15727 , n15628 , n15726 );
not ( n15728 , n15727 );
buf ( n15729 , n15728 );
nor ( n15730 , n15623 , n15729 );
nor ( n15731 , n15620 , n15730 );
not ( n15732 , n15731 );
buf ( n15733 , n13906 );
buf ( n15734 , n15733 );
not ( n15735 , n15734 );
not ( n15736 , n15572 );
not ( n15737 , n12983 );
and ( n15738 , n15736 , n15737 );
not ( n15739 , n277910 );
buf ( n15740 , n15430 );
not ( n15741 , n15740 );
buf ( n15742 , n15419 );
nand ( n15743 , n15741 , n15742 );
buf ( n15744 , n15743 );
buf ( n15745 , n15744 );
not ( n15746 , n15745 );
buf ( n15747 , n14970 );
buf ( n15748 , n15581 );
and ( n15749 , n15747 , n15748 );
buf ( n15750 , n15749 );
buf ( n15751 , n15750 );
not ( n15752 , n15751 );
buf ( n15753 , n15386 );
not ( n15754 , n15753 );
or ( n15755 , n15752 , n15754 );
buf ( n15756 , n15411 );
buf ( n15757 , n15581 );
and ( n15758 , n15756 , n15757 );
buf ( n15759 , n15424 );
nor ( n15760 , n15758 , n15759 );
buf ( n15761 , n15760 );
buf ( n15762 , n15761 );
nand ( n15763 , n15755 , n15762 );
buf ( n15764 , n15763 );
buf ( n15765 , n15764 );
not ( n15766 , n15765 );
or ( n15767 , n15746 , n15766 );
buf ( n15768 , n15764 );
buf ( n15769 , n15744 );
or ( n15770 , n15768 , n15769 );
nand ( n15771 , n15767 , n15770 );
buf ( n15772 , n15771 );
buf ( n15773 , n15772 );
not ( n15774 , n15773 );
or ( n15775 , n15739 , n15774 );
nand ( n15776 , n277352 , n9706 );
nand ( n15777 , n15775 , n15776 );
and ( n15778 , n14920 , n15777 );
nor ( n15779 , n15738 , n15778 );
not ( n15780 , n15779 );
buf ( n15781 , n15780 );
not ( n15782 , n15781 );
or ( n15783 , n15735 , n15782 );
not ( n15784 , n15734 );
not ( n15785 , n15781 );
nand ( n15786 , n15784 , n15785 );
nand ( n15787 , n15783 , n15786 );
not ( n15788 , n15787 );
and ( n15789 , n15618 , n15570 );
not ( n15790 , n15789 );
nand ( n15791 , n15788 , n15790 );
nand ( n15792 , n15732 , n15791 );
not ( n15793 , n15792 );
not ( n15794 , n15622 );
not ( n15795 , n15729 );
or ( n15796 , n15794 , n15795 );
not ( n15797 , n15729 );
nand ( n15798 , n15797 , n15623 );
nand ( n15799 , n15796 , n15798 );
buf ( n15800 , n13787 );
buf ( n15801 , n15800 );
not ( n15802 , n15801 );
not ( n15803 , n12823 );
not ( n15804 , n14919 );
or ( n15805 , n15803 , n15804 );
not ( n15806 , n277351 );
buf ( n15807 , n14960 );
not ( n15808 , n15807 );
buf ( n15809 , n15702 );
nand ( n15810 , n15808 , n15809 );
buf ( n15811 , n15810 );
buf ( n15812 , n15811 );
not ( n15813 , n15812 );
buf ( n15814 , n15387 );
not ( n15815 , n15814 );
or ( n15816 , n15813 , n15815 );
buf ( n15817 , n15387 );
buf ( n15818 , n15811 );
or ( n15819 , n15817 , n15818 );
nand ( n15820 , n15816 , n15819 );
buf ( n15821 , n15820 );
buf ( n15822 , n15821 );
not ( n15823 , n15822 );
or ( n15824 , n15806 , n15823 );
nand ( n15825 , n277603 , n9732 );
nand ( n15826 , n15824 , n15825 );
nand ( n15827 , n15572 , n15826 );
nand ( n15828 , n15805 , n15827 );
buf ( n15829 , n15828 );
nor ( n15830 , n15802 , n15829 );
or ( n15831 , n15799 , n15830 );
not ( n15832 , n15801 );
not ( n15833 , n15829 );
or ( n15834 , n15832 , n15833 );
not ( n15835 , n15829 );
nand ( n15836 , n15835 , n15802 );
nand ( n15837 , n15834 , n15836 );
buf ( n15838 , n13510 );
buf ( n15839 , n15838 );
buf ( n15840 , n15839 );
not ( n15841 , n15840 );
or ( n15842 , n15572 , n12864 );
not ( n15843 , n9431 );
buf ( n15844 , n15101 );
not ( n15845 , n15844 );
buf ( n15846 , n15142 );
nor ( n15847 , n15845 , n15846 );
buf ( n15848 , n15847 );
buf ( n15849 , n15848 );
buf ( n15850 , n15340 );
and ( n15851 , n15849 , n15850 );
buf ( n15852 , n15851 );
buf ( n15853 , n15852 );
not ( n15854 , n15853 );
buf ( n15855 , n15380 );
not ( n15856 , n15855 );
buf ( n15857 , n15668 );
nand ( n15858 , n15856 , n15857 );
buf ( n15859 , n15858 );
buf ( n15860 , n15859 );
not ( n15861 , n15860 );
or ( n15862 , n15854 , n15861 );
buf ( n15863 , n15636 );
not ( n15864 , n15863 );
buf ( n15865 , n15864 );
buf ( n15866 , n15865 );
buf ( n15867 , n15848 );
and ( n15868 , n15866 , n15867 );
buf ( n15869 , n15101 );
not ( n15870 , n15869 );
buf ( n15871 , n15287 );
buf ( n15872 , n15261 );
nand ( n15873 , n15871 , n15872 );
buf ( n15874 , n15873 );
buf ( n15875 , n15874 );
not ( n15876 , n15875 );
or ( n15877 , n15870 , n15876 );
buf ( n15878 , n15274 );
not ( n15879 , n15878 );
buf ( n15880 , n15879 );
buf ( n15881 , n15880 );
nand ( n15882 , n15877 , n15881 );
buf ( n15883 , n15882 );
buf ( n15884 , n15883 );
nor ( n15885 , n15868 , n15884 );
buf ( n15886 , n15885 );
buf ( n15887 , n15886 );
nand ( n15888 , n15862 , n15887 );
buf ( n15889 , n15888 );
buf ( n15890 , n15889 );
buf ( n15891 , n15094 );
buf ( n15892 , n15266 );
nand ( n15893 , n15891 , n15892 );
buf ( n15894 , n15893 );
buf ( n15895 , n15894 );
xnor ( n15896 , n15890 , n15895 );
buf ( n15897 , n15896 );
buf ( n15898 , n15897 );
not ( n15899 , n15898 );
or ( n15900 , n15843 , n15899 );
nand ( n15901 , n277817 , n9527 );
nand ( n15902 , n15900 , n15901 );
nand ( n15903 , n15522 , n15902 );
nand ( n15904 , n15842 , n15903 );
buf ( n15905 , n15904 );
nor ( n15906 , n15841 , n15905 );
or ( n15907 , n15837 , n15906 );
and ( n15908 , n15831 , n15907 );
nand ( n15909 , n15793 , n15908 );
not ( n15910 , n277910 );
buf ( n15911 , n15004 );
not ( n15912 , n15911 );
buf ( n15913 , n15472 );
nand ( n15914 , n15912 , n15913 );
buf ( n15915 , n15914 );
buf ( n15916 , n15915 );
not ( n15917 , n15916 );
buf ( n15918 , n14990 );
not ( n15919 , n15918 );
buf ( n15920 , n14997 );
nor ( n15921 , n15919 , n15920 );
buf ( n15922 , n15921 );
buf ( n15923 , n15922 );
buf ( n15924 , n14973 );
and ( n15925 , n15923 , n15924 );
buf ( n15926 , n15925 );
buf ( n15927 , n15926 );
not ( n15928 , n15927 );
buf ( n15929 , n15387 );
not ( n15930 , n15929 );
or ( n15931 , n15928 , n15930 );
buf ( n15932 , n15436 );
buf ( n15933 , n15922 );
and ( n15934 , n15932 , n15933 );
buf ( n15935 , n15458 );
not ( n15936 , n15935 );
buf ( n15937 , n15936 );
buf ( n15938 , n15937 );
buf ( n15939 , n14997 );
or ( n15940 , n15938 , n15939 );
buf ( n15941 , n15465 );
nand ( n15942 , n15940 , n15941 );
buf ( n15943 , n15942 );
buf ( n15944 , n15943 );
nor ( n15945 , n15934 , n15944 );
buf ( n15946 , n15945 );
buf ( n15947 , n15946 );
nand ( n15948 , n15931 , n15947 );
buf ( n15949 , n15948 );
buf ( n15950 , n15949 );
not ( n15951 , n15950 );
or ( n15952 , n15917 , n15951 );
buf ( n15953 , n15949 );
buf ( n15954 , n15915 );
or ( n15955 , n15953 , n15954 );
nand ( n15956 , n15952 , n15955 );
buf ( n15957 , n15956 );
buf ( n15958 , n15957 );
not ( n15959 , n15958 );
or ( n15960 , n15910 , n15959 );
nand ( n15961 , n277527 , n9688 );
nand ( n15962 , n15960 , n15961 );
and ( n15963 , n15572 , n15962 );
buf ( n15964 , n15963 );
not ( n15965 , n15964 );
buf ( n15966 , n13813 );
buf ( n15967 , n15966 );
not ( n15968 , n15967 );
or ( n15969 , n15965 , n15968 );
not ( n15970 , n15967 );
not ( n15971 , n15964 );
nand ( n15972 , n15970 , n15971 );
nand ( n15973 , n15969 , n15972 );
not ( n15974 , n277910 );
buf ( n15975 , n14997 );
not ( n15976 , n15975 );
buf ( n15977 , n15465 );
nand ( n15978 , n15976 , n15977 );
buf ( n15979 , n15978 );
buf ( n15980 , n15979 );
not ( n15981 , n15980 );
buf ( n15982 , n14973 );
buf ( n15983 , n14990 );
and ( n15984 , n15982 , n15983 );
buf ( n15985 , n15984 );
buf ( n15986 , n15985 );
not ( n15987 , n15986 );
buf ( n15988 , n15387 );
not ( n15989 , n15988 );
or ( n15990 , n15987 , n15989 );
buf ( n15991 , n15436 );
buf ( n15992 , n14990 );
and ( n15993 , n15991 , n15992 );
buf ( n15994 , n15458 );
nor ( n15995 , n15993 , n15994 );
buf ( n15996 , n15995 );
buf ( n15997 , n15996 );
nand ( n15998 , n15990 , n15997 );
buf ( n15999 , n15998 );
buf ( n16000 , n15999 );
not ( n16001 , n16000 );
or ( n16002 , n15981 , n16001 );
buf ( n16003 , n15999 );
buf ( n16004 , n15979 );
or ( n16005 , n16003 , n16004 );
nand ( n16006 , n16002 , n16005 );
buf ( n16007 , n16006 );
buf ( n16008 , n16007 );
not ( n16009 , n16008 );
or ( n16010 , n15974 , n16009 );
nand ( n16011 , n277603 , n9696 );
nand ( n16012 , n16010 , n16011 );
and ( n16013 , n14918 , n16012 );
buf ( n16014 , n16013 );
not ( n16015 , n16014 );
buf ( n16016 , n13883 );
buf ( n16017 , n16016 );
and ( n16018 , n16015 , n16017 );
nor ( n16019 , n15973 , n16018 );
not ( n16020 , n16019 );
not ( n16021 , n16014 );
not ( n16022 , n16017 );
or ( n16023 , n16021 , n16022 );
not ( n16024 , n16017 );
nand ( n16025 , n16024 , n16015 );
nand ( n16026 , n16023 , n16025 );
buf ( n16027 , n13836 );
buf ( n16028 , n16027 );
not ( n16029 , n277910 );
buf ( n16030 , n14973 );
buf ( n16031 , n14987 );
not ( n16032 , n16031 );
buf ( n16033 , n16032 );
buf ( n16034 , n16033 );
and ( n16035 , n16030 , n16034 );
buf ( n16036 , n16035 );
buf ( n16037 , n16036 );
not ( n16038 , n16037 );
buf ( n16039 , n15386 );
not ( n16040 , n16039 );
or ( n16041 , n16038 , n16040 );
buf ( n16042 , n15436 );
buf ( n16043 , n16033 );
and ( n16044 , n16042 , n16043 );
buf ( n16045 , n15443 );
nor ( n16046 , n16044 , n16045 );
buf ( n16047 , n16046 );
buf ( n16048 , n16047 );
nand ( n16049 , n16041 , n16048 );
buf ( n16050 , n16049 );
buf ( n16051 , n16050 );
buf ( n16052 , n15448 );
buf ( n16053 , n15455 );
nand ( n16054 , n16052 , n16053 );
buf ( n16055 , n16054 );
buf ( n16056 , n16055 );
not ( n16057 , n16056 );
buf ( n16058 , n16057 );
buf ( n16059 , n16058 );
and ( n16060 , n16051 , n16059 );
not ( n16061 , n16051 );
buf ( n16062 , n16055 );
and ( n16063 , n16061 , n16062 );
nor ( n16064 , n16060 , n16063 );
buf ( n16065 , n16064 );
buf ( n16066 , n16065 );
not ( n16067 , n16066 );
or ( n16068 , n16029 , n16067 );
nand ( n16069 , n277352 , n9671 );
nand ( n16070 , n16068 , n16069 );
nand ( n16071 , n15523 , n16070 );
not ( n16072 , n16071 );
buf ( n16073 , n16072 );
not ( n16074 , n16073 );
and ( n16075 , n16028 , n16074 );
or ( n16076 , n16026 , n16075 );
nand ( n16077 , n16020 , n16076 );
not ( n16078 , n16077 );
not ( n16079 , n16073 );
not ( n16080 , n16028 );
or ( n16081 , n16079 , n16080 );
not ( n16082 , n16028 );
nand ( n16083 , n16082 , n16074 );
nand ( n16084 , n16081 , n16083 );
buf ( n16085 , n13928 );
buf ( n16086 , n16085 );
not ( n16087 , n9433 );
buf ( n16088 , n15443 );
not ( n16089 , n16088 );
buf ( n16090 , n16033 );
nand ( n16091 , n16089 , n16090 );
buf ( n16092 , n16091 );
buf ( n16093 , n16092 );
not ( n16094 , n16093 );
buf ( n16095 , n14973 );
not ( n16096 , n16095 );
buf ( n16097 , n15386 );
not ( n16098 , n16097 );
or ( n16099 , n16096 , n16098 );
buf ( n16100 , n15436 );
not ( n16101 , n16100 );
buf ( n16102 , n16101 );
buf ( n16103 , n16102 );
nand ( n16104 , n16099 , n16103 );
buf ( n16105 , n16104 );
buf ( n16106 , n16105 );
not ( n16107 , n16106 );
or ( n16108 , n16094 , n16107 );
buf ( n16109 , n16105 );
buf ( n16110 , n16092 );
or ( n16111 , n16109 , n16110 );
nand ( n16112 , n16108 , n16111 );
buf ( n16113 , n16112 );
buf ( n16114 , n16113 );
not ( n16115 , n16114 );
or ( n16116 , n16087 , n16115 );
nand ( n16117 , n277352 , n9679 );
nand ( n16118 , n16116 , n16117 );
nand ( n16119 , n15629 , n16118 );
not ( n16120 , n16119 );
buf ( n16121 , n16120 );
not ( n16122 , n16121 );
and ( n16123 , n16086 , n16122 );
nor ( n16124 , n16084 , n16123 );
not ( n16125 , n16124 );
not ( n16126 , n16121 );
not ( n16127 , n16086 );
or ( n16128 , n16126 , n16127 );
not ( n16129 , n16086 );
nand ( n16130 , n16129 , n16122 );
nand ( n16131 , n16128 , n16130 );
not ( n16132 , n16131 );
and ( n16133 , n15785 , n15734 );
not ( n16134 , n16133 );
nand ( n16135 , n16132 , n16134 );
nand ( n16136 , n16125 , n16135 );
not ( n16137 , n16136 );
nand ( n16138 , n16078 , n16137 );
nor ( n16139 , n15909 , n16138 );
not ( n16140 , n16139 );
not ( n16141 , n15558 );
not ( n16142 , n15562 );
or ( n16143 , n16141 , n16142 );
not ( n16144 , n15562 );
nand ( n16145 , n15559 , n16144 );
nand ( n16146 , n16143 , n16145 );
and ( n16147 , n15967 , n15971 );
nor ( n16148 , n16146 , n16147 );
nor ( n16149 , n16140 , n16148 );
not ( n16150 , n16149 );
buf ( n16151 , n13466 );
buf ( n16152 , n16151 );
not ( n16153 , n16152 );
not ( n16154 , n16153 );
nand ( n16155 , n14915 , n14916 );
buf ( n16156 , n16155 );
not ( n16157 , n16156 );
not ( n16158 , n13004 );
and ( n16159 , n16157 , n16158 );
not ( n16160 , n277390 );
buf ( n16161 , n15062 );
buf ( n16162 , n15119 );
not ( n16163 , n16162 );
buf ( n16164 , n16163 );
buf ( n16165 , n16164 );
and ( n16166 , n16161 , n16165 );
buf ( n16167 , n16166 );
buf ( n16168 , n16167 );
not ( n16169 , n16168 );
buf ( n16170 , n15859 );
not ( n16171 , n16170 );
or ( n16172 , n16169 , n16171 );
buf ( n16173 , n15081 );
buf ( n16174 , n16164 );
and ( n16175 , n16173 , n16174 );
buf ( n16176 , n15314 );
nor ( n16177 , n16175 , n16176 );
buf ( n16178 , n16177 );
buf ( n16179 , n16178 );
nand ( n16180 , n16172 , n16179 );
buf ( n16181 , n16180 );
buf ( n16182 , n16181 );
buf ( n16183 , n15308 );
buf ( n16184 , n15321 );
nand ( n16185 , n16183 , n16184 );
buf ( n16186 , n16185 );
buf ( n16187 , n16186 );
not ( n16188 , n16187 );
buf ( n16189 , n16188 );
buf ( n16190 , n16189 );
and ( n16191 , n16182 , n16190 );
not ( n16192 , n16182 );
buf ( n16193 , n16186 );
and ( n16194 , n16192 , n16193 );
nor ( n16195 , n16191 , n16194 );
buf ( n16196 , n16195 );
buf ( n16197 , n16196 );
not ( n16198 , n16197 );
or ( n16199 , n16160 , n16198 );
nand ( n16200 , n277527 , n9535 );
nand ( n16201 , n16199 , n16200 );
and ( n16202 , n15624 , n16201 );
nor ( n16203 , n16159 , n16202 );
not ( n16204 , n16203 );
buf ( n16205 , n16204 );
not ( n16206 , n16205 );
not ( n16207 , n16206 );
or ( n16208 , n16154 , n16207 );
nand ( n16209 , n16205 , n16152 );
nand ( n16210 , n16208 , n16209 );
buf ( n16211 , n13483 );
buf ( n16212 , n16211 );
buf ( n16213 , n16212 );
or ( n16214 , n15572 , n13121 );
not ( n16215 , n277983 );
buf ( n16216 , n15062 );
not ( n16217 , n16216 );
buf ( n16218 , n15859 );
not ( n16219 , n16218 );
or ( n16220 , n16217 , n16219 );
buf ( n16221 , n15084 );
nand ( n16222 , n16220 , n16221 );
buf ( n16223 , n16222 );
buf ( n16224 , n16223 );
buf ( n16225 , n15314 );
not ( n16226 , n16225 );
buf ( n16227 , n16164 );
nand ( n16228 , n16226 , n16227 );
buf ( n16229 , n16228 );
buf ( n16230 , n16229 );
xnor ( n16231 , n16224 , n16230 );
buf ( n16232 , n16231 );
buf ( n16233 , n16232 );
not ( n16234 , n16233 );
or ( n16235 , n16215 , n16234 );
nand ( n16236 , n277817 , n9570 );
nand ( n16237 , n16235 , n16236 );
nand ( n16238 , n16156 , n16237 );
nand ( n16239 , n16214 , n16238 );
buf ( n16240 , n16239 );
buf ( n16241 , n16240 );
not ( n16242 , n16241 );
nand ( n16243 , n16213 , n16242 );
not ( n16244 , n16243 );
nor ( n16245 , n16210 , n16244 );
not ( n16246 , n16213 );
not ( n16247 , n16246 );
not ( n16248 , n16242 );
or ( n16249 , n16247 , n16248 );
nand ( n16250 , n16213 , n16241 );
nand ( n16251 , n16249 , n16250 );
or ( n16252 , n15522 , n13141 );
not ( n16253 , n277390 );
buf ( n16254 , n15052 );
buf ( n16255 , n15078 );
nand ( n16256 , n16254 , n16255 );
buf ( n16257 , n16256 );
buf ( n16258 , n16257 );
not ( n16259 , n16258 );
buf ( n16260 , n15059 );
not ( n16261 , n16260 );
buf ( n16262 , n15859 );
not ( n16263 , n16262 );
or ( n16264 , n16261 , n16263 );
buf ( n16265 , n15069 );
not ( n16266 , n16265 );
buf ( n16267 , n16266 );
buf ( n16268 , n16267 );
nand ( n16269 , n16264 , n16268 );
buf ( n16270 , n16269 );
buf ( n16271 , n16270 );
not ( n16272 , n16271 );
or ( n16273 , n16259 , n16272 );
buf ( n16274 , n16270 );
buf ( n16275 , n16257 );
or ( n16276 , n16274 , n16275 );
nand ( n16277 , n16273 , n16276 );
buf ( n16278 , n16277 );
buf ( n16279 , n16278 );
not ( n16280 , n16279 );
or ( n16281 , n16253 , n16280 );
not ( n16282 , n277350 );
not ( n16283 , n16282 );
nand ( n16284 , n16283 , n9509 );
nand ( n16285 , n16281 , n16284 );
nand ( n16286 , n16156 , n16285 );
nand ( n16287 , n16252 , n16286 );
buf ( n16288 , n16287 );
not ( n16289 , n16288 );
buf ( n16290 , n13622 );
buf ( n16291 , n16290 );
and ( n16292 , n16289 , n16291 );
nor ( n16293 , n16251 , n16292 );
nor ( n16294 , n16245 , n16293 );
buf ( n16295 , n13637 );
buf ( n16296 , n16295 );
buf ( n16297 , n16296 );
not ( n16298 , n16297 );
not ( n16299 , n16155 );
not ( n16300 , n16299 );
or ( n16301 , n16300 , n13155 );
not ( n16302 , n277910 );
buf ( n16303 , n15059 );
buf ( n16304 , n16267 );
nand ( n16305 , n16303 , n16304 );
buf ( n16306 , n16305 );
buf ( n16307 , n16306 );
not ( n16308 , n16307 );
buf ( n16309 , n15859 );
not ( n16310 , n16309 );
or ( n16311 , n16308 , n16310 );
buf ( n16312 , n15859 );
buf ( n16313 , n16306 );
or ( n16314 , n16312 , n16313 );
nand ( n16315 , n16311 , n16314 );
buf ( n16316 , n16315 );
buf ( n16317 , n16316 );
not ( n16318 , n16317 );
or ( n16319 , n16302 , n16318 );
nand ( n16320 , n277817 , n9517 );
nand ( n16321 , n16319 , n16320 );
nand ( n16322 , n16156 , n16321 );
nand ( n16323 , n16301 , n16322 );
buf ( n16324 , n16323 );
not ( n16325 , n16324 );
or ( n16326 , n16298 , n16325 );
not ( n16327 , n16324 );
not ( n16328 , n16297 );
nand ( n16329 , n16327 , n16328 );
nand ( n16330 , n16326 , n16329 );
buf ( n16331 , n13580 );
buf ( n16332 , n16331 );
buf ( n16333 , n16332 );
not ( n16334 , n16333 );
not ( n16335 , n277910 );
buf ( n16336 , n15374 );
not ( n16337 , n16336 );
buf ( n16338 , n15031 );
nand ( n16339 , n16337 , n16338 );
buf ( n16340 , n16339 );
buf ( n16341 , n16340 );
not ( n16342 , n16341 );
buf ( n16343 , n15165 );
buf ( n16344 , n15041 );
and ( n16345 , n16343 , n16344 );
buf ( n16346 , n16345 );
buf ( n16347 , n16346 );
not ( n16348 , n16347 );
buf ( n16349 , n15240 );
not ( n16350 , n16349 );
buf ( n16351 , n15227 );
not ( n16352 , n16351 );
or ( n16353 , n16350 , n16352 );
buf ( n16354 , n15191 );
not ( n16355 , n16354 );
buf ( n16356 , n16355 );
buf ( n16357 , n16356 );
nand ( n16358 , n16353 , n16357 );
buf ( n16359 , n16358 );
buf ( n16360 , n16359 );
not ( n16361 , n16360 );
or ( n16362 , n16348 , n16361 );
buf ( n16363 , n15359 );
buf ( n16364 , n15041 );
and ( n16365 , n16363 , n16364 );
buf ( n16366 , n15368 );
nor ( n16367 , n16365 , n16366 );
buf ( n16368 , n16367 );
buf ( n16369 , n16368 );
nand ( n16370 , n16362 , n16369 );
buf ( n16371 , n16370 );
buf ( n16372 , n16371 );
not ( n16373 , n16372 );
or ( n16374 , n16342 , n16373 );
buf ( n16375 , n16371 );
buf ( n16376 , n16340 );
or ( n16377 , n16375 , n16376 );
nand ( n16378 , n16374 , n16377 );
buf ( n16379 , n16378 );
buf ( n16380 , n16379 );
not ( n16381 , n16380 );
or ( n16382 , n16335 , n16381 );
nand ( n16383 , n277352 , n9552 );
nand ( n16384 , n16382 , n16383 );
not ( n16385 , n16384 );
not ( n16386 , n16156 );
or ( n16387 , n16385 , n16386 );
nand ( n16388 , n16299 , n12936 );
nand ( n16389 , n16387 , n16388 );
buf ( n16390 , n16389 );
nor ( n16391 , n16334 , n16390 );
nor ( n16392 , n16330 , n16391 );
not ( n16393 , n16291 );
not ( n16394 , n16393 );
not ( n16395 , n16289 );
or ( n16396 , n16394 , n16395 );
nand ( n16397 , n16288 , n16291 );
nand ( n16398 , n16396 , n16397 );
nor ( n16399 , n16324 , n16328 );
nor ( n16400 , n16398 , n16399 );
nor ( n16401 , n16392 , n16400 );
and ( n16402 , n16294 , n16401 );
not ( n16403 , n16333 );
not ( n16404 , n16390 );
nand ( n16405 , n16403 , n16404 );
nand ( n16406 , n16333 , n16390 );
nand ( n16407 , n16405 , n16406 );
not ( n16408 , n13019 );
not ( n16409 , n15521 );
or ( n16410 , n16408 , n16409 );
buf ( n16411 , n15165 );
not ( n16412 , n16411 );
buf ( n16413 , n16359 );
not ( n16414 , n16413 );
or ( n16415 , n16412 , n16414 );
buf ( n16416 , n15359 );
not ( n16417 , n16416 );
buf ( n16418 , n16417 );
buf ( n16419 , n16418 );
nand ( n16420 , n16415 , n16419 );
buf ( n16421 , n16420 );
buf ( n16422 , n16421 );
buf ( n16423 , n15368 );
not ( n16424 , n16423 );
buf ( n16425 , n15041 );
nand ( n16426 , n16424 , n16425 );
buf ( n16427 , n16426 );
buf ( n16428 , n16427 );
xnor ( n16429 , n16422 , n16428 );
buf ( n16430 , n16429 );
buf ( n16431 , n16430 );
not ( n16432 , n16431 );
or ( n16433 , n16432 , n9432 );
nand ( n16434 , n277352 , n9587 );
nand ( n16435 , n16433 , n16434 );
nand ( n16436 , n16300 , n16435 );
nand ( n16437 , n16410 , n16436 );
buf ( n16438 , n16437 );
buf ( n16439 , n13598 );
buf ( n16440 , n16439 );
buf ( n16441 , n16440 );
not ( n16442 , n16441 );
nor ( n16443 , n16438 , n16442 );
nor ( n16444 , n16407 , n16443 );
not ( n16445 , n16444 );
not ( n16446 , n16441 );
not ( n16447 , n16438 );
or ( n16448 , n16446 , n16447 );
not ( n16449 , n16438 );
nand ( n16450 , n16449 , n16442 );
nand ( n16451 , n16448 , n16450 );
not ( n16452 , n16156 );
not ( n16453 , n13033 );
not ( n16454 , n16453 );
and ( n16455 , n16452 , n16454 );
buf ( n16456 , n15159 );
not ( n16457 , n16456 );
buf ( n16458 , n16359 );
not ( n16459 , n16458 );
or ( n16460 , n16457 , n16459 );
buf ( n16461 , n15349 );
not ( n16462 , n16461 );
buf ( n16463 , n16462 );
buf ( n16464 , n16463 );
nand ( n16465 , n16460 , n16464 );
buf ( n16466 , n16465 );
buf ( n16467 , n16466 );
buf ( n16468 , n15152 );
buf ( n16469 , n15356 );
nand ( n16470 , n16468 , n16469 );
buf ( n16471 , n16470 );
buf ( n16472 , n16471 );
xnor ( n16473 , n16467 , n16472 );
buf ( n16474 , n16473 );
buf ( n16475 , n16474 );
not ( n16476 , n16475 );
or ( n16477 , n16476 , n277352 );
nand ( n16478 , n9432 , n9500 );
nand ( n16479 , n16477 , n16478 );
and ( n16480 , n15624 , n16479 );
nor ( n16481 , n16455 , n16480 );
not ( n16482 , n16481 );
buf ( n16483 , n16482 );
buf ( n16484 , n13684 );
buf ( n16485 , n16484 );
buf ( n16486 , n16485 );
not ( n16487 , n16486 );
nor ( n16488 , n16483 , n16487 );
nand ( n16489 , n16451 , n16488 );
not ( n16490 , n16489 );
and ( n16491 , n16445 , n16490 );
nand ( n16492 , n16407 , n16443 );
not ( n16493 , n16492 );
nor ( n16494 , n16491 , n16493 );
not ( n16495 , n16451 );
not ( n16496 , n16488 );
nand ( n16497 , n16495 , n16496 );
not ( n16498 , n16444 );
nand ( n16499 , n16497 , n16498 );
nand ( n16500 , n16494 , n16499 );
not ( n16501 , n15840 );
not ( n16502 , n16501 );
not ( n16503 , n15905 );
not ( n16504 , n16503 );
or ( n16505 , n16502 , n16504 );
nand ( n16506 , n15905 , n15840 );
nand ( n16507 , n16505 , n16506 );
buf ( n16508 , n13535 );
buf ( n16509 , n16508 );
buf ( n16510 , n16509 );
not ( n16511 , n16510 );
or ( n16512 , n15624 , n13190 );
not ( n16513 , n9431 );
buf ( n16514 , n15340 );
not ( n16515 , n16514 );
buf ( n16516 , n16515 );
buf ( n16517 , n16516 );
buf ( n16518 , n15142 );
nor ( n16519 , n16517 , n16518 );
buf ( n16520 , n16519 );
buf ( n16521 , n16520 );
not ( n16522 , n16521 );
buf ( n16523 , n15859 );
not ( n16524 , n16523 );
or ( n16525 , n16522 , n16524 );
buf ( n16526 , n15865 );
buf ( n16527 , n15142 );
not ( n16528 , n16527 );
buf ( n16529 , n16528 );
buf ( n16530 , n16529 );
and ( n16531 , n16526 , n16530 );
buf ( n16532 , n15874 );
nor ( n16533 , n16531 , n16532 );
buf ( n16534 , n16533 );
buf ( n16535 , n16534 );
nand ( n16536 , n16525 , n16535 );
buf ( n16537 , n16536 );
buf ( n16538 , n16537 );
buf ( n16539 , n15101 );
buf ( n16540 , n15880 );
nand ( n16541 , n16539 , n16540 );
buf ( n16542 , n16541 );
buf ( n16543 , n16542 );
xnor ( n16544 , n16538 , n16543 );
buf ( n16545 , n16544 );
buf ( n16546 , n16545 );
not ( n16547 , n16546 );
or ( n16548 , n16513 , n16547 );
nand ( n16549 , n277817 , n9562 );
nand ( n16550 , n16548 , n16549 );
nand ( n16551 , n15522 , n16550 );
nand ( n16552 , n16512 , n16551 );
buf ( n16553 , n16552 );
buf ( n16554 , n16553 );
nor ( n16555 , n16511 , n16554 );
nor ( n16556 , n16507 , n16555 );
not ( n16557 , n16554 );
not ( n16558 , n16557 );
not ( n16559 , n16511 );
or ( n16560 , n16558 , n16559 );
nand ( n16561 , n16554 , n16510 );
nand ( n16562 , n16560 , n16561 );
not ( n16563 , n15572 );
not ( n16564 , n13205 );
not ( n16565 , n16564 );
and ( n16566 , n16563 , n16565 );
not ( n16567 , n277390 );
buf ( n16568 , n16516 );
buf ( n16569 , n15139 );
not ( n16570 , n16569 );
buf ( n16571 , n16570 );
buf ( n16572 , n16571 );
nor ( n16573 , n16568 , n16572 );
buf ( n16574 , n16573 );
buf ( n16575 , n16574 );
not ( n16576 , n16575 );
buf ( n16577 , n15859 );
not ( n16578 , n16577 );
or ( n16579 , n16576 , n16578 );
buf ( n16580 , n15865 );
buf ( n16581 , n15139 );
and ( n16582 , n16580 , n16581 );
buf ( n16583 , n15284 );
nor ( n16584 , n16582 , n16583 );
buf ( n16585 , n16584 );
buf ( n16586 , n16585 );
nand ( n16587 , n16579 , n16586 );
buf ( n16588 , n16587 );
buf ( n16589 , n16588 );
buf ( n16590 , n15132 );
buf ( n16591 , n15261 );
nand ( n16592 , n16590 , n16591 );
buf ( n16593 , n16592 );
buf ( n16594 , n16593 );
not ( n16595 , n16594 );
buf ( n16596 , n16595 );
buf ( n16597 , n16596 );
and ( n16598 , n16589 , n16597 );
not ( n16599 , n16589 );
buf ( n16600 , n16593 );
and ( n16601 , n16599 , n16600 );
nor ( n16602 , n16598 , n16601 );
buf ( n16603 , n16602 );
buf ( n16604 , n16603 );
not ( n16605 , n16604 );
or ( n16606 , n16567 , n16605 );
nand ( n16607 , n277527 , n9544 );
nand ( n16608 , n16606 , n16607 );
and ( n16609 , n15629 , n16608 );
nor ( n16610 , n16566 , n16609 );
not ( n16611 , n16610 );
buf ( n16612 , n16611 );
buf ( n16613 , n13708 );
buf ( n16614 , n16613 );
buf ( n16615 , n16614 );
not ( n16616 , n16615 );
nor ( n16617 , n16612 , n16616 );
nor ( n16618 , n16562 , n16617 );
nor ( n16619 , n16556 , n16618 );
or ( n16620 , n15624 , n13173 );
not ( n16621 , n277390 );
buf ( n16622 , n15340 );
not ( n16623 , n16622 );
buf ( n16624 , n15859 );
not ( n16625 , n16624 );
or ( n16626 , n16623 , n16625 );
buf ( n16627 , n15636 );
nand ( n16628 , n16626 , n16627 );
buf ( n16629 , n16628 );
buf ( n16630 , n16629 );
buf ( n16631 , n15284 );
buf ( n16632 , n16571 );
nor ( n16633 , n16631 , n16632 );
buf ( n16634 , n16633 );
buf ( n16635 , n16634 );
xor ( n16636 , n16630 , n16635 );
buf ( n16637 , n16636 );
buf ( n16638 , n16637 );
not ( n16639 , n16638 );
or ( n16640 , n16621 , n16639 );
nand ( n16641 , n277817 , n9579 );
nand ( n16642 , n16640 , n16641 );
nand ( n16643 , n15522 , n16642 );
nand ( n16644 , n16620 , n16643 );
buf ( n16645 , n16644 );
buf ( n16646 , n16645 );
not ( n16647 , n16646 );
not ( n16648 , n16647 );
buf ( n16649 , n13726 );
buf ( n16650 , n16649 );
buf ( n16651 , n16650 );
not ( n16652 , n16651 );
not ( n16653 , n16652 );
or ( n16654 , n16648 , n16653 );
nand ( n16655 , n16646 , n16651 );
nand ( n16656 , n16654 , n16655 );
buf ( n16657 , n16205 );
nor ( n16658 , n16657 , n16153 );
nor ( n16659 , n16656 , n16658 );
not ( n16660 , n16616 );
not ( n16661 , n16612 );
not ( n16662 , n16661 );
or ( n16663 , n16660 , n16662 );
nand ( n16664 , n16612 , n16615 );
nand ( n16665 , n16663 , n16664 );
nor ( n16666 , n16646 , n16652 );
nor ( n16667 , n16665 , n16666 );
nor ( n16668 , n16659 , n16667 );
nand ( n16669 , n16402 , n16500 , n16619 , n16668 );
not ( n16670 , n16669 );
not ( n16671 , n16156 );
not ( n16672 , n13100 );
and ( n16673 , n16671 , n16672 );
and ( n16674 , n277350 , n9449 );
not ( n16675 , n277350 );
buf ( n16676 , n15217 );
not ( n16677 , n16676 );
buf ( n16678 , n15209 );
buf ( n16679 , n15224 );
nand ( n16680 , n16678 , n16679 );
buf ( n16681 , n16680 );
buf ( n16682 , n16681 );
not ( n16683 , n16682 );
or ( n16684 , n16677 , n16683 );
buf ( n16685 , n16681 );
buf ( n16686 , n15217 );
or ( n16687 , n16685 , n16686 );
nand ( n16688 , n16684 , n16687 );
buf ( n16689 , n16688 );
buf ( n16690 , n16689 );
and ( n16691 , n16675 , n16690 );
or ( n16692 , n16674 , n16691 );
and ( n16693 , n15572 , n16692 );
nor ( n16694 , n16673 , n16693 );
not ( n16695 , n16694 );
buf ( n16696 , n16695 );
not ( n16697 , n16696 );
not ( n16698 , n16697 );
buf ( n16699 , n14542 );
not ( n16700 , n16699 );
not ( n16701 , n16700 );
or ( n16702 , n16698 , n16701 );
nand ( n16703 , n16699 , n16696 );
nand ( n16704 , n16702 , n16703 );
buf ( n16705 , n14775 );
buf ( n16706 , n16705 );
nand ( n16707 , n16704 , n16706 );
not ( n16708 , n16706 );
or ( n16709 , n15629 , n13103 );
and ( n16710 , n277350 , n9440 );
not ( n16711 , n277350 );
buf ( n16712 , n15212 );
buf ( n16713 , n15214 );
xor ( n16714 , n16712 , n16713 );
buf ( n16715 , n16714 );
buf ( n16716 , n16715 );
and ( n16717 , n16711 , n16716 );
or ( n16718 , n16710 , n16717 );
nand ( n16719 , n15572 , n16718 );
nand ( n16720 , n16709 , n16719 );
buf ( n16721 , n16720 );
buf ( n16722 , n16721 );
not ( n16723 , n16722 );
nand ( n16724 , n16708 , n16723 );
nand ( n16725 , n16707 , n16724 );
not ( n16726 , n16704 );
nand ( n16727 , n16726 , n16708 );
not ( n16728 , n16156 );
not ( n16729 , n13084 );
not ( n16730 , n16729 );
and ( n16731 , n16728 , n16730 );
and ( n16732 , n277817 , n9470 );
not ( n16733 , n277817 );
buf ( n16734 , n15650 );
buf ( n16735 , n15640 );
nand ( n16736 , n16734 , n16735 );
buf ( n16737 , n16736 );
buf ( n16738 , n16737 );
not ( n16739 , n16738 );
buf ( n16740 , n15227 );
not ( n16741 , n16740 );
or ( n16742 , n16739 , n16741 );
buf ( n16743 , n15227 );
buf ( n16744 , n16737 );
or ( n16745 , n16743 , n16744 );
nand ( n16746 , n16742 , n16745 );
buf ( n16747 , n16746 );
buf ( n16748 , n16747 );
and ( n16749 , n16733 , n16748 );
or ( n16750 , n16732 , n16749 );
and ( n16751 , n15572 , n16750 );
nor ( n16752 , n16731 , n16751 );
not ( n16753 , n16752 );
buf ( n16754 , n16753 );
buf ( n16755 , n14564 );
or ( n16756 , n16754 , n16755 );
nand ( n16757 , n16755 , n16754 );
nand ( n16758 , n16756 , n16757 );
and ( n16759 , n16699 , n16697 );
or ( n16760 , n16758 , n16759 );
nand ( n16761 , n16725 , n16727 , n16760 );
not ( n16762 , n16761 );
buf ( n16763 , n13601 );
buf ( n16764 , n16763 );
buf ( n16765 , n13564 );
buf ( n16766 , n16765 );
buf ( n16767 , n16766 );
xor ( n16768 , n16764 , n16767 );
not ( n16769 , n13067 );
or ( n16770 , n16156 , n16769 );
not ( n16771 , n277351 );
buf ( n16772 , n15173 );
buf ( n16773 , n15188 );
nand ( n16774 , n16772 , n16773 );
buf ( n16775 , n16774 );
buf ( n16776 , n16775 );
not ( n16777 , n16776 );
buf ( n16778 , n15653 );
buf ( n16779 , n15640 );
nand ( n16780 , n16778 , n16779 );
buf ( n16781 , n16780 );
buf ( n16782 , n16781 );
not ( n16783 , n16782 );
or ( n16784 , n16777 , n16783 );
buf ( n16785 , n16781 );
buf ( n16786 , n16775 );
or ( n16787 , n16785 , n16786 );
nand ( n16788 , n16784 , n16787 );
buf ( n16789 , n16788 );
buf ( n16790 , n16789 );
not ( n16791 , n16790 );
or ( n16792 , n16771 , n16791 );
nand ( n16793 , n277817 , n9462 );
nand ( n16794 , n16792 , n16793 );
nand ( n16795 , n16156 , n16794 );
nand ( n16796 , n16770 , n16795 );
buf ( n16797 , n16796 );
not ( n16798 , n16797 );
xor ( n16799 , n16768 , n16798 );
not ( n16800 , n16755 );
nor ( n16801 , n16800 , n16754 );
nand ( n16802 , n16799 , n16801 );
nand ( n16803 , n16758 , n16759 );
and ( n16804 , n16802 , n16803 );
not ( n16805 , n16804 );
or ( n16806 , n16762 , n16805 );
not ( n16807 , n16486 );
not ( n16808 , n16483 );
or ( n16809 , n16807 , n16808 );
not ( n16810 , n16483 );
nand ( n16811 , n16810 , n16487 );
nand ( n16812 , n16809 , n16811 );
not ( n16813 , n16812 );
buf ( n16814 , n13659 );
not ( n16815 , n16814 );
not ( n16816 , n16815 );
buf ( n16817 , n16816 );
not ( n16818 , n16817 );
not ( n16819 , n16156 );
not ( n16820 , n13049 );
not ( n16821 , n16820 );
and ( n16822 , n16819 , n16821 );
not ( n16823 , n277390 );
buf ( n16824 , n15159 );
buf ( n16825 , n16463 );
nand ( n16826 , n16824 , n16825 );
buf ( n16827 , n16826 );
buf ( n16828 , n16827 );
not ( n16829 , n16828 );
buf ( n16830 , n16359 );
not ( n16831 , n16830 );
or ( n16832 , n16829 , n16831 );
buf ( n16833 , n16359 );
buf ( n16834 , n16827 );
or ( n16835 , n16833 , n16834 );
nand ( n16836 , n16832 , n16835 );
buf ( n16837 , n16836 );
buf ( n16838 , n16837 );
not ( n16839 , n16838 );
or ( n16840 , n16823 , n16839 );
nand ( n16841 , n277603 , n9492 );
nand ( n16842 , n16840 , n16841 );
and ( n16843 , n15572 , n16842 );
nor ( n16844 , n16822 , n16843 );
not ( n16845 , n16844 );
buf ( n16846 , n16845 );
nor ( n16847 , n16818 , n16846 );
not ( n16848 , n16847 );
nand ( n16849 , n16813 , n16848 );
xor ( n16850 , n16764 , n16767 );
and ( n16851 , n16850 , n16798 );
and ( n16852 , n16764 , n16767 );
or ( n16853 , n16851 , n16852 );
not ( n16854 , n16853 );
not ( n16855 , n16846 );
and ( n16856 , n16817 , n16855 );
not ( n16857 , n16817 );
and ( n16858 , n16857 , n16846 );
nor ( n16859 , n16856 , n16858 );
not ( n16860 , n16859 );
nand ( n16861 , n16854 , n16860 );
nand ( n16862 , n16849 , n16861 );
nor ( n16863 , n16801 , n16799 );
nor ( n16864 , n16862 , n16863 );
nand ( n16865 , n16806 , n16864 );
not ( n16866 , n16853 );
nor ( n16867 , n16866 , n16860 );
not ( n16868 , n16867 );
not ( n16869 , n16849 );
or ( n16870 , n16868 , n16869 );
buf ( n16871 , n16812 );
not ( n16872 , n16848 );
nand ( n16873 , n16871 , n16872 );
nand ( n16874 , n16870 , n16873 );
not ( n16875 , n16494 );
nor ( n16876 , n16874 , n16875 );
nand ( n16877 , n16865 , n16876 );
nand ( n16878 , n16670 , n16877 );
and ( n16879 , n16562 , n16617 );
not ( n16880 , n16879 );
not ( n16881 , n16556 );
not ( n16882 , n16881 );
or ( n16883 , n16880 , n16882 );
buf ( n16884 , n16507 );
buf ( n16885 , n16555 );
nand ( n16886 , n16884 , n16885 );
nand ( n16887 , n16883 , n16886 );
nand ( n16888 , n16656 , n16658 );
or ( n16889 , n16667 , n16888 );
nand ( n16890 , n16665 , n16666 );
nand ( n16891 , n16889 , n16890 );
nor ( n16892 , n16887 , n16891 );
not ( n16893 , n16892 );
not ( n16894 , n16400 );
and ( n16895 , n16330 , n16391 );
nand ( n16896 , n16894 , n16895 );
nand ( n16897 , n16210 , n16244 );
not ( n16898 , n16897 );
and ( n16899 , n16398 , n16399 );
nor ( n16900 , n16898 , n16899 );
nand ( n16901 , n16251 , n16292 );
nand ( n16902 , n16896 , n16900 , n16901 );
and ( n16903 , n16293 , n16897 );
nor ( n16904 , n16903 , n16245 );
nand ( n16905 , n16902 , n16904 , n16668 );
not ( n16906 , n16905 );
or ( n16907 , n16893 , n16906 );
not ( n16908 , n16887 );
not ( n16909 , n16619 );
nand ( n16910 , n16908 , n16909 );
nand ( n16911 , n16907 , n16910 );
nand ( n16912 , n16878 , n16911 );
buf ( n16913 , n16912 );
not ( n16914 , n16913 );
or ( n16915 , n16150 , n16914 );
not ( n16916 , n16148 );
not ( n16917 , n16916 );
nand ( n16918 , n15837 , n15906 );
not ( n16919 , n16918 );
nand ( n16920 , n15799 , n15830 );
not ( n16921 , n16920 );
or ( n16922 , n16919 , n16921 );
nand ( n16923 , n16922 , n15831 );
nor ( n16924 , n16923 , n15792 );
not ( n16925 , n16924 );
nand ( n16926 , n16026 , n16075 );
or ( n16927 , n16019 , n16926 );
nand ( n16928 , n15973 , n16018 );
nand ( n16929 , n16927 , n16928 );
nand ( n16930 , n16131 , n16133 );
or ( n16931 , n16124 , n16930 );
nand ( n16932 , n16084 , n16123 );
nand ( n16933 , n16931 , n16932 );
nor ( n16934 , n16929 , n16933 );
and ( n16935 , n15620 , n15730 );
and ( n16936 , n15791 , n16935 );
and ( n16937 , n15787 , n15789 );
nor ( n16938 , n16936 , n16937 );
nand ( n16939 , n16925 , n16934 , n16938 );
nand ( n16940 , n16934 , n16136 );
not ( n16941 , n16929 );
nand ( n16942 , n16941 , n16077 );
and ( n16943 , n16939 , n16940 , n16942 );
not ( n16944 , n16943 );
or ( n16945 , n16917 , n16944 );
nand ( n16946 , n16146 , n16147 );
nand ( n16947 , n16945 , n16946 );
not ( n16948 , n16947 );
nand ( n16949 , n16915 , n16948 );
not ( n16950 , n16949 );
or ( n16951 , n15568 , n16950 );
or ( n16952 , n16949 , n15567 );
nand ( n16953 , n16951 , n16952 );
buf ( n16954 , n16953 );
not ( n16955 , n14886 );
nor ( n16956 , n16955 , n14894 );
not ( n16957 , n16956 );
nand ( n16958 , n14895 , n16957 );
not ( n16959 , n16958 );
and ( n16960 , n14894 , n14905 );
not ( n16961 , n14894 );
and ( n16962 , n16961 , n14900 );
nor ( n16963 , n16960 , n16962 );
nand ( n16964 , n14831 , n16959 , n16963 );
not ( n16965 , n14858 );
not ( n16966 , n16965 );
nand ( n16967 , n14868 , n16966 , n14839 );
nor ( n16968 , n16964 , n16967 );
not ( n16969 , n16968 );
not ( n16970 , n16969 );
nand ( n16971 , n16954 , n16970 );
buf ( n16972 , n15509 );
buf ( n16973 , n15513 );
xor ( n16974 , n16972 , n16973 );
buf ( n16975 , n15560 );
buf ( n16976 , n16975 );
buf ( n16977 , n15557 );
and ( n16978 , n16976 , n16977 );
nor ( n16979 , n16974 , n16978 );
not ( n16980 , n16979 );
nand ( n16981 , n16974 , n16978 );
nand ( n16982 , n16980 , n16981 );
not ( n16983 , n16982 );
buf ( n16984 , n15728 );
not ( n16985 , n16984 );
not ( n16986 , n16985 );
buf ( n16987 , n15621 );
not ( n16988 , n16987 );
or ( n16989 , n16986 , n16988 );
not ( n16990 , n16987 );
nand ( n16991 , n16990 , n16984 );
nand ( n16992 , n16989 , n16991 );
buf ( n16993 , n15800 );
buf ( n16994 , n15828 );
and ( n16995 , n16993 , n16994 );
nor ( n16996 , n16992 , n16995 );
not ( n16997 , n16994 );
not ( n16998 , n16997 );
not ( n16999 , n16993 );
or ( n17000 , n16998 , n16999 );
not ( n17001 , n16993 );
nand ( n17002 , n16994 , n17001 );
nand ( n17003 , n17000 , n17002 );
buf ( n17004 , n15904 );
buf ( n17005 , n15838 );
and ( n17006 , n17004 , n17005 );
nor ( n17007 , n17003 , n17006 );
nor ( n17008 , n16996 , n17007 );
buf ( n17009 , n15613 );
not ( n17010 , n17009 );
buf ( n17011 , n15569 );
buf ( n17012 , n17011 );
not ( n17013 , n17012 );
not ( n17014 , n17013 );
or ( n17015 , n17010 , n17014 );
not ( n17016 , n17009 );
nand ( n17017 , n17016 , n17012 );
nand ( n17018 , n17015 , n17017 );
and ( n17019 , n16987 , n16984 );
nor ( n17020 , n17018 , n17019 );
buf ( n17021 , n15733 );
not ( n17022 , n17021 );
not ( n17023 , n17022 );
buf ( n17024 , n15780 );
not ( n17025 , n17024 );
or ( n17026 , n17023 , n17025 );
not ( n17027 , n17024 );
nand ( n17028 , n17027 , n17021 );
nand ( n17029 , n17026 , n17028 );
nand ( n17030 , n17012 , n17009 );
not ( n17031 , n17030 );
nor ( n17032 , n17029 , n17031 );
nor ( n17033 , n17020 , n17032 );
nand ( n17034 , n17008 , n17033 );
not ( n17035 , n17034 );
buf ( n17036 , n15963 );
not ( n17037 , n17036 );
buf ( n17038 , n15966 );
not ( n17039 , n17038 );
not ( n17040 , n17039 );
or ( n17041 , n17037 , n17040 );
not ( n17042 , n17036 );
nand ( n17043 , n17042 , n17038 );
nand ( n17044 , n17041 , n17043 );
buf ( n17045 , n16016 );
buf ( n17046 , n16013 );
nand ( n17047 , n17045 , n17046 );
not ( n17048 , n17047 );
nor ( n17049 , n17044 , n17048 );
not ( n17050 , n17046 );
not ( n17051 , n17050 );
not ( n17052 , n17045 );
or ( n17053 , n17051 , n17052 );
not ( n17054 , n17045 );
nand ( n17055 , n17054 , n17046 );
nand ( n17056 , n17053 , n17055 );
buf ( n17057 , n16027 );
buf ( n17058 , n16072 );
and ( n17059 , n17057 , n17058 );
nor ( n17060 , n17056 , n17059 );
nor ( n17061 , n17049 , n17060 );
not ( n17062 , n17061 );
not ( n17063 , n17058 );
not ( n17064 , n17057 );
not ( n17065 , n17064 );
or ( n17066 , n17063 , n17065 );
not ( n17067 , n17058 );
nand ( n17068 , n17057 , n17067 );
nand ( n17069 , n17066 , n17068 );
not ( n17070 , n16085 );
not ( n17071 , n17070 );
buf ( n17072 , n17071 );
buf ( n17073 , n16120 );
and ( n17074 , n17072 , n17073 );
nor ( n17075 , n17069 , n17074 );
not ( n17076 , n17075 );
not ( n17077 , n17073 );
not ( n17078 , n17072 );
not ( n17079 , n17078 );
or ( n17080 , n17077 , n17079 );
not ( n17081 , n17073 );
nand ( n17082 , n17081 , n17072 );
nand ( n17083 , n17080 , n17082 );
not ( n17084 , n17083 );
and ( n17085 , n17021 , n17024 );
not ( n17086 , n17085 );
nand ( n17087 , n17084 , n17086 );
nand ( n17088 , n17076 , n17087 );
nor ( n17089 , n17062 , n17088 );
nand ( n17090 , n17035 , n17089 );
not ( n17091 , n16976 );
nand ( n17092 , n17091 , n16977 );
not ( n17093 , n16977 );
nand ( n17094 , n17093 , n16976 );
nand ( n17095 , n17092 , n17094 );
and ( n17096 , n17038 , n17036 );
nor ( n17097 , n17095 , n17096 );
nor ( n17098 , n17090 , n17097 );
not ( n17099 , n17098 );
buf ( n17100 , n16613 );
buf ( n17101 , n16611 );
xor ( n17102 , n17100 , n17101 );
not ( n17103 , n17102 );
buf ( n17104 , n16644 );
buf ( n17105 , n16649 );
and ( n17106 , n17104 , n17105 );
not ( n17107 , n17106 );
nand ( n17108 , n17103 , n17107 );
not ( n17109 , n17105 );
not ( n17110 , n17104 );
not ( n17111 , n17110 );
or ( n17112 , n17109 , n17111 );
not ( n17113 , n17105 );
nand ( n17114 , n17104 , n17113 );
nand ( n17115 , n17112 , n17114 );
buf ( n17116 , n16151 );
buf ( n17117 , n16204 );
nand ( n17118 , n17116 , n17117 );
not ( n17119 , n17118 );
or ( n17120 , n17115 , n17119 );
and ( n17121 , n17108 , n17120 );
not ( n17122 , n17005 );
not ( n17123 , n17004 );
not ( n17124 , n17123 );
or ( n17125 , n17122 , n17124 );
not ( n17126 , n17005 );
nand ( n17127 , n17004 , n17126 );
nand ( n17128 , n17125 , n17127 );
buf ( n17129 , n16552 );
buf ( n17130 , n16508 );
nand ( n17131 , n17129 , n17130 );
not ( n17132 , n17131 );
nor ( n17133 , n17128 , n17132 );
not ( n17134 , n17130 );
not ( n17135 , n17134 );
not ( n17136 , n17129 );
or ( n17137 , n17135 , n17136 );
not ( n17138 , n17129 );
nand ( n17139 , n17138 , n17130 );
nand ( n17140 , n17137 , n17139 );
and ( n17141 , n17100 , n17101 );
nor ( n17142 , n17140 , n17141 );
nor ( n17143 , n17133 , n17142 );
nand ( n17144 , n17121 , n17143 );
buf ( n17145 , n16331 );
not ( n17146 , n17145 );
buf ( n17147 , n16389 );
not ( n17148 , n17147 );
not ( n17149 , n17148 );
or ( n17150 , n17146 , n17149 );
not ( n17151 , n17145 );
nand ( n17152 , n17151 , n17147 );
nand ( n17153 , n17150 , n17152 );
not ( n17154 , n17153 );
buf ( n17155 , n16439 );
buf ( n17156 , n16437 );
and ( n17157 , n17155 , n17156 );
not ( n17158 , n17157 );
nand ( n17159 , n17154 , n17158 );
not ( n17160 , n17159 );
not ( n17161 , n17155 );
not ( n17162 , n17156 );
not ( n17163 , n17162 );
or ( n17164 , n17161 , n17163 );
not ( n17165 , n17155 );
nand ( n17166 , n17165 , n17156 );
nand ( n17167 , n17164 , n17166 );
buf ( n17168 , n16482 );
buf ( n17169 , n16484 );
nand ( n17170 , n17168 , n17169 );
not ( n17171 , n17170 );
nand ( n17172 , n17167 , n17171 );
not ( n17173 , n17172 );
not ( n17174 , n17173 );
or ( n17175 , n17160 , n17174 );
or ( n17176 , n17154 , n17158 );
nand ( n17177 , n17175 , n17176 );
not ( n17178 , n17159 );
nor ( n17179 , n17167 , n17171 );
nor ( n17180 , n17178 , n17179 );
nor ( n17181 , n17177 , n17180 );
not ( n17182 , n17116 );
not ( n17183 , n17117 );
not ( n17184 , n17183 );
or ( n17185 , n17182 , n17184 );
not ( n17186 , n17116 );
nand ( n17187 , n17186 , n17117 );
nand ( n17188 , n17185 , n17187 );
buf ( n17189 , n16239 );
not ( n17190 , n17189 );
not ( n17191 , n17190 );
buf ( n17192 , n16211 );
and ( n17193 , n17191 , n17192 );
or ( n17194 , n17188 , n17193 );
not ( n17195 , n17192 );
not ( n17196 , n17190 );
or ( n17197 , n17195 , n17196 );
not ( n17198 , n17192 );
nand ( n17199 , n17189 , n17198 );
nand ( n17200 , n17197 , n17199 );
not ( n17201 , n17200 );
buf ( n17202 , n16290 );
buf ( n17203 , n17202 );
buf ( n17204 , n16287 );
and ( n17205 , n17203 , n17204 );
not ( n17206 , n17205 );
nand ( n17207 , n17201 , n17206 );
nand ( n17208 , n17194 , n17207 );
not ( n17209 , n17208 );
xor ( n17210 , n17203 , n17204 );
not ( n17211 , n17210 );
buf ( n17212 , n16323 );
buf ( n17213 , n16295 );
and ( n17214 , n17212 , n17213 );
not ( n17215 , n17214 );
nand ( n17216 , n17211 , n17215 );
not ( n17217 , n17216 );
not ( n17218 , n17213 );
not ( n17219 , n17212 );
not ( n17220 , n17219 );
or ( n17221 , n17218 , n17220 );
not ( n17222 , n17213 );
nand ( n17223 , n17212 , n17222 );
nand ( n17224 , n17221 , n17223 );
nand ( n17225 , n17145 , n17147 );
not ( n17226 , n17225 );
nor ( n17227 , n17224 , n17226 );
nor ( n17228 , n17217 , n17227 );
nand ( n17229 , n17209 , n17228 );
nor ( n17230 , n17144 , n17181 , n17229 );
not ( n17231 , n17230 );
buf ( n17232 , n16763 );
not ( n17233 , n17232 );
buf ( n17234 , n16765 );
not ( n17235 , n17234 );
not ( n17236 , n17235 );
or ( n17237 , n17233 , n17236 );
not ( n17238 , n17232 );
nand ( n17239 , n17234 , n17238 );
nand ( n17240 , n17237 , n17239 );
buf ( n17241 , n16796 );
and ( n17242 , n17240 , n17241 );
not ( n17243 , n17240 );
not ( n17244 , n17241 );
and ( n17245 , n17243 , n17244 );
nor ( n17246 , n17242 , n17245 );
not ( n17247 , n17246 );
buf ( n17248 , n14564 );
buf ( n17249 , n16753 );
and ( n17250 , n17248 , n17249 );
not ( n17251 , n17250 );
nand ( n17252 , n17247 , n17251 );
not ( n17253 , n17252 );
not ( n17254 , n17169 );
not ( n17255 , n17168 );
not ( n17256 , n17255 );
or ( n17257 , n17254 , n17256 );
not ( n17258 , n17169 );
nand ( n17259 , n17258 , n17168 );
nand ( n17260 , n17257 , n17259 );
buf ( n17261 , n16814 );
buf ( n17262 , n16845 );
nand ( n17263 , n17261 , n17262 );
not ( n17264 , n17263 );
nor ( n17265 , n17260 , n17264 );
not ( n17266 , n17265 );
not ( n17267 , n17238 );
not ( n17268 , n17235 );
or ( n17269 , n17267 , n17268 );
nand ( n17270 , n17269 , n17241 );
not ( n17271 , n17235 );
nand ( n17272 , n17271 , n17232 );
nand ( n17273 , n17270 , n17272 );
not ( n17274 , n17262 );
not ( n17275 , n17274 );
not ( n17276 , n17261 );
or ( n17277 , n17275 , n17276 );
not ( n17278 , n17261 );
nand ( n17279 , n17278 , n17262 );
nand ( n17280 , n17277 , n17279 );
or ( n17281 , n17273 , n17280 );
nand ( n17282 , n17266 , n17281 );
nor ( n17283 , n17253 , n17282 );
buf ( n17284 , n16695 );
not ( n17285 , n17284 );
buf ( n17286 , n14542 );
not ( n17287 , n17286 );
not ( n17288 , n17287 );
or ( n17289 , n17285 , n17288 );
not ( n17290 , n17284 );
nand ( n17291 , n17290 , n17286 );
nand ( n17292 , n17289 , n17291 );
buf ( n17293 , n14775 );
not ( n17294 , n17293 );
buf ( n17295 , n16720 );
not ( n17296 , n17295 );
nor ( n17297 , n17294 , n17296 );
nand ( n17298 , n17292 , n17297 );
not ( n17299 , n17298 );
not ( n17300 , n17249 );
not ( n17301 , n17248 );
not ( n17302 , n17301 );
or ( n17303 , n17300 , n17302 );
not ( n17304 , n17249 );
nand ( n17305 , n17304 , n17248 );
nand ( n17306 , n17303 , n17305 );
not ( n17307 , n17306 );
and ( n17308 , n17286 , n17284 );
not ( n17309 , n17308 );
nand ( n17310 , n17307 , n17309 );
nand ( n17311 , n17299 , n17310 );
nand ( n17312 , n17246 , n17250 );
buf ( n17313 , n17306 );
nand ( n17314 , n17313 , n17308 );
nand ( n17315 , n17311 , n17312 , n17314 );
nand ( n17316 , n17283 , n17315 );
nand ( n17317 , n17273 , n17280 );
not ( n17318 , n17317 );
not ( n17319 , n17318 );
not ( n17320 , n17266 );
or ( n17321 , n17319 , n17320 );
buf ( n17322 , n17260 );
buf ( n17323 , n17264 );
nand ( n17324 , n17322 , n17323 );
nand ( n17325 , n17321 , n17324 );
not ( n17326 , n17325 );
not ( n17327 , n17177 );
nand ( n17328 , n17326 , n17327 );
not ( n17329 , n17328 );
nand ( n17330 , n17316 , n17329 );
not ( n17331 , n17330 );
or ( n17332 , n17231 , n17331 );
nand ( n17333 , n17188 , n17193 );
nand ( n17334 , n17208 , n17333 );
nand ( n17335 , n17224 , n17226 );
not ( n17336 , n17335 );
nand ( n17337 , n17336 , n17216 );
nand ( n17338 , n17200 , n17205 );
nand ( n17339 , n17210 , n17214 );
and ( n17340 , n17338 , n17339 );
nand ( n17341 , n17337 , n17340 , n17333 );
nand ( n17342 , n17334 , n17341 );
not ( n17343 , n17342 );
not ( n17344 , n17144 );
and ( n17345 , n17343 , n17344 );
and ( n17346 , n17115 , n17119 );
not ( n17347 , n17346 );
not ( n17348 , n17108 );
or ( n17349 , n17347 , n17348 );
not ( n17350 , n17107 );
nand ( n17351 , n17350 , n17102 );
nand ( n17352 , n17349 , n17351 );
nand ( n17353 , n17352 , n17143 );
nand ( n17354 , n17140 , n17141 );
or ( n17355 , n17133 , n17354 );
nand ( n17356 , n17128 , n17132 );
nand ( n17357 , n17355 , n17356 );
not ( n17358 , n17357 );
nand ( n17359 , n17353 , n17358 );
nor ( n17360 , n17345 , n17359 );
nand ( n17361 , n17332 , n17360 );
buf ( n17362 , n17361 );
not ( n17363 , n17362 );
or ( n17364 , n17099 , n17363 );
nand ( n17365 , n17056 , n17059 );
or ( n17366 , n17049 , n17365 );
nand ( n17367 , n17044 , n17048 );
nand ( n17368 , n17366 , n17367 );
nand ( n17369 , n17083 , n17085 );
or ( n17370 , n17075 , n17369 );
nand ( n17371 , n17069 , n17074 );
nand ( n17372 , n17370 , n17371 );
nor ( n17373 , n17368 , n17372 );
and ( n17374 , n17373 , n17088 );
nor ( n17375 , n17368 , n17061 );
nor ( n17376 , n17374 , n17375 );
nand ( n17377 , n16992 , n16995 );
nand ( n17378 , n17003 , n17006 );
and ( n17379 , n17377 , n17378 );
nor ( n17380 , n17379 , n16996 );
nand ( n17381 , n17380 , n17033 );
not ( n17382 , n17032 );
nand ( n17383 , n17018 , n17019 );
not ( n17384 , n17383 );
and ( n17385 , n17382 , n17384 );
and ( n17386 , n17029 , n17031 );
nor ( n17387 , n17385 , n17386 );
nand ( n17388 , n17373 , n17381 , n17387 );
nand ( n17389 , n17376 , n17388 );
not ( n17390 , n17389 );
not ( n17391 , n17097 );
and ( n17392 , n17390 , n17391 );
nand ( n17393 , n17095 , n17096 );
not ( n17394 , n17393 );
nor ( n17395 , n17392 , n17394 );
nand ( n17396 , n17364 , n17395 );
not ( n17397 , n17396 );
or ( n17398 , n16983 , n17397 );
or ( n17399 , n17396 , n16982 );
nand ( n17400 , n17398 , n17399 );
buf ( n17401 , n17400 );
nor ( n17402 , n16958 , n16963 );
not ( n17403 , n17402 );
nor ( n17404 , n14869 , n17403 );
buf ( n17405 , n17404 );
and ( n17406 , n17401 , n17405 );
not ( n17407 , n14869 );
nand ( n17408 , n16956 , n14906 );
not ( n17409 , n17408 );
nand ( n17410 , n17407 , n17409 );
not ( n17411 , n17410 );
buf ( n17412 , n16845 );
buf ( n17413 , n16482 );
buf ( n17414 , n17413 );
or ( n17415 , n17412 , n17414 );
buf ( n17416 , n16389 );
buf ( n17417 , n17416 );
not ( n17418 , n17417 );
buf ( n17419 , n16437 );
buf ( n17420 , n17419 );
not ( n17421 , n17420 );
nand ( n17422 , n17418 , n17421 );
nor ( n17423 , n17415 , n17422 );
buf ( n17424 , n16721 );
buf ( n17425 , n16695 );
or ( n17426 , n17424 , n17425 );
buf ( n17427 , n16796 );
buf ( n17428 , n17427 );
not ( n17429 , n17428 );
buf ( n17430 , n16753 );
not ( n17431 , n17430 );
nand ( n17432 , n17429 , n17431 );
nor ( n17433 , n17426 , n17432 );
nand ( n17434 , n17423 , n17433 );
not ( n17435 , n17434 );
buf ( n17436 , n16287 );
buf ( n17437 , n17436 );
buf ( n17438 , n16323 );
buf ( n17439 , n17438 );
nor ( n17440 , n17437 , n17439 );
buf ( n17441 , n16240 );
buf ( n17442 , n17441 );
buf ( n17443 , n16204 );
buf ( n17444 , n17443 );
nor ( n17445 , n17442 , n17444 );
nand ( n17446 , n17440 , n17445 );
buf ( n17447 , n16611 );
buf ( n17448 , n17447 );
not ( n17449 , n17448 );
buf ( n17450 , n15904 );
buf ( n17451 , n17450 );
not ( n17452 , n17451 );
buf ( n17453 , n16645 );
buf ( n17454 , n17453 );
not ( n17455 , n17454 );
buf ( n17456 , n16553 );
buf ( n17457 , n17456 );
not ( n17458 , n17457 );
nand ( n17459 , n17449 , n17452 , n17455 , n17458 );
nor ( n17460 , n17446 , n17459 );
nand ( n17461 , n17435 , n17460 );
not ( n17462 , n17461 );
not ( n17463 , n17462 );
buf ( n17464 , n16072 );
buf ( n17465 , n17464 );
buf ( n17466 , n16120 );
buf ( n17467 , n17466 );
nor ( n17468 , n17465 , n17467 );
buf ( n17469 , n15828 );
buf ( n17470 , n17469 );
not ( n17471 , n17470 );
and ( n17472 , n17468 , n17471 );
buf ( n17473 , n15557 );
buf ( n17474 , n16013 );
buf ( n17475 , n17474 );
nor ( n17476 , n17473 , n17475 );
buf ( n17477 , n15780 );
buf ( n17478 , n17477 );
not ( n17479 , n17478 );
buf ( n17480 , n15728 );
buf ( n17481 , n17480 );
not ( n17482 , n17481 );
buf ( n17483 , n15963 );
buf ( n17484 , n17483 );
not ( n17485 , n17484 );
and ( n17486 , n17476 , n17479 , n17482 , n17485 );
buf ( n17487 , n15613 );
buf ( n17488 , n17487 );
not ( n17489 , n17488 );
nand ( n17490 , n17472 , n17486 , n17489 );
nor ( n17491 , n17463 , n17490 );
buf ( n17492 , n15509 );
or ( n17493 , n17491 , n17492 );
nand ( n17494 , n17491 , n17492 );
nand ( n17495 , n17493 , n17494 );
buf ( n17496 , n17495 );
nand ( n17497 , n17411 , n17496 );
not ( n17498 , n14869 );
nor ( n17499 , n16957 , n14900 );
nand ( n17500 , n17498 , n17499 );
buf ( n17501 , n17500 );
not ( n17502 , n17501 );
nand ( n17503 , n17502 , n15509 );
and ( n17504 , n13653 , n13555 );
nand ( n17505 , n17504 , n13677 );
not ( n17506 , n13592 );
nor ( n17507 , n17505 , n17506 );
nand ( n17508 , n17507 , n13574 );
not ( n17509 , n13631 );
nor ( n17510 , n17508 , n17509 );
nand ( n17511 , n17510 , n13617 );
not ( n17512 , n13476 );
nor ( n17513 , n17511 , n17512 );
nand ( n17514 , n17513 , n13458 );
not ( n17515 , n13714 );
nor ( n17516 , n17514 , n17515 );
nand ( n17517 , n17516 , n13699 );
not ( n17518 , n17517 );
nand ( n17519 , n17518 , n13526 );
not ( n17520 , n13490 );
nor ( n17521 , n17519 , n17520 );
nand ( n17522 , n17521 , n13770 );
not ( n17523 , n13745 );
nor ( n17524 , n17522 , n17523 );
nand ( n17525 , n17524 , n13856 );
not ( n17526 , n13896 );
nor ( n17527 , n17525 , n17526 );
nand ( n17528 , n17527 , n13910 );
not ( n17529 , n13827 );
nor ( n17530 , n17528 , n17529 );
and ( n17531 , n17530 , n13880 );
nand ( n17532 , n17531 , n13795 );
not ( n17533 , n13948 );
nor ( n17534 , n17532 , n17533 );
and ( n17535 , n17534 , n14002 );
not ( n17536 , n17534 );
not ( n17537 , n14001 );
and ( n17538 , n17536 , n17537 );
nor ( n17539 , n17535 , n17538 );
not ( n17540 , n14905 );
nand ( n17541 , n14900 , n17540 );
not ( n17542 , n14830 );
nor ( n17543 , n17541 , n17542 );
and ( n17544 , n16956 , n14827 , n17543 , n14839 );
buf ( n17545 , n17544 );
nand ( n17546 , n17539 , n17545 );
not ( n17547 , n14841 );
not ( n17548 , n14895 );
not ( n17549 , n14906 );
and ( n17550 , n17548 , n17549 );
not ( n17551 , n16957 );
not ( n17552 , n17541 );
and ( n17553 , n17551 , n17552 );
nor ( n17554 , n17553 , n16966 );
nor ( n17555 , n17550 , n17554 );
nor ( n17556 , n14894 , n14900 );
nor ( n17557 , n14906 , n17556 );
nand ( n17558 , n16958 , n17557 );
nand ( n17559 , n17558 , n14867 );
nand ( n17560 , n17547 , n17555 , n17559 );
not ( n17561 , n17560 );
not ( n17562 , n17561 );
nand ( n17563 , n17562 , n13990 );
nand ( n17564 , n17497 , n17503 , n17546 , n17563 );
nor ( n17565 , n17406 , n17564 );
and ( n17566 , n16971 , n17565 );
nand ( n17567 , n14910 , n17566 );
buf ( n17568 , n17567 );
buf ( n17569 , n17568 );
buf ( n17570 , RI210ccb90_257);
buf ( n17571 , n17570 );
not ( n17572 , n17571 );
buf ( n17573 , RI210c9b48_275);
not ( n17574 , n17573 );
not ( n17575 , n17574 );
not ( n17576 , n17575 );
buf ( n17577 , n17576 );
buf ( n17578 , n17577 );
not ( n17579 , n17578 );
or ( n17580 , n17572 , n17579 );
buf ( n17581 , n17571 );
not ( n17582 , n17581 );
not ( n17583 , n17582 );
buf ( n17584 , RI210cd658_251);
not ( n17585 , n17584 );
not ( n17586 , n17585 );
buf ( n17587 , n17586 );
buf ( n17588 , RI210cc140_262);
buf ( n17589 , n17588 );
buf ( n17590 , n17589 );
nor ( n17591 , n17587 , n17590 );
buf ( n17592 , RI210ca430_273);
buf ( n17593 , n17592 );
buf ( n17594 , n17593 );
buf ( n17595 , RI210c9ad0_276);
buf ( n17596 , n17595 );
buf ( n17597 , n17596 );
nor ( n17598 , n17594 , n17597 );
nand ( n17599 , n17591 , n17598 );
not ( n17600 , n17599 );
buf ( n17601 , RI210c91e8_278);
buf ( n17602 , n17601 );
buf ( n17603 , n17602 );
not ( n17604 , n17603 );
buf ( n17605 , RI210c9a58_277);
buf ( n17606 , n17605 );
buf ( n17607 , n17606 );
not ( n17608 , n17607 );
nand ( n17609 , n17604 , n17608 );
buf ( n17610 , RI210c2078_280);
buf ( n17611 , n17610 );
buf ( n17612 , n17611 );
not ( n17613 , n17612 );
buf ( n17614 , n17613 );
buf ( n17615 , RI210c9170_279);
buf ( n17616 , n17615 );
buf ( n17617 , n17616 );
not ( n17618 , n17617 );
buf ( n17619 , n17618 );
nand ( n17620 , n17614 , n17619 );
nor ( n17621 , n17609 , n17620 );
nand ( n17622 , n17600 , n17621 );
not ( n17623 , n17622 );
buf ( n17624 , RI210c07a0_282);
buf ( n17625 , n17624 );
buf ( n17626 , n17625 );
not ( n17627 , n17626 );
buf ( n17628 , RI210c0818_281);
buf ( n17629 , n17628 );
buf ( n17630 , n17629 );
not ( n17631 , n17630 );
nand ( n17632 , n17627 , n17631 );
buf ( n17633 , RI210cd568_253);
buf ( n17634 , n17633 );
buf ( n17635 , n17634 );
not ( n17636 , n17635 );
buf ( n17637 , n17636 );
buf ( n17638 , RI210cd5e0_252);
buf ( n17639 , n17638 );
buf ( n17640 , n17639 );
not ( n17641 , n17640 );
buf ( n17642 , n17641 );
nand ( n17643 , n17637 , n17642 );
nor ( n17644 , n17632 , n17643 );
buf ( n17645 , RI210ccc80_255);
buf ( n17646 , n17645 );
buf ( n17647 , n17646 );
not ( n17648 , n17647 );
buf ( n17649 , RI210cd4f0_254);
buf ( n17650 , n17649 );
buf ( n17651 , n17650 );
not ( n17652 , n17651 );
nand ( n17653 , n17648 , n17652 );
buf ( n17654 , RI210ccc08_256);
buf ( n17655 , n17654 );
buf ( n17656 , n17655 );
buf ( n17657 , n17656 );
nor ( n17658 , n17653 , n17657 );
and ( n17659 , n17644 , n17658 );
nand ( n17660 , n17623 , n17659 );
not ( n17661 , n17660 );
or ( n17662 , n17583 , n17661 );
nand ( n17663 , n17623 , n17659 );
or ( n17664 , n17663 , n17582 );
nand ( n17665 , n17662 , n17664 );
buf ( n17666 , n17665 );
not ( n17667 , n17575 );
not ( n17668 , n17667 );
nand ( n17669 , n17666 , n17668 );
nand ( n17670 , n17580 , n17669 );
not ( n17671 , n17670 );
not ( n17672 , n17578 );
not ( n17673 , n17672 );
nor ( n17674 , n17587 , n17590 );
nand ( n17675 , n17636 , n17613 );
nand ( n17676 , n17641 , n17618 );
nor ( n17677 , n17675 , n17676 );
nor ( n17678 , n17630 , n17607 );
nand ( n17679 , n17674 , n17677 , n17678 );
nor ( n17680 , n17581 , n17656 );
nor ( n17681 , n17651 , n17594 );
nor ( n17682 , n17626 , n17603 );
nor ( n17683 , n17647 , n17597 );
nand ( n17684 , n17680 , n17681 , n17682 , n17683 );
nor ( n17685 , n17679 , n17684 );
buf ( n17686 , n17685 );
buf ( n17687 , RI210cc2a8_259);
buf ( n17688 , n17687 );
buf ( n17689 , n17688 );
buf ( n17690 , RI210ccb18_258);
buf ( n17691 , n17690 );
buf ( n17692 , n17691 );
nor ( n17693 , n17689 , n17692 );
nand ( n17694 , n17686 , n17693 );
buf ( n17695 , RI210cc230_260);
buf ( n17696 , n17695 );
buf ( n17697 , n17696 );
not ( n17698 , n17697 );
xnor ( n17699 , n17694 , n17698 );
buf ( n17700 , n17699 );
not ( n17701 , n17700 );
or ( n17702 , n17673 , n17701 );
nand ( n17703 , n17578 , n17696 );
nand ( n17704 , n17702 , n17703 );
not ( n17705 , n17704 );
not ( n17706 , n17668 );
buf ( n17707 , n17689 );
not ( n17708 , n17707 );
not ( n17709 , n17692 );
nand ( n17710 , n17686 , n17709 );
not ( n17711 , n17710 );
not ( n17712 , n17711 );
or ( n17713 , n17708 , n17712 );
or ( n17714 , n17711 , n17707 );
nand ( n17715 , n17713 , n17714 );
buf ( n17716 , n17715 );
not ( n17717 , n17716 );
or ( n17718 , n17706 , n17717 );
nand ( n17719 , n17667 , n17688 );
nand ( n17720 , n17718 , n17719 );
not ( n17721 , n17720 );
not ( n17722 , n17691 );
not ( n17723 , n17578 );
or ( n17724 , n17722 , n17723 );
not ( n17725 , n17709 );
not ( n17726 , n17686 );
not ( n17727 , n17726 );
or ( n17728 , n17725 , n17727 );
or ( n17729 , n17726 , n17709 );
nand ( n17730 , n17728 , n17729 );
buf ( n17731 , n17730 );
not ( n17732 , n17667 );
nand ( n17733 , n17731 , n17732 );
nand ( n17734 , n17724 , n17733 );
not ( n17735 , n17734 );
and ( n17736 , n17671 , n17705 , n17721 , n17735 );
not ( n17737 , n17578 );
not ( n17738 , n17737 );
not ( n17739 , n17627 );
nand ( n17740 , n17600 , n17621 );
not ( n17741 , n17740 );
nand ( n17742 , n17741 , n17631 );
not ( n17743 , n17742 );
or ( n17744 , n17739 , n17743 );
nand ( n17745 , n17741 , n17631 );
or ( n17746 , n17745 , n17627 );
nand ( n17747 , n17744 , n17746 );
buf ( n17748 , n17747 );
not ( n17749 , n17748 );
or ( n17750 , n17738 , n17749 );
nand ( n17751 , n17578 , n17625 );
nand ( n17752 , n17750 , n17751 );
not ( n17753 , n17752 );
not ( n17754 , n17639 );
not ( n17755 , n17578 );
or ( n17756 , n17754 , n17755 );
not ( n17757 , n17667 );
not ( n17758 , n17642 );
not ( n17759 , n17632 );
nand ( n17760 , n17741 , n17759 );
not ( n17761 , n17760 );
or ( n17762 , n17758 , n17761 );
nand ( n17763 , n17623 , n17759 );
or ( n17764 , n17763 , n17642 );
nand ( n17765 , n17762 , n17764 );
buf ( n17766 , n17765 );
nand ( n17767 , n17757 , n17766 );
nand ( n17768 , n17756 , n17767 );
not ( n17769 , n17768 );
not ( n17770 , n17629 );
not ( n17771 , n17578 );
or ( n17772 , n17770 , n17771 );
not ( n17773 , n17578 );
and ( n17774 , n17631 , n17622 );
not ( n17775 , n17631 );
and ( n17776 , n17775 , n17623 );
or ( n17777 , n17774 , n17776 );
buf ( n17778 , n17777 );
nand ( n17779 , n17773 , n17778 );
nand ( n17780 , n17772 , n17779 );
buf ( n17781 , n17611 );
and ( n17782 , n17577 , n17781 );
not ( n17783 , n17577 );
not ( n17784 , n17614 );
not ( n17785 , n17619 );
nand ( n17786 , n17604 , n17608 );
nor ( n17787 , n17785 , n17786 );
nand ( n17788 , n17600 , n17787 );
not ( n17789 , n17788 );
or ( n17790 , n17784 , n17789 );
or ( n17791 , n17788 , n17614 );
nand ( n17792 , n17790 , n17791 );
buf ( n17793 , n17792 );
and ( n17794 , n17783 , n17793 );
or ( n17795 , n17782 , n17794 );
nor ( n17796 , n17780 , n17795 );
and ( n17797 , n17753 , n17769 , n17796 );
not ( n17798 , n17737 );
buf ( n17799 , RI210cb8d0_263);
buf ( n17800 , n17799 );
buf ( n17801 , n17800 );
buf ( n17802 , RI210cb858_264);
buf ( n17803 , n17802 );
buf ( n17804 , n17803 );
nor ( n17805 , n17801 , n17804 );
not ( n17806 , n17805 );
buf ( n17807 , RI210cc1b8_261);
buf ( n17808 , n17807 );
buf ( n17809 , n17808 );
buf ( n17810 , n17809 );
nor ( n17811 , n17810 , n17697 );
nand ( n17812 , n17811 , n17693 );
nor ( n17813 , n17806 , n17812 );
nand ( n17814 , n17686 , n17813 );
buf ( n17815 , RI210cb7e0_265);
buf ( n17816 , n17815 );
buf ( n17817 , n17816 );
not ( n17818 , n17817 );
xnor ( n17819 , n17814 , n17818 );
buf ( n17820 , n17819 );
not ( n17821 , n17820 );
or ( n17822 , n17798 , n17821 );
nand ( n17823 , n17578 , n17816 );
nand ( n17824 , n17822 , n17823 );
not ( n17825 , n17824 );
not ( n17826 , n17803 );
not ( n17827 , n17578 );
or ( n17828 , n17826 , n17827 );
buf ( n17829 , n17801 );
nor ( n17830 , n17812 , n17829 );
not ( n17831 , n17830 );
not ( n17832 , n17686 );
or ( n17833 , n17831 , n17832 );
not ( n17834 , n17804 );
nand ( n17835 , n17833 , n17834 );
not ( n17836 , n17684 );
buf ( n17837 , n17677 );
and ( n17838 , n17837 , n17693 );
and ( n17839 , n17678 , n17811 );
buf ( n17840 , n17587 );
buf ( n17841 , n17590 );
nor ( n17842 , n17840 , n17834 , n17829 , n17841 );
nand ( n17843 , n17836 , n17838 , n17839 , n17842 );
nand ( n17844 , n17835 , n17843 );
buf ( n17845 , n17844 );
nand ( n17846 , n17845 , n17672 );
nand ( n17847 , n17828 , n17846 );
not ( n17848 , n17737 );
not ( n17849 , n17829 );
nor ( n17850 , n17726 , n17812 );
not ( n17851 , n17850 );
or ( n17852 , n17849 , n17851 );
not ( n17853 , n17812 );
and ( n17854 , n17686 , n17853 );
or ( n17855 , n17854 , n17829 );
nand ( n17856 , n17852 , n17855 );
buf ( n17857 , n17856 );
not ( n17858 , n17857 );
or ( n17859 , n17848 , n17858 );
nand ( n17860 , n17667 , n17800 );
nand ( n17861 , n17859 , n17860 );
nor ( n17862 , n17847 , n17861 );
not ( n17863 , n17737 );
not ( n17864 , n17810 );
not ( n17865 , n17686 );
nand ( n17866 , n17693 , n17698 );
nor ( n17867 , n17865 , n17866 );
not ( n17868 , n17867 );
or ( n17869 , n17864 , n17868 );
not ( n17870 , n17686 );
nor ( n17871 , n17870 , n17866 );
or ( n17872 , n17871 , n17810 );
nand ( n17873 , n17869 , n17872 );
buf ( n17874 , n17873 );
not ( n17875 , n17874 );
or ( n17876 , n17863 , n17875 );
nand ( n17877 , n17578 , n17808 );
nand ( n17878 , n17876 , n17877 );
not ( n17879 , n17878 );
nand ( n17880 , n17825 , n17862 , n17879 );
not ( n17881 , n17880 );
nand ( n17882 , n17736 , n17797 , n17881 );
not ( n17883 , n17637 );
not ( n17884 , n17642 );
nor ( n17885 , n17884 , n17632 );
nand ( n17886 , n17741 , n17885 );
not ( n17887 , n17886 );
or ( n17888 , n17883 , n17887 );
nand ( n17889 , n17623 , n17885 );
or ( n17890 , n17889 , n17637 );
nand ( n17891 , n17888 , n17890 );
buf ( n17892 , n17891 );
nand ( n17893 , n17737 , n17892 );
nand ( n17894 , n17578 , n17634 );
nand ( n17895 , n17893 , n17894 );
not ( n17896 , n17895 );
not ( n17897 , n17655 );
not ( n17898 , n17667 );
or ( n17899 , n17897 , n17898 );
not ( n17900 , n17657 );
not ( n17901 , n17900 );
not ( n17902 , n17644 );
nor ( n17903 , n17902 , n17653 );
nand ( n17904 , n17741 , n17903 );
not ( n17905 , n17904 );
or ( n17906 , n17901 , n17905 );
nand ( n17907 , n17623 , n17903 );
or ( n17908 , n17907 , n17900 );
nand ( n17909 , n17906 , n17908 );
buf ( n17910 , n17909 );
nand ( n17911 , n17910 , n17668 );
nand ( n17912 , n17899 , n17911 );
not ( n17913 , n17912 );
not ( n17914 , n17646 );
not ( n17915 , n17578 );
or ( n17916 , n17914 , n17915 );
not ( n17917 , n17578 );
not ( n17918 , n17648 );
and ( n17919 , n17644 , n17652 );
nand ( n17920 , n17741 , n17919 );
not ( n17921 , n17920 );
or ( n17922 , n17918 , n17921 );
nand ( n17923 , n17741 , n17919 );
or ( n17924 , n17923 , n17648 );
nand ( n17925 , n17922 , n17924 );
buf ( n17926 , n17925 );
nand ( n17927 , n17917 , n17926 );
nand ( n17928 , n17916 , n17927 );
not ( n17929 , n17928 );
not ( n17930 , n17650 );
not ( n17931 , n17578 );
or ( n17932 , n17930 , n17931 );
not ( n17933 , n17652 );
nand ( n17934 , n17741 , n17644 );
not ( n17935 , n17934 );
or ( n17936 , n17933 , n17935 );
nand ( n17937 , n17623 , n17644 );
or ( n17938 , n17937 , n17652 );
nand ( n17939 , n17936 , n17938 );
buf ( n17940 , n17939 );
nand ( n17941 , n17940 , n17732 );
nand ( n17942 , n17932 , n17941 );
not ( n17943 , n17942 );
and ( n17944 , n17896 , n17913 , n17929 , n17943 );
not ( n17945 , n17737 );
buf ( n17946 , RI210cb768_266);
buf ( n17947 , n17946 );
buf ( n17948 , n17947 );
buf ( n17949 , n17948 );
not ( n17950 , n17949 );
nand ( n17951 , n17805 , n17818 );
not ( n17952 , n17951 );
nand ( n17953 , n17952 , n17853 );
nor ( n17954 , n17726 , n17953 );
not ( n17955 , n17954 );
or ( n17956 , n17950 , n17955 );
nor ( n17957 , n17812 , n17951 );
and ( n17958 , n17686 , n17957 );
or ( n17959 , n17958 , n17949 );
nand ( n17960 , n17956 , n17959 );
buf ( n17961 , n17960 );
not ( n17962 , n17961 );
or ( n17963 , n17945 , n17962 );
nand ( n17964 , n17578 , n17947 );
nand ( n17965 , n17963 , n17964 );
not ( n17966 , n17965 );
buf ( n17967 , RI210caef8_267);
buf ( n17968 , n17967 );
buf ( n17969 , n17968 );
and ( n17970 , n17667 , n17969 );
not ( n17971 , n17667 );
buf ( n17972 , n17968 );
buf ( n17973 , n17972 );
not ( n17974 , n17973 );
not ( n17975 , n17974 );
nor ( n17976 , n17804 , n17810 );
nor ( n17977 , n17817 , n17692 );
nor ( n17978 , n17689 , n17948 );
nor ( n17979 , n17697 , n17801 );
nand ( n17980 , n17976 , n17977 , n17978 , n17979 );
not ( n17981 , n17980 );
nand ( n17982 , n17686 , n17981 );
not ( n17983 , n17982 );
or ( n17984 , n17975 , n17983 );
nand ( n17985 , n17686 , n17981 );
or ( n17986 , n17985 , n17974 );
nand ( n17987 , n17984 , n17986 );
buf ( n17988 , n17987 );
and ( n17989 , n17971 , n17988 );
nor ( n17990 , n17970 , n17989 );
not ( n17991 , n17990 );
not ( n17992 , n17991 );
not ( n17993 , n17672 );
buf ( n17994 , RI210cae80_268);
buf ( n17995 , n17994 );
buf ( n17996 , n17995 );
buf ( n17997 , n17996 );
not ( n17998 , n17997 );
nor ( n17999 , n17801 , n17697 );
nor ( n18000 , n17809 , n17804 );
nand ( n18001 , n17977 , n17999 , n17978 , n18000 );
not ( n18002 , n18001 );
nand ( n18003 , n18002 , n17974 );
nor ( n18004 , n17865 , n18003 );
not ( n18005 , n18004 );
or ( n18006 , n17998 , n18005 );
nor ( n18007 , n17980 , n17973 );
and ( n18008 , n17686 , n18007 );
or ( n18009 , n18008 , n17997 );
nand ( n18010 , n18006 , n18009 );
buf ( n18011 , n18010 );
not ( n18012 , n18011 );
or ( n18013 , n17993 , n18012 );
nand ( n18014 , n17667 , n17995 );
nand ( n18015 , n18013 , n18014 );
not ( n18016 , n18015 );
not ( n18017 , n17668 );
buf ( n18018 , RI210cae08_269);
buf ( n18019 , n18018 );
buf ( n18020 , n18019 );
not ( n18021 , n18020 );
not ( n18022 , n18021 );
not ( n18023 , n18022 );
nor ( n18024 , n17996 , n17972 );
nand ( n18025 , n18002 , n18024 );
nor ( n18026 , n17865 , n18025 );
not ( n18027 , n18026 );
or ( n18028 , n18023 , n18027 );
not ( n18029 , n18024 );
nor ( n18030 , n18029 , n17980 );
and ( n18031 , n17686 , n18030 );
or ( n18032 , n18031 , n18022 );
nand ( n18033 , n18028 , n18032 );
buf ( n18034 , n18033 );
not ( n18035 , n18034 );
or ( n18036 , n18017 , n18035 );
nand ( n18037 , n17578 , n18019 );
nand ( n18038 , n18036 , n18037 );
not ( n18039 , n18038 );
nand ( n18040 , n17966 , n17992 , n18016 , n18039 );
not ( n18041 , n17575 );
buf ( n18042 , n17606 );
and ( n18043 , n18041 , n18042 );
not ( n18044 , n18041 );
not ( n18045 , n17608 );
not ( n18046 , n17599 );
or ( n18047 , n18045 , n18046 );
not ( n18048 , n17600 );
or ( n18049 , n18048 , n17608 );
nand ( n18050 , n18047 , n18049 );
buf ( n18051 , n18050 );
and ( n18052 , n18044 , n18051 );
nor ( n18053 , n18043 , n18052 );
not ( n18054 , n18053 );
buf ( n18055 , n17596 );
and ( n18056 , n17667 , n18055 );
not ( n18057 , n17667 );
not ( n18058 , n17597 );
not ( n18059 , n18058 );
not ( n18060 , n17674 );
not ( n18061 , n18060 );
not ( n18062 , n17594 );
nand ( n18063 , n18061 , n18062 );
not ( n18064 , n18063 );
or ( n18065 , n18059 , n18064 );
or ( n18066 , n18063 , n18058 );
nand ( n18067 , n18065 , n18066 );
buf ( n18068 , n18067 );
and ( n18069 , n18057 , n18068 );
nor ( n18070 , n18056 , n18069 );
not ( n18071 , n18070 );
nor ( n18072 , n18054 , n18071 );
buf ( n18073 , n17616 );
and ( n18074 , n17577 , n18073 );
not ( n18075 , n17577 );
not ( n18076 , n17619 );
not ( n18077 , n17786 );
nand ( n18078 , n18077 , n17600 );
not ( n18079 , n18078 );
or ( n18080 , n18076 , n18079 );
or ( n18081 , n18078 , n17619 );
nand ( n18082 , n18080 , n18081 );
buf ( n18083 , n18082 );
and ( n18084 , n18075 , n18083 );
nor ( n18085 , n18074 , n18084 );
not ( n18086 , n18085 );
not ( n18087 , n18086 );
not ( n18088 , n17604 );
nand ( n18089 , n17600 , n17608 );
not ( n18090 , n18089 );
or ( n18091 , n18088 , n18090 );
nand ( n18092 , n17600 , n17608 );
or ( n18093 , n18092 , n17604 );
nand ( n18094 , n18091 , n18093 );
buf ( n18095 , n18094 );
not ( n18096 , n18095 );
or ( n18097 , n18096 , n17667 );
buf ( n18098 , n17602 );
nand ( n18099 , n17577 , n18098 );
nand ( n18100 , n18097 , n18099 );
buf ( n18101 , n18100 );
not ( n18102 , n18101 );
not ( n18103 , n17575 );
not ( n18104 , n18062 );
not ( n18105 , n18060 );
or ( n18106 , n18104 , n18105 );
or ( n18107 , n18060 , n18062 );
nand ( n18108 , n18106 , n18107 );
buf ( n18109 , n18108 );
not ( n18110 , n18109 );
or ( n18111 , n18103 , n18110 );
buf ( n18112 , n17593 );
nand ( n18113 , n17576 , n18112 );
nand ( n18114 , n18111 , n18113 );
buf ( n18115 , n18114 );
not ( n18116 , n17575 );
not ( n18117 , n17841 );
not ( n18118 , n17840 );
not ( n18119 , n18118 );
or ( n18120 , n18117 , n18119 );
not ( n18121 , n17841 );
nand ( n18122 , n18121 , n17840 );
nand ( n18123 , n18120 , n18122 );
buf ( n18124 , n18123 );
not ( n18125 , n18124 );
or ( n18126 , n18116 , n18125 );
not ( n18127 , n17575 );
buf ( n18128 , n17589 );
nand ( n18129 , n18127 , n18128 );
nand ( n18130 , n18126 , n18129 );
buf ( n18131 , n18130 );
buf ( n18132 , n17586 );
not ( n18133 , n18132 );
not ( n18134 , n18133 );
buf ( n18135 , n18134 );
or ( n18136 , n18131 , n18135 );
nor ( n18137 , n18115 , n18136 );
nand ( n18138 , n18072 , n18087 , n18102 , n18137 );
nor ( n18139 , n18040 , n18138 );
nand ( n18140 , n17944 , n18139 );
or ( n18141 , n17882 , n18140 );
not ( n18142 , n17726 );
nor ( n18143 , n17972 , n17996 );
buf ( n18144 , RI210cad90_270);
buf ( n18145 , n18144 );
buf ( n18146 , n18145 );
nor ( n18147 , n18020 , n18146 );
nand ( n18148 , n18143 , n18147 );
not ( n18149 , n18148 );
buf ( n18150 , RI210ca4a8_272);
buf ( n18151 , n18150 );
buf ( n18152 , n18151 );
not ( n18153 , n18152 );
buf ( n18154 , RI210ca520_271);
buf ( n18155 , n18154 );
buf ( n18156 , n18155 );
not ( n18157 , n18156 );
nand ( n18158 , n18153 , n18157 );
buf ( n18159 , RI210ca3b8_274);
buf ( n18160 , n18159 );
buf ( n18161 , n18160 );
nor ( n18162 , n18158 , n18161 );
nand ( n18163 , n18149 , n18162 );
not ( n18164 , n17981 );
nor ( n18165 , n18163 , n18164 );
nand ( n18166 , n18142 , n18165 );
buf ( n18167 , n17575 );
buf ( n18168 , n18167 );
and ( n18169 , n18166 , n18168 );
not ( n18170 , n18166 );
not ( n18171 , n18168 );
and ( n18172 , n18170 , n18171 );
nor ( n18173 , n18169 , n18172 );
buf ( n18174 , n18173 );
nand ( n18175 , n18174 , n17668 );
not ( n18176 , n18175 );
nand ( n18177 , n18141 , n18176 );
buf ( n18178 , n18177 );
not ( n18179 , n18145 );
not ( n18180 , n17667 );
or ( n18181 , n18179 , n18180 );
nand ( n18182 , n18024 , n18021 );
nor ( n18183 , n18001 , n18182 );
nand ( n18184 , n17686 , n18183 );
not ( n18185 , n18146 );
xnor ( n18186 , n18184 , n18185 );
buf ( n18187 , n18186 );
nand ( n18188 , n18187 , n17672 );
nand ( n18189 , n18181 , n18188 );
not ( n18190 , n18189 );
or ( n18191 , n18178 , n18190 );
not ( n18192 , n18155 );
not ( n18193 , n17667 );
or ( n18194 , n18192 , n18193 );
and ( n18195 , n18061 , n17837 , n17678 );
nor ( n18196 , n17684 , n18148 );
nand ( n18197 , n18195 , n18196 , n18002 );
xnor ( n18198 , n18197 , n18157 );
buf ( n18199 , n18198 );
nand ( n18200 , n18199 , n17732 );
nand ( n18201 , n18194 , n18200 );
and ( n18202 , n18191 , n18201 );
not ( n18203 , n18191 );
not ( n18204 , n18201 );
and ( n18205 , n18203 , n18204 );
nor ( n18206 , n18202 , n18205 );
not ( n18207 , n18206 );
buf ( n18208 , n18207 );
buf ( n18209 , n18151 );
and ( n18210 , n17667 , n18209 );
not ( n18211 , n17667 );
not ( n18212 , n17726 );
nand ( n18213 , n18149 , n18157 );
nor ( n18214 , n18213 , n17980 );
nand ( n18215 , n18212 , n18214 );
and ( n18216 , n18215 , n18152 );
not ( n18217 , n18215 );
and ( n18218 , n18217 , n18153 );
nor ( n18219 , n18216 , n18218 );
buf ( n18220 , n18219 );
and ( n18221 , n18211 , n18220 );
nor ( n18222 , n18210 , n18221 );
not ( n18223 , n18222 );
not ( n18224 , n18223 );
nand ( n18225 , n17926 , n17672 );
nand ( n18226 , n17669 , n17911 , n18225 , n17733 );
not ( n18227 , n18226 );
nand ( n18228 , n17766 , n17732 );
nand ( n18229 , n17941 , n18228 );
and ( n18230 , n17577 , n17781 );
not ( n18231 , n17577 );
and ( n18232 , n18231 , n17793 );
nor ( n18233 , n18230 , n18232 );
nand ( n18234 , n18085 , n18233 );
not ( n18235 , n18234 );
not ( n18236 , n17578 );
nand ( n18237 , n18236 , n17778 );
nor ( n18238 , n18114 , n18130 );
nand ( n18239 , n18053 , n18070 , n18238 );
nor ( n18240 , n18239 , n18100 );
nand ( n18241 , n18235 , n18237 , n18240 );
nor ( n18242 , n18229 , n18241 );
nor ( n18243 , n17892 , n17748 );
nor ( n18244 , n17961 , n17820 );
nor ( n18245 , n17857 , n17700 );
and ( n18246 , n18243 , n17990 , n18244 , n18245 );
not ( n18247 , n18134 );
nand ( n18248 , n18247 , n18188 , n18200 , n17846 );
nor ( n18249 , n18011 , n17874 );
nor ( n18250 , n18034 , n17716 );
nand ( n18251 , n18249 , n18250 );
nor ( n18252 , n18248 , n18251 );
nand ( n18253 , n18227 , n18242 , n18246 , n18252 );
nand ( n18254 , n18253 , n18176 );
not ( n18255 , n18254 );
or ( n18256 , n18224 , n18255 );
or ( n18257 , n18254 , n18223 );
nand ( n18258 , n18256 , n18257 );
not ( n18259 , n18258 );
nor ( n18260 , n18222 , n18175 );
nand ( n18261 , n18253 , n18260 );
and ( n18262 , n17578 , n18160 );
not ( n18263 , n17578 );
not ( n18264 , n17726 );
not ( n18265 , n18158 );
nand ( n18266 , n18265 , n18149 );
nor ( n18267 , n18266 , n18164 );
nand ( n18268 , n18264 , n18267 );
xor ( n18269 , n18268 , n18161 );
buf ( n18270 , n18269 );
and ( n18271 , n18263 , n18270 );
nor ( n18272 , n18262 , n18271 );
not ( n18273 , n18272 );
and ( n18274 , n18261 , n18273 );
not ( n18275 , n18261 );
and ( n18276 , n18275 , n18272 );
nor ( n18277 , n18274 , n18276 );
buf ( n18278 , n18277 );
nor ( n18279 , n18259 , n18278 );
buf ( n18280 , n18279 );
buf ( n18281 , n18280 );
buf ( n18282 , RI210aeb90_395);
buf ( n18283 , n18282 );
nand ( n18284 , n18281 , n18283 );
nand ( n18285 , n18258 , n18278 );
buf ( n18286 , n18285 );
not ( n18287 , n18286 );
buf ( n18288 , RI210b43b0_360);
buf ( n18289 , n18288 );
nand ( n18290 , n18287 , n18289 );
not ( n18291 , n18258 );
nand ( n18292 , n18291 , n18278 );
buf ( n18293 , n18292 );
not ( n18294 , n18293 );
buf ( n18295 , RI210b7f38_335);
not ( n18296 , n18295 );
not ( n18297 , n18296 );
nand ( n18298 , n18294 , n18297 );
not ( n18299 , n18278 );
not ( n18300 , n18258 );
nand ( n18301 , n18299 , n18300 );
not ( n18302 , n18301 );
not ( n18303 , n18302 );
not ( n18304 , n18303 );
buf ( n18305 , RI210b2538_374);
buf ( n18306 , n18305 );
nand ( n18307 , n18304 , n18306 );
nand ( n18308 , n18284 , n18290 , n18298 , n18307 );
buf ( n18309 , n18308 );
and ( n18310 , n18208 , n18309 );
not ( n18311 , n18208 );
buf ( n18312 , RI210b5670_354);
not ( n18313 , n18312 );
not ( n18314 , n18313 );
not ( n18315 , n18314 );
not ( n18316 , n18294 );
or ( n18317 , n18315 , n18316 );
buf ( n18318 , RI21081aa0_439);
buf ( n18319 , n18318 );
nand ( n18320 , n18287 , n18319 );
nand ( n18321 , n18317 , n18320 );
not ( n18322 , n18321 );
buf ( n18323 , RI2107e878_458);
buf ( n18324 , n18323 );
and ( n18325 , n18281 , n18324 );
buf ( n18326 , RI210b07b0_386);
buf ( n18327 , n18326 );
and ( n18328 , n18304 , n18327 );
nor ( n18329 , n18325 , n18328 );
nand ( n18330 , n18322 , n18329 );
buf ( n18331 , n18330 );
buf ( n18332 , n18331 );
not ( n18333 , n18332 );
buf ( n18334 , RI210af478_393);
buf ( n18335 , n18334 );
nand ( n18336 , n18302 , n18335 );
not ( n18337 , n18286 );
buf ( n18338 , RI21080d80_445);
buf ( n18339 , n18338 );
nand ( n18340 , n18337 , n18339 );
nor ( n18341 , n18259 , n18278 );
not ( n18342 , n18341 );
not ( n18343 , n18342 );
buf ( n18344 , RI2107e698_462);
buf ( n18345 , n18344 );
nand ( n18346 , n18343 , n18345 );
nand ( n18347 , n18278 , n18300 );
not ( n18348 , n18347 );
buf ( n18349 , RI210834e0_427);
buf ( n18350 , n18349 );
nand ( n18351 , n18348 , n18350 );
nand ( n18352 , n18336 , n18340 , n18346 , n18351 );
buf ( n18353 , n18352 );
buf ( n18354 , n18353 );
buf ( n18355 , RI2107f3b8_456);
buf ( n18356 , n18355 );
not ( n18357 , n18356 );
not ( n18358 , n18302 );
or ( n18359 , n18357 , n18358 );
not ( n18360 , n18300 );
nand ( n18361 , n18278 , n18360 );
not ( n18362 , n18361 );
buf ( n18363 , RI21080f60_441);
buf ( n18364 , n18363 );
nand ( n18365 , n18362 , n18364 );
nand ( n18366 , n18359 , n18365 );
buf ( n18367 , RI210835d0_425);
buf ( n18368 , n18367 );
not ( n18369 , n18368 );
not ( n18370 , n18347 );
not ( n18371 , n18370 );
or ( n18372 , n18369 , n18371 );
buf ( n18373 , RI21084458_416);
buf ( n18374 , n18373 );
nand ( n18375 , n18341 , n18374 );
nand ( n18376 , n18372 , n18375 );
nor ( n18377 , n18366 , n18376 );
not ( n18378 , n18377 );
buf ( n18379 , n18378 );
buf ( n18380 , n18379 );
not ( n18381 , n18301 );
buf ( n18382 , RI210afdd8_390);
buf ( n18383 , n18382 );
nand ( n18384 , n18381 , n18383 );
not ( n18385 , n18361 );
buf ( n18386 , RI21080ee8_442);
buf ( n18387 , n18386 );
nand ( n18388 , n18385 , n18387 );
not ( n18389 , n18342 );
buf ( n18390 , RI2107e800_459);
buf ( n18391 , n18390 );
nand ( n18392 , n18389 , n18391 );
not ( n18393 , n18347 );
buf ( n18394 , RI210b4d10_357);
not ( n18395 , n18394 );
not ( n18396 , n18395 );
nand ( n18397 , n18393 , n18396 );
nand ( n18398 , n18384 , n18388 , n18392 , n18397 );
buf ( n18399 , n18398 );
buf ( n18400 , n18399 );
buf ( n18401 , RI210aec08_394);
buf ( n18402 , n18401 );
nand ( n18403 , n18302 , n18402 );
buf ( n18404 , RI210b25b0_373);
buf ( n18405 , n18404 );
nand ( n18406 , n18362 , n18405 );
buf ( n18407 , RI210843e0_417);
buf ( n18408 , n18407 );
nand ( n18409 , n18341 , n18408 );
buf ( n18410 , RI210b4428_359);
not ( n18411 , n18410 );
not ( n18412 , n18411 );
nand ( n18413 , n18370 , n18412 );
nand ( n18414 , n18403 , n18406 , n18409 , n18413 );
buf ( n18415 , n18414 );
buf ( n18416 , n18415 );
nand ( n18417 , n18354 , n18380 , n18400 , n18416 );
buf ( n18418 , n18417 );
buf ( n18419 , n18418 );
nand ( n18420 , n18299 , n18300 );
buf ( n18421 , n18420 );
buf ( n18422 , RI210b08a0_384);
not ( n18423 , n18422 );
not ( n18424 , n18423 );
not ( n18425 , n18424 );
nor ( n18426 , n18421 , n18425 );
buf ( n18427 , RI210b2f88_369);
not ( n18428 , n18427 );
not ( n18429 , n18428 );
not ( n18430 , n18429 );
nor ( n18431 , n18286 , n18430 );
nor ( n18432 , n18426 , n18431 );
buf ( n18433 , RI210b5760_352);
not ( n18434 , n18433 );
not ( n18435 , n18434 );
and ( n18436 , n18294 , n18435 );
not ( n18437 , n18280 );
buf ( n18438 , RI21084f98_414);
not ( n18439 , n18438 );
not ( n18440 , n18439 );
not ( n18441 , n18440 );
nor ( n18442 , n18437 , n18441 );
nor ( n18443 , n18436 , n18442 );
nand ( n18444 , n18432 , n18443 );
buf ( n18445 , n18444 );
buf ( n18446 , n18445 );
not ( n18447 , n18286 );
buf ( n18448 , RI210b2f10_370);
not ( n18449 , n18448 );
not ( n18450 , n18449 );
nand ( n18451 , n18447 , n18450 );
not ( n18452 , n18420 );
not ( n18453 , n18452 );
not ( n18454 , n18453 );
buf ( n18455 , RI210b0828_385);
not ( n18456 , n18455 );
not ( n18457 , n18456 );
nand ( n18458 , n18454 , n18457 );
buf ( n18459 , RI210b56e8_353);
not ( n18460 , n18459 );
not ( n18461 , n18460 );
nand ( n18462 , n18294 , n18461 );
nand ( n18463 , n18451 , n18458 , n18462 );
buf ( n18464 , n18463 );
buf ( n18465 , n18464 );
nand ( n18466 , n18446 , n18465 );
buf ( n18467 , n18466 );
buf ( n18468 , n18467 );
nor ( n18469 , n18419 , n18468 );
buf ( n18470 , n18469 );
buf ( n18471 , n18470 );
buf ( n18472 , RI210b3078_367);
not ( n18473 , n18472 );
not ( n18474 , n18473 );
and ( n18475 , n18447 , n18474 );
buf ( n18476 , RI210b1188_382);
not ( n18477 , n18476 );
not ( n18478 , n18477 );
not ( n18479 , n18478 );
nor ( n18480 , n18421 , n18479 );
nor ( n18481 , n18475 , n18480 );
buf ( n18482 , RI210b6048_350);
not ( n18483 , n18482 );
not ( n18484 , n18483 );
and ( n18485 , n18294 , n18484 );
buf ( n18486 , RI21085088_412);
buf ( n18487 , n18486 );
not ( n18488 , n18487 );
nor ( n18489 , n18437 , n18488 );
nor ( n18490 , n18485 , n18489 );
nand ( n18491 , n18481 , n18490 );
buf ( n18492 , n18491 );
buf ( n18493 , n18492 );
not ( n18494 , n18286 );
buf ( n18495 , RI210b3000_368);
not ( n18496 , n18495 );
not ( n18497 , n18496 );
not ( n18498 , n18497 );
not ( n18499 , n18498 );
and ( n18500 , n18494 , n18499 );
not ( n18501 , n18421 );
buf ( n18502 , RI210b0918_383);
not ( n18503 , n18502 );
not ( n18504 , n18503 );
and ( n18505 , n18501 , n18504 );
nor ( n18506 , n18500 , n18505 );
buf ( n18507 , RI21085010_413);
buf ( n18508 , n18507 );
not ( n18509 , n18508 );
nor ( n18510 , n18437 , n18509 );
buf ( n18511 , RI210b57d8_351);
not ( n18512 , n18511 );
not ( n18513 , n18512 );
not ( n18514 , n18513 );
nor ( n18515 , n18293 , n18514 );
nor ( n18516 , n18510 , n18515 );
nand ( n18517 , n18506 , n18516 );
buf ( n18518 , n18517 );
buf ( n18519 , n18518 );
nand ( n18520 , n18493 , n18519 );
buf ( n18521 , n18520 );
buf ( n18522 , n18521 );
not ( n18523 , n18280 );
buf ( n18524 , RI21085c40_409);
buf ( n18525 , n18524 );
not ( n18526 , n18525 );
nor ( n18527 , n18523 , n18526 );
buf ( n18528 , RI210b61b0_347);
not ( n18529 , n18528 );
not ( n18530 , n18529 );
not ( n18531 , n18530 );
nor ( n18532 , n18293 , n18531 );
nor ( n18533 , n18527 , n18532 );
not ( n18534 , n18452 );
buf ( n18535 , RI210b12f0_379);
buf ( n18536 , n18535 );
not ( n18537 , n18536 );
nor ( n18538 , n18534 , n18537 );
not ( n18539 , n18285 );
not ( n18540 , n18539 );
buf ( n18541 , RI210b39d8_364);
not ( n18542 , n18541 );
not ( n18543 , n18542 );
not ( n18544 , n18543 );
nor ( n18545 , n18540 , n18544 );
nor ( n18546 , n18538 , n18545 );
nand ( n18547 , n18533 , n18546 );
buf ( n18548 , n18547 );
buf ( n18549 , n18548 );
not ( n18550 , n18280 );
buf ( n18551 , RI21085cb8_408);
buf ( n18552 , n18551 );
not ( n18553 , n18552 );
nor ( n18554 , n18550 , n18553 );
buf ( n18555 , RI210b6a20_346);
not ( n18556 , n18555 );
not ( n18557 , n18556 );
not ( n18558 , n18557 );
nor ( n18559 , n18293 , n18558 );
nor ( n18560 , n18554 , n18559 );
buf ( n18561 , RI210b1b60_378);
not ( n18562 , n18561 );
not ( n18563 , n18562 );
not ( n18564 , n18563 );
nor ( n18565 , n18534 , n18564 );
buf ( n18566 , RI210b3a50_363);
not ( n18567 , n18566 );
not ( n18568 , n18567 );
not ( n18569 , n18568 );
nor ( n18570 , n18540 , n18569 );
nor ( n18571 , n18565 , n18570 );
nand ( n18572 , n18560 , n18571 );
buf ( n18573 , n18572 );
buf ( n18574 , n18573 );
nand ( n18575 , n18549 , n18574 );
buf ( n18576 , n18575 );
buf ( n18577 , n18576 );
nor ( n18578 , n18522 , n18577 );
buf ( n18579 , n18578 );
buf ( n18580 , n18579 );
nand ( n18581 , n18471 , n18580 );
buf ( n18582 , n18581 );
buf ( n18583 , n18582 );
not ( n18584 , n18293 );
buf ( n18585 , RI210b73f8_342);
not ( n18586 , n18585 );
not ( n18587 , n18586 );
not ( n18588 , n18587 );
not ( n18589 , n18588 );
and ( n18590 , n18584 , n18589 );
buf ( n18591 , RI21085e20_405);
buf ( n18592 , n18591 );
and ( n18593 , n18281 , n18592 );
nor ( n18594 , n18590 , n18593 );
buf ( n18595 , RI2107f520_453);
buf ( n18596 , n18595 );
not ( n18597 , n18596 );
nor ( n18598 , n18597 , n18534 );
buf ( n18599 , RI21081b90_437);
buf ( n18600 , n18599 );
not ( n18601 , n18600 );
nor ( n18602 , n18601 , n18540 );
nor ( n18603 , n18598 , n18602 );
nand ( n18604 , n18594 , n18603 );
buf ( n18605 , n18604 );
buf ( n18606 , n18605 );
not ( n18607 , n18293 );
buf ( n18608 , RI210836c0_423);
buf ( n18609 , n18608 );
not ( n18610 , n18609 );
not ( n18611 , n18610 );
and ( n18612 , n18607 , n18611 );
buf ( n18613 , RI21085e98_404);
buf ( n18614 , n18613 );
and ( n18615 , n18281 , n18614 );
nor ( n18616 , n18612 , n18615 );
not ( n18617 , n18539 );
not ( n18618 , n18617 );
buf ( n18619 , RI21081c08_436);
buf ( n18620 , n18619 );
not ( n18621 , n18620 );
not ( n18622 , n18621 );
and ( n18623 , n18618 , n18622 );
buf ( n18624 , RI210b1c50_376);
buf ( n18625 , n18624 );
and ( n18626 , n18501 , n18625 );
nor ( n18627 , n18623 , n18626 );
nand ( n18628 , n18616 , n18627 );
buf ( n18629 , n18628 );
buf ( n18630 , n18629 );
nand ( n18631 , n18606 , n18630 );
buf ( n18632 , n18631 );
buf ( n18633 , n18632 );
not ( n18634 , n18633 );
buf ( n18635 , n18634 );
buf ( n18636 , n18635 );
buf ( n18637 , RI210b1200_381);
buf ( n18638 , n18637 );
not ( n18639 , n18638 );
nor ( n18640 , n18421 , n18639 );
buf ( n18641 , RI210b38e8_366);
not ( n18642 , n18641 );
not ( n18643 , n18642 );
not ( n18644 , n18643 );
nor ( n18645 , n18286 , n18644 );
nor ( n18646 , n18640 , n18645 );
buf ( n18647 , RI210b60c0_349);
not ( n18648 , n18647 );
not ( n18649 , n18648 );
and ( n18650 , n18294 , n18649 );
not ( n18651 , n18280 );
buf ( n18652 , RI21085100_411);
buf ( n18653 , n18652 );
not ( n18654 , n18653 );
nor ( n18655 , n18651 , n18654 );
nor ( n18656 , n18650 , n18655 );
nand ( n18657 , n18646 , n18656 );
buf ( n18658 , n18657 );
buf ( n18659 , n18658 );
not ( n18660 , n18293 );
buf ( n18661 , RI210b6b10_344);
not ( n18662 , n18661 );
not ( n18663 , n18662 );
not ( n18664 , n18663 );
not ( n18665 , n18664 );
and ( n18666 , n18660 , n18665 );
buf ( n18667 , RI21085da8_406);
buf ( n18668 , n18667 );
and ( n18669 , n18281 , n18668 );
nor ( n18670 , n18666 , n18669 );
not ( n18671 , n18617 );
buf ( n18672 , RI210b4338_361);
not ( n18673 , n18672 );
not ( n18674 , n18673 );
not ( n18675 , n18674 );
not ( n18676 , n18675 );
and ( n18677 , n18671 , n18676 );
not ( n18678 , n18421 );
buf ( n18679 , RI2107f430_455);
buf ( n18680 , n18679 );
and ( n18681 , n18678 , n18680 );
nor ( n18682 , n18677 , n18681 );
nand ( n18683 , n18670 , n18682 );
buf ( n18684 , n18683 );
buf ( n18685 , n18684 );
and ( n18686 , n18659 , n18685 );
buf ( n18687 , n18686 );
buf ( n18688 , n18687 );
not ( n18689 , n18293 );
buf ( n18690 , RI210b7470_341);
not ( n18691 , n18690 );
not ( n18692 , n18691 );
not ( n18693 , n18692 );
not ( n18694 , n18693 );
and ( n18695 , n18689 , n18694 );
buf ( n18696 , RI21086a50_401);
buf ( n18697 , n18696 );
and ( n18698 , n18280 , n18697 );
nor ( n18699 , n18695 , n18698 );
buf ( n18700 , RI210800d8_450);
buf ( n18701 , n18700 );
not ( n18702 , n18701 );
nor ( n18703 , n18702 , n18534 );
buf ( n18704 , RI210827c0_433);
buf ( n18705 , n18704 );
not ( n18706 , n18705 );
nor ( n18707 , n18706 , n18540 );
nor ( n18708 , n18703 , n18707 );
nand ( n18709 , n18699 , n18708 );
buf ( n18710 , n18709 );
buf ( n18711 , n18710 );
not ( n18712 , n18293 );
buf ( n18713 , RI210b74e8_340);
not ( n18714 , n18713 );
not ( n18715 , n18714 );
not ( n18716 , n18715 );
not ( n18717 , n18716 );
and ( n18718 , n18712 , n18717 );
buf ( n18719 , RI21086ac8_400);
buf ( n18720 , n18719 );
and ( n18721 , n18280 , n18720 );
nor ( n18722 , n18718 , n18721 );
not ( n18723 , n18539 );
not ( n18724 , n18723 );
buf ( n18725 , RI21082838_432);
buf ( n18726 , n18725 );
not ( n18727 , n18726 );
not ( n18728 , n18727 );
and ( n18729 , n18724 , n18728 );
buf ( n18730 , RI21080150_449);
buf ( n18731 , n18730 );
and ( n18732 , n18501 , n18731 );
nor ( n18733 , n18729 , n18732 );
nand ( n18734 , n18722 , n18733 );
buf ( n18735 , n18734 );
buf ( n18736 , n18735 );
nand ( n18737 , n18711 , n18736 );
buf ( n18738 , n18737 );
buf ( n18739 , n18738 );
not ( n18740 , n18739 );
buf ( n18741 , n18740 );
buf ( n18742 , n18741 );
buf ( n18743 , RI210802b8_446);
buf ( n18744 , n18743 );
nand ( n18745 , n18452 , n18744 );
buf ( n18746 , RI210829a0_429);
buf ( n18747 , n18746 );
nand ( n18748 , n18539 , n18747 );
buf ( n18749 , RI21086e10_397);
buf ( n18750 , n18749 );
nand ( n18751 , n18280 , n18750 );
buf ( n18752 , RI210b7e48_337);
not ( n18753 , n18752 );
not ( n18754 , n18753 );
nand ( n18755 , n18370 , n18754 );
nand ( n18756 , n18745 , n18748 , n18751 , n18755 );
buf ( n18757 , n18756 );
buf ( n18758 , n18757 );
buf ( n18759 , RI210b1cc8_375);
buf ( n18760 , n18759 );
nand ( n18761 , n18302 , n18760 );
buf ( n18762 , RI21082a18_428);
buf ( n18763 , n18762 );
nand ( n18764 , n18362 , n18763 );
buf ( n18765 , RI210a63a0_396);
buf ( n18766 , n18765 );
nand ( n18767 , n18341 , n18766 );
buf ( n18768 , RI210b7ec0_336);
not ( n18769 , n18768 );
not ( n18770 , n18769 );
nand ( n18771 , n18370 , n18770 );
nand ( n18772 , n18761 , n18764 , n18767 , n18771 );
buf ( n18773 , n18772 );
buf ( n18774 , n18773 );
buf ( n18775 , n18774 );
nand ( n18776 , n18758 , n18775 );
buf ( n18777 , n18776 );
buf ( n18778 , n18777 );
not ( n18779 , n18778 );
buf ( n18780 , n18779 );
buf ( n18781 , n18780 );
nand ( n18782 , n18636 , n18688 , n18742 , n18781 );
buf ( n18783 , n18782 );
buf ( n18784 , n18783 );
nor ( n18785 , n18583 , n18784 );
buf ( n18786 , n18785 );
buf ( n18787 , n18786 );
buf ( n18788 , RI21085178_410);
buf ( n18789 , n18788 );
not ( n18790 , n18789 );
nor ( n18791 , n18437 , n18790 );
buf ( n18792 , RI210b6138_348);
not ( n18793 , n18792 );
not ( n18794 , n18793 );
not ( n18795 , n18794 );
nor ( n18796 , n18293 , n18795 );
nor ( n18797 , n18791 , n18796 );
buf ( n18798 , RI210b1278_380);
not ( n18799 , n18798 );
not ( n18800 , n18799 );
and ( n18801 , n18454 , n18800 );
buf ( n18802 , RI210b3960_365);
not ( n18803 , n18802 );
not ( n18804 , n18803 );
not ( n18805 , n18804 );
nor ( n18806 , n18286 , n18805 );
nor ( n18807 , n18801 , n18806 );
nand ( n18808 , n18797 , n18807 );
buf ( n18809 , n18808 );
buf ( n18810 , n18809 );
not ( n18811 , n18293 );
buf ( n18812 , RI210b6a98_345);
not ( n18813 , n18812 );
not ( n18814 , n18813 );
not ( n18815 , n18814 );
not ( n18816 , n18815 );
and ( n18817 , n18811 , n18816 );
buf ( n18818 , RI21085d30_407);
buf ( n18819 , n18818 );
and ( n18820 , n18281 , n18819 );
nor ( n18821 , n18817 , n18820 );
not ( n18822 , n18540 );
buf ( n18823 , RI210b42c0_362);
not ( n18824 , n18823 );
not ( n18825 , n18824 );
not ( n18826 , n18825 );
not ( n18827 , n18826 );
and ( n18828 , n18822 , n18827 );
buf ( n18829 , RI210b1bd8_377);
buf ( n18830 , n18829 );
and ( n18831 , n18678 , n18830 );
nor ( n18832 , n18828 , n18831 );
nand ( n18833 , n18821 , n18832 );
buf ( n18834 , n18833 );
buf ( n18835 , n18834 );
buf ( n18836 , RI210b26a0_371);
not ( n18837 , n18836 );
not ( n18838 , n18837 );
nand ( n18839 , n18447 , n18838 );
buf ( n18840 , RI210b4e00_355);
not ( n18841 , n18840 );
not ( n18842 , n18841 );
nand ( n18843 , n18294 , n18842 );
buf ( n18844 , RI210aff40_387);
not ( n18845 , n18844 );
not ( n18846 , n18845 );
nand ( n18847 , n18454 , n18846 );
nand ( n18848 , n18839 , n18843 , n18847 );
buf ( n18849 , n18848 );
buf ( n18850 , n18849 );
nand ( n18851 , n18810 , n18835 , n18850 );
buf ( n18852 , n18851 );
buf ( n18853 , n18852 );
not ( n18854 , n18853 );
not ( n18855 , n18293 );
buf ( n18856 , RI21083648_424);
buf ( n18857 , n18856 );
not ( n18858 , n18857 );
not ( n18859 , n18858 );
and ( n18860 , n18855 , n18859 );
buf ( n18861 , RI21084f20_415);
buf ( n18862 , n18861 );
and ( n18863 , n18280 , n18862 );
nor ( n18864 , n18860 , n18863 );
buf ( n18865 , RI210afe50_389);
buf ( n18866 , n18865 );
not ( n18867 , n18866 );
nor ( n18868 , n18867 , n18421 );
buf ( n18869 , RI21080fd8_440);
buf ( n18870 , n18869 );
not ( n18871 , n18870 );
nor ( n18872 , n18871 , n18286 );
nor ( n18873 , n18868 , n18872 );
nand ( n18874 , n18864 , n18873 );
buf ( n18875 , n18874 );
buf ( n18876 , n18875 );
buf ( n18877 , RI210af4f0_392);
buf ( n18878 , n18877 );
not ( n18879 , n18878 );
nor ( n18880 , n18879 , n18453 );
buf ( n18881 , RI21080df8_444);
buf ( n18882 , n18881 );
not ( n18883 , n18882 );
nor ( n18884 , n18540 , n18883 );
nor ( n18885 , n18880 , n18884 );
buf ( n18886 , RI2107e710_461);
buf ( n18887 , n18886 );
not ( n18888 , n18887 );
nor ( n18889 , n18550 , n18888 );
buf ( n18890 , RI21083558_426);
buf ( n18891 , n18890 );
not ( n18892 , n18891 );
nor ( n18893 , n18293 , n18892 );
nor ( n18894 , n18889 , n18893 );
nand ( n18895 , n18885 , n18894 );
buf ( n18896 , n18895 );
buf ( n18897 , n18896 );
buf ( n18898 , RI2107e788_460);
buf ( n18899 , n18898 );
not ( n18900 , n18899 );
nor ( n18901 , n18523 , n18900 );
buf ( n18902 , RI210b4c98_358);
buf ( n18903 , n18902 );
not ( n18904 , n18903 );
nor ( n18905 , n18293 , n18904 );
nor ( n18906 , n18901 , n18905 );
buf ( n18907 , RI210af568_391);
buf ( n18908 , n18907 );
not ( n18909 , n18908 );
nor ( n18910 , n18909 , n18421 );
buf ( n18911 , RI21080e70_443);
buf ( n18912 , n18911 );
not ( n18913 , n18912 );
nor ( n18914 , n18913 , n18723 );
nor ( n18915 , n18910 , n18914 );
nand ( n18916 , n18906 , n18915 );
buf ( n18917 , n18916 );
buf ( n18918 , n18917 );
buf ( n18919 , n18281 );
buf ( n18920 , n18919 );
buf ( n18921 , n18920 );
nand ( n18922 , n18876 , n18897 , n18918 , n18921 );
buf ( n18923 , n18922 );
buf ( n18924 , n18923 );
not ( n18925 , n18924 );
buf ( n18926 , n18925 );
buf ( n18927 , n18926 );
not ( n18928 , n18293 );
buf ( n18929 , RI21083738_422);
buf ( n18930 , n18929 );
not ( n18931 , n18930 );
not ( n18932 , n18931 );
and ( n18933 , n18928 , n18932 );
buf ( n18934 , RI21086960_403);
buf ( n18935 , n18934 );
and ( n18936 , n18281 , n18935 );
nor ( n18937 , n18933 , n18936 );
not ( n18938 , n18617 );
buf ( n18939 , RI21081c80_435);
buf ( n18940 , n18939 );
not ( n18941 , n18940 );
not ( n18942 , n18941 );
and ( n18943 , n18938 , n18942 );
buf ( n18944 , RI2107f598_452);
buf ( n18945 , n18944 );
and ( n18946 , n18678 , n18945 );
nor ( n18947 , n18943 , n18946 );
nand ( n18948 , n18937 , n18947 );
buf ( n18949 , n18948 );
buf ( n18950 , n18949 );
not ( n18951 , n18293 );
buf ( n18952 , RI21084200_421);
buf ( n18953 , n18952 );
not ( n18954 , n18953 );
not ( n18955 , n18954 );
and ( n18956 , n18951 , n18955 );
buf ( n18957 , RI210869d8_402);
buf ( n18958 , n18957 );
and ( n18959 , n18281 , n18958 );
nor ( n18960 , n18956 , n18959 );
not ( n18961 , n18617 );
buf ( n18962 , RI21081cf8_434);
buf ( n18963 , n18962 );
not ( n18964 , n18963 );
not ( n18965 , n18964 );
and ( n18966 , n18961 , n18965 );
buf ( n18967 , RI21080060_451);
buf ( n18968 , n18967 );
and ( n18969 , n18678 , n18968 );
nor ( n18970 , n18966 , n18969 );
nand ( n18971 , n18960 , n18970 );
buf ( n18972 , n18971 );
buf ( n18973 , n18972 );
nand ( n18974 , n18950 , n18973 );
buf ( n18975 , n18974 );
buf ( n18976 , n18975 );
not ( n18977 , n18976 );
buf ( n18978 , n18977 );
buf ( n18979 , n18978 );
not ( n18980 , n18540 );
buf ( n18981 , RI210828b0_431);
buf ( n18982 , n18981 );
not ( n18983 , n18982 );
not ( n18984 , n18983 );
and ( n18985 , n18980 , n18984 );
buf ( n18986 , RI210801c8_448);
buf ( n18987 , n18986 );
and ( n18988 , n18501 , n18987 );
nor ( n18989 , n18985 , n18988 );
buf ( n18990 , RI21086b40_399);
buf ( n18991 , n18990 );
not ( n18992 , n18991 );
nor ( n18993 , n18550 , n18992 );
buf ( n18994 , RI210b7560_339);
buf ( n18995 , n18994 );
buf ( n18996 , n18995 );
not ( n18997 , n18996 );
nor ( n18998 , n18293 , n18997 );
nor ( n18999 , n18993 , n18998 );
nand ( n19000 , n18989 , n18999 );
buf ( n19001 , n19000 );
buf ( n19002 , n19001 );
not ( n19003 , n18540 );
buf ( n19004 , RI21082928_430);
buf ( n19005 , n19004 );
not ( n19006 , n19005 );
not ( n19007 , n19006 );
and ( n19008 , n19003 , n19007 );
buf ( n19009 , RI21080240_447);
buf ( n19010 , n19009 );
and ( n19011 , n18501 , n19010 );
nor ( n19012 , n19008 , n19011 );
not ( n19013 , n18293 );
buf ( n19014 , RI210b7dd0_338);
buf ( n19015 , n19014 );
not ( n19016 , n19015 );
not ( n19017 , n19016 );
and ( n19018 , n19013 , n19017 );
buf ( n19019 , RI21086bb8_398);
buf ( n19020 , n19019 );
and ( n19021 , n18280 , n19020 );
nor ( n19022 , n19018 , n19021 );
nand ( n19023 , n19012 , n19022 );
buf ( n19024 , n19023 );
buf ( n19025 , n19024 );
nand ( n19026 , n19002 , n19025 );
buf ( n19027 , n19026 );
buf ( n19028 , n19027 );
not ( n19029 , n19028 );
buf ( n19030 , n19029 );
buf ( n19031 , n19030 );
nand ( n19032 , n18854 , n18927 , n18979 , n19031 );
buf ( n19033 , n19032 );
buf ( n19034 , n19033 );
not ( n19035 , n19034 );
buf ( n19036 , n19035 );
buf ( n19037 , n19036 );
nand ( n19038 , n18787 , n19037 );
buf ( n19039 , n19038 );
buf ( n19040 , n19039 );
buf ( n19041 , RI210b2628_372);
buf ( n19042 , n19041 );
not ( n19043 , n19042 );
not ( n19044 , n18447 );
or ( n19045 , n19043 , n19044 );
buf ( n19046 , RI210afec8_388);
buf ( n19047 , n19046 );
and ( n19048 , n18501 , n19047 );
buf ( n19049 , RI210b4d88_356);
buf ( n19050 , n19049 );
not ( n19051 , n19050 );
nor ( n19052 , n19051 , n18293 );
nor ( n19053 , n19048 , n19052 );
nand ( n19054 , n19045 , n19053 );
buf ( n19055 , n19054 );
buf ( n19056 , n19055 );
not ( n19057 , n19056 );
buf ( n19058 , n19057 );
buf ( n19059 , n19058 );
and ( n19060 , n19040 , n19059 );
not ( n19061 , n19040 );
buf ( n19062 , n19055 );
and ( n19063 , n19061 , n19062 );
nor ( n19064 , n19060 , n19063 );
buf ( n19065 , n19064 );
buf ( n19066 , n19065 );
and ( n19067 , n19066 , n18309 );
buf ( n19068 , n19067 );
buf ( n19069 , n19068 );
buf ( n19070 , RI210b6b88_343);
not ( n19071 , n19070 );
not ( n19072 , n19071 );
not ( n19073 , n19072 );
not ( n19074 , n18294 );
or ( n19075 , n19073 , n19074 );
buf ( n19076 , RI21081b18_438);
buf ( n19077 , n19076 );
nand ( n19078 , n18287 , n19077 );
nand ( n19079 , n19075 , n19078 );
not ( n19080 , n19079 );
not ( n19081 , n18303 );
buf ( n19082 , RI2107f4a8_454);
buf ( n19083 , n19082 );
not ( n19084 , n19083 );
not ( n19085 , n19084 );
and ( n19086 , n19081 , n19085 );
buf ( n19087 , RI2107f340_457);
buf ( n19088 , n19087 );
and ( n19089 , n18281 , n19088 );
nor ( n19090 , n19086 , n19089 );
nand ( n19091 , n19080 , n19090 );
buf ( n19092 , n19091 );
buf ( n19093 , n19092 );
buf ( n19094 , n19093 );
nand ( n19095 , n19069 , n19094 );
not ( n19096 , n19095 );
or ( n19097 , n18333 , n19096 );
or ( n19098 , n19095 , n18332 );
nand ( n19099 , n19097 , n19098 );
buf ( n19100 , n19099 );
and ( n19101 , n18311 , n19100 );
nor ( n19102 , n18310 , n19101 );
not ( n19103 , n17966 );
not ( n19104 , n19103 );
not ( n19105 , n18176 );
or ( n19106 , n19104 , n19105 );
nor ( n19107 , n17880 , n18138 );
nand ( n19108 , n19107 , n17944 , n17797 , n17736 );
nand ( n19109 , n19108 , n18176 );
nand ( n19110 , n19106 , n19109 );
buf ( n19111 , n17991 );
nand ( n19112 , n19110 , n19111 );
not ( n19113 , n19112 );
buf ( n19114 , n18015 );
and ( n19115 , n19113 , n19114 );
not ( n19116 , n19113 );
not ( n19117 , n19114 );
and ( n19118 , n19116 , n19117 );
nor ( n19119 , n19115 , n19118 );
and ( n19120 , n19110 , n19111 );
not ( n19121 , n19110 );
not ( n19122 , n19111 );
and ( n19123 , n19121 , n19122 );
nor ( n19124 , n19120 , n19123 );
and ( n19125 , n19119 , n19124 );
buf ( n19126 , n18038 );
not ( n19127 , n19126 );
nand ( n19128 , n19113 , n19114 );
not ( n19129 , n19128 );
or ( n19130 , n19127 , n19129 );
or ( n19131 , n19128 , n19126 );
nand ( n19132 , n19130 , n19131 );
and ( n19133 , n19125 , n19132 );
nor ( n19134 , n19133 , n275557 );
not ( n19135 , n19103 );
buf ( n19136 , n19109 );
not ( n19137 , n19136 );
or ( n19138 , n19135 , n19137 );
or ( n19139 , n19136 , n19103 );
nand ( n19140 , n19138 , n19139 );
not ( n19141 , n19140 );
nand ( n19142 , n19134 , n19141 );
not ( n19143 , n19142 );
buf ( n19144 , n19132 );
buf ( n19145 , RI210cdec8_250);
not ( n19146 , n19145 );
not ( n19147 , n19146 );
not ( n19148 , n19124 );
or ( n19149 , n19147 , n19148 );
not ( n19150 , n19124 );
buf ( n19151 , n19145 );
nand ( n19152 , n19150 , n19151 );
nand ( n19153 , n19149 , n19152 );
not ( n19154 , n19119 );
and ( n19155 , n19153 , n19154 );
buf ( n19156 , RI210bcdf8_303);
buf ( n19157 , n19156 );
nor ( n19158 , n19155 , n19157 );
and ( n19159 , n19144 , n19158 );
not ( n19160 , n19144 );
and ( n19161 , n19160 , n19154 );
nor ( n19162 , n19159 , n19161 );
nand ( n19163 , n19143 , n19162 );
not ( n19164 , n19163 );
or ( n19165 , n19152 , n19119 );
buf ( n19166 , RI210bd668_302);
not ( n19167 , n19166 );
nand ( n19168 , n19165 , n19167 );
nand ( n19169 , n19168 , n19144 );
not ( n19170 , n19151 );
not ( n19171 , n19144 );
or ( n19172 , n19170 , n19171 );
nand ( n19173 , n19172 , n19124 );
nand ( n19174 , n19169 , n19173 );
not ( n19175 , n19174 );
nand ( n19176 , n19164 , n19175 );
not ( n19177 , n19176 );
and ( n19178 , n18087 , n18102 , n18072 );
and ( n19179 , n19178 , n18137 );
nand ( n19180 , n17944 , n17736 , n17797 , n19179 );
nand ( n19181 , n19180 , n18176 );
buf ( n19182 , n17878 );
not ( n19183 , n19182 );
nor ( n19184 , n19181 , n19183 );
buf ( n19185 , n17861 );
nand ( n19186 , n19184 , n19185 );
buf ( n19187 , n17847 );
not ( n19188 , n19187 );
nor ( n19189 , n19186 , n19188 );
not ( n19190 , n19189 );
not ( n19191 , n17824 );
not ( n19192 , n19191 );
and ( n19193 , n19190 , n19192 );
and ( n19194 , n19189 , n19191 );
nor ( n19195 , n19193 , n19194 );
and ( n19196 , n19186 , n19187 );
not ( n19197 , n19186 );
and ( n19198 , n19197 , n19188 );
nor ( n19199 , n19196 , n19198 );
nor ( n19200 , n19195 , n19199 );
not ( n19201 , n19200 );
and ( n19202 , n19184 , n19185 );
not ( n19203 , n19184 );
not ( n19204 , n19185 );
and ( n19205 , n19203 , n19204 );
nor ( n19206 , n19202 , n19205 );
not ( n19207 , n19206 );
not ( n19208 , n19181 );
not ( n19209 , n19182 );
and ( n19210 , n19208 , n19209 );
and ( n19211 , n19181 , n19182 );
nor ( n19212 , n19210 , n19211 );
nand ( n19213 , n19207 , n19212 );
nor ( n19214 , n19201 , n19213 );
and ( n19215 , n19177 , n19214 );
not ( n19216 , n19215 );
or ( n19217 , n19102 , n19216 );
and ( n19218 , n19195 , n19206 );
and ( n19219 , n19218 , n19199 );
nand ( n19220 , n19177 , n19219 );
not ( n19221 , n19220 );
not ( n19222 , n18131 );
or ( n19223 , n17882 , n18140 );
nand ( n19224 , n19223 , n18176 );
not ( n19225 , n19224 );
not ( n19226 , n18189 );
and ( n19227 , n19225 , n19226 );
and ( n19228 , n18177 , n18189 );
nor ( n19229 , n19227 , n19228 );
and ( n19230 , n18201 , n18190 );
not ( n19231 , n18201 );
and ( n19232 , n19231 , n18189 );
nor ( n19233 , n19230 , n19232 );
and ( n19234 , n19229 , n19233 );
buf ( n19235 , n19234 );
not ( n19236 , n19235 );
or ( n19237 , n19222 , n19236 );
nor ( n19238 , n19224 , n18189 );
not ( n19239 , n19238 );
nand ( n19240 , n18177 , n18189 );
nand ( n19241 , n19239 , n19240 , n19233 );
buf ( n19242 , n19241 );
buf ( n19243 , n9436 );
buf ( n19244 , n19243 );
buf ( n19245 , n19244 );
buf ( n19246 , n11050 );
buf ( n19247 , n19246 );
and ( n19248 , n19245 , n19247 );
buf ( n19249 , n19248 );
buf ( n19250 , n19249 );
not ( n19251 , n19250 );
buf ( n19252 , n9445 );
buf ( n19253 , n19252 );
buf ( n19254 , n19253 );
buf ( n19255 , n10971 );
buf ( n19256 , n19255 );
or ( n19257 , n19254 , n19256 );
buf ( n19258 , n19257 );
buf ( n19259 , n19258 );
buf ( n19260 , n19253 );
buf ( n19261 , n19255 );
nand ( n19262 , n19260 , n19261 );
buf ( n19263 , n19262 );
buf ( n19264 , n19263 );
nand ( n19265 , n19259 , n19264 );
buf ( n19266 , n19265 );
buf ( n19267 , n19266 );
not ( n19268 , n19267 );
or ( n19269 , n19251 , n19268 );
buf ( n19270 , n19266 );
buf ( n19271 , n19249 );
or ( n19272 , n19270 , n19271 );
nand ( n19273 , n19269 , n19272 );
buf ( n19274 , n19273 );
buf ( n19275 , n19274 );
and ( n19276 , n277817 , n19275 );
not ( n19277 , n277817 );
buf ( n19278 , n19252 );
and ( n19279 , n19277 , n19278 );
or ( n19280 , n19276 , n19279 );
nand ( n19281 , n19242 , n19280 );
nand ( n19282 , n19237 , n19281 );
buf ( n19283 , n19282 );
buf ( n19284 , n19283 );
buf ( n19285 , n19284 );
buf ( n19286 , n19285 );
nand ( n19287 , n19221 , n19286 );
nand ( n19288 , n19195 , n19199 );
or ( n19289 , n19288 , n19213 );
not ( n19290 , n19289 );
nand ( n19291 , n19177 , n19290 );
not ( n19292 , n19291 );
buf ( n19293 , n19283 );
not ( n19294 , n18135 );
not ( n19295 , n19235 );
or ( n19296 , n19294 , n19295 );
buf ( n19297 , n19244 );
buf ( n19298 , n19246 );
xor ( n19299 , n19297 , n19298 );
buf ( n19300 , n19299 );
buf ( n19301 , n19300 );
and ( n19302 , n277350 , n19301 );
not ( n19303 , n277350 );
and ( n19304 , n19303 , n19243 );
or ( n19305 , n19302 , n19304 );
nand ( n19306 , n19242 , n19305 );
nand ( n19307 , n19296 , n19306 );
buf ( n19308 , n19307 );
buf ( n19309 , n19308 );
xor ( n19310 , n19293 , n19309 );
buf ( n19311 , n19310 );
not ( n19312 , n19311 );
not ( n19313 , n19312 );
and ( n19314 , n19292 , n19313 );
or ( n19315 , n19206 , n19212 );
nor ( n19316 , n19288 , n19315 );
nand ( n19317 , n19143 , n19316 );
not ( n19318 , n19317 );
and ( n19319 , n19318 , n19088 );
nor ( n19320 , n19314 , n19319 );
buf ( n19321 , n18309 );
not ( n19322 , n19321 );
buf ( n19323 , n19307 );
not ( n19324 , n19323 );
nand ( n19325 , n19322 , n19324 );
not ( n19326 , n19325 );
not ( n19327 , n19326 );
buf ( n19328 , n19282 );
not ( n19329 , n19328 );
not ( n19330 , n19329 );
buf ( n19331 , n19092 );
not ( n19332 , n19331 );
not ( n19333 , n19332 );
or ( n19334 , n19330 , n19333 );
nand ( n19335 , n19331 , n19328 );
nand ( n19336 , n19334 , n19335 );
nor ( n19337 , n19336 , n19321 );
buf ( n19338 , n19337 );
not ( n19339 , n19338 );
nand ( n19340 , n19336 , n19321 );
buf ( n19341 , n19340 );
nand ( n19342 , n19339 , n19341 );
not ( n19343 , n19342 );
or ( n19344 , n19327 , n19343 );
or ( n19345 , n19342 , n19326 );
nand ( n19346 , n19344 , n19345 );
buf ( n19347 , n19346 );
nor ( n19348 , n19195 , n19212 );
nor ( n19349 , n19218 , n19348 );
not ( n19350 , n19200 );
nand ( n19351 , n19350 , n19288 );
nor ( n19352 , n19349 , n19351 );
nand ( n19353 , n19177 , n19352 );
not ( n19354 , n19353 );
nand ( n19355 , n19347 , n19354 );
not ( n19356 , n19349 );
nor ( n19357 , n19356 , n19351 );
buf ( n19358 , n19357 );
nand ( n19359 , n19177 , n19358 );
not ( n19360 , n19359 );
buf ( n19361 , n18309 );
buf ( n19362 , n19307 );
nand ( n19363 , n19361 , n19362 );
not ( n19364 , n19363 );
buf ( n19365 , n19282 );
buf ( n19366 , n19092 );
xor ( n19367 , n19365 , n19366 );
not ( n19368 , n19367 );
or ( n19369 , n19364 , n19368 );
or ( n19370 , n19367 , n19363 );
nand ( n19371 , n19369 , n19370 );
buf ( n19372 , n19371 );
nand ( n19373 , n19360 , n19372 );
nand ( n19374 , n19287 , n19320 , n19355 , n19373 );
not ( n19375 , n19083 );
not ( n19376 , n19316 );
not ( n19377 , n19162 );
nand ( n19378 , n19376 , n19377 );
nand ( n19379 , n19200 , n19206 );
not ( n19380 , n19199 );
nand ( n19381 , n19348 , n19380 );
nand ( n19382 , n19143 , n19378 , n19379 , n19381 );
or ( n19383 , n19195 , n19207 );
nand ( n19384 , n19383 , n19315 );
and ( n19385 , n19351 , n19384 );
nor ( n19386 , n19385 , n19175 );
or ( n19387 , n19382 , n19386 );
not ( n19388 , n19387 );
nor ( n19389 , n19375 , n19388 );
nor ( n19390 , n19374 , n19389 );
nand ( n19391 , n19217 , n19390 );
buf ( n19392 , n19391 );
buf ( n19393 , n19392 );
buf ( n19394 , n18923 );
not ( n19395 , n19394 );
buf ( n19396 , n18399 );
buf ( n19397 , n19396 );
buf ( n19398 , n18379 );
nand ( n19399 , n19397 , n19398 );
buf ( n19400 , n19399 );
buf ( n19401 , n19400 );
not ( n19402 , n19401 );
buf ( n19403 , n19402 );
buf ( n19404 , n19403 );
nand ( n19405 , n19395 , n19404 );
buf ( n19406 , n19405 );
buf ( n19407 , n19406 );
not ( n19408 , n19407 );
buf ( n19409 , n19408 );
buf ( n19410 , n19409 );
buf ( n19411 , n18353 );
buf ( n19412 , n19411 );
buf ( n19413 , n19412 );
and ( n19414 , n19410 , n19413 );
buf ( n19415 , n19414 );
buf ( n19416 , n19415 );
buf ( n19417 , n18415 );
buf ( n19418 , n19417 );
and ( n19419 , n19416 , n19418 );
not ( n19420 , n19416 );
buf ( n19421 , n19417 );
not ( n19422 , n19421 );
buf ( n19423 , n19422 );
buf ( n19424 , n19423 );
and ( n19425 , n19420 , n19424 );
nor ( n19426 , n19419 , n19425 );
buf ( n19427 , n19426 );
buf ( n19428 , n19427 );
buf ( n19429 , n19428 );
and ( n19430 , n18208 , n19429 );
not ( n19431 , n18208 );
buf ( n19432 , n18757 );
buf ( n19433 , n19432 );
not ( n19434 , n19433 );
buf ( n19435 , n19409 );
buf ( n19436 , n19417 );
buf ( n19437 , n19411 );
nand ( n19438 , n19436 , n19437 );
buf ( n19439 , n19438 );
buf ( n19440 , n19439 );
buf ( n19441 , n18774 );
buf ( n19442 , n19441 );
not ( n19443 , n19442 );
buf ( n19444 , n19443 );
buf ( n19445 , n19444 );
nor ( n19446 , n19440 , n19445 );
buf ( n19447 , n19446 );
buf ( n19448 , n19447 );
nand ( n19449 , n19435 , n19448 );
buf ( n19450 , n19449 );
buf ( n19451 , n19450 );
not ( n19452 , n19451 );
or ( n19453 , n19434 , n19452 );
buf ( n19454 , n18926 );
buf ( n19455 , n19400 );
not ( n19456 , n19455 );
buf ( n19457 , n19456 );
buf ( n19458 , n19457 );
nand ( n19459 , n19454 , n19458 );
buf ( n19460 , n19459 );
buf ( n19461 , n19460 );
not ( n19462 , n19461 );
buf ( n19463 , n19462 );
buf ( n19464 , n19463 );
buf ( n19465 , n19447 );
nand ( n19466 , n19464 , n19465 );
buf ( n19467 , n19466 );
buf ( n19468 , n19467 );
buf ( n19469 , n19432 );
or ( n19470 , n19468 , n19469 );
nand ( n19471 , n19453 , n19470 );
buf ( n19472 , n19471 );
buf ( n19473 , n19472 );
buf ( n19474 , n19473 );
buf ( n19475 , n19474 );
not ( n19476 , n19475 );
buf ( n19477 , n19428 );
buf ( n19478 , n19477 );
not ( n19479 , n19478 );
buf ( n19480 , n19412 );
not ( n19481 , n19480 );
buf ( n19482 , n19409 );
not ( n19483 , n19482 );
buf ( n19484 , n19483 );
buf ( n19485 , n19484 );
not ( n19486 , n19485 );
or ( n19487 , n19481 , n19486 );
buf ( n19488 , n19412 );
not ( n19489 , n19488 );
buf ( n19490 , n19409 );
nand ( n19491 , n19489 , n19490 );
buf ( n19492 , n19491 );
buf ( n19493 , n19492 );
nand ( n19494 , n19487 , n19493 );
buf ( n19495 , n19494 );
buf ( n19496 , n19495 );
buf ( n19497 , n19496 );
buf ( n19498 , n18379 );
not ( n19499 , n19498 );
buf ( n19500 , n18875 );
buf ( n19501 , n19500 );
buf ( n19502 , n18920 );
nand ( n19503 , n19501 , n19502 );
buf ( n19504 , n19503 );
buf ( n19505 , n19504 );
not ( n19506 , n19505 );
or ( n19507 , n19499 , n19506 );
buf ( n19508 , n18379 );
not ( n19509 , n19508 );
buf ( n19510 , n18875 );
buf ( n19511 , n18920 );
nand ( n19512 , n19510 , n19511 );
buf ( n19513 , n19512 );
buf ( n19514 , n19513 );
not ( n19515 , n19514 );
buf ( n19516 , n19515 );
buf ( n19517 , n19516 );
nand ( n19518 , n19509 , n19517 );
buf ( n19519 , n19518 );
buf ( n19520 , n19519 );
nand ( n19521 , n19507 , n19520 );
buf ( n19522 , n19521 );
buf ( n19523 , n19522 );
buf ( n19524 , n19523 );
buf ( n19525 , n19504 );
buf ( n19526 , n19500 );
not ( n19527 , n19526 );
buf ( n19528 , n19527 );
buf ( n19529 , n19528 );
buf ( n19530 , n18920 );
not ( n19531 , n19530 );
buf ( n19532 , n19531 );
buf ( n19533 , n19532 );
nand ( n19534 , n19529 , n19533 );
buf ( n19535 , n19534 );
buf ( n19536 , n19535 );
and ( n19537 , n19525 , n19536 );
buf ( n19538 , n19537 );
buf ( n19539 , n19538 );
buf ( n19540 , n19539 );
and ( n19541 , n19093 , n18331 );
and ( n19542 , n19524 , n19540 , n19541 );
nand ( n19543 , n19497 , n19542 );
buf ( n19544 , n18896 );
buf ( n19545 , n19544 );
not ( n19546 , n19545 );
buf ( n19547 , n19513 );
not ( n19548 , n19547 );
buf ( n19549 , n19403 );
buf ( n19550 , n18917 );
buf ( n19551 , n19550 );
nand ( n19552 , n19548 , n19549 , n19551 );
buf ( n19553 , n19552 );
buf ( n19554 , n19553 );
not ( n19555 , n19554 );
or ( n19556 , n19546 , n19555 );
buf ( n19557 , n19553 );
buf ( n19558 , n19544 );
or ( n19559 , n19557 , n19558 );
nand ( n19560 , n19556 , n19559 );
buf ( n19561 , n19560 );
buf ( n19562 , n19561 );
buf ( n19563 , n19562 );
buf ( n19564 , n19516 );
buf ( n19565 , n18379 );
nand ( n19566 , n19564 , n19565 );
buf ( n19567 , n19566 );
buf ( n19568 , n19567 );
buf ( n19569 , n19396 );
buf ( n19570 , n19569 );
not ( n19571 , n19570 );
buf ( n19572 , n19571 );
buf ( n19573 , n19572 );
and ( n19574 , n19568 , n19573 );
not ( n19575 , n19568 );
buf ( n19576 , n19569 );
and ( n19577 , n19575 , n19576 );
nor ( n19578 , n19574 , n19577 );
buf ( n19579 , n19578 );
buf ( n19580 , n19579 );
buf ( n19581 , n19580 );
buf ( n19582 , n19504 );
buf ( n19583 , n19457 );
not ( n19584 , n19583 );
buf ( n19585 , n19584 );
buf ( n19586 , n19585 );
nor ( n19587 , n19582 , n19586 );
buf ( n19588 , n19587 );
buf ( n19589 , n19588 );
buf ( n19590 , n19550 );
and ( n19591 , n19589 , n19590 );
not ( n19592 , n19589 );
buf ( n19593 , n19550 );
not ( n19594 , n19593 );
buf ( n19595 , n19594 );
buf ( n19596 , n19595 );
and ( n19597 , n19592 , n19596 );
nor ( n19598 , n19591 , n19597 );
buf ( n19599 , n19598 );
buf ( n19600 , n19599 );
buf ( n19601 , n19600 );
nand ( n19602 , n19563 , n19581 , n19601 );
nor ( n19603 , n19543 , n19602 );
buf ( n19604 , n19603 );
nand ( n19605 , n19069 , n19604 );
nor ( n19606 , n19479 , n19605 );
buf ( n19607 , n19484 );
buf ( n19608 , n19439 );
nor ( n19609 , n19607 , n19608 );
buf ( n19610 , n19609 );
buf ( n19611 , n19610 );
buf ( n19612 , n19441 );
and ( n19613 , n19611 , n19612 );
not ( n19614 , n19611 );
buf ( n19615 , n19444 );
and ( n19616 , n19614 , n19615 );
nor ( n19617 , n19613 , n19616 );
buf ( n19618 , n19617 );
buf ( n19619 , n19618 );
buf ( n19620 , n19619 );
buf ( n19621 , n19620 );
nand ( n19622 , n19606 , n19621 );
not ( n19623 , n19622 );
or ( n19624 , n19476 , n19623 );
or ( n19625 , n19622 , n19475 );
nand ( n19626 , n19624 , n19625 );
buf ( n19627 , n19626 );
and ( n19628 , n19431 , n19627 );
nor ( n19629 , n19430 , n19628 );
not ( n19630 , n19142 );
nand ( n19631 , n19630 , n19174 );
nor ( n19632 , n19631 , n19377 );
nand ( n19633 , n19632 , n19214 );
buf ( n19634 , n19633 );
not ( n19635 , n19634 );
not ( n19636 , n19635 );
or ( n19637 , n19629 , n19636 );
nand ( n19638 , n19632 , n19352 );
not ( n19639 , n275557 );
and ( n19640 , n19633 , n19638 , n19639 );
not ( n19641 , n19219 );
not ( n19642 , n19632 );
or ( n19643 , n19641 , n19642 );
nand ( n19644 , n19643 , n19317 );
and ( n19645 , n19632 , n19290 );
nor ( n19646 , n19644 , n19645 );
nand ( n19647 , n19632 , n19357 );
and ( n19648 , n19640 , n19646 , n19647 );
not ( n19649 , n19648 );
not ( n19650 , n19649 );
not ( n19651 , n19650 );
not ( n19652 , n19651 );
and ( n19653 , n18862 , n18374 );
nand ( n19654 , n19653 , n18391 );
not ( n19655 , n18898 );
nor ( n19656 , n19654 , n19655 );
and ( n19657 , n19656 , n18887 );
nand ( n19658 , n19657 , n18345 );
not ( n19659 , n18407 );
nor ( n19660 , n19658 , n19659 );
not ( n19661 , n18765 );
and ( n19662 , n19660 , n19661 );
not ( n19663 , n19660 );
and ( n19664 , n19663 , n18766 );
nor ( n19665 , n19662 , n19664 );
not ( n19666 , n19665 );
and ( n19667 , n19652 , n19666 );
buf ( n19668 , n18773 );
buf ( n19669 , n19668 );
not ( n19670 , n19669 );
not ( n19671 , n17768 );
not ( n19672 , n19235 );
or ( n19673 , n19671 , n19672 );
not ( n19674 , n9432 );
buf ( n19675 , n9505 );
buf ( n19676 , n19675 );
buf ( n19677 , n11672 );
buf ( n19678 , n19677 );
or ( n19679 , n19676 , n19678 );
buf ( n19680 , n19679 );
buf ( n19681 , n19680 );
buf ( n19682 , n9513 );
buf ( n19683 , n19682 );
buf ( n19684 , n11592 );
buf ( n19685 , n19684 );
or ( n19686 , n19683 , n19685 );
buf ( n19687 , n19686 );
buf ( n19688 , n19687 );
and ( n19689 , n19681 , n19688 );
buf ( n19690 , n19689 );
buf ( n19691 , n19690 );
not ( n19692 , n19691 );
buf ( n19693 , n9548 );
buf ( n19694 , n19693 );
buf ( n19695 , n10830 );
buf ( n19696 , n19695 );
or ( n19697 , n19694 , n19696 );
buf ( n19698 , n19697 );
buf ( n19699 , n19698 );
buf ( n19700 , n10735 );
buf ( n19701 , n19700 );
not ( n19702 , n19701 );
buf ( n19703 , n9583 );
not ( n19704 , n19703 );
buf ( n19705 , n19704 );
buf ( n19706 , n19705 );
nand ( n19707 , n19702 , n19706 );
buf ( n19708 , n19707 );
buf ( n19709 , n19708 );
and ( n19710 , n19699 , n19709 );
buf ( n19711 , n19710 );
buf ( n19712 , n19711 );
not ( n19713 , n19712 );
buf ( n19714 , n9496 );
buf ( n19715 , n19714 );
buf ( n19716 , n10956 );
buf ( n19717 , n19716 );
or ( n19718 , n19715 , n19717 );
buf ( n19719 , n19718 );
buf ( n19720 , n19719 );
not ( n19721 , n19720 );
buf ( n19722 , n9488 );
buf ( n19723 , n19722 );
buf ( n19724 , n10846 );
buf ( n19725 , n19724 );
and ( n19726 , n19723 , n19725 );
buf ( n19727 , n19726 );
buf ( n19728 , n19727 );
not ( n19729 , n19728 );
or ( n19730 , n19721 , n19729 );
buf ( n19731 , n19714 );
buf ( n19732 , n19716 );
nand ( n19733 , n19731 , n19732 );
buf ( n19734 , n19733 );
buf ( n19735 , n19734 );
nand ( n19736 , n19730 , n19735 );
buf ( n19737 , n19736 );
buf ( n19738 , n19737 );
not ( n19739 , n19738 );
or ( n19740 , n19713 , n19739 );
buf ( n19741 , n19698 );
buf ( n19742 , n19700 );
not ( n19743 , n19742 );
buf ( n19744 , n19705 );
nor ( n19745 , n19743 , n19744 );
buf ( n19746 , n19745 );
buf ( n19747 , n19746 );
and ( n19748 , n19741 , n19747 );
buf ( n19749 , n19693 );
buf ( n19750 , n19695 );
and ( n19751 , n19749 , n19750 );
buf ( n19752 , n19751 );
buf ( n19753 , n19752 );
nor ( n19754 , n19748 , n19753 );
buf ( n19755 , n19754 );
buf ( n19756 , n19755 );
nand ( n19757 , n19740 , n19756 );
buf ( n19758 , n19757 );
buf ( n19759 , n19758 );
not ( n19760 , n19759 );
buf ( n19761 , n9466 );
buf ( n19762 , n19761 );
buf ( n19763 , n19762 );
buf ( n19764 , n11147 );
buf ( n19765 , n19764 );
and ( n19766 , n19763 , n19765 );
buf ( n19767 , n19766 );
buf ( n19768 , n19767 );
not ( n19769 , n19768 );
buf ( n19770 , n19769 );
buf ( n19771 , n19770 );
buf ( n19772 , n9458 );
buf ( n19773 , n19772 );
buf ( n19774 , n19773 );
buf ( n19775 , n11103 );
buf ( n19776 , n19775 );
nand ( n19777 , n19774 , n19776 );
buf ( n19778 , n19777 );
buf ( n19779 , n19778 );
and ( n19780 , n19771 , n19779 );
buf ( n19781 , n19780 );
buf ( n19782 , n19781 );
not ( n19783 , n19782 );
buf ( n19784 , n19258 );
not ( n19785 , n19784 );
buf ( n19786 , n19249 );
not ( n19787 , n19786 );
or ( n19788 , n19785 , n19787 );
buf ( n19789 , n19263 );
nand ( n19790 , n19788 , n19789 );
buf ( n19791 , n19790 );
buf ( n19792 , n19791 );
buf ( n19793 , n19762 );
buf ( n19794 , n19764 );
nor ( n19795 , n19793 , n19794 );
buf ( n19796 , n19795 );
buf ( n19797 , n19796 );
not ( n19798 , n19797 );
buf ( n19799 , n19798 );
buf ( n19800 , n19799 );
nand ( n19801 , n19792 , n19800 );
buf ( n19802 , n19801 );
buf ( n19803 , n19802 );
not ( n19804 , n19803 );
or ( n19805 , n19783 , n19804 );
buf ( n19806 , n19719 );
buf ( n19807 , n19722 );
buf ( n19808 , n19724 );
or ( n19809 , n19807 , n19808 );
buf ( n19810 , n19809 );
buf ( n19811 , n19810 );
nand ( n19812 , n19806 , n19811 );
buf ( n19813 , n19812 );
buf ( n19814 , n19813 );
not ( n19815 , n19814 );
buf ( n19816 , n19815 );
buf ( n19817 , n19816 );
buf ( n19818 , n19711 );
buf ( n19819 , n19778 );
buf ( n19820 , n19773 );
buf ( n19821 , n19775 );
nor ( n19822 , n19820 , n19821 );
buf ( n19823 , n19822 );
buf ( n19824 , n19823 );
nand ( n19825 , n19819 , n19824 );
buf ( n19826 , n19825 );
buf ( n19827 , n19826 );
and ( n19828 , n19817 , n19818 , n19827 );
buf ( n19829 , n19828 );
buf ( n19830 , n19829 );
nand ( n19831 , n19805 , n19830 );
buf ( n19832 , n19831 );
buf ( n19833 , n19832 );
nand ( n19834 , n19760 , n19833 );
buf ( n19835 , n19834 );
buf ( n19836 , n19835 );
not ( n19837 , n19836 );
or ( n19838 , n19692 , n19837 );
buf ( n19839 , n19682 );
buf ( n19840 , n19684 );
and ( n19841 , n19839 , n19840 );
buf ( n19842 , n19841 );
buf ( n19843 , n19842 );
not ( n19844 , n19843 );
buf ( n19845 , n19680 );
not ( n19846 , n19845 );
or ( n19847 , n19844 , n19846 );
buf ( n19848 , n19675 );
buf ( n19849 , n19677 );
nand ( n19850 , n19848 , n19849 );
buf ( n19851 , n19850 );
buf ( n19852 , n19851 );
nand ( n19853 , n19847 , n19852 );
buf ( n19854 , n19853 );
buf ( n19855 , n19854 );
not ( n19856 , n19855 );
buf ( n19857 , n19856 );
buf ( n19858 , n19857 );
nand ( n19859 , n19838 , n19858 );
buf ( n19860 , n19859 );
buf ( n19861 , n19860 );
buf ( n19862 , n9566 );
buf ( n19863 , n19862 );
buf ( n19864 , n11568 );
buf ( n19865 , n19864 );
and ( n19866 , n19863 , n19865 );
buf ( n19867 , n19866 );
buf ( n19868 , n19867 );
not ( n19869 , n19868 );
buf ( n19870 , n19862 );
buf ( n19871 , n19864 );
nor ( n19872 , n19870 , n19871 );
buf ( n19873 , n19872 );
buf ( n19874 , n19873 );
not ( n19875 , n19874 );
buf ( n19876 , n19875 );
buf ( n19877 , n19876 );
nand ( n19878 , n19869 , n19877 );
buf ( n19879 , n19878 );
buf ( n19880 , n19879 );
xnor ( n19881 , n19861 , n19880 );
buf ( n19882 , n19881 );
buf ( n19883 , n19882 );
not ( n19884 , n19883 );
or ( n19885 , n19674 , n19884 );
nand ( n19886 , n9433 , n9566 );
nand ( n19887 , n19885 , n19886 );
nand ( n19888 , n19242 , n19887 );
nand ( n19889 , n19673 , n19888 );
buf ( n19890 , n19889 );
not ( n19891 , n19890 );
or ( n19892 , n19670 , n19891 );
not ( n19893 , n19669 );
not ( n19894 , n19890 );
nand ( n19895 , n19893 , n19894 );
nand ( n19896 , n19892 , n19895 );
not ( n19897 , n277352 );
buf ( n19898 , n19680 );
buf ( n19899 , n19851 );
nand ( n19900 , n19898 , n19899 );
buf ( n19901 , n19900 );
buf ( n19902 , n19901 );
not ( n19903 , n19902 );
buf ( n19904 , n19687 );
not ( n19905 , n19904 );
buf ( n19906 , n19835 );
not ( n19907 , n19906 );
or ( n19908 , n19905 , n19907 );
buf ( n19909 , n19842 );
not ( n19910 , n19909 );
buf ( n19911 , n19910 );
buf ( n19912 , n19911 );
nand ( n19913 , n19908 , n19912 );
buf ( n19914 , n19913 );
buf ( n19915 , n19914 );
not ( n19916 , n19915 );
or ( n19917 , n19903 , n19916 );
buf ( n19918 , n19914 );
buf ( n19919 , n19901 );
or ( n19920 , n19918 , n19919 );
nand ( n19921 , n19917 , n19920 );
buf ( n19922 , n19921 );
buf ( n19923 , n19922 );
not ( n19924 , n19923 );
or ( n19925 , n19897 , n19924 );
nand ( n19926 , n277390 , n9505 );
nand ( n19927 , n19925 , n19926 );
not ( n19928 , n19927 );
not ( n19929 , n19242 );
or ( n19930 , n19928 , n19929 );
not ( n19931 , n17753 );
nand ( n19932 , n19235 , n19931 );
nand ( n19933 , n19930 , n19932 );
buf ( n19934 , n19933 );
not ( n19935 , n19934 );
not ( n19936 , n18414 );
not ( n19937 , n19936 );
buf ( n19938 , n19937 );
and ( n19939 , n19935 , n19938 );
nor ( n19940 , n19896 , n19939 );
not ( n19941 , n19940 );
nand ( n19942 , n19896 , n19939 );
nand ( n19943 , n19941 , n19942 );
not ( n19944 , n19943 );
not ( n19945 , n19938 );
not ( n19946 , n19934 );
or ( n19947 , n19945 , n19946 );
not ( n19948 , n19938 );
nand ( n19949 , n19948 , n19935 );
nand ( n19950 , n19947 , n19949 );
not ( n19951 , n19950 );
buf ( n19952 , n18352 );
buf ( n19953 , n19952 );
not ( n19954 , n19953 );
not ( n19955 , n17780 );
not ( n19956 , n19235 );
or ( n19957 , n19955 , n19956 );
not ( n19958 , n16283 );
buf ( n19959 , n19687 );
buf ( n19960 , n19911 );
nand ( n19961 , n19959 , n19960 );
buf ( n19962 , n19961 );
buf ( n19963 , n19962 );
not ( n19964 , n19963 );
buf ( n19965 , n19835 );
not ( n19966 , n19965 );
or ( n19967 , n19964 , n19966 );
buf ( n19968 , n19835 );
buf ( n19969 , n19962 );
or ( n19970 , n19968 , n19969 );
nand ( n19971 , n19967 , n19970 );
buf ( n19972 , n19971 );
buf ( n19973 , n19972 );
not ( n19974 , n19973 );
or ( n19975 , n19958 , n19974 );
nand ( n19976 , n9433 , n9513 );
nand ( n19977 , n19975 , n19976 );
nand ( n19978 , n19242 , n19977 );
nand ( n19979 , n19957 , n19978 );
buf ( n19980 , n19979 );
nor ( n19981 , n19954 , n19980 );
not ( n19982 , n19981 );
nand ( n19983 , n19951 , n19982 );
not ( n19984 , n19953 );
not ( n19985 , n19980 );
or ( n19986 , n19984 , n19985 );
not ( n19987 , n19980 );
not ( n19988 , n19953 );
nand ( n19989 , n19987 , n19988 );
nand ( n19990 , n19986 , n19989 );
not ( n19991 , n19990 );
buf ( n19992 , n18895 );
buf ( n19993 , n19992 );
not ( n19994 , n19993 );
not ( n19995 , n17795 );
not ( n19996 , n19235 );
or ( n19997 , n19995 , n19996 );
not ( n19998 , n9430 );
buf ( n19999 , n19752 );
not ( n20000 , n19999 );
buf ( n20001 , n19698 );
nand ( n20002 , n20000 , n20001 );
buf ( n20003 , n20002 );
buf ( n20004 , n20003 );
not ( n20005 , n20004 );
buf ( n20006 , n19816 );
buf ( n20007 , n19708 );
and ( n20008 , n20006 , n20007 );
buf ( n20009 , n20008 );
buf ( n20010 , n20009 );
not ( n20011 , n20010 );
buf ( n20012 , n19796 );
buf ( n20013 , n19823 );
nor ( n20014 , n20012 , n20013 );
buf ( n20015 , n20014 );
buf ( n20016 , n20015 );
not ( n20017 , n20016 );
buf ( n20018 , n19791 );
buf ( n20019 , n20018 );
not ( n20020 , n20019 );
or ( n20021 , n20017 , n20020 );
buf ( n20022 , n19773 );
buf ( n20023 , n19775 );
or ( n20024 , n20022 , n20023 );
buf ( n20025 , n20024 );
buf ( n20026 , n20025 );
not ( n20027 , n20026 );
buf ( n20028 , n19767 );
not ( n20029 , n20028 );
or ( n20030 , n20027 , n20029 );
buf ( n20031 , n19778 );
nand ( n20032 , n20030 , n20031 );
buf ( n20033 , n20032 );
buf ( n20034 , n20033 );
not ( n20035 , n20034 );
buf ( n20036 , n20035 );
buf ( n20037 , n20036 );
nand ( n20038 , n20021 , n20037 );
buf ( n20039 , n20038 );
buf ( n20040 , n20039 );
not ( n20041 , n20040 );
or ( n20042 , n20011 , n20041 );
buf ( n20043 , n19737 );
buf ( n20044 , n19708 );
and ( n20045 , n20043 , n20044 );
buf ( n20046 , n19746 );
nor ( n20047 , n20045 , n20046 );
buf ( n20048 , n20047 );
buf ( n20049 , n20048 );
nand ( n20050 , n20042 , n20049 );
buf ( n20051 , n20050 );
buf ( n20052 , n20051 );
not ( n20053 , n20052 );
or ( n20054 , n20005 , n20053 );
buf ( n20055 , n20051 );
buf ( n20056 , n20003 );
or ( n20057 , n20055 , n20056 );
nand ( n20058 , n20054 , n20057 );
buf ( n20059 , n20058 );
buf ( n20060 , n20059 );
not ( n20061 , n20060 );
or ( n20062 , n19998 , n20061 );
nand ( n20063 , n277390 , n9548 );
nand ( n20064 , n20062 , n20063 );
nand ( n20065 , n19242 , n20064 );
nand ( n20066 , n19997 , n20065 );
buf ( n20067 , n20066 );
nor ( n20068 , n19994 , n20067 );
not ( n20069 , n20068 );
nand ( n20070 , n19991 , n20069 );
and ( n20071 , n19983 , n20070 );
not ( n20072 , n20071 );
not ( n20073 , n20072 );
not ( n20074 , n20073 );
buf ( n20075 , n18919 );
not ( n20076 , n18071 );
not ( n20077 , n19235 );
or ( n20078 , n20076 , n20077 );
not ( n20079 , n19772 );
not ( n20080 , n16282 );
or ( n20081 , n20079 , n20080 );
buf ( n20082 , n20025 );
buf ( n20083 , n19778 );
nand ( n20084 , n20082 , n20083 );
buf ( n20085 , n20084 );
buf ( n20086 , n20085 );
not ( n20087 , n20086 );
buf ( n20088 , n19802 );
buf ( n20089 , n19770 );
nand ( n20090 , n20088 , n20089 );
buf ( n20091 , n20090 );
buf ( n20092 , n20091 );
not ( n20093 , n20092 );
or ( n20094 , n20087 , n20093 );
buf ( n20095 , n20091 );
buf ( n20096 , n20085 );
or ( n20097 , n20095 , n20096 );
nand ( n20098 , n20094 , n20097 );
buf ( n20099 , n20098 );
buf ( n20100 , n20099 );
not ( n20101 , n20100 );
or ( n20102 , n20101 , n277390 );
nand ( n20103 , n20081 , n20102 );
nand ( n20104 , n19242 , n20103 );
nand ( n20105 , n20078 , n20104 );
buf ( n20106 , n20105 );
not ( n20107 , n20106 );
xor ( n20108 , n20075 , n20107 );
buf ( n20109 , n18874 );
buf ( n20110 , n20109 );
and ( n20111 , n20108 , n20110 );
and ( n20112 , n20075 , n20107 );
or ( n20113 , n20111 , n20112 );
buf ( n20114 , n18378 );
buf ( n20115 , n20114 );
not ( n20116 , n20115 );
not ( n20117 , n18054 );
not ( n20118 , n19235 );
or ( n20119 , n20117 , n20118 );
not ( n20120 , n277352 );
buf ( n20121 , n19810 );
buf ( n20122 , n19727 );
not ( n20123 , n20122 );
buf ( n20124 , n20123 );
buf ( n20125 , n20124 );
nand ( n20126 , n20121 , n20125 );
buf ( n20127 , n20126 );
buf ( n20128 , n20127 );
not ( n20129 , n20128 );
buf ( n20130 , n20039 );
not ( n20131 , n20130 );
or ( n20132 , n20129 , n20131 );
buf ( n20133 , n20039 );
buf ( n20134 , n20127 );
or ( n20135 , n20133 , n20134 );
nand ( n20136 , n20132 , n20135 );
buf ( n20137 , n20136 );
buf ( n20138 , n20137 );
not ( n20139 , n20138 );
or ( n20140 , n20120 , n20139 );
nand ( n20141 , n277351 , n9488 );
nand ( n20142 , n20140 , n20141 );
nand ( n20143 , n19242 , n20142 );
nand ( n20144 , n20119 , n20143 );
buf ( n20145 , n20144 );
not ( n20146 , n20145 );
or ( n20147 , n20116 , n20146 );
not ( n20148 , n20115 );
not ( n20149 , n20145 );
nand ( n20150 , n20148 , n20149 );
nand ( n20151 , n20147 , n20150 );
and ( n20152 , n20113 , n20151 );
not ( n20153 , n20152 );
buf ( n20154 , n18398 );
buf ( n20155 , n20154 );
not ( n20156 , n20155 );
not ( n20157 , n18101 );
not ( n20158 , n19235 );
or ( n20159 , n20157 , n20158 );
not ( n20160 , n277603 );
buf ( n20161 , n19810 );
not ( n20162 , n20161 );
buf ( n20163 , n20039 );
not ( n20164 , n20163 );
or ( n20165 , n20162 , n20164 );
buf ( n20166 , n20124 );
nand ( n20167 , n20165 , n20166 );
buf ( n20168 , n20167 );
buf ( n20169 , n20168 );
buf ( n20170 , n19719 );
buf ( n20171 , n19734 );
nand ( n20172 , n20170 , n20171 );
buf ( n20173 , n20172 );
buf ( n20174 , n20173 );
xnor ( n20175 , n20169 , n20174 );
buf ( n20176 , n20175 );
buf ( n20177 , n20176 );
not ( n20178 , n20177 );
or ( n20179 , n20160 , n20178 );
nand ( n20180 , n16282 , n9496 );
nand ( n20181 , n20179 , n20180 );
nand ( n20182 , n19242 , n20181 );
nand ( n20183 , n20159 , n20182 );
buf ( n20184 , n20183 );
not ( n20185 , n20184 );
or ( n20186 , n20156 , n20185 );
not ( n20187 , n20184 );
not ( n20188 , n20155 );
nand ( n20189 , n20187 , n20188 );
nand ( n20190 , n20186 , n20189 );
not ( n20191 , n20190 );
nor ( n20192 , n20145 , n20148 );
not ( n20193 , n20192 );
nand ( n20194 , n20191 , n20193 );
not ( n20195 , n20194 );
or ( n20196 , n20153 , n20195 );
not ( n20197 , n20193 );
buf ( n20198 , n20190 );
nand ( n20199 , n20197 , n20198 );
nand ( n20200 , n20196 , n20199 );
not ( n20201 , n20067 );
not ( n20202 , n19993 );
or ( n20203 , n20201 , n20202 );
not ( n20204 , n20067 );
nand ( n20205 , n20204 , n19994 );
nand ( n20206 , n20203 , n20205 );
buf ( n20207 , n18916 );
buf ( n20208 , n20207 );
not ( n20209 , n20208 );
not ( n20210 , n18086 );
not ( n20211 , n19235 );
or ( n20212 , n20210 , n20211 );
not ( n20213 , n9430 );
buf ( n20214 , n19816 );
not ( n20215 , n20214 );
buf ( n20216 , n20039 );
not ( n20217 , n20216 );
or ( n20218 , n20215 , n20217 );
buf ( n20219 , n19737 );
not ( n20220 , n20219 );
buf ( n20221 , n20220 );
buf ( n20222 , n20221 );
nand ( n20223 , n20218 , n20222 );
buf ( n20224 , n20223 );
buf ( n20225 , n20224 );
buf ( n20226 , n19746 );
not ( n20227 , n20226 );
buf ( n20228 , n19708 );
nand ( n20229 , n20227 , n20228 );
buf ( n20230 , n20229 );
buf ( n20231 , n20230 );
xnor ( n20232 , n20225 , n20231 );
buf ( n20233 , n20232 );
buf ( n20234 , n20233 );
not ( n20235 , n20234 );
or ( n20236 , n20213 , n20235 );
nand ( n20237 , n16282 , n9583 );
nand ( n20238 , n20236 , n20237 );
nand ( n20239 , n19242 , n20238 );
nand ( n20240 , n20212 , n20239 );
buf ( n20241 , n20240 );
nor ( n20242 , n20209 , n20241 );
nor ( n20243 , n20206 , n20242 );
not ( n20244 , n20208 );
not ( n20245 , n20244 );
not ( n20246 , n20241 );
not ( n20247 , n20246 );
or ( n20248 , n20245 , n20247 );
nand ( n20249 , n20241 , n20208 );
nand ( n20250 , n20248 , n20249 );
nor ( n20251 , n20184 , n20188 );
nor ( n20252 , n20250 , n20251 );
nor ( n20253 , n20243 , n20252 );
buf ( n20254 , n20253 );
nand ( n20255 , n20200 , n20254 );
buf ( n20256 , n20251 );
nand ( n20257 , n20250 , n20256 );
or ( n20258 , n20243 , n20257 );
buf ( n20259 , n20206 );
buf ( n20260 , n20242 );
nand ( n20261 , n20259 , n20260 );
nand ( n20262 , n20258 , n20261 );
not ( n20263 , n20262 );
and ( n20264 , n20255 , n20263 );
not ( n20265 , n19321 );
nand ( n20266 , n20265 , n19324 );
not ( n20267 , n20266 );
not ( n20268 , n19340 );
or ( n20269 , n20267 , n20268 );
not ( n20270 , n18115 );
not ( n20271 , n19235 );
or ( n20272 , n20270 , n20271 );
not ( n20273 , n19761 );
not ( n20274 , n16282 );
or ( n20275 , n20273 , n20274 );
buf ( n20276 , n19799 );
buf ( n20277 , n19770 );
nand ( n20278 , n20276 , n20277 );
buf ( n20279 , n20278 );
buf ( n20280 , n20279 );
not ( n20281 , n20280 );
buf ( n20282 , n20018 );
not ( n20283 , n20282 );
or ( n20284 , n20281 , n20283 );
buf ( n20285 , n20018 );
buf ( n20286 , n20279 );
or ( n20287 , n20285 , n20286 );
nand ( n20288 , n20284 , n20287 );
buf ( n20289 , n20288 );
buf ( n20290 , n20289 );
nand ( n20291 , n20290 , n277817 );
nand ( n20292 , n20275 , n20291 );
nand ( n20293 , n19242 , n20292 );
nand ( n20294 , n20272 , n20293 );
buf ( n20295 , n20294 );
not ( n20296 , n20295 );
not ( n20297 , n20296 );
buf ( n20298 , n18330 );
not ( n20299 , n20298 );
not ( n20300 , n20299 );
or ( n20301 , n20297 , n20300 );
nand ( n20302 , n20298 , n20295 );
nand ( n20303 , n20301 , n20302 );
and ( n20304 , n19331 , n19329 );
nor ( n20305 , n20303 , n20304 );
nor ( n20306 , n19337 , n20305 );
nand ( n20307 , n20269 , n20306 );
not ( n20308 , n20307 );
not ( n20309 , n20308 );
xor ( n20310 , n20075 , n20107 );
xor ( n20311 , n20310 , n20110 );
not ( n20312 , n20311 );
not ( n20313 , n20298 );
nor ( n20314 , n20313 , n20295 );
not ( n20315 , n20314 );
nand ( n20316 , n20312 , n20315 );
not ( n20317 , n20316 );
not ( n20318 , n20317 );
not ( n20319 , n20318 );
or ( n20320 , n20309 , n20319 );
not ( n20321 , n20317 );
buf ( n20322 , n20303 );
nand ( n20323 , n20322 , n20304 );
not ( n20324 , n20323 );
and ( n20325 , n20321 , n20324 );
buf ( n20326 , n20311 );
nand ( n20327 , n20326 , n20314 );
not ( n20328 , n20327 );
nor ( n20329 , n20325 , n20328 );
nand ( n20330 , n20320 , n20329 );
not ( n20331 , n20113 );
not ( n20332 , n20151 );
nand ( n20333 , n20331 , n20332 );
and ( n20334 , n20194 , n20333 );
and ( n20335 , n20334 , n20254 );
nand ( n20336 , n20330 , n20335 );
nand ( n20337 , n20264 , n20336 );
not ( n20338 , n20337 );
or ( n20339 , n20074 , n20338 );
and ( n20340 , n19990 , n20068 );
not ( n20341 , n20340 );
not ( n20342 , n19983 );
or ( n20343 , n20341 , n20342 );
or ( n20344 , n19951 , n19982 );
nand ( n20345 , n20343 , n20344 );
not ( n20346 , n20345 );
nand ( n20347 , n20339 , n20346 );
not ( n20348 , n20347 );
or ( n20349 , n19944 , n20348 );
or ( n20350 , n20347 , n19943 );
nand ( n20351 , n20349 , n20350 );
buf ( n20352 , n20351 );
not ( n20353 , n19638 );
and ( n20354 , n20352 , n20353 );
nor ( n20355 , n19667 , n20354 );
buf ( n20356 , n19889 );
not ( n20357 , n20356 );
not ( n20358 , n20357 );
buf ( n20359 , n18773 );
not ( n20360 , n20359 );
or ( n20361 , n20358 , n20360 );
not ( n20362 , n20359 );
nand ( n20363 , n20356 , n20362 );
nand ( n20364 , n20361 , n20363 );
buf ( n20365 , n19933 );
not ( n20366 , n19936 );
buf ( n20367 , n20366 );
and ( n20368 , n20365 , n20367 );
or ( n20369 , n20364 , n20368 );
not ( n20370 , n20369 );
not ( n20371 , n20370 );
nand ( n20372 , n20364 , n20368 );
nand ( n20373 , n20371 , n20372 );
not ( n20374 , n20373 );
not ( n20375 , n20367 );
not ( n20376 , n20375 );
not ( n20377 , n20365 );
or ( n20378 , n20376 , n20377 );
not ( n20379 , n20365 );
nand ( n20380 , n20379 , n20367 );
nand ( n20381 , n20378 , n20380 );
not ( n20382 , n20381 );
buf ( n20383 , n19952 );
buf ( n20384 , n19979 );
and ( n20385 , n20383 , n20384 );
not ( n20386 , n20385 );
nand ( n20387 , n20382 , n20386 );
not ( n20388 , n20383 );
not ( n20389 , n20388 );
not ( n20390 , n20384 );
or ( n20391 , n20389 , n20390 );
not ( n20392 , n20384 );
nand ( n20393 , n20392 , n20383 );
nand ( n20394 , n20391 , n20393 );
not ( n20395 , n20394 );
buf ( n20396 , n20066 );
buf ( n20397 , n19992 );
and ( n20398 , n20396 , n20397 );
not ( n20399 , n20398 );
nand ( n20400 , n20395 , n20399 );
nand ( n20401 , n20387 , n20400 );
not ( n20402 , n20401 );
not ( n20403 , n20402 );
buf ( n20404 , n18919 );
buf ( n20405 , n20105 );
xor ( n20406 , n20404 , n20405 );
buf ( n20407 , n20109 );
xor ( n20408 , n20406 , n20407 );
buf ( n20409 , n20294 );
buf ( n20410 , n18330 );
and ( n20411 , n20409 , n20410 );
nor ( n20412 , n20408 , n20411 );
not ( n20413 , n20412 );
xor ( n20414 , n20409 , n20410 );
and ( n20415 , n19365 , n19366 );
nor ( n20416 , n20414 , n20415 );
not ( n20417 , n19363 );
nand ( n20418 , n20417 , n19367 );
nor ( n20419 , n20416 , n20418 );
nand ( n20420 , n20413 , n20419 );
nand ( n20421 , n20414 , n20415 );
not ( n20422 , n20421 );
nand ( n20423 , n20413 , n20422 );
nand ( n20424 , n20408 , n20411 );
nand ( n20425 , n20420 , n20423 , n20424 );
buf ( n20426 , n20183 );
not ( n20427 , n20426 );
buf ( n20428 , n20154 );
buf ( n20429 , n20428 );
not ( n20430 , n20429 );
not ( n20431 , n20430 );
or ( n20432 , n20427 , n20431 );
not ( n20433 , n20426 );
nand ( n20434 , n20433 , n20429 );
nand ( n20435 , n20432 , n20434 );
not ( n20436 , n20435 );
buf ( n20437 , n20114 );
buf ( n20438 , n20144 );
and ( n20439 , n20437 , n20438 );
not ( n20440 , n20439 );
nand ( n20441 , n20436 , n20440 );
xor ( n20442 , n20404 , n20405 );
and ( n20443 , n20442 , n20407 );
and ( n20444 , n20404 , n20405 );
or ( n20445 , n20443 , n20444 );
not ( n20446 , n20445 );
xor ( n20447 , n20437 , n20438 );
not ( n20448 , n20447 );
nand ( n20449 , n20446 , n20448 );
nand ( n20450 , n20441 , n20449 );
buf ( n20451 , n20240 );
not ( n20452 , n20451 );
not ( n20453 , n20452 );
buf ( n20454 , n20207 );
not ( n20455 , n20454 );
or ( n20456 , n20453 , n20455 );
not ( n20457 , n20454 );
nand ( n20458 , n20457 , n20451 );
nand ( n20459 , n20456 , n20458 );
not ( n20460 , n20459 );
and ( n20461 , n20426 , n20429 );
not ( n20462 , n20461 );
nand ( n20463 , n20460 , n20462 );
not ( n20464 , n20396 );
not ( n20465 , n20464 );
not ( n20466 , n20397 );
or ( n20467 , n20465 , n20466 );
not ( n20468 , n20397 );
nand ( n20469 , n20468 , n20396 );
nand ( n20470 , n20467 , n20469 );
nand ( n20471 , n20454 , n20451 );
not ( n20472 , n20471 );
nor ( n20473 , n20470 , n20472 );
not ( n20474 , n20473 );
nand ( n20475 , n20463 , n20474 );
nor ( n20476 , n20450 , n20475 );
nand ( n20477 , n20425 , n20476 );
not ( n20478 , n20475 );
not ( n20479 , n20478 );
not ( n20480 , n20445 );
nor ( n20481 , n20480 , n20448 );
not ( n20482 , n20481 );
not ( n20483 , n20441 );
or ( n20484 , n20482 , n20483 );
or ( n20485 , n20436 , n20440 );
nand ( n20486 , n20484 , n20485 );
not ( n20487 , n20486 );
or ( n20488 , n20479 , n20487 );
not ( n20489 , n20473 );
nand ( n20490 , n20459 , n20461 );
not ( n20491 , n20490 );
and ( n20492 , n20489 , n20491 );
nand ( n20493 , n20470 , n20472 );
not ( n20494 , n20493 );
nor ( n20495 , n20492 , n20494 );
not ( n20496 , n20495 );
not ( n20497 , n20496 );
nand ( n20498 , n20488 , n20497 );
not ( n20499 , n20498 );
nand ( n20500 , n20477 , n20499 );
not ( n20501 , n20500 );
or ( n20502 , n20403 , n20501 );
not ( n20503 , n20387 );
nand ( n20504 , n20394 , n20398 );
nor ( n20505 , n20503 , n20504 );
nand ( n20506 , n20381 , n20385 );
not ( n20507 , n20506 );
nor ( n20508 , n20505 , n20507 );
nand ( n20509 , n20502 , n20508 );
not ( n20510 , n20509 );
or ( n20511 , n20374 , n20510 );
or ( n20512 , n20509 , n20373 );
nand ( n20513 , n20511 , n20512 );
buf ( n20514 , n20513 );
not ( n20515 , n19647 );
and ( n20516 , n20514 , n20515 );
nor ( n20517 , n19639 , n19661 );
not ( n20518 , n20517 );
buf ( n20519 , n19889 );
buf ( n20520 , n20519 );
not ( n20521 , n20520 );
not ( n20522 , n20521 );
not ( n20523 , n20240 );
not ( n20524 , n20523 );
buf ( n20525 , n20524 );
not ( n20526 , n20066 );
not ( n20527 , n20526 );
buf ( n20528 , n20527 );
nor ( n20529 , n20525 , n20528 );
not ( n20530 , n20529 );
buf ( n20531 , n20183 );
buf ( n20532 , n20531 );
not ( n20533 , n20532 );
buf ( n20534 , n20144 );
buf ( n20535 , n20534 );
not ( n20536 , n20535 );
nand ( n20537 , n20533 , n20536 );
nor ( n20538 , n20530 , n20537 );
nor ( n20539 , n19309 , n19293 );
buf ( n20540 , n20294 );
buf ( n20541 , n20540 );
buf ( n20542 , n20105 );
buf ( n20543 , n20542 );
nor ( n20544 , n20541 , n20543 );
nand ( n20545 , n20539 , n20544 );
not ( n20546 , n20545 );
and ( n20547 , n20538 , n20546 );
buf ( n20548 , n19933 );
buf ( n20549 , n20548 );
buf ( n20550 , n19979 );
buf ( n20551 , n20550 );
nor ( n20552 , n20549 , n20551 );
nand ( n20553 , n20547 , n20552 );
not ( n20554 , n20553 );
or ( n20555 , n20522 , n20554 );
or ( n20556 , n20553 , n20521 );
nand ( n20557 , n20555 , n20556 );
buf ( n20558 , n20557 );
not ( n20559 , n19645 );
not ( n20560 , n20559 );
nand ( n20561 , n20558 , n20560 );
not ( n20562 , n19644 );
not ( n20563 , n20562 );
buf ( n20564 , n20519 );
buf ( n20565 , n20564 );
buf ( n20566 , n20565 );
nand ( n20567 , n20563 , n20566 );
nand ( n20568 , n20518 , n20561 , n20567 );
nor ( n20569 , n20516 , n20568 );
and ( n20570 , n20355 , n20569 );
nand ( n20571 , n19637 , n20570 );
buf ( n20572 , n20571 );
buf ( n20573 , n20572 );
buf ( n20574 , n275554 );
not ( n20575 , n275929 );
buf ( n20576 , n20575 );
buf ( n20577 , n20576 );
buf ( n20578 , n275554 );
not ( n20579 , n9063 );
not ( n20580 , n9171 );
nand ( n20581 , n20579 , n20580 );
nand ( n20582 , n11730 , n20581 );
and ( n20583 , n20582 , n275739 );
not ( n20584 , n20582 );
not ( n20585 , n9063 );
not ( n20586 , n20585 );
nand ( n20587 , n20586 , n9171 );
not ( n20588 , n20587 );
buf ( n20589 , n276324 );
not ( n20590 , n20589 );
buf ( n20591 , n11040 );
or ( n20592 , n20590 , n20591 );
nand ( n20593 , n20590 , n20591 );
nand ( n20594 , n20592 , n20593 );
buf ( n20595 , n20594 );
and ( n20596 , n20588 , n20595 );
buf ( n20597 , n276324 );
not ( n20598 , n20597 );
buf ( n20599 , n11018 );
or ( n20600 , n20598 , n20599 );
nand ( n20601 , n20598 , n20599 );
nand ( n20602 , n20600 , n20601 );
buf ( n20603 , n20602 );
not ( n20604 , n20603 );
not ( n20605 , n20580 );
or ( n20606 , n20604 , n20605 );
not ( n20607 , n275945 );
or ( n20608 , n20586 , n20607 );
nand ( n20609 , n20606 , n20608 );
nor ( n20610 , n20596 , n20609 );
and ( n20611 , n20584 , n20610 );
nor ( n20612 , n20583 , n20611 );
not ( n20613 , n9088 );
not ( n20614 , n20613 );
and ( n20615 , n9094 , n9099 );
nand ( n20616 , n20614 , n20615 );
not ( n20617 , n20616 );
nor ( n20618 , n20612 , n20617 );
buf ( n20619 , n11018 );
not ( n20620 , n20619 );
buf ( n20621 , n276325 );
or ( n20622 , n20620 , n20621 );
nand ( n20623 , n20621 , n20620 );
nand ( n20624 , n20622 , n20623 );
buf ( n20625 , n20624 );
not ( n20626 , n20625 );
not ( n20627 , n20581 );
nand ( n20628 , n20626 , n20627 );
buf ( n20629 , n11040 );
not ( n20630 , n20629 );
buf ( n20631 , n276325 );
or ( n20632 , n20630 , n20631 );
nand ( n20633 , n20631 , n20630 );
nand ( n20634 , n20632 , n20633 );
buf ( n20635 , n20634 );
not ( n20636 , n20635 );
nor ( n20637 , n9063 , n20580 );
nand ( n20638 , n20636 , n20637 );
nand ( n20639 , n20586 , n20607 );
nand ( n20640 , n20628 , n20638 , n20639 );
nand ( n20641 , n20640 , n20617 );
not ( n20642 , n9183 );
nand ( n20643 , n20642 , n9159 );
buf ( n20644 , n20643 );
not ( n20645 , n20644 );
nand ( n20646 , n20641 , n20645 );
or ( n20647 , n20618 , n20646 );
not ( n20648 , n11034 );
not ( n20649 , n9159 );
not ( n20650 , n20649 );
or ( n20651 , n20648 , n20650 );
not ( n20652 , n9184 );
nor ( n20653 , n20652 , n9411 );
not ( n20654 , n20653 );
or ( n20655 , n20654 , n275739 );
nand ( n20656 , n20651 , n20655 );
nand ( n20657 , n9411 , n9184 );
nor ( n20658 , n20610 , n20657 );
nor ( n20659 , n20656 , n20658 );
nand ( n20660 , n20647 , n20659 );
buf ( n20661 , n20660 );
buf ( n20662 , n20661 );
not ( n20663 , n14543 );
buf ( n20664 , n14778 );
not ( n20665 , n20664 );
not ( n20666 , n20665 );
or ( n20667 , n20663 , n20666 );
not ( n20668 , n14543 );
nand ( n20669 , n20664 , n20668 );
nand ( n20670 , n20667 , n20669 );
buf ( n20671 , n20670 );
not ( n20672 , n13373 );
nand ( n20673 , n20671 , n20672 );
or ( n20674 , n20673 , n14908 );
not ( n20675 , n17500 );
not ( n20676 , n17410 );
or ( n20677 , n20675 , n20676 );
buf ( n20678 , n16721 );
buf ( n20679 , n20678 );
buf ( n20680 , n20679 );
nand ( n20681 , n20677 , n20680 );
not ( n20682 , n17296 );
not ( n20683 , n17293 );
or ( n20684 , n20682 , n20683 );
or ( n20685 , n17293 , n17296 );
nand ( n20686 , n20684 , n20685 );
buf ( n20687 , n20686 );
and ( n20688 , n17404 , n20687 );
not ( n20689 , n14772 );
nor ( n20690 , n17561 , n20689 );
nor ( n20691 , n20688 , n20690 );
not ( n20692 , n16723 );
not ( n20693 , n16706 );
or ( n20694 , n20692 , n20693 );
or ( n20695 , n16706 , n16723 );
nand ( n20696 , n20694 , n20695 );
buf ( n20697 , n20696 );
and ( n20698 , n16968 , n20697 );
and ( n20699 , n17545 , n14761 );
nor ( n20700 , n20698 , n20699 );
and ( n20701 , n20681 , n20691 , n20700 );
nand ( n20702 , n20674 , n20701 );
buf ( n20703 , n20702 );
buf ( n20704 , n20703 );
not ( n20705 , n275929 );
buf ( n20706 , n20705 );
buf ( n20707 , n20706 );
not ( n20708 , n275929 );
buf ( n20709 , n20708 );
buf ( n20710 , n20709 );
not ( n20711 , n20672 );
buf ( n20712 , n20711 );
buf ( n20713 , n14404 );
and ( n20714 , n20712 , n20713 );
not ( n20715 , n20712 );
nand ( n20716 , n14276 , n14293 , n14212 );
nor ( n20717 , n14617 , n20716 );
buf ( n20718 , n20717 );
nand ( n20719 , n14778 , n20718 );
buf ( n20720 , n20719 );
buf ( n20721 , n14427 );
buf ( n20722 , n14185 );
buf ( n20723 , n14360 );
buf ( n20724 , n14080 );
nand ( n20725 , n20722 , n20723 , n20724 );
nor ( n20726 , n20721 , n20725 );
nand ( n20727 , n14132 , n14154 );
nor ( n20728 , n14252 , n20727 );
buf ( n20729 , n20728 );
nand ( n20730 , n20726 , n20729 );
nor ( n20731 , n20720 , n20730 );
buf ( n20732 , n14384 );
and ( n20733 , n20731 , n20732 );
not ( n20734 , n20731 );
not ( n20735 , n20732 );
and ( n20736 , n20734 , n20735 );
nor ( n20737 , n20733 , n20736 );
buf ( n20738 , n20737 );
and ( n20739 , n20715 , n20738 );
nor ( n20740 , n20714 , n20739 );
not ( n20741 , n14908 );
not ( n20742 , n20741 );
buf ( n20743 , n20742 );
or ( n20744 , n20740 , n20743 );
nand ( n20745 , n17076 , n17371 );
not ( n20746 , n20745 );
buf ( n20747 , n17034 );
not ( n20748 , n17087 );
nor ( n20749 , n20747 , n20748 );
not ( n20750 , n20749 );
not ( n20751 , n17362 );
or ( n20752 , n20750 , n20751 );
and ( n20753 , n17381 , n17387 );
or ( n20754 , n20753 , n20748 );
nand ( n20755 , n20754 , n17369 );
not ( n20756 , n20755 );
nand ( n20757 , n20752 , n20756 );
not ( n20758 , n20757 );
or ( n20759 , n20746 , n20758 );
or ( n20760 , n20757 , n20745 );
nand ( n20761 , n20759 , n20760 );
buf ( n20762 , n20761 );
buf ( n20763 , n17405 );
and ( n20764 , n20762 , n20763 );
not ( n20765 , n17545 );
not ( n20766 , n20765 );
and ( n20767 , n17528 , n13828 );
not ( n20768 , n17528 );
and ( n20769 , n20768 , n17529 );
nor ( n20770 , n20767 , n20769 );
not ( n20771 , n20770 );
and ( n20772 , n20766 , n20771 );
not ( n20773 , n17465 );
nor ( n20774 , n17481 , n17470 );
and ( n20775 , n20774 , n17489 , n17479 );
not ( n20776 , n17467 );
and ( n20777 , n17462 , n20775 , n20776 );
not ( n20778 , n20777 );
or ( n20779 , n20773 , n20778 );
or ( n20780 , n20777 , n17465 );
nand ( n20781 , n20779 , n20780 );
buf ( n20782 , n20781 );
and ( n20783 , n17411 , n20782 );
nor ( n20784 , n20772 , n20783 );
not ( n20785 , n17500 );
buf ( n20786 , n17464 );
buf ( n20787 , n20786 );
buf ( n20788 , n20787 );
nand ( n20789 , n20785 , n20788 );
nand ( n20790 , n17560 , n13823 );
nand ( n20791 , n20784 , n20789 , n20790 );
nor ( n20792 , n20764 , n20791 );
not ( n20793 , n16124 );
nand ( n20794 , n20793 , n16932 );
not ( n20795 , n20794 );
buf ( n20796 , n15909 );
not ( n20797 , n16135 );
nor ( n20798 , n20796 , n20797 );
not ( n20799 , n20798 );
not ( n20800 , n16913 );
or ( n20801 , n20799 , n20800 );
not ( n20802 , n16938 );
buf ( n20803 , n16924 );
nor ( n20804 , n20802 , n20803 );
or ( n20805 , n20804 , n20797 );
nand ( n20806 , n20805 , n16930 );
not ( n20807 , n20806 );
nand ( n20808 , n20801 , n20807 );
not ( n20809 , n20808 );
or ( n20810 , n20795 , n20809 );
or ( n20811 , n20808 , n20794 );
nand ( n20812 , n20810 , n20811 );
buf ( n20813 , n20812 );
nand ( n20814 , n20813 , n16970 );
and ( n20815 , n20792 , n20814 );
nand ( n20816 , n20744 , n20815 );
buf ( n20817 , n20816 );
buf ( n20818 , n20817 );
buf ( n20819 , n275554 );
buf ( n20820 , n14275 );
and ( n20821 , n13373 , n20820 );
not ( n20822 , n13373 );
not ( n20823 , n14213 );
not ( n20824 , n20823 );
buf ( n20825 , n14616 );
nand ( n20826 , n14777 , n20825 );
buf ( n20827 , n14514 );
not ( n20828 , n20827 );
nor ( n20829 , n20826 , n20828 );
buf ( n20830 , n14276 );
buf ( n20831 , n14487 );
and ( n20832 , n20830 , n20831 );
nand ( n20833 , n20829 , n20832 );
buf ( n20834 , n14449 );
not ( n20835 , n20834 );
nor ( n20836 , n20833 , n20835 );
buf ( n20837 , n20836 );
not ( n20838 , n20837 );
or ( n20839 , n20824 , n20838 );
or ( n20840 , n20837 , n20823 );
nand ( n20841 , n20839 , n20840 );
buf ( n20842 , n20841 );
and ( n20843 , n20822 , n20842 );
nor ( n20844 , n20821 , n20843 );
not ( n20845 , n20844 );
buf ( n20846 , n14895 );
not ( n20847 , n20846 );
and ( n20848 , n20845 , n20847 );
buf ( n20849 , n16293 );
not ( n20850 , n20849 );
nand ( n20851 , n20850 , n16901 );
not ( n20852 , n20851 );
not ( n20853 , n16401 );
nor ( n20854 , n16862 , n16499 );
not ( n20855 , n20854 );
not ( n20856 , n16863 );
not ( n20857 , n20856 );
not ( n20858 , n16761 );
not ( n20859 , n20858 );
or ( n20860 , n20857 , n20859 );
not ( n20861 , n16803 );
and ( n20862 , n20856 , n20861 );
not ( n20863 , n16802 );
nor ( n20864 , n20862 , n20863 );
nand ( n20865 , n20860 , n20864 );
not ( n20866 , n20865 );
or ( n20867 , n20855 , n20866 );
not ( n20868 , n16499 );
not ( n20869 , n20868 );
not ( n20870 , n16874 );
or ( n20871 , n20869 , n20870 );
not ( n20872 , n16875 );
nand ( n20873 , n20871 , n20872 );
not ( n20874 , n20873 );
nand ( n20875 , n20867 , n20874 );
not ( n20876 , n20875 );
or ( n20877 , n20853 , n20876 );
not ( n20878 , n16896 );
nor ( n20879 , n20878 , n16899 );
nand ( n20880 , n20877 , n20879 );
not ( n20881 , n20880 );
or ( n20882 , n20852 , n20881 );
or ( n20883 , n20880 , n20851 );
nand ( n20884 , n20882 , n20883 );
buf ( n20885 , n20884 );
and ( n20886 , n17556 , n16957 );
and ( n20887 , n14894 , n17540 );
nor ( n20888 , n20886 , n20887 );
not ( n20889 , n20888 );
nand ( n20890 , n20885 , n20889 );
buf ( n20891 , n17338 );
nand ( n20892 , n17207 , n20891 );
not ( n20893 , n20892 );
not ( n20894 , n17228 );
not ( n20895 , n17180 );
buf ( n20896 , n17282 );
nor ( n20897 , n20895 , n20896 );
not ( n20898 , n20897 );
not ( n20899 , n17314 );
nand ( n20900 , n20899 , n17252 );
not ( n20901 , n17311 );
nand ( n20902 , n17252 , n20901 );
buf ( n20903 , n17312 );
nand ( n20904 , n20900 , n20902 , n20903 );
not ( n20905 , n20904 );
or ( n20906 , n20898 , n20905 );
not ( n20907 , n17180 );
buf ( n20908 , n17325 );
not ( n20909 , n20908 );
or ( n20910 , n20907 , n20909 );
nand ( n20911 , n20910 , n17327 );
not ( n20912 , n20911 );
nand ( n20913 , n20906 , n20912 );
not ( n20914 , n20913 );
or ( n20915 , n20894 , n20914 );
buf ( n20916 , n17337 );
buf ( n20917 , n17339 );
and ( n20918 , n20916 , n20917 );
nand ( n20919 , n20915 , n20918 );
not ( n20920 , n20919 );
or ( n20921 , n20893 , n20920 );
or ( n20922 , n20919 , n20892 );
nand ( n20923 , n20921 , n20922 );
buf ( n20924 , n20923 );
buf ( n20925 , n17403 );
not ( n20926 , n20925 );
buf ( n20927 , n20926 );
nand ( n20928 , n20924 , n20927 );
not ( n20929 , n17440 );
buf ( n20930 , n17434 );
nor ( n20931 , n20929 , n20930 );
not ( n20932 , n17442 );
and ( n20933 , n20931 , n20932 );
not ( n20934 , n20931 );
and ( n20935 , n20934 , n17442 );
nor ( n20936 , n20933 , n20935 );
buf ( n20937 , n20936 );
and ( n20938 , n20937 , n17409 );
not ( n20939 , n17499 );
not ( n20940 , n20939 );
buf ( n20941 , n17441 );
buf ( n20942 , n20941 );
buf ( n20943 , n20942 );
and ( n20944 , n20940 , n20943 );
nor ( n20945 , n20938 , n20944 );
nand ( n20946 , n20890 , n20928 , n20945 );
nor ( n20947 , n20848 , n20946 );
nand ( n20948 , n17547 , n16965 , n14868 );
not ( n20949 , n20948 );
nand ( n20950 , n20949 , n17558 );
buf ( n20951 , n20950 );
or ( n20952 , n20947 , n20951 );
buf ( n20953 , n20950 );
nand ( n20954 , n20953 , n13481 );
nand ( n20955 , n20952 , n20954 );
buf ( n20956 , n20955 );
buf ( n20957 , n20956 );
not ( n20958 , n14824 );
nand ( n20959 , n14825 , n14837 , n14829 );
nor ( n20960 , n20958 , n20959 );
nand ( n20961 , n20960 , n14823 );
not ( n20962 , n20961 );
buf ( n20963 , n20962 );
buf ( n20964 , n20963 );
not ( n20965 , n275550 );
buf ( n20966 , n20965 );
buf ( n20967 , n20966 );
buf ( n20968 , n275554 );
buf ( n20969 , n275554 );
buf ( n20970 , n275554 );
and ( n20971 , n18208 , n19092 );
not ( n20972 , n18208 );
buf ( n20973 , n19540 );
not ( n20974 , n20973 );
not ( n20975 , n20974 );
buf ( n20976 , n19541 );
nand ( n20977 , n19069 , n20976 );
not ( n20978 , n20977 );
not ( n20979 , n20978 );
or ( n20980 , n20975 , n20979 );
or ( n20981 , n20978 , n20974 );
nand ( n20982 , n20980 , n20981 );
buf ( n20983 , n20982 );
and ( n20984 , n20972 , n20983 );
nor ( n20985 , n20971 , n20984 );
not ( n20986 , n20985 );
buf ( n20987 , n19200 );
and ( n20988 , n20986 , n20987 );
not ( n20989 , n20305 );
nand ( n20990 , n20989 , n20323 );
not ( n20991 , n20990 );
or ( n20992 , n19338 , n19325 );
nand ( n20993 , n20992 , n19341 );
not ( n20994 , n20993 );
or ( n20995 , n20991 , n20994 );
or ( n20996 , n20993 , n20990 );
nand ( n20997 , n20995 , n20996 );
buf ( n20998 , n20997 );
and ( n20999 , n19218 , n19288 );
nor ( n21000 , n20999 , n19348 );
not ( n21001 , n21000 );
nand ( n21002 , n20998 , n21001 );
not ( n21003 , n20418 );
not ( n21004 , n21003 );
not ( n21005 , n20416 );
nand ( n21006 , n21005 , n20421 );
not ( n21007 , n21006 );
or ( n21008 , n21004 , n21007 );
or ( n21009 , n21006 , n21003 );
nand ( n21010 , n21008 , n21009 );
buf ( n21011 , n21010 );
nand ( n21012 , n21011 , n19358 );
not ( n21013 , n20541 );
not ( n21014 , n20539 );
or ( n21015 , n21013 , n21014 );
or ( n21016 , n20539 , n20541 );
nand ( n21017 , n21015 , n21016 );
buf ( n21018 , n21017 );
and ( n21019 , n21018 , n19290 );
buf ( n21020 , n20540 );
buf ( n21021 , n21020 );
buf ( n21022 , n21021 );
and ( n21023 , n19219 , n21022 );
nor ( n21024 , n21019 , n21023 );
nand ( n21025 , n21002 , n21012 , n21024 );
nor ( n21026 , n20988 , n21025 );
not ( n21027 , n19631 );
not ( n21028 , n19385 );
and ( n21029 , n21027 , n21028 , n19377 );
not ( n21030 , n21029 );
or ( n21031 , n21026 , n21030 );
nand ( n21032 , n21030 , n18319 );
nand ( n21033 , n21031 , n21032 );
buf ( n21034 , n21033 );
buf ( n21035 , n21034 );
not ( n21036 , n275929 );
buf ( n21037 , n21036 );
buf ( n21038 , n21037 );
buf ( n21039 , n18208 );
buf ( n21040 , n19001 );
buf ( n21041 , n21040 );
not ( n21042 , n21041 );
buf ( n21043 , n18777 );
buf ( n21044 , n19439 );
nor ( n21045 , n21043 , n21044 );
buf ( n21046 , n21045 );
buf ( n21047 , n21046 );
buf ( n21048 , n19024 );
buf ( n21049 , n21048 );
nand ( n21050 , n21047 , n21049 );
buf ( n21051 , n21050 );
buf ( n21052 , n21051 );
not ( n21053 , n21052 );
buf ( n21054 , n21053 );
buf ( n21055 , n21054 );
buf ( n21056 , n19463 );
nand ( n21057 , n21055 , n21056 );
buf ( n21058 , n21057 );
buf ( n21059 , n21058 );
not ( n21060 , n21059 );
or ( n21061 , n21042 , n21060 );
buf ( n21062 , n19463 );
not ( n21063 , n21062 );
buf ( n21064 , n21063 );
buf ( n21065 , n21064 );
buf ( n21066 , n21051 );
nor ( n21067 , n21065 , n21066 );
buf ( n21068 , n21067 );
buf ( n21069 , n21068 );
buf ( n21070 , n21040 );
not ( n21071 , n21070 );
buf ( n21072 , n21071 );
buf ( n21073 , n21072 );
nand ( n21074 , n21069 , n21073 );
buf ( n21075 , n21074 );
buf ( n21076 , n21075 );
nand ( n21077 , n21061 , n21076 );
buf ( n21078 , n21077 );
buf ( n21079 , n21078 );
buf ( n21080 , n21079 );
and ( n21081 , n21039 , n21080 );
not ( n21082 , n21039 );
buf ( n21083 , n18710 );
buf ( n21084 , n21083 );
not ( n21085 , n21084 );
buf ( n21086 , n19460 );
not ( n21087 , n21086 );
buf ( n21088 , n21087 );
buf ( n21089 , n21088 );
buf ( n21090 , n21046 );
buf ( n21091 , n18735 );
buf ( n21092 , n21091 );
not ( n21093 , n21092 );
buf ( n21094 , n19027 );
nor ( n21095 , n21093 , n21094 );
buf ( n21096 , n21095 );
buf ( n21097 , n21096 );
and ( n21098 , n21090 , n21097 );
buf ( n21099 , n21098 );
buf ( n21100 , n21099 );
nand ( n21101 , n21089 , n21100 );
buf ( n21102 , n21101 );
buf ( n21103 , n21102 );
not ( n21104 , n21103 );
or ( n21105 , n21085 , n21104 );
buf ( n21106 , n21102 );
buf ( n21107 , n21083 );
or ( n21108 , n21106 , n21107 );
nand ( n21109 , n21105 , n21108 );
buf ( n21110 , n21109 );
buf ( n21111 , n21110 );
buf ( n21112 , n21111 );
buf ( n21113 , n21112 );
not ( n21114 , n21113 );
buf ( n21115 , n21079 );
and ( n21116 , n19603 , n21115 );
nand ( n21117 , n19620 , n19477 );
buf ( n21118 , n19460 );
not ( n21119 , n21118 );
buf ( n21120 , n21119 );
buf ( n21121 , n21120 );
buf ( n21122 , n21046 );
nand ( n21123 , n21121 , n21122 );
buf ( n21124 , n21123 );
buf ( n21125 , n21124 );
buf ( n21126 , n21048 );
not ( n21127 , n21126 );
buf ( n21128 , n21127 );
buf ( n21129 , n21128 );
and ( n21130 , n21125 , n21129 );
not ( n21131 , n21125 );
buf ( n21132 , n21048 );
and ( n21133 , n21131 , n21132 );
nor ( n21134 , n21130 , n21133 );
buf ( n21135 , n21134 );
buf ( n21136 , n21135 );
buf ( n21137 , n21136 );
nand ( n21138 , n21137 , n19474 );
nor ( n21139 , n21117 , n21138 );
nand ( n21140 , n21116 , n21139 );
not ( n21141 , n21140 );
buf ( n21142 , n21091 );
buf ( n21143 , n21142 );
not ( n21144 , n21143 );
buf ( n21145 , n21088 );
buf ( n21146 , n21046 );
buf ( n21147 , n19030 );
and ( n21148 , n21146 , n21147 );
buf ( n21149 , n21148 );
buf ( n21150 , n21149 );
nand ( n21151 , n21145 , n21150 );
buf ( n21152 , n21151 );
buf ( n21153 , n21152 );
not ( n21154 , n21153 );
or ( n21155 , n21144 , n21154 );
buf ( n21156 , n21152 );
buf ( n21157 , n21142 );
or ( n21158 , n21156 , n21157 );
nand ( n21159 , n21155 , n21158 );
buf ( n21160 , n21159 );
buf ( n21161 , n21160 );
buf ( n21162 , n21161 );
buf ( n21163 , n21162 );
nand ( n21164 , n19069 , n21141 , n21163 );
buf ( n21165 , n21164 );
not ( n21166 , n21165 );
or ( n21167 , n21114 , n21166 );
or ( n21168 , n21165 , n21113 );
nand ( n21169 , n21167 , n21168 );
buf ( n21170 , n21169 );
and ( n21171 , n21082 , n21170 );
nor ( n21172 , n21081 , n21171 );
not ( n21173 , n21172 );
buf ( n21174 , n20987 );
and ( n21175 , n21173 , n21174 );
not ( n21176 , n21001 );
not ( n21177 , n17912 );
not ( n21178 , n19235 );
or ( n21179 , n21177 , n21178 );
not ( n21180 , n277527 );
buf ( n21181 , n19690 );
buf ( n21182 , n9531 );
buf ( n21183 , n21182 );
buf ( n21184 , n21183 );
buf ( n21185 , n11512 );
buf ( n21186 , n21185 );
nor ( n21187 , n21184 , n21186 );
buf ( n21188 , n21187 );
buf ( n21189 , n21188 );
buf ( n21190 , n19873 );
nor ( n21191 , n21189 , n21190 );
buf ( n21192 , n21191 );
buf ( n21193 , n21192 );
and ( n21194 , n21181 , n21193 );
buf ( n21195 , n21194 );
buf ( n21196 , n21195 );
not ( n21197 , n21196 );
buf ( n21198 , n21197 );
buf ( n21199 , n21198 );
buf ( n21200 , n9540 );
buf ( n21201 , n21200 );
buf ( n21202 , n11452 );
buf ( n21203 , n21202 );
or ( n21204 , n21201 , n21203 );
buf ( n21205 , n21204 );
buf ( n21206 , n21205 );
buf ( n21207 , n9575 );
buf ( n21208 , n21207 );
buf ( n21209 , n11364 );
buf ( n21210 , n21209 );
or ( n21211 , n21208 , n21210 );
buf ( n21212 , n21211 );
buf ( n21213 , n21212 );
nand ( n21214 , n21206 , n21213 );
buf ( n21215 , n21214 );
buf ( n21216 , n21215 );
nor ( n21217 , n21199 , n21216 );
buf ( n21218 , n21217 );
buf ( n21219 , n21218 );
not ( n21220 , n21219 );
buf ( n21221 , n19835 );
not ( n21222 , n21221 );
or ( n21223 , n21220 , n21222 );
buf ( n21224 , n19854 );
buf ( n21225 , n21192 );
and ( n21226 , n21224 , n21225 );
buf ( n21227 , n21188 );
not ( n21228 , n21227 );
buf ( n21229 , n21228 );
buf ( n21230 , n21229 );
not ( n21231 , n21230 );
buf ( n21232 , n19867 );
not ( n21233 , n21232 );
or ( n21234 , n21231 , n21233 );
buf ( n21235 , n21183 );
buf ( n21236 , n21185 );
nand ( n21237 , n21235 , n21236 );
buf ( n21238 , n21237 );
buf ( n21239 , n21238 );
nand ( n21240 , n21234 , n21239 );
buf ( n21241 , n21240 );
buf ( n21242 , n21241 );
nor ( n21243 , n21226 , n21242 );
buf ( n21244 , n21243 );
buf ( n21245 , n21244 );
not ( n21246 , n21245 );
buf ( n21247 , n21246 );
buf ( n21248 , n21247 );
buf ( n21249 , n21215 );
not ( n21250 , n21249 );
buf ( n21251 , n21250 );
buf ( n21252 , n21251 );
and ( n21253 , n21248 , n21252 );
buf ( n21254 , n21205 );
buf ( n21255 , n21207 );
buf ( n21256 , n21209 );
and ( n21257 , n21255 , n21256 );
buf ( n21258 , n21257 );
buf ( n21259 , n21258 );
nand ( n21260 , n21254 , n21259 );
buf ( n21261 , n21260 );
buf ( n21262 , n21261 );
buf ( n21263 , n21200 );
buf ( n21264 , n21202 );
nand ( n21265 , n21263 , n21264 );
buf ( n21266 , n21265 );
buf ( n21267 , n21266 );
nand ( n21268 , n21262 , n21267 );
buf ( n21269 , n21268 );
buf ( n21270 , n21269 );
nor ( n21271 , n21253 , n21270 );
buf ( n21272 , n21271 );
buf ( n21273 , n21272 );
nand ( n21274 , n21223 , n21273 );
buf ( n21275 , n21274 );
buf ( n21276 , n21275 );
buf ( n21277 , n9558 );
buf ( n21278 , n21277 );
buf ( n21279 , n11236 );
buf ( n21280 , n21279 );
or ( n21281 , n21278 , n21280 );
buf ( n21282 , n21281 );
buf ( n21283 , n21282 );
buf ( n21284 , n21277 );
buf ( n21285 , n21279 );
and ( n21286 , n21284 , n21285 );
buf ( n21287 , n21286 );
buf ( n21288 , n21287 );
not ( n21289 , n21288 );
buf ( n21290 , n21289 );
buf ( n21291 , n21290 );
nand ( n21292 , n21283 , n21291 );
buf ( n21293 , n21292 );
buf ( n21294 , n21293 );
xnor ( n21295 , n21276 , n21294 );
buf ( n21296 , n21295 );
buf ( n21297 , n21296 );
not ( n21298 , n21297 );
or ( n21299 , n21180 , n21298 );
nand ( n21300 , n277351 , n9558 );
nand ( n21301 , n21299 , n21300 );
nand ( n21302 , n19242 , n21301 );
nand ( n21303 , n21179 , n21302 );
buf ( n21304 , n21303 );
not ( n21305 , n21304 );
not ( n21306 , n21305 );
buf ( n21307 , n18734 );
buf ( n21308 , n21307 );
not ( n21309 , n21308 );
not ( n21310 , n21309 );
or ( n21311 , n21306 , n21310 );
nand ( n21312 , n21308 , n21304 );
nand ( n21313 , n21311 , n21312 );
not ( n21314 , n17928 );
not ( n21315 , n19235 );
or ( n21316 , n21314 , n21315 );
not ( n21317 , n277527 );
buf ( n21318 , n21198 );
buf ( n21319 , n21212 );
not ( n21320 , n21319 );
buf ( n21321 , n21320 );
buf ( n21322 , n21321 );
nor ( n21323 , n21318 , n21322 );
buf ( n21324 , n21323 );
buf ( n21325 , n21324 );
not ( n21326 , n21325 );
buf ( n21327 , n19835 );
not ( n21328 , n21327 );
or ( n21329 , n21326 , n21328 );
buf ( n21330 , n21247 );
buf ( n21331 , n21212 );
and ( n21332 , n21330 , n21331 );
buf ( n21333 , n21258 );
nor ( n21334 , n21332 , n21333 );
buf ( n21335 , n21334 );
buf ( n21336 , n21335 );
nand ( n21337 , n21329 , n21336 );
buf ( n21338 , n21337 );
buf ( n21339 , n21338 );
buf ( n21340 , n21205 );
buf ( n21341 , n21266 );
nand ( n21342 , n21340 , n21341 );
buf ( n21343 , n21342 );
buf ( n21344 , n21343 );
xnor ( n21345 , n21339 , n21344 );
buf ( n21346 , n21345 );
buf ( n21347 , n21346 );
not ( n21348 , n21347 );
or ( n21349 , n21317 , n21348 );
nand ( n21350 , n277351 , n9540 );
nand ( n21351 , n21349 , n21350 );
nand ( n21352 , n19242 , n21351 );
nand ( n21353 , n21316 , n21352 );
buf ( n21354 , n21353 );
not ( n21355 , n21354 );
buf ( n21356 , n19000 );
buf ( n21357 , n21356 );
and ( n21358 , n21355 , n21357 );
nand ( n21359 , n21313 , n21358 );
not ( n21360 , n21359 );
not ( n21361 , n21360 );
nor ( n21362 , n21313 , n21358 );
not ( n21363 , n21362 );
nand ( n21364 , n21361 , n21363 );
not ( n21365 , n21364 );
buf ( n21366 , n18756 );
buf ( n21367 , n21366 );
not ( n21368 , n21367 );
not ( n21369 , n17895 );
not ( n21370 , n19235 );
or ( n21371 , n21369 , n21370 );
not ( n21372 , n277527 );
buf ( n21373 , n19690 );
buf ( n21374 , n19876 );
and ( n21375 , n21373 , n21374 );
buf ( n21376 , n21375 );
buf ( n21377 , n21376 );
not ( n21378 , n21377 );
buf ( n21379 , n19835 );
not ( n21380 , n21379 );
or ( n21381 , n21378 , n21380 );
buf ( n21382 , n19854 );
buf ( n21383 , n19876 );
and ( n21384 , n21382 , n21383 );
buf ( n21385 , n19867 );
nor ( n21386 , n21384 , n21385 );
buf ( n21387 , n21386 );
buf ( n21388 , n21387 );
nand ( n21389 , n21381 , n21388 );
buf ( n21390 , n21389 );
buf ( n21391 , n21390 );
buf ( n21392 , n21229 );
buf ( n21393 , n21238 );
nand ( n21394 , n21392 , n21393 );
buf ( n21395 , n21394 );
buf ( n21396 , n21395 );
xnor ( n21397 , n21391 , n21396 );
buf ( n21398 , n21397 );
buf ( n21399 , n21398 );
not ( n21400 , n21399 );
or ( n21401 , n21372 , n21400 );
nand ( n21402 , n277351 , n21182 );
nand ( n21403 , n21401 , n21402 );
nand ( n21404 , n19242 , n21403 );
nand ( n21405 , n21371 , n21404 );
buf ( n21406 , n21405 );
not ( n21407 , n21406 );
or ( n21408 , n21368 , n21407 );
not ( n21409 , n21367 );
not ( n21410 , n21406 );
nand ( n21411 , n21409 , n21410 );
nand ( n21412 , n21408 , n21411 );
and ( n21413 , n19894 , n19669 );
nor ( n21414 , n21412 , n21413 );
nor ( n21415 , n19940 , n21414 );
buf ( n21416 , n21415 );
nand ( n21417 , n20071 , n21416 );
buf ( n21418 , n19023 );
buf ( n21419 , n21418 );
not ( n21420 , n21419 );
not ( n21421 , n21420 );
not ( n21422 , n17942 );
not ( n21423 , n19235 );
or ( n21424 , n21422 , n21423 );
not ( n21425 , n9432 );
buf ( n21426 , n21195 );
not ( n21427 , n21426 );
buf ( n21428 , n19835 );
not ( n21429 , n21428 );
or ( n21430 , n21427 , n21429 );
buf ( n21431 , n21244 );
nand ( n21432 , n21430 , n21431 );
buf ( n21433 , n21432 );
buf ( n21434 , n21433 );
buf ( n21435 , n21258 );
buf ( n21436 , n21321 );
nor ( n21437 , n21435 , n21436 );
buf ( n21438 , n21437 );
buf ( n21439 , n21438 );
xor ( n21440 , n21434 , n21439 );
buf ( n21441 , n21440 );
buf ( n21442 , n21441 );
not ( n21443 , n21442 );
or ( n21444 , n21425 , n21443 );
nand ( n21445 , n9433 , n9575 );
nand ( n21446 , n21444 , n21445 );
nand ( n21447 , n19242 , n21446 );
nand ( n21448 , n21424 , n21447 );
buf ( n21449 , n21448 );
not ( n21450 , n21449 );
not ( n21451 , n21450 );
or ( n21452 , n21421 , n21451 );
nand ( n21453 , n21449 , n21419 );
nand ( n21454 , n21452 , n21453 );
nand ( n21455 , n21410 , n21367 );
not ( n21456 , n21455 );
nor ( n21457 , n21454 , n21456 );
not ( n21458 , n21457 );
not ( n21459 , n21355 );
not ( n21460 , n21357 );
not ( n21461 , n21460 );
or ( n21462 , n21459 , n21461 );
nand ( n21463 , n21357 , n21354 );
nand ( n21464 , n21462 , n21463 );
nand ( n21465 , n21450 , n21419 );
not ( n21466 , n21465 );
nor ( n21467 , n21464 , n21466 );
not ( n21468 , n21467 );
nand ( n21469 , n21458 , n21468 );
nor ( n21470 , n21417 , n21469 );
not ( n21471 , n21470 );
not ( n21472 , n20337 );
or ( n21473 , n21471 , n21472 );
not ( n21474 , n21469 );
not ( n21475 , n21474 );
not ( n21476 , n21416 );
not ( n21477 , n20345 );
or ( n21478 , n21476 , n21477 );
or ( n21479 , n21414 , n19942 );
buf ( n21480 , n21412 );
buf ( n21481 , n21413 );
nand ( n21482 , n21480 , n21481 );
nand ( n21483 , n21479 , n21482 );
not ( n21484 , n21483 );
nand ( n21485 , n21478 , n21484 );
not ( n21486 , n21485 );
or ( n21487 , n21475 , n21486 );
nand ( n21488 , n21454 , n21456 );
nand ( n21489 , n21464 , n21466 );
nand ( n21490 , n21488 , n21489 );
nand ( n21491 , n21490 , n21468 );
nand ( n21492 , n21487 , n21491 );
not ( n21493 , n21492 );
nand ( n21494 , n21473 , n21493 );
not ( n21495 , n21494 );
or ( n21496 , n21365 , n21495 );
or ( n21497 , n21494 , n21364 );
nand ( n21498 , n21496 , n21497 );
buf ( n21499 , n21498 );
not ( n21500 , n21499 );
or ( n21501 , n21176 , n21500 );
buf ( n21502 , n21303 );
not ( n21503 , n21502 );
buf ( n21504 , n21307 );
not ( n21505 , n21504 );
not ( n21506 , n21505 );
or ( n21507 , n21503 , n21506 );
not ( n21508 , n21502 );
nand ( n21509 , n21508 , n21504 );
nand ( n21510 , n21507 , n21509 );
buf ( n21511 , n21353 );
buf ( n21512 , n21356 );
and ( n21513 , n21511 , n21512 );
nor ( n21514 , n21510 , n21513 );
not ( n21515 , n21514 );
buf ( n21516 , n21510 );
buf ( n21517 , n21513 );
nand ( n21518 , n21516 , n21517 );
nand ( n21519 , n21515 , n21518 );
not ( n21520 , n21519 );
not ( n21521 , n21512 );
not ( n21522 , n21521 );
not ( n21523 , n21511 );
or ( n21524 , n21522 , n21523 );
not ( n21525 , n21511 );
nand ( n21526 , n21525 , n21512 );
nand ( n21527 , n21524 , n21526 );
not ( n21528 , n21527 );
buf ( n21529 , n21448 );
buf ( n21530 , n21418 );
and ( n21531 , n21529 , n21530 );
not ( n21532 , n21531 );
nand ( n21533 , n21528 , n21532 );
not ( n21534 , n21533 );
not ( n21535 , n21530 );
not ( n21536 , n21529 );
not ( n21537 , n21536 );
or ( n21538 , n21535 , n21537 );
not ( n21539 , n21530 );
nand ( n21540 , n21539 , n21529 );
nand ( n21541 , n21538 , n21540 );
buf ( n21542 , n21366 );
buf ( n21543 , n21405 );
nand ( n21544 , n21542 , n21543 );
not ( n21545 , n21544 );
nor ( n21546 , n21541 , n21545 );
nor ( n21547 , n21534 , n21546 );
not ( n21548 , n21547 );
not ( n21549 , n21543 );
not ( n21550 , n21549 );
not ( n21551 , n21542 );
or ( n21552 , n21550 , n21551 );
not ( n21553 , n21542 );
nand ( n21554 , n21553 , n21543 );
nand ( n21555 , n21552 , n21554 );
not ( n21556 , n21555 );
not ( n21557 , n20356 );
nor ( n21558 , n21557 , n20362 );
not ( n21559 , n21558 );
nand ( n21560 , n21556 , n21559 );
nand ( n21561 , n21560 , n20369 );
nor ( n21562 , n21561 , n20401 );
not ( n21563 , n21562 );
nor ( n21564 , n21548 , n21563 );
not ( n21565 , n21564 );
not ( n21566 , n20500 );
or ( n21567 , n21565 , n21566 );
nand ( n21568 , n20372 , n20506 );
or ( n21569 , n20505 , n21568 );
not ( n21570 , n21561 );
nand ( n21571 , n21569 , n21570 );
not ( n21572 , n21559 );
buf ( n21573 , n21555 );
nand ( n21574 , n21572 , n21573 );
nand ( n21575 , n21571 , n21574 );
buf ( n21576 , n21575 );
and ( n21577 , n21547 , n21576 );
and ( n21578 , n21541 , n21545 );
not ( n21579 , n21578 );
not ( n21580 , n21533 );
or ( n21581 , n21579 , n21580 );
not ( n21582 , n21532 );
buf ( n21583 , n21527 );
nand ( n21584 , n21582 , n21583 );
nand ( n21585 , n21581 , n21584 );
nor ( n21586 , n21577 , n21585 );
nand ( n21587 , n21567 , n21586 );
not ( n21588 , n21587 );
or ( n21589 , n21520 , n21588 );
or ( n21590 , n21587 , n21519 );
nand ( n21591 , n21589 , n21590 );
buf ( n21592 , n21591 );
and ( n21593 , n21592 , n19358 );
not ( n21594 , n19290 );
buf ( n21595 , n21303 );
buf ( n21596 , n21595 );
not ( n21597 , n21596 );
not ( n21598 , n21597 );
not ( n21599 , n20551 );
not ( n21600 , n20549 );
buf ( n21601 , n21405 );
buf ( n21602 , n21601 );
not ( n21603 , n21602 );
nand ( n21604 , n21599 , n21600 , n20521 , n21603 );
buf ( n21605 , n21604 );
not ( n21606 , n21605 );
buf ( n21607 , n21353 );
buf ( n21608 , n21607 );
buf ( n21609 , n21448 );
buf ( n21610 , n21609 );
nor ( n21611 , n21608 , n21610 );
and ( n21612 , n21606 , n21611 );
nand ( n21613 , n21612 , n20547 );
not ( n21614 , n21613 );
or ( n21615 , n21598 , n21614 );
or ( n21616 , n21613 , n21597 );
nand ( n21617 , n21615 , n21616 );
buf ( n21618 , n21617 );
not ( n21619 , n21618 );
or ( n21620 , n21594 , n21619 );
buf ( n21621 , n21595 );
buf ( n21622 , n21621 );
buf ( n21623 , n21622 );
buf ( n21624 , n21623 );
nand ( n21625 , n19219 , n21624 );
nand ( n21626 , n21620 , n21625 );
nor ( n21627 , n21593 , n21626 );
nand ( n21628 , n21501 , n21627 );
nor ( n21629 , n21175 , n21628 );
or ( n21630 , n21629 , n21030 );
nand ( n21631 , n21030 , n18726 );
nand ( n21632 , n21630 , n21631 );
buf ( n21633 , n21632 );
buf ( n21634 , n21633 );
buf ( n21635 , n275554 );
not ( n21636 , n275550 );
buf ( n21637 , n21636 );
buf ( n21638 , n21637 );
not ( n21639 , n275550 );
buf ( n21640 , n21639 );
buf ( n21641 , n21640 );
not ( n21642 , n275929 );
buf ( n21643 , n21642 );
buf ( n21644 , n21643 );
and ( n21645 , n20711 , n16705 );
not ( n21646 , n20711 );
buf ( n21647 , n14565 );
not ( n21648 , n21647 );
nand ( n21649 , n14778 , n14543 );
buf ( n21650 , n21649 );
not ( n21651 , n21650 );
or ( n21652 , n21648 , n21651 );
or ( n21653 , n21650 , n21647 );
nand ( n21654 , n21652 , n21653 );
buf ( n21655 , n21654 );
and ( n21656 , n21646 , n21655 );
nor ( n21657 , n21645 , n21656 );
not ( n21658 , n21657 );
not ( n21659 , n20846 );
and ( n21660 , n21658 , n21659 );
not ( n21661 , n20926 );
not ( n21662 , n17297 );
not ( n21663 , n21662 );
not ( n21664 , n17292 );
or ( n21665 , n21663 , n21664 );
or ( n21666 , n17292 , n21662 );
nand ( n21667 , n21665 , n21666 );
buf ( n21668 , n21667 );
not ( n21669 , n21668 );
or ( n21670 , n21661 , n21669 );
not ( n21671 , n16724 );
not ( n21672 , n21671 );
nand ( n21673 , n16727 , n16707 );
not ( n21674 , n21673 );
or ( n21675 , n21672 , n21674 );
or ( n21676 , n21673 , n21671 );
nand ( n21677 , n21675 , n21676 );
buf ( n21678 , n21677 );
and ( n21679 , n21678 , n20889 );
xor ( n21680 , n17424 , n17425 );
buf ( n21681 , n21680 );
and ( n21682 , n21681 , n17409 );
buf ( n21683 , n16695 );
buf ( n21684 , n21683 );
buf ( n21685 , n21684 );
and ( n21686 , n17499 , n21685 );
nor ( n21687 , n21682 , n21686 );
not ( n21688 , n21687 );
nor ( n21689 , n21679 , n21688 );
nand ( n21690 , n21670 , n21689 );
nor ( n21691 , n21660 , n21690 );
not ( n21692 , n16965 );
not ( n21693 , n14841 );
nand ( n21694 , n21693 , n14867 );
nor ( n21695 , n21692 , n21694 );
nand ( n21696 , n21695 , n17558 );
buf ( n21697 , n21696 );
or ( n21698 , n21691 , n21697 );
nand ( n21699 , n21696 , n14535 );
nand ( n21700 , n21698 , n21699 );
buf ( n21701 , n21700 );
buf ( n21702 , n21701 );
not ( n21703 , n275550 );
buf ( n21704 , n21703 );
buf ( n21705 , n21704 );
buf ( n21706 , n18923 );
not ( n21707 , n21706 );
buf ( n21708 , n18738 );
buf ( n21709 , n19027 );
nor ( n21710 , n21708 , n21709 );
buf ( n21711 , n21710 );
buf ( n21712 , n21711 );
buf ( n21713 , n18757 );
buf ( n21714 , n18774 );
nand ( n21715 , n21713 , n21714 );
buf ( n21716 , n21715 );
buf ( n21717 , n21716 );
buf ( n21718 , n18418 );
nor ( n21719 , n21717 , n21718 );
buf ( n21720 , n21719 );
buf ( n21721 , n21720 );
nand ( n21722 , n21707 , n21712 , n21721 );
buf ( n21723 , n21722 );
buf ( n21724 , n21723 );
not ( n21725 , n21724 );
buf ( n21726 , n21725 );
buf ( n21727 , n21726 );
buf ( n21728 , n18975 );
buf ( n21729 , n18632 );
nor ( n21730 , n21728 , n21729 );
buf ( n21731 , n21730 );
buf ( n21732 , n21731 );
not ( n21733 , n21732 );
buf ( n21734 , n21733 );
buf ( n21735 , n21734 );
buf ( n21736 , n18684 );
buf ( n21737 , n21736 );
not ( n21738 , n21737 );
buf ( n21739 , n21738 );
buf ( n21740 , n21739 );
nor ( n21741 , n21735 , n21740 );
buf ( n21742 , n21741 );
buf ( n21743 , n21742 );
nand ( n21744 , n21727 , n21743 );
buf ( n21745 , n21744 );
buf ( n21746 , n21745 );
buf ( n21747 , n18834 );
buf ( n21748 , n21747 );
not ( n21749 , n21748 );
buf ( n21750 , n21749 );
buf ( n21751 , n21750 );
and ( n21752 , n21746 , n21751 );
not ( n21753 , n21746 );
buf ( n21754 , n21747 );
and ( n21755 , n21753 , n21754 );
nor ( n21756 , n21752 , n21755 );
buf ( n21757 , n21756 );
buf ( n21758 , n21757 );
not ( n21759 , n21758 );
not ( n21760 , n21759 );
not ( n21761 , n21760 );
not ( n21762 , n19119 );
buf ( n21763 , n275556 );
not ( n21764 , n21763 );
nor ( n21765 , n21762 , n21764 );
nand ( n21766 , n19132 , n21765 );
not ( n21767 , n19140 );
nand ( n21768 , n21767 , n19124 );
or ( n21769 , n21766 , n21768 );
buf ( n21770 , n21769 );
or ( n21771 , n21761 , n21770 );
not ( n21772 , n21769 );
not ( n21773 , n21772 );
buf ( n21774 , n21773 );
nand ( n21775 , n21774 , n9671 );
nand ( n21776 , n21771 , n21775 );
buf ( n21777 , n21776 );
buf ( n21778 , n21777 );
buf ( n21779 , n275554 );
not ( n21780 , n275925 );
buf ( n21781 , n21780 );
buf ( n21782 , n21781 );
buf ( n21783 , n275554 );
not ( n21784 , n275550 );
buf ( n21785 , n21784 );
buf ( n21786 , n21785 );
not ( n21787 , n275550 );
buf ( n21788 , n21787 );
buf ( n21789 , n21788 );
not ( n21790 , n275550 );
buf ( n21791 , n21790 );
buf ( n21792 , n21791 );
buf ( n21793 , n275554 );
buf ( n21794 , n10772 );
buf ( n21795 , n21794 );
buf ( n21796 , n10739 );
buf ( n21797 , n21796 );
or ( n21798 , n21795 , n21797 );
buf ( n21799 , n21798 );
buf ( n21800 , n21799 );
not ( n21801 , n21800 );
buf ( n21802 , n21801 );
buf ( n21803 , n21802 );
not ( n21804 , n21803 );
buf ( n21805 , n21804 );
buf ( n21806 , n21805 );
not ( n21807 , n21806 );
buf ( n21808 , n10893 );
buf ( n21809 , n21808 );
buf ( n21810 , n10860 );
buf ( n21811 , n21810 );
and ( n21812 , n21809 , n21811 );
buf ( n21813 , n21812 );
buf ( n21814 , n21813 );
not ( n21815 , n21814 );
buf ( n21816 , n10921 );
not ( n21817 , n21816 );
buf ( n21818 , n21817 );
buf ( n21819 , n21818 );
buf ( n21820 , n10960 );
buf ( n21821 , n21820 );
not ( n21822 , n21821 );
buf ( n21823 , n21822 );
buf ( n21824 , n21823 );
nand ( n21825 , n21819 , n21824 );
buf ( n21826 , n21825 );
buf ( n21827 , n21826 );
not ( n21828 , n21827 );
or ( n21829 , n21815 , n21828 );
buf ( n21830 , n21818 );
not ( n21831 , n21830 );
buf ( n21832 , n21831 );
buf ( n21833 , n21832 );
buf ( n21834 , n21823 );
not ( n21835 , n21834 );
buf ( n21836 , n21835 );
buf ( n21837 , n21836 );
nand ( n21838 , n21833 , n21837 );
buf ( n21839 , n21838 );
buf ( n21840 , n21839 );
nand ( n21841 , n21829 , n21840 );
buf ( n21842 , n21841 );
buf ( n21843 , n21842 );
not ( n21844 , n21843 );
or ( n21845 , n21807 , n21844 );
buf ( n21846 , n21794 );
buf ( n21847 , n21796 );
and ( n21848 , n21846 , n21847 );
buf ( n21849 , n21848 );
buf ( n21850 , n21849 );
not ( n21851 , n21850 );
buf ( n21852 , n21851 );
buf ( n21853 , n21852 );
nand ( n21854 , n21845 , n21853 );
buf ( n21855 , n21854 );
buf ( n21856 , n21855 );
not ( n21857 , n21856 );
buf ( n21858 , n11097 );
buf ( n21859 , n21858 );
not ( n21860 , n21859 );
buf ( n21861 , n21860 );
buf ( n21862 , n21861 );
buf ( n21863 , n11122 );
buf ( n21864 , n21863 );
not ( n21865 , n21864 );
buf ( n21866 , n21865 );
buf ( n21867 , n21866 );
nand ( n21868 , n21862 , n21867 );
buf ( n21869 , n21868 );
buf ( n21870 , n21869 );
not ( n21871 , n21870 );
buf ( n21872 , n21858 );
buf ( n21873 , n21863 );
nand ( n21874 , n21872 , n21873 );
buf ( n21875 , n21874 );
buf ( n21876 , n21875 );
buf ( n21877 , n11141 );
buf ( n21878 , n21877 );
buf ( n21879 , n11161 );
buf ( n21880 , n21879 );
nand ( n21881 , n21878 , n21880 );
buf ( n21882 , n21881 );
buf ( n21883 , n21882 );
nand ( n21884 , n21876 , n21883 );
buf ( n21885 , n21884 );
buf ( n21886 , n21885 );
not ( n21887 , n21886 );
or ( n21888 , n21871 , n21887 );
buf ( n21889 , n21879 );
not ( n21890 , n21889 );
buf ( n21891 , n21890 );
buf ( n21892 , n21891 );
buf ( n21893 , n21877 );
not ( n21894 , n21893 );
buf ( n21895 , n21894 );
buf ( n21896 , n21895 );
nand ( n21897 , n21892 , n21896 );
buf ( n21898 , n21897 );
buf ( n21899 , n21898 );
buf ( n21900 , n21899 );
buf ( n21901 , n11045 );
buf ( n21902 , n21901 );
buf ( n21903 , n11062 );
buf ( n21904 , n21903 );
nand ( n21905 , n21902 , n21904 );
buf ( n21906 , n21905 );
buf ( n21907 , n21906 );
not ( n21908 , n21907 );
buf ( n21909 , n21908 );
buf ( n21910 , n21909 );
not ( n21911 , n21910 );
buf ( n21912 , n11009 );
buf ( n21913 , n21912 );
not ( n21914 , n21913 );
buf ( n21915 , n10984 );
buf ( n21916 , n21915 );
not ( n21917 , n21916 );
buf ( n21918 , n21917 );
buf ( n21919 , n21918 );
nand ( n21920 , n21914 , n21919 );
buf ( n21921 , n21920 );
buf ( n21922 , n21921 );
not ( n21923 , n21922 );
or ( n21924 , n21911 , n21923 );
buf ( n21925 , n21912 );
buf ( n21926 , n21915 );
nand ( n21927 , n21925 , n21926 );
buf ( n21928 , n21927 );
buf ( n21929 , n21928 );
nand ( n21930 , n21924 , n21929 );
buf ( n21931 , n21930 );
buf ( n21932 , n21931 );
buf ( n21933 , n21869 );
nand ( n21934 , n21900 , n21932 , n21933 );
buf ( n21935 , n21934 );
buf ( n21936 , n21935 );
nand ( n21937 , n21888 , n21936 );
buf ( n21938 , n21937 );
buf ( n21939 , n21938 );
buf ( n21940 , n21826 );
buf ( n21941 , n21940 );
buf ( n21942 , n21808 );
buf ( n21943 , n21810 );
or ( n21944 , n21942 , n21943 );
buf ( n21945 , n21944 );
buf ( n21946 , n21945 );
nand ( n21947 , n21941 , n21946 );
buf ( n21948 , n21947 );
buf ( n21949 , n21948 );
buf ( n21950 , n21802 );
nor ( n21951 , n21949 , n21950 );
buf ( n21952 , n21951 );
buf ( n21953 , n21952 );
nand ( n21954 , n21939 , n21953 );
buf ( n21955 , n21954 );
buf ( n21956 , n21955 );
nand ( n21957 , n21857 , n21956 );
buf ( n21958 , n21957 );
buf ( n21959 , n21958 );
buf ( n21960 , n10805 );
buf ( n21961 , n21960 );
not ( n21962 , n21961 );
buf ( n21963 , n10834 );
buf ( n21964 , n21963 );
not ( n21965 , n21964 );
buf ( n21966 , n21965 );
buf ( n21967 , n21966 );
nand ( n21968 , n21962 , n21967 );
buf ( n21969 , n21968 );
buf ( n21970 , n21969 );
buf ( n21971 , n21970 );
buf ( n21972 , n21966 );
not ( n21973 , n21972 );
buf ( n21974 , n21960 );
nand ( n21975 , n21973 , n21974 );
buf ( n21976 , n21975 );
buf ( n21977 , n21976 );
nand ( n21978 , n21971 , n21977 );
buf ( n21979 , n21978 );
buf ( n21980 , n21979 );
not ( n21981 , n21980 );
buf ( n21982 , n21981 );
buf ( n21983 , n21982 );
and ( n21984 , n21959 , n21983 );
not ( n21985 , n21959 );
buf ( n21986 , n21979 );
and ( n21987 , n21985 , n21986 );
nor ( n21988 , n21984 , n21987 );
buf ( n21989 , n21988 );
buf ( n21990 , n21989 );
not ( n21991 , n9152 );
or ( n21992 , n11728 , n21991 );
nand ( n21993 , n9130 , n12096 );
nand ( n21994 , n21992 , n21993 );
not ( n21995 , n9135 );
not ( n21996 , n9130 );
or ( n21997 , n21995 , n21996 );
nand ( n21998 , n21997 , n12686 );
buf ( n21999 , n21998 );
nor ( n22000 , n21994 , n21999 );
not ( n22001 , n22000 );
not ( n22002 , n22001 );
and ( n22003 , n21990 , n22002 );
and ( n22004 , n20581 , n20587 );
not ( n22005 , n9154 );
nand ( n22006 , n22004 , n22005 );
not ( n22007 , n22006 );
not ( n22008 , n22007 );
or ( n22009 , n22008 , n12340 );
not ( n22010 , n12686 );
nand ( n22011 , n22010 , n12679 );
buf ( n22012 , n22011 );
not ( n22013 , n22012 );
not ( n22014 , n22013 );
or ( n22015 , n22014 , n12128 );
nand ( n22016 , n22009 , n22015 );
nor ( n22017 , n22003 , n22016 );
buf ( n22018 , n10893 );
buf ( n22019 , n11010 );
nand ( n22020 , n22018 , n22019 );
buf ( n22021 , n11141 );
buf ( n22022 , n11097 );
nand ( n22023 , n22021 , n22022 );
nor ( n22024 , n22020 , n22023 );
not ( n22025 , n9366 );
nand ( n22026 , n22025 , n9372 );
not ( n22027 , n22026 );
not ( n22028 , n9399 );
or ( n22029 , n22027 , n22028 );
buf ( n22030 , n11045 );
nand ( n22031 , n22029 , n22030 );
not ( n22032 , n22031 );
buf ( n22033 , n22032 );
nand ( n22034 , n22024 , n22033 );
buf ( n22035 , n10773 );
buf ( n22036 , n10921 );
nand ( n22037 , n22035 , n22036 );
nor ( n22038 , n22034 , n22037 );
buf ( n22039 , n10806 );
not ( n22040 , n22039 );
not ( n22041 , n22040 );
nand ( n22042 , n22038 , n22041 );
buf ( n22043 , n11619 );
not ( n22044 , n22043 );
and ( n22045 , n22042 , n22044 );
not ( n22046 , n22042 );
and ( n22047 , n22046 , n22043 );
nor ( n22048 , n22045 , n22047 );
buf ( n22049 , n22048 );
not ( n22050 , n22004 );
nand ( n22051 , n22050 , n9155 );
not ( n22052 , n22051 );
nand ( n22053 , n22049 , n22052 );
not ( n22054 , n21998 );
nand ( n22055 , n22054 , n21994 );
buf ( n22056 , n22055 );
not ( n22057 , n22056 );
buf ( n22058 , n10806 );
not ( n22059 , n22058 );
not ( n22060 , n10835 );
buf ( n22061 , n22060 );
nand ( n22062 , n22059 , n22061 );
not ( n22063 , n22062 );
not ( n22064 , n22063 );
not ( n22065 , n22061 );
not ( n22066 , n22059 );
nand ( n22067 , n22065 , n22066 );
nand ( n22068 , n22064 , n22067 );
not ( n22069 , n22068 );
buf ( n22070 , n10773 );
not ( n22071 , n22070 );
buf ( n22072 , n10739 );
nand ( n22073 , n22071 , n22072 );
buf ( n22074 , n22073 );
not ( n22075 , n22074 );
buf ( n22076 , n10893 );
buf ( n22077 , n10860 );
not ( n22078 , n22077 );
and ( n22079 , n22076 , n22078 );
not ( n22080 , n22079 );
buf ( n22081 , n10921 );
not ( n22082 , n22081 );
buf ( n22083 , n10961 );
nand ( n22084 , n22082 , n22083 );
not ( n22085 , n22084 );
or ( n22086 , n22080 , n22085 );
not ( n22087 , n22083 );
nand ( n22088 , n22087 , n22081 );
nand ( n22089 , n22086 , n22088 );
not ( n22090 , n22089 );
or ( n22091 , n22075 , n22090 );
not ( n22092 , n22072 );
and ( n22093 , n22070 , n22092 );
not ( n22094 , n22093 );
nand ( n22095 , n22091 , n22094 );
not ( n22096 , n22095 );
buf ( n22097 , n11097 );
not ( n22098 , n22097 );
buf ( n22099 , n11122 );
nand ( n22100 , n22098 , n22099 );
not ( n22101 , n22100 );
buf ( n22102 , n11161 );
not ( n22103 , n22102 );
buf ( n22104 , n11141 );
nand ( n22105 , n22103 , n22104 );
not ( n22106 , n22099 );
nand ( n22107 , n22106 , n22097 );
nand ( n22108 , n22105 , n22107 );
not ( n22109 , n22108 );
or ( n22110 , n22101 , n22109 );
buf ( n22111 , n11009 );
not ( n22112 , n22111 );
buf ( n22113 , n10984 );
nand ( n22114 , n22112 , n22113 );
not ( n22115 , n22114 );
buf ( n22116 , n11045 );
not ( n22117 , n22116 );
buf ( n22118 , n11062 );
nand ( n22119 , n22117 , n22118 );
not ( n22120 , n22119 );
or ( n22121 , n22115 , n22120 );
not ( n22122 , n22113 );
nand ( n22123 , n22122 , n22111 );
nand ( n22124 , n22121 , n22123 );
not ( n22125 , n22104 );
nand ( n22126 , n22125 , n22102 );
nand ( n22127 , n22124 , n22126 , n22100 );
nand ( n22128 , n22110 , n22127 );
buf ( n22129 , n22128 );
not ( n22130 , n22076 );
nand ( n22131 , n22130 , n22077 );
nand ( n22132 , n22084 , n22131 );
not ( n22133 , n22074 );
nor ( n22134 , n22132 , n22133 );
nand ( n22135 , n22129 , n22134 );
nand ( n22136 , n22096 , n22135 );
not ( n22137 , n22136 );
or ( n22138 , n22069 , n22137 );
or ( n22139 , n22136 , n22068 );
nand ( n22140 , n22138 , n22139 );
buf ( n22141 , n22140 );
nand ( n22142 , n22057 , n22141 );
and ( n22143 , n22017 , n22053 , n22142 );
nor ( n22144 , n20643 , n9100 );
buf ( n22145 , n22144 );
buf ( n22146 , n22145 );
not ( n22147 , n9088 );
not ( n22148 , n9099 );
not ( n22149 , n22148 );
and ( n22150 , n22147 , n22149 );
nand ( n22151 , n9099 , n9162 );
nor ( n22152 , n9094 , n22151 );
nor ( n22153 , n22150 , n22152 );
nand ( n22154 , n22148 , n9163 );
nor ( n22155 , n9094 , n22154 );
nand ( n22156 , n9088 , n22155 );
buf ( n22157 , RI21077000_517);
not ( n22158 , n22157 );
not ( n22159 , n22158 );
nand ( n22160 , n22159 , n9088 );
nand ( n22161 , n22153 , n22156 , n22160 );
not ( n22162 , n22161 );
nand ( n22163 , n20613 , n9094 );
buf ( n22164 , RI21076538_518);
not ( n22165 , n22164 );
not ( n22166 , n22165 );
or ( n22167 , n22152 , n22166 );
nand ( n22168 , n22167 , n9088 );
nand ( n22169 , n22156 , n22163 , n22168 );
not ( n22170 , n22169 );
nand ( n22171 , n22146 , n22162 , n22170 );
not ( n22172 , n22171 );
not ( n22173 , n22172 );
not ( n22174 , n12686 );
not ( n22175 , n12376 );
or ( n22176 , n22174 , n22175 );
nand ( n22177 , n22176 , n12097 );
not ( n22178 , n12686 );
not ( n22179 , n9152 );
and ( n22180 , n22178 , n22179 );
nor ( n22181 , n22180 , n12111 );
nand ( n22182 , n12377 , n12105 );
nand ( n22183 , n12377 , n12108 );
nand ( n22184 , n22177 , n22181 , n22182 , n22183 );
not ( n22185 , n22184 );
or ( n22186 , n22173 , n22185 );
and ( n22187 , n22144 , n22161 );
nand ( n22188 , n22187 , n22169 );
not ( n22189 , n22188 );
nand ( n22190 , n12380 , n22189 );
nand ( n22191 , n22186 , n22190 );
buf ( n22192 , n22191 );
not ( n22193 , n22192 );
or ( n22194 , n22143 , n22193 );
not ( n22195 , n10795 );
or ( n22196 , n22192 , n22195 );
nand ( n22197 , n22194 , n22196 );
buf ( n22198 , n22197 );
buf ( n22199 , n22198 );
buf ( n22200 , n275554 );
not ( n22201 , n9433 );
buf ( n22202 , n15013 );
buf ( n22203 , n9744 );
buf ( n22204 , n22203 );
buf ( n22205 , n277605 );
buf ( n22206 , n22205 );
nor ( n22207 , n22204 , n22206 );
buf ( n22208 , n22207 );
buf ( n22209 , n22208 );
buf ( n22210 , n9752 );
buf ( n22211 , n22210 );
buf ( n22212 , n277529 );
buf ( n22213 , n22212 );
nor ( n22214 , n22211 , n22213 );
buf ( n22215 , n22214 );
buf ( n22216 , n22215 );
nor ( n22217 , n22209 , n22216 );
buf ( n22218 , n22217 );
buf ( n22219 , n22218 );
buf ( n22220 , n14927 );
buf ( n22221 , n15020 );
and ( n22222 , n22220 , n22221 );
buf ( n22223 , n22222 );
buf ( n22224 , n22223 );
and ( n22225 , n22219 , n22224 );
buf ( n22226 , n22225 );
buf ( n22227 , n22226 );
buf ( n22228 , n9787 );
buf ( n22229 , n22228 );
buf ( n22230 , n277408 );
buf ( n22231 , n22230 );
or ( n22232 , n22229 , n22231 );
buf ( n22233 , n22232 );
buf ( n22234 , n22233 );
and ( n22235 , n22227 , n22234 );
buf ( n22236 , n22235 );
buf ( n22237 , n22236 );
and ( n22238 , n22202 , n22237 );
buf ( n22239 , n22238 );
buf ( n22240 , n22239 );
not ( n22241 , n22240 );
buf ( n22242 , n15386 );
not ( n22243 , n22242 );
or ( n22244 , n22241 , n22243 );
buf ( n22245 , n15481 );
buf ( n22246 , n22236 );
and ( n22247 , n22245 , n22246 );
buf ( n22248 , n22233 );
not ( n22249 , n22248 );
buf ( n22250 , n14927 );
not ( n22251 , n22250 );
buf ( n22252 , n15488 );
not ( n22253 , n22252 );
or ( n22254 , n22251 , n22253 );
buf ( n22255 , n14932 );
nand ( n22256 , n22254 , n22255 );
buf ( n22257 , n22256 );
buf ( n22258 , n22257 );
not ( n22259 , n22258 );
buf ( n22260 , n22218 );
not ( n22261 , n22260 );
or ( n22262 , n22259 , n22261 );
buf ( n22263 , n22208 );
not ( n22264 , n22263 );
buf ( n22265 , n22210 );
buf ( n22266 , n22212 );
nand ( n22267 , n22265 , n22266 );
buf ( n22268 , n22267 );
buf ( n22269 , n22268 );
not ( n22270 , n22269 );
and ( n22271 , n22264 , n22270 );
buf ( n22272 , n22203 );
buf ( n22273 , n22205 );
and ( n22274 , n22272 , n22273 );
buf ( n22275 , n22274 );
buf ( n22276 , n22275 );
nor ( n22277 , n22271 , n22276 );
buf ( n22278 , n22277 );
buf ( n22279 , n22278 );
nand ( n22280 , n22262 , n22279 );
buf ( n22281 , n22280 );
buf ( n22282 , n22281 );
not ( n22283 , n22282 );
or ( n22284 , n22249 , n22283 );
buf ( n22285 , n22228 );
buf ( n22286 , n22230 );
nand ( n22287 , n22285 , n22286 );
buf ( n22288 , n22287 );
buf ( n22289 , n22288 );
nand ( n22290 , n22284 , n22289 );
buf ( n22291 , n22290 );
buf ( n22292 , n22291 );
nor ( n22293 , n22247 , n22292 );
buf ( n22294 , n22293 );
buf ( n22295 , n22294 );
nand ( n22296 , n22244 , n22295 );
buf ( n22297 , n22296 );
buf ( n22298 , n22297 );
buf ( n22299 , n9779 );
buf ( n22300 , n22299 );
buf ( n22301 , n277450 );
buf ( n22302 , n22301 );
nor ( n22303 , n22300 , n22302 );
buf ( n22304 , n22303 );
buf ( n22305 , n22304 );
buf ( n22306 , n22299 );
buf ( n22307 , n22301 );
and ( n22308 , n22306 , n22307 );
buf ( n22309 , n22308 );
buf ( n22310 , n22309 );
nor ( n22311 , n22305 , n22310 );
buf ( n22312 , n22311 );
buf ( n22313 , n22312 );
and ( n22314 , n22298 , n22313 );
not ( n22315 , n22298 );
buf ( n22316 , n22312 );
not ( n22317 , n22316 );
buf ( n22318 , n22317 );
buf ( n22319 , n22318 );
and ( n22320 , n22315 , n22319 );
nor ( n22321 , n22314 , n22320 );
buf ( n22322 , n22321 );
buf ( n22323 , n22322 );
not ( n22324 , n22323 );
or ( n22325 , n22201 , n22324 );
nand ( n22326 , n277352 , n9779 );
nand ( n22327 , n22325 , n22326 );
not ( n22328 , n22327 );
or ( n22329 , n22328 , n14830 );
nand ( n22330 , n14830 , n13388 );
nand ( n22331 , n22329 , n22330 );
buf ( n22332 , n22331 );
buf ( n22333 , n22332 );
buf ( n22334 , n275554 );
not ( n22335 , n275557 );
and ( n22336 , n22335 , n18273 );
not ( n22337 , n22335 );
not ( n22338 , n9432 );
buf ( n22339 , n9702 );
buf ( n22340 , n22339 );
buf ( n22341 , n278001 );
buf ( n22342 , n22341 );
nor ( n22343 , n22340 , n22342 );
buf ( n22344 , n22343 );
buf ( n22345 , n22344 );
buf ( n22346 , n9710 );
buf ( n22347 , n22346 );
buf ( n22348 , n277926 );
buf ( n22349 , n22348 );
nor ( n22350 , n22347 , n22349 );
buf ( n22351 , n22350 );
buf ( n22352 , n22351 );
nor ( n22353 , n22345 , n22352 );
buf ( n22354 , n22353 );
buf ( n22355 , n22354 );
buf ( n22356 , n9728 );
buf ( n22357 , n22356 );
buf ( n22358 , n10642 );
buf ( n22359 , n22358 );
nor ( n22360 , n22357 , n22359 );
buf ( n22361 , n22360 );
buf ( n22362 , n22361 );
buf ( n22363 , n9720 );
buf ( n22364 , n22363 );
buf ( n22365 , n278049 );
buf ( n22366 , n22365 );
nor ( n22367 , n22364 , n22366 );
buf ( n22368 , n22367 );
buf ( n22369 , n22368 );
nor ( n22370 , n22362 , n22369 );
buf ( n22371 , n22370 );
buf ( n22372 , n22371 );
and ( n22373 , n22355 , n22372 );
buf ( n22374 , n22373 );
buf ( n22375 , n22374 );
buf ( n22376 , n9667 );
buf ( n22377 , n22376 );
buf ( n22378 , n22377 );
buf ( n22379 , n277891 );
buf ( n22380 , n22379 );
nor ( n22381 , n22378 , n22380 );
buf ( n22382 , n22381 );
buf ( n22383 , n22382 );
buf ( n22384 , n9675 );
buf ( n22385 , n22384 );
buf ( n22386 , n277818 );
buf ( n22387 , n22386 );
nor ( n22388 , n22385 , n22387 );
buf ( n22389 , n22388 );
buf ( n22390 , n22389 );
nor ( n22391 , n22383 , n22390 );
buf ( n22392 , n22391 );
buf ( n22393 , n22392 );
buf ( n22394 , n9692 );
buf ( n22395 , n22394 );
buf ( n22396 , n277794 );
buf ( n22397 , n22396 );
nor ( n22398 , n22395 , n22397 );
buf ( n22399 , n22398 );
buf ( n22400 , n22399 );
buf ( n22401 , n9684 );
buf ( n22402 , n22401 );
buf ( n22403 , n277745 );
buf ( n22404 , n22403 );
nor ( n22405 , n22402 , n22404 );
buf ( n22406 , n22405 );
buf ( n22407 , n22406 );
nor ( n22408 , n22400 , n22407 );
buf ( n22409 , n22408 );
buf ( n22410 , n22409 );
and ( n22411 , n22393 , n22410 );
buf ( n22412 , n22411 );
buf ( n22413 , n22412 );
and ( n22414 , n22375 , n22413 );
buf ( n22415 , n22414 );
buf ( n22416 , n22415 );
buf ( n22417 , n9740 );
buf ( n22418 , n22417 );
buf ( n22419 , n277605 );
buf ( n22420 , n22419 );
nor ( n22421 , n22418 , n22420 );
buf ( n22422 , n22421 );
buf ( n22423 , n22422 );
buf ( n22424 , n9748 );
buf ( n22425 , n22424 );
buf ( n22426 , n277529 );
buf ( n22427 , n22426 );
nor ( n22428 , n22425 , n22427 );
buf ( n22429 , n22428 );
buf ( n22430 , n22429 );
nor ( n22431 , n22423 , n22430 );
buf ( n22432 , n22431 );
buf ( n22433 , n22432 );
buf ( n22434 , n9757 );
buf ( n22435 , n22434 );
buf ( n22436 , n277646 );
buf ( n22437 , n22436 );
or ( n22438 , n22435 , n22437 );
buf ( n22439 , n22438 );
buf ( n22440 , n22439 );
buf ( n22441 , n277692 );
buf ( n22442 , n22441 );
buf ( n22443 , n9765 );
buf ( n22444 , n22443 );
or ( n22445 , n22442 , n22444 );
buf ( n22446 , n22445 );
buf ( n22447 , n22446 );
and ( n22448 , n22440 , n22447 );
buf ( n22449 , n22448 );
buf ( n22450 , n22449 );
and ( n22451 , n22433 , n22450 );
buf ( n22452 , n22451 );
buf ( n22453 , n22452 );
buf ( n22454 , n9783 );
buf ( n22455 , n22454 );
buf ( n22456 , n277408 );
buf ( n22457 , n22456 );
or ( n22458 , n22455 , n22457 );
buf ( n22459 , n22458 );
buf ( n22460 , n22459 );
not ( n22461 , n22460 );
buf ( n22462 , n9775 );
buf ( n22463 , n22462 );
buf ( n22464 , n277450 );
buf ( n22465 , n22464 );
nor ( n22466 , n22463 , n22465 );
buf ( n22467 , n22466 );
buf ( n22468 , n22467 );
nor ( n22469 , n22461 , n22468 );
buf ( n22470 , n22469 );
buf ( n22471 , n22470 );
and ( n22472 , n22453 , n22471 );
buf ( n22473 , n22472 );
buf ( n22474 , n22473 );
and ( n22475 , n22416 , n22474 );
buf ( n22476 , n22475 );
buf ( n22477 , n22476 );
not ( n22478 , n22477 );
buf ( n22479 , n19711 );
not ( n22480 , n22479 );
buf ( n22481 , n19690 );
not ( n22482 , n22481 );
or ( n22483 , n22480 , n22482 );
buf ( n22484 , n19857 );
nand ( n22485 , n22483 , n22484 );
buf ( n22486 , n22485 );
buf ( n22487 , n22486 );
buf ( n22488 , n9523 );
buf ( n22489 , n22488 );
buf ( n22490 , n11329 );
buf ( n22491 , n22490 );
or ( n22492 , n22489 , n22491 );
buf ( n22493 , n22492 );
buf ( n22494 , n22493 );
buf ( n22495 , n21282 );
nand ( n22496 , n22494 , n22495 );
buf ( n22497 , n22496 );
buf ( n22498 , n22497 );
not ( n22499 , n22498 );
buf ( n22500 , n21192 );
nand ( n22501 , n22499 , n22500 );
buf ( n22502 , n22501 );
buf ( n22503 , n22502 );
buf ( n22504 , n21215 );
nor ( n22505 , n22503 , n22504 );
buf ( n22506 , n22505 );
buf ( n22507 , n22506 );
buf ( n22508 , n19816 );
not ( n22509 , n22508 );
buf ( n22510 , n20033 );
not ( n22511 , n22510 );
or ( n22512 , n22509 , n22511 );
buf ( n22513 , n19857 );
nand ( n22514 , n22512 , n22513 );
buf ( n22515 , n22514 );
buf ( n22516 , n22515 );
nand ( n22517 , n22487 , n22507 , n22516 );
buf ( n22518 , n22517 );
buf ( n22519 , n22518 );
buf ( n22520 , n19791 );
buf ( n22521 , n20015 );
and ( n22522 , n22520 , n22521 );
buf ( n22523 , n22522 );
buf ( n22524 , n22523 );
buf ( n22525 , n19690 );
buf ( n22526 , n19711 );
and ( n22527 , n22525 , n22526 );
buf ( n22528 , n22527 );
buf ( n22529 , n22528 );
buf ( n22530 , n22502 );
not ( n22531 , n22530 );
buf ( n22532 , n22531 );
buf ( n22533 , n22532 );
buf ( n22534 , n21215 );
buf ( n22535 , n19813 );
nor ( n22536 , n22534 , n22535 );
buf ( n22537 , n22536 );
buf ( n22538 , n22537 );
nand ( n22539 , n22524 , n22529 , n22533 , n22538 );
buf ( n22540 , n22539 );
buf ( n22541 , n22540 );
buf ( n22542 , n21266 );
buf ( n22543 , n22488 );
buf ( n22544 , n22490 );
nand ( n22545 , n22543 , n22544 );
buf ( n22546 , n22545 );
buf ( n22547 , n22546 );
nand ( n22548 , n22542 , n22547 );
buf ( n22549 , n22548 );
buf ( n22550 , n22549 );
buf ( n22551 , n21287 );
nor ( n22552 , n22550 , n22551 );
buf ( n22553 , n22552 );
buf ( n22554 , n22553 );
not ( n22555 , n22554 );
buf ( n22556 , n21261 );
not ( n22557 , n22556 );
or ( n22558 , n22555 , n22557 );
buf ( n22559 , n22497 );
buf ( n22560 , n22546 );
nand ( n22561 , n22559 , n22560 );
buf ( n22562 , n22561 );
buf ( n22563 , n22562 );
nand ( n22564 , n22558 , n22563 );
buf ( n22565 , n22564 );
buf ( n22566 , n22565 );
buf ( n22567 , n21205 );
buf ( n22568 , n22493 );
buf ( n22569 , n21212 );
buf ( n22570 , n21282 );
and ( n22571 , n22567 , n22568 , n22569 , n22570 );
buf ( n22572 , n22571 );
buf ( n22573 , n22572 );
buf ( n22574 , n21241 );
nand ( n22575 , n22573 , n22574 );
buf ( n22576 , n22575 );
buf ( n22577 , n22576 );
and ( n22578 , n22566 , n22577 );
buf ( n22579 , n22578 );
buf ( n22580 , n22579 );
buf ( n22581 , n22572 );
not ( n22582 , n22581 );
buf ( n22583 , n22582 );
buf ( n22584 , n22583 );
not ( n22585 , n22584 );
buf ( n22586 , n21195 );
buf ( n22587 , n19758 );
nand ( n22588 , n22585 , n22586 , n22587 );
buf ( n22589 , n22588 );
buf ( n22590 , n22589 );
nand ( n22591 , n22519 , n22541 , n22580 , n22590 );
buf ( n22592 , n22591 );
buf ( n22593 , n22592 );
buf ( n22594 , n22593 );
not ( n22595 , n22594 );
or ( n22596 , n22478 , n22595 );
buf ( n22597 , n22412 );
not ( n22598 , n22597 );
buf ( n22599 , n22356 );
buf ( n22600 , n22358 );
and ( n22601 , n22599 , n22600 );
buf ( n22602 , n22601 );
buf ( n22603 , n22602 );
buf ( n22604 , n22368 );
not ( n22605 , n22604 );
buf ( n22606 , n22605 );
buf ( n22607 , n22606 );
nand ( n22608 , n22603 , n22607 );
buf ( n22609 , n22608 );
buf ( n22610 , n22609 );
buf ( n22611 , n22363 );
buf ( n22612 , n22365 );
nand ( n22613 , n22611 , n22612 );
buf ( n22614 , n22613 );
buf ( n22615 , n22614 );
nand ( n22616 , n22610 , n22615 );
buf ( n22617 , n22616 );
buf ( n22618 , n22617 );
not ( n22619 , n22618 );
buf ( n22620 , n22354 );
not ( n22621 , n22620 );
or ( n22622 , n22619 , n22621 );
buf ( n22623 , n22344 );
not ( n22624 , n22623 );
buf ( n22625 , n22624 );
buf ( n22626 , n22625 );
buf ( n22627 , n22346 );
buf ( n22628 , n22348 );
and ( n22629 , n22627 , n22628 );
buf ( n22630 , n22629 );
buf ( n22631 , n22630 );
and ( n22632 , n22626 , n22631 );
buf ( n22633 , n22339 );
buf ( n22634 , n22341 );
and ( n22635 , n22633 , n22634 );
buf ( n22636 , n22635 );
buf ( n22637 , n22636 );
nor ( n22638 , n22632 , n22637 );
buf ( n22639 , n22638 );
buf ( n22640 , n22639 );
nand ( n22641 , n22622 , n22640 );
buf ( n22642 , n22641 );
buf ( n22643 , n22642 );
not ( n22644 , n22643 );
or ( n22645 , n22598 , n22644 );
buf ( n22646 , n22384 );
buf ( n22647 , n22386 );
and ( n22648 , n22646 , n22647 );
buf ( n22649 , n22648 );
buf ( n22650 , n22649 );
not ( n22651 , n22650 );
buf ( n22652 , n22382 );
not ( n22653 , n22652 );
buf ( n22654 , n22653 );
buf ( n22655 , n22654 );
not ( n22656 , n22655 );
or ( n22657 , n22651 , n22656 );
buf ( n22658 , n22377 );
buf ( n22659 , n22379 );
nand ( n22660 , n22658 , n22659 );
buf ( n22661 , n22660 );
buf ( n22662 , n22661 );
nand ( n22663 , n22657 , n22662 );
buf ( n22664 , n22663 );
buf ( n22665 , n22664 );
buf ( n22666 , n22409 );
and ( n22667 , n22665 , n22666 );
buf ( n22668 , n22394 );
buf ( n22669 , n22396 );
nand ( n22670 , n22668 , n22669 );
buf ( n22671 , n22670 );
buf ( n22672 , n22671 );
buf ( n22673 , n22406 );
or ( n22674 , n22672 , n22673 );
buf ( n22675 , n22401 );
buf ( n22676 , n22403 );
nand ( n22677 , n22675 , n22676 );
buf ( n22678 , n22677 );
buf ( n22679 , n22678 );
nand ( n22680 , n22674 , n22679 );
buf ( n22681 , n22680 );
buf ( n22682 , n22681 );
nor ( n22683 , n22667 , n22682 );
buf ( n22684 , n22683 );
buf ( n22685 , n22684 );
nand ( n22686 , n22645 , n22685 );
buf ( n22687 , n22686 );
buf ( n22688 , n22687 );
buf ( n22689 , n22473 );
and ( n22690 , n22688 , n22689 );
buf ( n22691 , n22470 );
not ( n22692 , n22691 );
buf ( n22693 , n22439 );
not ( n22694 , n22693 );
buf ( n22695 , n22443 );
buf ( n22696 , n22441 );
and ( n22697 , n22695 , n22696 );
buf ( n22698 , n22697 );
buf ( n22699 , n22698 );
not ( n22700 , n22699 );
or ( n22701 , n22694 , n22700 );
buf ( n22702 , n22434 );
buf ( n22703 , n22436 );
nand ( n22704 , n22702 , n22703 );
buf ( n22705 , n22704 );
buf ( n22706 , n22705 );
nand ( n22707 , n22701 , n22706 );
buf ( n22708 , n22707 );
buf ( n22709 , n22708 );
not ( n22710 , n22709 );
buf ( n22711 , n22432 );
not ( n22712 , n22711 );
or ( n22713 , n22710 , n22712 );
buf ( n22714 , n22422 );
not ( n22715 , n22714 );
buf ( n22716 , n22424 );
buf ( n22717 , n22426 );
nand ( n22718 , n22716 , n22717 );
buf ( n22719 , n22718 );
buf ( n22720 , n22719 );
not ( n22721 , n22720 );
and ( n22722 , n22715 , n22721 );
buf ( n22723 , n22417 );
buf ( n22724 , n22419 );
and ( n22725 , n22723 , n22724 );
buf ( n22726 , n22725 );
buf ( n22727 , n22726 );
nor ( n22728 , n22722 , n22727 );
buf ( n22729 , n22728 );
buf ( n22730 , n22729 );
nand ( n22731 , n22713 , n22730 );
buf ( n22732 , n22731 );
buf ( n22733 , n22732 );
not ( n22734 , n22733 );
or ( n22735 , n22692 , n22734 );
buf ( n22736 , n22467 );
not ( n22737 , n22736 );
buf ( n22738 , n22454 );
buf ( n22739 , n22456 );
nand ( n22740 , n22738 , n22739 );
buf ( n22741 , n22740 );
buf ( n22742 , n22741 );
not ( n22743 , n22742 );
and ( n22744 , n22737 , n22743 );
buf ( n22745 , n22462 );
buf ( n22746 , n22464 );
and ( n22747 , n22745 , n22746 );
buf ( n22748 , n22747 );
buf ( n22749 , n22748 );
nor ( n22750 , n22744 , n22749 );
buf ( n22751 , n22750 );
buf ( n22752 , n22751 );
nand ( n22753 , n22735 , n22752 );
buf ( n22754 , n22753 );
buf ( n22755 , n22754 );
nor ( n22756 , n22690 , n22755 );
buf ( n22757 , n22756 );
buf ( n22758 , n22757 );
nand ( n22759 , n22596 , n22758 );
buf ( n22760 , n22759 );
buf ( n22761 , n22760 );
buf ( n22762 , n277336 );
buf ( n22763 , n22762 );
buf ( n22764 , n277353 );
buf ( n22765 , n22764 );
nor ( n22766 , n22763 , n22765 );
buf ( n22767 , n22766 );
buf ( n22768 , n22767 );
not ( n22769 , n22768 );
buf ( n22770 , n22762 );
buf ( n22771 , n22764 );
nand ( n22772 , n22770 , n22771 );
buf ( n22773 , n22772 );
buf ( n22774 , n22773 );
nand ( n22775 , n22769 , n22774 );
buf ( n22776 , n22775 );
buf ( n22777 , n22776 );
not ( n22778 , n22777 );
buf ( n22779 , n22778 );
buf ( n22780 , n22779 );
and ( n22781 , n22761 , n22780 );
not ( n22782 , n22761 );
buf ( n22783 , n22776 );
and ( n22784 , n22782 , n22783 );
nor ( n22785 , n22781 , n22784 );
buf ( n22786 , n22785 );
buf ( n22787 , n22786 );
not ( n22788 , n22787 );
or ( n22789 , n22338 , n22788 );
nand ( n22790 , n277390 , n277336 );
nand ( n22791 , n22789 , n22790 );
and ( n22792 , n22337 , n22791 );
or ( n22793 , n22336 , n22792 );
buf ( n22794 , n22793 );
buf ( n22795 , n22794 );
buf ( n22796 , n275554 );
buf ( n22797 , n275554 );
buf ( n22798 , n18208 );
buf ( n22799 , n22798 );
buf ( n22800 , n19600 );
and ( n22801 , n22799 , n22800 );
not ( n22802 , n22799 );
buf ( n22803 , n19497 );
not ( n22804 , n22803 );
buf ( n22805 , n19542 );
nand ( n22806 , n19069 , n22805 );
not ( n22807 , n22806 );
not ( n22808 , n19602 );
nand ( n22809 , n22807 , n22808 );
not ( n22810 , n22809 );
or ( n22811 , n22804 , n22810 );
or ( n22812 , n22809 , n22803 );
nand ( n22813 , n22811 , n22812 );
buf ( n22814 , n22813 );
and ( n22815 , n22802 , n22814 );
nor ( n22816 , n22801 , n22815 );
not ( n22817 , n22816 );
and ( n22818 , n22817 , n20987 );
not ( n22819 , n19358 );
not ( n22820 , n20474 );
nor ( n22821 , n22820 , n20494 );
not ( n22822 , n22821 );
buf ( n22823 , n20425 );
not ( n22824 , n20463 );
nor ( n22825 , n22824 , n20450 );
and ( n22826 , n22823 , n22825 );
not ( n22827 , n20463 );
not ( n22828 , n20486 );
or ( n22829 , n22827 , n22828 );
nand ( n22830 , n22829 , n20490 );
nor ( n22831 , n22826 , n22830 );
not ( n22832 , n22831 );
or ( n22833 , n22822 , n22832 );
or ( n22834 , n22831 , n22821 );
nand ( n22835 , n22833 , n22834 );
buf ( n22836 , n22835 );
not ( n22837 , n22836 );
or ( n22838 , n22819 , n22837 );
not ( n22839 , n20243 );
nand ( n22840 , n22839 , n20261 );
not ( n22841 , n22840 );
buf ( n22842 , n20330 );
not ( n22843 , n22842 );
buf ( n22844 , n20334 );
not ( n22845 , n20252 );
nand ( n22846 , n22844 , n22845 );
or ( n22847 , n22843 , n22846 );
not ( n22848 , n22845 );
not ( n22849 , n20200 );
or ( n22850 , n22848 , n22849 );
nand ( n22851 , n22850 , n20257 );
not ( n22852 , n22851 );
nand ( n22853 , n22847 , n22852 );
not ( n22854 , n22853 );
or ( n22855 , n22841 , n22854 );
or ( n22856 , n22853 , n22840 );
nand ( n22857 , n22855 , n22856 );
buf ( n22858 , n22857 );
and ( n22859 , n22858 , n21001 );
not ( n22860 , n20525 );
not ( n22861 , n20537 );
nand ( n22862 , n22860 , n20546 , n22861 );
xor ( n22863 , n22862 , n20528 );
buf ( n22864 , n22863 );
not ( n22865 , n22864 );
or ( n22866 , n22865 , n19289 );
not ( n22867 , n19219 );
not ( n22868 , n20526 );
buf ( n22869 , n22868 );
buf ( n22870 , n22869 );
buf ( n22871 , n22870 );
not ( n22872 , n22871 );
or ( n22873 , n22867 , n22872 );
nand ( n22874 , n22866 , n22873 );
nor ( n22875 , n22859 , n22874 );
nand ( n22876 , n22838 , n22875 );
nor ( n22877 , n22818 , n22876 );
or ( n22878 , n22877 , n21030 );
nand ( n22879 , n21030 , n18882 );
nand ( n22880 , n22878 , n22879 );
buf ( n22881 , n22880 );
buf ( n22882 , n22881 );
not ( n22883 , n275925 );
buf ( n22884 , n22883 );
buf ( n22885 , n22884 );
buf ( n22886 , n275554 );
buf ( n22887 , n275554 );
not ( n22888 , n275929 );
buf ( n22889 , n22888 );
buf ( n22890 , n22889 );
not ( n22891 , n275929 );
buf ( n22892 , n22891 );
buf ( n22893 , n22892 );
not ( n22894 , n14896 );
not ( n22895 , n14840 );
or ( n22896 , n22894 , n22895 );
not ( n22897 , n14831 );
nand ( n22898 , n14838 , n14830 );
nand ( n22899 , n22897 , n22898 );
not ( n22900 , n13372 );
not ( n22901 , n14915 );
nor ( n22902 , n22900 , n22901 );
nand ( n22903 , n22899 , n22902 );
nand ( n22904 , n22896 , n22903 );
and ( n22905 , n22904 , n275878 );
nor ( n22906 , n14830 , n17515 );
nor ( n22907 , n22905 , n22906 );
not ( n22908 , n14895 );
not ( n22909 , n14831 );
or ( n22910 , n22908 , n22909 );
nand ( n22911 , n22910 , n22898 );
not ( n22912 , n22901 );
nor ( n22913 , n13373 , n22912 );
and ( n22914 , n22911 , n22913 );
buf ( n22915 , n13172 );
nand ( n22916 , n22914 , n22915 );
nor ( n22917 , n20672 , n22901 );
and ( n22918 , n22911 , n22917 );
buf ( n22919 , n22915 );
buf ( n22920 , n22919 );
buf ( n22921 , n13724 );
buf ( n22922 , n22921 );
nor ( n22923 , n22920 , n22922 );
buf ( n22924 , n22923 );
buf ( n22925 , n22924 );
not ( n22926 , n22925 );
buf ( n22927 , n22919 );
buf ( n22928 , n22921 );
nand ( n22929 , n22927 , n22928 );
buf ( n22930 , n22929 );
buf ( n22931 , n22930 );
nand ( n22932 , n22926 , n22931 );
buf ( n22933 , n22932 );
buf ( n22934 , n22933 );
not ( n22935 , n22934 );
buf ( n22936 , n12936 );
buf ( n22937 , n22936 );
buf ( n22938 , n22937 );
buf ( n22939 , n13568 );
buf ( n22940 , n22939 );
nor ( n22941 , n22938 , n22940 );
buf ( n22942 , n22941 );
buf ( n22943 , n22942 );
buf ( n22944 , n13019 );
buf ( n22945 , n22944 );
buf ( n22946 , n22945 );
buf ( n22947 , n13589 );
buf ( n22948 , n22947 );
nand ( n22949 , n22946 , n22948 );
buf ( n22950 , n22949 );
buf ( n22951 , n22950 );
or ( n22952 , n22943 , n22951 );
buf ( n22953 , n22937 );
buf ( n22954 , n22939 );
nand ( n22955 , n22953 , n22954 );
buf ( n22956 , n22955 );
buf ( n22957 , n22956 );
nand ( n22958 , n22952 , n22957 );
buf ( n22959 , n22958 );
buf ( n22960 , n22959 );
buf ( n22961 , n13033 );
buf ( n22962 , n22961 );
buf ( n22963 , n22962 );
buf ( n22964 , n13674 );
buf ( n22965 , n22964 );
nor ( n22966 , n22963 , n22965 );
buf ( n22967 , n22966 );
buf ( n22968 , n22967 );
buf ( n22969 , n13049 );
buf ( n22970 , n22969 );
buf ( n22971 , n22970 );
buf ( n22972 , n13649 );
buf ( n22973 , n22972 );
nand ( n22974 , n22971 , n22973 );
buf ( n22975 , n22974 );
buf ( n22976 , n22975 );
or ( n22977 , n22968 , n22976 );
buf ( n22978 , n22962 );
buf ( n22979 , n22964 );
nand ( n22980 , n22978 , n22979 );
buf ( n22981 , n22980 );
buf ( n22982 , n22981 );
nand ( n22983 , n22977 , n22982 );
buf ( n22984 , n22983 );
buf ( n22985 , n22984 );
nor ( n22986 , n22960 , n22985 );
buf ( n22987 , n22986 );
buf ( n22988 , n22987 );
buf ( n22989 , n22967 );
buf ( n22990 , n22970 );
buf ( n22991 , n22972 );
nor ( n22992 , n22990 , n22991 );
buf ( n22993 , n22992 );
buf ( n22994 , n22993 );
nor ( n22995 , n22989 , n22994 );
buf ( n22996 , n22995 );
buf ( n22997 , n22996 );
buf ( n22998 , n13067 );
buf ( n22999 , n22998 );
buf ( n23000 , n22999 );
buf ( n23001 , n13549 );
buf ( n23002 , n23001 );
nor ( n23003 , n23000 , n23002 );
buf ( n23004 , n23003 );
buf ( n23005 , n23004 );
buf ( n23006 , n14770 );
buf ( n23007 , n13101 );
and ( n23008 , n23006 , n23007 );
buf ( n23009 , n23008 );
buf ( n23010 , n23009 );
buf ( n23011 , n14535 );
xor ( n23012 , n23010 , n23011 );
buf ( n23013 , n13099 );
and ( n23014 , n23012 , n23013 );
and ( n23015 , n23010 , n23011 );
or ( n23016 , n23014 , n23015 );
buf ( n23017 , n23016 );
buf ( n23018 , n23017 );
buf ( n23019 , n13084 );
buf ( n23020 , n23019 );
buf ( n23021 , n14554 );
buf ( n23022 , n23021 );
or ( n23023 , n23020 , n23022 );
buf ( n23024 , n23023 );
buf ( n23025 , n23024 );
nand ( n23026 , n23018 , n23025 );
buf ( n23027 , n23026 );
buf ( n23028 , n23027 );
or ( n23029 , n23005 , n23028 );
buf ( n23030 , n23004 );
buf ( n23031 , n23019 );
buf ( n23032 , n23021 );
nand ( n23033 , n23031 , n23032 );
buf ( n23034 , n23033 );
buf ( n23035 , n23034 );
or ( n23036 , n23030 , n23035 );
buf ( n23037 , n22999 );
buf ( n23038 , n23001 );
nand ( n23039 , n23037 , n23038 );
buf ( n23040 , n23039 );
buf ( n23041 , n23040 );
nand ( n23042 , n23029 , n23036 , n23041 );
buf ( n23043 , n23042 );
buf ( n23044 , n23043 );
nand ( n23045 , n22997 , n23044 );
buf ( n23046 , n23045 );
buf ( n23047 , n23046 );
and ( n23048 , n22988 , n23047 );
buf ( n23049 , n22959 );
buf ( n23050 , n22942 );
buf ( n23051 , n22945 );
buf ( n23052 , n22947 );
nor ( n23053 , n23051 , n23052 );
buf ( n23054 , n23053 );
buf ( n23055 , n23054 );
nor ( n23056 , n23050 , n23055 );
buf ( n23057 , n23056 );
buf ( n23058 , n23057 );
or ( n23059 , n23049 , n23058 );
buf ( n23060 , n13120 );
buf ( n23061 , n23060 );
buf ( n23062 , n23061 );
buf ( n23063 , n13474 );
buf ( n23064 , n23063 );
or ( n23065 , n23062 , n23064 );
buf ( n23066 , n23065 );
buf ( n23067 , n23066 );
not ( n23068 , n23067 );
buf ( n23069 , n13003 );
buf ( n23070 , n23069 );
buf ( n23071 , n23070 );
buf ( n23072 , n13452 );
buf ( n23073 , n23072 );
nor ( n23074 , n23071 , n23073 );
buf ( n23075 , n23074 );
buf ( n23076 , n23075 );
nor ( n23077 , n23068 , n23076 );
buf ( n23078 , n23077 );
buf ( n23079 , n23078 );
buf ( n23080 , n13140 );
buf ( n23081 , n23080 );
buf ( n23082 , n23081 );
buf ( n23083 , n13614 );
buf ( n23084 , n23083 );
nor ( n23085 , n23082 , n23084 );
buf ( n23086 , n23085 );
buf ( n23087 , n23086 );
buf ( n23088 , n13154 );
buf ( n23089 , n23088 );
buf ( n23090 , n23089 );
buf ( n23091 , n13629 );
buf ( n23092 , n23091 );
nor ( n23093 , n23090 , n23092 );
buf ( n23094 , n23093 );
buf ( n23095 , n23094 );
nor ( n23096 , n23087 , n23095 );
buf ( n23097 , n23096 );
buf ( n23098 , n23097 );
nand ( n23099 , n23059 , n23079 , n23098 );
buf ( n23100 , n23099 );
buf ( n23101 , n23100 );
nor ( n23102 , n23048 , n23101 );
buf ( n23103 , n23102 );
buf ( n23104 , n23103 );
buf ( n23105 , n23075 );
buf ( n23106 , n23061 );
buf ( n23107 , n23063 );
nand ( n23108 , n23106 , n23107 );
buf ( n23109 , n23108 );
buf ( n23110 , n23109 );
or ( n23111 , n23105 , n23110 );
buf ( n23112 , n23078 );
buf ( n23113 , n23086 );
buf ( n23114 , n23089 );
buf ( n23115 , n23091 );
nand ( n23116 , n23114 , n23115 );
buf ( n23117 , n23116 );
buf ( n23118 , n23117 );
or ( n23119 , n23113 , n23118 );
buf ( n23120 , n23081 );
buf ( n23121 , n23083 );
nand ( n23122 , n23120 , n23121 );
buf ( n23123 , n23122 );
buf ( n23124 , n23123 );
nand ( n23125 , n23119 , n23124 );
buf ( n23126 , n23125 );
buf ( n23127 , n23126 );
nand ( n23128 , n23112 , n23127 );
buf ( n23129 , n23128 );
buf ( n23130 , n23129 );
buf ( n23131 , n23070 );
buf ( n23132 , n23072 );
nand ( n23133 , n23131 , n23132 );
buf ( n23134 , n23133 );
buf ( n23135 , n23134 );
nand ( n23136 , n23111 , n23130 , n23135 );
buf ( n23137 , n23136 );
buf ( n23138 , n23137 );
or ( n23139 , n23104 , n23138 );
buf ( n23140 , n23139 );
buf ( n23141 , n23140 );
not ( n23142 , n23141 );
or ( n23143 , n22935 , n23142 );
buf ( n23144 , n23140 );
buf ( n23145 , n22933 );
or ( n23146 , n23144 , n23145 );
nand ( n23147 , n23143 , n23146 );
buf ( n23148 , n23147 );
buf ( n23149 , n23148 );
nand ( n23150 , n22918 , n23149 );
and ( n23151 , n22900 , n22901 );
and ( n23152 , n22911 , n23151 );
buf ( n23153 , n22915 );
buf ( n23154 , n23153 );
buf ( n23155 , n13718 );
buf ( n23156 , n23155 );
nor ( n23157 , n23154 , n23156 );
buf ( n23158 , n23157 );
buf ( n23159 , n23158 );
not ( n23160 , n23159 );
buf ( n23161 , n23153 );
buf ( n23162 , n23155 );
nand ( n23163 , n23161 , n23162 );
buf ( n23164 , n23163 );
buf ( n23165 , n23164 );
nand ( n23166 , n23160 , n23165 );
buf ( n23167 , n23166 );
buf ( n23168 , n23167 );
not ( n23169 , n23168 );
buf ( n23170 , n22936 );
buf ( n23171 , n23170 );
buf ( n23172 , n13571 );
buf ( n23173 , n23172 );
nor ( n23174 , n23171 , n23173 );
buf ( n23175 , n23174 );
buf ( n23176 , n23175 );
buf ( n23177 , n22944 );
buf ( n23178 , n23177 );
buf ( n23179 , n13585 );
buf ( n23180 , n23179 );
nand ( n23181 , n23178 , n23180 );
buf ( n23182 , n23181 );
buf ( n23183 , n23182 );
or ( n23184 , n23176 , n23183 );
buf ( n23185 , n23170 );
buf ( n23186 , n23172 );
nand ( n23187 , n23185 , n23186 );
buf ( n23188 , n23187 );
buf ( n23189 , n23188 );
nand ( n23190 , n23184 , n23189 );
buf ( n23191 , n23190 );
buf ( n23192 , n23191 );
buf ( n23193 , n22961 );
buf ( n23194 , n23193 );
buf ( n23195 , n13670 );
buf ( n23196 , n23195 );
nor ( n23197 , n23194 , n23196 );
buf ( n23198 , n23197 );
buf ( n23199 , n23198 );
buf ( n23200 , n22969 );
buf ( n23201 , n23200 );
buf ( n23202 , n13645 );
buf ( n23203 , n23202 );
nand ( n23204 , n23201 , n23203 );
buf ( n23205 , n23204 );
buf ( n23206 , n23205 );
or ( n23207 , n23199 , n23206 );
buf ( n23208 , n23193 );
buf ( n23209 , n23195 );
nand ( n23210 , n23208 , n23209 );
buf ( n23211 , n23210 );
buf ( n23212 , n23211 );
nand ( n23213 , n23207 , n23212 );
buf ( n23214 , n23213 );
buf ( n23215 , n23214 );
nor ( n23216 , n23192 , n23215 );
buf ( n23217 , n23216 );
buf ( n23218 , n23217 );
buf ( n23219 , n23198 );
buf ( n23220 , n23200 );
buf ( n23221 , n23202 );
nor ( n23222 , n23220 , n23221 );
buf ( n23223 , n23222 );
buf ( n23224 , n23223 );
nor ( n23225 , n23219 , n23224 );
buf ( n23226 , n23225 );
buf ( n23227 , n23226 );
buf ( n23228 , n22998 );
buf ( n23229 , n23228 );
buf ( n23230 , n13546 );
buf ( n23231 , n23230 );
nor ( n23232 , n23229 , n23231 );
buf ( n23233 , n23232 );
buf ( n23234 , n23233 );
buf ( n23235 , n14773 );
buf ( n23236 , n13101 );
and ( n23237 , n23235 , n23236 );
buf ( n23238 , n23237 );
buf ( n23239 , n23238 );
buf ( n23240 , n14539 );
xor ( n23241 , n23239 , n23240 );
buf ( n23242 , n13099 );
and ( n23243 , n23241 , n23242 );
and ( n23244 , n23239 , n23240 );
or ( n23245 , n23243 , n23244 );
buf ( n23246 , n23245 );
buf ( n23247 , n23246 );
buf ( n23248 , n13084 );
buf ( n23249 , n23248 );
buf ( n23250 , n14550 );
buf ( n23251 , n23250 );
or ( n23252 , n23249 , n23251 );
buf ( n23253 , n23252 );
buf ( n23254 , n23253 );
nand ( n23255 , n23247 , n23254 );
buf ( n23256 , n23255 );
buf ( n23257 , n23256 );
or ( n23258 , n23234 , n23257 );
buf ( n23259 , n23233 );
buf ( n23260 , n23248 );
buf ( n23261 , n23250 );
nand ( n23262 , n23260 , n23261 );
buf ( n23263 , n23262 );
buf ( n23264 , n23263 );
or ( n23265 , n23259 , n23264 );
buf ( n23266 , n23228 );
buf ( n23267 , n23230 );
nand ( n23268 , n23266 , n23267 );
buf ( n23269 , n23268 );
buf ( n23270 , n23269 );
nand ( n23271 , n23258 , n23265 , n23270 );
buf ( n23272 , n23271 );
buf ( n23273 , n23272 );
nand ( n23274 , n23227 , n23273 );
buf ( n23275 , n23274 );
buf ( n23276 , n23275 );
and ( n23277 , n23218 , n23276 );
buf ( n23278 , n23191 );
buf ( n23279 , n23175 );
buf ( n23280 , n23177 );
buf ( n23281 , n23179 );
nor ( n23282 , n23280 , n23281 );
buf ( n23283 , n23282 );
buf ( n23284 , n23283 );
nor ( n23285 , n23279 , n23284 );
buf ( n23286 , n23285 );
buf ( n23287 , n23286 );
or ( n23288 , n23278 , n23287 );
buf ( n23289 , n23060 );
buf ( n23290 , n23289 );
buf ( n23291 , n13471 );
buf ( n23292 , n23291 );
or ( n23293 , n23290 , n23292 );
buf ( n23294 , n23293 );
buf ( n23295 , n23294 );
not ( n23296 , n23295 );
buf ( n23297 , n23069 );
buf ( n23298 , n23297 );
buf ( n23299 , n13446 );
buf ( n23300 , n23299 );
nor ( n23301 , n23298 , n23300 );
buf ( n23302 , n23301 );
buf ( n23303 , n23302 );
nor ( n23304 , n23296 , n23303 );
buf ( n23305 , n23304 );
buf ( n23306 , n23305 );
buf ( n23307 , n23080 );
buf ( n23308 , n23307 );
buf ( n23309 , n13611 );
buf ( n23310 , n23309 );
nor ( n23311 , n23308 , n23310 );
buf ( n23312 , n23311 );
buf ( n23313 , n23312 );
buf ( n23314 , n23088 );
buf ( n23315 , n23314 );
buf ( n23316 , n13626 );
buf ( n23317 , n23316 );
nor ( n23318 , n23315 , n23317 );
buf ( n23319 , n23318 );
buf ( n23320 , n23319 );
nor ( n23321 , n23313 , n23320 );
buf ( n23322 , n23321 );
buf ( n23323 , n23322 );
nand ( n23324 , n23288 , n23306 , n23323 );
buf ( n23325 , n23324 );
buf ( n23326 , n23325 );
nor ( n23327 , n23277 , n23326 );
buf ( n23328 , n23327 );
buf ( n23329 , n23328 );
buf ( n23330 , n23302 );
buf ( n23331 , n23289 );
buf ( n23332 , n23291 );
nand ( n23333 , n23331 , n23332 );
buf ( n23334 , n23333 );
buf ( n23335 , n23334 );
or ( n23336 , n23330 , n23335 );
buf ( n23337 , n23305 );
buf ( n23338 , n23312 );
buf ( n23339 , n23314 );
buf ( n23340 , n23316 );
nand ( n23341 , n23339 , n23340 );
buf ( n23342 , n23341 );
buf ( n23343 , n23342 );
or ( n23344 , n23338 , n23343 );
buf ( n23345 , n23307 );
buf ( n23346 , n23309 );
nand ( n23347 , n23345 , n23346 );
buf ( n23348 , n23347 );
buf ( n23349 , n23348 );
nand ( n23350 , n23344 , n23349 );
buf ( n23351 , n23350 );
buf ( n23352 , n23351 );
nand ( n23353 , n23337 , n23352 );
buf ( n23354 , n23353 );
buf ( n23355 , n23354 );
buf ( n23356 , n23297 );
buf ( n23357 , n23299 );
nand ( n23358 , n23356 , n23357 );
buf ( n23359 , n23358 );
buf ( n23360 , n23359 );
nand ( n23361 , n23336 , n23355 , n23360 );
buf ( n23362 , n23361 );
buf ( n23363 , n23362 );
or ( n23364 , n23329 , n23363 );
buf ( n23365 , n23364 );
buf ( n23366 , n23365 );
not ( n23367 , n23366 );
or ( n23368 , n23169 , n23367 );
buf ( n23369 , n23365 );
buf ( n23370 , n23167 );
or ( n23371 , n23369 , n23370 );
nand ( n23372 , n23368 , n23371 );
buf ( n23373 , n23372 );
buf ( n23374 , n23373 );
nand ( n23375 , n23152 , n23374 );
nand ( n23376 , n22907 , n22916 , n23150 , n23375 );
buf ( n23377 , n23376 );
buf ( n23378 , n23377 );
not ( n23379 , n277928 );
or ( n23380 , n23379 , n9158 );
not ( n23381 , n277906 );
or ( n23382 , n23381 , n9157 );
nand ( n23383 , n23380 , n23382 );
buf ( n23384 , n23383 );
buf ( n23385 , n23384 );
not ( n23386 , n13373 );
not ( n23387 , n23386 );
buf ( n23388 , n14426 );
not ( n23389 , n23388 );
and ( n23390 , n14777 , n20717 , n20728 );
nand ( n23391 , n23390 , n20724 );
buf ( n23392 , n23391 );
not ( n23393 , n23392 );
or ( n23394 , n23389 , n23393 );
or ( n23395 , n23392 , n23388 );
nand ( n23396 , n23394 , n23395 );
buf ( n23397 , n23396 );
not ( n23398 , n23397 );
or ( n23399 , n23387 , n23398 );
not ( n23400 , n23386 );
buf ( n23401 , n14227 );
nand ( n23402 , n23400 , n23401 );
nand ( n23403 , n23399 , n23402 );
not ( n23404 , n20846 );
and ( n23405 , n23403 , n23404 );
not ( n23406 , n20889 );
nand ( n23407 , n15831 , n16920 );
not ( n23408 , n23407 );
not ( n23409 , n15907 );
not ( n23410 , n16913 );
or ( n23411 , n23409 , n23410 );
buf ( n23412 , n16918 );
nand ( n23413 , n23411 , n23412 );
not ( n23414 , n23413 );
or ( n23415 , n23408 , n23414 );
or ( n23416 , n23413 , n23407 );
nand ( n23417 , n23415 , n23416 );
buf ( n23418 , n23417 );
not ( n23419 , n23418 );
or ( n23420 , n23406 , n23419 );
not ( n23421 , n16996 );
nand ( n23422 , n23421 , n17377 );
not ( n23423 , n23422 );
not ( n23424 , n17007 );
not ( n23425 , n23424 );
not ( n23426 , n17362 );
or ( n23427 , n23425 , n23426 );
nand ( n23428 , n23427 , n17378 );
not ( n23429 , n23428 );
or ( n23430 , n23423 , n23429 );
or ( n23431 , n23428 , n23422 );
nand ( n23432 , n23430 , n23431 );
buf ( n23433 , n23432 );
and ( n23434 , n23433 , n20927 );
not ( n23435 , n17409 );
buf ( n23436 , n17462 );
nand ( n23437 , n23436 , n17471 );
and ( n23438 , n23437 , n17481 );
not ( n23439 , n23437 );
and ( n23440 , n23439 , n17482 );
nor ( n23441 , n23438 , n23440 );
buf ( n23442 , n23441 );
not ( n23443 , n23442 );
or ( n23444 , n23435 , n23443 );
buf ( n23445 , n17480 );
buf ( n23446 , n23445 );
buf ( n23447 , n23446 );
nand ( n23448 , n20940 , n23447 );
nand ( n23449 , n23444 , n23448 );
nor ( n23450 , n23434 , n23449 );
nand ( n23451 , n23420 , n23450 );
nor ( n23452 , n23405 , n23451 );
or ( n23453 , n23452 , n20951 );
nand ( n23454 , n20953 , n13762 );
nand ( n23455 , n23453 , n23454 );
buf ( n23456 , n23455 );
buf ( n23457 , n23456 );
buf ( n23458 , n275554 );
and ( n23459 , n9158 , n9068 );
not ( n23460 , n9158 );
and ( n23461 , n23460 , n277694 );
or ( n23462 , n23459 , n23461 );
buf ( n23463 , n23462 );
buf ( n23464 , n23463 );
buf ( n23465 , n11543 );
buf ( n23466 , n23465 );
not ( n23467 , n23466 );
buf ( n23468 , n23467 );
buf ( n23469 , n23468 );
buf ( n23470 , n11573 );
buf ( n23471 , n23470 );
not ( n23472 , n23471 );
buf ( n23473 , n23472 );
buf ( n23474 , n23473 );
nand ( n23475 , n23469 , n23474 );
buf ( n23476 , n23475 );
buf ( n23477 , n23476 );
buf ( n23478 , n23465 );
buf ( n23479 , n23470 );
nand ( n23480 , n23478 , n23479 );
buf ( n23481 , n23480 );
buf ( n23482 , n23481 );
nand ( n23483 , n23477 , n23482 );
buf ( n23484 , n23483 );
buf ( n23485 , n23484 );
not ( n23486 , n23485 );
buf ( n23487 , n11619 );
buf ( n23488 , n23487 );
not ( n23489 , n23488 );
buf ( n23490 , n23489 );
buf ( n23491 , n23490 );
buf ( n23492 , n11596 );
buf ( n23493 , n23492 );
not ( n23494 , n23493 );
buf ( n23495 , n23494 );
buf ( n23496 , n23495 );
nand ( n23497 , n23491 , n23496 );
buf ( n23498 , n23497 );
buf ( n23499 , n23498 );
buf ( n23500 , n11649 );
buf ( n23501 , n23500 );
not ( n23502 , n23501 );
buf ( n23503 , n23502 );
buf ( n23504 , n23503 );
buf ( n23505 , n11677 );
buf ( n23506 , n23505 );
not ( n23507 , n23506 );
buf ( n23508 , n23507 );
buf ( n23509 , n23508 );
nand ( n23510 , n23504 , n23509 );
buf ( n23511 , n23510 );
buf ( n23512 , n23511 );
nand ( n23513 , n23499 , n23512 );
buf ( n23514 , n23513 );
buf ( n23515 , n23514 );
buf ( n23516 , n23515 );
not ( n23517 , n23516 );
buf ( n23518 , n23517 );
buf ( n23519 , n23518 );
not ( n23520 , n23519 );
buf ( n23521 , n21898 );
buf ( n23522 , n21906 );
buf ( n23523 , n21928 );
nand ( n23524 , n23522 , n23523 );
buf ( n23525 , n23524 );
buf ( n23526 , n23525 );
buf ( n23527 , n21921 );
nand ( n23528 , n23521 , n23526 , n23527 );
buf ( n23529 , n23528 );
buf ( n23530 , n23529 );
buf ( n23531 , n21885 );
not ( n23532 , n23531 );
buf ( n23533 , n23532 );
buf ( n23534 , n23533 );
nand ( n23535 , n23530 , n23534 );
buf ( n23536 , n23535 );
buf ( n23537 , n23536 );
buf ( n23538 , n21945 );
buf ( n23539 , n21826 );
buf ( n23540 , n21869 );
and ( n23541 , n23538 , n23539 , n23540 );
buf ( n23542 , n23541 );
buf ( n23543 , n23542 );
buf ( n23544 , n21799 );
buf ( n23545 , n21969 );
and ( n23546 , n23544 , n23545 );
buf ( n23547 , n23546 );
buf ( n23548 , n23547 );
nand ( n23549 , n23537 , n23543 , n23548 );
buf ( n23550 , n23549 );
buf ( n23551 , n23550 );
buf ( n23552 , n23547 );
buf ( n23553 , n21842 );
and ( n23554 , n23552 , n23553 );
buf ( n23555 , n21849 );
not ( n23556 , n23555 );
buf ( n23557 , n21969 );
not ( n23558 , n23557 );
or ( n23559 , n23556 , n23558 );
buf ( n23560 , n21976 );
nand ( n23561 , n23559 , n23560 );
buf ( n23562 , n23561 );
buf ( n23563 , n23562 );
nor ( n23564 , n23554 , n23563 );
buf ( n23565 , n23564 );
buf ( n23566 , n23565 );
nand ( n23567 , n23551 , n23566 );
buf ( n23568 , n23567 );
buf ( n23569 , n23568 );
not ( n23570 , n23569 );
or ( n23571 , n23520 , n23570 );
buf ( n23572 , n23487 );
buf ( n23573 , n23492 );
and ( n23574 , n23572 , n23573 );
buf ( n23575 , n23574 );
buf ( n23576 , n23575 );
buf ( n23577 , n23511 );
nand ( n23578 , n23576 , n23577 );
buf ( n23579 , n23578 );
buf ( n23580 , n23579 );
buf ( n23581 , n23500 );
buf ( n23582 , n23505 );
nand ( n23583 , n23581 , n23582 );
buf ( n23584 , n23583 );
buf ( n23585 , n23584 );
nand ( n23586 , n23580 , n23585 );
buf ( n23587 , n23586 );
buf ( n23588 , n23587 );
not ( n23589 , n23588 );
buf ( n23590 , n23589 );
buf ( n23591 , n23590 );
nand ( n23592 , n23571 , n23591 );
buf ( n23593 , n23592 );
buf ( n23594 , n23593 );
not ( n23595 , n23594 );
or ( n23596 , n23486 , n23595 );
buf ( n23597 , n23593 );
buf ( n23598 , n23484 );
or ( n23599 , n23597 , n23598 );
nand ( n23600 , n23596 , n23599 );
buf ( n23601 , n23600 );
buf ( n23602 , n23601 );
not ( n23603 , n22001 );
nand ( n23604 , n23602 , n23603 );
buf ( n23605 , n11543 );
not ( n23606 , n23605 );
buf ( n23607 , n11573 );
nand ( n23608 , n23606 , n23607 );
not ( n23609 , n23607 );
nand ( n23610 , n23609 , n23605 );
nand ( n23611 , n23608 , n23610 );
not ( n23612 , n23611 );
buf ( n23613 , n11619 );
not ( n23614 , n23613 );
buf ( n23615 , n11596 );
nand ( n23616 , n23614 , n23615 );
buf ( n23617 , n11649 );
not ( n23618 , n23617 );
buf ( n23619 , n11676 );
nand ( n23620 , n23618 , n23619 );
nand ( n23621 , n23616 , n23620 );
not ( n23622 , n23621 );
not ( n23623 , n23622 );
nand ( n23624 , n22073 , n22062 );
not ( n23625 , n23624 );
not ( n23626 , n23625 );
not ( n23627 , n22089 );
or ( n23628 , n23626 , n23627 );
not ( n23629 , n22062 );
not ( n23630 , n22093 );
or ( n23631 , n23629 , n23630 );
nand ( n23632 , n23631 , n22067 );
not ( n23633 , n23632 );
nand ( n23634 , n23628 , n23633 );
not ( n23635 , n23634 );
nor ( n23636 , n22132 , n23624 );
nand ( n23637 , n22129 , n23636 );
nand ( n23638 , n23635 , n23637 );
not ( n23639 , n23638 );
or ( n23640 , n23623 , n23639 );
not ( n23641 , n23615 );
and ( n23642 , n23613 , n23641 );
nand ( n23643 , n23642 , n23620 );
not ( n23644 , n23619 );
nand ( n23645 , n23644 , n23617 );
buf ( n23646 , n23645 );
nand ( n23647 , n23643 , n23646 );
not ( n23648 , n23647 );
nand ( n23649 , n23640 , n23648 );
not ( n23650 , n23649 );
or ( n23651 , n23612 , n23650 );
or ( n23652 , n23649 , n23611 );
nand ( n23653 , n23651 , n23652 );
buf ( n23654 , n23653 );
buf ( n23655 , n22057 );
nand ( n23656 , n23654 , n23655 );
buf ( n23657 , n11483 );
buf ( n23658 , n23657 );
not ( n23659 , n23658 );
buf ( n23660 , n11649 );
nand ( n23661 , n22039 , n22043 , n23660 );
nor ( n23662 , n22037 , n23661 );
buf ( n23663 , n11543 );
and ( n23664 , n22033 , n23663 );
nand ( n23665 , n22024 , n23662 , n23664 );
buf ( n23666 , n23665 );
not ( n23667 , n23666 );
or ( n23668 , n23659 , n23667 );
or ( n23669 , n23666 , n23658 );
nand ( n23670 , n23668 , n23669 );
buf ( n23671 , n23670 );
not ( n23672 , n22051 );
buf ( n23673 , n23672 );
and ( n23674 , n23671 , n23673 );
buf ( n23675 , n22006 );
buf ( n23676 , n11649 );
not ( n23677 , n23676 );
or ( n23678 , n23675 , n23677 );
not ( n23679 , n22012 );
not ( n23680 , n23679 );
or ( n23681 , n23680 , n12258 );
nand ( n23682 , n23678 , n23681 );
nor ( n23683 , n23674 , n23682 );
and ( n23684 , n23604 , n23656 , n23683 );
not ( n23685 , n22187 );
buf ( n23686 , n22169 );
nor ( n23687 , n23685 , n23686 );
not ( n23688 , n23687 );
nand ( n23689 , n22177 , n22181 , n22182 );
not ( n23690 , n12378 );
nor ( n23691 , n23689 , n23690 );
not ( n23692 , n23691 );
not ( n23693 , n23692 );
or ( n23694 , n23688 , n23693 );
nand ( n23695 , n22146 , n22162 , n23686 );
buf ( n23696 , n23695 );
not ( n23697 , n23696 );
not ( n23698 , n12108 );
not ( n23699 , n12377 );
or ( n23700 , n23698 , n23699 );
nand ( n23701 , n23700 , n9153 );
nand ( n23702 , n23697 , n23701 );
nand ( n23703 , n23694 , n23702 );
buf ( n23704 , n23703 );
not ( n23705 , n23704 );
buf ( n23706 , n23705 );
or ( n23707 , n23684 , n23706 );
not ( n23708 , n23704 );
nand ( n23709 , n23708 , n11538 );
nand ( n23710 , n23707 , n23709 );
buf ( n23711 , n23710 );
buf ( n23712 , n23711 );
buf ( n23713 , n275554 );
buf ( n23714 , n275554 );
buf ( n23715 , n275554 );
not ( n23716 , n20889 );
buf ( n23717 , n15731 );
nor ( n23718 , n23717 , n16935 );
not ( n23719 , n23718 );
buf ( n23720 , n16923 );
nand ( n23721 , n16878 , n16911 , n23720 );
not ( n23722 , n15908 );
nand ( n23723 , n23720 , n23722 );
nand ( n23724 , n23721 , n23723 );
not ( n23725 , n23724 );
or ( n23726 , n23719 , n23725 );
or ( n23727 , n23724 , n23718 );
nand ( n23728 , n23726 , n23727 );
buf ( n23729 , n23728 );
not ( n23730 , n23729 );
or ( n23731 , n23716 , n23730 );
buf ( n23732 , n17020 );
not ( n23733 , n23732 );
buf ( n23734 , n17383 );
nand ( n23735 , n23733 , n23734 );
not ( n23736 , n23735 );
and ( n23737 , n17342 , n17353 );
not ( n23738 , n17283 );
nand ( n23739 , n23738 , n17358 );
nor ( n23740 , n23739 , n17328 );
nand ( n23741 , n23737 , n23740 );
not ( n23742 , n17229 );
nor ( n23743 , n23742 , n17357 );
nand ( n23744 , n23737 , n23743 );
not ( n23745 , n17315 );
nand ( n23746 , n23745 , n17358 );
nor ( n23747 , n23746 , n17328 );
nand ( n23748 , n23737 , n23747 );
nand ( n23749 , n17342 , n17353 , n17181 , n17358 );
nand ( n23750 , n17353 , n17144 , n17358 );
and ( n23751 , n23749 , n23750 , n17008 );
nand ( n23752 , n23741 , n23744 , n23748 , n23751 );
not ( n23753 , n17380 );
nand ( n23754 , n23752 , n23753 );
not ( n23755 , n23754 );
or ( n23756 , n23736 , n23755 );
or ( n23757 , n23754 , n23735 );
nand ( n23758 , n23756 , n23757 );
buf ( n23759 , n23758 );
and ( n23760 , n23759 , n20927 );
not ( n23761 , n17409 );
nand ( n23762 , n17462 , n20774 );
xnor ( n23763 , n23762 , n17489 );
buf ( n23764 , n23763 );
not ( n23765 , n23764 );
or ( n23766 , n23761 , n23765 );
buf ( n23767 , n17487 );
buf ( n23768 , n23767 );
buf ( n23769 , n23768 );
nand ( n23770 , n20940 , n23769 );
nand ( n23771 , n23766 , n23770 );
nor ( n23772 , n23760 , n23771 );
nand ( n23773 , n23731 , n23772 );
buf ( n23774 , n14079 );
and ( n23775 , n13373 , n23774 );
not ( n23776 , n13373 );
not ( n23777 , n23388 );
nor ( n23778 , n23391 , n23777 );
not ( n23779 , n23778 );
not ( n23780 , n20722 );
and ( n23781 , n23779 , n23780 );
not ( n23782 , n23779 );
and ( n23783 , n23782 , n20722 );
nor ( n23784 , n23781 , n23783 );
buf ( n23785 , n23784 );
and ( n23786 , n23776 , n23785 );
nor ( n23787 , n23775 , n23786 );
buf ( n23788 , n14896 );
not ( n23789 , n23788 );
nor ( n23790 , n23787 , n23789 );
nor ( n23791 , n23773 , n23790 );
or ( n23792 , n23791 , n21697 );
nand ( n23793 , n21696 , n13849 );
nand ( n23794 , n23792 , n23793 );
buf ( n23795 , n23794 );
buf ( n23796 , n23795 );
not ( n23797 , n275550 );
buf ( n23798 , n23797 );
buf ( n23799 , n23798 );
not ( n23800 , n275929 );
buf ( n23801 , n23800 );
buf ( n23802 , n23801 );
not ( n23803 , n15902 );
or ( n23804 , n23803 , n14830 );
buf ( n23805 , n12863 );
not ( n23806 , n14830 );
not ( n23807 , n23806 );
nand ( n23808 , n23805 , n23807 );
nand ( n23809 , n23804 , n23808 );
buf ( n23810 , n23809 );
buf ( n23811 , n23810 );
not ( n23812 , n275550 );
buf ( n23813 , n23812 );
buf ( n23814 , n23813 );
buf ( n23815 , n275554 );
not ( n23816 , n275929 );
buf ( n23817 , n23816 );
buf ( n23818 , n23817 );
not ( n23819 , n275925 );
buf ( n23820 , n23819 );
buf ( n23821 , n23820 );
buf ( n23822 , n14336 );
and ( n23823 , n20711 , n23822 );
not ( n23824 , n20711 );
not ( n23825 , n14797 );
buf ( n23826 , n14782 );
not ( n23827 , n23826 );
not ( n23828 , n23827 );
or ( n23829 , n23825 , n23828 );
not ( n23830 , n23826 );
or ( n23831 , n23830 , n14797 );
nand ( n23832 , n23829 , n23831 );
buf ( n23833 , n23832 );
and ( n23834 , n23824 , n23833 );
nor ( n23835 , n23823 , n23834 );
not ( n23836 , n23835 );
and ( n23837 , n23836 , n23788 );
not ( n23838 , n20889 );
nand ( n23839 , n16916 , n16946 );
not ( n23840 , n23839 );
not ( n23841 , n16139 );
not ( n23842 , n16913 );
or ( n23843 , n23841 , n23842 );
not ( n23844 , n16943 );
nand ( n23845 , n23843 , n23844 );
not ( n23846 , n23845 );
or ( n23847 , n23840 , n23846 );
or ( n23848 , n23845 , n23839 );
nand ( n23849 , n23847 , n23848 );
buf ( n23850 , n23849 );
not ( n23851 , n23850 );
or ( n23852 , n23838 , n23851 );
not ( n23853 , n17097 );
nand ( n23854 , n23853 , n17393 );
not ( n23855 , n23854 );
not ( n23856 , n17090 );
not ( n23857 , n23856 );
not ( n23858 , n17362 );
or ( n23859 , n23857 , n23858 );
buf ( n23860 , n17389 );
nand ( n23861 , n23859 , n23860 );
not ( n23862 , n23861 );
or ( n23863 , n23855 , n23862 );
or ( n23864 , n23861 , n23854 );
nand ( n23865 , n23863 , n23864 );
buf ( n23866 , n23865 );
and ( n23867 , n23866 , n20926 );
not ( n23868 , n15557 );
not ( n23869 , n20940 );
or ( n23870 , n23868 , n23869 );
not ( n23871 , n17468 );
not ( n23872 , n17475 );
nand ( n23873 , n23872 , n17485 );
nor ( n23874 , n23871 , n23873 );
and ( n23875 , n20775 , n23874 );
not ( n23876 , n23875 );
nor ( n23877 , n17463 , n23876 );
or ( n23878 , n23877 , n17473 );
nand ( n23879 , n23877 , n17473 );
nand ( n23880 , n23878 , n23879 );
buf ( n23881 , n23880 );
nand ( n23882 , n23881 , n17409 );
nand ( n23883 , n23870 , n23882 );
nor ( n23884 , n23867 , n23883 );
nand ( n23885 , n23852 , n23884 );
nor ( n23886 , n23837 , n23885 );
buf ( n23887 , n20950 );
or ( n23888 , n23886 , n23887 );
nand ( n23889 , n23887 , n13955 );
nand ( n23890 , n23888 , n23889 );
buf ( n23891 , n23890 );
buf ( n23892 , n23891 );
and ( n23893 , n275557 , n19305 );
not ( n23894 , n275557 );
and ( n23895 , n23894 , n17586 );
or ( n23896 , n23893 , n23895 );
buf ( n23897 , n23896 );
buf ( n23898 , n23897 );
not ( n23899 , n275550 );
buf ( n23900 , n23899 );
buf ( n23901 , n23900 );
not ( n23902 , n275925 );
buf ( n23903 , n23902 );
buf ( n23904 , n23903 );
buf ( n23905 , n275554 );
not ( n23906 , n22798 );
not ( n23907 , n23906 );
buf ( n23908 , n18972 );
buf ( n23909 , n23908 );
not ( n23910 , n23909 );
buf ( n23911 , n23910 );
buf ( n23912 , n23911 );
not ( n23913 , n23912 );
buf ( n23914 , n21723 );
buf ( n23915 , n23914 );
not ( n23916 , n23915 );
buf ( n23917 , n23916 );
buf ( n23918 , n23917 );
not ( n23919 , n23918 );
or ( n23920 , n23913 , n23919 );
buf ( n23921 , n23911 );
not ( n23922 , n23921 );
buf ( n23923 , n23914 );
nand ( n23924 , n23922 , n23923 );
buf ( n23925 , n23924 );
buf ( n23926 , n23925 );
nand ( n23927 , n23920 , n23926 );
buf ( n23928 , n23927 );
buf ( n23929 , n23928 );
buf ( n23930 , n23929 );
not ( n23931 , n23930 );
not ( n23932 , n23931 );
and ( n23933 , n23907 , n23932 );
not ( n23934 , n23907 );
buf ( n23935 , n21726 );
buf ( n23936 , n18978 );
nand ( n23937 , n23935 , n23936 );
buf ( n23938 , n23937 );
buf ( n23939 , n23938 );
buf ( n23940 , n18629 );
buf ( n23941 , n23940 );
not ( n23942 , n23941 );
buf ( n23943 , n23942 );
buf ( n23944 , n23943 );
and ( n23945 , n23939 , n23944 );
not ( n23946 , n23939 );
buf ( n23947 , n23940 );
and ( n23948 , n23946 , n23947 );
nor ( n23949 , n23945 , n23948 );
buf ( n23950 , n23949 );
buf ( n23951 , n23950 );
buf ( n23952 , n23951 );
buf ( n23953 , n23952 );
not ( n23954 , n23953 );
buf ( n23955 , n23929 );
nand ( n23956 , n23955 , n21162 , n21112 );
not ( n23957 , n23956 );
and ( n23958 , n19069 , n23957 );
nand ( n23959 , n23958 , n21141 );
not ( n23960 , n23959 );
buf ( n23961 , n21726 );
buf ( n23962 , n23908 );
nand ( n23963 , n23961 , n23962 );
buf ( n23964 , n23963 );
buf ( n23965 , n23964 );
buf ( n23966 , n18949 );
buf ( n23967 , n23966 );
not ( n23968 , n23967 );
buf ( n23969 , n23968 );
buf ( n23970 , n23969 );
and ( n23971 , n23965 , n23970 );
not ( n23972 , n23965 );
buf ( n23973 , n23966 );
and ( n23974 , n23972 , n23973 );
nor ( n23975 , n23971 , n23974 );
buf ( n23976 , n23975 );
buf ( n23977 , n23976 );
buf ( n23978 , n23977 );
buf ( n23979 , n23978 );
not ( n23980 , n23979 );
not ( n23981 , n23980 );
nand ( n23982 , n23960 , n23981 );
not ( n23983 , n23982 );
or ( n23984 , n23954 , n23983 );
or ( n23985 , n23982 , n23953 );
nand ( n23986 , n23984 , n23985 );
buf ( n23987 , n23986 );
and ( n23988 , n23934 , n23987 );
nor ( n23989 , n23933 , n23988 );
not ( n23990 , n23989 );
not ( n23991 , n20987 );
not ( n23992 , n23991 );
and ( n23993 , n23990 , n23992 );
not ( n23994 , n21001 );
not ( n23995 , n17720 );
buf ( n23996 , n19235 );
not ( n23997 , n23996 );
or ( n23998 , n23995 , n23997 );
not ( n23999 , n277603 );
buf ( n24000 , n21244 );
buf ( n24001 , n19832 );
buf ( n24002 , n22565 );
not ( n24003 , n24002 );
buf ( n24004 , n24003 );
buf ( n24005 , n24004 );
buf ( n24006 , n19758 );
nor ( n24007 , n24005 , n24006 );
buf ( n24008 , n24007 );
buf ( n24009 , n24008 );
nand ( n24010 , n24000 , n24001 , n24009 );
buf ( n24011 , n24010 );
buf ( n24012 , n24011 );
buf ( n24013 , n21244 );
buf ( n24014 , n24004 );
buf ( n24015 , n21195 );
nor ( n24016 , n24014 , n24015 );
buf ( n24017 , n24016 );
buf ( n24018 , n24017 );
nand ( n24019 , n24013 , n24018 );
buf ( n24020 , n24019 );
buf ( n24021 , n24020 );
buf ( n24022 , n22565 );
buf ( n24023 , n22583 );
and ( n24024 , n24022 , n24023 );
buf ( n24025 , n22361 );
nor ( n24026 , n24024 , n24025 );
buf ( n24027 , n24026 );
buf ( n24028 , n24027 );
nand ( n24029 , n24012 , n24021 , n24028 );
buf ( n24030 , n24029 );
buf ( n24031 , n24030 );
buf ( n24032 , n22602 );
not ( n24033 , n24032 );
buf ( n24034 , n24033 );
buf ( n24035 , n24034 );
nand ( n24036 , n24031 , n24035 );
buf ( n24037 , n24036 );
buf ( n24038 , n24037 );
buf ( n24039 , n22606 );
buf ( n24040 , n22614 );
nand ( n24041 , n24039 , n24040 );
buf ( n24042 , n24041 );
buf ( n24043 , n24042 );
xnor ( n24044 , n24038 , n24043 );
buf ( n24045 , n24044 );
buf ( n24046 , n24045 );
not ( n24047 , n24046 );
or ( n24048 , n23999 , n24047 );
nand ( n24049 , n277351 , n9720 );
nand ( n24050 , n24048 , n24049 );
nand ( n24051 , n19242 , n24050 );
nand ( n24052 , n23998 , n24051 );
buf ( n24053 , n24052 );
not ( n24054 , n24053 );
buf ( n24055 , n18948 );
buf ( n24056 , n24055 );
not ( n24057 , n24056 );
or ( n24058 , n24054 , n24057 );
not ( n24059 , n24056 );
not ( n24060 , n24053 );
nand ( n24061 , n24059 , n24060 );
nand ( n24062 , n24058 , n24061 );
not ( n24063 , n17734 );
not ( n24064 , n23996 );
or ( n24065 , n24063 , n24064 );
not ( n24066 , n277603 );
buf ( n24067 , n22361 );
not ( n24068 , n24067 );
buf ( n24069 , n24034 );
nand ( n24070 , n24068 , n24069 );
buf ( n24071 , n24070 );
buf ( n24072 , n24071 );
not ( n24073 , n24072 );
buf ( n24074 , n22593 );
not ( n24075 , n24074 );
or ( n24076 , n24073 , n24075 );
buf ( n24077 , n22592 );
buf ( n24078 , n24071 );
or ( n24079 , n24077 , n24078 );
nand ( n24080 , n24076 , n24079 );
buf ( n24081 , n24080 );
buf ( n24082 , n24081 );
not ( n24083 , n24082 );
or ( n24084 , n24066 , n24083 );
nand ( n24085 , n277390 , n9728 );
nand ( n24086 , n24084 , n24085 );
nand ( n24087 , n19242 , n24086 );
nand ( n24088 , n24065 , n24087 );
buf ( n24089 , n24088 );
not ( n24090 , n24089 );
buf ( n24091 , n18971 );
buf ( n24092 , n24091 );
and ( n24093 , n24090 , n24092 );
nor ( n24094 , n24062 , n24093 );
not ( n24095 , n24094 );
nand ( n24096 , n24062 , n24093 );
nand ( n24097 , n24095 , n24096 );
not ( n24098 , n24097 );
not ( n24099 , n24089 );
not ( n24100 , n24092 );
or ( n24101 , n24099 , n24100 );
not ( n24102 , n24092 );
nand ( n24103 , n24102 , n24090 );
nand ( n24104 , n24101 , n24103 );
not ( n24105 , n17671 );
not ( n24106 , n24105 );
not ( n24107 , n19235 );
or ( n24108 , n24106 , n24107 );
not ( n24109 , n277527 );
buf ( n24110 , n21282 );
not ( n24111 , n24110 );
buf ( n24112 , n21215 );
nor ( n24113 , n24111 , n24112 );
buf ( n24114 , n24113 );
buf ( n24115 , n24114 );
buf ( n24116 , n21195 );
and ( n24117 , n24115 , n24116 );
buf ( n24118 , n24117 );
buf ( n24119 , n24118 );
not ( n24120 , n24119 );
buf ( n24121 , n19835 );
not ( n24122 , n24121 );
or ( n24123 , n24120 , n24122 );
buf ( n24124 , n21247 );
buf ( n24125 , n24114 );
and ( n24126 , n24124 , n24125 );
buf ( n24127 , n21282 );
not ( n24128 , n24127 );
buf ( n24129 , n21269 );
not ( n24130 , n24129 );
or ( n24131 , n24128 , n24130 );
buf ( n24132 , n21290 );
nand ( n24133 , n24131 , n24132 );
buf ( n24134 , n24133 );
buf ( n24135 , n24134 );
nor ( n24136 , n24126 , n24135 );
buf ( n24137 , n24136 );
buf ( n24138 , n24137 );
nand ( n24139 , n24123 , n24138 );
buf ( n24140 , n24139 );
buf ( n24141 , n24140 );
buf ( n24142 , n22493 );
buf ( n24143 , n22546 );
nand ( n24144 , n24142 , n24143 );
buf ( n24145 , n24144 );
buf ( n24146 , n24145 );
xnor ( n24147 , n24141 , n24146 );
buf ( n24148 , n24147 );
buf ( n24149 , n24148 );
not ( n24150 , n24149 );
or ( n24151 , n24109 , n24150 );
nand ( n24152 , n277351 , n9523 );
nand ( n24153 , n24151 , n24152 );
nand ( n24154 , n19242 , n24153 );
nand ( n24155 , n24108 , n24154 );
buf ( n24156 , n24155 );
not ( n24157 , n24156 );
buf ( n24158 , n18709 );
buf ( n24159 , n24158 );
and ( n24160 , n24157 , n24159 );
or ( n24161 , n24104 , n24160 );
not ( n24162 , n24161 );
nor ( n24163 , n20345 , n20262 );
nand ( n24164 , n24163 , n20255 );
not ( n24165 , n24164 );
not ( n24166 , n21362 );
not ( n24167 , n24157 );
not ( n24168 , n24159 );
not ( n24169 , n24168 );
or ( n24170 , n24167 , n24169 );
nand ( n24171 , n24159 , n24156 );
nand ( n24172 , n24170 , n24171 );
nand ( n24173 , n21305 , n21308 );
not ( n24174 , n24173 );
nor ( n24175 , n24172 , n24174 );
not ( n24176 , n24175 );
nand ( n24177 , n24166 , n24176 );
nor ( n24178 , n21469 , n24177 );
nand ( n24179 , n24178 , n21416 );
nor ( n24180 , n20345 , n20071 );
nor ( n24181 , n24179 , n24180 );
not ( n24182 , n24181 );
or ( n24183 , n24165 , n24182 );
nand ( n24184 , n19340 , n19325 );
nand ( n24185 , n20306 , n24184 );
nand ( n24186 , n20326 , n20314 );
nand ( n24187 , n24185 , n24186 , n20323 );
and ( n24188 , n20316 , n20253 , n21415 );
nand ( n24189 , n24187 , n24188 );
nor ( n24190 , n24175 , n21467 );
nor ( n24191 , n21457 , n21362 );
nand ( n24192 , n24190 , n20334 , n24191 , n20071 );
nor ( n24193 , n24189 , n24192 );
and ( n24194 , n24190 , n21490 , n21363 );
or ( n24195 , n24175 , n21359 );
nand ( n24196 , n24172 , n24174 );
nand ( n24197 , n24195 , n24196 );
nor ( n24198 , n24194 , n24197 );
nand ( n24199 , n24178 , n21483 );
nand ( n24200 , n24198 , n24199 );
nor ( n24201 , n24193 , n24200 );
nand ( n24202 , n24183 , n24201 );
not ( n24203 , n24202 );
not ( n24204 , n24203 );
not ( n24205 , n24204 );
or ( n24206 , n24162 , n24205 );
nand ( n24207 , n24104 , n24160 );
nand ( n24208 , n24206 , n24207 );
not ( n24209 , n24208 );
or ( n24210 , n24098 , n24209 );
or ( n24211 , n24208 , n24097 );
nand ( n24212 , n24210 , n24211 );
buf ( n24213 , n24212 );
not ( n24214 , n24213 );
or ( n24215 , n23994 , n24214 );
buf ( n24216 , n24088 );
not ( n24217 , n24216 );
not ( n24218 , n24217 );
buf ( n24219 , n24091 );
not ( n24220 , n24219 );
or ( n24221 , n24218 , n24220 );
not ( n24222 , n24219 );
nand ( n24223 , n24222 , n24216 );
nand ( n24224 , n24221 , n24223 );
buf ( n24225 , n24158 );
buf ( n24226 , n24155 );
and ( n24227 , n24225 , n24226 );
or ( n24228 , n24224 , n24227 );
not ( n24229 , n24228 );
not ( n24230 , n24225 );
not ( n24231 , n24230 );
not ( n24232 , n24226 );
or ( n24233 , n24231 , n24232 );
not ( n24234 , n24226 );
nand ( n24235 , n24234 , n24225 );
nand ( n24236 , n24233 , n24235 );
not ( n24237 , n24236 );
and ( n24238 , n21504 , n21502 );
not ( n24239 , n24238 );
nand ( n24240 , n24237 , n24239 );
not ( n24241 , n24240 );
nor ( n24242 , n21514 , n24241 );
not ( n24243 , n24242 );
not ( n24244 , n21585 );
or ( n24245 , n24243 , n24244 );
nand ( n24246 , n24236 , n24238 );
not ( n24247 , n24246 );
nor ( n24248 , n24241 , n21518 );
nor ( n24249 , n24247 , n24248 );
nand ( n24250 , n24245 , n24249 );
not ( n24251 , n24250 );
or ( n24252 , n24229 , n24251 );
nand ( n24253 , n24224 , n24227 );
nand ( n24254 , n24252 , n24253 );
not ( n24255 , n24254 );
nor ( n24256 , n21546 , n21514 );
and ( n24257 , n24256 , n21533 , n24240 );
nand ( n24258 , n21575 , n24257 );
not ( n24259 , n24258 );
nor ( n24260 , n20486 , n20496 );
not ( n24261 , n24260 );
not ( n24262 , n20424 );
nor ( n24263 , n20419 , n20422 );
not ( n24264 , n24263 );
or ( n24265 , n24262 , n24264 );
nor ( n24266 , n20450 , n20412 );
nand ( n24267 , n24265 , n24266 );
not ( n24268 , n24267 );
or ( n24269 , n24261 , n24268 );
nand ( n24270 , n20495 , n20475 );
and ( n24271 , n24270 , n24257 , n21562 );
nand ( n24272 , n24269 , n24271 );
not ( n24273 , n24272 );
or ( n24274 , n24259 , n24273 );
nand ( n24275 , n24274 , n24228 );
nand ( n24276 , n24255 , n24275 );
buf ( n24277 , n24052 );
not ( n24278 , n24277 );
not ( n24279 , n24278 );
buf ( n24280 , n24055 );
not ( n24281 , n24280 );
or ( n24282 , n24279 , n24281 );
not ( n24283 , n24280 );
nand ( n24284 , n24283 , n24277 );
nand ( n24285 , n24282 , n24284 );
and ( n24286 , n24219 , n24216 );
nor ( n24287 , n24285 , n24286 );
not ( n24288 , n24287 );
nand ( n24289 , n24285 , n24286 );
nand ( n24290 , n24288 , n24289 );
not ( n24291 , n24290 );
and ( n24292 , n24276 , n24291 );
not ( n24293 , n24276 );
and ( n24294 , n24293 , n24290 );
nor ( n24295 , n24292 , n24294 );
buf ( n24296 , n24295 );
and ( n24297 , n24296 , n19358 );
not ( n24298 , n19290 );
buf ( n24299 , n24052 );
buf ( n24300 , n24299 );
not ( n24301 , n24300 );
not ( n24302 , n24301 );
buf ( n24303 , n24088 );
buf ( n24304 , n24303 );
not ( n24305 , n24304 );
nor ( n24306 , n21610 , n21596 );
buf ( n24307 , n24155 );
buf ( n24308 , n24307 );
nor ( n24309 , n21608 , n24308 );
nand ( n24310 , n20529 , n24306 , n24309 );
nor ( n24311 , n21604 , n24310 );
nor ( n24312 , n20545 , n20537 );
nand ( n24313 , n24311 , n24312 );
not ( n24314 , n24313 );
nand ( n24315 , n24305 , n24314 );
not ( n24316 , n24315 );
or ( n24317 , n24302 , n24316 );
or ( n24318 , n24315 , n24301 );
nand ( n24319 , n24317 , n24318 );
buf ( n24320 , n24319 );
not ( n24321 , n24320 );
or ( n24322 , n24298 , n24321 );
buf ( n24323 , n24299 );
buf ( n24324 , n24323 );
buf ( n24325 , n24324 );
nand ( n24326 , n19219 , n24325 );
nand ( n24327 , n24322 , n24326 );
nor ( n24328 , n24297 , n24327 );
nand ( n24329 , n24215 , n24328 );
nor ( n24330 , n23993 , n24329 );
or ( n24331 , n24330 , n21030 );
nand ( n24332 , n21030 , n18940 );
nand ( n24333 , n24331 , n24332 );
buf ( n24334 , n24333 );
buf ( n24335 , n24334 );
buf ( n24336 , n275554 );
nand ( n24337 , n275736 , n275762 );
not ( n24338 , n24337 );
not ( n24339 , n275759 );
or ( n24340 , n24338 , n24339 );
or ( n24341 , n275759 , n24337 );
nand ( n24342 , n24340 , n24341 );
buf ( n24343 , n24342 );
buf ( n24344 , n24343 );
not ( n24345 , n275625 );
nand ( n24346 , n24345 , n275852 );
not ( n24347 , n24346 );
not ( n24348 , n275847 );
or ( n24349 , n24348 , n275644 );
nand ( n24350 , n24349 , n275850 );
not ( n24351 , n24350 );
or ( n24352 , n24347 , n24351 );
or ( n24353 , n24350 , n24346 );
nand ( n24354 , n24352 , n24353 );
buf ( n24355 , n24354 );
buf ( n24356 , n24355 );
or ( n24357 , n20844 , n20743 );
nand ( n24358 , n20885 , n16970 );
nand ( n24359 , n20924 , n17405 );
nand ( n24360 , n17411 , n20937 );
nand ( n24361 , n20785 , n20943 );
nand ( n24362 , n17562 , n13471 );
and ( n24363 , n17511 , n17512 );
not ( n24364 , n17511 );
and ( n24365 , n24364 , n13477 );
nor ( n24366 , n24363 , n24365 );
nand ( n24367 , n17545 , n24366 );
and ( n24368 , n24360 , n24361 , n24362 , n24367 );
and ( n24369 , n24358 , n24359 , n24368 );
nand ( n24370 , n24357 , n24369 );
buf ( n24371 , n24370 );
buf ( n24372 , n24371 );
not ( n24373 , n275925 );
buf ( n24374 , n24373 );
buf ( n24375 , n24374 );
buf ( n24376 , n275554 );
not ( n24377 , n275929 );
buf ( n24378 , n24377 );
buf ( n24379 , n24378 );
buf ( n24380 , n275554 );
buf ( n24381 , n275554 );
buf ( n24382 , n275554 );
not ( n24383 , n275929 );
buf ( n24384 , n24383 );
buf ( n24385 , n24384 );
buf ( n24386 , n19523 );
and ( n24387 , n22799 , n24386 );
not ( n24388 , n22799 );
buf ( n24389 , n19601 );
not ( n24390 , n24389 );
buf ( n24391 , n19581 );
and ( n24392 , n22805 , n24391 );
nand ( n24393 , n19069 , n24392 );
not ( n24394 , n24393 );
or ( n24395 , n24390 , n24394 );
or ( n24396 , n24393 , n24389 );
nand ( n24397 , n24395 , n24396 );
buf ( n24398 , n24397 );
and ( n24399 , n24388 , n24398 );
nor ( n24400 , n24387 , n24399 );
not ( n24401 , n24400 );
and ( n24402 , n24401 , n21174 );
not ( n24403 , n19358 );
nand ( n24404 , n20441 , n20485 );
not ( n24405 , n24404 );
not ( n24406 , n22823 );
not ( n24407 , n20449 );
or ( n24408 , n24406 , n24407 );
not ( n24409 , n20481 );
nand ( n24410 , n24408 , n24409 );
not ( n24411 , n24410 );
or ( n24412 , n24405 , n24411 );
or ( n24413 , n24410 , n24404 );
nand ( n24414 , n24412 , n24413 );
buf ( n24415 , n24414 );
not ( n24416 , n24415 );
or ( n24417 , n24403 , n24416 );
nand ( n24418 , n20194 , n20199 );
not ( n24419 , n24418 );
not ( n24420 , n20333 );
not ( n24421 , n22842 );
or ( n24422 , n24420 , n24421 );
not ( n24423 , n20152 );
nand ( n24424 , n24422 , n24423 );
not ( n24425 , n24424 );
or ( n24426 , n24419 , n24425 );
or ( n24427 , n24424 , n24418 );
nand ( n24428 , n24426 , n24427 );
buf ( n24429 , n24428 );
and ( n24430 , n24429 , n21001 );
not ( n24431 , n20532 );
nor ( n24432 , n20545 , n20535 );
not ( n24433 , n24432 );
or ( n24434 , n24431 , n24433 );
or ( n24435 , n24432 , n20532 );
nand ( n24436 , n24434 , n24435 );
buf ( n24437 , n24436 );
not ( n24438 , n24437 );
or ( n24439 , n24438 , n19289 );
not ( n24440 , n19219 );
buf ( n24441 , n20531 );
buf ( n24442 , n24441 );
not ( n24443 , n24442 );
or ( n24444 , n24440 , n24443 );
nand ( n24445 , n24439 , n24444 );
nor ( n24446 , n24430 , n24445 );
nand ( n24447 , n24417 , n24446 );
nor ( n24448 , n24402 , n24447 );
nand ( n24449 , n19143 , n19377 , n19175 );
or ( n24450 , n24449 , n19385 );
or ( n24451 , n24448 , n24450 );
buf ( n24452 , n24450 );
nand ( n24453 , n24452 , n18396 );
nand ( n24454 , n24451 , n24453 );
buf ( n24455 , n24454 );
buf ( n24456 , n24455 );
and ( n24457 , n13374 , n14795 );
not ( n24458 , n13374 );
not ( n24459 , n14798 );
nand ( n24460 , n24459 , n14058 );
buf ( n24461 , n13743 );
buf ( n24462 , n14014 );
buf ( n24463 , n14009 );
buf ( n24464 , n14045 );
nand ( n24465 , n24463 , n24464 );
buf ( n24466 , n24465 );
buf ( n24467 , n24466 );
nor ( n24468 , n24462 , n24467 );
buf ( n24469 , n24468 );
buf ( n24470 , n24469 );
nand ( n24471 , n24461 , n24470 );
buf ( n24472 , n24471 );
buf ( n24473 , n24472 );
buf ( n24474 , n14719 );
buf ( n24475 , n24474 );
not ( n24476 , n24475 );
buf ( n24477 , n24476 );
buf ( n24478 , n24477 );
and ( n24479 , n24473 , n24478 );
not ( n24480 , n24473 );
buf ( n24481 , n24474 );
and ( n24482 , n24480 , n24481 );
nor ( n24483 , n24479 , n24482 );
buf ( n24484 , n24483 );
buf ( n24485 , n24484 );
buf ( n24486 , n24485 );
not ( n24487 , n24486 );
and ( n24488 , n24460 , n24487 );
not ( n24489 , n24460 );
and ( n24490 , n24489 , n24486 );
nor ( n24491 , n24488 , n24490 );
buf ( n24492 , n24491 );
and ( n24493 , n24458 , n24492 );
nor ( n24494 , n24457 , n24493 );
not ( n24495 , n24494 );
and ( n24496 , n24495 , n23788 );
not ( n24497 , n20889 );
not ( n24498 , n16282 );
buf ( n24499 , n22215 );
not ( n24500 , n24499 );
buf ( n24501 , n22268 );
nand ( n24502 , n24500 , n24501 );
buf ( n24503 , n24502 );
buf ( n24504 , n24503 );
not ( n24505 , n24504 );
buf ( n24506 , n15387 );
buf ( n24507 , n15013 );
buf ( n24508 , n22223 );
and ( n24509 , n24507 , n24508 );
buf ( n24510 , n24509 );
buf ( n24511 , n24510 );
nand ( n24512 , n24506 , n24511 );
buf ( n24513 , n24512 );
buf ( n24514 , n24513 );
buf ( n24515 , n15481 );
buf ( n24516 , n22223 );
and ( n24517 , n24515 , n24516 );
buf ( n24518 , n22257 );
nor ( n24519 , n24517 , n24518 );
buf ( n24520 , n24519 );
buf ( n24521 , n24520 );
nand ( n24522 , n24514 , n24521 );
buf ( n24523 , n24522 );
buf ( n24524 , n24523 );
not ( n24525 , n24524 );
or ( n24526 , n24505 , n24525 );
buf ( n24527 , n24523 );
buf ( n24528 , n24503 );
or ( n24529 , n24527 , n24528 );
nand ( n24530 , n24526 , n24529 );
buf ( n24531 , n24530 );
buf ( n24532 , n24531 );
not ( n24533 , n24532 );
or ( n24534 , n24498 , n24533 );
nand ( n24535 , n277352 , n9752 );
nand ( n24536 , n24534 , n24535 );
nand ( n24537 , n15523 , n24536 );
not ( n24538 , n24537 );
buf ( n24539 , n24538 );
not ( n24540 , n24539 );
buf ( n24541 , n14043 );
buf ( n24542 , n24541 );
buf ( n24543 , n24542 );
not ( n24544 , n24543 );
or ( n24545 , n24540 , n24544 );
not ( n24546 , n24539 );
not ( n24547 , n24543 );
nand ( n24548 , n24546 , n24547 );
nand ( n24549 , n24545 , n24548 );
and ( n24550 , n15518 , n15514 );
or ( n24551 , n24549 , n24550 );
nand ( n24552 , n24549 , n24550 );
nand ( n24553 , n24551 , n24552 );
not ( n24554 , n24553 );
nor ( n24555 , n15564 , n16148 );
not ( n24556 , n24555 );
nor ( n24557 , n16140 , n24556 );
not ( n24558 , n24557 );
not ( n24559 , n16913 );
or ( n24560 , n24558 , n24559 );
not ( n24561 , n24555 );
not ( n24562 , n16943 );
or ( n24563 , n24561 , n24562 );
or ( n24564 , n15564 , n16946 );
nand ( n24565 , n24564 , n15566 );
not ( n24566 , n24565 );
nand ( n24567 , n24563 , n24566 );
not ( n24568 , n24567 );
nand ( n24569 , n24560 , n24568 );
not ( n24570 , n24569 );
or ( n24571 , n24554 , n24570 );
or ( n24572 , n24569 , n24553 );
nand ( n24573 , n24571 , n24572 );
buf ( n24574 , n24573 );
not ( n24575 , n24574 );
or ( n24576 , n24497 , n24575 );
buf ( n24577 , n24542 );
not ( n24578 , n24577 );
buf ( n24579 , n24538 );
nand ( n24580 , n24578 , n24579 );
not ( n24581 , n24579 );
nand ( n24582 , n24581 , n24577 );
nand ( n24583 , n24580 , n24582 );
and ( n24584 , n16972 , n16973 );
nor ( n24585 , n24583 , n24584 );
not ( n24586 , n24585 );
nand ( n24587 , n24583 , n24584 );
nand ( n24588 , n24586 , n24587 );
not ( n24589 , n24588 );
nor ( n24590 , n17097 , n16979 );
not ( n24591 , n24590 );
nor ( n24592 , n17090 , n24591 );
not ( n24593 , n24592 );
not ( n24594 , n17362 );
or ( n24595 , n24593 , n24594 );
not ( n24596 , n17389 );
not ( n24597 , n24591 );
and ( n24598 , n24596 , n24597 );
or ( n24599 , n16979 , n17393 );
nand ( n24600 , n24599 , n16981 );
nor ( n24601 , n24598 , n24600 );
nand ( n24602 , n24595 , n24601 );
not ( n24603 , n24602 );
or ( n24604 , n24589 , n24603 );
or ( n24605 , n24602 , n24588 );
nand ( n24606 , n24604 , n24605 );
buf ( n24607 , n24606 );
and ( n24608 , n24607 , n20926 );
and ( n24609 , n20774 , n17489 );
and ( n24610 , n17462 , n24609 );
nor ( n24611 , n17492 , n17484 );
and ( n24612 , n17468 , n17476 , n24611 , n17479 );
nand ( n24613 , n24610 , n24612 );
buf ( n24614 , n24538 );
not ( n24615 , n24614 );
xnor ( n24616 , n24613 , n24615 );
buf ( n24617 , n24616 );
nand ( n24618 , n24617 , n17409 );
nand ( n24619 , n20940 , n24538 );
nand ( n24620 , n24618 , n24619 );
nor ( n24621 , n24608 , n24620 );
nand ( n24622 , n24576 , n24621 );
nor ( n24623 , n24496 , n24622 );
or ( n24624 , n24623 , n23887 );
nand ( n24625 , n20953 , n14039 );
nand ( n24626 , n24624 , n24625 );
buf ( n24627 , n24626 );
buf ( n24628 , n24627 );
buf ( n24629 , n275554 );
buf ( n24630 , n275554 );
not ( n24631 , n19094 );
not ( n24632 , n19069 );
not ( n24633 , n24632 );
or ( n24634 , n24631 , n24633 );
not ( n24635 , n19094 );
nand ( n24636 , n19069 , n24635 );
nand ( n24637 , n24634 , n24636 );
buf ( n24638 , n24637 );
nand ( n24639 , n24638 , n23906 );
or ( n24640 , n24639 , n19216 );
not ( n24641 , n19291 );
not ( n24642 , n19220 );
or ( n24643 , n24641 , n24642 );
buf ( n24644 , n19308 );
buf ( n24645 , n24644 );
buf ( n24646 , n24645 );
nand ( n24647 , n24643 , n24646 );
not ( n24648 , n19324 );
not ( n24649 , n19321 );
or ( n24650 , n24648 , n24649 );
or ( n24651 , n19321 , n19324 );
nand ( n24652 , n24650 , n24651 );
buf ( n24653 , n24652 );
and ( n24654 , n19354 , n24653 );
and ( n24655 , n19318 , n18283 );
nor ( n24656 , n24654 , n24655 );
not ( n24657 , n19362 );
not ( n24658 , n24657 );
not ( n24659 , n19361 );
or ( n24660 , n24658 , n24659 );
or ( n24661 , n19361 , n24657 );
nand ( n24662 , n24660 , n24661 );
buf ( n24663 , n24662 );
nand ( n24664 , n19360 , n24663 );
nand ( n24665 , n19387 , n18306 );
and ( n24666 , n24647 , n24656 , n24664 , n24665 );
nand ( n24667 , n24640 , n24666 );
buf ( n24668 , n24667 );
buf ( n24669 , n24668 );
buf ( n24670 , n275554 );
buf ( n24671 , n275554 );
buf ( n24672 , n14580 );
and ( n24673 , n13373 , n24672 );
not ( n24674 , n13373 );
not ( n24675 , n20827 );
buf ( n24676 , n20826 );
not ( n24677 , n24676 );
or ( n24678 , n24675 , n24677 );
or ( n24679 , n24676 , n20827 );
nand ( n24680 , n24678 , n24679 );
buf ( n24681 , n24680 );
and ( n24682 , n24674 , n24681 );
nor ( n24683 , n24673 , n24682 );
not ( n24684 , n24683 );
not ( n24685 , n23789 );
and ( n24686 , n24684 , n24685 );
nand ( n24687 , n16497 , n16489 );
not ( n24688 , n24687 );
not ( n24689 , n16874 );
buf ( n24690 , n16865 );
nand ( n24691 , n24689 , n24690 );
not ( n24692 , n24691 );
or ( n24693 , n24688 , n24692 );
or ( n24694 , n24691 , n24687 );
nand ( n24695 , n24693 , n24694 );
buf ( n24696 , n24695 );
nand ( n24697 , n24696 , n20889 );
not ( n24698 , n17179 );
buf ( n24699 , n17172 );
nand ( n24700 , n24698 , n24699 );
not ( n24701 , n24700 );
buf ( n24702 , n20908 );
not ( n24703 , n24702 );
buf ( n24704 , n17316 );
nand ( n24705 , n24703 , n24704 );
not ( n24706 , n24705 );
or ( n24707 , n24701 , n24706 );
or ( n24708 , n24705 , n24700 );
nand ( n24709 , n24707 , n24708 );
buf ( n24710 , n24709 );
not ( n24711 , n20925 );
nand ( n24712 , n24710 , n24711 );
not ( n24713 , n17420 );
not ( n24714 , n17433 );
nor ( n24715 , n24714 , n17415 );
not ( n24716 , n24715 );
or ( n24717 , n24713 , n24716 );
or ( n24718 , n24715 , n17420 );
nand ( n24719 , n24717 , n24718 );
buf ( n24720 , n24719 );
and ( n24721 , n24720 , n17409 );
buf ( n24722 , n17419 );
buf ( n24723 , n24722 );
buf ( n24724 , n24723 );
and ( n24725 , n20940 , n24724 );
nor ( n24726 , n24721 , n24725 );
nand ( n24727 , n24697 , n24712 , n24726 );
nor ( n24728 , n24686 , n24727 );
or ( n24729 , n24728 , n21696 );
nand ( n24730 , n21696 , n13589 );
nand ( n24731 , n24729 , n24730 );
buf ( n24732 , n24731 );
buf ( n24733 , n24732 );
and ( n24734 , n17562 , n14675 );
not ( n24735 , n17562 );
buf ( n24736 , n14759 );
buf ( n24737 , n24736 );
buf ( n24738 , n24737 );
not ( n24739 , n24738 );
not ( n24740 , n14798 );
or ( n24741 , n24739 , n24740 );
buf ( n24742 , n13743 );
buf ( n24743 , n14014 );
buf ( n24744 , n14722 );
not ( n24745 , n24744 );
buf ( n24746 , n14009 );
nand ( n24747 , n24745 , n24746 );
buf ( n24748 , n24747 );
buf ( n24749 , n24748 );
nor ( n24750 , n24743 , n24749 );
buf ( n24751 , n24750 );
buf ( n24752 , n24751 );
nand ( n24753 , n24742 , n24752 );
buf ( n24754 , n24753 );
buf ( n24755 , n24754 );
buf ( n24756 , n14650 );
buf ( n24757 , n24756 );
not ( n24758 , n24757 );
buf ( n24759 , n24758 );
buf ( n24760 , n24759 );
and ( n24761 , n24755 , n24760 );
not ( n24762 , n24755 );
buf ( n24763 , n24756 );
and ( n24764 , n24762 , n24763 );
nor ( n24765 , n24761 , n24764 );
buf ( n24766 , n24765 );
buf ( n24767 , n24766 );
buf ( n24768 , n24767 );
buf ( n24769 , n13743 );
buf ( n24770 , n14014 );
buf ( n24771 , n24748 );
buf ( n24772 , n24759 );
nor ( n24773 , n24770 , n24771 , n24772 );
buf ( n24774 , n24773 );
buf ( n24775 , n24774 );
nand ( n24776 , n24769 , n24775 );
buf ( n24777 , n24776 );
buf ( n24778 , n24777 );
buf ( n24779 , n14665 );
buf ( n24780 , n24779 );
not ( n24781 , n24780 );
buf ( n24782 , n24781 );
buf ( n24783 , n24782 );
and ( n24784 , n24778 , n24783 );
not ( n24785 , n24778 );
buf ( n24786 , n24779 );
and ( n24787 , n24785 , n24786 );
nor ( n24788 , n24784 , n24787 );
buf ( n24789 , n24788 );
buf ( n24790 , n24789 );
buf ( n24791 , n24790 );
and ( n24792 , n24768 , n24791 );
buf ( n24793 , n14684 );
buf ( n24794 , n24793 );
not ( n24795 , n24794 );
buf ( n24796 , n14158 );
buf ( n24797 , n24748 );
buf ( n24798 , n13935 );
buf ( n24799 , n14668 );
nor ( n24800 , n24797 , n24798 , n24799 );
buf ( n24801 , n24800 );
buf ( n24802 , n24801 );
nand ( n24803 , n24796 , n24802 );
buf ( n24804 , n24803 );
buf ( n24805 , n24804 );
not ( n24806 , n24805 );
or ( n24807 , n24795 , n24806 );
buf ( n24808 , n24804 );
buf ( n24809 , n24793 );
or ( n24810 , n24808 , n24809 );
nand ( n24811 , n24807 , n24810 );
buf ( n24812 , n24811 );
buf ( n24813 , n24812 );
buf ( n24814 , n24813 );
buf ( n24815 , n24814 );
buf ( n24816 , n24815 );
nand ( n24817 , n24792 , n24816 );
and ( n24818 , n24817 , n24738 );
not ( n24819 , n24738 );
not ( n24820 , n14059 );
or ( n24821 , n24819 , n24820 );
nand ( n24822 , n24487 , n24738 );
nand ( n24823 , n24821 , n24822 );
nor ( n24824 , n24818 , n24823 );
nand ( n24825 , n24741 , n24824 );
not ( n24826 , n24825 );
not ( n24827 , n24738 );
nand ( n24828 , n24827 , n14058 , n24486 );
nor ( n24829 , n24817 , n24828 );
nand ( n24830 , n14799 , n24829 );
nand ( n24831 , n24826 , n24830 );
buf ( n24832 , n24831 );
or ( n24833 , n13373 , n14847 );
buf ( n24834 , n15523 );
nand ( n24835 , n24833 , n24834 );
and ( n24836 , n23788 , n24835 );
nand ( n24837 , n24832 , n24836 );
not ( n24838 , n277910 );
buf ( n24839 , n22208 );
buf ( n24840 , n22275 );
or ( n24841 , n24839 , n24840 );
buf ( n24842 , n24841 );
buf ( n24843 , n24842 );
not ( n24844 , n24843 );
buf ( n24845 , n15013 );
buf ( n24846 , n22223 );
not ( n24847 , n24846 );
buf ( n24848 , n22215 );
nor ( n24849 , n24847 , n24848 );
buf ( n24850 , n24849 );
buf ( n24851 , n24850 );
and ( n24852 , n24845 , n24851 );
buf ( n24853 , n24852 );
buf ( n24854 , n24853 );
not ( n24855 , n24854 );
buf ( n24856 , n15387 );
not ( n24857 , n24856 );
or ( n24858 , n24855 , n24857 );
buf ( n24859 , n15481 );
buf ( n24860 , n24850 );
and ( n24861 , n24859 , n24860 );
buf ( n24862 , n22257 );
not ( n24863 , n24862 );
buf ( n24864 , n24863 );
buf ( n24865 , n24864 );
buf ( n24866 , n22215 );
or ( n24867 , n24865 , n24866 );
buf ( n24868 , n22268 );
nand ( n24869 , n24867 , n24868 );
buf ( n24870 , n24869 );
buf ( n24871 , n24870 );
nor ( n24872 , n24861 , n24871 );
buf ( n24873 , n24872 );
buf ( n24874 , n24873 );
nand ( n24875 , n24858 , n24874 );
buf ( n24876 , n24875 );
buf ( n24877 , n24876 );
not ( n24878 , n24877 );
or ( n24879 , n24844 , n24878 );
buf ( n24880 , n24876 );
buf ( n24881 , n24842 );
or ( n24882 , n24880 , n24881 );
nand ( n24883 , n24879 , n24882 );
buf ( n24884 , n24883 );
buf ( n24885 , n24884 );
not ( n24886 , n24885 );
or ( n24887 , n24838 , n24886 );
nand ( n24888 , n277527 , n9744 );
nand ( n24889 , n24887 , n24888 );
nand ( n24890 , n14920 , n24889 );
not ( n24891 , n24890 );
buf ( n24892 , n24891 );
not ( n24893 , n24892 );
not ( n24894 , n17473 );
not ( n24895 , n17492 );
nand ( n24896 , n24893 , n24894 , n24895 , n24615 );
not ( n24897 , n24896 );
not ( n24898 , n277910 );
buf ( n24899 , n22233 );
buf ( n24900 , n22288 );
nand ( n24901 , n24899 , n24900 );
buf ( n24902 , n24901 );
buf ( n24903 , n24902 );
not ( n24904 , n24903 );
buf ( n24905 , n15013 );
buf ( n24906 , n22226 );
and ( n24907 , n24905 , n24906 );
buf ( n24908 , n24907 );
buf ( n24909 , n24908 );
not ( n24910 , n24909 );
buf ( n24911 , n15387 );
not ( n24912 , n24911 );
or ( n24913 , n24910 , n24912 );
buf ( n24914 , n15481 );
buf ( n24915 , n22226 );
and ( n24916 , n24914 , n24915 );
buf ( n24917 , n22281 );
nor ( n24918 , n24916 , n24917 );
buf ( n24919 , n24918 );
buf ( n24920 , n24919 );
nand ( n24921 , n24913 , n24920 );
buf ( n24922 , n24921 );
buf ( n24923 , n24922 );
not ( n24924 , n24923 );
or ( n24925 , n24904 , n24924 );
buf ( n24926 , n24922 );
buf ( n24927 , n24902 );
or ( n24928 , n24926 , n24927 );
nand ( n24929 , n24925 , n24928 );
buf ( n24930 , n24929 );
buf ( n24931 , n24930 );
not ( n24932 , n24931 );
or ( n24933 , n24898 , n24932 );
nand ( n24934 , n277352 , n9787 );
nand ( n24935 , n24933 , n24934 );
nand ( n24936 , n24834 , n24935 );
not ( n24937 , n24936 );
buf ( n24938 , n24937 );
and ( n24939 , n24834 , n22327 );
buf ( n24940 , n24939 );
nor ( n24941 , n24938 , n24940 );
nand ( n24942 , n24897 , n24941 );
nor ( n24943 , n23876 , n24942 );
nand ( n24944 , n23436 , n24943 );
not ( n24945 , n16282 );
buf ( n24946 , n15013 );
buf ( n24947 , n22226 );
buf ( n24948 , n22233 );
not ( n24949 , n24948 );
buf ( n24950 , n22304 );
nor ( n24951 , n24949 , n24950 );
buf ( n24952 , n24951 );
buf ( n24953 , n24952 );
and ( n24954 , n24947 , n24953 );
buf ( n24955 , n24954 );
buf ( n24956 , n24955 );
and ( n24957 , n24946 , n24956 );
buf ( n24958 , n24957 );
buf ( n24959 , n24958 );
not ( n24960 , n24959 );
buf ( n24961 , n15387 );
not ( n24962 , n24961 );
or ( n24963 , n24960 , n24962 );
buf ( n24964 , n15481 );
buf ( n24965 , n24955 );
and ( n24966 , n24964 , n24965 );
buf ( n24967 , n24952 );
not ( n24968 , n24967 );
buf ( n24969 , n22281 );
not ( n24970 , n24969 );
or ( n24971 , n24968 , n24970 );
buf ( n24972 , n22304 );
not ( n24973 , n24972 );
buf ( n24974 , n22288 );
not ( n24975 , n24974 );
and ( n24976 , n24973 , n24975 );
buf ( n24977 , n22309 );
nor ( n24978 , n24976 , n24977 );
buf ( n24979 , n24978 );
buf ( n24980 , n24979 );
nand ( n24981 , n24971 , n24980 );
buf ( n24982 , n24981 );
buf ( n24983 , n24982 );
nor ( n24984 , n24966 , n24983 );
buf ( n24985 , n24984 );
buf ( n24986 , n24985 );
nand ( n24987 , n24963 , n24986 );
buf ( n24988 , n24987 );
buf ( n24989 , n24988 );
buf ( n24990 , n277340 );
buf ( n24991 , n24990 );
buf ( n24992 , n277353 );
buf ( n24993 , n24992 );
nor ( n24994 , n24991 , n24993 );
buf ( n24995 , n24994 );
buf ( n24996 , n24995 );
not ( n24997 , n24996 );
buf ( n24998 , n24990 );
buf ( n24999 , n24992 );
nand ( n25000 , n24998 , n24999 );
buf ( n25001 , n25000 );
buf ( n25002 , n25001 );
nand ( n25003 , n24997 , n25002 );
buf ( n25004 , n25003 );
buf ( n25005 , n25004 );
not ( n25006 , n25005 );
buf ( n25007 , n25006 );
buf ( n25008 , n25007 );
and ( n25009 , n24989 , n25008 );
not ( n25010 , n24989 );
buf ( n25011 , n25004 );
and ( n25012 , n25010 , n25011 );
nor ( n25013 , n25009 , n25012 );
buf ( n25014 , n25013 );
buf ( n25015 , n25014 );
not ( n25016 , n25015 );
or ( n25017 , n24945 , n25016 );
nand ( n25018 , n277603 , n277340 );
nand ( n25019 , n25017 , n25018 );
and ( n25020 , n24834 , n25019 );
buf ( n25021 , n25020 );
and ( n25022 , n24944 , n25021 );
not ( n25023 , n24944 );
not ( n25024 , n25021 );
and ( n25025 , n25023 , n25024 );
nor ( n25026 , n25022 , n25025 );
buf ( n25027 , n25026 );
and ( n25028 , n25027 , n17409 );
and ( n25029 , n20940 , n25020 );
nor ( n25030 , n25028 , n25029 );
and ( n25031 , n24837 , n25030 );
and ( n25032 , n24735 , n25031 );
nor ( n25033 , n24734 , n25032 );
buf ( n25034 , n25033 );
buf ( n25035 , n25034 );
buf ( n25036 , n275554 );
not ( n25037 , n275549 );
not ( n25038 , n25037 );
buf ( n25039 , n25038 );
buf ( n25040 , n25039 );
not ( n25041 , n275925 );
buf ( n25042 , n25041 );
buf ( n25043 , n25042 );
buf ( n25044 , n275554 );
nand ( n25045 , n19140 , n19639 );
nand ( n25046 , n19200 , n25045 );
not ( n25047 , n19134 );
nand ( n25048 , n25047 , n25045 );
buf ( n25049 , n19242 );
not ( n25050 , n25049 );
not ( n25051 , n25050 );
and ( n25052 , n25046 , n25048 , n25051 );
not ( n25053 , n18189 );
not ( n25054 , n18178 );
or ( n25055 , n25053 , n25054 );
or ( n25056 , n18178 , n18189 );
nand ( n25057 , n25055 , n25056 );
nand ( n25058 , n25052 , n25057 );
not ( n25059 , n21766 );
and ( n25060 , n19124 , n19141 );
nand ( n25061 , n25059 , n25060 );
and ( n25062 , n25058 , n25061 );
nor ( n25063 , n25062 , n18208 );
buf ( n25064 , n25063 );
buf ( n25065 , n17670 );
not ( n25066 , n25065 );
not ( n25067 , n25066 );
nand ( n25068 , n25064 , n25067 );
buf ( n25069 , n25065 );
buf ( n25070 , n25069 );
buf ( n25071 , n18701 );
buf ( n25072 , n25071 );
nand ( n25073 , n25070 , n25072 );
buf ( n25074 , n25073 );
buf ( n25075 , n25074 );
not ( n25076 , n25075 );
buf ( n25077 , n25069 );
buf ( n25078 , n25071 );
nor ( n25079 , n25077 , n25078 );
buf ( n25080 , n25079 );
buf ( n25081 , n25080 );
nor ( n25082 , n25076 , n25081 );
buf ( n25083 , n25082 );
buf ( n25084 , n25083 );
not ( n25085 , n25084 );
buf ( n25086 , n17895 );
buf ( n25087 , n25086 );
buf ( n25088 , n25087 );
buf ( n25089 , n25088 );
buf ( n25090 , n18744 );
buf ( n25091 , n25090 );
nor ( n25092 , n25089 , n25091 );
buf ( n25093 , n25092 );
buf ( n25094 , n25093 );
buf ( n25095 , n17768 );
buf ( n25096 , n25095 );
buf ( n25097 , n25096 );
buf ( n25098 , n25097 );
buf ( n25099 , n25098 );
buf ( n25100 , n18760 );
buf ( n25101 , n25100 );
nor ( n25102 , n25099 , n25101 );
buf ( n25103 , n25102 );
buf ( n25104 , n25103 );
nor ( n25105 , n25094 , n25104 );
buf ( n25106 , n25105 );
buf ( n25107 , n25106 );
buf ( n25108 , n17752 );
buf ( n25109 , n25108 );
buf ( n25110 , n25109 );
buf ( n25111 , n25110 );
buf ( n25112 , n18402 );
buf ( n25113 , n25112 );
or ( n25114 , n25111 , n25113 );
buf ( n25115 , n25114 );
buf ( n25116 , n25115 );
not ( n25117 , n25116 );
buf ( n25118 , n17780 );
buf ( n25119 , n25118 );
buf ( n25120 , n25119 );
buf ( n25121 , n25120 );
buf ( n25122 , n18335 );
buf ( n25123 , n25122 );
nor ( n25124 , n25121 , n25123 );
buf ( n25125 , n25124 );
buf ( n25126 , n25125 );
nor ( n25127 , n25117 , n25126 );
buf ( n25128 , n25127 );
buf ( n25129 , n25128 );
and ( n25130 , n25107 , n25129 );
buf ( n25131 , n25130 );
buf ( n25132 , n25131 );
buf ( n25133 , n17795 );
buf ( n25134 , n25133 );
buf ( n25135 , n25134 );
buf ( n25136 , n18878 );
buf ( n25137 , n25136 );
nor ( n25138 , n25135 , n25137 );
buf ( n25139 , n25138 );
buf ( n25140 , n25139 );
buf ( n25141 , n18086 );
buf ( n25142 , n25141 );
buf ( n25143 , n25142 );
buf ( n25144 , n25143 );
buf ( n25145 , n18908 );
buf ( n25146 , n25145 );
nor ( n25147 , n25144 , n25146 );
buf ( n25148 , n25147 );
buf ( n25149 , n25148 );
nor ( n25150 , n25140 , n25149 );
buf ( n25151 , n25150 );
buf ( n25152 , n25151 );
not ( n25153 , n25152 );
not ( n25154 , n18101 );
not ( n25155 , n25154 );
buf ( n25156 , n25155 );
buf ( n25157 , n25156 );
buf ( n25158 , n18383 );
buf ( n25159 , n25158 );
nor ( n25160 , n25157 , n25159 );
buf ( n25161 , n25160 );
buf ( n25162 , n25161 );
buf ( n25163 , n18054 );
buf ( n25164 , n25163 );
buf ( n25165 , n25164 );
buf ( n25166 , n25165 );
buf ( n25167 , n18356 );
buf ( n25168 , n25167 );
nor ( n25169 , n25166 , n25168 );
buf ( n25170 , n25169 );
buf ( n25171 , n25170 );
nor ( n25172 , n25162 , n25171 );
buf ( n25173 , n25172 );
buf ( n25174 , n25173 );
buf ( n25175 , n18071 );
buf ( n25176 , n25175 );
buf ( n25177 , n18866 );
buf ( n25178 , n25177 );
nor ( n25179 , n25176 , n25178 );
buf ( n25180 , n25179 );
buf ( n25181 , n25180 );
buf ( n25182 , n18306 );
not ( n25183 , n18133 );
buf ( n25184 , n25183 );
buf ( n25185 , n25184 );
and ( n25186 , n25182 , n25185 );
buf ( n25187 , n25186 );
buf ( n25188 , n25187 );
buf ( n25189 , n19083 );
xor ( n25190 , n25188 , n25189 );
buf ( n25191 , n18131 );
and ( n25192 , n25190 , n25191 );
and ( n25193 , n25188 , n25189 );
or ( n25194 , n25192 , n25193 );
buf ( n25195 , n25194 );
buf ( n25196 , n25195 );
buf ( n25197 , n18115 );
buf ( n25198 , n25197 );
buf ( n25199 , n18327 );
buf ( n25200 , n25199 );
or ( n25201 , n25198 , n25200 );
buf ( n25202 , n25201 );
buf ( n25203 , n25202 );
nand ( n25204 , n25196 , n25203 );
buf ( n25205 , n25204 );
buf ( n25206 , n25205 );
or ( n25207 , n25181 , n25206 );
buf ( n25208 , n25180 );
buf ( n25209 , n25197 );
buf ( n25210 , n25199 );
nand ( n25211 , n25209 , n25210 );
buf ( n25212 , n25211 );
buf ( n25213 , n25212 );
or ( n25214 , n25208 , n25213 );
buf ( n25215 , n25175 );
buf ( n25216 , n25177 );
nand ( n25217 , n25215 , n25216 );
buf ( n25218 , n25217 );
buf ( n25219 , n25218 );
nand ( n25220 , n25207 , n25214 , n25219 );
buf ( n25221 , n25220 );
buf ( n25222 , n25221 );
and ( n25223 , n25174 , n25222 );
buf ( n25224 , n25223 );
buf ( n25225 , n25224 );
not ( n25226 , n25225 );
or ( n25227 , n25153 , n25226 );
buf ( n25228 , n25151 );
buf ( n25229 , n25161 );
buf ( n25230 , n25165 );
buf ( n25231 , n25167 );
nand ( n25232 , n25230 , n25231 );
buf ( n25233 , n25232 );
buf ( n25234 , n25233 );
or ( n25235 , n25229 , n25234 );
buf ( n25236 , n25156 );
buf ( n25237 , n25158 );
nand ( n25238 , n25236 , n25237 );
buf ( n25239 , n25238 );
buf ( n25240 , n25239 );
nand ( n25241 , n25235 , n25240 );
buf ( n25242 , n25241 );
buf ( n25243 , n25242 );
and ( n25244 , n25228 , n25243 );
buf ( n25245 , n25139 );
buf ( n25246 , n25143 );
buf ( n25247 , n25145 );
nand ( n25248 , n25246 , n25247 );
buf ( n25249 , n25248 );
buf ( n25250 , n25249 );
or ( n25251 , n25245 , n25250 );
buf ( n25252 , n25134 );
buf ( n25253 , n25136 );
nand ( n25254 , n25252 , n25253 );
buf ( n25255 , n25254 );
buf ( n25256 , n25255 );
nand ( n25257 , n25251 , n25256 );
buf ( n25258 , n25257 );
buf ( n25259 , n25258 );
nor ( n25260 , n25244 , n25259 );
buf ( n25261 , n25260 );
buf ( n25262 , n25261 );
nand ( n25263 , n25227 , n25262 );
buf ( n25264 , n25263 );
buf ( n25265 , n25264 );
buf ( n25266 , n17928 );
buf ( n25267 , n25266 );
buf ( n25268 , n25267 );
buf ( n25269 , n25268 );
buf ( n25270 , n18987 );
buf ( n25271 , n25270 );
nor ( n25272 , n25269 , n25271 );
buf ( n25273 , n25272 );
buf ( n25274 , n25273 );
buf ( n25275 , n17942 );
buf ( n25276 , n25275 );
buf ( n25277 , n25276 );
buf ( n25278 , n25277 );
buf ( n25279 , n19010 );
buf ( n25280 , n25279 );
nor ( n25281 , n25278 , n25280 );
buf ( n25282 , n25281 );
buf ( n25283 , n25282 );
nor ( n25284 , n25274 , n25283 );
buf ( n25285 , n25284 );
buf ( n25286 , n25285 );
buf ( n25287 , n17912 );
buf ( n25288 , n25287 );
buf ( n25289 , n25288 );
buf ( n25290 , n25289 );
buf ( n25291 , n18731 );
buf ( n25292 , n25291 );
nor ( n25293 , n25290 , n25292 );
buf ( n25294 , n25293 );
buf ( n25295 , n25294 );
not ( n25296 , n25295 );
buf ( n25297 , n25296 );
buf ( n25298 , n25297 );
and ( n25299 , n25286 , n25298 );
buf ( n25300 , n25299 );
buf ( n25301 , n25300 );
and ( n25302 , n25132 , n25265 , n25301 );
buf ( n25303 , n25300 );
not ( n25304 , n25303 );
buf ( n25305 , n25093 );
buf ( n25306 , n25098 );
buf ( n25307 , n25100 );
nand ( n25308 , n25306 , n25307 );
buf ( n25309 , n25308 );
buf ( n25310 , n25309 );
or ( n25311 , n25305 , n25310 );
buf ( n25312 , n25106 );
buf ( n25313 , n25120 );
buf ( n25314 , n25122 );
nand ( n25315 , n25313 , n25314 );
buf ( n25316 , n25315 );
buf ( n25317 , n25316 );
not ( n25318 , n25317 );
buf ( n25319 , n25115 );
nand ( n25320 , n25318 , n25319 );
buf ( n25321 , n25320 );
buf ( n25322 , n25321 );
buf ( n25323 , n25110 );
buf ( n25324 , n25112 );
nand ( n25325 , n25323 , n25324 );
buf ( n25326 , n25325 );
buf ( n25327 , n25326 );
nand ( n25328 , n25322 , n25327 );
buf ( n25329 , n25328 );
buf ( n25330 , n25329 );
nand ( n25331 , n25312 , n25330 );
buf ( n25332 , n25331 );
buf ( n25333 , n25332 );
buf ( n25334 , n25088 );
buf ( n25335 , n25090 );
nand ( n25336 , n25334 , n25335 );
buf ( n25337 , n25336 );
buf ( n25338 , n25337 );
nand ( n25339 , n25311 , n25333 , n25338 );
buf ( n25340 , n25339 );
buf ( n25341 , n25340 );
not ( n25342 , n25341 );
or ( n25343 , n25304 , n25342 );
buf ( n25344 , n25273 );
buf ( n25345 , n25277 );
buf ( n25346 , n25279 );
nand ( n25347 , n25345 , n25346 );
buf ( n25348 , n25347 );
buf ( n25349 , n25348 );
or ( n25350 , n25344 , n25349 );
buf ( n25351 , n25268 );
buf ( n25352 , n25270 );
nand ( n25353 , n25351 , n25352 );
buf ( n25354 , n25353 );
buf ( n25355 , n25354 );
nand ( n25356 , n25350 , n25355 );
buf ( n25357 , n25356 );
buf ( n25358 , n25357 );
buf ( n25359 , n25297 );
and ( n25360 , n25358 , n25359 );
buf ( n25361 , n25289 );
buf ( n25362 , n25291 );
nand ( n25363 , n25361 , n25362 );
buf ( n25364 , n25363 );
buf ( n25365 , n25364 );
not ( n25366 , n25365 );
buf ( n25367 , n25366 );
buf ( n25368 , n25367 );
nor ( n25369 , n25360 , n25368 );
buf ( n25370 , n25369 );
buf ( n25371 , n25370 );
nand ( n25372 , n25343 , n25371 );
buf ( n25373 , n25372 );
buf ( n25374 , n25373 );
nor ( n25375 , n25302 , n25374 );
buf ( n25376 , n25375 );
buf ( n25377 , n25376 );
not ( n25378 , n25377 );
or ( n25379 , n25085 , n25378 );
buf ( n25380 , n25376 );
buf ( n25381 , n25083 );
or ( n25382 , n25380 , n25381 );
nand ( n25383 , n25379 , n25382 );
buf ( n25384 , n25383 );
buf ( n25385 , n25384 );
not ( n25386 , n25385 );
nand ( n25387 , n18207 , n25057 );
not ( n25388 , n25387 );
nand ( n25389 , n25052 , n25388 );
nor ( n25390 , n25386 , n25389 );
not ( n25391 , n19200 );
not ( n25392 , n19143 );
or ( n25393 , n25391 , n25392 );
not ( n25394 , n25051 );
nand ( n25395 , n25048 , n25394 );
nand ( n25396 , n25393 , n25395 );
buf ( n25397 , n25396 );
nand ( n25398 , n25397 , n275562 );
not ( n25399 , n25061 );
nor ( n25400 , n18206 , n25057 );
nand ( n25401 , n25399 , n25400 );
not ( n25402 , n25401 );
buf ( n25403 , n25065 );
buf ( n25404 , n25403 );
buf ( n25405 , n18705 );
buf ( n25406 , n25405 );
nand ( n25407 , n25404 , n25406 );
buf ( n25408 , n25407 );
buf ( n25409 , n25408 );
not ( n25410 , n25409 );
buf ( n25411 , n25403 );
buf ( n25412 , n25405 );
nor ( n25413 , n25411 , n25412 );
buf ( n25414 , n25413 );
buf ( n25415 , n25414 );
nor ( n25416 , n25410 , n25415 );
buf ( n25417 , n25416 );
buf ( n25418 , n25417 );
not ( n25419 , n25418 );
buf ( n25420 , n25087 );
buf ( n25421 , n25420 );
buf ( n25422 , n18747 );
buf ( n25423 , n25422 );
nor ( n25424 , n25421 , n25423 );
buf ( n25425 , n25424 );
buf ( n25426 , n25425 );
buf ( n25427 , n25096 );
buf ( n25428 , n25427 );
buf ( n25429 , n18763 );
buf ( n25430 , n25429 );
nor ( n25431 , n25428 , n25430 );
buf ( n25432 , n25431 );
buf ( n25433 , n25432 );
nor ( n25434 , n25426 , n25433 );
buf ( n25435 , n25434 );
buf ( n25436 , n25435 );
buf ( n25437 , n25109 );
buf ( n25438 , n25437 );
buf ( n25439 , n18405 );
buf ( n25440 , n25439 );
or ( n25441 , n25438 , n25440 );
buf ( n25442 , n25441 );
buf ( n25443 , n25442 );
not ( n25444 , n25443 );
buf ( n25445 , n25118 );
buf ( n25446 , n25445 );
buf ( n25447 , n18339 );
buf ( n25448 , n25447 );
nor ( n25449 , n25446 , n25448 );
buf ( n25450 , n25449 );
buf ( n25451 , n25450 );
nor ( n25452 , n25444 , n25451 );
buf ( n25453 , n25452 );
buf ( n25454 , n25453 );
and ( n25455 , n25436 , n25454 );
buf ( n25456 , n25455 );
buf ( n25457 , n25456 );
not ( n25458 , n25141 );
not ( n25459 , n25458 );
buf ( n25460 , n25459 );
buf ( n25461 , n25460 );
buf ( n25462 , n18912 );
buf ( n25463 , n25462 );
nor ( n25464 , n25461 , n25463 );
buf ( n25465 , n25464 );
buf ( n25466 , n25465 );
buf ( n25467 , n25133 );
buf ( n25468 , n25467 );
buf ( n25469 , n18882 );
buf ( n25470 , n25469 );
nor ( n25471 , n25468 , n25470 );
buf ( n25472 , n25471 );
buf ( n25473 , n25472 );
nor ( n25474 , n25466 , n25473 );
buf ( n25475 , n25474 );
buf ( n25476 , n25475 );
not ( n25477 , n25476 );
not ( n25478 , n25154 );
buf ( n25479 , n25478 );
buf ( n25480 , n25479 );
buf ( n25481 , n18387 );
buf ( n25482 , n25481 );
nor ( n25483 , n25480 , n25482 );
buf ( n25484 , n25483 );
buf ( n25485 , n25484 );
buf ( n25486 , n25163 );
buf ( n25487 , n25486 );
buf ( n25488 , n18364 );
buf ( n25489 , n25488 );
nor ( n25490 , n25487 , n25489 );
buf ( n25491 , n25490 );
buf ( n25492 , n25491 );
nor ( n25493 , n25485 , n25492 );
buf ( n25494 , n25493 );
buf ( n25495 , n25494 );
buf ( n25496 , n18071 );
buf ( n25497 , n25496 );
buf ( n25498 , n18870 );
buf ( n25499 , n25498 );
nor ( n25500 , n25497 , n25499 );
buf ( n25501 , n25500 );
buf ( n25502 , n25501 );
buf ( n25503 , n18289 );
buf ( n25504 , n18132 );
and ( n25505 , n25503 , n25504 );
buf ( n25506 , n25505 );
buf ( n25507 , n25506 );
buf ( n25508 , n19077 );
xor ( n25509 , n25507 , n25508 );
buf ( n25510 , n18131 );
and ( n25511 , n25509 , n25510 );
and ( n25512 , n25507 , n25508 );
or ( n25513 , n25511 , n25512 );
buf ( n25514 , n25513 );
buf ( n25515 , n25514 );
buf ( n25516 , n18319 );
buf ( n25517 , n25516 );
buf ( n25518 , n18115 );
buf ( n25519 , n25518 );
or ( n25520 , n25517 , n25519 );
buf ( n25521 , n25520 );
buf ( n25522 , n25521 );
nand ( n25523 , n25515 , n25522 );
buf ( n25524 , n25523 );
buf ( n25525 , n25524 );
or ( n25526 , n25502 , n25525 );
buf ( n25527 , n25501 );
buf ( n25528 , n25518 );
buf ( n25529 , n25516 );
nand ( n25530 , n25528 , n25529 );
buf ( n25531 , n25530 );
buf ( n25532 , n25531 );
or ( n25533 , n25527 , n25532 );
buf ( n25534 , n25496 );
buf ( n25535 , n25498 );
nand ( n25536 , n25534 , n25535 );
buf ( n25537 , n25536 );
buf ( n25538 , n25537 );
nand ( n25539 , n25526 , n25533 , n25538 );
buf ( n25540 , n25539 );
buf ( n25541 , n25540 );
nand ( n25542 , n25495 , n25541 );
buf ( n25543 , n25542 );
buf ( n25544 , n25543 );
not ( n25545 , n25544 );
buf ( n25546 , n25545 );
buf ( n25547 , n25546 );
not ( n25548 , n25547 );
or ( n25549 , n25477 , n25548 );
buf ( n25550 , n25484 );
buf ( n25551 , n25486 );
buf ( n25552 , n25488 );
nand ( n25553 , n25551 , n25552 );
buf ( n25554 , n25553 );
buf ( n25555 , n25554 );
or ( n25556 , n25550 , n25555 );
buf ( n25557 , n25479 );
buf ( n25558 , n25481 );
nand ( n25559 , n25557 , n25558 );
buf ( n25560 , n25559 );
buf ( n25561 , n25560 );
nand ( n25562 , n25556 , n25561 );
buf ( n25563 , n25562 );
buf ( n25564 , n25563 );
buf ( n25565 , n25475 );
and ( n25566 , n25564 , n25565 );
buf ( n25567 , n25472 );
buf ( n25568 , n25460 );
buf ( n25569 , n25462 );
nand ( n25570 , n25568 , n25569 );
buf ( n25571 , n25570 );
buf ( n25572 , n25571 );
or ( n25573 , n25567 , n25572 );
buf ( n25574 , n25467 );
buf ( n25575 , n25469 );
nand ( n25576 , n25574 , n25575 );
buf ( n25577 , n25576 );
buf ( n25578 , n25577 );
nand ( n25579 , n25573 , n25578 );
buf ( n25580 , n25579 );
buf ( n25581 , n25580 );
nor ( n25582 , n25566 , n25581 );
buf ( n25583 , n25582 );
buf ( n25584 , n25583 );
nand ( n25585 , n25549 , n25584 );
buf ( n25586 , n25585 );
buf ( n25587 , n25586 );
not ( n25588 , n25266 );
not ( n25589 , n25588 );
buf ( n25590 , n25589 );
buf ( n25591 , n25590 );
buf ( n25592 , n18982 );
buf ( n25593 , n25592 );
nor ( n25594 , n25591 , n25593 );
buf ( n25595 , n25594 );
buf ( n25596 , n25595 );
buf ( n25597 , n25275 );
buf ( n25598 , n25597 );
buf ( n25599 , n25598 );
buf ( n25600 , n19005 );
buf ( n25601 , n25600 );
nor ( n25602 , n25599 , n25601 );
buf ( n25603 , n25602 );
buf ( n25604 , n25603 );
nor ( n25605 , n25596 , n25604 );
buf ( n25606 , n25605 );
buf ( n25607 , n25606 );
not ( n25608 , n25287 );
not ( n25609 , n25608 );
buf ( n25610 , n25609 );
buf ( n25611 , n25610 );
buf ( n25612 , n18726 );
buf ( n25613 , n25612 );
nor ( n25614 , n25611 , n25613 );
buf ( n25615 , n25614 );
buf ( n25616 , n25615 );
not ( n25617 , n25616 );
buf ( n25618 , n25617 );
buf ( n25619 , n25618 );
and ( n25620 , n25607 , n25619 );
buf ( n25621 , n25620 );
buf ( n25622 , n25621 );
and ( n25623 , n25457 , n25587 , n25622 );
buf ( n25624 , n25621 );
not ( n25625 , n25624 );
buf ( n25626 , n25445 );
buf ( n25627 , n25447 );
nand ( n25628 , n25626 , n25627 );
buf ( n25629 , n25628 );
buf ( n25630 , n25629 );
not ( n25631 , n25630 );
buf ( n25632 , n25442 );
nand ( n25633 , n25631 , n25632 );
buf ( n25634 , n25633 );
buf ( n25635 , n25634 );
buf ( n25636 , n25437 );
buf ( n25637 , n25439 );
nand ( n25638 , n25636 , n25637 );
buf ( n25639 , n25638 );
buf ( n25640 , n25639 );
nand ( n25641 , n25635 , n25640 );
buf ( n25642 , n25641 );
buf ( n25643 , n25642 );
not ( n25644 , n25643 );
buf ( n25645 , n25435 );
not ( n25646 , n25645 );
or ( n25647 , n25644 , n25646 );
buf ( n25648 , n25425 );
not ( n25649 , n25648 );
buf ( n25650 , n25427 );
buf ( n25651 , n25429 );
nand ( n25652 , n25650 , n25651 );
buf ( n25653 , n25652 );
buf ( n25654 , n25653 );
not ( n25655 , n25654 );
and ( n25656 , n25649 , n25655 );
buf ( n25657 , n25420 );
buf ( n25658 , n25422 );
and ( n25659 , n25657 , n25658 );
buf ( n25660 , n25659 );
buf ( n25661 , n25660 );
nor ( n25662 , n25656 , n25661 );
buf ( n25663 , n25662 );
buf ( n25664 , n25663 );
nand ( n25665 , n25647 , n25664 );
buf ( n25666 , n25665 );
buf ( n25667 , n25666 );
not ( n25668 , n25667 );
or ( n25669 , n25625 , n25668 );
buf ( n25670 , n25595 );
buf ( n25671 , n25598 );
buf ( n25672 , n25600 );
nand ( n25673 , n25671 , n25672 );
buf ( n25674 , n25673 );
buf ( n25675 , n25674 );
or ( n25676 , n25670 , n25675 );
buf ( n25677 , n25590 );
buf ( n25678 , n25592 );
nand ( n25679 , n25677 , n25678 );
buf ( n25680 , n25679 );
buf ( n25681 , n25680 );
nand ( n25682 , n25676 , n25681 );
buf ( n25683 , n25682 );
buf ( n25684 , n25683 );
buf ( n25685 , n25618 );
and ( n25686 , n25684 , n25685 );
buf ( n25687 , n25610 );
buf ( n25688 , n25612 );
nand ( n25689 , n25687 , n25688 );
buf ( n25690 , n25689 );
buf ( n25691 , n25690 );
not ( n25692 , n25691 );
buf ( n25693 , n25692 );
buf ( n25694 , n25693 );
nor ( n25695 , n25686 , n25694 );
buf ( n25696 , n25695 );
buf ( n25697 , n25696 );
nand ( n25698 , n25669 , n25697 );
buf ( n25699 , n25698 );
buf ( n25700 , n25699 );
nor ( n25701 , n25623 , n25700 );
buf ( n25702 , n25701 );
buf ( n25703 , n25702 );
not ( n25704 , n25703 );
or ( n25705 , n25419 , n25704 );
buf ( n25706 , n25702 );
buf ( n25707 , n25417 );
or ( n25708 , n25706 , n25707 );
nand ( n25709 , n25705 , n25708 );
buf ( n25710 , n25709 );
buf ( n25711 , n25710 );
and ( n25712 , n25402 , n25711 );
not ( n25713 , n18696 );
nor ( n25714 , n19639 , n25713 );
nor ( n25715 , n25712 , n25714 );
or ( n25716 , n25061 , n25387 );
not ( n25717 , n25716 );
not ( n25718 , n25066 );
buf ( n25719 , n25718 );
buf ( n25720 , n25719 );
buf ( n25721 , n18701 );
buf ( n25722 , n25721 );
nand ( n25723 , n25720 , n25722 );
buf ( n25724 , n25723 );
buf ( n25725 , n25724 );
not ( n25726 , n25725 );
buf ( n25727 , n25719 );
buf ( n25728 , n25721 );
nor ( n25729 , n25727 , n25728 );
buf ( n25730 , n25729 );
buf ( n25731 , n25730 );
nor ( n25732 , n25726 , n25731 );
buf ( n25733 , n25732 );
buf ( n25734 , n25733 );
not ( n25735 , n25734 );
buf ( n25736 , n25086 );
buf ( n25737 , n25736 );
buf ( n25738 , n18744 );
buf ( n25739 , n25738 );
or ( n25740 , n25737 , n25739 );
buf ( n25741 , n25740 );
buf ( n25742 , n25741 );
buf ( n25743 , n18760 );
buf ( n25744 , n25743 );
buf ( n25745 , n25095 );
buf ( n25746 , n25745 );
or ( n25747 , n25744 , n25746 );
buf ( n25748 , n25747 );
buf ( n25749 , n25748 );
and ( n25750 , n25742 , n25749 );
buf ( n25751 , n25750 );
buf ( n25752 , n25751 );
buf ( n25753 , n25108 );
buf ( n25754 , n25753 );
buf ( n25755 , n25754 );
buf ( n25756 , n18402 );
buf ( n25757 , n25756 );
or ( n25758 , n25755 , n25757 );
buf ( n25759 , n25758 );
buf ( n25760 , n25759 );
not ( n25761 , n25760 );
buf ( n25762 , n25119 );
buf ( n25763 , n25762 );
buf ( n25764 , n18335 );
buf ( n25765 , n25764 );
nor ( n25766 , n25763 , n25765 );
buf ( n25767 , n25766 );
buf ( n25768 , n25767 );
nor ( n25769 , n25761 , n25768 );
buf ( n25770 , n25769 );
buf ( n25771 , n25770 );
and ( n25772 , n25752 , n25771 );
buf ( n25773 , n25772 );
buf ( n25774 , n25773 );
buf ( n25775 , n25142 );
buf ( n25776 , n25775 );
buf ( n25777 , n18908 );
buf ( n25778 , n25777 );
nor ( n25779 , n25776 , n25778 );
buf ( n25780 , n25779 );
buf ( n25781 , n25780 );
not ( n25782 , n25133 );
not ( n25783 , n25782 );
buf ( n25784 , n25783 );
buf ( n25785 , n25784 );
buf ( n25786 , n18878 );
buf ( n25787 , n25786 );
nor ( n25788 , n25785 , n25787 );
buf ( n25789 , n25788 );
buf ( n25790 , n25789 );
nor ( n25791 , n25781 , n25790 );
buf ( n25792 , n25791 );
buf ( n25793 , n25792 );
not ( n25794 , n25793 );
buf ( n25795 , n25478 );
buf ( n25796 , n25795 );
buf ( n25797 , n18383 );
buf ( n25798 , n25797 );
nor ( n25799 , n25796 , n25798 );
buf ( n25800 , n25799 );
buf ( n25801 , n25800 );
buf ( n25802 , n25163 );
buf ( n25803 , n25802 );
buf ( n25804 , n18356 );
buf ( n25805 , n25804 );
nor ( n25806 , n25803 , n25805 );
buf ( n25807 , n25806 );
buf ( n25808 , n25807 );
nor ( n25809 , n25801 , n25808 );
buf ( n25810 , n25809 );
buf ( n25811 , n25810 );
buf ( n25812 , n18071 );
buf ( n25813 , n25812 );
buf ( n25814 , n18866 );
buf ( n25815 , n25814 );
nor ( n25816 , n25813 , n25815 );
buf ( n25817 , n25816 );
buf ( n25818 , n25817 );
buf ( n25819 , n18306 );
buf ( n25820 , n18132 );
and ( n25821 , n25819 , n25820 );
buf ( n25822 , n25821 );
buf ( n25823 , n25822 );
buf ( n25824 , n19083 );
xor ( n25825 , n25823 , n25824 );
buf ( n25826 , n18131 );
and ( n25827 , n25825 , n25826 );
and ( n25828 , n25823 , n25824 );
or ( n25829 , n25827 , n25828 );
buf ( n25830 , n25829 );
buf ( n25831 , n25830 );
buf ( n25832 , n18115 );
buf ( n25833 , n25832 );
buf ( n25834 , n18327 );
buf ( n25835 , n25834 );
or ( n25836 , n25833 , n25835 );
buf ( n25837 , n25836 );
buf ( n25838 , n25837 );
nand ( n25839 , n25831 , n25838 );
buf ( n25840 , n25839 );
buf ( n25841 , n25840 );
or ( n25842 , n25818 , n25841 );
buf ( n25843 , n25817 );
buf ( n25844 , n25832 );
buf ( n25845 , n25834 );
nand ( n25846 , n25844 , n25845 );
buf ( n25847 , n25846 );
buf ( n25848 , n25847 );
or ( n25849 , n25843 , n25848 );
buf ( n25850 , n25812 );
buf ( n25851 , n25814 );
nand ( n25852 , n25850 , n25851 );
buf ( n25853 , n25852 );
buf ( n25854 , n25853 );
nand ( n25855 , n25842 , n25849 , n25854 );
buf ( n25856 , n25855 );
buf ( n25857 , n25856 );
nand ( n25858 , n25811 , n25857 );
buf ( n25859 , n25858 );
buf ( n25860 , n25859 );
not ( n25861 , n25860 );
buf ( n25862 , n25861 );
buf ( n25863 , n25862 );
not ( n25864 , n25863 );
or ( n25865 , n25794 , n25864 );
buf ( n25866 , n25800 );
buf ( n25867 , n25802 );
buf ( n25868 , n25804 );
nand ( n25869 , n25867 , n25868 );
buf ( n25870 , n25869 );
buf ( n25871 , n25870 );
or ( n25872 , n25866 , n25871 );
buf ( n25873 , n25795 );
buf ( n25874 , n25797 );
nand ( n25875 , n25873 , n25874 );
buf ( n25876 , n25875 );
buf ( n25877 , n25876 );
nand ( n25878 , n25872 , n25877 );
buf ( n25879 , n25878 );
buf ( n25880 , n25879 );
buf ( n25881 , n25792 );
and ( n25882 , n25880 , n25881 );
buf ( n25883 , n25789 );
buf ( n25884 , n25775 );
buf ( n25885 , n25777 );
nand ( n25886 , n25884 , n25885 );
buf ( n25887 , n25886 );
buf ( n25888 , n25887 );
or ( n25889 , n25883 , n25888 );
buf ( n25890 , n25784 );
buf ( n25891 , n25786 );
nand ( n25892 , n25890 , n25891 );
buf ( n25893 , n25892 );
buf ( n25894 , n25893 );
nand ( n25895 , n25889 , n25894 );
buf ( n25896 , n25895 );
buf ( n25897 , n25896 );
nor ( n25898 , n25882 , n25897 );
buf ( n25899 , n25898 );
buf ( n25900 , n25899 );
nand ( n25901 , n25865 , n25900 );
buf ( n25902 , n25901 );
buf ( n25903 , n25902 );
not ( n25904 , n25588 );
buf ( n25905 , n25904 );
buf ( n25906 , n25905 );
buf ( n25907 , n18987 );
buf ( n25908 , n25907 );
nor ( n25909 , n25906 , n25908 );
buf ( n25910 , n25909 );
buf ( n25911 , n25910 );
buf ( n25912 , n25597 );
buf ( n25913 , n25912 );
buf ( n25914 , n19010 );
buf ( n25915 , n25914 );
nor ( n25916 , n25913 , n25915 );
buf ( n25917 , n25916 );
buf ( n25918 , n25917 );
nor ( n25919 , n25911 , n25918 );
buf ( n25920 , n25919 );
buf ( n25921 , n25920 );
not ( n25922 , n25608 );
buf ( n25923 , n25922 );
buf ( n25924 , n25923 );
buf ( n25925 , n18731 );
buf ( n25926 , n25925 );
nor ( n25927 , n25924 , n25926 );
buf ( n25928 , n25927 );
buf ( n25929 , n25928 );
not ( n25930 , n25929 );
buf ( n25931 , n25930 );
buf ( n25932 , n25931 );
and ( n25933 , n25921 , n25932 );
buf ( n25934 , n25933 );
buf ( n25935 , n25934 );
and ( n25936 , n25774 , n25903 , n25935 );
buf ( n25937 , n25934 );
not ( n25938 , n25937 );
buf ( n25939 , n25751 );
buf ( n25940 , n25762 );
buf ( n25941 , n25764 );
nand ( n25942 , n25940 , n25941 );
buf ( n25943 , n25942 );
buf ( n25944 , n25943 );
not ( n25945 , n25944 );
buf ( n25946 , n25759 );
nand ( n25947 , n25945 , n25946 );
buf ( n25948 , n25947 );
buf ( n25949 , n25948 );
buf ( n25950 , n25754 );
buf ( n25951 , n25756 );
nand ( n25952 , n25950 , n25951 );
buf ( n25953 , n25952 );
buf ( n25954 , n25953 );
nand ( n25955 , n25949 , n25954 );
buf ( n25956 , n25955 );
buf ( n25957 , n25956 );
nand ( n25958 , n25939 , n25957 );
buf ( n25959 , n25958 );
buf ( n25960 , n25959 );
buf ( n25961 , n25745 );
buf ( n25962 , n25743 );
nand ( n25963 , n25961 , n25962 );
buf ( n25964 , n25963 );
buf ( n25965 , n25964 );
not ( n25966 , n25965 );
buf ( n25967 , n25741 );
nand ( n25968 , n25966 , n25967 );
buf ( n25969 , n25968 );
buf ( n25970 , n25969 );
buf ( n25971 , n25736 );
buf ( n25972 , n25738 );
nand ( n25973 , n25971 , n25972 );
buf ( n25974 , n25973 );
buf ( n25975 , n25974 );
nand ( n25976 , n25960 , n25970 , n25975 );
buf ( n25977 , n25976 );
buf ( n25978 , n25977 );
not ( n25979 , n25978 );
or ( n25980 , n25938 , n25979 );
buf ( n25981 , n25910 );
buf ( n25982 , n25912 );
buf ( n25983 , n25914 );
nand ( n25984 , n25982 , n25983 );
buf ( n25985 , n25984 );
buf ( n25986 , n25985 );
or ( n25987 , n25981 , n25986 );
buf ( n25988 , n25905 );
buf ( n25989 , n25907 );
nand ( n25990 , n25988 , n25989 );
buf ( n25991 , n25990 );
buf ( n25992 , n25991 );
nand ( n25993 , n25987 , n25992 );
buf ( n25994 , n25993 );
buf ( n25995 , n25994 );
buf ( n25996 , n25931 );
and ( n25997 , n25995 , n25996 );
buf ( n25998 , n25923 );
buf ( n25999 , n25925 );
nand ( n26000 , n25998 , n25999 );
buf ( n26001 , n26000 );
buf ( n26002 , n26001 );
not ( n26003 , n26002 );
buf ( n26004 , n26003 );
buf ( n26005 , n26004 );
nor ( n26006 , n25997 , n26005 );
buf ( n26007 , n26006 );
buf ( n26008 , n26007 );
nand ( n26009 , n25980 , n26008 );
buf ( n26010 , n26009 );
buf ( n26011 , n26010 );
nor ( n26012 , n25936 , n26011 );
buf ( n26013 , n26012 );
buf ( n26014 , n26013 );
not ( n26015 , n26014 );
or ( n26016 , n25735 , n26015 );
buf ( n26017 , n26013 );
buf ( n26018 , n25733 );
or ( n26019 , n26017 , n26018 );
nand ( n26020 , n26016 , n26019 );
buf ( n26021 , n26020 );
buf ( n26022 , n26021 );
nand ( n26023 , n25717 , n26022 );
nand ( n26024 , n25398 , n25715 , n26023 );
nor ( n26025 , n25390 , n26024 );
nand ( n26026 , n25052 , n25400 );
not ( n26027 , n26026 );
buf ( n26028 , n25067 );
buf ( n26029 , n26028 );
buf ( n26030 , n18705 );
buf ( n26031 , n26030 );
nand ( n26032 , n26029 , n26031 );
buf ( n26033 , n26032 );
buf ( n26034 , n26033 );
not ( n26035 , n26034 );
buf ( n26036 , n26028 );
buf ( n26037 , n26030 );
nor ( n26038 , n26036 , n26037 );
buf ( n26039 , n26038 );
buf ( n26040 , n26039 );
nor ( n26041 , n26035 , n26040 );
buf ( n26042 , n26041 );
buf ( n26043 , n26042 );
not ( n26044 , n26043 );
buf ( n26045 , n25096 );
buf ( n26046 , n26045 );
buf ( n26047 , n18763 );
buf ( n26048 , n26047 );
or ( n26049 , n26046 , n26048 );
buf ( n26050 , n26049 );
buf ( n26051 , n26050 );
not ( n26052 , n26051 );
buf ( n26053 , n25086 );
buf ( n26054 , n26053 );
buf ( n26055 , n18747 );
buf ( n26056 , n26055 );
nor ( n26057 , n26054 , n26056 );
buf ( n26058 , n26057 );
buf ( n26059 , n26058 );
nor ( n26060 , n26052 , n26059 );
buf ( n26061 , n26060 );
buf ( n26062 , n26061 );
buf ( n26063 , n25753 );
buf ( n26064 , n26063 );
buf ( n26065 , n18405 );
buf ( n26066 , n26065 );
nor ( n26067 , n26064 , n26066 );
buf ( n26068 , n26067 );
buf ( n26069 , n26068 );
buf ( n26070 , n25119 );
buf ( n26071 , n26070 );
buf ( n26072 , n18339 );
buf ( n26073 , n26072 );
nor ( n26074 , n26071 , n26073 );
buf ( n26075 , n26074 );
buf ( n26076 , n26075 );
nor ( n26077 , n26069 , n26076 );
buf ( n26078 , n26077 );
buf ( n26079 , n26078 );
and ( n26080 , n26062 , n26079 );
buf ( n26081 , n26080 );
buf ( n26082 , n26081 );
not ( n26083 , n25782 );
buf ( n26084 , n26083 );
buf ( n26085 , n26084 );
buf ( n26086 , n18882 );
buf ( n26087 , n26086 );
nor ( n26088 , n26085 , n26087 );
buf ( n26089 , n26088 );
buf ( n26090 , n26089 );
not ( n26091 , n25458 );
buf ( n26092 , n26091 );
buf ( n26093 , n26092 );
buf ( n26094 , n18912 );
buf ( n26095 , n26094 );
nor ( n26096 , n26093 , n26095 );
buf ( n26097 , n26096 );
buf ( n26098 , n26097 );
nor ( n26099 , n26090 , n26098 );
buf ( n26100 , n26099 );
buf ( n26101 , n26100 );
not ( n26102 , n26101 );
not ( n26103 , n25154 );
buf ( n26104 , n26103 );
buf ( n26105 , n26104 );
buf ( n26106 , n18387 );
buf ( n26107 , n26106 );
nor ( n26108 , n26105 , n26107 );
buf ( n26109 , n26108 );
buf ( n26110 , n26109 );
buf ( n26111 , n25164 );
buf ( n26112 , n26111 );
buf ( n26113 , n18364 );
buf ( n26114 , n26113 );
nor ( n26115 , n26112 , n26114 );
buf ( n26116 , n26115 );
buf ( n26117 , n26116 );
nor ( n26118 , n26110 , n26117 );
buf ( n26119 , n26118 );
buf ( n26120 , n26119 );
buf ( n26121 , n18071 );
buf ( n26122 , n26121 );
buf ( n26123 , n18870 );
buf ( n26124 , n26123 );
nor ( n26125 , n26122 , n26124 );
buf ( n26126 , n26125 );
buf ( n26127 , n26126 );
buf ( n26128 , n18289 );
buf ( n26129 , n18134 );
buf ( n26130 , n26129 );
and ( n26131 , n26128 , n26130 );
buf ( n26132 , n26131 );
buf ( n26133 , n26132 );
buf ( n26134 , n19077 );
xor ( n26135 , n26133 , n26134 );
buf ( n26136 , n18131 );
and ( n26137 , n26135 , n26136 );
and ( n26138 , n26133 , n26134 );
or ( n26139 , n26137 , n26138 );
buf ( n26140 , n26139 );
buf ( n26141 , n26140 );
buf ( n26142 , n18115 );
buf ( n26143 , n26142 );
buf ( n26144 , n18319 );
buf ( n26145 , n26144 );
or ( n26146 , n26143 , n26145 );
buf ( n26147 , n26146 );
buf ( n26148 , n26147 );
nand ( n26149 , n26141 , n26148 );
buf ( n26150 , n26149 );
buf ( n26151 , n26150 );
or ( n26152 , n26127 , n26151 );
buf ( n26153 , n26126 );
buf ( n26154 , n26142 );
buf ( n26155 , n26144 );
nand ( n26156 , n26154 , n26155 );
buf ( n26157 , n26156 );
buf ( n26158 , n26157 );
or ( n26159 , n26153 , n26158 );
buf ( n26160 , n26121 );
buf ( n26161 , n26123 );
nand ( n26162 , n26160 , n26161 );
buf ( n26163 , n26162 );
buf ( n26164 , n26163 );
nand ( n26165 , n26152 , n26159 , n26164 );
buf ( n26166 , n26165 );
buf ( n26167 , n26166 );
nand ( n26168 , n26120 , n26167 );
buf ( n26169 , n26168 );
buf ( n26170 , n26169 );
not ( n26171 , n26170 );
buf ( n26172 , n26171 );
buf ( n26173 , n26172 );
not ( n26174 , n26173 );
or ( n26175 , n26102 , n26174 );
buf ( n26176 , n26109 );
buf ( n26177 , n26111 );
buf ( n26178 , n26113 );
nand ( n26179 , n26177 , n26178 );
buf ( n26180 , n26179 );
buf ( n26181 , n26180 );
or ( n26182 , n26176 , n26181 );
buf ( n26183 , n26104 );
buf ( n26184 , n26106 );
nand ( n26185 , n26183 , n26184 );
buf ( n26186 , n26185 );
buf ( n26187 , n26186 );
nand ( n26188 , n26182 , n26187 );
buf ( n26189 , n26188 );
buf ( n26190 , n26189 );
buf ( n26191 , n26100 );
and ( n26192 , n26190 , n26191 );
buf ( n26193 , n26089 );
buf ( n26194 , n26092 );
buf ( n26195 , n26094 );
nand ( n26196 , n26194 , n26195 );
buf ( n26197 , n26196 );
buf ( n26198 , n26197 );
or ( n26199 , n26193 , n26198 );
buf ( n26200 , n26084 );
buf ( n26201 , n26086 );
nand ( n26202 , n26200 , n26201 );
buf ( n26203 , n26202 );
buf ( n26204 , n26203 );
nand ( n26205 , n26199 , n26204 );
buf ( n26206 , n26205 );
buf ( n26207 , n26206 );
nor ( n26208 , n26192 , n26207 );
buf ( n26209 , n26208 );
buf ( n26210 , n26209 );
nand ( n26211 , n26175 , n26210 );
buf ( n26212 , n26211 );
buf ( n26213 , n26212 );
buf ( n26214 , n25267 );
buf ( n26215 , n26214 );
buf ( n26216 , n18982 );
buf ( n26217 , n26216 );
nor ( n26218 , n26215 , n26217 );
buf ( n26219 , n26218 );
buf ( n26220 , n26219 );
buf ( n26221 , n25276 );
buf ( n26222 , n26221 );
buf ( n26223 , n19005 );
buf ( n26224 , n26223 );
nor ( n26225 , n26222 , n26224 );
buf ( n26226 , n26225 );
buf ( n26227 , n26226 );
nor ( n26228 , n26220 , n26227 );
buf ( n26229 , n26228 );
buf ( n26230 , n26229 );
not ( n26231 , n25288 );
not ( n26232 , n26231 );
buf ( n26233 , n26232 );
buf ( n26234 , n26233 );
buf ( n26235 , n18726 );
buf ( n26236 , n26235 );
nor ( n26237 , n26234 , n26236 );
buf ( n26238 , n26237 );
buf ( n26239 , n26238 );
not ( n26240 , n26239 );
buf ( n26241 , n26240 );
buf ( n26242 , n26241 );
and ( n26243 , n26230 , n26242 );
buf ( n26244 , n26243 );
buf ( n26245 , n26244 );
and ( n26246 , n26082 , n26213 , n26245 );
buf ( n26247 , n26244 );
not ( n26248 , n26247 );
buf ( n26249 , n26058 );
buf ( n26250 , n26045 );
buf ( n26251 , n26047 );
nand ( n26252 , n26250 , n26251 );
buf ( n26253 , n26252 );
buf ( n26254 , n26253 );
or ( n26255 , n26249 , n26254 );
buf ( n26256 , n26061 );
buf ( n26257 , n26068 );
buf ( n26258 , n26070 );
buf ( n26259 , n26072 );
nand ( n26260 , n26258 , n26259 );
buf ( n26261 , n26260 );
buf ( n26262 , n26261 );
or ( n26263 , n26257 , n26262 );
buf ( n26264 , n26063 );
buf ( n26265 , n26065 );
nand ( n26266 , n26264 , n26265 );
buf ( n26267 , n26266 );
buf ( n26268 , n26267 );
nand ( n26269 , n26263 , n26268 );
buf ( n26270 , n26269 );
buf ( n26271 , n26270 );
nand ( n26272 , n26256 , n26271 );
buf ( n26273 , n26272 );
buf ( n26274 , n26273 );
buf ( n26275 , n26053 );
buf ( n26276 , n26055 );
nand ( n26277 , n26275 , n26276 );
buf ( n26278 , n26277 );
buf ( n26279 , n26278 );
nand ( n26280 , n26255 , n26274 , n26279 );
buf ( n26281 , n26280 );
buf ( n26282 , n26281 );
not ( n26283 , n26282 );
or ( n26284 , n26248 , n26283 );
buf ( n26285 , n26219 );
buf ( n26286 , n26221 );
buf ( n26287 , n26223 );
nand ( n26288 , n26286 , n26287 );
buf ( n26289 , n26288 );
buf ( n26290 , n26289 );
or ( n26291 , n26285 , n26290 );
buf ( n26292 , n26214 );
buf ( n26293 , n26216 );
nand ( n26294 , n26292 , n26293 );
buf ( n26295 , n26294 );
buf ( n26296 , n26295 );
nand ( n26297 , n26291 , n26296 );
buf ( n26298 , n26297 );
buf ( n26299 , n26298 );
buf ( n26300 , n26241 );
and ( n26301 , n26299 , n26300 );
buf ( n26302 , n26233 );
buf ( n26303 , n26235 );
nand ( n26304 , n26302 , n26303 );
buf ( n26305 , n26304 );
buf ( n26306 , n26305 );
not ( n26307 , n26306 );
buf ( n26308 , n26307 );
buf ( n26309 , n26308 );
nor ( n26310 , n26301 , n26309 );
buf ( n26311 , n26310 );
buf ( n26312 , n26311 );
nand ( n26313 , n26284 , n26312 );
buf ( n26314 , n26313 );
buf ( n26315 , n26314 );
nor ( n26316 , n26246 , n26315 );
buf ( n26317 , n26316 );
buf ( n26318 , n26317 );
not ( n26319 , n26318 );
or ( n26320 , n26044 , n26319 );
buf ( n26321 , n26317 );
buf ( n26322 , n26042 );
or ( n26323 , n26321 , n26322 );
nand ( n26324 , n26320 , n26323 );
buf ( n26325 , n26324 );
buf ( n26326 , n26325 );
nand ( n26327 , n26027 , n26326 );
nand ( n26328 , n25068 , n26025 , n26327 );
buf ( n26329 , n26328 );
buf ( n26330 , n26329 );
not ( n26331 , n275550 );
buf ( n26332 , n26331 );
buf ( n26333 , n26332 );
not ( n26334 , n275550 );
buf ( n26335 , n26334 );
buf ( n26336 , n26335 );
buf ( n26337 , n275554 );
or ( n26338 , n21657 , n14909 );
nand ( n26339 , n17411 , n21681 );
not ( n26340 , n17561 );
not ( n26341 , n14538 );
not ( n26342 , n26341 );
and ( n26343 , n26340 , n26342 );
and ( n26344 , n17405 , n21668 );
nor ( n26345 , n26343 , n26344 );
nand ( n26346 , n17502 , n21685 );
not ( n26347 , n20765 );
not ( n26348 , n14527 );
not ( n26349 , n26348 );
and ( n26350 , n26347 , n26349 );
and ( n26351 , n21678 , n16968 );
nor ( n26352 , n26350 , n26351 );
and ( n26353 , n26339 , n26345 , n26346 , n26352 );
nand ( n26354 , n26338 , n26353 );
buf ( n26355 , n26354 );
buf ( n26356 , n26355 );
nand ( n26357 , n14867 , n14858 , n14839 );
not ( n26358 , n26357 );
nand ( n26359 , n14906 , n14830 );
not ( n26360 , n26359 );
nand ( n26361 , n26360 , n14827 );
nor ( n26362 , n26361 , n14895 );
nand ( n26363 , n26358 , n26362 );
buf ( n26364 , n26363 );
buf ( n26365 , n26364 );
or ( n26366 , n20740 , n26365 );
nor ( n26367 , n16964 , n26357 );
not ( n26368 , n26367 );
buf ( n26369 , n26368 );
not ( n26370 , n26369 );
nand ( n26371 , n20813 , n26370 );
nor ( n26372 , n26357 , n22897 );
nand ( n26373 , n26372 , n17402 );
not ( n26374 , n26373 );
nand ( n26375 , n20762 , n26374 );
not ( n26376 , n17499 );
not ( n26377 , n26372 );
or ( n26378 , n26376 , n26377 );
not ( n26379 , n17544 );
nand ( n26380 , n26378 , n26379 );
not ( n26381 , n26358 );
not ( n26382 , n26361 );
nand ( n26383 , n26382 , n16956 );
nor ( n26384 , n26381 , n26383 );
nor ( n26385 , n26380 , n26384 );
not ( n26386 , n17542 );
nand ( n26387 , n26363 , n26386 );
nor ( n26388 , n26367 , n26387 );
nand ( n26389 , n26385 , n26388 , n26373 );
buf ( n26390 , n26389 );
nor ( n26391 , n26390 , n20770 );
not ( n26392 , n26384 );
not ( n26393 , n26392 );
nand ( n26394 , n20782 , n26393 );
buf ( n26395 , n26380 );
nand ( n26396 , n26395 , n20788 );
nand ( n26397 , n17542 , n13828 );
nand ( n26398 , n26394 , n26396 , n26397 );
nor ( n26399 , n26391 , n26398 );
and ( n26400 , n26371 , n26375 , n26399 );
nand ( n26401 , n26366 , n26400 );
buf ( n26402 , n26401 );
buf ( n26403 , n26402 );
not ( n26404 , n10832 );
not ( n26405 , n9157 );
or ( n26406 , n26404 , n26405 );
not ( n26407 , n10809 );
not ( n26408 , n26407 );
or ( n26409 , n9157 , n26408 );
nand ( n26410 , n26406 , n26409 );
buf ( n26411 , n26410 );
buf ( n26412 , n26411 );
buf ( n26413 , n275554 );
buf ( n26414 , n275554 );
buf ( n26415 , n275554 );
not ( n26416 , n11454 );
or ( n26417 , n26416 , n9158 );
not ( n26418 , n11432 );
or ( n26419 , n26418 , n9157 );
nand ( n26420 , n26417 , n26419 );
buf ( n26421 , n26420 );
buf ( n26422 , n26421 );
buf ( n26423 , n14292 );
and ( n26424 , n13373 , n26423 );
not ( n26425 , n13373 );
buf ( n26426 , n14251 );
not ( n26427 , n26426 );
nor ( n26428 , n20719 , n26427 );
buf ( n26429 , n26428 );
buf ( n26430 , n14154 );
and ( n26431 , n26429 , n26430 );
not ( n26432 , n26429 );
not ( n26433 , n26430 );
and ( n26434 , n26432 , n26433 );
nor ( n26435 , n26431 , n26434 );
buf ( n26436 , n26435 );
and ( n26437 , n26425 , n26436 );
nor ( n26438 , n26424 , n26437 );
not ( n26439 , n26438 );
not ( n26440 , n23789 );
and ( n26441 , n26439 , n26440 );
not ( n26442 , n16667 );
nand ( n26443 , n26442 , n16890 );
not ( n26444 , n26443 );
not ( n26445 , n16402 );
buf ( n26446 , n16659 );
nor ( n26447 , n26445 , n26446 );
not ( n26448 , n26447 );
not ( n26449 , n20875 );
or ( n26450 , n26448 , n26449 );
nand ( n26451 , n16902 , n16904 );
not ( n26452 , n26451 );
not ( n26453 , n26446 );
and ( n26454 , n26452 , n26453 );
not ( n26455 , n16888 );
nor ( n26456 , n26454 , n26455 );
nand ( n26457 , n26450 , n26456 );
not ( n26458 , n26457 );
or ( n26459 , n26444 , n26458 );
or ( n26460 , n26457 , n26443 );
nand ( n26461 , n26459 , n26460 );
buf ( n26462 , n26461 );
nand ( n26463 , n26462 , n20889 );
nand ( n26464 , n17108 , n17351 );
not ( n26465 , n26464 );
not ( n26466 , n17120 );
nor ( n26467 , n17229 , n26466 );
not ( n26468 , n26467 );
not ( n26469 , n20913 );
or ( n26470 , n26468 , n26469 );
and ( n26471 , n17333 , n20917 );
nand ( n26472 , n20916 , n26471 , n20891 );
nand ( n26473 , n17334 , n26472 );
not ( n26474 , n26473 );
not ( n26475 , n26466 );
and ( n26476 , n26474 , n26475 );
nor ( n26477 , n26476 , n17346 );
nand ( n26478 , n26470 , n26477 );
not ( n26479 , n26478 );
or ( n26480 , n26465 , n26479 );
or ( n26481 , n26478 , n26464 );
nand ( n26482 , n26480 , n26481 );
buf ( n26483 , n26482 );
nand ( n26484 , n26483 , n20927 );
not ( n26485 , n17448 );
not ( n26486 , n20930 );
not ( n26487 , n17446 );
and ( n26488 , n26486 , n26487 , n17455 );
not ( n26489 , n26488 );
or ( n26490 , n26485 , n26489 );
or ( n26491 , n26488 , n17448 );
nand ( n26492 , n26490 , n26491 );
buf ( n26493 , n26492 );
and ( n26494 , n26493 , n17409 );
buf ( n26495 , n17447 );
buf ( n26496 , n26495 );
buf ( n26497 , n26496 );
buf ( n26498 , n26497 );
and ( n26499 , n20940 , n26498 );
nor ( n26500 , n26494 , n26499 );
nand ( n26501 , n26463 , n26484 , n26500 );
nor ( n26502 , n26441 , n26501 );
or ( n26503 , n26502 , n20950 );
nand ( n26504 , n20950 , n13704 );
nand ( n26505 , n26503 , n26504 );
buf ( n26506 , n26505 );
buf ( n26507 , n26506 );
not ( n26508 , n275550 );
buf ( n26509 , n26508 );
buf ( n26510 , n26509 );
or ( n26511 , n24728 , n20950 );
nand ( n26512 , n20950 , n13596 );
nand ( n26513 , n26511 , n26512 );
buf ( n26514 , n26513 );
buf ( n26515 , n26514 );
buf ( n26516 , n21039 );
and ( n26517 , n26516 , n21760 );
not ( n26518 , n26516 );
buf ( n26519 , n21726 );
buf ( n26520 , n21734 );
buf ( n26521 , n18834 );
buf ( n26522 , n18684 );
nand ( n26523 , n26521 , n26522 );
buf ( n26524 , n26523 );
buf ( n26525 , n26524 );
not ( n26526 , n26525 );
buf ( n26527 , n26526 );
buf ( n26528 , n26527 );
buf ( n26529 , n18573 );
buf ( n26530 , n26529 );
nand ( n26531 , n26528 , n26530 );
buf ( n26532 , n26531 );
buf ( n26533 , n26532 );
nor ( n26534 , n26520 , n26533 );
buf ( n26535 , n26534 );
buf ( n26536 , n26535 );
nand ( n26537 , n26519 , n26536 );
buf ( n26538 , n26537 );
buf ( n26539 , n26538 );
buf ( n26540 , n18548 );
buf ( n26541 , n26540 );
not ( n26542 , n26541 );
buf ( n26543 , n26542 );
buf ( n26544 , n26543 );
and ( n26545 , n26539 , n26544 );
not ( n26546 , n26539 );
buf ( n26547 , n26540 );
and ( n26548 , n26546 , n26547 );
nor ( n26549 , n26545 , n26548 );
buf ( n26550 , n26549 );
buf ( n26551 , n26550 );
buf ( n26552 , n26551 );
buf ( n26553 , n26552 );
buf ( n26554 , n19069 );
not ( n26555 , n21138 );
not ( n26556 , n21117 );
nand ( n26557 , n26555 , n26556 );
buf ( n26558 , n21726 );
buf ( n26559 , n21734 );
buf ( n26560 , n26527 );
not ( n26561 , n26560 );
buf ( n26562 , n26561 );
buf ( n26563 , n26562 );
nor ( n26564 , n26559 , n26563 );
buf ( n26565 , n26564 );
buf ( n26566 , n26565 );
nand ( n26567 , n26558 , n26566 );
buf ( n26568 , n26567 );
buf ( n26569 , n26568 );
buf ( n26570 , n26529 );
not ( n26571 , n26570 );
buf ( n26572 , n26571 );
buf ( n26573 , n26572 );
and ( n26574 , n26569 , n26573 );
not ( n26575 , n26569 );
buf ( n26576 , n26529 );
and ( n26577 , n26575 , n26576 );
nor ( n26578 , n26574 , n26577 );
buf ( n26579 , n26578 );
buf ( n26580 , n26579 );
buf ( n26581 , n26580 );
nand ( n26582 , n19603 , n26581 );
nor ( n26583 , n26557 , n26582 );
buf ( n26584 , n21734 );
not ( n26585 , n26584 );
buf ( n26586 , n21726 );
nand ( n26587 , n26585 , n26586 );
buf ( n26588 , n26587 );
buf ( n26589 , n26588 );
buf ( n26590 , n21739 );
and ( n26591 , n26589 , n26590 );
not ( n26592 , n26589 );
buf ( n26593 , n21736 );
and ( n26594 , n26592 , n26593 );
nor ( n26595 , n26591 , n26594 );
buf ( n26596 , n26595 );
buf ( n26597 , n26596 );
buf ( n26598 , n26597 );
nand ( n26599 , n26598 , n23952 , n21115 );
nor ( n26600 , n23956 , n26599 );
nand ( n26601 , n26583 , n26600 );
not ( n26602 , n26601 );
buf ( n26603 , n21726 );
buf ( n26604 , n18978 );
not ( n26605 , n26604 );
buf ( n26606 , n26605 );
buf ( n26607 , n26606 );
buf ( n26608 , n23943 );
nor ( n26609 , n26607 , n26608 );
buf ( n26610 , n26609 );
buf ( n26611 , n26610 );
nand ( n26612 , n26603 , n26611 );
buf ( n26613 , n26612 );
buf ( n26614 , n26613 );
buf ( n26615 , n18605 );
buf ( n26616 , n26615 );
not ( n26617 , n26616 );
buf ( n26618 , n26617 );
buf ( n26619 , n26618 );
and ( n26620 , n26614 , n26619 );
not ( n26621 , n26614 );
buf ( n26622 , n26615 );
and ( n26623 , n26621 , n26622 );
nor ( n26624 , n26620 , n26623 );
buf ( n26625 , n26624 );
buf ( n26626 , n26625 );
buf ( n26627 , n26626 );
buf ( n26628 , n21758 );
nand ( n26629 , n23978 , n26627 , n26628 );
buf ( n26630 , n26629 );
not ( n26631 , n26630 );
and ( n26632 , n26554 , n26602 , n26631 );
xor ( n26633 , n26553 , n26632 );
buf ( n26634 , n26633 );
and ( n26635 , n26518 , n26634 );
nor ( n26636 , n26517 , n26635 );
not ( n26637 , n26636 );
buf ( n26638 , n20987 );
and ( n26639 , n26637 , n26638 );
not ( n26640 , n21001 );
not ( n26641 , n277603 );
buf ( n26642 , n22399 );
not ( n26643 , n26642 );
buf ( n26644 , n22671 );
nand ( n26645 , n26643 , n26644 );
buf ( n26646 , n26645 );
buf ( n26647 , n26646 );
not ( n26648 , n26647 );
buf ( n26649 , n22374 );
buf ( n26650 , n22392 );
and ( n26651 , n26649 , n26650 );
buf ( n26652 , n26651 );
buf ( n26653 , n26652 );
not ( n26654 , n26653 );
buf ( n26655 , n22593 );
not ( n26656 , n26655 );
or ( n26657 , n26654 , n26656 );
buf ( n26658 , n22642 );
buf ( n26659 , n22392 );
and ( n26660 , n26658 , n26659 );
buf ( n26661 , n22664 );
nor ( n26662 , n26660 , n26661 );
buf ( n26663 , n26662 );
buf ( n26664 , n26663 );
nand ( n26665 , n26657 , n26664 );
buf ( n26666 , n26665 );
buf ( n26667 , n26666 );
not ( n26668 , n26667 );
or ( n26669 , n26648 , n26668 );
buf ( n26670 , n26666 );
buf ( n26671 , n26646 );
or ( n26672 , n26670 , n26671 );
nand ( n26673 , n26669 , n26672 );
buf ( n26674 , n26673 );
buf ( n26675 , n26674 );
not ( n26676 , n26675 );
or ( n26677 , n26641 , n26676 );
nand ( n26678 , n277351 , n9692 );
nand ( n26679 , n26677 , n26678 );
and ( n26680 , n19242 , n26679 );
buf ( n26681 , n26680 );
not ( n26682 , n26681 );
buf ( n26683 , n18572 );
buf ( n26684 , n26683 );
not ( n26685 , n26684 );
or ( n26686 , n26682 , n26685 );
not ( n26687 , n26681 );
not ( n26688 , n26684 );
nand ( n26689 , n26687 , n26688 );
nand ( n26690 , n26686 , n26689 );
buf ( n26691 , n18833 );
buf ( n26692 , n26691 );
not ( n26693 , n277527 );
buf ( n26694 , n22374 );
buf ( n26695 , n22389 );
not ( n26696 , n26695 );
buf ( n26697 , n26696 );
buf ( n26698 , n26697 );
and ( n26699 , n26694 , n26698 );
buf ( n26700 , n26699 );
buf ( n26701 , n26700 );
not ( n26702 , n26701 );
buf ( n26703 , n22592 );
not ( n26704 , n26703 );
or ( n26705 , n26702 , n26704 );
buf ( n26706 , n22642 );
buf ( n26707 , n26697 );
and ( n26708 , n26706 , n26707 );
buf ( n26709 , n22649 );
nor ( n26710 , n26708 , n26709 );
buf ( n26711 , n26710 );
buf ( n26712 , n26711 );
nand ( n26713 , n26705 , n26712 );
buf ( n26714 , n26713 );
buf ( n26715 , n26714 );
buf ( n26716 , n22654 );
buf ( n26717 , n22661 );
nand ( n26718 , n26716 , n26717 );
buf ( n26719 , n26718 );
buf ( n26720 , n26719 );
xnor ( n26721 , n26715 , n26720 );
buf ( n26722 , n26721 );
buf ( n26723 , n26722 );
not ( n26724 , n26723 );
or ( n26725 , n26693 , n26724 );
nand ( n26726 , n277983 , n22376 );
nand ( n26727 , n26725 , n26726 );
nand ( n26728 , n19242 , n26727 );
not ( n26729 , n26728 );
buf ( n26730 , n26729 );
not ( n26731 , n26730 );
and ( n26732 , n26692 , n26731 );
or ( n26733 , n26690 , n26732 );
nand ( n26734 , n26690 , n26732 );
nand ( n26735 , n26733 , n26734 );
not ( n26736 , n26735 );
not ( n26737 , n17879 );
not ( n26738 , n26737 );
not ( n26739 , n23996 );
or ( n26740 , n26738 , n26739 );
not ( n26741 , n16283 );
buf ( n26742 , n22636 );
not ( n26743 , n26742 );
buf ( n26744 , n22625 );
nand ( n26745 , n26743 , n26744 );
buf ( n26746 , n26745 );
buf ( n26747 , n26746 );
not ( n26748 , n26747 );
buf ( n26749 , n22371 );
buf ( n26750 , n22351 );
not ( n26751 , n26750 );
buf ( n26752 , n26751 );
buf ( n26753 , n26752 );
and ( n26754 , n26749 , n26753 );
buf ( n26755 , n26754 );
buf ( n26756 , n26755 );
not ( n26757 , n26756 );
buf ( n26758 , n22592 );
not ( n26759 , n26758 );
or ( n26760 , n26757 , n26759 );
buf ( n26761 , n22617 );
buf ( n26762 , n26752 );
and ( n26763 , n26761 , n26762 );
buf ( n26764 , n22630 );
nor ( n26765 , n26763 , n26764 );
buf ( n26766 , n26765 );
buf ( n26767 , n26766 );
nand ( n26768 , n26760 , n26767 );
buf ( n26769 , n26768 );
buf ( n26770 , n26769 );
not ( n26771 , n26770 );
or ( n26772 , n26748 , n26771 );
buf ( n26773 , n26769 );
buf ( n26774 , n26746 );
or ( n26775 , n26773 , n26774 );
nand ( n26776 , n26772 , n26775 );
buf ( n26777 , n26776 );
buf ( n26778 , n26777 );
not ( n26779 , n26778 );
or ( n26780 , n26741 , n26779 );
nand ( n26781 , n277983 , n9702 );
nand ( n26782 , n26780 , n26781 );
nand ( n26783 , n19242 , n26782 );
nand ( n26784 , n26740 , n26783 );
buf ( n26785 , n26784 );
not ( n26786 , n26785 );
not ( n26787 , n26786 );
buf ( n26788 , n18604 );
buf ( n26789 , n26788 );
not ( n26790 , n26789 );
not ( n26791 , n26790 );
or ( n26792 , n26787 , n26791 );
nand ( n26793 , n26789 , n26785 );
nand ( n26794 , n26792 , n26793 );
buf ( n26795 , n18628 );
buf ( n26796 , n26795 );
buf ( n26797 , n26796 );
not ( n26798 , n26797 );
not ( n26799 , n17704 );
not ( n26800 , n23996 );
or ( n26801 , n26799 , n26800 );
not ( n26802 , n277527 );
buf ( n26803 , n22630 );
not ( n26804 , n26803 );
buf ( n26805 , n26752 );
nand ( n26806 , n26804 , n26805 );
buf ( n26807 , n26806 );
buf ( n26808 , n26807 );
not ( n26809 , n26808 );
buf ( n26810 , n22371 );
not ( n26811 , n26810 );
buf ( n26812 , n22592 );
not ( n26813 , n26812 );
or ( n26814 , n26811 , n26813 );
buf ( n26815 , n22617 );
not ( n26816 , n26815 );
buf ( n26817 , n26816 );
buf ( n26818 , n26817 );
nand ( n26819 , n26814 , n26818 );
buf ( n26820 , n26819 );
buf ( n26821 , n26820 );
not ( n26822 , n26821 );
or ( n26823 , n26809 , n26822 );
buf ( n26824 , n26820 );
buf ( n26825 , n26807 );
or ( n26826 , n26824 , n26825 );
nand ( n26827 , n26823 , n26826 );
buf ( n26828 , n26827 );
buf ( n26829 , n26828 );
not ( n26830 , n26829 );
or ( n26831 , n26802 , n26830 );
nand ( n26832 , n277351 , n9710 );
nand ( n26833 , n26831 , n26832 );
nand ( n26834 , n19242 , n26833 );
nand ( n26835 , n26801 , n26834 );
buf ( n26836 , n26835 );
nor ( n26837 , n26798 , n26836 );
nor ( n26838 , n26794 , n26837 );
not ( n26839 , n26836 );
not ( n26840 , n26839 );
not ( n26841 , n26797 );
not ( n26842 , n26841 );
or ( n26843 , n26840 , n26842 );
nand ( n26844 , n26797 , n26836 );
nand ( n26845 , n26843 , n26844 );
and ( n26846 , n24056 , n24060 );
nor ( n26847 , n26845 , n26846 );
nor ( n26848 , n26838 , n26847 );
not ( n26849 , n26848 );
not ( n26850 , n24094 );
nand ( n26851 , n26850 , n24161 );
nor ( n26852 , n26849 , n26851 );
not ( n26853 , n26852 );
not ( n26854 , n26730 );
not ( n26855 , n26692 );
or ( n26856 , n26854 , n26855 );
or ( n26857 , n26730 , n26692 );
nand ( n26858 , n26856 , n26857 );
not ( n26859 , n18683 );
not ( n26860 , n26859 );
buf ( n26861 , n26860 );
not ( n26862 , n277527 );
buf ( n26863 , n22649 );
not ( n26864 , n26863 );
buf ( n26865 , n26697 );
nand ( n26866 , n26864 , n26865 );
buf ( n26867 , n26866 );
buf ( n26868 , n26867 );
not ( n26869 , n26868 );
buf ( n26870 , n22374 );
not ( n26871 , n26870 );
buf ( n26872 , n22592 );
not ( n26873 , n26872 );
or ( n26874 , n26871 , n26873 );
buf ( n26875 , n22642 );
not ( n26876 , n26875 );
buf ( n26877 , n26876 );
buf ( n26878 , n26877 );
nand ( n26879 , n26874 , n26878 );
buf ( n26880 , n26879 );
buf ( n26881 , n26880 );
not ( n26882 , n26881 );
or ( n26883 , n26869 , n26882 );
buf ( n26884 , n26880 );
buf ( n26885 , n26867 );
or ( n26886 , n26884 , n26885 );
nand ( n26887 , n26883 , n26886 );
buf ( n26888 , n26887 );
buf ( n26889 , n26888 );
not ( n26890 , n26889 );
or ( n26891 , n26862 , n26890 );
nand ( n26892 , n277390 , n9675 );
nand ( n26893 , n26891 , n26892 );
nand ( n26894 , n19242 , n26893 );
not ( n26895 , n26894 );
buf ( n26896 , n26895 );
not ( n26897 , n26896 );
and ( n26898 , n26861 , n26897 );
nor ( n26899 , n26858 , n26898 );
not ( n26900 , n26899 );
not ( n26901 , n26896 );
not ( n26902 , n26861 );
or ( n26903 , n26901 , n26902 );
not ( n26904 , n26896 );
not ( n26905 , n26861 );
nand ( n26906 , n26904 , n26905 );
nand ( n26907 , n26903 , n26906 );
not ( n26908 , n26907 );
and ( n26909 , n26786 , n26789 );
not ( n26910 , n26909 );
nand ( n26911 , n26908 , n26910 );
nand ( n26912 , n26900 , n26911 );
nor ( n26913 , n26853 , n26912 );
not ( n26914 , n26913 );
not ( n26915 , n24203 );
not ( n26916 , n26915 );
or ( n26917 , n26914 , n26916 );
not ( n26918 , n26912 );
not ( n26919 , n26918 );
or ( n26920 , n24094 , n24207 );
nand ( n26921 , n26920 , n24096 );
nand ( n26922 , n26921 , n26848 );
buf ( n26923 , n26922 );
nand ( n26924 , n26845 , n26846 );
nor ( n26925 , n26838 , n26924 );
and ( n26926 , n26794 , n26837 );
nor ( n26927 , n26925 , n26926 );
nand ( n26928 , n26923 , n26927 );
not ( n26929 , n26928 );
or ( n26930 , n26919 , n26929 );
nand ( n26931 , n26907 , n26909 );
or ( n26932 , n26899 , n26931 );
nand ( n26933 , n26858 , n26898 );
nand ( n26934 , n26932 , n26933 );
buf ( n26935 , n26934 );
not ( n26936 , n26935 );
nand ( n26937 , n26930 , n26936 );
not ( n26938 , n26937 );
nand ( n26939 , n26917 , n26938 );
not ( n26940 , n26939 );
or ( n26941 , n26736 , n26940 );
or ( n26942 , n26939 , n26735 );
nand ( n26943 , n26941 , n26942 );
buf ( n26944 , n26943 );
not ( n26945 , n26944 );
or ( n26946 , n26640 , n26945 );
buf ( n26947 , n26680 );
not ( n26948 , n26947 );
buf ( n26949 , n26683 );
not ( n26950 , n26949 );
not ( n26951 , n26950 );
or ( n26952 , n26948 , n26951 );
not ( n26953 , n26947 );
nand ( n26954 , n26953 , n26949 );
nand ( n26955 , n26952 , n26954 );
buf ( n26956 , n26691 );
buf ( n26957 , n26729 );
and ( n26958 , n26956 , n26957 );
nor ( n26959 , n26955 , n26958 );
not ( n26960 , n26959 );
nand ( n26961 , n26955 , n26958 );
nand ( n26962 , n26960 , n26961 );
not ( n26963 , n26962 );
buf ( n26964 , n26784 );
not ( n26965 , n26964 );
not ( n26966 , n26965 );
buf ( n26967 , n26788 );
not ( n26968 , n26967 );
or ( n26969 , n26966 , n26968 );
not ( n26970 , n26967 );
nand ( n26971 , n26970 , n26964 );
nand ( n26972 , n26969 , n26971 );
buf ( n26973 , n26795 );
buf ( n26974 , n26835 );
nand ( n26975 , n26973 , n26974 );
not ( n26976 , n26975 );
nor ( n26977 , n26972 , n26976 );
not ( n26978 , n26974 );
not ( n26979 , n26978 );
not ( n26980 , n26973 );
or ( n26981 , n26979 , n26980 );
not ( n26982 , n26973 );
nand ( n26983 , n26982 , n26974 );
nand ( n26984 , n26981 , n26983 );
and ( n26985 , n24280 , n24277 );
nor ( n26986 , n26984 , n26985 );
nor ( n26987 , n26977 , n26986 );
not ( n26988 , n26987 );
nand ( n26989 , n24288 , n24228 );
nor ( n26990 , n26988 , n26989 );
not ( n26991 , n26990 );
buf ( n26992 , n26895 );
not ( n26993 , n26992 );
not ( n26994 , n26859 );
buf ( n26995 , n26994 );
not ( n26996 , n26995 );
not ( n26997 , n26996 );
or ( n26998 , n26993 , n26997 );
not ( n26999 , n26992 );
nand ( n27000 , n26999 , n26995 );
nand ( n27001 , n26998 , n27000 );
and ( n27002 , n26964 , n26967 );
nor ( n27003 , n27001 , n27002 );
not ( n27004 , n26957 );
not ( n27005 , n26956 );
not ( n27006 , n27005 );
or ( n27007 , n27004 , n27006 );
not ( n27008 , n26957 );
nand ( n27009 , n26956 , n27008 );
nand ( n27010 , n27007 , n27009 );
and ( n27011 , n26995 , n26992 );
nor ( n27012 , n27010 , n27011 );
nor ( n27013 , n27003 , n27012 );
not ( n27014 , n27013 );
nor ( n27015 , n26991 , n27014 );
not ( n27016 , n27015 );
not ( n27017 , n24250 );
nand ( n27018 , n24258 , n27017 );
not ( n27019 , n27018 );
nand ( n27020 , n27019 , n24272 );
not ( n27021 , n27020 );
or ( n27022 , n27016 , n27021 );
and ( n27023 , n26984 , n26985 );
not ( n27024 , n26977 );
and ( n27025 , n27023 , n27024 );
and ( n27026 , n26972 , n26976 );
nor ( n27027 , n27025 , n27026 );
not ( n27028 , n27027 );
not ( n27029 , n27028 );
or ( n27030 , n24287 , n24253 );
nand ( n27031 , n27030 , n24289 );
and ( n27032 , n27031 , n26987 );
not ( n27033 , n27032 );
nand ( n27034 , n27029 , n27033 );
and ( n27035 , n27013 , n27034 );
nand ( n27036 , n27001 , n27002 );
or ( n27037 , n27012 , n27036 );
nand ( n27038 , n27010 , n27011 );
nand ( n27039 , n27037 , n27038 );
nor ( n27040 , n27035 , n27039 );
nand ( n27041 , n27022 , n27040 );
not ( n27042 , n27041 );
or ( n27043 , n26963 , n27042 );
or ( n27044 , n27041 , n26962 );
nand ( n27045 , n27043 , n27044 );
buf ( n27046 , n27045 );
and ( n27047 , n27046 , n19358 );
buf ( n27048 , n26680 );
buf ( n27049 , n27048 );
buf ( n27050 , n27049 );
not ( n27051 , n27050 );
not ( n27052 , n19219 );
or ( n27053 , n27051 , n27052 );
buf ( n27054 , n27048 );
not ( n27055 , n27054 );
not ( n27056 , n27055 );
nor ( n27057 , n24300 , n24304 );
buf ( n27058 , n26835 );
buf ( n27059 , n27058 );
not ( n27060 , n26784 );
not ( n27061 , n27060 );
buf ( n27062 , n27061 );
nor ( n27063 , n27059 , n27062 );
and ( n27064 , n27057 , n27063 );
not ( n27065 , n27064 );
buf ( n27066 , n26729 );
buf ( n27067 , n27066 );
not ( n27068 , n27067 );
buf ( n27069 , n26895 );
buf ( n27070 , n27069 );
not ( n27071 , n27070 );
nand ( n27072 , n27068 , n27071 );
nor ( n27073 , n27065 , n27072 );
nand ( n27074 , n24314 , n27073 );
not ( n27075 , n27074 );
or ( n27076 , n27056 , n27075 );
or ( n27077 , n27074 , n27055 );
nand ( n27078 , n27076 , n27077 );
buf ( n27079 , n27078 );
nand ( n27080 , n27079 , n19290 );
nand ( n27081 , n27053 , n27080 );
nor ( n27082 , n27047 , n27081 );
nand ( n27083 , n26946 , n27082 );
nor ( n27084 , n26639 , n27083 );
or ( n27085 , n27084 , n21030 );
nand ( n27086 , n21030 , n18568 );
nand ( n27087 , n27085 , n27086 );
buf ( n27088 , n27087 );
buf ( n27089 , n27088 );
not ( n27090 , n275929 );
buf ( n27091 , n27090 );
buf ( n27092 , n27091 );
buf ( n27093 , n275554 );
not ( n27094 , n275925 );
buf ( n27095 , n27094 );
buf ( n27096 , n27095 );
buf ( n27097 , n275554 );
buf ( n27098 , n14448 );
and ( n27099 , n20711 , n27098 );
not ( n27100 , n20711 );
not ( n27101 , n14293 );
not ( n27102 , n27101 );
nand ( n27103 , n20836 , n14213 );
not ( n27104 , n27103 );
not ( n27105 , n27104 );
or ( n27106 , n27102 , n27105 );
not ( n27107 , n27103 );
or ( n27108 , n27107 , n27101 );
nand ( n27109 , n27106 , n27108 );
buf ( n27110 , n27109 );
and ( n27111 , n27100 , n27110 );
nor ( n27112 , n27099 , n27111 );
not ( n27113 , n27112 );
and ( n27114 , n27113 , n26440 );
not ( n27115 , n16245 );
nand ( n27116 , n27115 , n16897 );
not ( n27117 , n27116 );
not ( n27118 , n16401 );
nor ( n27119 , n27118 , n20849 );
not ( n27120 , n27119 );
not ( n27121 , n20875 );
or ( n27122 , n27120 , n27121 );
or ( n27123 , n20879 , n20849 );
nand ( n27124 , n27123 , n16901 );
not ( n27125 , n27124 );
nand ( n27126 , n27122 , n27125 );
not ( n27127 , n27126 );
or ( n27128 , n27117 , n27127 );
or ( n27129 , n27126 , n27116 );
nand ( n27130 , n27128 , n27129 );
buf ( n27131 , n27130 );
nand ( n27132 , n27131 , n20889 );
nand ( n27133 , n17194 , n17333 );
not ( n27134 , n27133 );
not ( n27135 , n17228 );
not ( n27136 , n17207 );
nor ( n27137 , n27135 , n27136 );
not ( n27138 , n27137 );
not ( n27139 , n20913 );
or ( n27140 , n27138 , n27139 );
or ( n27141 , n20918 , n27136 );
nand ( n27142 , n27141 , n20891 );
not ( n27143 , n27142 );
nand ( n27144 , n27140 , n27143 );
not ( n27145 , n27144 );
or ( n27146 , n27134 , n27145 );
or ( n27147 , n27144 , n27133 );
nand ( n27148 , n27146 , n27147 );
buf ( n27149 , n27148 );
nand ( n27150 , n27149 , n20927 );
nand ( n27151 , n20931 , n20932 );
not ( n27152 , n17444 );
nor ( n27153 , n27151 , n27152 );
not ( n27154 , n27153 );
nand ( n27155 , n27151 , n27152 );
nand ( n27156 , n27154 , n27155 );
buf ( n27157 , n27156 );
and ( n27158 , n27157 , n17409 );
buf ( n27159 , n17443 );
buf ( n27160 , n27159 );
buf ( n27161 , n27160 );
and ( n27162 , n17499 , n27161 );
nor ( n27163 , n27158 , n27162 );
nand ( n27164 , n27132 , n27150 , n27163 );
nor ( n27165 , n27114 , n27164 );
or ( n27166 , n27165 , n20950 );
nand ( n27167 , n20953 , n13464 );
nand ( n27168 , n27166 , n27167 );
buf ( n27169 , n27168 );
buf ( n27170 , n27169 );
not ( n27171 , n275549 );
not ( n27172 , n27171 );
buf ( n27173 , n27172 );
buf ( n27174 , n27173 );
not ( n27175 , n275929 );
buf ( n27176 , n27175 );
buf ( n27177 , n27176 );
not ( n27178 , n278066 );
buf ( n27179 , n23708 );
not ( n27180 , n27179 );
or ( n27181 , n27178 , n27180 );
buf ( n27182 , n10627 );
not ( n27183 , n27182 );
buf ( n27184 , n10647 );
nand ( n27185 , n27183 , n27184 );
nor ( n27186 , n27183 , n27184 );
not ( n27187 , n27186 );
nand ( n27188 , n27185 , n27187 );
not ( n27189 , n27188 );
nor ( n27190 , n22089 , n23632 );
not ( n27191 , n27190 );
not ( n27192 , n22108 );
not ( n27193 , n27192 );
not ( n27194 , n22119 );
nand ( n27195 , n27194 , n22123 );
buf ( n27196 , n22114 );
nand ( n27197 , n22126 , n27195 , n27196 );
not ( n27198 , n27197 );
or ( n27199 , n27193 , n27198 );
not ( n27200 , n22100 );
nor ( n27201 , n22132 , n27200 );
nand ( n27202 , n27199 , n27201 );
not ( n27203 , n27202 );
or ( n27204 , n27191 , n27203 );
buf ( n27205 , n11483 );
not ( n27206 , n27205 );
buf ( n27207 , n11516 );
nand ( n27208 , n27206 , n27207 );
nand ( n27209 , n23608 , n27208 );
nor ( n27210 , n27209 , n23621 );
buf ( n27211 , n11421 );
buf ( n27212 , n27211 );
not ( n27213 , n27212 );
buf ( n27214 , n11457 );
nand ( n27215 , n27213 , n27214 );
buf ( n27216 , n11396 );
not ( n27217 , n27216 );
buf ( n27218 , n11368 );
nand ( n27219 , n27217 , n27218 );
buf ( n27220 , n11262 );
not ( n27221 , n27220 );
buf ( n27222 , n11240 );
nand ( n27223 , n27221 , n27222 );
buf ( n27224 , n11295 );
not ( n27225 , n27224 );
buf ( n27226 , n11333 );
nand ( n27227 , n27225 , n27226 );
and ( n27228 , n27215 , n27219 , n27223 , n27227 );
not ( n27229 , n22073 );
and ( n27230 , n27229 , n22067 );
nor ( n27231 , n27230 , n22063 );
and ( n27232 , n27210 , n27228 , n27231 );
nand ( n27233 , n27204 , n27232 );
not ( n27234 , n27207 );
nand ( n27235 , n27205 , n27234 );
and ( n27236 , n23610 , n27235 , n23645 );
nand ( n27237 , n27236 , n23643 );
buf ( n27238 , n27235 );
nand ( n27239 , n27209 , n27238 );
nand ( n27240 , n27237 , n27239 , n27228 );
not ( n27241 , n27216 );
nor ( n27242 , n27241 , n27218 );
not ( n27243 , n27242 );
not ( n27244 , n27215 );
or ( n27245 , n27243 , n27244 );
not ( n27246 , n27214 );
buf ( n27247 , n27212 );
nand ( n27248 , n27246 , n27247 );
nand ( n27249 , n27245 , n27248 );
not ( n27250 , n27227 );
not ( n27251 , n27223 );
nor ( n27252 , n27250 , n27251 );
nand ( n27253 , n27249 , n27252 );
not ( n27254 , n27220 );
nor ( n27255 , n27254 , n27222 );
and ( n27256 , n27255 , n27227 );
nor ( n27257 , n27225 , n27226 );
nor ( n27258 , n27256 , n27257 );
and ( n27259 , n27240 , n27253 , n27258 );
nand ( n27260 , n27233 , n27259 );
not ( n27261 , n27260 );
or ( n27262 , n27189 , n27261 );
or ( n27263 , n27260 , n27188 );
nand ( n27264 , n27262 , n27263 );
buf ( n27265 , n27264 );
not ( n27266 , n22056 );
nand ( n27267 , n27265 , n27266 );
buf ( n27268 , n10627 );
buf ( n27269 , n27268 );
buf ( n27270 , n10647 );
buf ( n27271 , n27270 );
and ( n27272 , n27269 , n27271 );
buf ( n27273 , n27272 );
buf ( n27274 , n27273 );
not ( n27275 , n27274 );
buf ( n27276 , n27275 );
buf ( n27277 , n27276 );
buf ( n27278 , n27268 );
buf ( n27279 , n27270 );
or ( n27280 , n27278 , n27279 );
buf ( n27281 , n27280 );
buf ( n27282 , n27281 );
nand ( n27283 , n27277 , n27282 );
buf ( n27284 , n27283 );
buf ( n27285 , n27284 );
not ( n27286 , n27285 );
buf ( n27287 , n21842 );
buf ( n27288 , n23562 );
nor ( n27289 , n27287 , n27288 );
buf ( n27290 , n27289 );
buf ( n27291 , n27290 );
not ( n27292 , n27291 );
buf ( n27293 , n23542 );
buf ( n27294 , n23536 );
nand ( n27295 , n27293 , n27294 );
buf ( n27296 , n27295 );
buf ( n27297 , n27296 );
not ( n27298 , n27297 );
or ( n27299 , n27292 , n27298 );
buf ( n27300 , n23476 );
buf ( n27301 , n11483 );
buf ( n27302 , n27301 );
not ( n27303 , n27302 );
buf ( n27304 , n27303 );
buf ( n27305 , n27304 );
buf ( n27306 , n11516 );
buf ( n27307 , n27306 );
not ( n27308 , n27307 );
buf ( n27309 , n27308 );
buf ( n27310 , n27309 );
nand ( n27311 , n27305 , n27310 );
buf ( n27312 , n27311 );
buf ( n27313 , n27312 );
nand ( n27314 , n27300 , n27313 );
buf ( n27315 , n27314 );
buf ( n27316 , n27315 );
buf ( n27317 , n23514 );
nor ( n27318 , n27316 , n27317 );
buf ( n27319 , n27318 );
buf ( n27320 , n27319 );
buf ( n27321 , n21802 );
buf ( n27322 , n21976 );
and ( n27323 , n27321 , n27322 );
buf ( n27324 , n21970 );
not ( n27325 , n27324 );
buf ( n27326 , n27325 );
buf ( n27327 , n27326 );
nor ( n27328 , n27323 , n27327 );
buf ( n27329 , n27328 );
buf ( n27330 , n27329 );
buf ( n27331 , n27211 );
buf ( n27332 , n27331 );
not ( n27333 , n27332 );
buf ( n27334 , n27333 );
buf ( n27335 , n27334 );
buf ( n27336 , n11457 );
buf ( n27337 , n27336 );
not ( n27338 , n27337 );
buf ( n27339 , n27338 );
buf ( n27340 , n27339 );
nand ( n27341 , n27335 , n27340 );
buf ( n27342 , n27341 );
buf ( n27343 , n27342 );
buf ( n27344 , n11396 );
not ( n27345 , n27344 );
buf ( n27346 , n27345 );
buf ( n27347 , n27346 );
buf ( n27348 , n11368 );
buf ( n27349 , n27348 );
not ( n27350 , n27349 );
buf ( n27351 , n27350 );
buf ( n27352 , n27351 );
nand ( n27353 , n27347 , n27352 );
buf ( n27354 , n27353 );
buf ( n27355 , n27354 );
buf ( n27356 , n11262 );
buf ( n27357 , n27356 );
not ( n27358 , n27357 );
buf ( n27359 , n27358 );
buf ( n27360 , n27359 );
buf ( n27361 , n11240 );
buf ( n27362 , n27361 );
not ( n27363 , n27362 );
buf ( n27364 , n27363 );
buf ( n27365 , n27364 );
nand ( n27366 , n27360 , n27365 );
buf ( n27367 , n27366 );
buf ( n27368 , n27367 );
buf ( n27369 , n11295 );
buf ( n27370 , n27369 );
not ( n27371 , n27370 );
buf ( n27372 , n27371 );
buf ( n27373 , n27372 );
buf ( n27374 , n11333 );
buf ( n27375 , n27374 );
not ( n27376 , n27375 );
buf ( n27377 , n27376 );
buf ( n27378 , n27377 );
nand ( n27379 , n27373 , n27378 );
buf ( n27380 , n27379 );
buf ( n27381 , n27380 );
and ( n27382 , n27343 , n27355 , n27368 , n27381 );
buf ( n27383 , n27382 );
buf ( n27384 , n27383 );
and ( n27385 , n27320 , n27330 , n27384 );
buf ( n27386 , n27385 );
buf ( n27387 , n27386 );
nand ( n27388 , n27299 , n27387 );
buf ( n27389 , n27388 );
buf ( n27390 , n27389 );
buf ( n27391 , n27315 );
buf ( n27392 , n27301 );
buf ( n27393 , n27306 );
nand ( n27394 , n27392 , n27393 );
buf ( n27395 , n27394 );
buf ( n27396 , n27395 );
nand ( n27397 , n27391 , n27396 );
buf ( n27398 , n27397 );
buf ( n27399 , n27398 );
not ( n27400 , n27399 );
buf ( n27401 , n27383 );
not ( n27402 , n27401 );
buf ( n27403 , n27402 );
buf ( n27404 , n27403 );
nor ( n27405 , n27400 , n27404 );
buf ( n27406 , n27405 );
buf ( n27407 , n27406 );
buf ( n27408 , n23481 );
buf ( n27409 , n27395 );
buf ( n27410 , n23584 );
and ( n27411 , n27408 , n27409 , n27410 );
buf ( n27412 , n27411 );
buf ( n27413 , n27412 );
buf ( n27414 , n23579 );
nand ( n27415 , n27413 , n27414 );
buf ( n27416 , n27415 );
buf ( n27417 , n27416 );
and ( n27418 , n27407 , n27417 );
buf ( n27419 , n27367 );
not ( n27420 , n27419 );
buf ( n27421 , n27420 );
buf ( n27422 , n27421 );
buf ( n27423 , n27380 );
not ( n27424 , n27423 );
buf ( n27425 , n27424 );
buf ( n27426 , n27425 );
nor ( n27427 , n27422 , n27426 );
buf ( n27428 , n27427 );
buf ( n27429 , n27428 );
not ( n27430 , n27429 );
buf ( n27431 , n27346 );
buf ( n27432 , n27351 );
nor ( n27433 , n27431 , n27432 );
buf ( n27434 , n27433 );
buf ( n27435 , n27434 );
not ( n27436 , n27435 );
buf ( n27437 , n27342 );
not ( n27438 , n27437 );
or ( n27439 , n27436 , n27438 );
buf ( n27440 , n27331 );
buf ( n27441 , n27336 );
nand ( n27442 , n27440 , n27441 );
buf ( n27443 , n27442 );
buf ( n27444 , n27443 );
nand ( n27445 , n27439 , n27444 );
buf ( n27446 , n27445 );
buf ( n27447 , n27446 );
not ( n27448 , n27447 );
or ( n27449 , n27430 , n27448 );
buf ( n27450 , n27425 );
buf ( n27451 , n27356 );
buf ( n27452 , n27364 );
not ( n27453 , n27452 );
buf ( n27454 , n27453 );
buf ( n27455 , n27454 );
nand ( n27456 , n27451 , n27455 );
buf ( n27457 , n27456 );
buf ( n27458 , n27457 );
or ( n27459 , n27450 , n27458 );
buf ( n27460 , n27372 );
buf ( n27461 , n27377 );
or ( n27462 , n27460 , n27461 );
buf ( n27463 , n27462 );
buf ( n27464 , n27463 );
nand ( n27465 , n27459 , n27464 );
buf ( n27466 , n27465 );
buf ( n27467 , n27466 );
not ( n27468 , n27467 );
buf ( n27469 , n27468 );
buf ( n27470 , n27469 );
nand ( n27471 , n27449 , n27470 );
buf ( n27472 , n27471 );
buf ( n27473 , n27472 );
nor ( n27474 , n27418 , n27473 );
buf ( n27475 , n27474 );
buf ( n27476 , n27475 );
nand ( n27477 , n27390 , n27476 );
buf ( n27478 , n27477 );
buf ( n27479 , n27478 );
buf ( n27480 , n27479 );
not ( n27481 , n27480 );
or ( n27482 , n27286 , n27481 );
buf ( n27483 , n27479 );
buf ( n27484 , n27284 );
or ( n27485 , n27483 , n27484 );
nand ( n27486 , n27482 , n27485 );
buf ( n27487 , n27486 );
buf ( n27488 , n27487 );
buf ( n27489 , n22002 );
nand ( n27490 , n27488 , n27489 );
buf ( n27491 , n278025 );
buf ( n27492 , n27491 );
not ( n27493 , n27492 );
not ( n27494 , n27493 );
buf ( n27495 , n22033 );
buf ( n27496 , n11396 );
buf ( n27497 , n11295 );
nand ( n27498 , n27496 , n23660 , n27497 );
buf ( n27499 , n11421 );
nand ( n27500 , n22043 , n23663 , n23657 , n27499 );
nor ( n27501 , n27498 , n27500 );
buf ( n27502 , n10627 );
nand ( n27503 , n27495 , n27501 , n27502 );
not ( n27504 , n22036 );
not ( n27505 , n22035 );
nor ( n27506 , n27504 , n27505 );
nand ( n27507 , n22039 , n22021 );
nor ( n27508 , n22020 , n27507 );
buf ( n27509 , n11262 );
and ( n27510 , n22022 , n27509 );
nand ( n27511 , n27506 , n27508 , n27510 );
nor ( n27512 , n27503 , n27511 );
buf ( n27513 , n27512 );
not ( n27514 , n27513 );
or ( n27515 , n27494 , n27514 );
or ( n27516 , n27513 , n27493 );
nand ( n27517 , n27515 , n27516 );
buf ( n27518 , n27517 );
and ( n27519 , n27518 , n22052 );
buf ( n27520 , n22007 );
not ( n27521 , n27520 );
or ( n27522 , n27521 , n12174 );
or ( n27523 , n23680 , n12291 );
nand ( n27524 , n27522 , n27523 );
nor ( n27525 , n27519 , n27524 );
and ( n27526 , n27267 , n27490 , n27525 );
or ( n27527 , n27526 , n27179 );
nand ( n27528 , n27181 , n27527 );
buf ( n27529 , n27528 );
buf ( n27530 , n27529 );
buf ( n27531 , n275554 );
buf ( n27532 , n21945 );
buf ( n27533 , n21813 );
not ( n27534 , n27533 );
buf ( n27535 , n27534 );
buf ( n27536 , n27535 );
nand ( n27537 , n27532 , n27536 );
buf ( n27538 , n27537 );
buf ( n27539 , n27538 );
not ( n27540 , n27539 );
buf ( n27541 , n21869 );
not ( n27542 , n27541 );
buf ( n27543 , n21885 );
not ( n27544 , n27543 );
or ( n27545 , n27542 , n27544 );
buf ( n27546 , n21935 );
nand ( n27547 , n27545 , n27546 );
buf ( n27548 , n27547 );
buf ( n27549 , n27548 );
not ( n27550 , n27549 );
or ( n27551 , n27540 , n27550 );
buf ( n27552 , n21945 );
buf ( n27553 , n27535 );
nand ( n27554 , n27552 , n27553 );
buf ( n27555 , n27554 );
buf ( n27556 , n27555 );
buf ( n27557 , n27548 );
or ( n27558 , n27556 , n27557 );
nand ( n27559 , n27551 , n27558 );
buf ( n27560 , n27559 );
buf ( n27561 , n27560 );
and ( n27562 , n27561 , n22002 );
not ( n27563 , n12189 );
not ( n27564 , n22007 );
or ( n27565 , n27563 , n27564 );
nand ( n27566 , n23679 , n12233 );
nand ( n27567 , n27565 , n27566 );
nor ( n27568 , n27562 , n27567 );
buf ( n27569 , n22034 );
buf ( n27570 , n22036 );
not ( n27571 , n27570 );
and ( n27572 , n27569 , n27571 );
not ( n27573 , n27569 );
and ( n27574 , n27573 , n27570 );
nor ( n27575 , n27572 , n27574 );
buf ( n27576 , n27575 );
nand ( n27577 , n27576 , n23672 );
buf ( n27578 , n22131 );
not ( n27579 , n22079 );
nand ( n27580 , n27578 , n27579 );
not ( n27581 , n27580 );
not ( n27582 , n22128 );
or ( n27583 , n27581 , n27582 );
or ( n27584 , n22128 , n27580 );
nand ( n27585 , n27583 , n27584 );
buf ( n27586 , n27585 );
nand ( n27587 , n27586 , n22057 );
and ( n27588 , n27568 , n27577 , n27587 );
not ( n27589 , n22191 );
buf ( n27590 , n27589 );
or ( n27591 , n27588 , n27590 );
not ( n27592 , n10868 );
or ( n27593 , n22192 , n27592 );
nand ( n27594 , n27591 , n27593 );
buf ( n27595 , n27594 );
buf ( n27596 , n27595 );
buf ( n27597 , n275554 );
buf ( n27598 , n275554 );
buf ( n27599 , n275554 );
not ( n27600 , n275550 );
buf ( n27601 , n27600 );
buf ( n27602 , n27601 );
buf ( n27603 , n275554 );
not ( n27604 , n275929 );
buf ( n27605 , n27604 );
buf ( n27606 , n27605 );
not ( n27607 , n275550 );
buf ( n27608 , n27607 );
buf ( n27609 , n27608 );
not ( n27610 , n19629 );
and ( n27611 , n27610 , n21174 );
not ( n27612 , n21001 );
not ( n27613 , n20352 );
or ( n27614 , n27612 , n27613 );
and ( n27615 , n20514 , n19358 );
not ( n27616 , n19290 );
not ( n27617 , n20558 );
or ( n27618 , n27616 , n27617 );
not ( n27619 , n24440 );
nand ( n27620 , n27619 , n20566 );
nand ( n27621 , n27618 , n27620 );
nor ( n27622 , n27615 , n27621 );
nand ( n27623 , n27614 , n27622 );
nor ( n27624 , n27611 , n27623 );
or ( n27625 , n27624 , n21030 );
nand ( n27626 , n21030 , n18763 );
nand ( n27627 , n27625 , n27626 );
buf ( n27628 , n27627 );
buf ( n27629 , n27628 );
not ( n27630 , n275550 );
buf ( n27631 , n27630 );
buf ( n27632 , n27631 );
buf ( n27633 , n275554 );
buf ( n27634 , n275554 );
buf ( n27635 , n275554 );
not ( n27636 , n275550 );
buf ( n27637 , n27636 );
buf ( n27638 , n27637 );
or ( n27639 , n27588 , n23708 );
not ( n27640 , n23703 );
buf ( n27641 , n27640 );
nand ( n27642 , n27641 , n10881 );
nand ( n27643 , n27639 , n27642 );
buf ( n27644 , n27643 );
buf ( n27645 , n27644 );
or ( n27646 , n24623 , n21697 );
buf ( n27647 , n21696 );
nand ( n27648 , n27647 , n14025 );
nand ( n27649 , n27646 , n27648 );
buf ( n27650 , n27649 );
buf ( n27651 , n27650 );
not ( n27652 , n275550 );
buf ( n27653 , n27652 );
buf ( n27654 , n27653 );
not ( n27655 , n275929 );
buf ( n27656 , n27655 );
buf ( n27657 , n27656 );
not ( n27658 , n275550 );
buf ( n27659 , n27658 );
buf ( n27660 , n27659 );
buf ( n27661 , n275554 );
buf ( n27662 , n275554 );
not ( n27663 , n13254 );
not ( n27664 , n14830 );
not ( n27665 , n27664 );
not ( n27666 , n27665 );
or ( n27667 , n27663 , n27666 );
not ( n27668 , n15507 );
or ( n27669 , n27668 , n27665 );
nand ( n27670 , n27667 , n27669 );
buf ( n27671 , n27670 );
buf ( n27672 , n27671 );
not ( n27673 , n275550 );
buf ( n27674 , n27673 );
buf ( n27675 , n27674 );
and ( n27676 , n14830 , n13084 );
not ( n27677 , n14830 );
and ( n27678 , n27677 , n16750 );
or ( n27679 , n27676 , n27678 );
buf ( n27680 , n27679 );
buf ( n27681 , n27680 );
buf ( n27682 , n275554 );
buf ( n27683 , n275554 );
buf ( n27684 , n275554 );
buf ( n27685 , n14211 );
and ( n27686 , n20711 , n27685 );
not ( n27687 , n20711 );
not ( n27688 , n26426 );
buf ( n27689 , n20720 );
not ( n27690 , n27689 );
or ( n27691 , n27688 , n27690 );
or ( n27692 , n27689 , n26426 );
nand ( n27693 , n27691 , n27692 );
buf ( n27694 , n27693 );
and ( n27695 , n27687 , n27694 );
nor ( n27696 , n27686 , n27695 );
not ( n27697 , n27696 );
and ( n27698 , n27697 , n23404 );
not ( n27699 , n20889 );
not ( n27700 , n26446 );
nand ( n27701 , n27700 , n16888 );
not ( n27702 , n27701 );
not ( n27703 , n16402 );
not ( n27704 , n20875 );
or ( n27705 , n27703 , n27704 );
nand ( n27706 , n27705 , n26451 );
not ( n27707 , n27706 );
or ( n27708 , n27702 , n27707 );
or ( n27709 , n27706 , n27701 );
nand ( n27710 , n27708 , n27709 );
buf ( n27711 , n27710 );
not ( n27712 , n27711 );
or ( n27713 , n27699 , n27712 );
or ( n27714 , n17346 , n26466 );
not ( n27715 , n27714 );
not ( n27716 , n23742 );
not ( n27717 , n20913 );
or ( n27718 , n27716 , n27717 );
nand ( n27719 , n27718 , n26473 );
not ( n27720 , n27719 );
or ( n27721 , n27715 , n27720 );
or ( n27722 , n27719 , n27714 );
nand ( n27723 , n27721 , n27722 );
buf ( n27724 , n27723 );
and ( n27725 , n27724 , n24711 );
buf ( n27726 , n17453 );
buf ( n27727 , n27726 );
buf ( n27728 , n27727 );
not ( n27729 , n27728 );
not ( n27730 , n20940 );
or ( n27731 , n27729 , n27730 );
nand ( n27732 , n26486 , n26487 );
and ( n27733 , n27732 , n17454 );
not ( n27734 , n27732 );
and ( n27735 , n27734 , n17455 );
nor ( n27736 , n27733 , n27735 );
buf ( n27737 , n27736 );
nand ( n27738 , n27737 , n17409 );
nand ( n27739 , n27731 , n27738 );
nor ( n27740 , n27725 , n27739 );
nand ( n27741 , n27713 , n27740 );
nor ( n27742 , n27698 , n27741 );
or ( n27743 , n27742 , n20950 );
nand ( n27744 , n20953 , n13721 );
nand ( n27745 , n27743 , n27744 );
buf ( n27746 , n27745 );
buf ( n27747 , n27746 );
buf ( n27748 , n275554 );
not ( n27749 , n275929 );
buf ( n27750 , n27749 );
buf ( n27751 , n27750 );
not ( n27752 , n275925 );
buf ( n27753 , n27752 );
buf ( n27754 , n27753 );
buf ( n27755 , n275554 );
buf ( n27756 , n21726 );
buf ( n27757 , n21731 );
buf ( n27758 , n26524 );
buf ( n27759 , n18576 );
nor ( n27760 , n27758 , n27759 );
buf ( n27761 , n27760 );
buf ( n27762 , n27761 );
nand ( n27763 , n27757 , n27762 );
buf ( n27764 , n27763 );
buf ( n27765 , n27764 );
not ( n27766 , n27765 );
buf ( n27767 , n27766 );
buf ( n27768 , n27767 );
nand ( n27769 , n27756 , n27768 );
buf ( n27770 , n27769 );
buf ( n27771 , n27770 );
buf ( n27772 , n18809 );
not ( n27773 , n27772 );
buf ( n27774 , n27773 );
buf ( n27775 , n27774 );
and ( n27776 , n27771 , n27775 );
not ( n27777 , n27771 );
buf ( n27778 , n18809 );
and ( n27779 , n27777 , n27778 );
nor ( n27780 , n27776 , n27779 );
buf ( n27781 , n27780 );
buf ( n27782 , n27781 );
buf ( n27783 , n27782 );
and ( n27784 , n26516 , n27783 );
not ( n27785 , n26516 );
buf ( n27786 , n23914 );
not ( n27787 , n27786 );
buf ( n27788 , n27764 );
buf ( n27789 , n18658 );
buf ( n27790 , n18809 );
nand ( n27791 , n27789 , n27790 );
buf ( n27792 , n27791 );
buf ( n27793 , n27792 );
not ( n27794 , n27793 );
buf ( n27795 , n27794 );
buf ( n27796 , n27795 );
not ( n27797 , n27796 );
buf ( n27798 , n27797 );
buf ( n27799 , n27798 );
nor ( n27800 , n27788 , n27799 );
buf ( n27801 , n27800 );
buf ( n27802 , n27801 );
nand ( n27803 , n27787 , n27802 );
buf ( n27804 , n27803 );
buf ( n27805 , n27804 );
buf ( n27806 , n18492 );
buf ( n27807 , n27806 );
xnor ( n27808 , n27805 , n27807 );
buf ( n27809 , n27808 );
buf ( n27810 , n27809 );
buf ( n27811 , n27810 );
buf ( n27812 , n27811 );
not ( n27813 , n27812 );
buf ( n27814 , n27782 );
nand ( n27815 , n27814 , n26552 );
nor ( n27816 , n27815 , n26629 );
nand ( n27817 , n19069 , n27816 );
nor ( n27818 , n27817 , n26601 );
buf ( n27819 , n23914 );
not ( n27820 , n27819 );
buf ( n27821 , n27764 );
buf ( n27822 , n27774 );
nor ( n27823 , n27821 , n27822 );
buf ( n27824 , n27823 );
buf ( n27825 , n27824 );
nand ( n27826 , n27820 , n27825 );
buf ( n27827 , n27826 );
buf ( n27828 , n27827 );
buf ( n27829 , n18658 );
xnor ( n27830 , n27828 , n27829 );
buf ( n27831 , n27830 );
buf ( n27832 , n27831 );
buf ( n27833 , n27832 );
buf ( n27834 , n27833 );
nand ( n27835 , n27818 , n27834 );
buf ( n27836 , n27835 );
not ( n27837 , n27836 );
or ( n27838 , n27813 , n27837 );
or ( n27839 , n27812 , n27836 );
nand ( n27840 , n27838 , n27839 );
buf ( n27841 , n27840 );
and ( n27842 , n27785 , n27841 );
nor ( n27843 , n27784 , n27842 );
not ( n27844 , n27843 );
buf ( n27845 , n21174 );
and ( n27846 , n27844 , n27845 );
not ( n27847 , n9432 );
buf ( n27848 , n22439 );
buf ( n27849 , n22705 );
nand ( n27850 , n27848 , n27849 );
buf ( n27851 , n27850 );
buf ( n27852 , n27851 );
not ( n27853 , n27852 );
buf ( n27854 , n22415 );
buf ( n27855 , n22446 );
and ( n27856 , n27854 , n27855 );
buf ( n27857 , n27856 );
buf ( n27858 , n27857 );
not ( n27859 , n27858 );
buf ( n27860 , n22593 );
not ( n27861 , n27860 );
or ( n27862 , n27859 , n27861 );
buf ( n27863 , n22687 );
buf ( n27864 , n22446 );
and ( n27865 , n27863 , n27864 );
buf ( n27866 , n22698 );
nor ( n27867 , n27865 , n27866 );
buf ( n27868 , n27867 );
buf ( n27869 , n27868 );
nand ( n27870 , n27862 , n27869 );
buf ( n27871 , n27870 );
buf ( n27872 , n27871 );
not ( n27873 , n27872 );
or ( n27874 , n27853 , n27873 );
buf ( n27875 , n27871 );
buf ( n27876 , n27851 );
or ( n27877 , n27875 , n27876 );
nand ( n27878 , n27874 , n27877 );
buf ( n27879 , n27878 );
buf ( n27880 , n27879 );
not ( n27881 , n27880 );
or ( n27882 , n27847 , n27881 );
nand ( n27883 , n277390 , n9757 );
nand ( n27884 , n27882 , n27883 );
and ( n27885 , n19242 , n27884 );
buf ( n27886 , n27885 );
not ( n27887 , n27886 );
buf ( n27888 , n18657 );
buf ( n27889 , n27888 );
not ( n27890 , n27889 );
or ( n27891 , n27887 , n27890 );
not ( n27892 , n27889 );
not ( n27893 , n27886 );
nand ( n27894 , n27892 , n27893 );
nand ( n27895 , n27891 , n27894 );
not ( n27896 , n27895 );
buf ( n27897 , n18808 );
buf ( n27898 , n27897 );
not ( n27899 , n277603 );
buf ( n27900 , n22698 );
not ( n27901 , n27900 );
buf ( n27902 , n22446 );
nand ( n27903 , n27901 , n27902 );
buf ( n27904 , n27903 );
buf ( n27905 , n27904 );
not ( n27906 , n27905 );
buf ( n27907 , n22415 );
not ( n27908 , n27907 );
buf ( n27909 , n22593 );
not ( n27910 , n27909 );
or ( n27911 , n27908 , n27910 );
buf ( n27912 , n22687 );
not ( n27913 , n27912 );
buf ( n27914 , n27913 );
buf ( n27915 , n27914 );
nand ( n27916 , n27911 , n27915 );
buf ( n27917 , n27916 );
buf ( n27918 , n27917 );
not ( n27919 , n27918 );
or ( n27920 , n27906 , n27919 );
buf ( n27921 , n27917 );
buf ( n27922 , n27904 );
or ( n27923 , n27921 , n27922 );
nand ( n27924 , n27920 , n27923 );
buf ( n27925 , n27924 );
buf ( n27926 , n27925 );
not ( n27927 , n27926 );
or ( n27928 , n27899 , n27927 );
nand ( n27929 , n277351 , n9765 );
nand ( n27930 , n27928 , n27929 );
nand ( n27931 , n25049 , n27930 );
not ( n27932 , n27931 );
buf ( n27933 , n27932 );
not ( n27934 , n27933 );
and ( n27935 , n27898 , n27934 );
not ( n27936 , n27935 );
nand ( n27937 , n27896 , n27936 );
not ( n27938 , n27937 );
not ( n27939 , n27938 );
nand ( n27940 , n27895 , n27935 );
nand ( n27941 , n27939 , n27940 );
not ( n27942 , n27941 );
not ( n27943 , n277603 );
buf ( n27944 , n22406 );
not ( n27945 , n27944 );
buf ( n27946 , n22678 );
nand ( n27947 , n27945 , n27946 );
buf ( n27948 , n27947 );
buf ( n27949 , n27948 );
not ( n27950 , n27949 );
buf ( n27951 , n22392 );
not ( n27952 , n27951 );
buf ( n27953 , n22399 );
nor ( n27954 , n27952 , n27953 );
buf ( n27955 , n27954 );
buf ( n27956 , n27955 );
buf ( n27957 , n22374 );
and ( n27958 , n27956 , n27957 );
buf ( n27959 , n27958 );
buf ( n27960 , n27959 );
not ( n27961 , n27960 );
buf ( n27962 , n22593 );
not ( n27963 , n27962 );
or ( n27964 , n27961 , n27963 );
buf ( n27965 , n22642 );
buf ( n27966 , n27955 );
and ( n27967 , n27965 , n27966 );
buf ( n27968 , n22664 );
not ( n27969 , n27968 );
buf ( n27970 , n27969 );
buf ( n27971 , n27970 );
buf ( n27972 , n22399 );
or ( n27973 , n27971 , n27972 );
buf ( n27974 , n22671 );
nand ( n27975 , n27973 , n27974 );
buf ( n27976 , n27975 );
buf ( n27977 , n27976 );
nor ( n27978 , n27967 , n27977 );
buf ( n27979 , n27978 );
buf ( n27980 , n27979 );
nand ( n27981 , n27964 , n27980 );
buf ( n27982 , n27981 );
buf ( n27983 , n27982 );
not ( n27984 , n27983 );
or ( n27985 , n27950 , n27984 );
buf ( n27986 , n27982 );
buf ( n27987 , n27948 );
or ( n27988 , n27986 , n27987 );
nand ( n27989 , n27985 , n27988 );
buf ( n27990 , n27989 );
buf ( n27991 , n27990 );
not ( n27992 , n27991 );
or ( n27993 , n27943 , n27992 );
nand ( n27994 , n277390 , n9684 );
nand ( n27995 , n27993 , n27994 );
nand ( n27996 , n19242 , n27995 );
not ( n27997 , n27996 );
buf ( n27998 , n27997 );
not ( n27999 , n27998 );
buf ( n28000 , n18547 );
buf ( n28001 , n28000 );
not ( n28002 , n28001 );
or ( n28003 , n27999 , n28002 );
not ( n28004 , n27998 );
not ( n28005 , n28001 );
nand ( n28006 , n28004 , n28005 );
nand ( n28007 , n28003 , n28006 );
not ( n28008 , n26681 );
and ( n28009 , n26684 , n28008 );
nor ( n28010 , n28007 , n28009 );
not ( n28011 , n28010 );
nand ( n28012 , n28011 , n26733 );
nor ( n28013 , n28012 , n26912 );
nand ( n28014 , n26852 , n28013 );
not ( n28015 , n27933 );
not ( n28016 , n27898 );
or ( n28017 , n28015 , n28016 );
or ( n28018 , n27898 , n27933 );
nand ( n28019 , n28017 , n28018 );
not ( n28020 , n27998 );
and ( n28021 , n28001 , n28020 );
nor ( n28022 , n28019 , n28021 );
buf ( n28023 , n28022 );
nor ( n28024 , n28014 , n28023 );
not ( n28025 , n28024 );
not ( n28026 , n24204 );
or ( n28027 , n28025 , n28026 );
or ( n28028 , n28010 , n26734 );
nand ( n28029 , n28007 , n28009 );
nand ( n28030 , n28028 , n28029 );
nor ( n28031 , n28030 , n26934 );
nand ( n28032 , n28031 , n26922 , n26927 );
nand ( n28033 , n28031 , n26912 );
not ( n28034 , n28030 );
nand ( n28035 , n28034 , n28012 );
and ( n28036 , n28032 , n28033 , n28035 );
not ( n28037 , n28036 );
not ( n28038 , n28037 );
not ( n28039 , n28023 );
and ( n28040 , n28038 , n28039 );
nand ( n28041 , n28019 , n28021 );
not ( n28042 , n28041 );
nor ( n28043 , n28040 , n28042 );
nand ( n28044 , n28027 , n28043 );
not ( n28045 , n28044 );
or ( n28046 , n27942 , n28045 );
or ( n28047 , n28044 , n27941 );
nand ( n28048 , n28046 , n28047 );
buf ( n28049 , n28048 );
nand ( n28050 , n28049 , n21001 );
buf ( n28051 , n27885 );
buf ( n28052 , n27888 );
buf ( n28053 , n28052 );
xor ( n28054 , n28051 , n28053 );
buf ( n28055 , n27897 );
buf ( n28056 , n28055 );
buf ( n28057 , n27932 );
nand ( n28058 , n28056 , n28057 );
not ( n28059 , n28058 );
nor ( n28060 , n28054 , n28059 );
not ( n28061 , n28060 );
nand ( n28062 , n28054 , n28059 );
nand ( n28063 , n28061 , n28062 );
not ( n28064 , n28063 );
buf ( n28065 , n27997 );
not ( n28066 , n28065 );
buf ( n28067 , n28000 );
not ( n28068 , n28067 );
not ( n28069 , n28068 );
or ( n28070 , n28066 , n28069 );
not ( n28071 , n28065 );
nand ( n28072 , n28071 , n28067 );
nand ( n28073 , n28070 , n28072 );
and ( n28074 , n26949 , n26947 );
nor ( n28075 , n28073 , n28074 );
nor ( n28076 , n28075 , n26959 );
not ( n28077 , n28076 );
nor ( n28078 , n28077 , n27014 );
nand ( n28079 , n26990 , n28078 );
not ( n28080 , n28057 );
not ( n28081 , n28056 );
not ( n28082 , n28081 );
or ( n28083 , n28080 , n28082 );
not ( n28084 , n28057 );
nand ( n28085 , n28084 , n28056 );
nand ( n28086 , n28083 , n28085 );
buf ( n28087 , n28065 );
and ( n28088 , n28067 , n28087 );
nor ( n28089 , n28086 , n28088 );
nor ( n28090 , n28079 , n28089 );
not ( n28091 , n28090 );
nand ( n28092 , n27019 , n24272 );
not ( n28093 , n28092 );
or ( n28094 , n28091 , n28093 );
not ( n28095 , n28089 );
not ( n28096 , n28095 );
or ( n28097 , n28075 , n26961 );
nand ( n28098 , n28073 , n28074 );
nand ( n28099 , n28097 , n28098 );
nor ( n28100 , n27039 , n28099 );
nand ( n28101 , n28100 , n27027 );
not ( n28102 , n28101 );
not ( n28103 , n27032 );
and ( n28104 , n28102 , n28103 );
not ( n28105 , n28100 );
or ( n28106 , n28105 , n27013 );
or ( n28107 , n28099 , n28076 );
nand ( n28108 , n28106 , n28107 );
nor ( n28109 , n28104 , n28108 );
not ( n28110 , n28109 );
or ( n28111 , n28096 , n28110 );
nand ( n28112 , n28086 , n28088 );
nand ( n28113 , n28111 , n28112 );
not ( n28114 , n28113 );
nand ( n28115 , n28094 , n28114 );
not ( n28116 , n28115 );
or ( n28117 , n28064 , n28116 );
or ( n28118 , n28115 , n28063 );
nand ( n28119 , n28117 , n28118 );
buf ( n28120 , n28119 );
nand ( n28121 , n28120 , n19358 );
buf ( n28122 , n27885 );
not ( n28123 , n28122 );
buf ( n28124 , n24313 );
nor ( n28125 , n27072 , n24304 );
buf ( n28126 , n27932 );
nor ( n28127 , n28126 , n27054 );
not ( n28128 , n27062 );
buf ( n28129 , n27997 );
buf ( n28130 , n28129 );
not ( n28131 , n28130 );
and ( n28132 , n28127 , n28128 , n28131 );
not ( n28133 , n27059 );
nand ( n28134 , n28125 , n28132 , n28133 , n24301 );
nor ( n28135 , n28124 , n28134 );
not ( n28136 , n28135 );
or ( n28137 , n28123 , n28136 );
or ( n28138 , n28135 , n28122 );
nand ( n28139 , n28137 , n28138 );
buf ( n28140 , n28139 );
and ( n28141 , n28140 , n19290 );
and ( n28142 , n27619 , n27885 );
nor ( n28143 , n28141 , n28142 );
nand ( n28144 , n28050 , n28121 , n28143 );
nor ( n28145 , n27846 , n28144 );
buf ( n28146 , n24450 );
or ( n28147 , n28145 , n28146 );
not ( n28148 , n18648 );
nand ( n28149 , n28148 , n24450 );
nand ( n28150 , n28147 , n28149 );
buf ( n28151 , n28150 );
buf ( n28152 , n28151 );
not ( n28153 , n275550 );
buf ( n28154 , n28153 );
buf ( n28155 , n28154 );
not ( n28156 , n22169 );
not ( n28157 , n22145 );
or ( n28158 , n28156 , n28157 );
or ( n28159 , n22145 , n22165 );
nand ( n28160 , n28158 , n28159 );
buf ( n28161 , n28160 );
buf ( n28162 , n28161 );
not ( n28163 , n275925 );
buf ( n28164 , n28163 );
buf ( n28165 , n28164 );
not ( n28166 , n275929 );
buf ( n28167 , n28166 );
buf ( n28168 , n28167 );
buf ( n28169 , n275554 );
buf ( n28170 , n275554 );
buf ( n28171 , n275554 );
not ( n28172 , n275929 );
buf ( n28173 , n28172 );
buf ( n28174 , n28173 );
not ( n28175 , n275550 );
buf ( n28176 , n28175 );
buf ( n28177 , n28176 );
buf ( n28178 , n275554 );
or ( n28179 , n23691 , n23695 );
and ( n28180 , n23701 , n23687 );
and ( n28181 , n22010 , n22145 , n12105 );
nor ( n28182 , n28180 , n28181 );
nand ( n28183 , n28179 , n28182 );
buf ( n28184 , n28183 );
not ( n28185 , n28184 );
nor ( n28186 , n28185 , n22056 );
nand ( n28187 , n22123 , n27196 );
buf ( n28188 , n27194 );
and ( n28189 , n28187 , n28188 );
not ( n28190 , n28187 );
not ( n28191 , n28188 );
and ( n28192 , n28190 , n28191 );
nor ( n28193 , n28189 , n28192 );
buf ( n28194 , n28193 );
nand ( n28195 , n28186 , n28194 );
and ( n28196 , n28184 , n22000 );
buf ( n28197 , n21928 );
buf ( n28198 , n21921 );
nand ( n28199 , n28197 , n28198 );
buf ( n28200 , n28199 );
buf ( n28201 , n28200 );
buf ( n28202 , n21909 );
buf ( n28203 , n28202 );
not ( n28204 , n28203 );
buf ( n28205 , n28204 );
buf ( n28206 , n28205 );
and ( n28207 , n28201 , n28206 );
not ( n28208 , n28201 );
buf ( n28209 , n28202 );
and ( n28210 , n28208 , n28209 );
nor ( n28211 , n28207 , n28210 );
buf ( n28212 , n28211 );
buf ( n28213 , n28212 );
nand ( n28214 , n28196 , n28213 );
and ( n28215 , n28195 , n28214 );
not ( n28216 , n28184 );
nor ( n28217 , n28216 , n22051 );
not ( n28218 , n28217 );
not ( n28219 , n28218 );
buf ( n28220 , n22019 );
nand ( n28221 , n22033 , n28220 );
buf ( n28222 , n28221 );
not ( n28223 , n22021 );
and ( n28224 , n28222 , n28223 );
not ( n28225 , n28222 );
and ( n28226 , n28225 , n22021 );
nor ( n28227 , n28224 , n28226 );
buf ( n28228 , n28227 );
nand ( n28229 , n28219 , n28228 );
nand ( n28230 , n28184 , n22007 );
not ( n28231 , n28230 );
and ( n28232 , n28231 , n12318 );
buf ( n28233 , n28184 );
not ( n28234 , n10990 );
or ( n28235 , n28233 , n28234 );
buf ( n28236 , n28181 );
nand ( n28237 , n28236 , n11006 );
nand ( n28238 , n28235 , n28237 );
nor ( n28239 , n28232 , n28238 );
nand ( n28240 , n28184 , n23679 );
buf ( n28241 , n28240 );
not ( n28242 , n28241 );
nand ( n28243 , n28242 , n12141 );
nand ( n28244 , n28215 , n28229 , n28239 , n28243 );
buf ( n28245 , n28244 );
buf ( n28246 , n28245 );
not ( n28247 , n20961 );
not ( n28248 , n28247 );
buf ( n28249 , n14525 );
not ( n28250 , n28249 );
or ( n28251 , n28248 , n28250 );
not ( n28252 , n28247 );
nand ( n28253 , n28252 , n9458 );
nand ( n28254 , n28251 , n28253 );
buf ( n28255 , n28254 );
buf ( n28256 , n28255 );
buf ( n28257 , n275554 );
buf ( n28258 , n27342 );
buf ( n28259 , n27443 );
nand ( n28260 , n28258 , n28259 );
buf ( n28261 , n28260 );
buf ( n28262 , n28261 );
not ( n28263 , n28262 );
buf ( n28264 , n27319 );
not ( n28265 , n28264 );
buf ( n28266 , n28265 );
buf ( n28267 , n28266 );
buf ( n28268 , n27354 );
buf ( n28269 , n28268 );
not ( n28270 , n28269 );
buf ( n28271 , n28270 );
buf ( n28272 , n28271 );
nor ( n28273 , n28267 , n28272 );
buf ( n28274 , n28273 );
buf ( n28275 , n28274 );
not ( n28276 , n28275 );
buf ( n28277 , n23568 );
not ( n28278 , n28277 );
or ( n28279 , n28276 , n28278 );
buf ( n28280 , n27416 );
buf ( n28281 , n27398 );
nand ( n28282 , n28280 , n28281 );
buf ( n28283 , n28282 );
buf ( n28284 , n28283 );
not ( n28285 , n28284 );
buf ( n28286 , n28271 );
not ( n28287 , n28286 );
and ( n28288 , n28285 , n28287 );
buf ( n28289 , n27434 );
nor ( n28290 , n28288 , n28289 );
buf ( n28291 , n28290 );
buf ( n28292 , n28291 );
nand ( n28293 , n28279 , n28292 );
buf ( n28294 , n28293 );
buf ( n28295 , n28294 );
not ( n28296 , n28295 );
or ( n28297 , n28263 , n28296 );
buf ( n28298 , n28294 );
buf ( n28299 , n28261 );
or ( n28300 , n28298 , n28299 );
nand ( n28301 , n28297 , n28300 );
buf ( n28302 , n28301 );
buf ( n28303 , n28302 );
nand ( n28304 , n28233 , n22000 );
buf ( n28305 , n28304 );
not ( n28306 , n28305 );
nand ( n28307 , n28303 , n28306 );
nand ( n28308 , n27215 , n27248 );
not ( n28309 , n28308 );
buf ( n28310 , n27219 );
not ( n28311 , n28310 );
not ( n28312 , n27210 );
nor ( n28313 , n28311 , n28312 );
not ( n28314 , n28313 );
not ( n28315 , n23638 );
or ( n28316 , n28314 , n28315 );
nand ( n28317 , n27237 , n27239 );
not ( n28318 , n28317 );
and ( n28319 , n28318 , n28310 );
nor ( n28320 , n28319 , n27242 );
nand ( n28321 , n28316 , n28320 );
not ( n28322 , n28321 );
or ( n28323 , n28309 , n28322 );
or ( n28324 , n28321 , n28308 );
nand ( n28325 , n28323 , n28324 );
buf ( n28326 , n28325 );
not ( n28327 , n28184 );
nor ( n28328 , n28327 , n22056 );
not ( n28329 , n28328 );
not ( n28330 , n28329 );
nand ( n28331 , n28326 , n28330 );
not ( n28332 , n28218 );
not ( n28333 , n27509 );
not ( n28334 , n28333 );
not ( n28335 , n23658 );
nor ( n28336 , n23665 , n28335 );
buf ( n28337 , n27496 );
nand ( n28338 , n28336 , n28337 );
buf ( n28339 , n27499 );
not ( n28340 , n28339 );
nor ( n28341 , n28338 , n28340 );
not ( n28342 , n28341 );
or ( n28343 , n28334 , n28342 );
not ( n28344 , n28333 );
not ( n28345 , n28344 );
or ( n28346 , n28341 , n28345 );
nand ( n28347 , n28343 , n28346 );
buf ( n28348 , n28347 );
and ( n28349 , n28332 , n28348 );
not ( n28350 , n28241 );
and ( n28351 , n28350 , n12353 );
nor ( n28352 , n28349 , n28351 );
and ( n28353 , n28231 , n12219 );
buf ( n28354 , n28233 );
or ( n28355 , n28354 , n11410 );
not ( n28356 , n28236 );
not ( n28357 , n28356 );
nand ( n28358 , n28357 , n11404 );
nand ( n28359 , n28355 , n28358 );
nor ( n28360 , n28353 , n28359 );
nand ( n28361 , n28307 , n28331 , n28352 , n28360 );
buf ( n28362 , n28361 );
buf ( n28363 , n28362 );
buf ( n28364 , n275554 );
buf ( n28365 , n275554 );
buf ( n28366 , n27434 );
not ( n28367 , n28366 );
buf ( n28368 , n28268 );
nand ( n28369 , n28367 , n28368 );
buf ( n28370 , n28369 );
buf ( n28371 , n28370 );
not ( n28372 , n28371 );
buf ( n28373 , n28266 );
not ( n28374 , n28373 );
buf ( n28375 , n28374 );
buf ( n28376 , n28375 );
not ( n28377 , n28376 );
buf ( n28378 , n23568 );
not ( n28379 , n28378 );
or ( n28380 , n28377 , n28379 );
buf ( n28381 , n28283 );
not ( n28382 , n28381 );
buf ( n28383 , n28382 );
buf ( n28384 , n28383 );
not ( n28385 , n28384 );
buf ( n28386 , n28385 );
buf ( n28387 , n28386 );
nand ( n28388 , n28380 , n28387 );
buf ( n28389 , n28388 );
buf ( n28390 , n28389 );
not ( n28391 , n28390 );
or ( n28392 , n28372 , n28391 );
buf ( n28393 , n28389 );
buf ( n28394 , n28370 );
or ( n28395 , n28393 , n28394 );
nand ( n28396 , n28392 , n28395 );
buf ( n28397 , n28396 );
buf ( n28398 , n28397 );
not ( n28399 , n22189 );
not ( n28400 , n11741 );
not ( n28401 , n12111 );
or ( n28402 , n28400 , n28401 );
nand ( n28403 , n28402 , n22182 );
not ( n28404 , n28403 );
or ( n28405 , n28399 , n28404 );
nand ( n28406 , n23690 , n22172 );
nand ( n28407 , n28405 , n28406 );
buf ( n28408 , n28407 );
nand ( n28409 , n28398 , n28408 );
not ( n28410 , n27242 );
nand ( n28411 , n28410 , n28310 );
not ( n28412 , n28411 );
not ( n28413 , n28312 );
not ( n28414 , n28413 );
not ( n28415 , n23634 );
nand ( n28416 , n22129 , n23636 );
nand ( n28417 , n28415 , n28416 );
not ( n28418 , n28417 );
or ( n28419 , n28414 , n28418 );
not ( n28420 , n28318 );
nand ( n28421 , n28419 , n28420 );
not ( n28422 , n28421 );
or ( n28423 , n28412 , n28422 );
or ( n28424 , n28421 , n28411 );
nand ( n28425 , n28423 , n28424 );
buf ( n28426 , n28425 );
nor ( n28427 , n22055 , n22188 );
buf ( n28428 , n28427 );
not ( n28429 , n28428 );
not ( n28430 , n28429 );
nand ( n28431 , n28426 , n28430 );
xnor ( n28432 , n28338 , n28339 );
buf ( n28433 , n28432 );
nand ( n28434 , n22005 , n22172 );
not ( n28435 , n28434 );
not ( n28436 , n22004 );
nand ( n28437 , n28435 , n28436 );
not ( n28438 , n28437 );
not ( n28439 , n28438 );
not ( n28440 , n28439 );
nand ( n28441 , n28433 , n28440 );
not ( n28442 , n22055 );
or ( n28443 , n28403 , n28442 );
nand ( n28444 , n28443 , n22189 );
nand ( n28445 , n12380 , n22172 );
not ( n28446 , n22011 );
not ( n28447 , n22188 );
and ( n28448 , n28446 , n28447 );
nor ( n28449 , n28448 , n28181 );
nand ( n28450 , n28444 , n28445 , n28449 , n9159 );
not ( n28451 , n28450 );
nand ( n28452 , n28451 , n11392 );
nor ( n28453 , n28434 , n28436 );
not ( n28454 , n28453 );
not ( n28455 , n28454 );
buf ( n28456 , n12239 );
and ( n28457 , n28455 , n28456 );
not ( n28458 , n28449 );
not ( n28459 , n28458 );
or ( n28460 , n28459 , n12221 );
nand ( n28461 , n20649 , n9298 );
nand ( n28462 , n28460 , n28461 );
nor ( n28463 , n28457 , n28462 );
and ( n28464 , n28441 , n28452 , n28463 );
nand ( n28465 , n28409 , n28431 , n28464 );
buf ( n28466 , n28465 );
buf ( n28467 , n28466 );
not ( n28468 , n275550 );
buf ( n28469 , n28468 );
buf ( n28470 , n28469 );
buf ( n28471 , n275554 );
not ( n28472 , n275925 );
buf ( n28473 , n28472 );
buf ( n28474 , n28473 );
nand ( n28475 , n25063 , n19182 );
buf ( n28476 , n19182 );
buf ( n28477 , n28476 );
buf ( n28478 , n28477 );
not ( n28479 , n28478 );
buf ( n28480 , n18596 );
buf ( n28481 , n28480 );
not ( n28482 , n28481 );
and ( n28483 , n28479 , n28482 );
buf ( n28484 , n28477 );
buf ( n28485 , n28480 );
and ( n28486 , n28484 , n28485 );
nor ( n28487 , n28483 , n28486 );
buf ( n28488 , n28487 );
buf ( n28489 , n28488 );
not ( n28490 , n28489 );
buf ( n28491 , n25258 );
buf ( n28492 , n25242 );
nor ( n28493 , n28491 , n28492 );
buf ( n28494 , n28493 );
buf ( n28495 , n28494 );
buf ( n28496 , n25224 );
not ( n28497 , n28496 );
buf ( n28498 , n28497 );
buf ( n28499 , n28498 );
and ( n28500 , n28495 , n28499 );
buf ( n28501 , n25258 );
buf ( n28502 , n25151 );
or ( n28503 , n28501 , n28502 );
buf ( n28504 , n25106 );
buf ( n28505 , n25128 );
nand ( n28506 , n28503 , n28504 , n28505 );
buf ( n28507 , n28506 );
buf ( n28508 , n28507 );
nor ( n28509 , n28500 , n28508 );
buf ( n28510 , n28509 );
buf ( n28511 , n28510 );
buf ( n28512 , n25340 );
or ( n28513 , n28511 , n28512 );
buf ( n28514 , n28513 );
buf ( n28515 , n28514 );
buf ( n28516 , n25080 );
buf ( n28517 , n25294 );
nor ( n28518 , n28516 , n28517 );
buf ( n28519 , n28518 );
buf ( n28520 , n28519 );
buf ( n28521 , n25285 );
and ( n28522 , n28520 , n28521 );
buf ( n28523 , n28522 );
buf ( n28524 , n28523 );
buf ( n28525 , n17720 );
not ( n28526 , n28525 );
not ( n28527 , n28526 );
buf ( n28528 , n28527 );
buf ( n28529 , n28528 );
buf ( n28530 , n18945 );
buf ( n28531 , n28530 );
nor ( n28532 , n28529 , n28531 );
buf ( n28533 , n28532 );
buf ( n28534 , n28533 );
buf ( n28535 , n17734 );
not ( n28536 , n28535 );
not ( n28537 , n28536 );
buf ( n28538 , n28537 );
buf ( n28539 , n28538 );
buf ( n28540 , n18968 );
buf ( n28541 , n28540 );
nor ( n28542 , n28539 , n28541 );
buf ( n28543 , n28542 );
buf ( n28544 , n28543 );
or ( n28545 , n28534 , n28544 );
buf ( n28546 , n28545 );
buf ( n28547 , n28546 );
buf ( n28548 , n17704 );
not ( n28549 , n28548 );
not ( n28550 , n28549 );
buf ( n28551 , n28550 );
buf ( n28552 , n28551 );
buf ( n28553 , n18625 );
buf ( n28554 , n28553 );
nor ( n28555 , n28552 , n28554 );
buf ( n28556 , n28555 );
buf ( n28557 , n28556 );
nor ( n28558 , n28547 , n28557 );
buf ( n28559 , n28558 );
buf ( n28560 , n28559 );
and ( n28561 , n28515 , n28524 , n28560 );
buf ( n28562 , n28519 );
buf ( n28563 , n25357 );
and ( n28564 , n28562 , n28563 );
buf ( n28565 , n25080 );
buf ( n28566 , n25364 );
or ( n28567 , n28565 , n28566 );
buf ( n28568 , n25074 );
nand ( n28569 , n28567 , n28568 );
buf ( n28570 , n28569 );
buf ( n28571 , n28570 );
nor ( n28572 , n28564 , n28571 );
buf ( n28573 , n28572 );
buf ( n28574 , n28573 );
buf ( n28575 , n28559 );
not ( n28576 , n28575 );
buf ( n28577 , n28576 );
buf ( n28578 , n28577 );
or ( n28579 , n28574 , n28578 );
buf ( n28580 , n28556 );
buf ( n28581 , n28533 );
not ( n28582 , n28581 );
buf ( n28583 , n28538 );
buf ( n28584 , n28540 );
nand ( n28585 , n28583 , n28584 );
buf ( n28586 , n28585 );
buf ( n28587 , n28586 );
not ( n28588 , n28587 );
and ( n28589 , n28582 , n28588 );
buf ( n28590 , n28528 );
buf ( n28591 , n28530 );
and ( n28592 , n28590 , n28591 );
buf ( n28593 , n28592 );
buf ( n28594 , n28593 );
nor ( n28595 , n28589 , n28594 );
buf ( n28596 , n28595 );
buf ( n28597 , n28596 );
or ( n28598 , n28580 , n28597 );
buf ( n28599 , n28551 );
buf ( n28600 , n28553 );
nand ( n28601 , n28599 , n28600 );
buf ( n28602 , n28601 );
buf ( n28603 , n28602 );
nand ( n28604 , n28579 , n28598 , n28603 );
buf ( n28605 , n28604 );
buf ( n28606 , n28605 );
nor ( n28607 , n28561 , n28606 );
buf ( n28608 , n28607 );
buf ( n28609 , n28608 );
not ( n28610 , n28609 );
or ( n28611 , n28490 , n28610 );
buf ( n28612 , n28608 );
buf ( n28613 , n28488 );
or ( n28614 , n28612 , n28613 );
nand ( n28615 , n28611 , n28614 );
buf ( n28616 , n28615 );
buf ( n28617 , n28616 );
not ( n28618 , n28617 );
nor ( n28619 , n28618 , n25389 );
nand ( n28620 , n25396 , n9416 );
buf ( n28621 , n28476 );
buf ( n28622 , n28621 );
not ( n28623 , n28622 );
buf ( n28624 , n18600 );
buf ( n28625 , n28624 );
not ( n28626 , n28625 );
and ( n28627 , n28623 , n28626 );
buf ( n28628 , n28621 );
buf ( n28629 , n28624 );
and ( n28630 , n28628 , n28629 );
nor ( n28631 , n28627 , n28630 );
buf ( n28632 , n28631 );
buf ( n28633 , n28632 );
not ( n28634 , n28633 );
buf ( n28635 , n25563 );
buf ( n28636 , n25580 );
nor ( n28637 , n28635 , n28636 );
buf ( n28638 , n28637 );
buf ( n28639 , n28638 );
buf ( n28640 , n25543 );
and ( n28641 , n28639 , n28640 );
buf ( n28642 , n25580 );
buf ( n28643 , n25475 );
or ( n28644 , n28642 , n28643 );
buf ( n28645 , n25435 );
buf ( n28646 , n25453 );
nand ( n28647 , n28644 , n28645 , n28646 );
buf ( n28648 , n28647 );
buf ( n28649 , n28648 );
nor ( n28650 , n28641 , n28649 );
buf ( n28651 , n28650 );
buf ( n28652 , n28651 );
buf ( n28653 , n25666 );
or ( n28654 , n28652 , n28653 );
buf ( n28655 , n28654 );
buf ( n28656 , n28655 );
buf ( n28657 , n25414 );
buf ( n28658 , n25615 );
nor ( n28659 , n28657 , n28658 );
buf ( n28660 , n28659 );
buf ( n28661 , n28660 );
buf ( n28662 , n25606 );
nand ( n28663 , n28661 , n28662 );
buf ( n28664 , n28663 );
buf ( n28665 , n28664 );
not ( n28666 , n28665 );
buf ( n28667 , n28666 );
buf ( n28668 , n28667 );
buf ( n28669 , n28548 );
buf ( n28670 , n28669 );
buf ( n28671 , n28670 );
buf ( n28672 , n18620 );
buf ( n28673 , n28672 );
nor ( n28674 , n28671 , n28673 );
buf ( n28675 , n28674 );
buf ( n28676 , n28675 );
not ( n28677 , n28676 );
not ( n28678 , n28526 );
buf ( n28679 , n28678 );
buf ( n28680 , n28679 );
buf ( n28681 , n18940 );
buf ( n28682 , n28681 );
nor ( n28683 , n28680 , n28682 );
buf ( n28684 , n28683 );
buf ( n28685 , n28684 );
buf ( n28686 , n28535 );
buf ( n28687 , n28686 );
buf ( n28688 , n18963 );
buf ( n28689 , n28688 );
nor ( n28690 , n28687 , n28689 );
buf ( n28691 , n28690 );
buf ( n28692 , n28691 );
nor ( n28693 , n28685 , n28692 );
buf ( n28694 , n28693 );
buf ( n28695 , n28694 );
nand ( n28696 , n28677 , n28695 );
buf ( n28697 , n28696 );
buf ( n28698 , n28697 );
not ( n28699 , n28698 );
buf ( n28700 , n28699 );
buf ( n28701 , n28700 );
and ( n28702 , n28656 , n28668 , n28701 );
buf ( n28703 , n28660 );
buf ( n28704 , n25683 );
and ( n28705 , n28703 , n28704 );
buf ( n28706 , n25414 );
buf ( n28707 , n25690 );
or ( n28708 , n28706 , n28707 );
buf ( n28709 , n25408 );
nand ( n28710 , n28708 , n28709 );
buf ( n28711 , n28710 );
buf ( n28712 , n28711 );
nor ( n28713 , n28705 , n28712 );
buf ( n28714 , n28713 );
buf ( n28715 , n28714 );
buf ( n28716 , n28697 );
or ( n28717 , n28715 , n28716 );
buf ( n28718 , n28675 );
buf ( n28719 , n28684 );
buf ( n28720 , n28686 );
buf ( n28721 , n28688 );
nand ( n28722 , n28720 , n28721 );
buf ( n28723 , n28722 );
buf ( n28724 , n28723 );
or ( n28725 , n28719 , n28724 );
buf ( n28726 , n28679 );
buf ( n28727 , n28681 );
nand ( n28728 , n28726 , n28727 );
buf ( n28729 , n28728 );
buf ( n28730 , n28729 );
nand ( n28731 , n28725 , n28730 );
buf ( n28732 , n28731 );
buf ( n28733 , n28732 );
not ( n28734 , n28733 );
buf ( n28735 , n28734 );
buf ( n28736 , n28735 );
or ( n28737 , n28718 , n28736 );
buf ( n28738 , n28670 );
buf ( n28739 , n28672 );
nand ( n28740 , n28738 , n28739 );
buf ( n28741 , n28740 );
buf ( n28742 , n28741 );
nand ( n28743 , n28717 , n28737 , n28742 );
buf ( n28744 , n28743 );
buf ( n28745 , n28744 );
nor ( n28746 , n28702 , n28745 );
buf ( n28747 , n28746 );
buf ( n28748 , n28747 );
not ( n28749 , n28748 );
or ( n28750 , n28634 , n28749 );
buf ( n28751 , n28747 );
buf ( n28752 , n28632 );
or ( n28753 , n28751 , n28752 );
nand ( n28754 , n28750 , n28753 );
buf ( n28755 , n28754 );
buf ( n28756 , n28755 );
and ( n28757 , n25402 , n28756 );
not ( n28758 , n18591 );
nor ( n28759 , n19639 , n28758 );
nor ( n28760 , n28757 , n28759 );
not ( n28761 , n25716 );
buf ( n28762 , n28476 );
buf ( n28763 , n28762 );
not ( n28764 , n28763 );
buf ( n28765 , n18596 );
buf ( n28766 , n28765 );
not ( n28767 , n28766 );
and ( n28768 , n28764 , n28767 );
buf ( n28769 , n28762 );
buf ( n28770 , n28765 );
and ( n28771 , n28769 , n28770 );
nor ( n28772 , n28768 , n28771 );
buf ( n28773 , n28772 );
buf ( n28774 , n28773 );
not ( n28775 , n28774 );
buf ( n28776 , n25879 );
buf ( n28777 , n25896 );
nor ( n28778 , n28776 , n28777 );
buf ( n28779 , n28778 );
buf ( n28780 , n28779 );
buf ( n28781 , n25859 );
and ( n28782 , n28780 , n28781 );
buf ( n28783 , n25896 );
buf ( n28784 , n25792 );
or ( n28785 , n28783 , n28784 );
buf ( n28786 , n25751 );
buf ( n28787 , n25770 );
nand ( n28788 , n28785 , n28786 , n28787 );
buf ( n28789 , n28788 );
buf ( n28790 , n28789 );
nor ( n28791 , n28782 , n28790 );
buf ( n28792 , n28791 );
buf ( n28793 , n28792 );
buf ( n28794 , n25977 );
or ( n28795 , n28793 , n28794 );
buf ( n28796 , n28795 );
buf ( n28797 , n28796 );
buf ( n28798 , n25730 );
buf ( n28799 , n25928 );
nor ( n28800 , n28798 , n28799 );
buf ( n28801 , n28800 );
buf ( n28802 , n28801 );
buf ( n28803 , n25920 );
nand ( n28804 , n28802 , n28803 );
buf ( n28805 , n28804 );
buf ( n28806 , n28805 );
not ( n28807 , n28806 );
buf ( n28808 , n28807 );
buf ( n28809 , n28808 );
buf ( n28810 , n28669 );
buf ( n28811 , n28810 );
buf ( n28812 , n18625 );
buf ( n28813 , n28812 );
nor ( n28814 , n28811 , n28813 );
buf ( n28815 , n28814 );
buf ( n28816 , n28815 );
not ( n28817 , n28816 );
buf ( n28818 , n28525 );
buf ( n28819 , n28818 );
buf ( n28820 , n28819 );
buf ( n28821 , n18945 );
buf ( n28822 , n28821 );
nor ( n28823 , n28820 , n28822 );
buf ( n28824 , n28823 );
buf ( n28825 , n28824 );
not ( n28826 , n28536 );
buf ( n28827 , n28826 );
buf ( n28828 , n28827 );
buf ( n28829 , n18968 );
buf ( n28830 , n28829 );
nor ( n28831 , n28828 , n28830 );
buf ( n28832 , n28831 );
buf ( n28833 , n28832 );
nor ( n28834 , n28825 , n28833 );
buf ( n28835 , n28834 );
buf ( n28836 , n28835 );
nand ( n28837 , n28817 , n28836 );
buf ( n28838 , n28837 );
buf ( n28839 , n28838 );
not ( n28840 , n28839 );
buf ( n28841 , n28840 );
buf ( n28842 , n28841 );
and ( n28843 , n28797 , n28809 , n28842 );
buf ( n28844 , n28801 );
buf ( n28845 , n25994 );
and ( n28846 , n28844 , n28845 );
buf ( n28847 , n25730 );
buf ( n28848 , n26001 );
or ( n28849 , n28847 , n28848 );
buf ( n28850 , n25724 );
nand ( n28851 , n28849 , n28850 );
buf ( n28852 , n28851 );
buf ( n28853 , n28852 );
nor ( n28854 , n28846 , n28853 );
buf ( n28855 , n28854 );
buf ( n28856 , n28855 );
buf ( n28857 , n28838 );
or ( n28858 , n28856 , n28857 );
buf ( n28859 , n28815 );
buf ( n28860 , n28824 );
buf ( n28861 , n28827 );
buf ( n28862 , n28829 );
nand ( n28863 , n28861 , n28862 );
buf ( n28864 , n28863 );
buf ( n28865 , n28864 );
or ( n28866 , n28860 , n28865 );
buf ( n28867 , n28819 );
buf ( n28868 , n28821 );
nand ( n28869 , n28867 , n28868 );
buf ( n28870 , n28869 );
buf ( n28871 , n28870 );
nand ( n28872 , n28866 , n28871 );
buf ( n28873 , n28872 );
buf ( n28874 , n28873 );
not ( n28875 , n28874 );
buf ( n28876 , n28875 );
buf ( n28877 , n28876 );
or ( n28878 , n28859 , n28877 );
buf ( n28879 , n28810 );
buf ( n28880 , n28812 );
nand ( n28881 , n28879 , n28880 );
buf ( n28882 , n28881 );
buf ( n28883 , n28882 );
nand ( n28884 , n28858 , n28878 , n28883 );
buf ( n28885 , n28884 );
buf ( n28886 , n28885 );
nor ( n28887 , n28843 , n28886 );
buf ( n28888 , n28887 );
buf ( n28889 , n28888 );
not ( n28890 , n28889 );
or ( n28891 , n28775 , n28890 );
buf ( n28892 , n28888 );
buf ( n28893 , n28773 );
or ( n28894 , n28892 , n28893 );
nand ( n28895 , n28891 , n28894 );
buf ( n28896 , n28895 );
buf ( n28897 , n28896 );
nand ( n28898 , n28761 , n28897 );
nand ( n28899 , n28620 , n28760 , n28898 );
nor ( n28900 , n28619 , n28899 );
buf ( n28901 , n28476 );
buf ( n28902 , n28901 );
not ( n28903 , n28902 );
buf ( n28904 , n18600 );
buf ( n28905 , n28904 );
not ( n28906 , n28905 );
and ( n28907 , n28903 , n28906 );
buf ( n28908 , n28901 );
buf ( n28909 , n28904 );
and ( n28910 , n28908 , n28909 );
nor ( n28911 , n28907 , n28910 );
buf ( n28912 , n28911 );
buf ( n28913 , n28912 );
not ( n28914 , n28913 );
buf ( n28915 , n26206 );
buf ( n28916 , n26189 );
nor ( n28917 , n28915 , n28916 );
buf ( n28918 , n28917 );
buf ( n28919 , n28918 );
buf ( n28920 , n26169 );
and ( n28921 , n28919 , n28920 );
buf ( n28922 , n26206 );
buf ( n28923 , n26100 );
or ( n28924 , n28922 , n28923 );
buf ( n28925 , n26061 );
buf ( n28926 , n26078 );
nand ( n28927 , n28924 , n28925 , n28926 );
buf ( n28928 , n28927 );
buf ( n28929 , n28928 );
nor ( n28930 , n28921 , n28929 );
buf ( n28931 , n28930 );
buf ( n28932 , n28931 );
buf ( n28933 , n26281 );
or ( n28934 , n28932 , n28933 );
buf ( n28935 , n28934 );
buf ( n28936 , n28935 );
buf ( n28937 , n26039 );
buf ( n28938 , n26238 );
nor ( n28939 , n28937 , n28938 );
buf ( n28940 , n28939 );
buf ( n28941 , n28940 );
buf ( n28942 , n26229 );
nand ( n28943 , n28941 , n28942 );
buf ( n28944 , n28943 );
buf ( n28945 , n28944 );
not ( n28946 , n28945 );
buf ( n28947 , n28946 );
buf ( n28948 , n28947 );
buf ( n28949 , n28527 );
buf ( n28950 , n28949 );
buf ( n28951 , n28950 );
buf ( n28952 , n18940 );
buf ( n28953 , n28952 );
nor ( n28954 , n28951 , n28953 );
buf ( n28955 , n28954 );
buf ( n28956 , n28955 );
not ( n28957 , n28536 );
buf ( n28958 , n28957 );
buf ( n28959 , n28958 );
buf ( n28960 , n28959 );
buf ( n28961 , n18963 );
buf ( n28962 , n28961 );
nor ( n28963 , n28960 , n28962 );
buf ( n28964 , n28963 );
buf ( n28965 , n28964 );
or ( n28966 , n28956 , n28965 );
buf ( n28967 , n28966 );
buf ( n28968 , n28967 );
buf ( n28969 , n28550 );
buf ( n28970 , n28969 );
buf ( n28971 , n28970 );
buf ( n28972 , n18620 );
buf ( n28973 , n28972 );
nor ( n28974 , n28971 , n28973 );
buf ( n28975 , n28974 );
buf ( n28976 , n28975 );
nor ( n28977 , n28968 , n28976 );
buf ( n28978 , n28977 );
buf ( n28979 , n28978 );
and ( n28980 , n28936 , n28948 , n28979 );
buf ( n28981 , n28940 );
buf ( n28982 , n26298 );
and ( n28983 , n28981 , n28982 );
buf ( n28984 , n26039 );
buf ( n28985 , n26305 );
or ( n28986 , n28984 , n28985 );
buf ( n28987 , n26033 );
nand ( n28988 , n28986 , n28987 );
buf ( n28989 , n28988 );
buf ( n28990 , n28989 );
nor ( n28991 , n28983 , n28990 );
buf ( n28992 , n28991 );
buf ( n28993 , n28992 );
buf ( n28994 , n28978 );
not ( n28995 , n28994 );
buf ( n28996 , n28995 );
buf ( n28997 , n28996 );
or ( n28998 , n28993 , n28997 );
buf ( n28999 , n28975 );
buf ( n29000 , n28955 );
not ( n29001 , n29000 );
buf ( n29002 , n28959 );
buf ( n29003 , n28961 );
nand ( n29004 , n29002 , n29003 );
buf ( n29005 , n29004 );
buf ( n29006 , n29005 );
not ( n29007 , n29006 );
and ( n29008 , n29001 , n29007 );
buf ( n29009 , n28950 );
buf ( n29010 , n28952 );
and ( n29011 , n29009 , n29010 );
buf ( n29012 , n29011 );
buf ( n29013 , n29012 );
nor ( n29014 , n29008 , n29013 );
buf ( n29015 , n29014 );
buf ( n29016 , n29015 );
or ( n29017 , n28999 , n29016 );
buf ( n29018 , n28970 );
buf ( n29019 , n28972 );
nand ( n29020 , n29018 , n29019 );
buf ( n29021 , n29020 );
buf ( n29022 , n29021 );
nand ( n29023 , n28998 , n29017 , n29022 );
buf ( n29024 , n29023 );
buf ( n29025 , n29024 );
nor ( n29026 , n28980 , n29025 );
buf ( n29027 , n29026 );
buf ( n29028 , n29027 );
not ( n29029 , n29028 );
or ( n29030 , n28914 , n29029 );
buf ( n29031 , n29027 );
buf ( n29032 , n28912 );
or ( n29033 , n29031 , n29032 );
nand ( n29034 , n29030 , n29033 );
buf ( n29035 , n29034 );
buf ( n29036 , n29035 );
nand ( n29037 , n26027 , n29036 );
nand ( n29038 , n28475 , n28900 , n29037 );
buf ( n29039 , n29038 );
buf ( n29040 , n29039 );
buf ( n29041 , n275554 );
buf ( n29042 , n14425 );
not ( n29043 , n29042 );
not ( n29044 , n28247 );
or ( n29045 , n29043 , n29044 );
buf ( n29046 , n28252 );
nand ( n29047 , n29046 , n9710 );
nand ( n29048 , n29045 , n29047 );
buf ( n29049 , n29048 );
buf ( n29050 , n29049 );
not ( n29051 , n275550 );
buf ( n29052 , n29051 );
buf ( n29053 , n29052 );
not ( n29054 , n275550 );
buf ( n29055 , n29054 );
buf ( n29056 , n29055 );
buf ( n29057 , n14153 );
not ( n29058 , n29057 );
or ( n29059 , n29058 , n29046 );
nand ( n29060 , n28252 , n9558 );
nand ( n29061 , n29059 , n29060 );
buf ( n29062 , n29061 );
buf ( n29063 , n29062 );
not ( n29064 , n275925 );
buf ( n29065 , n29064 );
buf ( n29066 , n29065 );
or ( n29067 , n19629 , n19216 );
and ( n29068 , n20514 , n19360 );
not ( n29069 , n19317 );
not ( n29070 , n19665 );
and ( n29071 , n29069 , n29070 );
and ( n29072 , n19221 , n20566 );
nor ( n29073 , n29071 , n29072 );
nor ( n29074 , n19176 , n19289 );
buf ( n29075 , n29074 );
nand ( n29076 , n20558 , n29075 );
nand ( n29077 , n19387 , n18760 );
nand ( n29078 , n29073 , n29076 , n29077 );
nor ( n29079 , n29068 , n29078 );
nand ( n29080 , n20352 , n19354 );
and ( n29081 , n29079 , n29080 );
nand ( n29082 , n29067 , n29081 );
buf ( n29083 , n29082 );
buf ( n29084 , n29083 );
buf ( n29085 , n275554 );
buf ( n29086 , n275554 );
not ( n29087 , n275929 );
buf ( n29088 , n29087 );
buf ( n29089 , n29088 );
not ( n29090 , n275550 );
buf ( n29091 , n29090 );
buf ( n29092 , n29091 );
not ( n29093 , n275550 );
buf ( n29094 , n29093 );
buf ( n29095 , n29094 );
buf ( n29096 , n275554 );
not ( n29097 , n275929 );
buf ( n29098 , n29097 );
buf ( n29099 , n29098 );
not ( n29100 , n275929 );
buf ( n29101 , n29100 );
buf ( n29102 , n29101 );
buf ( n29103 , n275554 );
not ( n29104 , n16642 );
or ( n29105 , n29104 , n14830 );
nand ( n29106 , n22915 , n23807 );
nand ( n29107 , n29105 , n29106 );
buf ( n29108 , n29107 );
buf ( n29109 , n29108 );
buf ( n29110 , n23951 );
not ( n29111 , n29110 );
or ( n29112 , n29111 , n21770 );
nand ( n29113 , n21774 , n9714 );
nand ( n29114 , n29112 , n29113 );
buf ( n29115 , n29114 );
buf ( n29116 , n29115 );
not ( n29117 , n22089 );
nand ( n29118 , n27202 , n29117 );
not ( n29119 , n29118 );
buf ( n29120 , n22074 );
nand ( n29121 , n29120 , n22094 );
not ( n29122 , n29121 );
or ( n29123 , n29119 , n29122 );
or ( n29124 , n29118 , n29121 );
nand ( n29125 , n29123 , n29124 );
buf ( n29126 , n29125 );
and ( n29127 , n29126 , n22057 );
not ( n29128 , n12264 );
not ( n29129 , n22007 );
or ( n29130 , n29128 , n29129 );
nand ( n29131 , n22013 , n10740 );
nand ( n29132 , n29130 , n29131 );
nor ( n29133 , n29127 , n29132 );
and ( n29134 , n22038 , n22041 );
not ( n29135 , n22038 );
and ( n29136 , n29135 , n22040 );
nor ( n29137 , n29134 , n29136 );
buf ( n29138 , n29137 );
nand ( n29139 , n29138 , n22052 );
buf ( n29140 , n21842 );
not ( n29141 , n29140 );
buf ( n29142 , n27296 );
nand ( n29143 , n29141 , n29142 );
buf ( n29144 , n29143 );
buf ( n29145 , n29144 );
buf ( n29146 , n21805 );
buf ( n29147 , n21852 );
nand ( n29148 , n29146 , n29147 );
buf ( n29149 , n29148 );
buf ( n29150 , n29149 );
xnor ( n29151 , n29145 , n29150 );
buf ( n29152 , n29151 );
buf ( n29153 , n29152 );
nand ( n29154 , n29153 , n22002 );
nand ( n29155 , n29133 , n29139 , n29154 );
not ( n29156 , n29155 );
or ( n29157 , n29156 , n23708 );
nand ( n29158 , n27641 , n10765 );
nand ( n29159 , n29157 , n29158 );
buf ( n29160 , n29159 );
buf ( n29161 , n29160 );
buf ( n29162 , n28437 );
not ( n29163 , n29162 );
nand ( n29164 , n27576 , n29163 );
and ( n29165 , n27561 , n28408 );
and ( n29166 , n27586 , n28428 );
nor ( n29167 , n29165 , n29166 );
not ( n29168 , n28450 );
not ( n29169 , n10888 );
nand ( n29170 , n29168 , n29169 );
buf ( n29171 , n28453 );
not ( n29172 , n29171 );
not ( n29173 , n29172 );
not ( n29174 , n12190 );
and ( n29175 , n29173 , n29174 );
or ( n29176 , n28459 , n12234 );
nand ( n29177 , n20649 , n9285 );
nand ( n29178 , n29176 , n29177 );
nor ( n29179 , n29175 , n29178 );
nand ( n29180 , n29164 , n29167 , n29170 , n29179 );
buf ( n29181 , n29180 );
buf ( n29182 , n29181 );
not ( n29183 , n275929 );
buf ( n29184 , n29183 );
buf ( n29185 , n29184 );
not ( n29186 , n275929 );
buf ( n29187 , n29186 );
buf ( n29188 , n29187 );
buf ( n29189 , n21931 );
buf ( n29190 , n29189 );
not ( n29191 , n29190 );
buf ( n29192 , n21899 );
buf ( n29193 , n21882 );
buf ( n29194 , n29193 );
nand ( n29195 , n29192 , n29194 );
buf ( n29196 , n29195 );
buf ( n29197 , n29196 );
not ( n29198 , n29197 );
or ( n29199 , n29191 , n29198 );
buf ( n29200 , n29196 );
buf ( n29201 , n29189 );
or ( n29202 , n29200 , n29201 );
nand ( n29203 , n29199 , n29202 );
buf ( n29204 , n29203 );
buf ( n29205 , n29204 );
nand ( n29206 , n29205 , n28407 );
buf ( n29207 , n22124 );
not ( n29208 , n29207 );
not ( n29209 , n22102 );
nand ( n29210 , n29209 , n22104 );
nand ( n29211 , n29210 , n22126 );
not ( n29212 , n29211 );
or ( n29213 , n29208 , n29212 );
or ( n29214 , n29207 , n29211 );
nand ( n29215 , n29213 , n29214 );
buf ( n29216 , n29215 );
nand ( n29217 , n29216 , n28427 );
nand ( n29218 , n28458 , n12280 );
and ( n29219 , n29206 , n29217 , n29218 );
not ( n29220 , n28454 );
not ( n29221 , n12143 );
and ( n29222 , n29220 , n29221 );
buf ( n29223 , n22022 );
not ( n29224 , n29223 );
not ( n29225 , n29224 );
nor ( n29226 , n28221 , n28223 );
not ( n29227 , n29226 );
or ( n29228 , n29225 , n29227 );
or ( n29229 , n29226 , n29224 );
nand ( n29230 , n29228 , n29229 );
buf ( n29231 , n29230 );
and ( n29232 , n29231 , n28438 );
nor ( n29233 , n29222 , n29232 );
nand ( n29234 , n28450 , n9159 );
nand ( n29235 , n29234 , n11137 );
nand ( n29236 , n29219 , n29233 , n29235 );
buf ( n29237 , n29236 );
buf ( n29238 , n29237 );
buf ( n29239 , n275554 );
and ( n29240 , n22904 , n275702 );
not ( n29241 , n14545 );
not ( n29242 , n17542 );
or ( n29243 , n29241 , n29242 );
buf ( n29244 , n13102 );
buf ( n29245 , n29244 );
buf ( n29246 , n14773 );
xor ( n29247 , n29245 , n29246 );
buf ( n29248 , n29247 );
buf ( n29249 , n29248 );
and ( n29250 , n23151 , n29249 );
buf ( n29251 , n29244 );
buf ( n29252 , n14770 );
xor ( n29253 , n29251 , n29252 );
buf ( n29254 , n29253 );
buf ( n29255 , n29254 );
nand ( n29256 , n22912 , n29255 );
and ( n29257 , n13373 , n29256 );
buf ( n29258 , n12742 );
not ( n29259 , n29258 );
and ( n29260 , n13372 , n29259 );
nor ( n29261 , n29257 , n29260 );
nor ( n29262 , n29250 , n29261 );
or ( n29263 , n29044 , n29262 );
nand ( n29264 , n29243 , n29263 );
nor ( n29265 , n29240 , n29264 );
nand ( n29266 , n22914 , n13084 );
buf ( n29267 , n23017 );
not ( n29268 , n29267 );
buf ( n29269 , n23034 );
buf ( n29270 , n23024 );
nand ( n29271 , n29269 , n29270 );
buf ( n29272 , n29271 );
buf ( n29273 , n29272 );
not ( n29274 , n29273 );
or ( n29275 , n29268 , n29274 );
buf ( n29276 , n29272 );
buf ( n29277 , n23017 );
or ( n29278 , n29276 , n29277 );
nand ( n29279 , n29275 , n29278 );
buf ( n29280 , n29279 );
buf ( n29281 , n29280 );
nand ( n29282 , n22918 , n29281 );
buf ( n29283 , n23246 );
not ( n29284 , n29283 );
buf ( n29285 , n23263 );
buf ( n29286 , n23253 );
nand ( n29287 , n29285 , n29286 );
buf ( n29288 , n29287 );
buf ( n29289 , n29288 );
not ( n29290 , n29289 );
or ( n29291 , n29284 , n29290 );
buf ( n29292 , n29288 );
buf ( n29293 , n23246 );
or ( n29294 , n29292 , n29293 );
nand ( n29295 , n29291 , n29294 );
buf ( n29296 , n29295 );
buf ( n29297 , n29296 );
nand ( n29298 , n23152 , n29297 );
nand ( n29299 , n29265 , n29266 , n29282 , n29298 );
buf ( n29300 , n29299 );
buf ( n29301 , n29300 );
not ( n29302 , n275550 );
buf ( n29303 , n29302 );
buf ( n29304 , n29303 );
not ( n29305 , n275929 );
buf ( n29306 , n29305 );
buf ( n29307 , n29306 );
buf ( n29308 , n275554 );
buf ( n29309 , n275554 );
buf ( n29310 , n275554 );
not ( n29311 , n14532 );
not ( n29312 , n20950 );
or ( n29313 , n29311 , n29312 );
or ( n29314 , n21691 , n23887 );
nand ( n29315 , n29313 , n29314 );
buf ( n29316 , n29315 );
buf ( n29317 , n29316 );
not ( n29318 , n275550 );
buf ( n29319 , n29318 );
buf ( n29320 , n29319 );
buf ( n29321 , n23511 );
buf ( n29322 , n23584 );
nand ( n29323 , n29321 , n29322 );
buf ( n29324 , n29323 );
buf ( n29325 , n29324 );
not ( n29326 , n29325 );
buf ( n29327 , n23498 );
not ( n29328 , n29327 );
buf ( n29329 , n23568 );
not ( n29330 , n29329 );
or ( n29331 , n29328 , n29330 );
buf ( n29332 , n23575 );
not ( n29333 , n29332 );
buf ( n29334 , n29333 );
buf ( n29335 , n29334 );
nand ( n29336 , n29331 , n29335 );
buf ( n29337 , n29336 );
buf ( n29338 , n29337 );
not ( n29339 , n29338 );
or ( n29340 , n29326 , n29339 );
buf ( n29341 , n29337 );
buf ( n29342 , n29324 );
or ( n29343 , n29341 , n29342 );
nand ( n29344 , n29340 , n29343 );
buf ( n29345 , n29344 );
buf ( n29346 , n29345 );
nand ( n29347 , n29346 , n23603 );
nand ( n29348 , n23620 , n23646 );
not ( n29349 , n29348 );
not ( n29350 , n23616 );
not ( n29351 , n28417 );
or ( n29352 , n29350 , n29351 );
not ( n29353 , n23642 );
nand ( n29354 , n29352 , n29353 );
not ( n29355 , n29354 );
or ( n29356 , n29349 , n29355 );
or ( n29357 , n29354 , n29348 );
nand ( n29358 , n29356 , n29357 );
buf ( n29359 , n29358 );
nand ( n29360 , n29359 , n23655 );
not ( n29361 , n23663 );
not ( n29362 , n29361 );
not ( n29363 , n23662 );
nor ( n29364 , n29363 , n27569 );
not ( n29365 , n29364 );
or ( n29366 , n29362 , n29365 );
or ( n29367 , n29364 , n29361 );
nand ( n29368 , n29366 , n29367 );
buf ( n29369 , n29368 );
not ( n29370 , n23672 );
not ( n29371 , n29370 );
and ( n29372 , n29369 , n29371 );
or ( n29373 , n22008 , n12270 );
or ( n29374 , n23680 , n12131 );
nand ( n29375 , n29373 , n29374 );
nor ( n29376 , n29372 , n29375 );
and ( n29377 , n29347 , n29360 , n29376 );
or ( n29378 , n29377 , n22193 );
buf ( n29379 , n27590 );
not ( n29380 , n29379 );
or ( n29381 , n29380 , n11631 );
nand ( n29382 , n29378 , n29381 );
buf ( n29383 , n29382 );
buf ( n29384 , n29383 );
buf ( n29385 , n275554 );
buf ( n29386 , n275554 );
buf ( n29387 , n275554 );
not ( n29388 , n275550 );
buf ( n29389 , n29388 );
buf ( n29390 , n29389 );
not ( n29391 , n275925 );
buf ( n29392 , n29391 );
buf ( n29393 , n29392 );
not ( n29394 , n19473 );
not ( n29395 , n29394 );
and ( n29396 , n22799 , n29395 );
not ( n29397 , n22799 );
buf ( n29398 , n21115 );
not ( n29399 , n29398 );
not ( n29400 , n24632 );
nand ( n29401 , n19604 , n26555 , n26556 );
not ( n29402 , n29401 );
nand ( n29403 , n29400 , n29402 );
not ( n29404 , n29403 );
or ( n29405 , n29399 , n29404 );
or ( n29406 , n29398 , n29403 );
nand ( n29407 , n29405 , n29406 );
buf ( n29408 , n29407 );
and ( n29409 , n29397 , n29408 );
nor ( n29410 , n29396 , n29409 );
not ( n29411 , n29410 );
and ( n29412 , n29411 , n21174 );
not ( n29413 , n21001 );
or ( n29414 , n21454 , n21456 );
nand ( n29415 , n29414 , n21488 );
not ( n29416 , n29415 );
not ( n29417 , n21417 );
not ( n29418 , n29417 );
not ( n29419 , n20337 );
or ( n29420 , n29418 , n29419 );
not ( n29421 , n21485 );
nand ( n29422 , n29420 , n29421 );
not ( n29423 , n29422 );
or ( n29424 , n29416 , n29423 );
or ( n29425 , n29422 , n29415 );
nand ( n29426 , n29424 , n29425 );
buf ( n29427 , n29426 );
not ( n29428 , n29427 );
or ( n29429 , n29413 , n29428 );
not ( n29430 , n21546 );
not ( n29431 , n21578 );
nand ( n29432 , n29430 , n29431 );
not ( n29433 , n29432 );
nor ( n29434 , n21561 , n20401 );
not ( n29435 , n29434 );
not ( n29436 , n20500 );
or ( n29437 , n29435 , n29436 );
not ( n29438 , n21576 );
nand ( n29439 , n29437 , n29438 );
not ( n29440 , n29439 );
or ( n29441 , n29433 , n29440 );
or ( n29442 , n29439 , n29432 );
nand ( n29443 , n29441 , n29442 );
buf ( n29444 , n29443 );
and ( n29445 , n29444 , n19358 );
not ( n29446 , n19290 );
not ( n29447 , n21610 );
not ( n29448 , n29447 );
nand ( n29449 , n20547 , n21606 );
not ( n29450 , n29449 );
or ( n29451 , n29448 , n29450 );
or ( n29452 , n29449 , n29447 );
nand ( n29453 , n29451 , n29452 );
buf ( n29454 , n29453 );
not ( n29455 , n29454 );
or ( n29456 , n29446 , n29455 );
buf ( n29457 , n21609 );
buf ( n29458 , n29457 );
buf ( n29459 , n29458 );
nand ( n29460 , n27619 , n29459 );
nand ( n29461 , n29456 , n29460 );
nor ( n29462 , n29445 , n29461 );
nand ( n29463 , n29429 , n29462 );
nor ( n29464 , n29412 , n29463 );
or ( n29465 , n29464 , n21030 );
nand ( n29466 , n21030 , n19005 );
nand ( n29467 , n29465 , n29466 );
buf ( n29468 , n29467 );
buf ( n29469 , n29468 );
or ( n29470 , n23989 , n19634 );
not ( n29471 , n19647 );
and ( n29472 , n24296 , n29471 );
and ( n29473 , n19660 , n18766 );
nand ( n29474 , n29473 , n18750 );
not ( n29475 , n19019 );
nor ( n29476 , n29474 , n29475 );
nand ( n29477 , n29476 , n18991 );
not ( n29478 , n18719 );
nor ( n29479 , n29477 , n29478 );
nand ( n29480 , n29479 , n18697 );
not ( n29481 , n18957 );
nor ( n29482 , n29480 , n29481 );
not ( n29483 , n18934 );
and ( n29484 , n29482 , n29483 );
not ( n29485 , n29482 );
and ( n29486 , n29485 , n18935 );
nor ( n29487 , n29484 , n29486 );
not ( n29488 , n29487 );
not ( n29489 , n29488 );
not ( n29490 , n19648 );
or ( n29491 , n29489 , n29490 );
not ( n29492 , n20559 );
nand ( n29493 , n24320 , n29492 );
not ( n29494 , n20562 );
nand ( n29495 , n29494 , n24325 );
nor ( n29496 , n19639 , n29483 );
not ( n29497 , n29496 );
and ( n29498 , n29493 , n29495 , n29497 );
nand ( n29499 , n29491 , n29498 );
nor ( n29500 , n29472 , n29499 );
nand ( n29501 , n24213 , n20353 );
and ( n29502 , n29500 , n29501 );
nand ( n29503 , n29470 , n29502 );
buf ( n29504 , n29503 );
buf ( n29505 , n29504 );
buf ( n29506 , n21136 );
and ( n29507 , n18208 , n29506 );
not ( n29508 , n18208 );
not ( n29509 , n21163 );
nand ( n29510 , n19069 , n21141 );
not ( n29511 , n29510 );
or ( n29512 , n29509 , n29511 );
or ( n29513 , n29510 , n21163 );
nand ( n29514 , n29512 , n29513 );
buf ( n29515 , n29514 );
and ( n29516 , n29508 , n29515 );
nor ( n29517 , n29507 , n29516 );
or ( n29518 , n29517 , n19216 );
nand ( n29519 , n21533 , n21584 );
not ( n29520 , n29519 );
nor ( n29521 , n21563 , n21546 );
not ( n29522 , n29521 );
not ( n29523 , n20500 );
or ( n29524 , n29522 , n29523 );
not ( n29525 , n29430 );
not ( n29526 , n21576 );
or ( n29527 , n29525 , n29526 );
nand ( n29528 , n29527 , n29431 );
not ( n29529 , n29528 );
nand ( n29530 , n29524 , n29529 );
not ( n29531 , n29530 );
or ( n29532 , n29520 , n29531 );
or ( n29533 , n29530 , n29519 );
nand ( n29534 , n29532 , n29533 );
buf ( n29535 , n29534 );
and ( n29536 , n29535 , n19360 );
not ( n29537 , n19318 );
not ( n29538 , n29537 );
not ( n29539 , n18990 );
and ( n29540 , n29476 , n29539 );
not ( n29541 , n29476 );
and ( n29542 , n29541 , n18991 );
nor ( n29543 , n29540 , n29542 );
not ( n29544 , n29543 );
and ( n29545 , n29538 , n29544 );
buf ( n29546 , n21607 );
buf ( n29547 , n29546 );
buf ( n29548 , n29547 );
and ( n29549 , n19221 , n29548 );
nor ( n29550 , n29545 , n29549 );
not ( n29551 , n21608 );
and ( n29552 , n20547 , n21606 , n29447 );
not ( n29553 , n29552 );
or ( n29554 , n29551 , n29553 );
or ( n29555 , n29552 , n21608 );
nand ( n29556 , n29554 , n29555 );
buf ( n29557 , n29556 );
nand ( n29558 , n29557 , n29075 );
nand ( n29559 , n19387 , n18987 );
nand ( n29560 , n29550 , n29558 , n29559 );
nor ( n29561 , n29536 , n29560 );
nand ( n29562 , n21468 , n21489 );
not ( n29563 , n29562 );
not ( n29564 , n29414 );
nor ( n29565 , n29564 , n21417 );
not ( n29566 , n29565 );
not ( n29567 , n20337 );
or ( n29568 , n29566 , n29567 );
not ( n29569 , n29414 );
not ( n29570 , n21485 );
or ( n29571 , n29569 , n29570 );
nand ( n29572 , n29571 , n21488 );
not ( n29573 , n29572 );
nand ( n29574 , n29568 , n29573 );
not ( n29575 , n29574 );
or ( n29576 , n29563 , n29575 );
or ( n29577 , n29574 , n29562 );
nand ( n29578 , n29576 , n29577 );
buf ( n29579 , n29578 );
nand ( n29580 , n29579 , n19354 );
and ( n29581 , n29561 , n29580 );
nand ( n29582 , n29518 , n29581 );
buf ( n29583 , n29582 );
buf ( n29584 , n29583 );
buf ( n29585 , n275554 );
not ( n29586 , n275550 );
buf ( n29587 , n29586 );
buf ( n29588 , n29587 );
buf ( n29589 , n275554 );
not ( n29590 , n275925 );
buf ( n29591 , n29590 );
buf ( n29592 , n29591 );
not ( n29593 , n275925 );
buf ( n29594 , n29593 );
buf ( n29595 , n29594 );
and ( n29596 , n27179 , n277957 );
not ( n29597 , n27179 );
not ( n29598 , n27489 );
not ( n29599 , n29598 );
not ( n29600 , n29599 );
buf ( n29601 , n277977 );
buf ( n29602 , n29601 );
not ( n29603 , n29602 );
buf ( n29604 , n278005 );
buf ( n29605 , n29604 );
not ( n29606 , n29605 );
buf ( n29607 , n29606 );
buf ( n29608 , n29607 );
nand ( n29609 , n29603 , n29608 );
buf ( n29610 , n29609 );
buf ( n29611 , n29610 );
buf ( n29612 , n29607 );
not ( n29613 , n29612 );
buf ( n29614 , n29601 );
nand ( n29615 , n29613 , n29614 );
buf ( n29616 , n29615 );
buf ( n29617 , n29616 );
nand ( n29618 , n29611 , n29617 );
buf ( n29619 , n29618 );
buf ( n29620 , n29619 );
not ( n29621 , n29620 );
buf ( n29622 , n277951 );
buf ( n29623 , n29622 );
not ( n29624 , n29623 );
buf ( n29625 , n29624 );
buf ( n29626 , n29625 );
buf ( n29627 , n277930 );
buf ( n29628 , n29627 );
not ( n29629 , n29628 );
buf ( n29630 , n29629 );
buf ( n29631 , n29630 );
nand ( n29632 , n29626 , n29631 );
buf ( n29633 , n29632 );
buf ( n29634 , n29633 );
buf ( n29635 , n29634 );
not ( n29636 , n29635 );
buf ( n29637 , n27281 );
buf ( n29638 , n278025 );
buf ( n29639 , n29638 );
not ( n29640 , n29639 );
buf ( n29641 , n29640 );
buf ( n29642 , n29641 );
buf ( n29643 , n278054 );
buf ( n29644 , n29643 );
not ( n29645 , n29644 );
buf ( n29646 , n29645 );
buf ( n29647 , n29646 );
nand ( n29648 , n29642 , n29647 );
buf ( n29649 , n29648 );
buf ( n29650 , n29649 );
nand ( n29651 , n29637 , n29650 );
buf ( n29652 , n29651 );
buf ( n29653 , n29652 );
nor ( n29654 , n29636 , n29653 );
buf ( n29655 , n29654 );
buf ( n29656 , n29655 );
not ( n29657 , n29656 );
buf ( n29658 , n27479 );
not ( n29659 , n29658 );
or ( n29660 , n29657 , n29659 );
buf ( n29661 , n29634 );
not ( n29662 , n29661 );
buf ( n29663 , n29649 );
not ( n29664 , n29663 );
buf ( n29665 , n27273 );
not ( n29666 , n29665 );
or ( n29667 , n29664 , n29666 );
buf ( n29668 , n29638 );
buf ( n29669 , n29643 );
nand ( n29670 , n29668 , n29669 );
buf ( n29671 , n29670 );
buf ( n29672 , n29671 );
nand ( n29673 , n29667 , n29672 );
buf ( n29674 , n29673 );
buf ( n29675 , n29674 );
not ( n29676 , n29675 );
or ( n29677 , n29662 , n29676 );
buf ( n29678 , n29622 );
buf ( n29679 , n29627 );
and ( n29680 , n29678 , n29679 );
buf ( n29681 , n29680 );
buf ( n29682 , n29681 );
not ( n29683 , n29682 );
buf ( n29684 , n29683 );
buf ( n29685 , n29684 );
nand ( n29686 , n29677 , n29685 );
buf ( n29687 , n29686 );
buf ( n29688 , n29687 );
not ( n29689 , n29688 );
buf ( n29690 , n29689 );
buf ( n29691 , n29690 );
nand ( n29692 , n29660 , n29691 );
buf ( n29693 , n29692 );
buf ( n29694 , n29693 );
not ( n29695 , n29694 );
or ( n29696 , n29621 , n29695 );
buf ( n29697 , n29693 );
buf ( n29698 , n29619 );
or ( n29699 , n29697 , n29698 );
nand ( n29700 , n29696 , n29699 );
buf ( n29701 , n29700 );
buf ( n29702 , n29701 );
not ( n29703 , n29702 );
or ( n29704 , n29600 , n29703 );
buf ( n29705 , n277977 );
not ( n29706 , n29705 );
buf ( n29707 , n278005 );
nand ( n29708 , n29706 , n29707 );
not ( n29709 , n29707 );
nand ( n29710 , n29709 , n29705 );
nand ( n29711 , n29708 , n29710 );
not ( n29712 , n29711 );
buf ( n29713 , n277951 );
not ( n29714 , n29713 );
buf ( n29715 , n277930 );
nand ( n29716 , n29714 , n29715 );
buf ( n29717 , n29716 );
not ( n29718 , n29717 );
buf ( n29719 , n278025 );
not ( n29720 , n29719 );
buf ( n29721 , n278054 );
nand ( n29722 , n29720 , n29721 );
buf ( n29723 , n29722 );
nand ( n29724 , n27185 , n29723 );
buf ( n29725 , n29724 );
nor ( n29726 , n29718 , n29725 );
not ( n29727 , n29726 );
nand ( n29728 , n27233 , n27259 );
not ( n29729 , n29728 );
or ( n29730 , n29727 , n29729 );
not ( n29731 , n29722 );
not ( n29732 , n27186 );
or ( n29733 , n29731 , n29732 );
not ( n29734 , n29721 );
nand ( n29735 , n29734 , n29719 );
nand ( n29736 , n29733 , n29735 );
nand ( n29737 , n29736 , n29717 );
not ( n29738 , n29715 );
and ( n29739 , n29713 , n29738 );
not ( n29740 , n29739 );
and ( n29741 , n29737 , n29740 );
nand ( n29742 , n29730 , n29741 );
not ( n29743 , n29742 );
or ( n29744 , n29712 , n29743 );
or ( n29745 , n29742 , n29711 );
nand ( n29746 , n29744 , n29745 );
buf ( n29747 , n29746 );
and ( n29748 , n29747 , n23655 );
not ( n29749 , n22052 );
buf ( n29750 , n277842 );
not ( n29751 , n29750 );
not ( n29752 , n29751 );
nand ( n29753 , n27512 , n27492 );
buf ( n29754 , n277951 );
buf ( n29755 , n29754 );
buf ( n29756 , n277977 );
nand ( n29757 , n29755 , n29756 );
nor ( n29758 , n29753 , n29757 );
buf ( n29759 , n29758 );
not ( n29760 , n29759 );
or ( n29761 , n29752 , n29760 );
or ( n29762 , n29759 , n29751 );
nand ( n29763 , n29761 , n29762 );
buf ( n29764 , n29763 );
not ( n29765 , n29764 );
or ( n29766 , n29749 , n29765 );
and ( n29767 , n27520 , n12355 );
not ( n29768 , n22014 );
and ( n29769 , n29768 , n12156 );
nor ( n29770 , n29767 , n29769 );
nand ( n29771 , n29766 , n29770 );
nor ( n29772 , n29748 , n29771 );
nand ( n29773 , n29704 , n29772 );
and ( n29774 , n29597 , n29773 );
or ( n29775 , n29596 , n29774 );
buf ( n29776 , n29775 );
buf ( n29777 , n29776 );
buf ( n29778 , n23914 );
not ( n29779 , n29778 );
buf ( n29780 , n27764 );
buf ( n29781 , n27795 );
buf ( n29782 , n27806 );
nand ( n29783 , n29781 , n29782 );
buf ( n29784 , n29783 );
buf ( n29785 , n29784 );
nor ( n29786 , n29780 , n29785 );
buf ( n29787 , n29786 );
buf ( n29788 , n29787 );
nand ( n29789 , n29779 , n29788 );
buf ( n29790 , n29789 );
buf ( n29791 , n29790 );
buf ( n29792 , n18518 );
xnor ( n29793 , n29791 , n29792 );
buf ( n29794 , n29793 );
buf ( n29795 , n29794 );
and ( n29796 , n26516 , n29795 );
not ( n29797 , n26516 );
buf ( n29798 , n23914 );
not ( n29799 , n29798 );
buf ( n29800 , n27764 );
buf ( n29801 , n18521 );
buf ( n29802 , n27792 );
nor ( n29803 , n29801 , n29802 );
buf ( n29804 , n29803 );
buf ( n29805 , n29804 );
buf ( n29806 , n18445 );
buf ( n29807 , n29806 );
nand ( n29808 , n29805 , n29807 );
buf ( n29809 , n29808 );
buf ( n29810 , n29809 );
nor ( n29811 , n29800 , n29810 );
buf ( n29812 , n29811 );
buf ( n29813 , n29812 );
nand ( n29814 , n29799 , n29813 );
buf ( n29815 , n29814 );
buf ( n29816 , n29815 );
buf ( n29817 , n18464 );
xnor ( n29818 , n29816 , n29817 );
buf ( n29819 , n29818 );
buf ( n29820 , n29819 );
buf ( n29821 , n29820 );
buf ( n29822 , n29821 );
not ( n29823 , n29822 );
buf ( n29824 , n29795 );
nand ( n29825 , n27833 , n27811 , n29824 );
not ( n29826 , n26600 );
nor ( n29827 , n29825 , n29826 );
not ( n29828 , n26583 );
buf ( n29829 , n27815 );
nor ( n29830 , n29828 , n29829 , n26630 );
and ( n29831 , n29827 , n29830 , n26554 );
buf ( n29832 , n23914 );
buf ( n29833 , n27767 );
buf ( n29834 , n29804 );
nand ( n29835 , n29833 , n29834 );
buf ( n29836 , n29835 );
buf ( n29837 , n29836 );
nor ( n29838 , n29832 , n29837 );
buf ( n29839 , n29838 );
buf ( n29840 , n29839 );
buf ( n29841 , n29806 );
not ( n29842 , n29841 );
buf ( n29843 , n29842 );
buf ( n29844 , n29843 );
nor ( n29845 , n29840 , n29844 );
buf ( n29846 , n29845 );
buf ( n29847 , n29846 );
not ( n29848 , n29847 );
buf ( n29849 , n29839 );
buf ( n29850 , n29843 );
nand ( n29851 , n29849 , n29850 );
buf ( n29852 , n29851 );
buf ( n29853 , n29852 );
nand ( n29854 , n29848 , n29853 );
buf ( n29855 , n29854 );
buf ( n29856 , n29855 );
buf ( n29857 , n29856 );
nand ( n29858 , n29831 , n29857 );
not ( n29859 , n29858 );
or ( n29860 , n29823 , n29859 );
or ( n29861 , n29858 , n29822 );
nand ( n29862 , n29860 , n29861 );
buf ( n29863 , n29862 );
and ( n29864 , n29797 , n29863 );
nor ( n29865 , n29796 , n29864 );
not ( n29866 , n19635 );
or ( n29867 , n29865 , n29866 );
not ( n29868 , n277527 );
buf ( n29869 , n22422 );
buf ( n29870 , n22726 );
or ( n29871 , n29869 , n29870 );
buf ( n29872 , n29871 );
buf ( n29873 , n29872 );
not ( n29874 , n29873 );
buf ( n29875 , n22415 );
buf ( n29876 , n22449 );
not ( n29877 , n29876 );
buf ( n29878 , n22429 );
nor ( n29879 , n29877 , n29878 );
buf ( n29880 , n29879 );
buf ( n29881 , n29880 );
and ( n29882 , n29875 , n29881 );
buf ( n29883 , n29882 );
buf ( n29884 , n29883 );
not ( n29885 , n29884 );
buf ( n29886 , n22593 );
not ( n29887 , n29886 );
or ( n29888 , n29885 , n29887 );
buf ( n29889 , n22687 );
buf ( n29890 , n29880 );
and ( n29891 , n29889 , n29890 );
buf ( n29892 , n22708 );
not ( n29893 , n29892 );
buf ( n29894 , n29893 );
buf ( n29895 , n29894 );
buf ( n29896 , n22429 );
or ( n29897 , n29895 , n29896 );
buf ( n29898 , n22719 );
nand ( n29899 , n29897 , n29898 );
buf ( n29900 , n29899 );
buf ( n29901 , n29900 );
nor ( n29902 , n29891 , n29901 );
buf ( n29903 , n29902 );
buf ( n29904 , n29903 );
nand ( n29905 , n29888 , n29904 );
buf ( n29906 , n29905 );
buf ( n29907 , n29906 );
not ( n29908 , n29907 );
or ( n29909 , n29874 , n29908 );
buf ( n29910 , n29906 );
buf ( n29911 , n29872 );
or ( n29912 , n29910 , n29911 );
nand ( n29913 , n29909 , n29912 );
buf ( n29914 , n29913 );
buf ( n29915 , n29914 );
not ( n29916 , n29915 );
or ( n29917 , n29868 , n29916 );
nand ( n29918 , n277390 , n9740 );
nand ( n29919 , n29917 , n29918 );
and ( n29920 , n25049 , n29919 );
buf ( n29921 , n29920 );
not ( n29922 , n29921 );
buf ( n29923 , n18517 );
buf ( n29924 , n29923 );
and ( n29925 , n29922 , n29924 );
not ( n29926 , n277527 );
buf ( n29927 , n22459 );
buf ( n29928 , n22741 );
nand ( n29929 , n29927 , n29928 );
buf ( n29930 , n29929 );
buf ( n29931 , n29930 );
not ( n29932 , n29931 );
buf ( n29933 , n22415 );
buf ( n29934 , n22452 );
and ( n29935 , n29933 , n29934 );
buf ( n29936 , n29935 );
buf ( n29937 , n29936 );
not ( n29938 , n29937 );
buf ( n29939 , n22593 );
not ( n29940 , n29939 );
or ( n29941 , n29938 , n29940 );
buf ( n29942 , n22687 );
buf ( n29943 , n22452 );
and ( n29944 , n29942 , n29943 );
buf ( n29945 , n22732 );
nor ( n29946 , n29944 , n29945 );
buf ( n29947 , n29946 );
buf ( n29948 , n29947 );
nand ( n29949 , n29941 , n29948 );
buf ( n29950 , n29949 );
buf ( n29951 , n29950 );
not ( n29952 , n29951 );
or ( n29953 , n29932 , n29952 );
buf ( n29954 , n29950 );
buf ( n29955 , n29930 );
or ( n29956 , n29954 , n29955 );
nand ( n29957 , n29953 , n29956 );
buf ( n29958 , n29957 );
buf ( n29959 , n29958 );
not ( n29960 , n29959 );
or ( n29961 , n29926 , n29960 );
nand ( n29962 , n277390 , n9783 );
nand ( n29963 , n29961 , n29962 );
and ( n29964 , n25049 , n29963 );
buf ( n29965 , n29964 );
not ( n29966 , n29965 );
buf ( n29967 , n18444 );
buf ( n29968 , n29967 );
buf ( n29969 , n29968 );
xor ( n29970 , n29966 , n29969 );
or ( n29971 , n29925 , n29970 );
nand ( n29972 , n29970 , n29925 );
nand ( n29973 , n29971 , n29972 );
not ( n29974 , n29973 );
xor ( n29975 , n29922 , n29924 );
not ( n29976 , n29975 );
buf ( n29977 , n18491 );
buf ( n29978 , n29977 );
not ( n29979 , n277603 );
buf ( n29980 , n22429 );
not ( n29981 , n29980 );
buf ( n29982 , n22719 );
nand ( n29983 , n29981 , n29982 );
buf ( n29984 , n29983 );
buf ( n29985 , n29984 );
not ( n29986 , n29985 );
buf ( n29987 , n22593 );
buf ( n29988 , n22415 );
buf ( n29989 , n22449 );
and ( n29990 , n29988 , n29989 );
buf ( n29991 , n29990 );
buf ( n29992 , n29991 );
nand ( n29993 , n29987 , n29992 );
buf ( n29994 , n29993 );
buf ( n29995 , n29994 );
buf ( n29996 , n22687 );
buf ( n29997 , n22449 );
and ( n29998 , n29996 , n29997 );
buf ( n29999 , n22708 );
nor ( n30000 , n29998 , n29999 );
buf ( n30001 , n30000 );
buf ( n30002 , n30001 );
nand ( n30003 , n29995 , n30002 );
buf ( n30004 , n30003 );
buf ( n30005 , n30004 );
not ( n30006 , n30005 );
or ( n30007 , n29986 , n30006 );
buf ( n30008 , n30004 );
buf ( n30009 , n29984 );
or ( n30010 , n30008 , n30009 );
nand ( n30011 , n30007 , n30010 );
buf ( n30012 , n30011 );
buf ( n30013 , n30012 );
not ( n30014 , n30013 );
or ( n30015 , n29979 , n30014 );
nand ( n30016 , n9433 , n9748 );
nand ( n30017 , n30015 , n30016 );
nand ( n30018 , n25049 , n30017 );
not ( n30019 , n30018 );
buf ( n30020 , n30019 );
not ( n30021 , n30020 );
and ( n30022 , n29978 , n30021 );
not ( n30023 , n30022 );
nand ( n30024 , n29976 , n30023 );
not ( n30025 , n30020 );
not ( n30026 , n29978 );
or ( n30027 , n30025 , n30026 );
not ( n30028 , n29978 );
nand ( n30029 , n30028 , n30021 );
nand ( n30030 , n30027 , n30029 );
not ( n30031 , n30030 );
not ( n30032 , n27889 );
nor ( n30033 , n30032 , n27886 );
not ( n30034 , n30033 );
nand ( n30035 , n30031 , n30034 );
nand ( n30036 , n30024 , n30035 );
not ( n30037 , n28022 );
nand ( n30038 , n30037 , n27937 );
nor ( n30039 , n30036 , n30038 );
not ( n30040 , n30039 );
nor ( n30041 , n28014 , n30040 );
not ( n30042 , n30041 );
not ( n30043 , n24203 );
not ( n30044 , n30043 );
or ( n30045 , n30042 , n30044 );
not ( n30046 , n28037 );
not ( n30047 , n30040 );
and ( n30048 , n30046 , n30047 );
not ( n30049 , n30036 );
not ( n30050 , n30049 );
or ( n30051 , n27938 , n28041 );
nand ( n30052 , n30051 , n27940 );
not ( n30053 , n30052 );
or ( n30054 , n30050 , n30053 );
not ( n30055 , n30024 );
not ( n30056 , n30055 );
nand ( n30057 , n30030 , n30033 );
not ( n30058 , n30057 );
and ( n30059 , n30056 , n30058 );
or ( n30060 , n29976 , n30023 );
not ( n30061 , n30060 );
nor ( n30062 , n30059 , n30061 );
nand ( n30063 , n30054 , n30062 );
nor ( n30064 , n30048 , n30063 );
nand ( n30065 , n30045 , n30064 );
not ( n30066 , n30065 );
or ( n30067 , n29974 , n30066 );
or ( n30068 , n30065 , n29973 );
nand ( n30069 , n30067 , n30068 );
buf ( n30070 , n30069 );
nand ( n30071 , n30070 , n20353 );
buf ( n30072 , n29964 );
buf ( n30073 , n30072 );
buf ( n30074 , n29968 );
xor ( n30075 , n30073 , n30074 );
buf ( n30076 , n29920 );
buf ( n30077 , n30076 );
buf ( n30078 , n29923 );
buf ( n30079 , n30078 );
and ( n30080 , n30077 , n30079 );
or ( n30081 , n30075 , n30080 );
nand ( n30082 , n30075 , n30080 );
nand ( n30083 , n30081 , n30082 );
not ( n30084 , n30083 );
xor ( n30085 , n30077 , n30079 );
buf ( n30086 , n29977 );
buf ( n30087 , n30086 );
buf ( n30088 , n30019 );
and ( n30089 , n30087 , n30088 );
nor ( n30090 , n30085 , n30089 );
not ( n30091 , n30088 );
not ( n30092 , n30091 );
not ( n30093 , n30087 );
or ( n30094 , n30092 , n30093 );
not ( n30095 , n30087 );
nand ( n30096 , n30095 , n30088 );
nand ( n30097 , n30094 , n30096 );
and ( n30098 , n28051 , n28053 );
nor ( n30099 , n30097 , n30098 );
nor ( n30100 , n30090 , n30099 );
nor ( n30101 , n28060 , n28089 );
and ( n30102 , n30100 , n30101 );
not ( n30103 , n30102 );
nor ( n30104 , n30103 , n28079 );
not ( n30105 , n30104 );
not ( n30106 , n28092 );
or ( n30107 , n30105 , n30106 );
not ( n30108 , n30102 );
not ( n30109 , n28109 );
or ( n30110 , n30108 , n30109 );
not ( n30111 , n30100 );
or ( n30112 , n28060 , n28112 );
nand ( n30113 , n30112 , n28062 );
not ( n30114 , n30113 );
or ( n30115 , n30111 , n30114 );
not ( n30116 , n30090 );
nand ( n30117 , n30097 , n30098 );
not ( n30118 , n30117 );
and ( n30119 , n30116 , n30118 );
and ( n30120 , n30085 , n30089 );
nor ( n30121 , n30119 , n30120 );
nand ( n30122 , n30115 , n30121 );
not ( n30123 , n30122 );
nand ( n30124 , n30110 , n30123 );
not ( n30125 , n30124 );
nand ( n30126 , n30107 , n30125 );
not ( n30127 , n30126 );
or ( n30128 , n30084 , n30127 );
or ( n30129 , n30126 , n30083 );
nand ( n30130 , n30128 , n30129 );
buf ( n30131 , n30130 );
not ( n30132 , n19647 );
nand ( n30133 , n30131 , n30132 );
not ( n30134 , n18439 );
nand ( n30135 , n29482 , n18935 );
not ( n30136 , n18613 );
nor ( n30137 , n30135 , n30136 );
nand ( n30138 , n30137 , n18592 );
not ( n30139 , n18667 );
nor ( n30140 , n30138 , n30139 );
and ( n30141 , n30140 , n18819 );
nand ( n30142 , n30141 , n18552 );
not ( n30143 , n18524 );
nor ( n30144 , n30142 , n30143 );
and ( n30145 , n30144 , n18789 );
nand ( n30146 , n30145 , n18653 );
not ( n30147 , n18486 );
nor ( n30148 , n30146 , n30147 );
and ( n30149 , n30148 , n18508 );
not ( n30150 , n30149 );
or ( n30151 , n30134 , n30150 );
or ( n30152 , n30149 , n18439 );
nand ( n30153 , n30151 , n30152 );
and ( n30154 , n30153 , n19650 );
buf ( n30155 , n30072 );
buf ( n30156 , n30155 );
not ( n30157 , n30156 );
nand ( n30158 , n28131 , n27055 );
nor ( n30159 , n30158 , n27072 );
and ( n30160 , n27064 , n30159 );
not ( n30161 , n28122 );
buf ( n30162 , n30019 );
buf ( n30163 , n30076 );
nor ( n30164 , n30162 , n30163 );
not ( n30165 , n28126 );
nand ( n30166 , n30161 , n30164 , n30165 );
not ( n30167 , n30166 );
nand ( n30168 , n30160 , n30167 );
nor ( n30169 , n28124 , n30168 );
not ( n30170 , n30169 );
or ( n30171 , n30157 , n30170 );
or ( n30172 , n30169 , n30156 );
nand ( n30173 , n30171 , n30172 );
buf ( n30174 , n30173 );
nand ( n30175 , n30174 , n20560 );
buf ( n30176 , n30155 );
buf ( n30177 , n30176 );
nand ( n30178 , n29494 , n30177 );
not ( n30179 , n19639 );
nand ( n30180 , n30179 , n18440 );
nand ( n30181 , n30175 , n30178 , n30180 );
nor ( n30182 , n30154 , n30181 );
and ( n30183 , n30071 , n30133 , n30182 );
nand ( n30184 , n29867 , n30183 );
buf ( n30185 , n30184 );
buf ( n30186 , n30185 );
not ( n30187 , n277603 );
buf ( n30188 , n22415 );
buf ( n30189 , n22452 );
buf ( n30190 , n22459 );
and ( n30191 , n30189 , n30190 );
buf ( n30192 , n30191 );
buf ( n30193 , n30192 );
and ( n30194 , n30188 , n30193 );
buf ( n30195 , n30194 );
buf ( n30196 , n30195 );
not ( n30197 , n30196 );
buf ( n30198 , n22592 );
not ( n30199 , n30198 );
or ( n30200 , n30197 , n30199 );
buf ( n30201 , n22687 );
buf ( n30202 , n30192 );
and ( n30203 , n30201 , n30202 );
buf ( n30204 , n22459 );
not ( n30205 , n30204 );
buf ( n30206 , n22732 );
not ( n30207 , n30206 );
or ( n30208 , n30205 , n30207 );
buf ( n30209 , n22741 );
nand ( n30210 , n30208 , n30209 );
buf ( n30211 , n30210 );
buf ( n30212 , n30211 );
nor ( n30213 , n30203 , n30212 );
buf ( n30214 , n30213 );
buf ( n30215 , n30214 );
nand ( n30216 , n30200 , n30215 );
buf ( n30217 , n30216 );
buf ( n30218 , n30217 );
buf ( n30219 , n22467 );
buf ( n30220 , n22748 );
nor ( n30221 , n30219 , n30220 );
buf ( n30222 , n30221 );
buf ( n30223 , n30222 );
and ( n30224 , n30218 , n30223 );
not ( n30225 , n30218 );
buf ( n30226 , n30222 );
not ( n30227 , n30226 );
buf ( n30228 , n30227 );
buf ( n30229 , n30228 );
and ( n30230 , n30225 , n30229 );
nor ( n30231 , n30224 , n30230 );
buf ( n30232 , n30231 );
buf ( n30233 , n30232 );
not ( n30234 , n30233 );
or ( n30235 , n30187 , n30234 );
nand ( n30236 , n277983 , n9775 );
nand ( n30237 , n30235 , n30236 );
not ( n30238 , n30237 );
or ( n30239 , n30238 , n22335 );
nand ( n30240 , n18223 , n22335 );
nand ( n30241 , n30239 , n30240 );
buf ( n30242 , n30241 );
buf ( n30243 , n30242 );
and ( n30244 , n13374 , n24485 );
not ( n30245 , n13374 );
not ( n30246 , n14798 );
and ( n30247 , n14058 , n24486 , n24768 );
nand ( n30248 , n30246 , n30247 );
not ( n30249 , n24791 );
and ( n30250 , n30248 , n30249 );
not ( n30251 , n30248 );
and ( n30252 , n30251 , n24791 );
nor ( n30253 , n30250 , n30252 );
buf ( n30254 , n30253 );
and ( n30255 , n30245 , n30254 );
nor ( n30256 , n30244 , n30255 );
not ( n30257 , n30256 );
and ( n30258 , n30257 , n23788 );
not ( n30259 , n20889 );
buf ( n30260 , n24937 );
not ( n30261 , n30260 );
buf ( n30262 , n14649 );
buf ( n30263 , n30262 );
not ( n30264 , n30263 );
or ( n30265 , n30261 , n30264 );
not ( n30266 , n30260 );
not ( n30267 , n30263 );
nand ( n30268 , n30266 , n30267 );
nand ( n30269 , n30265 , n30268 );
buf ( n30270 , n14718 );
buf ( n30271 , n30270 );
buf ( n30272 , n30271 );
buf ( n30273 , n24891 );
not ( n30274 , n30273 );
and ( n30275 , n30272 , n30274 );
nor ( n30276 , n30269 , n30275 );
not ( n30277 , n30276 );
nand ( n30278 , n30269 , n30275 );
nand ( n30279 , n30277 , n30278 );
not ( n30280 , n30279 );
not ( n30281 , n24551 );
not ( n30282 , n30273 );
not ( n30283 , n30272 );
or ( n30284 , n30282 , n30283 );
not ( n30285 , n30272 );
nand ( n30286 , n30285 , n30274 );
nand ( n30287 , n30284 , n30286 );
not ( n30288 , n24543 );
nor ( n30289 , n30288 , n24539 );
nor ( n30290 , n30287 , n30289 );
nor ( n30291 , n30281 , n30290 );
nand ( n30292 , n30291 , n24555 );
nor ( n30293 , n16140 , n30292 );
not ( n30294 , n30293 );
not ( n30295 , n16913 );
or ( n30296 , n30294 , n30295 );
not ( n30297 , n30292 );
not ( n30298 , n30297 );
not ( n30299 , n16943 );
or ( n30300 , n30298 , n30299 );
not ( n30301 , n30291 );
not ( n30302 , n24565 );
or ( n30303 , n30301 , n30302 );
not ( n30304 , n30290 );
not ( n30305 , n24552 );
and ( n30306 , n30304 , n30305 );
and ( n30307 , n30287 , n30289 );
nor ( n30308 , n30306 , n30307 );
nand ( n30309 , n30303 , n30308 );
not ( n30310 , n30309 );
nand ( n30311 , n30300 , n30310 );
not ( n30312 , n30311 );
nand ( n30313 , n30296 , n30312 );
not ( n30314 , n30313 );
or ( n30315 , n30280 , n30314 );
or ( n30316 , n30313 , n30279 );
nand ( n30317 , n30315 , n30316 );
buf ( n30318 , n30317 );
not ( n30319 , n30318 );
or ( n30320 , n30259 , n30319 );
buf ( n30321 , n24937 );
buf ( n30322 , n30262 );
buf ( n30323 , n30322 );
xor ( n30324 , n30321 , n30323 );
buf ( n30325 , n24891 );
buf ( n30326 , n30270 );
buf ( n30327 , n30326 );
and ( n30328 , n30325 , n30327 );
or ( n30329 , n30324 , n30328 );
nand ( n30330 , n30324 , n30328 );
nand ( n30331 , n30329 , n30330 );
not ( n30332 , n30331 );
xor ( n30333 , n30325 , n30327 );
and ( n30334 , n24577 , n24579 );
nor ( n30335 , n30333 , n30334 );
nor ( n30336 , n30335 , n24585 );
and ( n30337 , n30336 , n24590 );
not ( n30338 , n30337 );
nor ( n30339 , n17090 , n30338 );
not ( n30340 , n30339 );
not ( n30341 , n17362 );
or ( n30342 , n30340 , n30341 );
not ( n30343 , n17389 );
not ( n30344 , n30338 );
and ( n30345 , n30343 , n30344 );
not ( n30346 , n30336 );
not ( n30347 , n24600 );
or ( n30348 , n30346 , n30347 );
not ( n30349 , n30335 );
not ( n30350 , n24587 );
and ( n30351 , n30349 , n30350 );
and ( n30352 , n30333 , n30334 );
nor ( n30353 , n30351 , n30352 );
nand ( n30354 , n30348 , n30353 );
nor ( n30355 , n30345 , n30354 );
nand ( n30356 , n30342 , n30355 );
not ( n30357 , n30356 );
or ( n30358 , n30332 , n30357 );
or ( n30359 , n30356 , n30331 );
nand ( n30360 , n30358 , n30359 );
buf ( n30361 , n30360 );
and ( n30362 , n30361 , n20926 );
not ( n30363 , n24937 );
not ( n30364 , n20940 );
or ( n30365 , n30363 , n30364 );
not ( n30366 , n24938 );
not ( n30367 , n23436 );
nand ( n30368 , n23875 , n24897 );
nor ( n30369 , n30367 , n30368 );
not ( n30370 , n30369 );
or ( n30371 , n30366 , n30370 );
or ( n30372 , n30369 , n24938 );
nand ( n30373 , n30371 , n30372 );
buf ( n30374 , n30373 );
nand ( n30375 , n30374 , n17409 );
nand ( n30376 , n30365 , n30375 );
nor ( n30377 , n30362 , n30376 );
nand ( n30378 , n30320 , n30377 );
nor ( n30379 , n30258 , n30378 );
or ( n30380 , n30379 , n21697 );
nand ( n30381 , n21696 , n14635 );
nand ( n30382 , n30380 , n30381 );
buf ( n30383 , n30382 );
buf ( n30384 , n30383 );
not ( n30385 , n275929 );
buf ( n30386 , n30385 );
buf ( n30387 , n30386 );
buf ( n30388 , n275554 );
buf ( n30389 , n275554 );
buf ( n30390 , n275554 );
buf ( n30391 , n275554 );
buf ( n30392 , n27380 );
buf ( n30393 , n27463 );
nand ( n30394 , n30392 , n30393 );
buf ( n30395 , n30394 );
buf ( n30396 , n30395 );
not ( n30397 , n30396 );
buf ( n30398 , n27342 );
buf ( n30399 , n27354 );
nand ( n30400 , n30398 , n30399 );
buf ( n30401 , n30400 );
buf ( n30402 , n30401 );
not ( n30403 , n30402 );
buf ( n30404 , n27421 );
not ( n30405 , n30404 );
buf ( n30406 , n30405 );
buf ( n30407 , n30406 );
nand ( n30408 , n30403 , n30407 );
buf ( n30409 , n30408 );
buf ( n30410 , n30409 );
buf ( n30411 , n28266 );
nor ( n30412 , n30410 , n30411 );
buf ( n30413 , n30412 );
buf ( n30414 , n30413 );
not ( n30415 , n30414 );
buf ( n30416 , n23568 );
not ( n30417 , n30416 );
or ( n30418 , n30415 , n30417 );
buf ( n30419 , n28383 );
buf ( n30420 , n30409 );
not ( n30421 , n30420 );
buf ( n30422 , n30421 );
buf ( n30423 , n30422 );
and ( n30424 , n30419 , n30423 );
buf ( n30425 , n30406 );
not ( n30426 , n30425 );
buf ( n30427 , n27446 );
not ( n30428 , n30427 );
or ( n30429 , n30426 , n30428 );
buf ( n30430 , n27457 );
buf ( n30431 , n30430 );
nand ( n30432 , n30429 , n30431 );
buf ( n30433 , n30432 );
buf ( n30434 , n30433 );
nor ( n30435 , n30424 , n30434 );
buf ( n30436 , n30435 );
buf ( n30437 , n30436 );
nand ( n30438 , n30418 , n30437 );
buf ( n30439 , n30438 );
buf ( n30440 , n30439 );
not ( n30441 , n30440 );
or ( n30442 , n30397 , n30441 );
buf ( n30443 , n30439 );
buf ( n30444 , n30395 );
or ( n30445 , n30443 , n30444 );
nand ( n30446 , n30442 , n30445 );
buf ( n30447 , n30446 );
buf ( n30448 , n30447 );
nand ( n30449 , n30448 , n23603 );
not ( n30450 , n27257 );
nand ( n30451 , n30450 , n27227 );
not ( n30452 , n30451 );
nand ( n30453 , n27215 , n27219 );
or ( n30454 , n30453 , n27251 );
nor ( n30455 , n30454 , n28312 );
not ( n30456 , n30455 );
not ( n30457 , n28417 );
or ( n30458 , n30456 , n30457 );
not ( n30459 , n30454 );
and ( n30460 , n28318 , n30459 );
not ( n30461 , n27223 );
not ( n30462 , n27249 );
or ( n30463 , n30461 , n30462 );
not ( n30464 , n27255 );
nand ( n30465 , n30463 , n30464 );
nor ( n30466 , n30460 , n30465 );
nand ( n30467 , n30458 , n30466 );
not ( n30468 , n30467 );
or ( n30469 , n30452 , n30468 );
or ( n30470 , n30467 , n30451 );
nand ( n30471 , n30469 , n30470 );
buf ( n30472 , n30471 );
nand ( n30473 , n30472 , n23655 );
not ( n30474 , n27502 );
not ( n30475 , n30474 );
nor ( n30476 , n22040 , n28333 );
nand ( n30477 , n22024 , n27506 , n30476 );
not ( n30478 , n30477 );
not ( n30479 , n30478 );
nand ( n30480 , n27501 , n22033 );
not ( n30481 , n30480 );
not ( n30482 , n30481 );
nor ( n30483 , n30479 , n30482 );
not ( n30484 , n30483 );
or ( n30485 , n30475 , n30484 );
or ( n30486 , n30483 , n30474 );
nand ( n30487 , n30485 , n30486 );
buf ( n30488 , n30487 );
and ( n30489 , n30488 , n23673 );
or ( n30490 , n23675 , n12208 );
not ( n30491 , n12153 );
or ( n30492 , n23680 , n30491 );
nand ( n30493 , n30490 , n30492 );
nor ( n30494 , n30489 , n30493 );
and ( n30495 , n30449 , n30473 , n30494 );
or ( n30496 , n30495 , n23706 );
nand ( n30497 , n23708 , n11290 );
nand ( n30498 , n30496 , n30497 );
buf ( n30499 , n30498 );
buf ( n30500 , n30499 );
buf ( n30501 , n275554 );
not ( n30502 , n275929 );
buf ( n30503 , n30502 );
buf ( n30504 , n30503 );
buf ( n30505 , n275554 );
buf ( n30506 , n19562 );
not ( n30507 , n30506 );
or ( n30508 , n30507 , n21770 );
nand ( n30509 , n21774 , n9552 );
nand ( n30510 , n30508 , n30509 );
buf ( n30511 , n30510 );
buf ( n30512 , n30511 );
and ( n30513 , n22904 , n275610 );
nor ( n30514 , n14830 , n17509 );
nor ( n30515 , n30513 , n30514 );
nand ( n30516 , n22914 , n23088 );
buf ( n30517 , n23094 );
not ( n30518 , n30517 );
buf ( n30519 , n23117 );
nand ( n30520 , n30518 , n30519 );
buf ( n30521 , n30520 );
buf ( n30522 , n30521 );
not ( n30523 , n30522 );
buf ( n30524 , n23057 );
not ( n30525 , n30524 );
buf ( n30526 , n23046 );
not ( n30527 , n30526 );
buf ( n30528 , n30527 );
buf ( n30529 , n30528 );
not ( n30530 , n30529 );
or ( n30531 , n30525 , n30530 );
buf ( n30532 , n22984 );
buf ( n30533 , n23057 );
and ( n30534 , n30532 , n30533 );
buf ( n30535 , n22959 );
nor ( n30536 , n30534 , n30535 );
buf ( n30537 , n30536 );
buf ( n30538 , n30537 );
nand ( n30539 , n30531 , n30538 );
buf ( n30540 , n30539 );
buf ( n30541 , n30540 );
not ( n30542 , n30541 );
or ( n30543 , n30523 , n30542 );
buf ( n30544 , n30540 );
buf ( n30545 , n30521 );
or ( n30546 , n30544 , n30545 );
nand ( n30547 , n30543 , n30546 );
buf ( n30548 , n30547 );
buf ( n30549 , n30548 );
nand ( n30550 , n22918 , n30549 );
buf ( n30551 , n23319 );
not ( n30552 , n30551 );
buf ( n30553 , n23342 );
nand ( n30554 , n30552 , n30553 );
buf ( n30555 , n30554 );
buf ( n30556 , n30555 );
not ( n30557 , n30556 );
buf ( n30558 , n23286 );
not ( n30559 , n30558 );
buf ( n30560 , n23275 );
not ( n30561 , n30560 );
buf ( n30562 , n30561 );
buf ( n30563 , n30562 );
not ( n30564 , n30563 );
or ( n30565 , n30559 , n30564 );
buf ( n30566 , n23214 );
buf ( n30567 , n23286 );
and ( n30568 , n30566 , n30567 );
buf ( n30569 , n23191 );
nor ( n30570 , n30568 , n30569 );
buf ( n30571 , n30570 );
buf ( n30572 , n30571 );
nand ( n30573 , n30565 , n30572 );
buf ( n30574 , n30573 );
buf ( n30575 , n30574 );
not ( n30576 , n30575 );
or ( n30577 , n30557 , n30576 );
buf ( n30578 , n30574 );
buf ( n30579 , n30555 );
or ( n30580 , n30578 , n30579 );
nand ( n30581 , n30577 , n30580 );
buf ( n30582 , n30581 );
buf ( n30583 , n30582 );
nand ( n30584 , n23152 , n30583 );
nand ( n30585 , n30515 , n30516 , n30550 , n30584 );
buf ( n30586 , n30585 );
buf ( n30587 , n30586 );
buf ( n30588 , n275554 );
not ( n30589 , n275925 );
buf ( n30590 , n30589 );
buf ( n30591 , n30590 );
not ( n30592 , n275925 );
buf ( n30593 , n30592 );
buf ( n30594 , n30593 );
buf ( n30595 , n275554 );
not ( n30596 , n275929 );
buf ( n30597 , n30596 );
buf ( n30598 , n30597 );
buf ( n30599 , n19539 );
and ( n30600 , n22798 , n30599 );
not ( n30601 , n22798 );
not ( n30602 , n24391 );
nand ( n30603 , n19069 , n22805 );
not ( n30604 , n30603 );
or ( n30605 , n30602 , n30604 );
or ( n30606 , n30603 , n24391 );
nand ( n30607 , n30605 , n30606 );
buf ( n30608 , n30607 );
and ( n30609 , n30601 , n30608 );
nor ( n30610 , n30600 , n30609 );
or ( n30611 , n30610 , n29866 );
not ( n30612 , n19649 );
and ( n30613 , n18374 , n18862 );
not ( n30614 , n18374 );
not ( n30615 , n18862 );
and ( n30616 , n30614 , n30615 );
nor ( n30617 , n30613 , n30616 );
nand ( n30618 , n30612 , n30617 );
nor ( n30619 , n24420 , n20152 );
and ( n30620 , n30619 , n22842 );
not ( n30621 , n30619 );
and ( n30622 , n30621 , n22843 );
nor ( n30623 , n30620 , n30622 );
buf ( n30624 , n30623 );
and ( n30625 , n30624 , n20353 );
buf ( n30626 , n20534 );
buf ( n30627 , n30626 );
buf ( n30628 , n30627 );
not ( n30629 , n30628 );
or ( n30630 , n20562 , n30629 );
and ( n30631 , n20545 , n20535 );
not ( n30632 , n20545 );
and ( n30633 , n30632 , n20536 );
nor ( n30634 , n30631 , n30633 );
buf ( n30635 , n30634 );
not ( n30636 , n30635 );
or ( n30637 , n20559 , n30636 );
not ( n30638 , n18374 );
nor ( n30639 , n30638 , n19639 );
not ( n30640 , n30639 );
nand ( n30641 , n30630 , n30637 , n30640 );
nor ( n30642 , n30625 , n30641 );
nor ( n30643 , n24407 , n20481 );
not ( n30644 , n30643 );
not ( n30645 , n24406 );
or ( n30646 , n30644 , n30645 );
or ( n30647 , n24406 , n30643 );
nand ( n30648 , n30646 , n30647 );
buf ( n30649 , n30648 );
nand ( n30650 , n30649 , n20515 );
and ( n30651 , n30618 , n30642 , n30650 );
nand ( n30652 , n30611 , n30651 );
buf ( n30653 , n30652 );
buf ( n30654 , n30653 );
not ( n30655 , n29517 );
and ( n30656 , n30655 , n21174 );
not ( n30657 , n21001 );
not ( n30658 , n29579 );
or ( n30659 , n30657 , n30658 );
and ( n30660 , n29535 , n19358 );
not ( n30661 , n19290 );
not ( n30662 , n29557 );
or ( n30663 , n30661 , n30662 );
nand ( n30664 , n19219 , n29548 );
nand ( n30665 , n30663 , n30664 );
nor ( n30666 , n30660 , n30665 );
nand ( n30667 , n30659 , n30666 );
nor ( n30668 , n30656 , n30667 );
or ( n30669 , n30668 , n24450 );
nand ( n30670 , n24450 , n18995 );
nand ( n30671 , n30669 , n30670 );
buf ( n30672 , n30671 );
buf ( n30673 , n30672 );
buf ( n30674 , n275554 );
buf ( n30675 , n27312 );
buf ( n30676 , n27395 );
nand ( n30677 , n30675 , n30676 );
buf ( n30678 , n30677 );
buf ( n30679 , n30678 );
not ( n30680 , n30679 );
buf ( n30681 , n23476 );
not ( n30682 , n30681 );
buf ( n30683 , n23515 );
nor ( n30684 , n30682 , n30683 );
buf ( n30685 , n30684 );
buf ( n30686 , n30685 );
not ( n30687 , n30686 );
buf ( n30688 , n23568 );
not ( n30689 , n30688 );
or ( n30690 , n30687 , n30689 );
buf ( n30691 , n23476 );
not ( n30692 , n30691 );
buf ( n30693 , n23587 );
not ( n30694 , n30693 );
or ( n30695 , n30692 , n30694 );
buf ( n30696 , n23481 );
nand ( n30697 , n30695 , n30696 );
buf ( n30698 , n30697 );
buf ( n30699 , n30698 );
not ( n30700 , n30699 );
buf ( n30701 , n30700 );
buf ( n30702 , n30701 );
nand ( n30703 , n30690 , n30702 );
buf ( n30704 , n30703 );
buf ( n30705 , n30704 );
not ( n30706 , n30705 );
or ( n30707 , n30680 , n30706 );
buf ( n30708 , n30704 );
buf ( n30709 , n30678 );
or ( n30710 , n30708 , n30709 );
nand ( n30711 , n30707 , n30710 );
buf ( n30712 , n30711 );
buf ( n30713 , n30712 );
nand ( n30714 , n30713 , n27489 );
nand ( n30715 , n27208 , n27238 );
not ( n30716 , n30715 );
not ( n30717 , n23608 );
nor ( n30718 , n30717 , n23621 );
not ( n30719 , n30718 );
not ( n30720 , n28417 );
or ( n30721 , n30719 , n30720 );
not ( n30722 , n23608 );
not ( n30723 , n23647 );
or ( n30724 , n30722 , n30723 );
nand ( n30725 , n30724 , n23610 );
not ( n30726 , n30725 );
nand ( n30727 , n30721 , n30726 );
not ( n30728 , n30727 );
or ( n30729 , n30716 , n30728 );
or ( n30730 , n30727 , n30715 );
nand ( n30731 , n30729 , n30730 );
buf ( n30732 , n30731 );
nand ( n30733 , n30732 , n23655 );
not ( n30734 , n28337 );
not ( n30735 , n30734 );
buf ( n30736 , n28336 );
not ( n30737 , n30736 );
or ( n30738 , n30735 , n30737 );
or ( n30739 , n30736 , n30734 );
nand ( n30740 , n30738 , n30739 );
buf ( n30741 , n30740 );
and ( n30742 , n30741 , n23673 );
not ( n30743 , n12255 );
or ( n30744 , n23675 , n30743 );
or ( n30745 , n23680 , n12240 );
nand ( n30746 , n30744 , n30745 );
nor ( n30747 , n30742 , n30746 );
and ( n30748 , n30714 , n30733 , n30747 );
or ( n30749 , n30748 , n23706 );
nand ( n30750 , n23708 , n11467 );
nand ( n30751 , n30749 , n30750 );
buf ( n30752 , n30751 );
buf ( n30753 , n30752 );
buf ( n30754 , n275554 );
buf ( n30755 , n275554 );
buf ( n30756 , n275554 );
not ( n30757 , n275929 );
buf ( n30758 , n30757 );
buf ( n30759 , n30758 );
buf ( n30760 , n275554 );
buf ( n30761 , n275554 );
buf ( n30762 , n275554 );
not ( n30763 , n275925 );
buf ( n30764 , n30763 );
buf ( n30765 , n30764 );
not ( n30766 , n275929 );
buf ( n30767 , n30766 );
buf ( n30768 , n30767 );
not ( n30769 , n275550 );
buf ( n30770 , n30769 );
buf ( n30771 , n30770 );
buf ( n30772 , n275554 );
not ( n30773 , n275929 );
buf ( n30774 , n30773 );
buf ( n30775 , n30774 );
not ( n30776 , n14056 );
or ( n30777 , n30776 , n29046 );
nand ( n30778 , n29044 , n9748 );
nand ( n30779 , n30777 , n30778 );
buf ( n30780 , n30779 );
buf ( n30781 , n30780 );
not ( n30782 , n275929 );
buf ( n30783 , n30782 );
buf ( n30784 , n30783 );
buf ( n30785 , n275554 );
buf ( n30786 , n275554 );
not ( n30787 , n275929 );
buf ( n30788 , n30787 );
buf ( n30789 , n30788 );
and ( n30790 , n22193 , n277753 );
not ( n30791 , n22193 );
not ( n30792 , n29599 );
buf ( n30793 , n277775 );
buf ( n30794 , n30793 );
buf ( n30795 , n277798 );
buf ( n30796 , n30795 );
or ( n30797 , n30794 , n30796 );
buf ( n30798 , n30797 );
buf ( n30799 , n30798 );
buf ( n30800 , n30793 );
buf ( n30801 , n30795 );
and ( n30802 , n30800 , n30801 );
buf ( n30803 , n30802 );
buf ( n30804 , n30803 );
not ( n30805 , n30804 );
buf ( n30806 , n30805 );
buf ( n30807 , n30806 );
nand ( n30808 , n30799 , n30807 );
buf ( n30809 , n30808 );
buf ( n30810 , n30809 );
not ( n30811 , n30810 );
buf ( n30812 , n29610 );
buf ( n30813 , n29633 );
and ( n30814 , n30812 , n30813 );
buf ( n30815 , n30814 );
buf ( n30816 , n30815 );
not ( n30817 , n30816 );
buf ( n30818 , n29652 );
nor ( n30819 , n30817 , n30818 );
buf ( n30820 , n30819 );
buf ( n30821 , n30820 );
not ( n30822 , n30821 );
buf ( n30823 , n30822 );
buf ( n30824 , n30823 );
buf ( n30825 , n277842 );
buf ( n30826 , n30825 );
buf ( n30827 , n277822 );
buf ( n30828 , n30827 );
or ( n30829 , n30826 , n30828 );
buf ( n30830 , n30829 );
buf ( n30831 , n30830 );
buf ( n30832 , n277896 );
buf ( n30833 , n30832 );
buf ( n30834 , n277872 );
buf ( n30835 , n30834 );
or ( n30836 , n30833 , n30835 );
buf ( n30837 , n30836 );
buf ( n30838 , n30837 );
nand ( n30839 , n30831 , n30838 );
buf ( n30840 , n30839 );
buf ( n30841 , n30840 );
nor ( n30842 , n30824 , n30841 );
buf ( n30843 , n30842 );
buf ( n30844 , n30843 );
not ( n30845 , n30844 );
buf ( n30846 , n27479 );
not ( n30847 , n30846 );
or ( n30848 , n30845 , n30847 );
buf ( n30849 , n30840 );
not ( n30850 , n30849 );
buf ( n30851 , n29674 );
not ( n30852 , n30851 );
buf ( n30853 , n30815 );
not ( n30854 , n30853 );
or ( n30855 , n30852 , n30854 );
buf ( n30856 , n29681 );
not ( n30857 , n30856 );
buf ( n30858 , n29610 );
not ( n30859 , n30858 );
or ( n30860 , n30857 , n30859 );
buf ( n30861 , n29616 );
nand ( n30862 , n30860 , n30861 );
buf ( n30863 , n30862 );
buf ( n30864 , n30863 );
not ( n30865 , n30864 );
buf ( n30866 , n30865 );
buf ( n30867 , n30866 );
nand ( n30868 , n30855 , n30867 );
buf ( n30869 , n30868 );
buf ( n30870 , n30869 );
nand ( n30871 , n30850 , n30870 );
buf ( n30872 , n30871 );
buf ( n30873 , n30872 );
not ( n30874 , n30873 );
buf ( n30875 , n30825 );
buf ( n30876 , n30827 );
nand ( n30877 , n30875 , n30876 );
buf ( n30878 , n30877 );
buf ( n30879 , n30878 );
not ( n30880 , n30879 );
buf ( n30881 , n30837 );
nand ( n30882 , n30880 , n30881 );
buf ( n30883 , n30882 );
buf ( n30884 , n30883 );
buf ( n30885 , n30834 );
buf ( n30886 , n30832 );
nand ( n30887 , n30885 , n30886 );
buf ( n30888 , n30887 );
buf ( n30889 , n30888 );
nand ( n30890 , n30884 , n30889 );
buf ( n30891 , n30890 );
buf ( n30892 , n30891 );
nor ( n30893 , n30874 , n30892 );
buf ( n30894 , n30893 );
buf ( n30895 , n30894 );
nand ( n30896 , n30848 , n30895 );
buf ( n30897 , n30896 );
buf ( n30898 , n30897 );
not ( n30899 , n30898 );
or ( n30900 , n30811 , n30899 );
buf ( n30901 , n30897 );
buf ( n30902 , n30809 );
or ( n30903 , n30901 , n30902 );
nand ( n30904 , n30900 , n30903 );
buf ( n30905 , n30904 );
buf ( n30906 , n30905 );
not ( n30907 , n30906 );
or ( n30908 , n30792 , n30907 );
buf ( n30909 , n277775 );
not ( n30910 , n30909 );
buf ( n30911 , n277798 );
nand ( n30912 , n30910 , n30911 );
not ( n30913 , n30912 );
not ( n30914 , n30909 );
nor ( n30915 , n30914 , n30911 );
or ( n30916 , n30913 , n30915 );
not ( n30917 , n30916 );
buf ( n30918 , n277842 );
not ( n30919 , n30918 );
buf ( n30920 , n277822 );
nand ( n30921 , n30919 , n30920 );
buf ( n30922 , n277872 );
not ( n30923 , n30922 );
buf ( n30924 , n277896 );
nand ( n30925 , n30923 , n30924 );
nand ( n30926 , n30921 , n30925 );
not ( n30927 , n30926 );
not ( n30928 , n30927 );
and ( n30929 , n29708 , n29716 );
not ( n30930 , n30929 );
nor ( n30931 , n30930 , n29724 );
not ( n30932 , n30931 );
nor ( n30933 , n30928 , n30932 );
not ( n30934 , n30933 );
not ( n30935 , n29728 );
or ( n30936 , n30934 , n30935 );
not ( n30937 , n29736 );
not ( n30938 , n30929 );
or ( n30939 , n30937 , n30938 );
not ( n30940 , n29739 );
not ( n30941 , n29708 );
or ( n30942 , n30940 , n30941 );
nand ( n30943 , n30942 , n29710 );
not ( n30944 , n30943 );
nand ( n30945 , n30939 , n30944 );
nand ( n30946 , n30945 , n30927 );
not ( n30947 , n30946 );
not ( n30948 , n30920 );
nand ( n30949 , n30948 , n30918 );
not ( n30950 , n30949 );
nand ( n30951 , n30950 , n30925 );
not ( n30952 , n30924 );
nand ( n30953 , n30952 , n30922 );
nand ( n30954 , n30951 , n30953 );
nor ( n30955 , n30947 , n30954 );
nand ( n30956 , n30936 , n30955 );
not ( n30957 , n30956 );
or ( n30958 , n30917 , n30957 );
or ( n30959 , n30956 , n30916 );
nand ( n30960 , n30958 , n30959 );
buf ( n30961 , n30960 );
buf ( n30962 , n27266 );
and ( n30963 , n30961 , n30962 );
not ( n30964 , n23673 );
buf ( n30965 , n277717 );
not ( n30966 , n30965 );
not ( n30967 , n30966 );
not ( n30968 , n30482 );
nand ( n30969 , n29754 , n27502 );
buf ( n30970 , n30969 );
buf ( n30971 , n277775 );
buf ( n30972 , n30971 );
nand ( n30973 , n27492 , n30972 );
nor ( n30974 , n30970 , n30973 );
not ( n30975 , n29756 );
buf ( n30976 , n277872 );
not ( n30977 , n30976 );
nor ( n30978 , n29751 , n30975 , n30977 );
buf ( n30979 , n30978 );
nand ( n30980 , n30974 , n30979 );
nor ( n30981 , n27511 , n30980 );
nand ( n30982 , n30968 , n30981 );
not ( n30983 , n30982 );
not ( n30984 , n30983 );
or ( n30985 , n30967 , n30984 );
or ( n30986 , n30983 , n30966 );
nand ( n30987 , n30985 , n30986 );
buf ( n30988 , n30987 );
not ( n30989 , n30988 );
or ( n30990 , n30964 , n30989 );
and ( n30991 , n27520 , n12185 );
and ( n30992 , n22013 , n12370 );
nor ( n30993 , n30991 , n30992 );
nand ( n30994 , n30990 , n30993 );
nor ( n30995 , n30963 , n30994 );
nand ( n30996 , n30908 , n30995 );
and ( n30997 , n30791 , n30996 );
or ( n30998 , n30790 , n30997 );
buf ( n30999 , n30998 );
buf ( n31000 , n30999 );
not ( n31001 , n275925 );
buf ( n31002 , n31001 );
buf ( n31003 , n31002 );
nand ( n31004 , n28213 , n22000 );
not ( n31005 , n22056 );
nand ( n31006 , n28194 , n31005 );
not ( n31007 , n22012 );
nand ( n31008 , n31007 , n12141 );
and ( n31009 , n31004 , n31006 , n31008 );
nand ( n31010 , n28228 , n23672 );
nand ( n31011 , n22007 , n12318 );
nand ( n31012 , n31009 , n31010 , n31011 );
not ( n31013 , n31012 );
or ( n31014 , n31013 , n27589 );
or ( n31015 , n22191 , n11002 );
nand ( n31016 , n31014 , n31015 );
buf ( n31017 , n31016 );
buf ( n31018 , n31017 );
not ( n31019 , n275925 );
buf ( n31020 , n31019 );
buf ( n31021 , n31020 );
not ( n31022 , n26091 );
not ( n31023 , n22335 );
or ( n31024 , n31022 , n31023 );
nand ( n31025 , n20238 , n275557 );
nand ( n31026 , n31024 , n31025 );
buf ( n31027 , n31026 );
buf ( n31028 , n31027 );
not ( n31029 , n275929 );
buf ( n31030 , n31029 );
buf ( n31031 , n31030 );
buf ( n31032 , n275554 );
buf ( n31033 , n275554 );
not ( n31034 , n275929 );
buf ( n31035 , n31034 );
buf ( n31036 , n31035 );
not ( n31037 , n275550 );
buf ( n31038 , n31037 );
buf ( n31039 , n31038 );
not ( n31040 , n26597 );
not ( n31041 , n31040 );
and ( n31042 , n26516 , n31041 );
not ( n31043 , n26516 );
buf ( n31044 , n26581 );
not ( n31045 , n31044 );
not ( n31046 , n29403 );
not ( n31047 , n26631 );
nor ( n31048 , n29826 , n31047 );
nand ( n31049 , n31046 , n31048 );
not ( n31050 , n31049 );
or ( n31051 , n31045 , n31050 );
or ( n31052 , n31049 , n31044 );
nand ( n31053 , n31051 , n31052 );
buf ( n31054 , n31053 );
and ( n31055 , n31043 , n31054 );
nor ( n31056 , n31042 , n31055 );
or ( n31057 , n31056 , n19634 );
not ( n31058 , n27012 );
nand ( n31059 , n31058 , n27038 );
not ( n31060 , n31059 );
nor ( n31061 , n26991 , n27003 );
not ( n31062 , n31061 );
not ( n31063 , n27020 );
or ( n31064 , n31062 , n31063 );
not ( n31065 , n27003 );
not ( n31066 , n31065 );
not ( n31067 , n27034 );
or ( n31068 , n31066 , n31067 );
nand ( n31069 , n31068 , n27036 );
not ( n31070 , n31069 );
nand ( n31071 , n31064 , n31070 );
not ( n31072 , n31071 );
or ( n31073 , n31060 , n31072 );
or ( n31074 , n31071 , n31059 );
nand ( n31075 , n31073 , n31074 );
buf ( n31076 , n31075 );
and ( n31077 , n31076 , n29471 );
not ( n31078 , n18818 );
not ( n31079 , n31078 );
not ( n31080 , n30140 );
or ( n31081 , n31079 , n31080 );
or ( n31082 , n30140 , n31078 );
nand ( n31083 , n31081 , n31082 );
not ( n31084 , n31083 );
not ( n31085 , n30612 );
or ( n31086 , n31084 , n31085 );
not ( n31087 , n27068 );
nor ( n31088 , n27065 , n27070 );
nand ( n31089 , n24314 , n31088 );
not ( n31090 , n31089 );
or ( n31091 , n31087 , n31090 );
or ( n31092 , n31089 , n27068 );
nand ( n31093 , n31091 , n31092 );
buf ( n31094 , n31093 );
not ( n31095 , n20559 );
nand ( n31096 , n31094 , n31095 );
buf ( n31097 , n27066 );
buf ( n31098 , n31097 );
nand ( n31099 , n20563 , n31098 );
nand ( n31100 , n30179 , n18819 );
and ( n31101 , n31096 , n31099 , n31100 );
nand ( n31102 , n31086 , n31101 );
nor ( n31103 , n31077 , n31102 );
not ( n31104 , n26899 );
nand ( n31105 , n31104 , n26933 );
not ( n31106 , n31105 );
not ( n31107 , n26911 );
nor ( n31108 , n31107 , n26853 );
not ( n31109 , n31108 );
not ( n31110 , n26915 );
or ( n31111 , n31109 , n31110 );
not ( n31112 , n26911 );
not ( n31113 , n26928 );
or ( n31114 , n31112 , n31113 );
nand ( n31115 , n31114 , n26931 );
not ( n31116 , n31115 );
nand ( n31117 , n31111 , n31116 );
not ( n31118 , n31117 );
or ( n31119 , n31106 , n31118 );
or ( n31120 , n31117 , n31105 );
nand ( n31121 , n31119 , n31120 );
buf ( n31122 , n31121 );
nand ( n31123 , n31122 , n20353 );
and ( n31124 , n31103 , n31123 );
nand ( n31125 , n31057 , n31124 );
buf ( n31126 , n31125 );
buf ( n31127 , n31126 );
buf ( n31128 , n275554 );
buf ( n31129 , n275554 );
not ( n31130 , n20672 );
not ( n31131 , n20724 );
not ( n31132 , n23390 );
not ( n31133 , n31132 );
or ( n31134 , n31131 , n31133 );
or ( n31135 , n31132 , n20724 );
nand ( n31136 , n31134 , n31135 );
buf ( n31137 , n31136 );
not ( n31138 , n31137 );
or ( n31139 , n31130 , n31138 );
buf ( n31140 , n14131 );
nand ( n31141 , n31140 , n13373 );
nand ( n31142 , n31139 , n31141 );
not ( n31143 , n31142 );
or ( n31144 , n31143 , n26364 );
nand ( n31145 , n15907 , n23412 );
not ( n31146 , n31145 );
not ( n31147 , n16913 );
or ( n31148 , n31146 , n31147 );
buf ( n31149 , n16913 );
or ( n31150 , n31149 , n31145 );
nand ( n31151 , n31148 , n31150 );
buf ( n31152 , n31151 );
nand ( n31153 , n31152 , n26370 );
nand ( n31154 , n23424 , n17378 );
not ( n31155 , n31154 );
not ( n31156 , n17362 );
or ( n31157 , n31155 , n31156 );
buf ( n31158 , n17362 );
or ( n31159 , n31158 , n31154 );
nand ( n31160 , n31157 , n31159 );
buf ( n31161 , n31160 );
nand ( n31162 , n31161 , n26374 );
not ( n31163 , n17470 );
not ( n31164 , n23436 );
or ( n31165 , n31163 , n31164 );
not ( n31166 , n17463 );
or ( n31167 , n31166 , n17470 );
nand ( n31168 , n31165 , n31167 );
buf ( n31169 , n31168 );
nand ( n31170 , n31169 , n26393 );
buf ( n31171 , n17469 );
buf ( n31172 , n31171 );
not ( n31173 , n31172 );
not ( n31174 , n31173 );
nand ( n31175 , n26395 , n31174 );
not ( n31176 , n13769 );
nor ( n31177 , n26386 , n31176 );
not ( n31178 , n31177 );
and ( n31179 , n31170 , n31175 , n31178 );
not ( n31180 , n26390 );
and ( n31181 , n17521 , n13770 );
not ( n31182 , n17521 );
and ( n31183 , n31182 , n31176 );
nor ( n31184 , n31181 , n31183 );
nand ( n31185 , n31180 , n31184 );
and ( n31186 , n31153 , n31162 , n31179 , n31185 );
nand ( n31187 , n31144 , n31186 );
buf ( n31188 , n31187 );
buf ( n31189 , n31188 );
buf ( n31190 , n275554 );
not ( n31191 , n275925 );
buf ( n31192 , n31191 );
buf ( n31193 , n31192 );
not ( n31194 , n275925 );
buf ( n31195 , n31194 );
buf ( n31196 , n31195 );
nand ( n31197 , n25064 , n25164 );
buf ( n31198 , n25170 );
not ( n31199 , n31198 );
buf ( n31200 , n25233 );
nand ( n31201 , n31199 , n31200 );
buf ( n31202 , n31201 );
buf ( n31203 , n31202 );
not ( n31204 , n31203 );
buf ( n31205 , n25221 );
not ( n31206 , n31205 );
or ( n31207 , n31204 , n31206 );
buf ( n31208 , n25221 );
buf ( n31209 , n31202 );
or ( n31210 , n31208 , n31209 );
nand ( n31211 , n31207 , n31210 );
buf ( n31212 , n31211 );
buf ( n31213 , n31212 );
not ( n31214 , n31213 );
nor ( n31215 , n31214 , n25389 );
nand ( n31216 , n25397 , n275787 );
buf ( n31217 , n25554 );
not ( n31218 , n31217 );
buf ( n31219 , n25491 );
nor ( n31220 , n31218 , n31219 );
buf ( n31221 , n31220 );
buf ( n31222 , n31221 );
not ( n31223 , n31222 );
buf ( n31224 , n25540 );
not ( n31225 , n31224 );
buf ( n31226 , n31225 );
buf ( n31227 , n31226 );
not ( n31228 , n31227 );
or ( n31229 , n31223 , n31228 );
buf ( n31230 , n31226 );
buf ( n31231 , n31221 );
or ( n31232 , n31230 , n31231 );
nand ( n31233 , n31229 , n31232 );
buf ( n31234 , n31233 );
buf ( n31235 , n31234 );
and ( n31236 , n25402 , n31235 );
nor ( n31237 , n31236 , n30639 );
buf ( n31238 , n25870 );
not ( n31239 , n31238 );
buf ( n31240 , n25807 );
nor ( n31241 , n31239 , n31240 );
buf ( n31242 , n31241 );
buf ( n31243 , n31242 );
not ( n31244 , n31243 );
buf ( n31245 , n25856 );
not ( n31246 , n31245 );
buf ( n31247 , n31246 );
buf ( n31248 , n31247 );
not ( n31249 , n31248 );
or ( n31250 , n31244 , n31249 );
buf ( n31251 , n31247 );
buf ( n31252 , n31242 );
or ( n31253 , n31251 , n31252 );
nand ( n31254 , n31250 , n31253 );
buf ( n31255 , n31254 );
buf ( n31256 , n31255 );
nand ( n31257 , n25717 , n31256 );
nand ( n31258 , n31216 , n31237 , n31257 );
nor ( n31259 , n31215 , n31258 );
buf ( n31260 , n26180 );
not ( n31261 , n31260 );
buf ( n31262 , n26116 );
nor ( n31263 , n31261 , n31262 );
buf ( n31264 , n31263 );
buf ( n31265 , n31264 );
not ( n31266 , n31265 );
buf ( n31267 , n26166 );
not ( n31268 , n31267 );
buf ( n31269 , n31268 );
buf ( n31270 , n31269 );
not ( n31271 , n31270 );
or ( n31272 , n31266 , n31271 );
buf ( n31273 , n31269 );
buf ( n31274 , n31264 );
or ( n31275 , n31273 , n31274 );
nand ( n31276 , n31272 , n31275 );
buf ( n31277 , n31276 );
buf ( n31278 , n31277 );
nand ( n31279 , n26027 , n31278 );
nand ( n31280 , n31197 , n31259 , n31279 );
buf ( n31281 , n31280 );
buf ( n31282 , n31281 );
not ( n31283 , n275929 );
buf ( n31284 , n31283 );
buf ( n31285 , n31284 );
buf ( n31286 , n275554 );
buf ( n31287 , n275554 );
not ( n31288 , n275925 );
buf ( n31289 , n31288 );
buf ( n31290 , n31289 );
not ( n31291 , n23386 );
not ( n31292 , n20723 );
and ( n31293 , n23778 , n20722 );
buf ( n31294 , n14405 );
nand ( n31295 , n31293 , n31294 );
not ( n31296 , n31295 );
or ( n31297 , n31292 , n31296 );
or ( n31298 , n31295 , n20723 );
nand ( n31299 , n31297 , n31298 );
buf ( n31300 , n31299 );
not ( n31301 , n31300 );
or ( n31302 , n31291 , n31301 );
buf ( n31303 , n14184 );
not ( n31304 , n23386 );
nand ( n31305 , n31303 , n31304 );
nand ( n31306 , n31302 , n31305 );
not ( n31307 , n31306 );
or ( n31308 , n31307 , n20743 );
nand ( n31309 , n17087 , n17369 );
not ( n31310 , n31309 );
not ( n31311 , n20747 );
not ( n31312 , n31311 );
not ( n31313 , n17362 );
or ( n31314 , n31312 , n31313 );
nand ( n31315 , n31314 , n20753 );
not ( n31316 , n31315 );
or ( n31317 , n31310 , n31316 );
or ( n31318 , n31315 , n31309 );
nand ( n31319 , n31317 , n31318 );
buf ( n31320 , n31319 );
and ( n31321 , n20763 , n31320 );
nand ( n31322 , n23436 , n20775 );
and ( n31323 , n31322 , n17467 );
not ( n31324 , n31322 );
and ( n31325 , n31324 , n20776 );
nor ( n31326 , n31323 , n31325 );
buf ( n31327 , n31326 );
nand ( n31328 , n17411 , n31327 );
buf ( n31329 , n17466 );
buf ( n31330 , n31329 );
not ( n31331 , n31330 );
not ( n31332 , n31331 );
nand ( n31333 , n20785 , n31332 );
nand ( n31334 , n17560 , n13920 );
and ( n31335 , n17527 , n13910 );
not ( n31336 , n17527 );
not ( n31337 , n13909 );
and ( n31338 , n31336 , n31337 );
nor ( n31339 , n31335 , n31338 );
nand ( n31340 , n17545 , n31339 );
nand ( n31341 , n31328 , n31333 , n31334 , n31340 );
nor ( n31342 , n31321 , n31341 );
not ( n31343 , n20797 );
nand ( n31344 , n31343 , n16930 );
not ( n31345 , n31344 );
not ( n31346 , n20796 );
not ( n31347 , n31346 );
not ( n31348 , n16913 );
or ( n31349 , n31347 , n31348 );
buf ( n31350 , n20804 );
nand ( n31351 , n31349 , n31350 );
not ( n31352 , n31351 );
or ( n31353 , n31345 , n31352 );
or ( n31354 , n31351 , n31344 );
nand ( n31355 , n31353 , n31354 );
buf ( n31356 , n31355 );
nand ( n31357 , n31356 , n16970 );
and ( n31358 , n31342 , n31357 );
nand ( n31359 , n31308 , n31358 );
buf ( n31360 , n31359 );
buf ( n31361 , n31360 );
not ( n31362 , n275550 );
buf ( n31363 , n31362 );
buf ( n31364 , n31363 );
buf ( n31365 , n275554 );
not ( n31366 , n275550 );
buf ( n31367 , n31366 );
buf ( n31368 , n31367 );
not ( n31369 , n275550 );
buf ( n31370 , n31369 );
buf ( n31371 , n31370 );
not ( n31372 , n275550 );
buf ( n31373 , n31372 );
buf ( n31374 , n31373 );
buf ( n31375 , n275554 );
buf ( n31376 , n275554 );
buf ( n31377 , n275554 );
not ( n31378 , n275929 );
buf ( n31379 , n31378 );
buf ( n31380 , n31379 );
not ( n31381 , n275550 );
buf ( n31382 , n31381 );
buf ( n31383 , n31382 );
buf ( n31384 , n275554 );
not ( n31385 , n275929 );
buf ( n31386 , n31385 );
buf ( n31387 , n31386 );
not ( n31388 , n275550 );
buf ( n31389 , n31388 );
buf ( n31390 , n31389 );
buf ( n31391 , n275554 );
buf ( n31392 , n29684 );
buf ( n31393 , n29634 );
nand ( n31394 , n31392 , n31393 );
buf ( n31395 , n31394 );
buf ( n31396 , n31395 );
not ( n31397 , n31396 );
buf ( n31398 , n29652 );
not ( n31399 , n31398 );
buf ( n31400 , n31399 );
buf ( n31401 , n31400 );
not ( n31402 , n31401 );
buf ( n31403 , n27479 );
not ( n31404 , n31403 );
or ( n31405 , n31402 , n31404 );
buf ( n31406 , n29674 );
not ( n31407 , n31406 );
buf ( n31408 , n31407 );
buf ( n31409 , n31408 );
nand ( n31410 , n31405 , n31409 );
buf ( n31411 , n31410 );
buf ( n31412 , n31411 );
not ( n31413 , n31412 );
or ( n31414 , n31397 , n31413 );
buf ( n31415 , n31411 );
buf ( n31416 , n31395 );
or ( n31417 , n31415 , n31416 );
nand ( n31418 , n31414 , n31417 );
buf ( n31419 , n31418 );
buf ( n31420 , n31419 );
not ( n31421 , n28306 );
not ( n31422 , n31421 );
nand ( n31423 , n31420 , n31422 );
nand ( n31424 , n29717 , n29740 );
not ( n31425 , n31424 );
not ( n31426 , n29725 );
not ( n31427 , n31426 );
not ( n31428 , n29728 );
or ( n31429 , n31427 , n31428 );
not ( n31430 , n29736 );
nand ( n31431 , n31429 , n31430 );
not ( n31432 , n31431 );
or ( n31433 , n31425 , n31432 );
or ( n31434 , n31431 , n31424 );
nand ( n31435 , n31433 , n31434 );
buf ( n31436 , n31435 );
not ( n31437 , n28329 );
nand ( n31438 , n31436 , n31437 );
not ( n31439 , n30975 );
not ( n31440 , n29755 );
buf ( n31441 , n29753 );
nor ( n31442 , n31440 , n31441 );
not ( n31443 , n31442 );
or ( n31444 , n31439 , n31443 );
or ( n31445 , n31442 , n30975 );
nand ( n31446 , n31444 , n31445 );
buf ( n31447 , n31446 );
buf ( n31448 , n28218 );
not ( n31449 , n31448 );
nand ( n31450 , n31447 , n31449 );
not ( n31451 , n28230 );
and ( n31452 , n31451 , n12294 );
buf ( n31453 , n28233 );
not ( n31454 , n277933 );
or ( n31455 , n31453 , n31454 );
nand ( n31456 , n28236 , n277941 );
nand ( n31457 , n31455 , n31456 );
nor ( n31458 , n31452 , n31457 );
not ( n31459 , n28241 );
buf ( n31460 , n31459 );
nand ( n31461 , n31460 , n12357 );
and ( n31462 , n31450 , n31458 , n31461 );
nand ( n31463 , n31423 , n31438 , n31462 );
buf ( n31464 , n31463 );
buf ( n31465 , n31464 );
buf ( n31466 , n275554 );
not ( n31467 , n22904 );
not ( n31468 , n31467 );
and ( n31469 , n31468 , n275571 );
nor ( n31470 , n14830 , n17520 );
nor ( n31471 , n31469 , n31470 );
nand ( n31472 , n22914 , n23805 );
buf ( n31473 , n23805 );
buf ( n31474 , n31473 );
buf ( n31475 , n13501 );
buf ( n31476 , n31475 );
nand ( n31477 , n31474 , n31476 );
buf ( n31478 , n31477 );
buf ( n31479 , n31478 );
not ( n31480 , n31479 );
buf ( n31481 , n31473 );
buf ( n31482 , n31475 );
nor ( n31483 , n31481 , n31482 );
buf ( n31484 , n31483 );
buf ( n31485 , n31484 );
nor ( n31486 , n31480 , n31485 );
buf ( n31487 , n31486 );
buf ( n31488 , n31487 );
not ( n31489 , n31488 );
buf ( n31490 , n23078 );
buf ( n31491 , n23097 );
and ( n31492 , n31490 , n31491 );
buf ( n31493 , n31492 );
buf ( n31494 , n31493 );
buf ( n31495 , n30540 );
buf ( n31496 , n13205 );
buf ( n31497 , n31496 );
buf ( n31498 , n31497 );
buf ( n31499 , n13689 );
buf ( n31500 , n31499 );
nor ( n31501 , n31498 , n31500 );
buf ( n31502 , n31501 );
buf ( n31503 , n31502 );
buf ( n31504 , n22924 );
nor ( n31505 , n31503 , n31504 );
buf ( n31506 , n31505 );
buf ( n31507 , n31506 );
buf ( n31508 , n13189 );
buf ( n31509 , n31508 );
buf ( n31510 , n31509 );
buf ( n31511 , n13517 );
buf ( n31512 , n31511 );
nor ( n31513 , n31510 , n31512 );
buf ( n31514 , n31513 );
buf ( n31515 , n31514 );
not ( n31516 , n31515 );
buf ( n31517 , n31516 );
buf ( n31518 , n31517 );
and ( n31519 , n31507 , n31518 );
buf ( n31520 , n31519 );
buf ( n31521 , n31520 );
and ( n31522 , n31494 , n31495 , n31521 );
buf ( n31523 , n31520 );
not ( n31524 , n31523 );
buf ( n31525 , n23137 );
not ( n31526 , n31525 );
or ( n31527 , n31524 , n31526 );
buf ( n31528 , n31502 );
buf ( n31529 , n22930 );
or ( n31530 , n31528 , n31529 );
buf ( n31531 , n31497 );
buf ( n31532 , n31499 );
nand ( n31533 , n31531 , n31532 );
buf ( n31534 , n31533 );
buf ( n31535 , n31534 );
nand ( n31536 , n31530 , n31535 );
buf ( n31537 , n31536 );
buf ( n31538 , n31537 );
buf ( n31539 , n31517 );
and ( n31540 , n31538 , n31539 );
buf ( n31541 , n31509 );
buf ( n31542 , n31511 );
nand ( n31543 , n31541 , n31542 );
buf ( n31544 , n31543 );
buf ( n31545 , n31544 );
not ( n31546 , n31545 );
buf ( n31547 , n31546 );
buf ( n31548 , n31547 );
nor ( n31549 , n31540 , n31548 );
buf ( n31550 , n31549 );
buf ( n31551 , n31550 );
nand ( n31552 , n31527 , n31551 );
buf ( n31553 , n31552 );
buf ( n31554 , n31553 );
nor ( n31555 , n31522 , n31554 );
buf ( n31556 , n31555 );
buf ( n31557 , n31556 );
not ( n31558 , n31557 );
or ( n31559 , n31489 , n31558 );
buf ( n31560 , n31556 );
buf ( n31561 , n31487 );
or ( n31562 , n31560 , n31561 );
nand ( n31563 , n31559 , n31562 );
buf ( n31564 , n31563 );
buf ( n31565 , n31564 );
nand ( n31566 , n22918 , n31565 );
buf ( n31567 , n23805 );
buf ( n31568 , n31567 );
buf ( n31569 , n13495 );
buf ( n31570 , n31569 );
nand ( n31571 , n31568 , n31570 );
buf ( n31572 , n31571 );
buf ( n31573 , n31572 );
not ( n31574 , n31573 );
buf ( n31575 , n31567 );
buf ( n31576 , n31569 );
nor ( n31577 , n31575 , n31576 );
buf ( n31578 , n31577 );
buf ( n31579 , n31578 );
nor ( n31580 , n31574 , n31579 );
buf ( n31581 , n31580 );
buf ( n31582 , n31581 );
not ( n31583 , n31582 );
buf ( n31584 , n23305 );
buf ( n31585 , n23322 );
and ( n31586 , n31584 , n31585 );
buf ( n31587 , n31586 );
buf ( n31588 , n31587 );
buf ( n31589 , n30574 );
buf ( n31590 , n31496 );
buf ( n31591 , n31590 );
buf ( n31592 , n13695 );
buf ( n31593 , n31592 );
nor ( n31594 , n31591 , n31593 );
buf ( n31595 , n31594 );
buf ( n31596 , n31595 );
buf ( n31597 , n23158 );
nor ( n31598 , n31596 , n31597 );
buf ( n31599 , n31598 );
buf ( n31600 , n31599 );
buf ( n31601 , n31508 );
buf ( n31602 , n31601 );
buf ( n31603 , n13522 );
buf ( n31604 , n31603 );
nor ( n31605 , n31602 , n31604 );
buf ( n31606 , n31605 );
buf ( n31607 , n31606 );
not ( n31608 , n31607 );
buf ( n31609 , n31608 );
buf ( n31610 , n31609 );
and ( n31611 , n31600 , n31610 );
buf ( n31612 , n31611 );
buf ( n31613 , n31612 );
and ( n31614 , n31588 , n31589 , n31613 );
buf ( n31615 , n31612 );
not ( n31616 , n31615 );
buf ( n31617 , n23362 );
not ( n31618 , n31617 );
or ( n31619 , n31616 , n31618 );
buf ( n31620 , n31595 );
buf ( n31621 , n23164 );
or ( n31622 , n31620 , n31621 );
buf ( n31623 , n31590 );
buf ( n31624 , n31592 );
nand ( n31625 , n31623 , n31624 );
buf ( n31626 , n31625 );
buf ( n31627 , n31626 );
nand ( n31628 , n31622 , n31627 );
buf ( n31629 , n31628 );
buf ( n31630 , n31629 );
buf ( n31631 , n31609 );
and ( n31632 , n31630 , n31631 );
buf ( n31633 , n31601 );
buf ( n31634 , n31603 );
nand ( n31635 , n31633 , n31634 );
buf ( n31636 , n31635 );
buf ( n31637 , n31636 );
not ( n31638 , n31637 );
buf ( n31639 , n31638 );
buf ( n31640 , n31639 );
nor ( n31641 , n31632 , n31640 );
buf ( n31642 , n31641 );
buf ( n31643 , n31642 );
nand ( n31644 , n31619 , n31643 );
buf ( n31645 , n31644 );
buf ( n31646 , n31645 );
nor ( n31647 , n31614 , n31646 );
buf ( n31648 , n31647 );
buf ( n31649 , n31648 );
not ( n31650 , n31649 );
or ( n31651 , n31583 , n31650 );
buf ( n31652 , n31648 );
buf ( n31653 , n31581 );
or ( n31654 , n31652 , n31653 );
nand ( n31655 , n31651 , n31654 );
buf ( n31656 , n31655 );
buf ( n31657 , n31656 );
nand ( n31658 , n23152 , n31657 );
nand ( n31659 , n31471 , n31472 , n31566 , n31658 );
buf ( n31660 , n31659 );
buf ( n31661 , n31660 );
buf ( n31662 , n275554 );
not ( n31663 , n275929 );
buf ( n31664 , n31663 );
buf ( n31665 , n31664 );
buf ( n31666 , n275554 );
not ( n31667 , n275550 );
buf ( n31668 , n31667 );
buf ( n31669 , n31668 );
not ( n31670 , n275925 );
buf ( n31671 , n31670 );
buf ( n31672 , n31671 );
buf ( n31673 , n275554 );
and ( n31674 , n9158 , n9120 );
not ( n31675 , n9158 );
and ( n31676 , n31675 , n277893 );
or ( n31677 , n31674 , n31676 );
buf ( n31678 , n31677 );
buf ( n31679 , n31678 );
buf ( n31680 , RI21a12988_75);
not ( n31681 , n31680 );
not ( n31682 , n31681 );
buf ( n31683 , n31682 );
buf ( n31684 , RI210bf468_289);
not ( n31685 , n31684 );
not ( n31686 , n31685 );
buf ( n31687 , n31686 );
xor ( n31688 , n31683 , n31687 );
buf ( n31689 , RI21078ab8_504);
not ( n31690 , n31689 );
not ( n31691 , n31690 );
buf ( n31692 , n31691 );
not ( n31693 , n31692 );
xor ( n31694 , n31688 , n31693 );
xor ( n31695 , n275563 , n275568 );
and ( n31696 , n31695 , n275572 );
and ( n31697 , n275563 , n275568 );
or ( n31698 , n31696 , n31697 );
nand ( n31699 , n31694 , n31698 );
not ( n31700 , n31699 );
nor ( n31701 , n31694 , n31698 );
nor ( n31702 , n31700 , n31701 );
not ( n31703 , n31702 );
nor ( n31704 , n275590 , n275914 );
and ( n31705 , n275901 , n31704 );
and ( n31706 , n275862 , n31705 );
not ( n31707 , n275914 );
and ( n31708 , n275906 , n31707 );
nor ( n31709 , n31708 , n275916 );
or ( n31710 , n31709 , n275590 );
nand ( n31711 , n31710 , n275592 );
nor ( n31712 , n31706 , n31711 );
not ( n31713 , n31712 );
or ( n31714 , n31703 , n31713 );
or ( n31715 , n31712 , n31702 );
nand ( n31716 , n31714 , n31715 );
buf ( n31717 , n31716 );
buf ( n31718 , n31717 );
not ( n31719 , n22192 );
and ( n31720 , n31719 , n277945 );
not ( n31721 , n31719 );
not ( n31722 , n29599 );
not ( n31723 , n31420 );
or ( n31724 , n31722 , n31723 );
and ( n31725 , n31436 , n23655 );
not ( n31726 , n22052 );
not ( n31727 , n31447 );
or ( n31728 , n31726 , n31727 );
and ( n31729 , n27520 , n12294 );
and ( n31730 , n23679 , n12357 );
nor ( n31731 , n31729 , n31730 );
nand ( n31732 , n31728 , n31731 );
nor ( n31733 , n31725 , n31732 );
nand ( n31734 , n31724 , n31733 );
and ( n31735 , n31721 , n31734 );
or ( n31736 , n31720 , n31735 );
buf ( n31737 , n31736 );
buf ( n31738 , n31737 );
buf ( n31739 , n275554 );
buf ( n31740 , n275554 );
nand ( n31741 , n29226 , n29223 );
not ( n31742 , n22018 );
xor ( n31743 , n31741 , n31742 );
buf ( n31744 , n31743 );
and ( n31745 , n31744 , n28438 );
not ( n31746 , n29171 );
nor ( n31747 , n31746 , n12282 );
nor ( n31748 , n31745 , n31747 );
buf ( n31749 , n21869 );
buf ( n31750 , n21875 );
nand ( n31751 , n31749 , n31750 );
buf ( n31752 , n31751 );
buf ( n31753 , n31752 );
not ( n31754 , n31753 );
buf ( n31755 , n23529 );
buf ( n31756 , n29193 );
nand ( n31757 , n31755 , n31756 );
buf ( n31758 , n31757 );
buf ( n31759 , n31758 );
not ( n31760 , n31759 );
or ( n31761 , n31754 , n31760 );
buf ( n31762 , n31758 );
buf ( n31763 , n31752 );
or ( n31764 , n31762 , n31763 );
nand ( n31765 , n31761 , n31764 );
buf ( n31766 , n31765 );
buf ( n31767 , n31766 );
and ( n31768 , n31767 , n28408 );
not ( n31769 , n27200 );
buf ( n31770 , n22107 );
nand ( n31771 , n31769 , n31770 );
not ( n31772 , n31771 );
buf ( n31773 , n27197 );
buf ( n31774 , n29210 );
nand ( n31775 , n31773 , n31774 );
not ( n31776 , n31775 );
or ( n31777 , n31772 , n31776 );
or ( n31778 , n31775 , n31771 );
nand ( n31779 , n31777 , n31778 );
buf ( n31780 , n31779 );
and ( n31781 , n31780 , n28428 );
nor ( n31782 , n31768 , n31781 );
not ( n31783 , n28450 );
not ( n31784 , n10885 );
nand ( n31785 , n31783 , n31784 );
and ( n31786 , n28458 , n12192 );
nand ( n31787 , n20649 , n9287 );
not ( n31788 , n31787 );
nor ( n31789 , n31786 , n31788 );
nand ( n31790 , n31748 , n31782 , n31785 , n31789 );
buf ( n31791 , n31790 );
buf ( n31792 , n31791 );
buf ( n31793 , n277554 );
buf ( n31794 , n31793 );
not ( n31795 , n31794 );
buf ( n31796 , n31795 );
buf ( n31797 , n31796 );
buf ( n31798 , n277533 );
buf ( n31799 , n31798 );
not ( n31800 , n31799 );
buf ( n31801 , n31800 );
buf ( n31802 , n31801 );
nand ( n31803 , n31797 , n31802 );
buf ( n31804 , n31803 );
buf ( n31805 , n31804 );
buf ( n31806 , n31793 );
buf ( n31807 , n31798 );
nand ( n31808 , n31806 , n31807 );
buf ( n31809 , n31808 );
buf ( n31810 , n31809 );
nand ( n31811 , n31805 , n31810 );
buf ( n31812 , n31811 );
buf ( n31813 , n31812 );
not ( n31814 , n31813 );
buf ( n31815 , n277717 );
buf ( n31816 , n31815 );
buf ( n31817 , n31816 );
buf ( n31818 , n277749 );
buf ( n31819 , n31818 );
or ( n31820 , n31817 , n31819 );
buf ( n31821 , n30793 );
not ( n31822 , n31821 );
buf ( n31823 , n30795 );
not ( n31824 , n31823 );
and ( n31825 , n31822 , n31824 );
buf ( n31826 , n30840 );
nor ( n31827 , n31825 , n31826 );
buf ( n31828 , n31827 );
buf ( n31829 , n31828 );
nand ( n31830 , n31820 , n31829 );
buf ( n31831 , n31830 );
buf ( n31832 , n31831 );
not ( n31833 , n31832 );
buf ( n31834 , n31833 );
buf ( n31835 , n31834 );
buf ( n31836 , n30820 );
nand ( n31837 , n31835 , n31836 );
buf ( n31838 , n31837 );
buf ( n31839 , n31838 );
buf ( n31840 , n11789 );
buf ( n31841 , n31840 );
not ( n31842 , n31841 );
buf ( n31843 , n31842 );
buf ( n31844 , n31843 );
buf ( n31845 , n277696 );
buf ( n31846 , n31845 );
not ( n31847 , n31846 );
buf ( n31848 , n31847 );
buf ( n31849 , n31848 );
nand ( n31850 , n31844 , n31849 );
buf ( n31851 , n31850 );
buf ( n31852 , n31851 );
buf ( n31853 , n277649 );
buf ( n31854 , n31853 );
buf ( n31855 , n277628 );
buf ( n31856 , n31855 );
or ( n31857 , n31854 , n31856 );
buf ( n31858 , n31857 );
buf ( n31859 , n31858 );
nand ( n31860 , n31852 , n31859 );
buf ( n31861 , n31860 );
buf ( n31862 , n31861 );
nor ( n31863 , n31839 , n31862 );
buf ( n31864 , n31863 );
buf ( n31865 , n31864 );
not ( n31866 , n31865 );
buf ( n31867 , n27479 );
not ( n31868 , n31867 );
or ( n31869 , n31866 , n31868 );
buf ( n31870 , n31861 );
not ( n31871 , n31870 );
buf ( n31872 , n31871 );
buf ( n31873 , n31872 );
not ( n31874 , n31873 );
buf ( n31875 , n30869 );
not ( n31876 , n31875 );
buf ( n31877 , n31834 );
not ( n31878 , n31877 );
or ( n31879 , n31876 , n31878 );
buf ( n31880 , n30891 );
not ( n31881 , n31880 );
buf ( n31882 , n31816 );
not ( n31883 , n31882 );
buf ( n31884 , n31883 );
buf ( n31885 , n31884 );
buf ( n31886 , n31818 );
not ( n31887 , n31886 );
buf ( n31888 , n31887 );
buf ( n31889 , n31888 );
nand ( n31890 , n31885 , n31889 );
buf ( n31891 , n31890 );
buf ( n31892 , n31891 );
buf ( n31893 , n30798 );
and ( n31894 , n31892 , n31893 );
buf ( n31895 , n31894 );
buf ( n31896 , n31895 );
not ( n31897 , n31896 );
or ( n31898 , n31881 , n31897 );
buf ( n31899 , n30803 );
not ( n31900 , n31899 );
buf ( n31901 , n31891 );
not ( n31902 , n31901 );
or ( n31903 , n31900 , n31902 );
buf ( n31904 , n31816 );
buf ( n31905 , n31818 );
nand ( n31906 , n31904 , n31905 );
buf ( n31907 , n31906 );
buf ( n31908 , n31907 );
nand ( n31909 , n31903 , n31908 );
buf ( n31910 , n31909 );
buf ( n31911 , n31910 );
not ( n31912 , n31911 );
buf ( n31913 , n31912 );
buf ( n31914 , n31913 );
nand ( n31915 , n31898 , n31914 );
buf ( n31916 , n31915 );
buf ( n31917 , n31916 );
not ( n31918 , n31917 );
buf ( n31919 , n31918 );
buf ( n31920 , n31919 );
nand ( n31921 , n31879 , n31920 );
buf ( n31922 , n31921 );
buf ( n31923 , n31922 );
not ( n31924 , n31923 );
or ( n31925 , n31874 , n31924 );
buf ( n31926 , n31858 );
not ( n31927 , n31926 );
buf ( n31928 , n31840 );
buf ( n31929 , n31845 );
and ( n31930 , n31928 , n31929 );
buf ( n31931 , n31930 );
buf ( n31932 , n31931 );
not ( n31933 , n31932 );
or ( n31934 , n31927 , n31933 );
buf ( n31935 , n31855 );
buf ( n31936 , n31853 );
nand ( n31937 , n31935 , n31936 );
buf ( n31938 , n31937 );
buf ( n31939 , n31938 );
nand ( n31940 , n31934 , n31939 );
buf ( n31941 , n31940 );
buf ( n31942 , n31941 );
not ( n31943 , n31942 );
buf ( n31944 , n31943 );
buf ( n31945 , n31944 );
nand ( n31946 , n31925 , n31945 );
buf ( n31947 , n31946 );
buf ( n31948 , n31947 );
not ( n31949 , n31948 );
buf ( n31950 , n31949 );
buf ( n31951 , n31950 );
nand ( n31952 , n31869 , n31951 );
buf ( n31953 , n31952 );
buf ( n31954 , n31953 );
not ( n31955 , n31954 );
or ( n31956 , n31814 , n31955 );
buf ( n31957 , n31953 );
buf ( n31958 , n31812 );
or ( n31959 , n31957 , n31958 );
nand ( n31960 , n31956 , n31959 );
buf ( n31961 , n31960 );
buf ( n31962 , n31961 );
nand ( n31963 , n31962 , n31422 );
buf ( n31964 , n277554 );
not ( n31965 , n31964 );
buf ( n31966 , n277533 );
nand ( n31967 , n31965 , n31966 );
not ( n31968 , n31966 );
nand ( n31969 , n31968 , n31964 );
nand ( n31970 , n31967 , n31969 );
not ( n31971 , n31970 );
buf ( n31972 , n31815 );
not ( n31973 , n31972 );
buf ( n31974 , n277749 );
nand ( n31975 , n31973 , n31974 );
nand ( n31976 , n31975 , n30912 );
nor ( n31977 , n31976 , n30926 );
and ( n31978 , n31977 , n30931 );
not ( n31979 , n31978 );
buf ( n31980 , n277676 );
not ( n31981 , n31980 );
buf ( n31982 , n277696 );
nand ( n31983 , n31981 , n31982 );
buf ( n31984 , n277628 );
not ( n31985 , n31984 );
buf ( n31986 , n277649 );
nand ( n31987 , n31985 , n31986 );
nand ( n31988 , n31983 , n31987 );
nor ( n31989 , n31979 , n31988 );
not ( n31990 , n31989 );
not ( n31991 , n27260 );
or ( n31992 , n31990 , n31991 );
not ( n31993 , n31988 );
not ( n31994 , n31993 );
not ( n31995 , n30945 );
not ( n31996 , n31977 );
or ( n31997 , n31995 , n31996 );
not ( n31998 , n30954 );
not ( n31999 , n31976 );
not ( n32000 , n31999 );
or ( n32001 , n31998 , n32000 );
not ( n32002 , n30915 );
not ( n32003 , n31975 );
or ( n32004 , n32002 , n32003 );
not ( n32005 , n31974 );
nand ( n32006 , n32005 , n31972 );
nand ( n32007 , n32004 , n32006 );
not ( n32008 , n32007 );
nand ( n32009 , n32001 , n32008 );
not ( n32010 , n32009 );
nand ( n32011 , n31997 , n32010 );
not ( n32012 , n32011 );
or ( n32013 , n31994 , n32012 );
not ( n32014 , n31987 );
nor ( n32015 , n31981 , n31982 );
not ( n32016 , n32015 );
or ( n32017 , n32014 , n32016 );
not ( n32018 , n31986 );
nand ( n32019 , n32018 , n31984 );
nand ( n32020 , n32017 , n32019 );
not ( n32021 , n32020 );
nand ( n32022 , n32013 , n32021 );
not ( n32023 , n32022 );
nand ( n32024 , n31992 , n32023 );
not ( n32025 , n32024 );
or ( n32026 , n31971 , n32025 );
or ( n32027 , n32024 , n31970 );
nand ( n32028 , n32026 , n32027 );
buf ( n32029 , n32028 );
nand ( n32030 , n32029 , n28330 );
buf ( n32031 , n12168 );
buf ( n32032 , n32031 );
not ( n32033 , n32032 );
not ( n32034 , n32033 );
buf ( n32035 , n277676 );
nand ( n32036 , n30971 , n32035 );
nand ( n32037 , n27491 , n30965 );
nor ( n32038 , n30969 , n32036 , n32037 );
nand ( n32039 , n32038 , n30978 );
not ( n32040 , n32039 );
buf ( n32041 , n277628 );
and ( n32042 , n30481 , n30478 , n32040 , n32041 );
buf ( n32043 , n277554 );
nand ( n32044 , n32042 , n32043 );
not ( n32045 , n32044 );
buf ( n32046 , n32045 );
not ( n32047 , n32046 );
or ( n32048 , n32034 , n32047 );
or ( n32049 , n32046 , n32033 );
nand ( n32050 , n32048 , n32049 );
buf ( n32051 , n32050 );
nand ( n32052 , n32051 , n31449 );
not ( n32053 , n31451 );
not ( n32054 , n32053 );
buf ( n32055 , n277628 );
and ( n32056 , n32054 , n32055 );
not ( n32057 , n277544 );
not ( n32058 , n32057 );
not ( n32059 , n28357 );
or ( n32060 , n32058 , n32059 );
buf ( n32061 , n28233 );
or ( n32062 , n32061 , n277538 );
nand ( n32063 , n32060 , n32062 );
nor ( n32064 , n32056 , n32063 );
nand ( n32065 , n31460 , n277533 );
and ( n32066 , n32052 , n32064 , n32065 );
nand ( n32067 , n31963 , n32030 , n32066 );
buf ( n32068 , n32067 );
buf ( n32069 , n32068 );
not ( n32070 , n275550 );
buf ( n32071 , n32070 );
buf ( n32072 , n32071 );
not ( n32073 , n19635 );
buf ( n32074 , n32073 );
or ( n32075 , n21172 , n32074 );
not ( n32076 , n19649 );
and ( n32077 , n29477 , n18720 );
not ( n32078 , n29477 );
and ( n32079 , n32078 , n29478 );
nor ( n32080 , n32077 , n32079 );
not ( n32081 , n32080 );
and ( n32082 , n32076 , n32081 );
and ( n32083 , n21499 , n20353 );
nor ( n32084 , n32082 , n32083 );
and ( n32085 , n21592 , n20515 );
nor ( n32086 , n19639 , n29478 );
not ( n32087 , n32086 );
nand ( n32088 , n21618 , n20560 );
nand ( n32089 , n29494 , n21624 );
nand ( n32090 , n32087 , n32088 , n32089 );
nor ( n32091 , n32085 , n32090 );
and ( n32092 , n32084 , n32091 );
nand ( n32093 , n32075 , n32092 );
buf ( n32094 , n32093 );
buf ( n32095 , n32094 );
or ( n32096 , n23791 , n20950 );
nand ( n32097 , n20950 , n13853 );
nand ( n32098 , n32096 , n32097 );
buf ( n32099 , n32098 );
buf ( n32100 , n32099 );
buf ( n32101 , n275554 );
not ( n32102 , n275925 );
buf ( n32103 , n32102 );
buf ( n32104 , n32103 );
not ( n32105 , n275929 );
buf ( n32106 , n32105 );
buf ( n32107 , n32106 );
buf ( n32108 , n275554 );
and ( n32109 , n31719 , n277548 );
not ( n32110 , n31719 );
not ( n32111 , n29599 );
not ( n32112 , n31962 );
or ( n32113 , n32111 , n32112 );
and ( n32114 , n32029 , n30962 );
not ( n32115 , n23673 );
not ( n32116 , n32051 );
or ( n32117 , n32115 , n32116 );
and ( n32118 , n27520 , n32055 );
and ( n32119 , n22013 , n277533 );
nor ( n32120 , n32118 , n32119 );
nand ( n32121 , n32117 , n32120 );
nor ( n32122 , n32114 , n32121 );
nand ( n32123 , n32113 , n32122 );
and ( n32124 , n32110 , n32123 );
or ( n32125 , n32109 , n32124 );
buf ( n32126 , n32125 );
buf ( n32127 , n32126 );
not ( n32128 , n275929 );
buf ( n32129 , n32128 );
buf ( n32130 , n32129 );
buf ( n32131 , n14513 );
and ( n32132 , n20711 , n32131 );
not ( n32133 , n20711 );
buf ( n32134 , n14515 );
not ( n32135 , n32134 );
not ( n32136 , n32135 );
buf ( n32137 , n14600 );
not ( n32138 , n32137 );
buf ( n32139 , n14581 );
not ( n32140 , n32139 );
buf ( n32141 , n14615 );
nand ( n32142 , n14567 , n32141 );
nor ( n32143 , n32140 , n32142 );
nand ( n32144 , n14778 , n32143 );
nor ( n32145 , n32138 , n32144 );
not ( n32146 , n32145 );
or ( n32147 , n32136 , n32146 );
nand ( n32148 , n32147 , n20830 );
nor ( n32149 , n32134 , n20830 );
nand ( n32150 , n32145 , n32149 );
nand ( n32151 , n32148 , n32150 );
buf ( n32152 , n32151 );
and ( n32153 , n32133 , n32152 );
nor ( n32154 , n32132 , n32153 );
or ( n32155 , n32154 , n26364 );
not ( n32156 , n16895 );
not ( n32157 , n16392 );
nand ( n32158 , n32156 , n32157 );
not ( n32159 , n32158 );
not ( n32160 , n20875 );
or ( n32161 , n32159 , n32160 );
or ( n32162 , n32158 , n20875 );
nand ( n32163 , n32161 , n32162 );
buf ( n32164 , n32163 );
nand ( n32165 , n32164 , n26370 );
not ( n32166 , n17227 );
and ( n32167 , n32166 , n17335 );
not ( n32168 , n32167 );
not ( n32169 , n20913 );
not ( n32170 , n32169 );
or ( n32171 , n32168 , n32170 );
or ( n32172 , n32169 , n32167 );
nand ( n32173 , n32171 , n32172 );
buf ( n32174 , n32173 );
nand ( n32175 , n32174 , n26374 );
not ( n32176 , n26390 );
and ( n32177 , n17508 , n17509 );
not ( n32178 , n17508 );
and ( n32179 , n32178 , n13632 );
nor ( n32180 , n32177 , n32179 );
nand ( n32181 , n32176 , n32180 );
not ( n32182 , n17439 );
not ( n32183 , n26486 );
or ( n32184 , n32182 , n32183 );
or ( n32185 , n26486 , n17439 );
nand ( n32186 , n32184 , n32185 );
buf ( n32187 , n32186 );
not ( n32188 , n26392 );
nand ( n32189 , n32187 , n32188 );
buf ( n32190 , n17438 );
buf ( n32191 , n32190 );
buf ( n32192 , n32191 );
nand ( n32193 , n26395 , n32192 );
not ( n32194 , n30514 );
and ( n32195 , n32189 , n32193 , n32194 );
and ( n32196 , n32165 , n32175 , n32181 , n32195 );
nand ( n32197 , n32155 , n32196 );
buf ( n32198 , n32197 );
buf ( n32199 , n32198 );
not ( n32200 , n25019 );
or ( n32201 , n32200 , n23807 );
nand ( n32202 , n13434 , n14830 );
nand ( n32203 , n32201 , n32202 );
buf ( n32204 , n32203 );
buf ( n32205 , n32204 );
nand ( n32206 , n275717 , n275766 );
not ( n32207 , n32206 );
not ( n32208 , n275763 );
or ( n32209 , n32207 , n32208 );
or ( n32210 , n275763 , n32206 );
nand ( n32211 , n32209 , n32210 );
buf ( n32212 , n32211 );
buf ( n32213 , n32212 );
not ( n32214 , n22057 );
not ( n32215 , n31780 );
or ( n32216 , n32214 , n32215 );
nand ( n32217 , n31744 , n22052 );
nand ( n32218 , n32216 , n32217 );
not ( n32219 , n22002 );
not ( n32220 , n31767 );
or ( n32221 , n32219 , n32220 );
not ( n32222 , n22006 );
not ( n32223 , n12282 );
and ( n32224 , n32222 , n32223 );
and ( n32225 , n23679 , n12192 );
nor ( n32226 , n32224 , n32225 );
nand ( n32227 , n32221 , n32226 );
nor ( n32228 , n32218 , n32227 );
or ( n32229 , n32228 , n23705 );
nand ( n32230 , n23705 , n11090 );
nand ( n32231 , n32229 , n32230 );
buf ( n32232 , n32231 );
buf ( n32233 , n32232 );
or ( n32234 , n24400 , n19216 );
nand ( n32235 , n24415 , n19360 );
nand ( n32236 , n24429 , n19354 );
not ( n32237 , n18391 );
not ( n32238 , n19653 );
not ( n32239 , n32238 );
or ( n32240 , n32237 , n32239 );
or ( n32241 , n32238 , n18391 );
nand ( n32242 , n32240 , n32241 );
not ( n32243 , n32242 );
not ( n32244 , n19318 );
or ( n32245 , n32243 , n32244 );
or ( n32246 , n19291 , n24438 );
nand ( n32247 , n32245 , n32246 );
nand ( n32248 , n19177 , n19219 );
nor ( n32249 , n32248 , n24443 );
not ( n32250 , n18383 );
nor ( n32251 , n32250 , n19388 );
nor ( n32252 , n32247 , n32249 , n32251 );
and ( n32253 , n32235 , n32236 , n32252 );
nand ( n32254 , n32234 , n32253 );
buf ( n32255 , n32254 );
buf ( n32256 , n32255 );
buf ( n32257 , n275554 );
buf ( n32258 , n275554 );
and ( n32259 , n22335 , n18131 );
not ( n32260 , n22335 );
and ( n32261 , n32260 , n19280 );
or ( n32262 , n32259 , n32261 );
buf ( n32263 , n32262 );
buf ( n32264 , n32263 );
not ( n32265 , n20672 );
xor ( n32266 , n31293 , n31294 );
buf ( n32267 , n32266 );
not ( n32268 , n32267 );
or ( n32269 , n32265 , n32268 );
nand ( n32270 , n29042 , n31304 );
nand ( n32271 , n32269 , n32270 );
not ( n32272 , n32271 );
or ( n32273 , n32272 , n26365 );
not ( n32274 , n16937 );
nand ( n32275 , n32274 , n15791 );
not ( n32276 , n32275 );
nor ( n32277 , n23722 , n23717 );
not ( n32278 , n32277 );
not ( n32279 , n16913 );
or ( n32280 , n32278 , n32279 );
not ( n32281 , n23720 );
not ( n32282 , n23717 );
and ( n32283 , n32281 , n32282 );
nor ( n32284 , n32283 , n16935 );
nand ( n32285 , n32280 , n32284 );
not ( n32286 , n32285 );
or ( n32287 , n32276 , n32286 );
or ( n32288 , n32285 , n32275 );
nand ( n32289 , n32287 , n32288 );
buf ( n32290 , n32289 );
nand ( n32291 , n32290 , n26370 );
or ( n32292 , n17386 , n17032 );
not ( n32293 , n32292 );
not ( n32294 , n17008 );
nor ( n32295 , n32294 , n23732 );
not ( n32296 , n32295 );
not ( n32297 , n17362 );
or ( n32298 , n32296 , n32297 );
not ( n32299 , n23753 );
not ( n32300 , n23732 );
and ( n32301 , n32299 , n32300 );
not ( n32302 , n23734 );
nor ( n32303 , n32301 , n32302 );
nand ( n32304 , n32298 , n32303 );
not ( n32305 , n32304 );
or ( n32306 , n32293 , n32305 );
or ( n32307 , n32304 , n32292 );
nand ( n32308 , n32306 , n32307 );
buf ( n32309 , n32308 );
nand ( n32310 , n32309 , n26374 );
and ( n32311 , n17525 , n13897 );
not ( n32312 , n17525 );
and ( n32313 , n32312 , n17526 );
nor ( n32314 , n32311 , n32313 );
nor ( n32315 , n26390 , n32314 );
nor ( n32316 , n14830 , n17526 );
not ( n32317 , n32316 );
not ( n32318 , n17478 );
not ( n32319 , n24610 );
or ( n32320 , n32318 , n32319 );
or ( n32321 , n24610 , n17478 );
nand ( n32322 , n32320 , n32321 );
buf ( n32323 , n32322 );
nand ( n32324 , n32323 , n26393 );
buf ( n32325 , n17477 );
buf ( n32326 , n32325 );
buf ( n32327 , n32326 );
nand ( n32328 , n26395 , n32327 );
nand ( n32329 , n32317 , n32324 , n32328 );
nor ( n32330 , n32315 , n32329 );
and ( n32331 , n32291 , n32310 , n32330 );
nand ( n32332 , n32273 , n32331 );
buf ( n32333 , n32332 );
buf ( n32334 , n32333 );
or ( n32335 , n32154 , n14908 );
nand ( n32336 , n32164 , n16968 );
nand ( n32337 , n32174 , n17405 );
not ( n32338 , n32187 );
not ( n32339 , n17410 );
not ( n32340 , n32339 );
or ( n32341 , n32338 , n32340 );
nand ( n32342 , n17545 , n32180 );
nand ( n32343 , n32341 , n32342 );
not ( n32344 , n32192 );
nor ( n32345 , n32344 , n17500 );
not ( n32346 , n13625 );
nor ( n32347 , n17561 , n32346 );
nor ( n32348 , n32343 , n32345 , n32347 );
and ( n32349 , n32336 , n32337 , n32348 );
nand ( n32350 , n32335 , n32349 );
buf ( n32351 , n32350 );
buf ( n32352 , n32351 );
buf ( n32353 , n14486 );
not ( n32354 , n32353 );
not ( n32355 , n32354 );
and ( n32356 , n20712 , n32355 );
not ( n32357 , n20712 );
not ( n32358 , n20834 );
buf ( n32359 , n20833 );
not ( n32360 , n32359 );
or ( n32361 , n32358 , n32360 );
or ( n32362 , n32359 , n20834 );
nand ( n32363 , n32361 , n32362 );
buf ( n32364 , n32363 );
and ( n32365 , n32357 , n32364 );
nor ( n32366 , n32356 , n32365 );
not ( n32367 , n32366 );
and ( n32368 , n32367 , n23404 );
or ( n32369 , n16899 , n16400 );
not ( n32370 , n32369 );
not ( n32371 , n32157 );
not ( n32372 , n20875 );
or ( n32373 , n32371 , n32372 );
not ( n32374 , n16895 );
nand ( n32375 , n32373 , n32374 );
not ( n32376 , n32375 );
or ( n32377 , n32370 , n32376 );
or ( n32378 , n32375 , n32369 );
nand ( n32379 , n32377 , n32378 );
buf ( n32380 , n32379 );
nand ( n32381 , n32380 , n20889 );
not ( n32382 , n17217 );
nand ( n32383 , n32382 , n20917 );
not ( n32384 , n32383 );
not ( n32385 , n32166 );
not ( n32386 , n20913 );
or ( n32387 , n32385 , n32386 );
nand ( n32388 , n32387 , n17335 );
not ( n32389 , n32388 );
or ( n32390 , n32384 , n32389 );
or ( n32391 , n32388 , n32383 );
nand ( n32392 , n32390 , n32391 );
buf ( n32393 , n32392 );
nand ( n32394 , n32393 , n24711 );
not ( n32395 , n17437 );
nor ( n32396 , n20930 , n17439 );
not ( n32397 , n32396 );
or ( n32398 , n32395 , n32397 );
or ( n32399 , n32396 , n17437 );
nand ( n32400 , n32398 , n32399 );
buf ( n32401 , n32400 );
and ( n32402 , n32401 , n17409 );
buf ( n32403 , n17436 );
buf ( n32404 , n32403 );
buf ( n32405 , n32404 );
and ( n32406 , n17499 , n32405 );
nor ( n32407 , n32402 , n32406 );
nand ( n32408 , n32381 , n32394 , n32407 );
nor ( n32409 , n32368 , n32408 );
or ( n32410 , n32409 , n27647 );
nand ( n32411 , n21696 , n13614 );
nand ( n32412 , n32410 , n32411 );
buf ( n32413 , n32412 );
buf ( n32414 , n32413 );
buf ( n32415 , n275554 );
nand ( n32416 , n25064 , n26083 );
buf ( n32417 , n25255 );
not ( n32418 , n32417 );
buf ( n32419 , n25139 );
nor ( n32420 , n32418 , n32419 );
buf ( n32421 , n32420 );
buf ( n32422 , n32421 );
not ( n32423 , n32422 );
buf ( n32424 , n25173 );
buf ( n32425 , n25221 );
buf ( n32426 , n25148 );
not ( n32427 , n32426 );
buf ( n32428 , n32427 );
buf ( n32429 , n32428 );
and ( n32430 , n32424 , n32425 , n32429 );
buf ( n32431 , n32428 );
not ( n32432 , n32431 );
buf ( n32433 , n25242 );
not ( n32434 , n32433 );
or ( n32435 , n32432 , n32434 );
buf ( n32436 , n25249 );
nand ( n32437 , n32435 , n32436 );
buf ( n32438 , n32437 );
buf ( n32439 , n32438 );
nor ( n32440 , n32430 , n32439 );
buf ( n32441 , n32440 );
buf ( n32442 , n32441 );
not ( n32443 , n32442 );
or ( n32444 , n32423 , n32443 );
buf ( n32445 , n32441 );
buf ( n32446 , n32421 );
or ( n32447 , n32445 , n32446 );
nand ( n32448 , n32444 , n32447 );
buf ( n32449 , n32448 );
buf ( n32450 , n32449 );
not ( n32451 , n32450 );
nor ( n32452 , n32451 , n25389 );
nand ( n32453 , n25397 , n275633 );
buf ( n32454 , n25577 );
not ( n32455 , n32454 );
buf ( n32456 , n25472 );
nor ( n32457 , n32455 , n32456 );
buf ( n32458 , n32457 );
buf ( n32459 , n32458 );
not ( n32460 , n32459 );
buf ( n32461 , n25494 );
buf ( n32462 , n25540 );
buf ( n32463 , n25465 );
not ( n32464 , n32463 );
buf ( n32465 , n32464 );
buf ( n32466 , n32465 );
and ( n32467 , n32461 , n32462 , n32466 );
buf ( n32468 , n32465 );
not ( n32469 , n32468 );
buf ( n32470 , n25560 );
buf ( n32471 , n25554 );
and ( n32472 , n32470 , n32471 );
buf ( n32473 , n25484 );
nor ( n32474 , n32472 , n32473 );
buf ( n32475 , n32474 );
buf ( n32476 , n32475 );
not ( n32477 , n32476 );
or ( n32478 , n32469 , n32477 );
buf ( n32479 , n25571 );
nand ( n32480 , n32478 , n32479 );
buf ( n32481 , n32480 );
buf ( n32482 , n32481 );
nor ( n32483 , n32467 , n32482 );
buf ( n32484 , n32483 );
buf ( n32485 , n32484 );
not ( n32486 , n32485 );
or ( n32487 , n32460 , n32486 );
buf ( n32488 , n32484 );
buf ( n32489 , n32458 );
or ( n32490 , n32488 , n32489 );
nand ( n32491 , n32487 , n32490 );
buf ( n32492 , n32491 );
buf ( n32493 , n32492 );
and ( n32494 , n25402 , n32493 );
not ( n32495 , n18887 );
nor ( n32496 , n32495 , n19639 );
nor ( n32497 , n32494 , n32496 );
buf ( n32498 , n25893 );
not ( n32499 , n32498 );
buf ( n32500 , n25789 );
nor ( n32501 , n32499 , n32500 );
buf ( n32502 , n32501 );
buf ( n32503 , n32502 );
not ( n32504 , n32503 );
buf ( n32505 , n25810 );
buf ( n32506 , n25856 );
buf ( n32507 , n25780 );
not ( n32508 , n32507 );
buf ( n32509 , n32508 );
buf ( n32510 , n32509 );
and ( n32511 , n32505 , n32506 , n32510 );
buf ( n32512 , n32509 );
not ( n32513 , n32512 );
buf ( n32514 , n25876 );
buf ( n32515 , n25870 );
and ( n32516 , n32514 , n32515 );
buf ( n32517 , n25800 );
nor ( n32518 , n32516 , n32517 );
buf ( n32519 , n32518 );
buf ( n32520 , n32519 );
not ( n32521 , n32520 );
or ( n32522 , n32513 , n32521 );
buf ( n32523 , n25887 );
nand ( n32524 , n32522 , n32523 );
buf ( n32525 , n32524 );
buf ( n32526 , n32525 );
nor ( n32527 , n32511 , n32526 );
buf ( n32528 , n32527 );
buf ( n32529 , n32528 );
not ( n32530 , n32529 );
or ( n32531 , n32504 , n32530 );
buf ( n32532 , n32528 );
buf ( n32533 , n32502 );
or ( n32534 , n32532 , n32533 );
nand ( n32535 , n32531 , n32534 );
buf ( n32536 , n32535 );
buf ( n32537 , n32536 );
nand ( n32538 , n25717 , n32537 );
nand ( n32539 , n32453 , n32497 , n32538 );
nor ( n32540 , n32452 , n32539 );
buf ( n32541 , n26203 );
not ( n32542 , n32541 );
buf ( n32543 , n26089 );
nor ( n32544 , n32542 , n32543 );
buf ( n32545 , n32544 );
buf ( n32546 , n32545 );
not ( n32547 , n32546 );
buf ( n32548 , n26119 );
buf ( n32549 , n26166 );
buf ( n32550 , n26097 );
not ( n32551 , n32550 );
buf ( n32552 , n32551 );
buf ( n32553 , n32552 );
and ( n32554 , n32548 , n32549 , n32553 );
buf ( n32555 , n32552 );
not ( n32556 , n32555 );
buf ( n32557 , n26189 );
not ( n32558 , n32557 );
or ( n32559 , n32556 , n32558 );
buf ( n32560 , n26197 );
nand ( n32561 , n32559 , n32560 );
buf ( n32562 , n32561 );
buf ( n32563 , n32562 );
nor ( n32564 , n32554 , n32563 );
buf ( n32565 , n32564 );
buf ( n32566 , n32565 );
not ( n32567 , n32566 );
or ( n32568 , n32547 , n32567 );
buf ( n32569 , n32565 );
buf ( n32570 , n32545 );
or ( n32571 , n32569 , n32570 );
nand ( n32572 , n32568 , n32571 );
buf ( n32573 , n32572 );
buf ( n32574 , n32573 );
nand ( n32575 , n26027 , n32574 );
nand ( n32576 , n32416 , n32540 , n32575 );
buf ( n32577 , n32576 );
buf ( n32578 , n32577 );
not ( n32579 , n14855 );
or ( n32580 , n14840 , n32579 );
nand ( n32581 , n32580 , n14859 );
buf ( n32582 , n32581 );
buf ( n32583 , n32582 );
not ( n32584 , n275550 );
buf ( n32585 , n32584 );
buf ( n32586 , n32585 );
not ( n32587 , n275550 );
buf ( n32588 , n32587 );
buf ( n32589 , n32588 );
not ( n32590 , n275550 );
buf ( n32591 , n32590 );
buf ( n32592 , n32591 );
not ( n32593 , n275550 );
buf ( n32594 , n32593 );
buf ( n32595 , n32594 );
not ( n32596 , n275550 );
buf ( n32597 , n32596 );
buf ( n32598 , n32597 );
buf ( n32599 , n275554 );
nand ( n32600 , n29346 , n28306 );
nand ( n32601 , n29359 , n28330 );
and ( n32602 , n28332 , n29369 );
and ( n32603 , n28350 , n12130 );
nor ( n32604 , n32602 , n32603 );
not ( n32605 , n12270 );
and ( n32606 , n28231 , n32605 );
or ( n32607 , n28354 , n11625 );
not ( n32608 , n11644 );
nand ( n32609 , n28357 , n32608 );
nand ( n32610 , n32607 , n32609 );
nor ( n32611 , n32606 , n32610 );
nand ( n32612 , n32600 , n32601 , n32604 , n32611 );
buf ( n32613 , n32612 );
buf ( n32614 , n32613 );
buf ( n32615 , n275554 );
buf ( n32616 , n275554 );
buf ( n32617 , n14383 );
and ( n32618 , n20712 , n32617 );
not ( n32619 , n20712 );
buf ( n32620 , n14779 );
and ( n32621 , n32620 , n14781 );
not ( n32622 , n32620 );
and ( n32623 , n32622 , n14780 );
nor ( n32624 , n32621 , n32623 );
buf ( n32625 , n32624 );
and ( n32626 , n32619 , n32625 );
nor ( n32627 , n32618 , n32626 );
not ( n32628 , n32627 );
not ( n32629 , n23789 );
and ( n32630 , n32628 , n32629 );
not ( n32631 , n20889 );
not ( n32632 , n16019 );
nand ( n32633 , n32632 , n16928 );
not ( n32634 , n32633 );
nand ( n32635 , n16137 , n16076 );
nor ( n32636 , n20796 , n32635 );
not ( n32637 , n32636 );
not ( n32638 , n16913 );
or ( n32639 , n32637 , n32638 );
not ( n32640 , n20804 );
not ( n32641 , n32635 );
and ( n32642 , n32640 , n32641 );
not ( n32643 , n16076 );
not ( n32644 , n16933 );
or ( n32645 , n32643 , n32644 );
nand ( n32646 , n32645 , n16926 );
nor ( n32647 , n32642 , n32646 );
nand ( n32648 , n32639 , n32647 );
not ( n32649 , n32648 );
or ( n32650 , n32634 , n32649 );
or ( n32651 , n32648 , n32633 );
nand ( n32652 , n32650 , n32651 );
buf ( n32653 , n32652 );
not ( n32654 , n32653 );
or ( n32655 , n32631 , n32654 );
not ( n32656 , n17049 );
nand ( n32657 , n32656 , n17367 );
not ( n32658 , n32657 );
not ( n32659 , n17088 );
not ( n32660 , n17060 );
nand ( n32661 , n32659 , n32660 );
nor ( n32662 , n20747 , n32661 );
not ( n32663 , n32662 );
not ( n32664 , n17362 );
or ( n32665 , n32663 , n32664 );
not ( n32666 , n20753 );
not ( n32667 , n32661 );
and ( n32668 , n32666 , n32667 );
not ( n32669 , n32660 );
not ( n32670 , n17372 );
or ( n32671 , n32669 , n32670 );
nand ( n32672 , n32671 , n17365 );
nor ( n32673 , n32668 , n32672 );
nand ( n32674 , n32665 , n32673 );
not ( n32675 , n32674 );
or ( n32676 , n32658 , n32675 );
or ( n32677 , n32674 , n32657 );
nand ( n32678 , n32676 , n32677 );
buf ( n32679 , n32678 );
and ( n32680 , n32679 , n20926 );
not ( n32681 , n17409 );
not ( n32682 , n17484 );
nor ( n32683 , n23871 , n17475 );
and ( n32684 , n17462 , n20775 , n32683 );
not ( n32685 , n32684 );
or ( n32686 , n32682 , n32685 );
or ( n32687 , n32684 , n17484 );
nand ( n32688 , n32686 , n32687 );
buf ( n32689 , n32688 );
not ( n32690 , n32689 );
or ( n32691 , n32681 , n32690 );
buf ( n32692 , n17483 );
buf ( n32693 , n32692 );
buf ( n32694 , n32693 );
nand ( n32695 , n17499 , n32694 );
nand ( n32696 , n32691 , n32695 );
nor ( n32697 , n32680 , n32696 );
nand ( n32698 , n32655 , n32697 );
nor ( n32699 , n32630 , n32698 );
or ( n32700 , n32699 , n21697 );
nand ( n32701 , n21696 , n13800 );
nand ( n32702 , n32700 , n32701 );
buf ( n32703 , n32702 );
buf ( n32704 , n32703 );
buf ( n32705 , n275554 );
buf ( n32706 , n275554 );
buf ( n32707 , n275554 );
not ( n32708 , n26727 );
or ( n32709 , n32708 , n22335 );
or ( n32710 , n275557 , n19188 );
nand ( n32711 , n32709 , n32710 );
buf ( n32712 , n32711 );
buf ( n32713 , n32712 );
not ( n32714 , n275925 );
buf ( n32715 , n32714 );
buf ( n32716 , n32715 );
buf ( n32717 , n275554 );
buf ( n32718 , n275554 );
nand ( n32719 , n28398 , n23603 );
nand ( n32720 , n28426 , n27266 );
and ( n32721 , n28433 , n29371 );
not ( n32722 , n22007 );
not ( n32723 , n28456 );
or ( n32724 , n32722 , n32723 );
or ( n32725 , n22014 , n12221 );
nand ( n32726 , n32724 , n32725 );
nor ( n32727 , n32721 , n32726 );
and ( n32728 , n32719 , n32720 , n32727 );
or ( n32729 , n32728 , n27179 );
nand ( n32730 , n23708 , n11372 );
nand ( n32731 , n32729 , n32730 );
buf ( n32732 , n32731 );
buf ( n32733 , n32732 );
not ( n32734 , n275856 );
nor ( n32735 , n32734 , n275665 );
not ( n32736 , n32735 );
and ( n32737 , n275847 , n275645 );
nor ( n32738 , n32737 , n275853 );
not ( n32739 , n32738 );
or ( n32740 , n32736 , n32739 );
or ( n32741 , n32738 , n32735 );
nand ( n32742 , n32740 , n32741 );
buf ( n32743 , n32742 );
buf ( n32744 , n32743 );
buf ( n32745 , n275554 );
not ( n32746 , n275550 );
buf ( n32747 , n32746 );
buf ( n32748 , n32747 );
buf ( n32749 , n275554 );
nand ( n32750 , n28303 , n28408 );
not ( n32751 , n28429 );
nand ( n32752 , n28326 , n32751 );
nand ( n32753 , n28348 , n28440 );
nand ( n32754 , n28451 , n11404 );
not ( n32755 , n29172 );
and ( n32756 , n32755 , n12219 );
not ( n32757 , n28458 );
or ( n32758 , n32757 , n12360 );
nand ( n32759 , n20649 , n9317 );
nand ( n32760 , n32758 , n32759 );
nor ( n32761 , n32756 , n32760 );
and ( n32762 , n32753 , n32754 , n32761 );
nand ( n32763 , n32750 , n32752 , n32762 );
buf ( n32764 , n32763 );
buf ( n32765 , n32764 );
not ( n32766 , n275929 );
buf ( n32767 , n32766 );
buf ( n32768 , n32767 );
not ( n32769 , n19072 );
not ( n32770 , n24450 );
or ( n32771 , n32769 , n32770 );
not ( n32772 , n19102 );
and ( n32773 , n32772 , n20987 );
not ( n32774 , n19358 );
not ( n32775 , n19372 );
or ( n32776 , n32774 , n32775 );
and ( n32777 , n19347 , n21001 );
not ( n32778 , n19286 );
not ( n32779 , n19219 );
or ( n32780 , n32778 , n32779 );
or ( n32781 , n19312 , n19289 );
nand ( n32782 , n32780 , n32781 );
nor ( n32783 , n32777 , n32782 );
nand ( n32784 , n32776 , n32783 );
nor ( n32785 , n32773 , n32784 );
or ( n32786 , n32785 , n24450 );
nand ( n32787 , n32771 , n32786 );
buf ( n32788 , n32787 );
buf ( n32789 , n32788 );
buf ( n32790 , n12226 );
buf ( n32791 , n277386 );
nand ( n32792 , n32790 , n32791 );
not ( n32793 , n32031 );
nor ( n32794 , n32792 , n32793 );
buf ( n32795 , n11748 );
not ( n32796 , n32795 );
not ( n32797 , n32043 );
nor ( n32798 , n32796 , n32797 );
nand ( n32799 , n32794 , n32798 );
not ( n32800 , n32799 );
not ( n32801 , n32039 );
and ( n32802 , n32801 , n30478 , n30481 , n32041 );
nand ( n32803 , n32800 , n32802 );
buf ( n32804 , n12322 );
buf ( n32805 , n32804 );
not ( n32806 , n32805 );
and ( n32807 , n32803 , n32806 );
not ( n32808 , n32803 );
and ( n32809 , n32808 , n32805 );
nor ( n32810 , n32807 , n32809 );
buf ( n32811 , n32810 );
buf ( n32812 , n11728 );
not ( n32813 , n32812 );
nor ( n32814 , n32811 , n32813 );
not ( n32815 , n21999 );
or ( n32816 , n32814 , n32815 );
nand ( n32817 , n32816 , n12118 );
and ( n32818 , n20627 , n32813 );
not ( n32819 , n32813 );
and ( n32820 , n20581 , n32819 );
nor ( n32821 , n32818 , n32820 );
not ( n32822 , n32821 );
not ( n32823 , n20588 );
and ( n32824 , n32822 , n32823 );
or ( n32825 , n12688 , n12118 );
nand ( n32826 , n32825 , n12679 );
nor ( n32827 , n32824 , n32826 );
nand ( n32828 , n32817 , n32827 );
not ( n32829 , n277497 );
not ( n32830 , n32813 );
or ( n32831 , n32829 , n32830 );
nand ( n32832 , n32819 , n9172 );
nand ( n32833 , n32831 , n32832 );
nand ( n32834 , n23704 , n32833 );
or ( n32835 , n32828 , n32834 );
buf ( n32836 , n9377 );
nand ( n32837 , n27641 , n32836 );
nand ( n32838 , n32835 , n32837 );
buf ( n32839 , n32838 );
buf ( n32840 , n32839 );
not ( n32841 , n29506 );
or ( n32842 , n32841 , n21770 );
nand ( n32843 , n21774 , n9579 );
nand ( n32844 , n32842 , n32843 );
buf ( n32845 , n32844 );
buf ( n32846 , n32845 );
not ( n32847 , n275925 );
buf ( n32848 , n32847 );
buf ( n32849 , n32848 );
not ( n32850 , n275925 );
buf ( n32851 , n32850 );
buf ( n32852 , n32851 );
buf ( n32853 , n275554 );
buf ( n32854 , n275554 );
buf ( n32855 , n275554 );
buf ( n32856 , n275554 );
buf ( n32857 , n275554 );
not ( n32858 , n275929 );
buf ( n32859 , n32858 );
buf ( n32860 , n32859 );
buf ( n32861 , n275554 );
not ( n32862 , n275929 );
buf ( n32863 , n32862 );
buf ( n32864 , n32863 );
buf ( n32865 , n275554 );
buf ( n32866 , n275554 );
not ( n32867 , n275929 );
buf ( n32868 , n32867 );
buf ( n32869 , n32868 );
buf ( n32870 , n275554 );
buf ( n32871 , n275554 );
not ( n32872 , n22335 );
not ( n32873 , n28549 );
not ( n32874 , n32873 );
or ( n32875 , n32872 , n32874 );
not ( n32876 , n26833 );
or ( n32877 , n32876 , n22335 );
nand ( n32878 , n32875 , n32877 );
buf ( n32879 , n32878 );
buf ( n32880 , n32879 );
not ( n32881 , n275929 );
buf ( n32882 , n32881 );
buf ( n32883 , n32882 );
or ( n32884 , n27696 , n26364 );
nand ( n32885 , n27711 , n26370 );
nand ( n32886 , n27724 , n26374 );
and ( n32887 , n17514 , n17515 );
not ( n32888 , n17514 );
and ( n32889 , n32888 , n13715 );
nor ( n32890 , n32887 , n32889 );
nand ( n32891 , n31180 , n32890 );
nand ( n32892 , n27737 , n26393 );
nand ( n32893 , n26395 , n27728 );
not ( n32894 , n22906 );
and ( n32895 , n32892 , n32893 , n32894 );
and ( n32896 , n32885 , n32886 , n32891 , n32895 );
nand ( n32897 , n32884 , n32896 );
buf ( n32898 , n32897 );
buf ( n32899 , n32898 );
not ( n32900 , n20740 );
not ( n32901 , n20846 );
and ( n32902 , n32900 , n32901 );
not ( n32903 , n20889 );
not ( n32904 , n20813 );
or ( n32905 , n32903 , n32904 );
and ( n32906 , n20762 , n24711 );
not ( n32907 , n17409 );
not ( n32908 , n20782 );
or ( n32909 , n32907 , n32908 );
nand ( n32910 , n17499 , n20788 );
nand ( n32911 , n32909 , n32910 );
nor ( n32912 , n32906 , n32911 );
nand ( n32913 , n32905 , n32912 );
nor ( n32914 , n32902 , n32913 );
or ( n32915 , n32914 , n23887 );
nand ( n32916 , n20950 , n13832 );
nand ( n32917 , n32915 , n32916 );
buf ( n32918 , n32917 );
buf ( n32919 , n32918 );
buf ( n32920 , n275554 );
not ( n32921 , n275929 );
buf ( n32922 , n32921 );
buf ( n32923 , n32922 );
buf ( n32924 , n275554 );
not ( n32925 , n275925 );
buf ( n32926 , n32925 );
buf ( n32927 , n32926 );
not ( n32928 , n23386 );
not ( n32929 , n32139 );
not ( n32930 , n32142 );
nand ( n32931 , n32930 , n20664 );
not ( n32932 , n32931 );
or ( n32933 , n32929 , n32932 );
or ( n32934 , n32931 , n32139 );
nand ( n32935 , n32933 , n32934 );
buf ( n32936 , n32935 );
not ( n32937 , n32936 );
or ( n32938 , n32928 , n32937 );
nand ( n32939 , n28249 , n13373 );
nand ( n32940 , n32938 , n32939 );
not ( n32941 , n32940 );
or ( n32942 , n32941 , n26364 );
buf ( n32943 , n20865 );
buf ( n32944 , n16861 );
not ( n32945 , n16867 );
nand ( n32946 , n32944 , n32945 );
xnor ( n32947 , n32943 , n32946 );
buf ( n32948 , n32947 );
nand ( n32949 , n32948 , n26370 );
buf ( n32950 , n20904 );
buf ( n32951 , n17281 );
buf ( n32952 , n17317 );
nand ( n32953 , n32951 , n32952 );
xnor ( n32954 , n32950 , n32953 );
buf ( n32955 , n32954 );
nand ( n32956 , n32955 , n26374 );
buf ( n32957 , n16845 );
buf ( n32958 , n32957 );
nand ( n32959 , n26395 , n32958 );
buf ( n32960 , n17412 );
and ( n32961 , n32960 , n24714 );
not ( n32962 , n32960 );
and ( n32963 , n32962 , n17433 );
nor ( n32964 , n32961 , n32963 );
buf ( n32965 , n32964 );
and ( n32966 , n26393 , n32965 );
not ( n32967 , n13652 );
nor ( n32968 , n14830 , n32967 );
nor ( n32969 , n32966 , n32968 );
nand ( n32970 , n32949 , n32956 , n32959 , n32969 );
and ( n32971 , n32967 , n13555 );
not ( n32972 , n13554 );
and ( n32973 , n13653 , n32972 );
nor ( n32974 , n32971 , n32973 );
nor ( n32975 , n26390 , n32974 );
nor ( n32976 , n32970 , n32975 );
nand ( n32977 , n32942 , n32976 );
buf ( n32978 , n32977 );
buf ( n32979 , n32978 );
buf ( n32980 , n14359 );
and ( n32981 , n20712 , n32980 );
not ( n32982 , n20712 );
nand ( n32983 , n20731 , n20732 );
buf ( n32984 , n14337 );
not ( n32985 , n32984 );
and ( n32986 , n32983 , n32985 );
not ( n32987 , n32983 );
and ( n32988 , n32987 , n32984 );
nor ( n32989 , n32986 , n32988 );
buf ( n32990 , n32989 );
and ( n32991 , n32982 , n32990 );
nor ( n32992 , n32981 , n32991 );
or ( n32993 , n32992 , n26365 );
nand ( n32994 , n16076 , n16926 );
not ( n32995 , n32994 );
nor ( n32996 , n20796 , n16136 );
not ( n32997 , n32996 );
not ( n32998 , n16913 );
or ( n32999 , n32997 , n32998 );
not ( n33000 , n20804 );
not ( n33001 , n16136 );
and ( n33002 , n33000 , n33001 );
nor ( n33003 , n33002 , n16933 );
nand ( n33004 , n32999 , n33003 );
not ( n33005 , n33004 );
or ( n33006 , n32995 , n33005 );
or ( n33007 , n32994 , n33004 );
nand ( n33008 , n33006 , n33007 );
buf ( n33009 , n33008 );
nand ( n33010 , n33009 , n26370 );
nand ( n33011 , n32660 , n17365 );
not ( n33012 , n33011 );
nor ( n33013 , n20747 , n17088 );
not ( n33014 , n33013 );
not ( n33015 , n17362 );
or ( n33016 , n33014 , n33015 );
not ( n33017 , n20753 );
not ( n33018 , n17088 );
and ( n33019 , n33017 , n33018 );
nor ( n33020 , n33019 , n17372 );
nand ( n33021 , n33016 , n33020 );
not ( n33022 , n33021 );
or ( n33023 , n33012 , n33022 );
or ( n33024 , n33021 , n33011 );
nand ( n33025 , n33023 , n33024 );
buf ( n33026 , n33025 );
nand ( n33027 , n33026 , n26374 );
not ( n33028 , n13879 );
and ( n33029 , n17530 , n33028 );
not ( n33030 , n17530 );
and ( n33031 , n33030 , n13880 );
nor ( n33032 , n33029 , n33031 );
nor ( n33033 , n26390 , n33032 );
nand ( n33034 , n20775 , n17468 );
nor ( n33035 , n17463 , n33034 );
or ( n33036 , n33035 , n17475 );
nand ( n33037 , n33035 , n17475 );
nand ( n33038 , n33036 , n33037 );
buf ( n33039 , n33038 );
nand ( n33040 , n33039 , n26393 );
buf ( n33041 , n17474 );
buf ( n33042 , n33041 );
not ( n33043 , n33042 );
not ( n33044 , n33043 );
nand ( n33045 , n26395 , n33044 );
nand ( n33046 , n17542 , n13880 );
nand ( n33047 , n33040 , n33045 , n33046 );
nor ( n33048 , n33033 , n33047 );
and ( n33049 , n33010 , n33027 , n33048 );
nand ( n33050 , n32993 , n33049 );
buf ( n33051 , n33050 );
buf ( n33052 , n33051 );
buf ( n33053 , n275554 );
buf ( n33054 , n275554 );
buf ( n33055 , n275554 );
not ( n33056 , n22798 );
not ( n33057 , n33056 );
and ( n33058 , n33057 , n29110 );
not ( n33059 , n33057 );
buf ( n33060 , n26598 );
not ( n33061 , n33060 );
not ( n33062 , n33061 );
not ( n33063 , n23958 );
not ( n33064 , n23979 );
not ( n33065 , n26627 );
not ( n33066 , n33065 );
nand ( n33067 , n23953 , n33066 );
nor ( n33068 , n33064 , n33067 );
nand ( n33069 , n21141 , n33068 );
nor ( n33070 , n33063 , n33069 );
not ( n33071 , n33070 );
or ( n33072 , n33062 , n33071 );
or ( n33073 , n33070 , n33061 );
nand ( n33074 , n33072 , n33073 );
buf ( n33075 , n33074 );
and ( n33076 , n33059 , n33075 );
nor ( n33077 , n33058 , n33076 );
or ( n33078 , n33077 , n19634 );
not ( n33079 , n27026 );
nand ( n33080 , n33079 , n27024 );
not ( n33081 , n33080 );
buf ( n33082 , n26986 );
nor ( n33083 , n26989 , n33082 );
not ( n33084 , n33083 );
not ( n33085 , n27020 );
or ( n33086 , n33084 , n33085 );
not ( n33087 , n33082 );
not ( n33088 , n33087 );
not ( n33089 , n27031 );
or ( n33090 , n33088 , n33089 );
not ( n33091 , n27023 );
nand ( n33092 , n33090 , n33091 );
not ( n33093 , n33092 );
nand ( n33094 , n33086 , n33093 );
not ( n33095 , n33094 );
or ( n33096 , n33081 , n33095 );
or ( n33097 , n33094 , n33080 );
nand ( n33098 , n33096 , n33097 );
buf ( n33099 , n33098 );
and ( n33100 , n29471 , n33099 );
and ( n33101 , n30137 , n28758 );
not ( n33102 , n30137 );
and ( n33103 , n33102 , n18592 );
nor ( n33104 , n33101 , n33103 );
not ( n33105 , n33104 );
not ( n33106 , n33105 );
not ( n33107 , n30612 );
or ( n33108 , n33106 , n33107 );
not ( n33109 , n28128 );
and ( n33110 , n27057 , n28133 );
nand ( n33111 , n24314 , n33110 );
not ( n33112 , n33111 );
or ( n33113 , n33109 , n33112 );
or ( n33114 , n33111 , n28128 );
nand ( n33115 , n33113 , n33114 );
buf ( n33116 , n33115 );
nand ( n33117 , n33116 , n31095 );
not ( n33118 , n27060 );
buf ( n33119 , n33118 );
buf ( n33120 , n33119 );
nand ( n33121 , n20563 , n33120 );
not ( n33122 , n28759 );
and ( n33123 , n33117 , n33121 , n33122 );
nand ( n33124 , n33108 , n33123 );
nor ( n33125 , n33100 , n33124 );
or ( n33126 , n26926 , n26838 );
not ( n33127 , n33126 );
nor ( n33128 , n26851 , n26847 );
not ( n33129 , n33128 );
not ( n33130 , n24204 );
or ( n33131 , n33129 , n33130 );
not ( n33132 , n26847 );
not ( n33133 , n33132 );
not ( n33134 , n26921 );
or ( n33135 , n33133 , n33134 );
nand ( n33136 , n33135 , n26924 );
not ( n33137 , n33136 );
nand ( n33138 , n33131 , n33137 );
not ( n33139 , n33138 );
or ( n33140 , n33127 , n33139 );
or ( n33141 , n33138 , n33126 );
nand ( n33142 , n33140 , n33141 );
buf ( n33143 , n33142 );
nand ( n33144 , n33143 , n20353 );
and ( n33145 , n33125 , n33144 );
nand ( n33146 , n33078 , n33145 );
buf ( n33147 , n33146 );
buf ( n33148 , n33147 );
not ( n33149 , n275550 );
buf ( n33150 , n33149 );
buf ( n33151 , n33150 );
buf ( n33152 , n275554 );
not ( n33153 , n275550 );
buf ( n33154 , n33153 );
buf ( n33155 , n33154 );
or ( n33156 , n29865 , n19216 );
not ( n33157 , n19353 );
nand ( n33158 , n30070 , n33157 );
nand ( n33159 , n30131 , n19360 );
nand ( n33160 , n30153 , n19318 );
nand ( n33161 , n30174 , n29075 );
not ( n33162 , n32248 );
nand ( n33163 , n33162 , n30177 );
nand ( n33164 , n19387 , n18424 );
and ( n33165 , n33160 , n33161 , n33163 , n33164 );
and ( n33166 , n33158 , n33159 , n33165 );
nand ( n33167 , n33156 , n33166 );
buf ( n33168 , n33167 );
buf ( n33169 , n33168 );
not ( n33170 , n275550 );
buf ( n33171 , n33170 );
buf ( n33172 , n33171 );
buf ( n33173 , n275554 );
not ( n33174 , n275929 );
buf ( n33175 , n33174 );
buf ( n33176 , n33175 );
not ( n33177 , n275925 );
buf ( n33178 , n33177 );
buf ( n33179 , n33178 );
buf ( n33180 , n275554 );
buf ( n33181 , n275554 );
buf ( n33182 , n275554 );
not ( n33183 , n29865 );
and ( n33184 , n33183 , n27845 );
not ( n33185 , n21001 );
not ( n33186 , n30070 );
or ( n33187 , n33185 , n33186 );
and ( n33188 , n30131 , n19358 );
not ( n33189 , n30177 );
not ( n33190 , n19219 );
or ( n33191 , n33189 , n33190 );
nand ( n33192 , n30174 , n19290 );
nand ( n33193 , n33191 , n33192 );
nor ( n33194 , n33188 , n33193 );
nand ( n33195 , n33187 , n33194 );
nor ( n33196 , n33184 , n33195 );
or ( n33197 , n33196 , n21030 );
nand ( n33198 , n21030 , n18429 );
nand ( n33199 , n33197 , n33198 );
buf ( n33200 , n33199 );
buf ( n33201 , n33200 );
buf ( n33202 , n275554 );
not ( n33203 , n275550 );
buf ( n33204 , n33203 );
buf ( n33205 , n33204 );
not ( n33206 , n275550 );
buf ( n33207 , n33206 );
buf ( n33208 , n33207 );
not ( n33209 , n21001 );
nand ( n33210 , n33132 , n26924 );
not ( n33211 , n33210 );
not ( n33212 , n26851 );
not ( n33213 , n33212 );
not ( n33214 , n24202 );
or ( n33215 , n33213 , n33214 );
not ( n33216 , n26921 );
nand ( n33217 , n33215 , n33216 );
not ( n33218 , n33217 );
or ( n33219 , n33211 , n33218 );
or ( n33220 , n33217 , n33210 );
nand ( n33221 , n33219 , n33220 );
buf ( n33222 , n33221 );
not ( n33223 , n33222 );
or ( n33224 , n33209 , n33223 );
nor ( n33225 , n33082 , n27023 );
not ( n33226 , n33225 );
nor ( n33227 , n24250 , n27031 );
nand ( n33228 , n24272 , n33227 , n24258 );
not ( n33229 , n27031 );
nand ( n33230 , n33229 , n26989 );
nand ( n33231 , n33228 , n33230 );
not ( n33232 , n33231 );
or ( n33233 , n33226 , n33232 );
or ( n33234 , n33231 , n33225 );
nand ( n33235 , n33233 , n33234 );
buf ( n33236 , n33235 );
and ( n33237 , n33236 , n19358 );
not ( n33238 , n19290 );
not ( n33239 , n28133 );
nand ( n33240 , n24314 , n27057 );
not ( n33241 , n33240 );
or ( n33242 , n33239 , n33241 );
or ( n33243 , n33240 , n28133 );
nand ( n33244 , n33242 , n33243 );
buf ( n33245 , n33244 );
not ( n33246 , n33245 );
or ( n33247 , n33238 , n33246 );
buf ( n33248 , n27058 );
not ( n33249 , n33248 );
not ( n33250 , n33249 );
nand ( n33251 , n19219 , n33250 );
nand ( n33252 , n33247 , n33251 );
nor ( n33253 , n33237 , n33252 );
nand ( n33254 , n33224 , n33253 );
not ( n33255 , n23977 );
not ( n33256 , n33255 );
and ( n33257 , n22798 , n33256 );
not ( n33258 , n22798 );
not ( n33259 , n33066 );
not ( n33260 , n29510 );
or ( n33261 , n33259 , n33260 );
and ( n33262 , n23978 , n23952 );
nand ( n33263 , n33262 , n23957 );
nand ( n33264 , n33065 , n29398 );
nor ( n33265 , n33263 , n29401 , n33264 );
and ( n33266 , n26554 , n33265 );
and ( n33267 , n33263 , n33066 );
nor ( n33268 , n33266 , n33267 );
nand ( n33269 , n33261 , n33268 );
buf ( n33270 , n33269 );
and ( n33271 , n33258 , n33270 );
nor ( n33272 , n33257 , n33271 );
nor ( n33273 , n33272 , n23991 );
nor ( n33274 , n33254 , n33273 );
or ( n33275 , n33274 , n24450 );
nand ( n33276 , n24450 , n18609 );
nand ( n33277 , n33275 , n33276 );
buf ( n33278 , n33277 );
buf ( n33279 , n33278 );
not ( n33280 , n275550 );
buf ( n33281 , n33280 );
buf ( n33282 , n33281 );
not ( n33283 , n275929 );
buf ( n33284 , n33283 );
buf ( n33285 , n33284 );
buf ( n33286 , n275554 );
buf ( n33287 , n275554 );
not ( n33288 , n275550 );
buf ( n33289 , n33288 );
buf ( n33290 , n33289 );
not ( n33291 , n275929 );
buf ( n33292 , n33291 );
buf ( n33293 , n33292 );
buf ( n33294 , n275554 );
buf ( n33295 , n275554 );
not ( n33296 , n26580 );
not ( n33297 , n33296 );
not ( n33298 , n33297 );
or ( n33299 , n33298 , n21774 );
nand ( n33300 , n21774 , n9696 );
nand ( n33301 , n33299 , n33300 );
buf ( n33302 , n33301 );
buf ( n33303 , n33302 );
buf ( n33304 , n275554 );
not ( n33305 , n275925 );
buf ( n33306 , n33305 );
buf ( n33307 , n33306 );
not ( n33308 , n275929 );
buf ( n33309 , n33308 );
buf ( n33310 , n33309 );
not ( n33311 , n275929 );
buf ( n33312 , n33311 );
buf ( n33313 , n33312 );
not ( n33314 , n275929 );
buf ( n33315 , n33314 );
buf ( n33316 , n33315 );
not ( n33317 , n275925 );
buf ( n33318 , n33317 );
buf ( n33319 , n33318 );
buf ( n33320 , n12226 );
buf ( n33321 , n33320 );
buf ( n33322 , n277453 );
buf ( n33323 , n33322 );
xor ( n33324 , n33321 , n33323 );
not ( n33325 , n33324 );
buf ( n33326 , n12415 );
buf ( n33327 , n277609 );
not ( n33328 , n33327 );
nor ( n33329 , n33326 , n33328 );
not ( n33330 , n33329 );
nand ( n33331 , n33330 , n31967 );
nor ( n33332 , n33331 , n31988 );
buf ( n33333 , n277386 );
not ( n33334 , n33333 );
buf ( n33335 , n277411 );
nand ( n33336 , n33334 , n33335 );
and ( n33337 , n33332 , n33336 );
and ( n33338 , n31978 , n33337 );
not ( n33339 , n33338 );
not ( n33340 , n27260 );
or ( n33341 , n33339 , n33340 );
not ( n33342 , n33337 );
not ( n33343 , n32011 );
or ( n33344 , n33342 , n33343 );
not ( n33345 , n33336 );
not ( n33346 , n32020 );
not ( n33347 , n33331 );
not ( n33348 , n33347 );
or ( n33349 , n33346 , n33348 );
not ( n33350 , n33329 );
not ( n33351 , n31969 );
and ( n33352 , n33350 , n33351 );
not ( n33353 , n33326 );
nor ( n33354 , n33353 , n33327 );
nor ( n33355 , n33352 , n33354 );
nand ( n33356 , n33349 , n33355 );
not ( n33357 , n33356 );
or ( n33358 , n33345 , n33357 );
not ( n33359 , n33335 );
nand ( n33360 , n33359 , n33333 );
nand ( n33361 , n33358 , n33360 );
not ( n33362 , n33361 );
nand ( n33363 , n33344 , n33362 );
not ( n33364 , n33363 );
nand ( n33365 , n33341 , n33364 );
not ( n33366 , n33365 );
or ( n33367 , n33325 , n33366 );
or ( n33368 , n33365 , n33324 );
nand ( n33369 , n33367 , n33368 );
buf ( n33370 , n33369 );
nand ( n33371 , n33370 , n31437 );
buf ( n33372 , n33322 );
buf ( n33373 , n33372 );
not ( n33374 , n33373 );
buf ( n33375 , n33320 );
buf ( n33376 , n33375 );
not ( n33377 , n33376 );
or ( n33378 , n33374 , n33377 );
buf ( n33379 , n33375 );
buf ( n33380 , n33372 );
or ( n33381 , n33379 , n33380 );
nand ( n33382 , n33378 , n33381 );
buf ( n33383 , n33382 );
buf ( n33384 , n33383 );
not ( n33385 , n33384 );
buf ( n33386 , n11774 );
buf ( n33387 , n33386 );
buf ( n33388 , n277609 );
buf ( n33389 , n33388 );
nor ( n33390 , n33387 , n33389 );
buf ( n33391 , n33390 );
buf ( n33392 , n33391 );
not ( n33393 , n33392 );
buf ( n33394 , n31804 );
nand ( n33395 , n33393 , n33394 );
buf ( n33396 , n33395 );
buf ( n33397 , n33396 );
buf ( n33398 , n31861 );
nor ( n33399 , n33397 , n33398 );
buf ( n33400 , n33399 );
buf ( n33401 , n33400 );
buf ( n33402 , n277411 );
buf ( n33403 , n33402 );
buf ( n33404 , n277386 );
buf ( n33405 , n33404 );
or ( n33406 , n33403 , n33405 );
buf ( n33407 , n33406 );
buf ( n33408 , n33407 );
and ( n33409 , n33401 , n33408 );
buf ( n33410 , n33409 );
buf ( n33411 , n33410 );
not ( n33412 , n33411 );
buf ( n33413 , n31838 );
nor ( n33414 , n33412 , n33413 );
buf ( n33415 , n33414 );
buf ( n33416 , n33415 );
not ( n33417 , n33416 );
buf ( n33418 , n27479 );
not ( n33419 , n33418 );
or ( n33420 , n33417 , n33419 );
buf ( n33421 , n33410 );
buf ( n33422 , n31922 );
and ( n33423 , n33421 , n33422 );
buf ( n33424 , n33407 );
not ( n33425 , n33424 );
buf ( n33426 , n31941 );
not ( n33427 , n33426 );
buf ( n33428 , n33396 );
not ( n33429 , n33428 );
buf ( n33430 , n33429 );
buf ( n33431 , n33430 );
not ( n33432 , n33431 );
or ( n33433 , n33427 , n33432 );
buf ( n33434 , n33391 );
not ( n33435 , n33434 );
buf ( n33436 , n31809 );
not ( n33437 , n33436 );
and ( n33438 , n33435 , n33437 );
buf ( n33439 , n33386 );
buf ( n33440 , n33388 );
and ( n33441 , n33439 , n33440 );
buf ( n33442 , n33441 );
buf ( n33443 , n33442 );
nor ( n33444 , n33438 , n33443 );
buf ( n33445 , n33444 );
buf ( n33446 , n33445 );
nand ( n33447 , n33433 , n33446 );
buf ( n33448 , n33447 );
buf ( n33449 , n33448 );
not ( n33450 , n33449 );
or ( n33451 , n33425 , n33450 );
buf ( n33452 , n33404 );
buf ( n33453 , n33402 );
nand ( n33454 , n33452 , n33453 );
buf ( n33455 , n33454 );
buf ( n33456 , n33455 );
nand ( n33457 , n33451 , n33456 );
buf ( n33458 , n33457 );
buf ( n33459 , n33458 );
nor ( n33460 , n33423 , n33459 );
buf ( n33461 , n33460 );
buf ( n33462 , n33461 );
nand ( n33463 , n33420 , n33462 );
buf ( n33464 , n33463 );
buf ( n33465 , n33464 );
not ( n33466 , n33465 );
or ( n33467 , n33385 , n33466 );
buf ( n33468 , n33464 );
buf ( n33469 , n33383 );
or ( n33470 , n33468 , n33469 );
nand ( n33471 , n33467 , n33470 );
buf ( n33472 , n33471 );
buf ( n33473 , n33472 );
nand ( n33474 , n33473 , n31422 );
not ( n33475 , n277453 );
not ( n33476 , n31460 );
or ( n33477 , n33475 , n33476 );
not ( n33478 , n32796 );
nor ( n33479 , n32792 , n33478 );
not ( n33480 , n33479 );
nand ( n33481 , n32045 , n32032 );
not ( n33482 , n33481 );
not ( n33483 , n33482 );
or ( n33484 , n33480 , n33483 );
not ( n33485 , n32794 );
not ( n33486 , n32045 );
or ( n33487 , n33485 , n33486 );
nand ( n33488 , n33487 , n33478 );
nand ( n33489 , n33484 , n33488 );
buf ( n33490 , n33489 );
nand ( n33491 , n20586 , n9163 );
nand ( n33492 , n33490 , n33491 );
or ( n33493 , n33492 , n28218 );
nand ( n33494 , n33477 , n33493 );
not ( n33495 , n28231 );
or ( n33496 , n33495 , n12160 );
not ( n33497 , n31453 );
not ( n33498 , n277423 );
and ( n33499 , n33497 , n33498 );
nand ( n33500 , n28236 , n9367 );
not ( n33501 , n33500 );
nor ( n33502 , n33499 , n33501 );
nand ( n33503 , n33496 , n33502 );
nor ( n33504 , n33494 , n33503 );
nand ( n33505 , n33371 , n33474 , n33504 );
buf ( n33506 , n33505 );
buf ( n33507 , n33506 );
buf ( n33508 , n275554 );
not ( n33509 , n13300 );
not ( n33510 , n27665 );
or ( n33511 , n33509 , n33510 );
not ( n33512 , n15555 );
or ( n33513 , n33512 , n27665 );
nand ( n33514 , n33511 , n33513 );
buf ( n33515 , n33514 );
buf ( n33516 , n33515 );
not ( n33517 , n22007 );
not ( n33518 , n12142 );
or ( n33519 , n33517 , n33518 );
not ( n33520 , n22051 );
nand ( n33521 , n33520 , n29231 );
nand ( n33522 , n33519 , n33521 );
nand ( n33523 , n29205 , n22000 );
nand ( n33524 , n29216 , n31005 );
nand ( n33525 , n22013 , n12280 );
nand ( n33526 , n33523 , n33524 , n33525 );
nor ( n33527 , n33522 , n33526 );
or ( n33528 , n33527 , n27640 );
nand ( n33529 , n27640 , n11130 );
nand ( n33530 , n33528 , n33529 );
buf ( n33531 , n33530 );
buf ( n33532 , n33531 );
not ( n33533 , n24639 );
not ( n33534 , n19201 );
and ( n33535 , n33533 , n33534 );
not ( n33536 , n19358 );
not ( n33537 , n24663 );
or ( n33538 , n33536 , n33537 );
nand ( n33539 , n19289 , n24440 );
and ( n33540 , n33539 , n24646 );
and ( n33541 , n24653 , n21001 );
nor ( n33542 , n33540 , n33541 );
nand ( n33543 , n33538 , n33542 );
nor ( n33544 , n33535 , n33543 );
or ( n33545 , n33544 , n24450 );
not ( n33546 , n24450 );
or ( n33547 , n33546 , n18296 );
nand ( n33548 , n33545 , n33547 );
buf ( n33549 , n33548 );
buf ( n33550 , n33549 );
buf ( n33551 , n275554 );
buf ( n33552 , n275554 );
buf ( n33553 , n275554 );
buf ( n33554 , n275554 );
buf ( n33555 , n275554 );
or ( n33556 , n27084 , n28146 );
nand ( n33557 , n24450 , n18557 );
nand ( n33558 , n33556 , n33557 );
buf ( n33559 , n33558 );
buf ( n33560 , n33559 );
buf ( n33561 , n275554 );
and ( n33562 , n31719 , n277653 );
not ( n33563 , n31719 );
not ( n33564 , n29599 );
buf ( n33565 , n31851 );
buf ( n33566 , n31931 );
not ( n33567 , n33566 );
buf ( n33568 , n33567 );
buf ( n33569 , n33568 );
nand ( n33570 , n33565 , n33569 );
buf ( n33571 , n33570 );
buf ( n33572 , n33571 );
not ( n33573 , n33572 );
buf ( n33574 , n31838 );
not ( n33575 , n33574 );
buf ( n33576 , n33575 );
buf ( n33577 , n33576 );
not ( n33578 , n33577 );
buf ( n33579 , n27479 );
not ( n33580 , n33579 );
or ( n33581 , n33578 , n33580 );
buf ( n33582 , n31922 );
not ( n33583 , n33582 );
buf ( n33584 , n33583 );
buf ( n33585 , n33584 );
nand ( n33586 , n33581 , n33585 );
buf ( n33587 , n33586 );
buf ( n33588 , n33587 );
not ( n33589 , n33588 );
or ( n33590 , n33573 , n33589 );
buf ( n33591 , n33587 );
buf ( n33592 , n33571 );
or ( n33593 , n33591 , n33592 );
nand ( n33594 , n33590 , n33593 );
buf ( n33595 , n33594 );
buf ( n33596 , n33595 );
not ( n33597 , n33596 );
or ( n33598 , n33564 , n33597 );
not ( n33599 , n31983 );
or ( n33600 , n33599 , n32015 );
not ( n33601 , n33600 );
not ( n33602 , n31978 );
not ( n33603 , n27260 );
or ( n33604 , n33602 , n33603 );
not ( n33605 , n32011 );
nand ( n33606 , n33604 , n33605 );
not ( n33607 , n33606 );
or ( n33608 , n33601 , n33607 );
or ( n33609 , n33606 , n33600 );
nand ( n33610 , n33608 , n33609 );
buf ( n33611 , n33610 );
and ( n33612 , n33611 , n23655 );
not ( n33613 , n23673 );
not ( n33614 , n32041 );
not ( n33615 , n33614 );
and ( n33616 , n30483 , n32801 );
not ( n33617 , n33616 );
or ( n33618 , n33615 , n33617 );
or ( n33619 , n33616 , n33614 );
nand ( n33620 , n33618 , n33619 );
buf ( n33621 , n33620 );
not ( n33622 , n33621 );
or ( n33623 , n33613 , n33622 );
and ( n33624 , n27520 , n12302 );
and ( n33625 , n22013 , n277696 );
nor ( n33626 , n33624 , n33625 );
nand ( n33627 , n33623 , n33626 );
nor ( n33628 , n33612 , n33627 );
nand ( n33629 , n33598 , n33628 );
and ( n33630 , n33563 , n33629 );
or ( n33631 , n33562 , n33630 );
buf ( n33632 , n33631 );
buf ( n33633 , n33632 );
and ( n33634 , n31468 , n275677 );
not ( n33635 , n13457 );
nor ( n33636 , n14830 , n33635 );
nor ( n33637 , n33634 , n33636 );
nand ( n33638 , n22914 , n23069 );
buf ( n33639 , n23134 );
not ( n33640 , n33639 );
buf ( n33641 , n23075 );
nor ( n33642 , n33640 , n33641 );
buf ( n33643 , n33642 );
buf ( n33644 , n33643 );
not ( n33645 , n33644 );
buf ( n33646 , n30540 );
buf ( n33647 , n23097 );
buf ( n33648 , n23066 );
and ( n33649 , n33646 , n33647 , n33648 );
buf ( n33650 , n23066 );
not ( n33651 , n33650 );
buf ( n33652 , n23126 );
not ( n33653 , n33652 );
or ( n33654 , n33651 , n33653 );
buf ( n33655 , n23109 );
nand ( n33656 , n33654 , n33655 );
buf ( n33657 , n33656 );
buf ( n33658 , n33657 );
nor ( n33659 , n33649 , n33658 );
buf ( n33660 , n33659 );
buf ( n33661 , n33660 );
not ( n33662 , n33661 );
or ( n33663 , n33645 , n33662 );
buf ( n33664 , n33660 );
buf ( n33665 , n33643 );
or ( n33666 , n33664 , n33665 );
nand ( n33667 , n33663 , n33666 );
buf ( n33668 , n33667 );
buf ( n33669 , n33668 );
nand ( n33670 , n22918 , n33669 );
buf ( n33671 , n23359 );
not ( n33672 , n33671 );
buf ( n33673 , n23302 );
nor ( n33674 , n33672 , n33673 );
buf ( n33675 , n33674 );
buf ( n33676 , n33675 );
not ( n33677 , n33676 );
buf ( n33678 , n30574 );
buf ( n33679 , n23322 );
buf ( n33680 , n23294 );
and ( n33681 , n33678 , n33679 , n33680 );
buf ( n33682 , n23294 );
not ( n33683 , n33682 );
buf ( n33684 , n23351 );
not ( n33685 , n33684 );
or ( n33686 , n33683 , n33685 );
buf ( n33687 , n23334 );
nand ( n33688 , n33686 , n33687 );
buf ( n33689 , n33688 );
buf ( n33690 , n33689 );
nor ( n33691 , n33681 , n33690 );
buf ( n33692 , n33691 );
buf ( n33693 , n33692 );
not ( n33694 , n33693 );
or ( n33695 , n33677 , n33694 );
buf ( n33696 , n33692 );
buf ( n33697 , n33675 );
or ( n33698 , n33696 , n33697 );
nand ( n33699 , n33695 , n33698 );
buf ( n33700 , n33699 );
buf ( n33701 , n33700 );
nand ( n33702 , n23152 , n33701 );
nand ( n33703 , n33637 , n33638 , n33670 , n33702 );
buf ( n33704 , n33703 );
buf ( n33705 , n33704 );
not ( n33706 , n277648 );
or ( n33707 , n33706 , n9158 );
nand ( n33708 , n9078 , n9158 );
nand ( n33709 , n33707 , n33708 );
buf ( n33710 , n33709 );
buf ( n33711 , n33710 );
and ( n33712 , n26516 , n26551 );
not ( n33713 , n26516 );
not ( n33714 , n27834 );
buf ( n33715 , n27818 );
not ( n33716 , n33715 );
not ( n33717 , n33716 );
or ( n33718 , n33714 , n33717 );
or ( n33719 , n33716 , n27834 );
nand ( n33720 , n33718 , n33719 );
buf ( n33721 , n33720 );
and ( n33722 , n33713 , n33721 );
nor ( n33723 , n33712 , n33722 );
or ( n33724 , n33723 , n32074 );
nand ( n33725 , n28095 , n28112 );
not ( n33726 , n33725 );
not ( n33727 , n28079 );
not ( n33728 , n33727 );
not ( n33729 , n27020 );
or ( n33730 , n33728 , n33729 );
not ( n33731 , n28109 );
nand ( n33732 , n33730 , n33731 );
not ( n33733 , n33732 );
or ( n33734 , n33726 , n33733 );
or ( n33735 , n33732 , n33725 );
nand ( n33736 , n33734 , n33735 );
buf ( n33737 , n33736 );
and ( n33738 , n33737 , n20515 );
not ( n33739 , n18788 );
and ( n33740 , n30144 , n33739 );
not ( n33741 , n30144 );
and ( n33742 , n33741 , n18789 );
nor ( n33743 , n33740 , n33742 );
not ( n33744 , n33743 );
not ( n33745 , n33744 );
not ( n33746 , n19650 );
or ( n33747 , n33745 , n33746 );
not ( n33748 , n30165 );
nand ( n33749 , n24314 , n30160 );
not ( n33750 , n33749 );
or ( n33751 , n33748 , n33750 );
or ( n33752 , n33749 , n30165 );
nand ( n33753 , n33751 , n33752 );
buf ( n33754 , n33753 );
nand ( n33755 , n33754 , n29492 );
nand ( n33756 , n20563 , n27932 );
nand ( n33757 , n30179 , n18789 );
and ( n33758 , n33755 , n33756 , n33757 );
nand ( n33759 , n33747 , n33758 );
nor ( n33760 , n33738 , n33759 );
not ( n33761 , n28023 );
nand ( n33762 , n33761 , n28041 );
not ( n33763 , n33762 );
not ( n33764 , n28014 );
not ( n33765 , n33764 );
not ( n33766 , n26915 );
or ( n33767 , n33765 , n33766 );
nand ( n33768 , n33767 , n28037 );
not ( n33769 , n33768 );
or ( n33770 , n33763 , n33769 );
or ( n33771 , n33768 , n33762 );
nand ( n33772 , n33770 , n33771 );
buf ( n33773 , n33772 );
nand ( n33774 , n33773 , n20353 );
and ( n33775 , n33760 , n33774 );
nand ( n33776 , n33724 , n33775 );
buf ( n33777 , n33776 );
buf ( n33778 , n33777 );
not ( n33779 , n275929 );
buf ( n33780 , n33779 );
buf ( n33781 , n33780 );
not ( n33782 , n275925 );
buf ( n33783 , n33782 );
buf ( n33784 , n33783 );
not ( n33785 , n33056 );
not ( n33786 , n23981 );
not ( n33787 , n23959 );
or ( n33788 , n33786 , n33787 );
or ( n33789 , n23959 , n23981 );
nand ( n33790 , n33788 , n33789 );
buf ( n33791 , n33790 );
not ( n33792 , n33791 );
or ( n33793 , n33785 , n33792 );
buf ( n33794 , n21111 );
nand ( n33795 , n33794 , n22798 );
nand ( n33796 , n33793 , n33795 );
not ( n33797 , n33796 );
or ( n33798 , n33797 , n19216 );
nand ( n33799 , n24161 , n24207 );
not ( n33800 , n33799 );
not ( n33801 , n30043 );
or ( n33802 , n33800 , n33801 );
or ( n33803 , n30043 , n33799 );
nand ( n33804 , n33802 , n33803 );
buf ( n33805 , n33804 );
not ( n33806 , n33805 );
not ( n33807 , n33806 );
not ( n33808 , n19353 );
and ( n33809 , n33807 , n33808 );
not ( n33810 , n19360 );
nand ( n33811 , n24228 , n24253 );
not ( n33812 , n33811 );
not ( n33813 , n28092 );
or ( n33814 , n33812 , n33813 );
or ( n33815 , n28092 , n33811 );
nand ( n33816 , n33814 , n33815 );
buf ( n33817 , n33816 );
not ( n33818 , n33817 );
or ( n33819 , n33810 , n33818 );
not ( n33820 , n24304 );
not ( n33821 , n28124 );
not ( n33822 , n33821 );
or ( n33823 , n33820 , n33822 );
or ( n33824 , n33821 , n24304 );
nand ( n33825 , n33823 , n33824 );
buf ( n33826 , n33825 );
nand ( n33827 , n33826 , n29075 );
not ( n33828 , n29537 );
and ( n33829 , n29480 , n18958 );
not ( n33830 , n29480 );
and ( n33831 , n33830 , n29481 );
nor ( n33832 , n33829 , n33831 );
not ( n33833 , n33832 );
and ( n33834 , n33828 , n33833 );
buf ( n33835 , n24303 );
buf ( n33836 , n33835 );
buf ( n33837 , n33836 );
and ( n33838 , n19221 , n33837 );
nor ( n33839 , n33834 , n33838 );
not ( n33840 , n19388 );
nand ( n33841 , n33840 , n18968 );
and ( n33842 , n33827 , n33839 , n33841 );
nand ( n33843 , n33819 , n33842 );
nor ( n33844 , n33809 , n33843 );
nand ( n33845 , n33798 , n33844 );
buf ( n33846 , n33845 );
buf ( n33847 , n33846 );
not ( n33848 , n14861 );
or ( n33849 , n17547 , n33848 );
nand ( n33850 , n33849 , n21694 );
buf ( n33851 , n33850 );
buf ( n33852 , n33851 );
not ( n33853 , n275929 );
buf ( n33854 , n33853 );
buf ( n33855 , n33854 );
not ( n33856 , n275550 );
buf ( n33857 , n33856 );
buf ( n33858 , n33857 );
not ( n33859 , n275550 );
buf ( n33860 , n33859 );
buf ( n33861 , n33860 );
buf ( n33862 , n275554 );
buf ( n33863 , n275554 );
nand ( n33864 , n28213 , n28407 );
nand ( n33865 , n28194 , n28427 );
nand ( n33866 , n28458 , n12141 );
and ( n33867 , n33864 , n33865 , n33866 );
nand ( n33868 , n28228 , n28438 );
nand ( n33869 , n29234 , n11006 );
nand ( n33870 , n28453 , n12318 );
nand ( n33871 , n33867 , n33868 , n33869 , n33870 );
buf ( n33872 , n33871 );
buf ( n33873 , n33872 );
nand ( n33874 , n23602 , n28306 );
not ( n33875 , n28329 );
nand ( n33876 , n23654 , n33875 );
and ( n33877 , n31449 , n23671 );
and ( n33878 , n28350 , n12257 );
nor ( n33879 , n33877 , n33878 );
and ( n33880 , n28231 , n23676 );
or ( n33881 , n28354 , n11521 );
not ( n33882 , n11535 );
nand ( n33883 , n28357 , n33882 );
nand ( n33884 , n33881 , n33883 );
nor ( n33885 , n33880 , n33884 );
nand ( n33886 , n33874 , n33876 , n33879 , n33885 );
buf ( n33887 , n33886 );
buf ( n33888 , n33887 );
and ( n33889 , n13374 , n14056 );
not ( n33890 , n13374 );
nand ( n33891 , n14797 , n14058 , n24486 );
not ( n33892 , n33891 );
nand ( n33893 , n33892 , n23826 );
not ( n33894 , n24768 );
and ( n33895 , n33893 , n33894 );
not ( n33896 , n33893 );
and ( n33897 , n33896 , n24768 );
nor ( n33898 , n33895 , n33897 );
buf ( n33899 , n33898 );
and ( n33900 , n33890 , n33899 );
nor ( n33901 , n33889 , n33900 );
or ( n33902 , n33901 , n14909 );
or ( n33903 , n30290 , n30307 );
not ( n33904 , n33903 );
not ( n33905 , n24551 );
nor ( n33906 , n33905 , n24556 );
not ( n33907 , n33906 );
nor ( n33908 , n33907 , n16140 );
not ( n33909 , n33908 );
not ( n33910 , n16913 );
or ( n33911 , n33909 , n33910 );
not ( n33912 , n33906 );
not ( n33913 , n16943 );
or ( n33914 , n33912 , n33913 );
not ( n33915 , n24551 );
not ( n33916 , n24565 );
or ( n33917 , n33915 , n33916 );
nand ( n33918 , n33917 , n24552 );
not ( n33919 , n33918 );
nand ( n33920 , n33914 , n33919 );
not ( n33921 , n33920 );
nand ( n33922 , n33911 , n33921 );
not ( n33923 , n33922 );
or ( n33924 , n33904 , n33923 );
or ( n33925 , n33922 , n33903 );
nand ( n33926 , n33924 , n33925 );
buf ( n33927 , n33926 );
nand ( n33928 , n33927 , n16970 );
or ( n33929 , n30335 , n30352 );
not ( n33930 , n33929 );
nand ( n33931 , n24590 , n24586 );
nor ( n33932 , n17090 , n33931 );
not ( n33933 , n33932 );
not ( n33934 , n17362 );
or ( n33935 , n33933 , n33934 );
not ( n33936 , n17389 );
not ( n33937 , n33931 );
and ( n33938 , n33936 , n33937 );
not ( n33939 , n24586 );
not ( n33940 , n24600 );
or ( n33941 , n33939 , n33940 );
nand ( n33942 , n33941 , n24587 );
nor ( n33943 , n33938 , n33942 );
nand ( n33944 , n33935 , n33943 );
not ( n33945 , n33944 );
or ( n33946 , n33930 , n33945 );
or ( n33947 , n33944 , n33929 );
nand ( n33948 , n33946 , n33947 );
buf ( n33949 , n33948 );
and ( n33950 , n33949 , n17405 );
nand ( n33951 , n17534 , n14002 );
not ( n33952 , n14033 );
nor ( n33953 , n33951 , n33952 );
and ( n33954 , n33953 , n14714 );
not ( n33955 , n33953 );
not ( n33956 , n14713 );
and ( n33957 , n33955 , n33956 );
nor ( n33958 , n33954 , n33957 );
nand ( n33959 , n33958 , n17545 );
not ( n33960 , n23873 );
nand ( n33961 , n17489 , n24615 , n24895 );
nor ( n33962 , n33961 , n17478 , n17481 , n17473 );
nand ( n33963 , n33960 , n17472 , n33962 );
nor ( n33964 , n17463 , n33963 );
or ( n33965 , n33964 , n24892 );
nand ( n33966 , n33964 , n24892 );
nand ( n33967 , n33965 , n33966 );
buf ( n33968 , n33967 );
nand ( n33969 , n32339 , n33968 );
nand ( n33970 , n20785 , n24891 );
nand ( n33971 , n17562 , n14700 );
nand ( n33972 , n33959 , n33969 , n33970 , n33971 );
nor ( n33973 , n33950 , n33972 );
and ( n33974 , n33928 , n33973 );
nand ( n33975 , n33902 , n33974 );
buf ( n33976 , n33975 );
buf ( n33977 , n33976 );
buf ( n33978 , n275554 );
buf ( n33979 , n275554 );
buf ( n33980 , n18330 );
and ( n33981 , n22798 , n33980 );
not ( n33982 , n22798 );
buf ( n33983 , n19524 );
not ( n33984 , n33983 );
nand ( n33985 , n20978 , n20973 );
not ( n33986 , n33985 );
or ( n33987 , n33984 , n33986 );
not ( n33988 , n20974 );
nand ( n33989 , n20978 , n33988 );
or ( n33990 , n33989 , n33983 );
nand ( n33991 , n33987 , n33990 );
buf ( n33992 , n33991 );
and ( n33993 , n33982 , n33992 );
nor ( n33994 , n33981 , n33993 );
not ( n33995 , n33994 );
and ( n33996 , n33995 , n20987 );
not ( n33997 , n21001 );
not ( n33998 , n20328 );
buf ( n33999 , n20318 );
nand ( n34000 , n33998 , n33999 );
not ( n34001 , n34000 );
not ( n34002 , n20308 );
nand ( n34003 , n34002 , n20323 );
not ( n34004 , n34003 );
or ( n34005 , n34001 , n34004 );
or ( n34006 , n34003 , n34000 );
nand ( n34007 , n34005 , n34006 );
buf ( n34008 , n34007 );
not ( n34009 , n34008 );
or ( n34010 , n33997 , n34009 );
not ( n34011 , n24263 );
not ( n34012 , n34011 );
nand ( n34013 , n20413 , n20424 );
not ( n34014 , n34013 );
or ( n34015 , n34012 , n34014 );
or ( n34016 , n34013 , n34011 );
nand ( n34017 , n34015 , n34016 );
buf ( n34018 , n34017 );
and ( n34019 , n34018 , n19358 );
not ( n34020 , n19290 );
not ( n34021 , n20541 );
nand ( n34022 , n34021 , n20539 );
xor ( n34023 , n34022 , n20543 );
buf ( n34024 , n34023 );
not ( n34025 , n34024 );
or ( n34026 , n34020 , n34025 );
buf ( n34027 , n20542 );
buf ( n34028 , n34027 );
buf ( n34029 , n34028 );
not ( n34030 , n34029 );
or ( n34031 , n24440 , n34030 );
nand ( n34032 , n34026 , n34031 );
nor ( n34033 , n34019 , n34032 );
nand ( n34034 , n34010 , n34033 );
nor ( n34035 , n33996 , n34034 );
or ( n34036 , n34035 , n24450 );
nand ( n34037 , n24450 , n18857 );
nand ( n34038 , n34036 , n34037 );
buf ( n34039 , n34038 );
buf ( n34040 , n34039 );
buf ( n34041 , n23498 );
buf ( n34042 , n29334 );
nand ( n34043 , n34041 , n34042 );
buf ( n34044 , n34043 );
buf ( n34045 , n34044 );
not ( n34046 , n34045 );
buf ( n34047 , n23568 );
not ( n34048 , n34047 );
or ( n34049 , n34046 , n34048 );
buf ( n34050 , n23568 );
buf ( n34051 , n34044 );
or ( n34052 , n34050 , n34051 );
nand ( n34053 , n34049 , n34052 );
buf ( n34054 , n34053 );
buf ( n34055 , n34054 );
nand ( n34056 , n34055 , n28306 );
nand ( n34057 , n23616 , n29353 );
not ( n34058 , n34057 );
not ( n34059 , n23638 );
or ( n34060 , n34058 , n34059 );
or ( n34061 , n23638 , n34057 );
nand ( n34062 , n34060 , n34061 );
buf ( n34063 , n34062 );
nand ( n34064 , n34063 , n33875 );
buf ( n34065 , n23660 );
not ( n34066 , n34065 );
not ( n34067 , n34066 );
nor ( n34068 , n22042 , n22044 );
not ( n34069 , n34068 );
or ( n34070 , n34067 , n34069 );
or ( n34071 , n34068 , n34066 );
nand ( n34072 , n34070 , n34071 );
buf ( n34073 , n34072 );
and ( n34074 , n28219 , n34073 );
and ( n34075 , n28242 , n12271 );
nor ( n34076 , n34074 , n34075 );
and ( n34077 , n31451 , n12126 );
or ( n34078 , n31453 , n11601 );
nand ( n34079 , n28236 , n11607 );
nand ( n34080 , n34078 , n34079 );
nor ( n34081 , n34077 , n34080 );
nand ( n34082 , n34056 , n34064 , n34076 , n34081 );
buf ( n34083 , n34082 );
buf ( n34084 , n34083 );
not ( n34085 , n275550 );
buf ( n34086 , n34085 );
buf ( n34087 , n34086 );
not ( n34088 , n275550 );
buf ( n34089 , n34088 );
buf ( n34090 , n34089 );
buf ( n34091 , n275554 );
buf ( n34092 , n14250 );
not ( n34093 , n34092 );
or ( n34094 , n34093 , n28252 );
nand ( n34095 , n29044 , n9540 );
nand ( n34096 , n34094 , n34095 );
buf ( n34097 , n34096 );
buf ( n34098 , n34097 );
not ( n34099 , n275550 );
buf ( n34100 , n34099 );
buf ( n34101 , n34100 );
buf ( n34102 , n275554 );
or ( n34103 , n24639 , n19634 );
not ( n34104 , n19648 );
nand ( n34105 , n34104 , n19639 );
nand ( n34106 , n34105 , n18283 );
not ( n34107 , n24646 );
nor ( n34108 , n34107 , n19646 );
not ( n34109 , n24653 );
nor ( n34110 , n34109 , n19638 );
not ( n34111 , n24663 );
nor ( n34112 , n34111 , n19647 );
nor ( n34113 , n34108 , n34110 , n34112 );
nand ( n34114 , n34103 , n34106 , n34113 );
buf ( n34115 , n34114 );
buf ( n34116 , n34115 );
and ( n34117 , n21030 , n19042 );
not ( n34118 , n21030 );
not ( n34119 , n33716 );
not ( n34120 , n34119 );
nand ( n34121 , n29821 , n29857 );
not ( n34122 , n34121 );
buf ( n34123 , n18849 );
not ( n34124 , n34123 );
buf ( n34125 , n34124 );
buf ( n34126 , n34125 );
not ( n34127 , n34126 );
buf ( n34128 , n29804 );
buf ( n34129 , n18467 );
not ( n34130 , n34129 );
buf ( n34131 , n34130 );
buf ( n34132 , n34131 );
and ( n34133 , n34128 , n34132 );
buf ( n34134 , n34133 );
buf ( n34135 , n34134 );
buf ( n34136 , n27767 );
nand ( n34137 , n34135 , n34136 );
buf ( n34138 , n34137 );
buf ( n34139 , n34138 );
buf ( n34140 , n23914 );
nor ( n34141 , n34139 , n34140 );
buf ( n34142 , n34141 );
buf ( n34143 , n34142 );
not ( n34144 , n34143 );
or ( n34145 , n34127 , n34144 );
buf ( n34146 , n34142 );
buf ( n34147 , n34125 );
or ( n34148 , n34146 , n34147 );
nand ( n34149 , n34145 , n34148 );
buf ( n34150 , n34149 );
buf ( n34151 , n34150 );
buf ( n34152 , n34151 );
not ( n34153 , n34152 );
not ( n34154 , n34153 );
buf ( n34155 , n34154 );
nand ( n34156 , n34122 , n34155 );
buf ( n34157 , n19066 );
buf ( n34158 , n34157 );
buf ( n34159 , n34158 );
nor ( n34160 , n34156 , n29825 , n34159 );
not ( n34161 , n34160 );
or ( n34162 , n34120 , n34161 );
not ( n34163 , n34156 );
not ( n34164 , n34163 );
buf ( n34165 , n29831 );
not ( n34166 , n34165 );
or ( n34167 , n34164 , n34166 );
nand ( n34168 , n34167 , n34159 );
nand ( n34169 , n34162 , n34168 );
buf ( n34170 , n34169 );
or ( n34171 , n18208 , n19151 );
nand ( n34172 , n34171 , n25051 );
and ( n34173 , n20987 , n34172 );
nand ( n34174 , n34170 , n34173 );
buf ( n34175 , n277457 );
buf ( n34176 , n34175 );
not ( n34177 , n34176 );
buf ( n34178 , n277495 );
buf ( n34179 , n34178 );
not ( n34180 , n34179 );
and ( n34181 , n34177 , n34180 );
buf ( n34182 , n34175 );
buf ( n34183 , n34178 );
and ( n34184 , n34182 , n34183 );
nor ( n34185 , n34181 , n34184 );
buf ( n34186 , n34185 );
buf ( n34187 , n34186 );
not ( n34188 , n34187 );
buf ( n34189 , n22592 );
buf ( n34190 , n22415 );
buf ( n34191 , n22452 );
buf ( n34192 , n22470 );
not ( n34193 , n34192 );
buf ( n34194 , n22767 );
nor ( n34195 , n34193 , n34194 );
buf ( n34196 , n34195 );
buf ( n34197 , n34196 );
and ( n34198 , n34191 , n34197 );
buf ( n34199 , n34198 );
buf ( n34200 , n34199 );
and ( n34201 , n34190 , n34200 );
buf ( n34202 , n34201 );
buf ( n34203 , n34202 );
and ( n34204 , n34189 , n34203 );
buf ( n34205 , n34199 );
not ( n34206 , n34205 );
buf ( n34207 , n22687 );
not ( n34208 , n34207 );
or ( n34209 , n34206 , n34208 );
buf ( n34210 , n22732 );
buf ( n34211 , n34196 );
and ( n34212 , n34210 , n34211 );
buf ( n34213 , n22751 );
buf ( n34214 , n22767 );
or ( n34215 , n34213 , n34214 );
buf ( n34216 , n22773 );
nand ( n34217 , n34215 , n34216 );
buf ( n34218 , n34217 );
buf ( n34219 , n34218 );
nor ( n34220 , n34212 , n34219 );
buf ( n34221 , n34220 );
buf ( n34222 , n34221 );
nand ( n34223 , n34209 , n34222 );
buf ( n34224 , n34223 );
buf ( n34225 , n34224 );
nor ( n34226 , n34204 , n34225 );
buf ( n34227 , n34226 );
buf ( n34228 , n34227 );
not ( n34229 , n34228 );
or ( n34230 , n34188 , n34229 );
buf ( n34231 , n34227 );
buf ( n34232 , n34186 );
or ( n34233 , n34231 , n34232 );
nand ( n34234 , n34230 , n34233 );
buf ( n34235 , n34234 );
buf ( n34236 , n34235 );
not ( n34237 , n34236 );
or ( n34238 , n34237 , n277910 );
nand ( n34239 , n277983 , n277457 );
nand ( n34240 , n34238 , n34239 );
and ( n34241 , n25049 , n34240 );
buf ( n34242 , n34241 );
not ( n34243 , n34242 );
and ( n34244 , n25051 , n22791 );
buf ( n34245 , n34244 );
not ( n34246 , n34245 );
and ( n34247 , n25049 , n30237 );
buf ( n34248 , n34247 );
not ( n34249 , n34248 );
not ( n34250 , n34249 );
buf ( n34251 , n34250 );
nor ( n34252 , n30156 , n34251 );
nand ( n34253 , n34246 , n30160 , n34252 , n30167 );
nor ( n34254 , n28124 , n34253 );
not ( n34255 , n34254 );
or ( n34256 , n34243 , n34255 );
or ( n34257 , n34254 , n34242 );
nand ( n34258 , n34256 , n34257 );
buf ( n34259 , n34258 );
and ( n34260 , n34259 , n19290 );
and ( n34261 , n19219 , n34241 );
nor ( n34262 , n34260 , n34261 );
nand ( n34263 , n34174 , n34262 );
and ( n34264 , n34118 , n34263 );
or ( n34265 , n34117 , n34264 );
buf ( n34266 , n34265 );
buf ( n34267 , n34266 );
not ( n34268 , n275929 );
buf ( n34269 , n34268 );
buf ( n34270 , n34269 );
or ( n34271 , n22816 , n32073 );
and ( n34272 , n22858 , n20353 );
or ( n34273 , n20562 , n22872 );
or ( n34274 , n20559 , n22865 );
not ( n34275 , n32496 );
nand ( n34276 , n34273 , n34274 , n34275 );
nor ( n34277 , n34272 , n34276 );
nand ( n34278 , n22836 , n20515 );
not ( n34279 , n18887 );
not ( n34280 , n19656 );
not ( n34281 , n34280 );
or ( n34282 , n34279 , n34281 );
or ( n34283 , n34280 , n18887 );
nand ( n34284 , n34282 , n34283 );
nand ( n34285 , n19650 , n34284 );
and ( n34286 , n34277 , n34278 , n34285 );
nand ( n34287 , n34271 , n34286 );
buf ( n34288 , n34287 );
buf ( n34289 , n34288 );
buf ( n34290 , n275554 );
and ( n34291 , n23706 , n277758 );
not ( n34292 , n23706 );
and ( n34293 , n34292 , n30996 );
or ( n34294 , n34291 , n34293 );
buf ( n34295 , n34294 );
buf ( n34296 , n34295 );
not ( n34297 , n275550 );
buf ( n34298 , n34297 );
buf ( n34299 , n34298 );
not ( n34300 , n28408 );
buf ( n34301 , n34300 );
not ( n34302 , n34301 );
not ( n34303 , n34302 );
not ( n34304 , n30906 );
or ( n34305 , n34303 , n34304 );
and ( n34306 , n30961 , n28430 );
not ( n34307 , n29162 );
nand ( n34308 , n30988 , n34307 );
nand ( n34309 , n28451 , n277771 );
nand ( n34310 , n29171 , n12185 );
not ( n34311 , n32757 );
and ( n34312 , n34311 , n12370 );
not ( n34313 , n9159 );
and ( n34314 , n34313 , n9274 );
nor ( n34315 , n34312 , n34314 );
and ( n34316 , n34310 , n34315 );
nand ( n34317 , n34308 , n34309 , n34316 );
nor ( n34318 , n34306 , n34317 );
nand ( n34319 , n34305 , n34318 );
buf ( n34320 , n34319 );
buf ( n34321 , n34320 );
buf ( n34322 , n275554 );
buf ( n34323 , n30406 );
buf ( n34324 , n30430 );
nand ( n34325 , n34323 , n34324 );
buf ( n34326 , n34325 );
buf ( n34327 , n34326 );
not ( n34328 , n34327 );
buf ( n34329 , n28266 );
buf ( n34330 , n30401 );
buf ( n34331 , n34330 );
nor ( n34332 , n34329 , n34331 );
buf ( n34333 , n34332 );
buf ( n34334 , n34333 );
not ( n34335 , n34334 );
buf ( n34336 , n23568 );
not ( n34337 , n34336 );
or ( n34338 , n34335 , n34337 );
buf ( n34339 , n28383 );
buf ( n34340 , n34330 );
not ( n34341 , n34340 );
buf ( n34342 , n34341 );
buf ( n34343 , n34342 );
and ( n34344 , n34339 , n34343 );
buf ( n34345 , n27446 );
nor ( n34346 , n34344 , n34345 );
buf ( n34347 , n34346 );
buf ( n34348 , n34347 );
nand ( n34349 , n34338 , n34348 );
buf ( n34350 , n34349 );
buf ( n34351 , n34350 );
not ( n34352 , n34351 );
or ( n34353 , n34328 , n34352 );
buf ( n34354 , n34350 );
buf ( n34355 , n34326 );
or ( n34356 , n34354 , n34355 );
nand ( n34357 , n34353 , n34356 );
buf ( n34358 , n34357 );
buf ( n34359 , n34358 );
nand ( n34360 , n34359 , n28408 );
nand ( n34361 , n27223 , n30464 );
not ( n34362 , n34361 );
buf ( n34363 , n30453 );
nor ( n34364 , n28312 , n34363 );
not ( n34365 , n34364 );
not ( n34366 , n23638 );
or ( n34367 , n34365 , n34366 );
not ( n34368 , n34363 );
and ( n34369 , n28318 , n34368 );
nor ( n34370 , n34369 , n27249 );
nand ( n34371 , n34367 , n34370 );
not ( n34372 , n34371 );
or ( n34373 , n34362 , n34372 );
or ( n34374 , n34371 , n34361 );
nand ( n34375 , n34373 , n34374 );
buf ( n34376 , n34375 );
nand ( n34377 , n34376 , n28430 );
nand ( n34378 , n28344 , n28339 );
nor ( n34379 , n34378 , n30734 );
nand ( n34380 , n28336 , n34379 );
buf ( n34381 , n27497 );
xnor ( n34382 , n34380 , n34381 );
buf ( n34383 , n34382 );
nand ( n34384 , n34383 , n28440 );
nand ( n34385 , n28451 , n11246 );
and ( n34386 , n28455 , n12351 );
not ( n34387 , n12205 );
or ( n34388 , n28459 , n34387 );
nand ( n34389 , n20649 , n9303 );
nand ( n34390 , n34388 , n34389 );
nor ( n34391 , n34386 , n34390 );
and ( n34392 , n34384 , n34385 , n34391 );
nand ( n34393 , n34360 , n34377 , n34392 );
buf ( n34394 , n34393 );
buf ( n34395 , n34394 );
buf ( n34396 , n275554 );
not ( n34397 , n275550 );
buf ( n34398 , n34397 );
buf ( n34399 , n34398 );
nand ( n34400 , n24792 , n24486 );
not ( n34401 , n24816 );
nand ( n34402 , n34401 , n14797 , n14058 );
nor ( n34403 , n34400 , n34402 );
not ( n34404 , n34403 );
not ( n34405 , n23826 );
or ( n34406 , n34404 , n34405 );
and ( n34407 , n23827 , n24816 );
not ( n34408 , n24816 );
not ( n34409 , n34400 );
or ( n34410 , n34408 , n34409 );
not ( n34411 , n34401 );
not ( n34412 , n14797 );
and ( n34413 , n34411 , n34412 );
and ( n34414 , n14059 , n24816 );
nor ( n34415 , n34413 , n34414 );
nand ( n34416 , n34410 , n34415 );
nor ( n34417 , n34407 , n34416 );
nand ( n34418 , n34406 , n34417 );
buf ( n34419 , n34418 );
and ( n34420 , n34419 , n24835 );
not ( n34421 , n24767 );
nor ( n34422 , n34421 , n23386 );
nor ( n34423 , n34420 , n34422 );
not ( n34424 , n34423 );
and ( n34425 , n34424 , n26440 );
not ( n34426 , n20889 );
nor ( n34427 , n30267 , n30260 );
not ( n34428 , n34427 );
buf ( n34429 , n24939 );
not ( n34430 , n34429 );
buf ( n34431 , n14664 );
buf ( n34432 , n34431 );
buf ( n34433 , n34432 );
not ( n34434 , n34433 );
or ( n34435 , n34430 , n34434 );
or ( n34436 , n34433 , n34429 );
nand ( n34437 , n34435 , n34436 );
not ( n34438 , n34437 );
or ( n34439 , n34428 , n34438 );
or ( n34440 , n34427 , n34437 );
nand ( n34441 , n34439 , n34440 );
not ( n34442 , n34441 );
nor ( n34443 , n30292 , n30276 );
and ( n34444 , n16139 , n34443 );
not ( n34445 , n34444 );
not ( n34446 , n16913 );
or ( n34447 , n34445 , n34446 );
not ( n34448 , n34443 );
not ( n34449 , n16943 );
or ( n34450 , n34448 , n34449 );
not ( n34451 , n30277 );
not ( n34452 , n30309 );
or ( n34453 , n34451 , n34452 );
nand ( n34454 , n34453 , n30278 );
not ( n34455 , n34454 );
nand ( n34456 , n34450 , n34455 );
not ( n34457 , n34456 );
nand ( n34458 , n34447 , n34457 );
not ( n34459 , n34458 );
or ( n34460 , n34442 , n34459 );
or ( n34461 , n34458 , n34441 );
nand ( n34462 , n34460 , n34461 );
buf ( n34463 , n34462 );
not ( n34464 , n34463 );
or ( n34465 , n34426 , n34464 );
buf ( n34466 , n24939 );
not ( n34467 , n34466 );
buf ( n34468 , n34432 );
not ( n34469 , n34468 );
not ( n34470 , n34469 );
or ( n34471 , n34467 , n34470 );
or ( n34472 , n34469 , n34466 );
nand ( n34473 , n34471 , n34472 );
not ( n34474 , n34473 );
and ( n34475 , n30321 , n30323 );
not ( n34476 , n34475 );
or ( n34477 , n34474 , n34476 );
or ( n34478 , n34475 , n34473 );
nand ( n34479 , n34477 , n34478 );
not ( n34480 , n34479 );
nand ( n34481 , n30337 , n30329 );
nor ( n34482 , n17090 , n34481 );
not ( n34483 , n34482 );
not ( n34484 , n17362 );
or ( n34485 , n34483 , n34484 );
not ( n34486 , n17389 );
not ( n34487 , n34481 );
and ( n34488 , n34486 , n34487 );
not ( n34489 , n30329 );
not ( n34490 , n30354 );
or ( n34491 , n34489 , n34490 );
nand ( n34492 , n34491 , n30330 );
nor ( n34493 , n34488 , n34492 );
nand ( n34494 , n34485 , n34493 );
not ( n34495 , n34494 );
or ( n34496 , n34480 , n34495 );
or ( n34497 , n34494 , n34479 );
nand ( n34498 , n34496 , n34497 );
buf ( n34499 , n34498 );
and ( n34500 , n34499 , n24711 );
not ( n34501 , n17409 );
not ( n34502 , n24940 );
nor ( n34503 , n24896 , n24938 );
nand ( n34504 , n23875 , n34503 );
nor ( n34505 , n17463 , n34504 );
not ( n34506 , n34505 );
or ( n34507 , n34502 , n34506 );
or ( n34508 , n34505 , n24940 );
nand ( n34509 , n34507 , n34508 );
buf ( n34510 , n34509 );
not ( n34511 , n34510 );
or ( n34512 , n34501 , n34511 );
nand ( n34513 , n20940 , n24939 );
nand ( n34514 , n34512 , n34513 );
nor ( n34515 , n34500 , n34514 );
nand ( n34516 , n34465 , n34515 );
nor ( n34517 , n34425 , n34516 );
or ( n34518 , n34517 , n20951 );
nand ( n34519 , n20950 , n14662 );
nand ( n34520 , n34518 , n34519 );
buf ( n34521 , n34520 );
buf ( n34522 , n34521 );
buf ( n34523 , n275554 );
buf ( n34524 , n275554 );
buf ( n34525 , n12823 );
not ( n34526 , n34525 );
not ( n34527 , n14830 );
or ( n34528 , n34526 , n34527 );
not ( n34529 , n15826 );
or ( n34530 , n34529 , n23807 );
nand ( n34531 , n34528 , n34530 );
buf ( n34532 , n34531 );
buf ( n34533 , n34532 );
not ( n34534 , n275929 );
buf ( n34535 , n34534 );
buf ( n34536 , n34535 );
and ( n34537 , n9158 , n9021 );
not ( n34538 , n9158 );
and ( n34539 , n34538 , n277497 );
or ( n34540 , n34537 , n34539 );
buf ( n34541 , n34540 );
buf ( n34542 , n34541 );
nand ( n34543 , n25064 , n18115 );
not ( n34544 , n25389 );
buf ( n34545 , n25195 );
not ( n34546 , n34545 );
buf ( n34547 , n25212 );
buf ( n34548 , n25202 );
nand ( n34549 , n34547 , n34548 );
buf ( n34550 , n34549 );
buf ( n34551 , n34550 );
not ( n34552 , n34551 );
or ( n34553 , n34546 , n34552 );
buf ( n34554 , n34550 );
buf ( n34555 , n25195 );
or ( n34556 , n34554 , n34555 );
nand ( n34557 , n34553 , n34556 );
buf ( n34558 , n34557 );
buf ( n34559 , n34558 );
and ( n34560 , n34544 , n34559 );
not ( n34561 , n275706 );
not ( n34562 , n25396 );
or ( n34563 , n34561 , n34562 );
buf ( n34564 , n25514 );
not ( n34565 , n34564 );
buf ( n34566 , n25531 );
buf ( n34567 , n25521 );
nand ( n34568 , n34566 , n34567 );
buf ( n34569 , n34568 );
buf ( n34570 , n34569 );
not ( n34571 , n34570 );
or ( n34572 , n34565 , n34571 );
buf ( n34573 , n34569 );
buf ( n34574 , n25514 );
or ( n34575 , n34573 , n34574 );
nand ( n34576 , n34572 , n34575 );
buf ( n34577 , n34576 );
buf ( n34578 , n34577 );
and ( n34579 , n25402 , n34578 );
buf ( n34580 , n25830 );
not ( n34581 , n34580 );
buf ( n34582 , n25847 );
buf ( n34583 , n25837 );
nand ( n34584 , n34582 , n34583 );
buf ( n34585 , n34584 );
buf ( n34586 , n34585 );
not ( n34587 , n34586 );
or ( n34588 , n34581 , n34587 );
buf ( n34589 , n34585 );
buf ( n34590 , n25830 );
or ( n34591 , n34589 , n34590 );
nand ( n34592 , n34588 , n34591 );
buf ( n34593 , n34592 );
buf ( n34594 , n34593 );
not ( n34595 , n34594 );
not ( n34596 , n28761 );
or ( n34597 , n34595 , n34596 );
nand ( n34598 , n275557 , n18324 );
nand ( n34599 , n34597 , n34598 );
nor ( n34600 , n34579 , n34599 );
nand ( n34601 , n34563 , n34600 );
nor ( n34602 , n34560 , n34601 );
buf ( n34603 , n26140 );
not ( n34604 , n34603 );
buf ( n34605 , n26157 );
buf ( n34606 , n26147 );
nand ( n34607 , n34605 , n34606 );
buf ( n34608 , n34607 );
buf ( n34609 , n34608 );
not ( n34610 , n34609 );
or ( n34611 , n34604 , n34610 );
buf ( n34612 , n34608 );
buf ( n34613 , n26140 );
or ( n34614 , n34612 , n34613 );
nand ( n34615 , n34611 , n34614 );
buf ( n34616 , n34615 );
buf ( n34617 , n34616 );
nand ( n34618 , n26027 , n34617 );
nand ( n34619 , n34543 , n34602 , n34618 );
buf ( n34620 , n34619 );
buf ( n34621 , n34620 );
buf ( n34622 , n275554 );
buf ( n34623 , n14614 );
and ( n34624 , n13373 , n34623 );
not ( n34625 , n13373 );
not ( n34626 , n32137 );
buf ( n34627 , n32144 );
not ( n34628 , n34627 );
or ( n34629 , n34626 , n34628 );
or ( n34630 , n34627 , n32137 );
nand ( n34631 , n34629 , n34630 );
buf ( n34632 , n34631 );
and ( n34633 , n34625 , n34632 );
nor ( n34634 , n34624 , n34633 );
not ( n34635 , n34634 );
not ( n34636 , n20846 );
and ( n34637 , n34635 , n34636 );
nand ( n34638 , n16849 , n16873 );
not ( n34639 , n34638 );
not ( n34640 , n32944 );
not ( n34641 , n32943 );
or ( n34642 , n34640 , n34641 );
nand ( n34643 , n34642 , n32945 );
not ( n34644 , n34643 );
or ( n34645 , n34639 , n34644 );
or ( n34646 , n34643 , n34638 );
nand ( n34647 , n34645 , n34646 );
buf ( n34648 , n34647 );
nand ( n34649 , n34648 , n20889 );
not ( n34650 , n32951 );
not ( n34651 , n32950 );
or ( n34652 , n34650 , n34651 );
nand ( n34653 , n34652 , n32952 );
nand ( n34654 , n17266 , n17324 );
xnor ( n34655 , n34653 , n34654 );
buf ( n34656 , n34655 );
nand ( n34657 , n34656 , n20926 );
not ( n34658 , n17414 );
nor ( n34659 , n24714 , n32960 );
not ( n34660 , n34659 );
or ( n34661 , n34658 , n34660 );
or ( n34662 , n34659 , n17414 );
nand ( n34663 , n34661 , n34662 );
buf ( n34664 , n34663 );
and ( n34665 , n34664 , n17409 );
buf ( n34666 , n17413 );
buf ( n34667 , n34666 );
buf ( n34668 , n34667 );
and ( n34669 , n20940 , n34668 );
nor ( n34670 , n34665 , n34669 );
nand ( n34671 , n34649 , n34657 , n34670 );
nor ( n34672 , n34637 , n34671 );
not ( n34673 , n21696 );
not ( n34674 , n34673 );
or ( n34675 , n34672 , n34674 );
nand ( n34676 , n27647 , n13674 );
nand ( n34677 , n34675 , n34676 );
buf ( n34678 , n34677 );
buf ( n34679 , n34678 );
not ( n34680 , n13562 );
not ( n34681 , n20950 );
or ( n34682 , n34680 , n34681 );
and ( n34683 , n20711 , n14564 );
not ( n34684 , n20711 );
not ( n34685 , n21647 );
nor ( n34686 , n21649 , n34685 );
buf ( n34687 , n14526 );
nand ( n34688 , n34686 , n34687 );
not ( n34689 , n32141 );
and ( n34690 , n34688 , n34689 );
not ( n34691 , n34688 );
and ( n34692 , n34691 , n32141 );
nor ( n34693 , n34690 , n34692 );
buf ( n34694 , n34693 );
and ( n34695 , n34684 , n34694 );
nor ( n34696 , n34683 , n34695 );
not ( n34697 , n34696 );
not ( n34698 , n23789 );
and ( n34699 , n34697 , n34698 );
not ( n34700 , n20889 );
not ( n34701 , n20858 );
nand ( n34702 , n34701 , n16803 );
not ( n34703 , n20863 );
nand ( n34704 , n34703 , n20856 );
xnor ( n34705 , n34702 , n34704 );
buf ( n34706 , n34705 );
not ( n34707 , n34706 );
or ( n34708 , n34700 , n34707 );
not ( n34709 , n20901 );
nand ( n34710 , n34709 , n17314 );
not ( n34711 , n34710 );
nand ( n34712 , n17252 , n20903 );
not ( n34713 , n34712 );
or ( n34714 , n34711 , n34713 );
or ( n34715 , n34712 , n34710 );
nand ( n34716 , n34714 , n34715 );
buf ( n34717 , n34716 );
and ( n34718 , n34717 , n20926 );
buf ( n34719 , n17427 );
buf ( n34720 , n34719 );
not ( n34721 , n34720 );
buf ( n34722 , n34721 );
not ( n34723 , n34722 );
not ( n34724 , n34723 );
not ( n34725 , n17499 );
or ( n34726 , n34724 , n34725 );
not ( n34727 , n17428 );
not ( n34728 , n17426 );
and ( n34729 , n17431 , n34728 );
not ( n34730 , n34729 );
or ( n34731 , n34727 , n34730 );
or ( n34732 , n34729 , n17428 );
nand ( n34733 , n34731 , n34732 );
buf ( n34734 , n34733 );
nand ( n34735 , n34734 , n17409 );
nand ( n34736 , n34726 , n34735 );
nor ( n34737 , n34718 , n34736 );
nand ( n34738 , n34708 , n34737 );
nor ( n34739 , n34699 , n34738 );
or ( n34740 , n34739 , n20950 );
nand ( n34741 , n34682 , n34740 );
buf ( n34742 , n34741 );
buf ( n34743 , n34742 );
not ( n34744 , n275550 );
buf ( n34745 , n34744 );
buf ( n34746 , n34745 );
or ( n34747 , n31013 , n27640 );
nand ( n34748 , n27640 , n10996 );
nand ( n34749 , n34747 , n34748 );
buf ( n34750 , n34749 );
buf ( n34751 , n34750 );
not ( n34752 , n275550 );
buf ( n34753 , n34752 );
buf ( n34754 , n34753 );
buf ( n34755 , n275554 );
not ( n34756 , n34302 );
buf ( n34757 , n33442 );
buf ( n34758 , n33391 );
or ( n34759 , n34757 , n34758 );
buf ( n34760 , n34759 );
buf ( n34761 , n34760 );
not ( n34762 , n34761 );
buf ( n34763 , n31804 );
not ( n34764 , n34763 );
buf ( n34765 , n31861 );
nor ( n34766 , n34764 , n34765 );
buf ( n34767 , n34766 );
buf ( n34768 , n34767 );
not ( n34769 , n34768 );
buf ( n34770 , n31838 );
nor ( n34771 , n34769 , n34770 );
buf ( n34772 , n34771 );
buf ( n34773 , n34772 );
not ( n34774 , n34773 );
buf ( n34775 , n27479 );
not ( n34776 , n34775 );
or ( n34777 , n34774 , n34776 );
buf ( n34778 , n34767 );
not ( n34779 , n34778 );
buf ( n34780 , n31922 );
not ( n34781 , n34780 );
or ( n34782 , n34779 , n34781 );
buf ( n34783 , n31804 );
not ( n34784 , n34783 );
buf ( n34785 , n31941 );
not ( n34786 , n34785 );
or ( n34787 , n34784 , n34786 );
buf ( n34788 , n31809 );
nand ( n34789 , n34787 , n34788 );
buf ( n34790 , n34789 );
buf ( n34791 , n34790 );
not ( n34792 , n34791 );
buf ( n34793 , n34792 );
buf ( n34794 , n34793 );
nand ( n34795 , n34782 , n34794 );
buf ( n34796 , n34795 );
buf ( n34797 , n34796 );
not ( n34798 , n34797 );
buf ( n34799 , n34798 );
buf ( n34800 , n34799 );
nand ( n34801 , n34777 , n34800 );
buf ( n34802 , n34801 );
buf ( n34803 , n34802 );
not ( n34804 , n34803 );
or ( n34805 , n34762 , n34804 );
buf ( n34806 , n34802 );
buf ( n34807 , n34760 );
or ( n34808 , n34806 , n34807 );
nand ( n34809 , n34805 , n34808 );
buf ( n34810 , n34809 );
buf ( n34811 , n34810 );
not ( n34812 , n34811 );
or ( n34813 , n34756 , n34812 );
or ( n34814 , n33354 , n33329 );
not ( n34815 , n34814 );
not ( n34816 , n31967 );
nor ( n34817 , n34816 , n31988 );
and ( n34818 , n31978 , n34817 );
not ( n34819 , n34818 );
not ( n34820 , n27260 );
or ( n34821 , n34819 , n34820 );
not ( n34822 , n34817 );
not ( n34823 , n32011 );
or ( n34824 , n34822 , n34823 );
not ( n34825 , n31967 );
not ( n34826 , n32020 );
or ( n34827 , n34825 , n34826 );
nand ( n34828 , n34827 , n31969 );
not ( n34829 , n34828 );
nand ( n34830 , n34824 , n34829 );
not ( n34831 , n34830 );
nand ( n34832 , n34821 , n34831 );
not ( n34833 , n34832 );
or ( n34834 , n34815 , n34833 );
or ( n34835 , n34832 , n34814 );
nand ( n34836 , n34834 , n34835 );
buf ( n34837 , n34836 );
and ( n34838 , n34837 , n28430 );
buf ( n34839 , n32791 );
and ( n34840 , n34839 , n33481 );
not ( n34841 , n34839 );
and ( n34842 , n34841 , n33482 );
or ( n34843 , n34840 , n34842 );
buf ( n34844 , n34843 );
nand ( n34845 , n34844 , n34307 );
nand ( n34846 , n28451 , n277573 );
and ( n34847 , n32755 , n277554 );
not ( n34848 , n28459 );
and ( n34849 , n34848 , n277609 );
and ( n34850 , n34313 , n9360 );
nor ( n34851 , n34847 , n34849 , n34850 );
nand ( n34852 , n34845 , n34846 , n34851 );
nor ( n34853 , n34838 , n34852 );
nand ( n34854 , n34813 , n34853 );
buf ( n34855 , n34854 );
buf ( n34856 , n34855 );
and ( n34857 , n20711 , n34092 );
not ( n34858 , n20711 );
buf ( n34859 , n14132 );
not ( n34860 , n34859 );
nand ( n34861 , n26428 , n26430 );
buf ( n34862 , n34861 );
not ( n34863 , n34862 );
or ( n34864 , n34860 , n34863 );
or ( n34865 , n34862 , n34859 );
nand ( n34866 , n34864 , n34865 );
buf ( n34867 , n34866 );
and ( n34868 , n34858 , n34867 );
nor ( n34869 , n34857 , n34868 );
or ( n34870 , n34869 , n26364 );
not ( n34871 , n16618 );
not ( n34872 , n16879 );
nand ( n34873 , n34871 , n34872 );
not ( n34874 , n34873 );
not ( n34875 , n16668 );
nor ( n34876 , n34875 , n26445 );
not ( n34877 , n34876 );
not ( n34878 , n20875 );
or ( n34879 , n34877 , n34878 );
not ( n34880 , n16891 );
and ( n34881 , n16905 , n34880 );
nand ( n34882 , n34879 , n34881 );
not ( n34883 , n34882 );
or ( n34884 , n34874 , n34883 );
or ( n34885 , n34882 , n34873 );
nand ( n34886 , n34884 , n34885 );
buf ( n34887 , n34886 );
nand ( n34888 , n34887 , n26370 );
not ( n34889 , n17142 );
nand ( n34890 , n34889 , n17354 );
not ( n34891 , n34890 );
not ( n34892 , n17121 );
nor ( n34893 , n17229 , n34892 );
not ( n34894 , n34893 );
not ( n34895 , n20913 );
or ( n34896 , n34894 , n34895 );
not ( n34897 , n26473 );
not ( n34898 , n34892 );
and ( n34899 , n34897 , n34898 );
nor ( n34900 , n34899 , n17352 );
nand ( n34901 , n34896 , n34900 );
not ( n34902 , n34901 );
or ( n34903 , n34891 , n34902 );
or ( n34904 , n34901 , n34890 );
nand ( n34905 , n34903 , n34904 );
buf ( n34906 , n34905 );
nand ( n34907 , n34906 , n26374 );
not ( n34908 , n13525 );
and ( n34909 , n17517 , n34908 );
not ( n34910 , n17517 );
and ( n34911 , n34910 , n13526 );
nor ( n34912 , n34909 , n34911 );
nand ( n34913 , n31180 , n34912 );
not ( n34914 , n17457 );
nor ( n34915 , n17448 , n17454 );
nand ( n34916 , n26487 , n34915 );
nor ( n34917 , n34916 , n20930 );
not ( n34918 , n34917 );
or ( n34919 , n34914 , n34918 );
or ( n34920 , n34917 , n17457 );
nand ( n34921 , n34919 , n34920 );
buf ( n34922 , n34921 );
nand ( n34923 , n34922 , n26393 );
buf ( n34924 , n17456 );
buf ( n34925 , n34924 );
buf ( n34926 , n34925 );
not ( n34927 , n34926 );
not ( n34928 , n34927 );
nand ( n34929 , n26395 , n34928 );
nor ( n34930 , n14830 , n34908 );
not ( n34931 , n34930 );
and ( n34932 , n34923 , n34929 , n34931 );
and ( n34933 , n34888 , n34907 , n34913 , n34932 );
nand ( n34934 , n34870 , n34933 );
buf ( n34935 , n34934 );
buf ( n34936 , n34935 );
not ( n34937 , n275929 );
buf ( n34938 , n34937 );
buf ( n34939 , n34938 );
buf ( n34940 , n275554 );
and ( n34941 , n22335 , n18176 );
not ( n34942 , n22335 );
and ( n34943 , n34942 , n34240 );
or ( n34944 , n34941 , n34943 );
buf ( n34945 , n34944 );
buf ( n34946 , n34945 );
not ( n34947 , n275929 );
buf ( n34948 , n34947 );
buf ( n34949 , n34948 );
and ( n34950 , n23706 , n277621 );
not ( n34951 , n23706 );
not ( n34952 , n29599 );
buf ( n34953 , n31858 );
buf ( n34954 , n31938 );
nand ( n34955 , n34953 , n34954 );
buf ( n34956 , n34955 );
buf ( n34957 , n34956 );
not ( n34958 , n34957 );
buf ( n34959 , n31838 );
buf ( n34960 , n31851 );
not ( n34961 , n34960 );
buf ( n34962 , n34961 );
buf ( n34963 , n34962 );
nor ( n34964 , n34959 , n34963 );
buf ( n34965 , n34964 );
buf ( n34966 , n34965 );
not ( n34967 , n34966 );
buf ( n34968 , n27479 );
not ( n34969 , n34968 );
or ( n34970 , n34967 , n34969 );
buf ( n34971 , n30883 );
buf ( n34972 , n33568 );
buf ( n34973 , n30888 );
and ( n34974 , n34972 , n34973 );
buf ( n34975 , n34974 );
buf ( n34976 , n34975 );
nand ( n34977 , n34971 , n34976 );
buf ( n34978 , n34977 );
buf ( n34979 , n34978 );
buf ( n34980 , n31910 );
nor ( n34981 , n34979 , n34980 );
buf ( n34982 , n34981 );
buf ( n34983 , n34982 );
not ( n34984 , n34983 );
buf ( n34985 , n30872 );
not ( n34986 , n34985 );
or ( n34987 , n34984 , n34986 );
buf ( n34988 , n31895 );
not ( n34989 , n34988 );
buf ( n34990 , n34989 );
buf ( n34991 , n34990 );
buf ( n34992 , n31913 );
buf ( n34993 , n33568 );
and ( n34994 , n34991 , n34992 , n34993 );
buf ( n34995 , n34962 );
nor ( n34996 , n34994 , n34995 );
buf ( n34997 , n34996 );
buf ( n34998 , n34997 );
nand ( n34999 , n34987 , n34998 );
buf ( n35000 , n34999 );
buf ( n35001 , n35000 );
nand ( n35002 , n34970 , n35001 );
buf ( n35003 , n35002 );
buf ( n35004 , n35003 );
not ( n35005 , n35004 );
or ( n35006 , n34958 , n35005 );
buf ( n35007 , n35003 );
buf ( n35008 , n34956 );
or ( n35009 , n35007 , n35008 );
nand ( n35010 , n35006 , n35009 );
buf ( n35011 , n35010 );
buf ( n35012 , n35011 );
not ( n35013 , n35012 );
or ( n35014 , n34952 , n35013 );
nand ( n35015 , n31987 , n32019 );
not ( n35016 , n35015 );
nor ( n35017 , n31979 , n33599 );
not ( n35018 , n35017 );
not ( n35019 , n27260 );
or ( n35020 , n35018 , n35019 );
not ( n35021 , n32015 );
and ( n35022 , n35021 , n30953 );
nand ( n35023 , n30951 , n35022 );
nor ( n35024 , n35023 , n32007 );
not ( n35025 , n35024 );
not ( n35026 , n30946 );
or ( n35027 , n35025 , n35026 );
not ( n35028 , n31999 );
and ( n35029 , n32008 , n35028 , n35021 );
nor ( n35030 , n35029 , n33599 );
nand ( n35031 , n35027 , n35030 );
nand ( n35032 , n35020 , n35031 );
not ( n35033 , n35032 );
or ( n35034 , n35016 , n35033 );
or ( n35035 , n35032 , n35015 );
nand ( n35036 , n35034 , n35035 );
buf ( n35037 , n35036 );
and ( n35038 , n35037 , n23655 );
not ( n35039 , n23673 );
buf ( n35040 , n32802 );
or ( n35041 , n35040 , n32797 );
nand ( n35042 , n35040 , n32797 );
nand ( n35043 , n35041 , n35042 );
buf ( n35044 , n35043 );
not ( n35045 , n35044 );
or ( n35046 , n35039 , n35045 );
and ( n35047 , n27520 , n12198 );
and ( n35048 , n22013 , n12365 );
nor ( n35049 , n35047 , n35048 );
nand ( n35050 , n35046 , n35049 );
nor ( n35051 , n35038 , n35050 );
nand ( n35052 , n35014 , n35051 );
and ( n35053 , n34951 , n35052 );
or ( n35054 , n34950 , n35053 );
buf ( n35055 , n35054 );
buf ( n35056 , n35055 );
nand ( n35057 , n33473 , n29599 );
nand ( n35058 , n33370 , n30962 );
not ( n35059 , n33492 );
not ( n35060 , n23673 );
not ( n35061 , n35060 );
and ( n35062 , n35059 , n35061 );
not ( n35063 , n277453 );
not ( n35064 , n29768 );
or ( n35065 , n35063 , n35064 );
or ( n35066 , n32722 , n12160 );
nand ( n35067 , n35065 , n35066 );
nor ( n35068 , n35062 , n35067 );
and ( n35069 , n35057 , n35058 , n35068 );
or ( n35070 , n35069 , n22193 );
buf ( n35071 , n22192 );
buf ( n35072 , n35071 );
not ( n35073 , n277420 );
or ( n35074 , n35072 , n35073 );
nand ( n35075 , n35070 , n35074 );
buf ( n35076 , n35075 );
buf ( n35077 , n35076 );
not ( n35078 , n275925 );
buf ( n35079 , n35078 );
buf ( n35080 , n35079 );
not ( n35081 , n275929 );
buf ( n35082 , n35081 );
buf ( n35083 , n35082 );
not ( n35084 , n275550 );
buf ( n35085 , n35084 );
buf ( n35086 , n35085 );
buf ( n35087 , n275554 );
not ( n35088 , n275550 );
buf ( n35089 , n35088 );
buf ( n35090 , n35089 );
not ( n35091 , n275550 );
buf ( n35092 , n35091 );
buf ( n35093 , n35092 );
buf ( n35094 , n275554 );
nand ( n35095 , n30448 , n28408 );
nand ( n35096 , n30472 , n32751 );
nand ( n35097 , n30488 , n29163 );
nand ( n35098 , n28451 , n11283 );
and ( n35099 , n28455 , n12207 );
or ( n35100 , n28459 , n30491 );
nand ( n35101 , n20649 , n9300 );
nand ( n35102 , n35100 , n35101 );
nor ( n35103 , n35099 , n35102 );
and ( n35104 , n35097 , n35098 , n35103 );
nand ( n35105 , n35095 , n35096 , n35104 );
buf ( n35106 , n35105 );
buf ( n35107 , n35106 );
buf ( n35108 , n23080 );
and ( n35109 , n14830 , n35108 );
not ( n35110 , n14830 );
and ( n35111 , n35110 , n16285 );
or ( n35112 , n35109 , n35111 );
buf ( n35113 , n35112 );
buf ( n35114 , n35113 );
not ( n35115 , n275925 );
buf ( n35116 , n35115 );
buf ( n35117 , n35116 );
not ( n35118 , n275929 );
buf ( n35119 , n35118 );
buf ( n35120 , n35119 );
buf ( n35121 , n19580 );
and ( n35122 , n22799 , n35121 );
not ( n35123 , n22799 );
not ( n35124 , n19563 );
not ( n35125 , n35124 );
not ( n35126 , n24389 );
nor ( n35127 , n24393 , n35126 );
not ( n35128 , n35127 );
or ( n35129 , n35125 , n35128 );
or ( n35130 , n35127 , n35124 );
nand ( n35131 , n35129 , n35130 );
buf ( n35132 , n35131 );
and ( n35133 , n35123 , n35132 );
nor ( n35134 , n35122 , n35133 );
or ( n35135 , n35134 , n19216 );
not ( n35136 , n19360 );
nand ( n35137 , n20463 , n20490 );
not ( n35138 , n35137 );
not ( n35139 , n20486 );
nand ( n35140 , n35139 , n24267 );
not ( n35141 , n35140 );
or ( n35142 , n35138 , n35141 );
or ( n35143 , n35140 , n35137 );
nand ( n35144 , n35142 , n35143 );
buf ( n35145 , n35144 );
not ( n35146 , n35145 );
or ( n35147 , n35136 , n35146 );
nand ( n35148 , n19387 , n18908 );
nand ( n35149 , n35147 , n35148 );
not ( n35150 , n19353 );
not ( n35151 , n35150 );
nand ( n35152 , n22845 , n20257 );
not ( n35153 , n35152 );
not ( n35154 , n22844 );
not ( n35155 , n33999 );
nor ( n35156 , n35154 , n35155 );
not ( n35157 , n35156 );
not ( n35158 , n24187 );
or ( n35159 , n35157 , n35158 );
not ( n35160 , n20200 );
nand ( n35161 , n35159 , n35160 );
not ( n35162 , n35161 );
or ( n35163 , n35153 , n35162 );
or ( n35164 , n35161 , n35152 );
nand ( n35165 , n35163 , n35164 );
buf ( n35166 , n35165 );
not ( n35167 , n35166 );
or ( n35168 , n35151 , n35167 );
not ( n35169 , n18899 );
not ( n35170 , n19654 );
or ( n35171 , n35169 , n35170 );
or ( n35172 , n19654 , n18899 );
nand ( n35173 , n35171 , n35172 );
not ( n35174 , n35173 );
not ( n35175 , n19318 );
or ( n35176 , n35174 , n35175 );
not ( n35177 , n20525 );
not ( n35178 , n24312 );
or ( n35179 , n35177 , n35178 );
or ( n35180 , n24312 , n20525 );
nand ( n35181 , n35179 , n35180 );
buf ( n35182 , n35181 );
not ( n35183 , n35182 );
or ( n35184 , n19291 , n35183 );
nand ( n35185 , n35176 , n35184 );
not ( n35186 , n20523 );
buf ( n35187 , n35186 );
buf ( n35188 , n35187 );
not ( n35189 , n35188 );
nor ( n35190 , n32248 , n35189 );
nor ( n35191 , n35185 , n35190 );
nand ( n35192 , n35168 , n35191 );
nor ( n35193 , n35149 , n35192 );
nand ( n35194 , n35135 , n35193 );
buf ( n35195 , n35194 );
buf ( n35196 , n35195 );
buf ( n35197 , n275554 );
buf ( n35198 , n275554 );
not ( n35199 , n33723 );
and ( n35200 , n35199 , n27845 );
not ( n35201 , n21001 );
not ( n35202 , n33773 );
or ( n35203 , n35201 , n35202 );
and ( n35204 , n33737 , n19358 );
not ( n35205 , n27932 );
not ( n35206 , n19219 );
or ( n35207 , n35205 , n35206 );
nand ( n35208 , n33754 , n19290 );
nand ( n35209 , n35207 , n35208 );
nor ( n35210 , n35204 , n35209 );
nand ( n35211 , n35203 , n35210 );
nor ( n35212 , n35200 , n35211 );
or ( n35213 , n35212 , n21030 );
nand ( n35214 , n21030 , n18804 );
nand ( n35215 , n35213 , n35214 );
buf ( n35216 , n35215 );
buf ( n35217 , n35216 );
not ( n35218 , n275550 );
buf ( n35219 , n35218 );
buf ( n35220 , n35219 );
buf ( n35221 , n275554 );
buf ( n35222 , n275554 );
or ( n35223 , n27112 , n20743 );
nand ( n35224 , n27131 , n16968 );
nand ( n35225 , n27149 , n17405 );
nand ( n35226 , n17411 , n27157 );
nand ( n35227 , n20785 , n27161 );
nand ( n35228 , n17562 , n13446 );
and ( n35229 , n17513 , n13458 );
not ( n35230 , n17513 );
and ( n35231 , n35230 , n33635 );
nor ( n35232 , n35229 , n35231 );
nand ( n35233 , n17545 , n35232 );
and ( n35234 , n35226 , n35227 , n35228 , n35233 );
and ( n35235 , n35224 , n35225 , n35234 );
nand ( n35236 , n35223 , n35235 );
buf ( n35237 , n35236 );
buf ( n35238 , n35237 );
not ( n35239 , n275925 );
buf ( n35240 , n35239 );
buf ( n35241 , n35240 );
not ( n35242 , n275550 );
buf ( n35243 , n35242 );
buf ( n35244 , n35243 );
buf ( n35245 , n275554 );
not ( n35246 , n275929 );
buf ( n35247 , n35246 );
buf ( n35248 , n35247 );
not ( n35249 , n275929 );
buf ( n35250 , n35249 );
buf ( n35251 , n35250 );
nand ( n35252 , n25064 , n25267 );
buf ( n35253 , n25273 );
not ( n35254 , n35253 );
buf ( n35255 , n25354 );
nand ( n35256 , n35254 , n35255 );
buf ( n35257 , n35256 );
buf ( n35258 , n35257 );
not ( n35259 , n35258 );
buf ( n35260 , n25340 );
not ( n35261 , n35260 );
buf ( n35262 , n35261 );
buf ( n35263 , n35262 );
buf ( n35264 , n25282 );
or ( n35265 , n35263 , n35264 );
buf ( n35266 , n25282 );
not ( n35267 , n35266 );
buf ( n35268 , n25131 );
buf ( n35269 , n25264 );
nand ( n35270 , n35267 , n35268 , n35269 );
buf ( n35271 , n35270 );
buf ( n35272 , n35271 );
buf ( n35273 , n25348 );
nand ( n35274 , n35265 , n35272 , n35273 );
buf ( n35275 , n35274 );
buf ( n35276 , n35275 );
not ( n35277 , n35276 );
or ( n35278 , n35259 , n35277 );
buf ( n35279 , n35275 );
buf ( n35280 , n35257 );
or ( n35281 , n35279 , n35280 );
nand ( n35282 , n35278 , n35281 );
buf ( n35283 , n35282 );
buf ( n35284 , n35283 );
not ( n35285 , n35284 );
nor ( n35286 , n35285 , n25389 );
nand ( n35287 , n25397 , n275868 );
buf ( n35288 , n25595 );
not ( n35289 , n35288 );
buf ( n35290 , n25680 );
nand ( n35291 , n35289 , n35290 );
buf ( n35292 , n35291 );
buf ( n35293 , n35292 );
not ( n35294 , n35293 );
buf ( n35295 , n25666 );
not ( n35296 , n35295 );
buf ( n35297 , n35296 );
buf ( n35298 , n35297 );
buf ( n35299 , n25603 );
or ( n35300 , n35298 , n35299 );
buf ( n35301 , n25603 );
not ( n35302 , n35301 );
buf ( n35303 , n25456 );
buf ( n35304 , n25586 );
nand ( n35305 , n35302 , n35303 , n35304 );
buf ( n35306 , n35305 );
buf ( n35307 , n35306 );
buf ( n35308 , n25674 );
nand ( n35309 , n35300 , n35307 , n35308 );
buf ( n35310 , n35309 );
buf ( n35311 , n35310 );
not ( n35312 , n35311 );
or ( n35313 , n35294 , n35312 );
buf ( n35314 , n35310 );
buf ( n35315 , n35292 );
or ( n35316 , n35314 , n35315 );
nand ( n35317 , n35313 , n35316 );
buf ( n35318 , n35317 );
buf ( n35319 , n35318 );
and ( n35320 , n25402 , n35319 );
nor ( n35321 , n19639 , n29539 );
nor ( n35322 , n35320 , n35321 );
buf ( n35323 , n25910 );
not ( n35324 , n35323 );
buf ( n35325 , n25991 );
nand ( n35326 , n35324 , n35325 );
buf ( n35327 , n35326 );
buf ( n35328 , n35327 );
not ( n35329 , n35328 );
buf ( n35330 , n25977 );
not ( n35331 , n35330 );
buf ( n35332 , n35331 );
buf ( n35333 , n35332 );
buf ( n35334 , n25917 );
or ( n35335 , n35333 , n35334 );
buf ( n35336 , n25917 );
not ( n35337 , n35336 );
buf ( n35338 , n25773 );
buf ( n35339 , n25902 );
nand ( n35340 , n35337 , n35338 , n35339 );
buf ( n35341 , n35340 );
buf ( n35342 , n35341 );
buf ( n35343 , n25985 );
nand ( n35344 , n35335 , n35342 , n35343 );
buf ( n35345 , n35344 );
buf ( n35346 , n35345 );
not ( n35347 , n35346 );
or ( n35348 , n35329 , n35347 );
buf ( n35349 , n35345 );
buf ( n35350 , n35327 );
or ( n35351 , n35349 , n35350 );
nand ( n35352 , n35348 , n35351 );
buf ( n35353 , n35352 );
buf ( n35354 , n35353 );
nand ( n35355 , n25717 , n35354 );
nand ( n35356 , n35287 , n35322 , n35355 );
nor ( n35357 , n35286 , n35356 );
buf ( n35358 , n26219 );
not ( n35359 , n35358 );
buf ( n35360 , n26295 );
nand ( n35361 , n35359 , n35360 );
buf ( n35362 , n35361 );
buf ( n35363 , n35362 );
not ( n35364 , n35363 );
buf ( n35365 , n26281 );
not ( n35366 , n35365 );
buf ( n35367 , n35366 );
buf ( n35368 , n35367 );
buf ( n35369 , n26226 );
or ( n35370 , n35368 , n35369 );
buf ( n35371 , n26226 );
not ( n35372 , n35371 );
buf ( n35373 , n26081 );
buf ( n35374 , n26212 );
nand ( n35375 , n35372 , n35373 , n35374 );
buf ( n35376 , n35375 );
buf ( n35377 , n35376 );
buf ( n35378 , n26289 );
nand ( n35379 , n35370 , n35377 , n35378 );
buf ( n35380 , n35379 );
buf ( n35381 , n35380 );
not ( n35382 , n35381 );
or ( n35383 , n35364 , n35382 );
buf ( n35384 , n35380 );
buf ( n35385 , n35362 );
or ( n35386 , n35384 , n35385 );
nand ( n35387 , n35383 , n35386 );
buf ( n35388 , n35387 );
buf ( n35389 , n35388 );
nand ( n35390 , n26027 , n35389 );
nand ( n35391 , n35252 , n35357 , n35390 );
buf ( n35392 , n35391 );
buf ( n35393 , n35392 );
not ( n35394 , n24386 );
or ( n35395 , n35394 , n21774 );
nand ( n35396 , n21770 , n9492 );
nand ( n35397 , n35395 , n35396 );
buf ( n35398 , n35397 );
buf ( n35399 , n35398 );
and ( n35400 , n26516 , n27832 );
not ( n35401 , n26516 );
not ( n35402 , n27835 );
nand ( n35403 , n35402 , n27812 );
buf ( n35404 , n29824 );
not ( n35405 , n35404 );
and ( n35406 , n35403 , n35405 );
not ( n35407 , n35403 );
and ( n35408 , n35407 , n35404 );
nor ( n35409 , n35406 , n35408 );
buf ( n35410 , n35409 );
and ( n35411 , n35401 , n35410 );
nor ( n35412 , n35400 , n35411 );
not ( n35413 , n35412 );
and ( n35414 , n35413 , n26638 );
not ( n35415 , n21001 );
nand ( n35416 , n30035 , n30057 );
not ( n35417 , n35416 );
nor ( n35418 , n28014 , n30038 );
not ( n35419 , n35418 );
not ( n35420 , n30043 );
or ( n35421 , n35419 , n35420 );
not ( n35422 , n28037 );
not ( n35423 , n30038 );
and ( n35424 , n35422 , n35423 );
nor ( n35425 , n35424 , n30052 );
nand ( n35426 , n35421 , n35425 );
not ( n35427 , n35426 );
or ( n35428 , n35417 , n35427 );
or ( n35429 , n35426 , n35416 );
nand ( n35430 , n35428 , n35429 );
buf ( n35431 , n35430 );
not ( n35432 , n35431 );
or ( n35433 , n35415 , n35432 );
not ( n35434 , n30099 );
nand ( n35435 , n35434 , n30117 );
not ( n35436 , n35435 );
not ( n35437 , n30101 );
nor ( n35438 , n28079 , n35437 );
not ( n35439 , n35438 );
not ( n35440 , n28092 );
or ( n35441 , n35439 , n35440 );
not ( n35442 , n30101 );
not ( n35443 , n28109 );
or ( n35444 , n35442 , n35443 );
not ( n35445 , n30113 );
nand ( n35446 , n35444 , n35445 );
not ( n35447 , n35446 );
nand ( n35448 , n35441 , n35447 );
not ( n35449 , n35448 );
or ( n35450 , n35436 , n35449 );
or ( n35451 , n35448 , n35435 );
nand ( n35452 , n35450 , n35451 );
buf ( n35453 , n35452 );
and ( n35454 , n35453 , n19358 );
not ( n35455 , n30019 );
not ( n35456 , n27619 );
or ( n35457 , n35455 , n35456 );
not ( n35458 , n30162 );
not ( n35459 , n27072 );
nor ( n35460 , n28122 , n28130 );
nand ( n35461 , n28127 , n35459 , n35460 , n28128 );
nor ( n35462 , n33111 , n35461 );
not ( n35463 , n35462 );
or ( n35464 , n35458 , n35463 );
or ( n35465 , n35462 , n30162 );
nand ( n35466 , n35464 , n35465 );
buf ( n35467 , n35466 );
nand ( n35468 , n35467 , n19290 );
nand ( n35469 , n35457 , n35468 );
nor ( n35470 , n35454 , n35469 );
nand ( n35471 , n35433 , n35470 );
nor ( n35472 , n35414 , n35471 );
not ( n35473 , n33546 );
or ( n35474 , n35472 , n35473 );
nand ( n35475 , n28146 , n18484 );
nand ( n35476 , n35474 , n35475 );
buf ( n35477 , n35476 );
buf ( n35478 , n35477 );
not ( n35479 , n275550 );
buf ( n35480 , n35479 );
buf ( n35481 , n35480 );
buf ( n35482 , n275554 );
not ( n35483 , n275929 );
buf ( n35484 , n35483 );
buf ( n35485 , n35484 );
not ( n35486 , n16237 );
or ( n35487 , n35486 , n23807 );
buf ( n35488 , n23060 );
nand ( n35489 , n35488 , n23807 );
nand ( n35490 , n35487 , n35489 );
buf ( n35491 , n35490 );
buf ( n35492 , n35491 );
buf ( n35493 , n275554 );
not ( n35494 , n275929 );
buf ( n35495 , n35494 );
buf ( n35496 , n35495 );
not ( n35497 , n275929 );
buf ( n35498 , n35497 );
buf ( n35499 , n35498 );
not ( n35500 , n275550 );
buf ( n35501 , n35500 );
buf ( n35502 , n35501 );
not ( n35503 , n275925 );
buf ( n35504 , n35503 );
buf ( n35505 , n35504 );
not ( n35506 , n275925 );
buf ( n35507 , n35506 );
buf ( n35508 , n35507 );
not ( n35509 , n275925 );
buf ( n35510 , n35509 );
buf ( n35511 , n35510 );
buf ( n35512 , n275554 );
not ( n35513 , n275925 );
buf ( n35514 , n35513 );
buf ( n35515 , n35514 );
or ( n35516 , n33274 , n21030 );
nand ( n35517 , n21030 , n18620 );
nand ( n35518 , n35516 , n35517 );
buf ( n35519 , n35518 );
buf ( n35520 , n35519 );
not ( n35521 , n275929 );
buf ( n35522 , n35521 );
buf ( n35523 , n35522 );
nand ( n35524 , n34359 , n28306 );
nand ( n35525 , n34376 , n28330 );
and ( n35526 , n31449 , n34383 );
and ( n35527 , n28350 , n12205 );
nor ( n35528 , n35526 , n35527 );
and ( n35529 , n28231 , n12351 );
or ( n35530 , n28354 , n11251 );
nand ( n35531 , n28357 , n11246 );
nand ( n35532 , n35530 , n35531 );
nor ( n35533 , n35529 , n35532 );
nand ( n35534 , n35524 , n35525 , n35528 , n35533 );
buf ( n35535 , n35534 );
buf ( n35536 , n35535 );
not ( n35537 , n275550 );
buf ( n35538 , n35537 );
buf ( n35539 , n35538 );
buf ( n35540 , n275554 );
buf ( n35541 , n275554 );
buf ( n35542 , n275554 );
buf ( n35543 , n275554 );
not ( n35544 , n275550 );
buf ( n35545 , n35544 );
buf ( n35546 , n35545 );
not ( n35547 , n275929 );
buf ( n35548 , n35547 );
buf ( n35549 , n35548 );
and ( n35550 , n17547 , n14896 );
and ( n35551 , n22899 , n22902 );
nor ( n35552 , n35550 , n35551 );
not ( n35553 , n35552 );
not ( n35554 , n275721 );
not ( n35555 , n35554 );
and ( n35556 , n35553 , n35555 );
and ( n35557 , n17542 , n14528 );
nor ( n35558 , n35556 , n35557 );
xor ( n35559 , n23010 , n23011 );
xor ( n35560 , n35559 , n23013 );
buf ( n35561 , n35560 );
buf ( n35562 , n35561 );
nand ( n35563 , n22918 , n35562 );
nand ( n35564 , n22914 , n13099 );
xor ( n35565 , n23239 , n23240 );
xor ( n35566 , n35565 , n23242 );
buf ( n35567 , n35566 );
buf ( n35568 , n35567 );
nand ( n35569 , n23152 , n35568 );
nand ( n35570 , n35558 , n35563 , n35564 , n35569 );
buf ( n35571 , n35570 );
buf ( n35572 , n35571 );
not ( n35573 , n275929 );
buf ( n35574 , n35573 );
buf ( n35575 , n35574 );
buf ( n35576 , n275554 );
or ( n35577 , n23931 , n21774 );
nand ( n35578 , n21774 , n9732 );
nand ( n35579 , n35577 , n35578 );
buf ( n35580 , n35579 );
buf ( n35581 , n35580 );
buf ( n35582 , n275554 );
not ( n35583 , n275550 );
buf ( n35584 , n35583 );
buf ( n35585 , n35584 );
buf ( n35586 , n275554 );
and ( n35587 , n31468 , n275769 );
not ( n35588 , n13676 );
nor ( n35589 , n14830 , n35588 );
nor ( n35590 , n35587 , n35589 );
buf ( n35591 , n22967 );
not ( n35592 , n35591 );
buf ( n35593 , n22981 );
nand ( n35594 , n35592 , n35593 );
buf ( n35595 , n35594 );
buf ( n35596 , n35595 );
not ( n35597 , n35596 );
buf ( n35598 , n23043 );
not ( n35599 , n35598 );
buf ( n35600 , n35599 );
buf ( n35601 , n35600 );
buf ( n35602 , n22993 );
or ( n35603 , n35601 , n35602 );
buf ( n35604 , n22975 );
nand ( n35605 , n35603 , n35604 );
buf ( n35606 , n35605 );
buf ( n35607 , n35606 );
not ( n35608 , n35607 );
or ( n35609 , n35597 , n35608 );
buf ( n35610 , n35606 );
buf ( n35611 , n35595 );
or ( n35612 , n35610 , n35611 );
nand ( n35613 , n35609 , n35612 );
buf ( n35614 , n35613 );
buf ( n35615 , n35614 );
nand ( n35616 , n22918 , n35615 );
nand ( n35617 , n22914 , n22961 );
buf ( n35618 , n23198 );
not ( n35619 , n35618 );
buf ( n35620 , n23211 );
nand ( n35621 , n35619 , n35620 );
buf ( n35622 , n35621 );
buf ( n35623 , n35622 );
not ( n35624 , n35623 );
buf ( n35625 , n23272 );
not ( n35626 , n35625 );
buf ( n35627 , n35626 );
buf ( n35628 , n35627 );
buf ( n35629 , n23223 );
or ( n35630 , n35628 , n35629 );
buf ( n35631 , n23205 );
nand ( n35632 , n35630 , n35631 );
buf ( n35633 , n35632 );
buf ( n35634 , n35633 );
not ( n35635 , n35634 );
or ( n35636 , n35624 , n35635 );
buf ( n35637 , n35633 );
buf ( n35638 , n35622 );
or ( n35639 , n35637 , n35638 );
nand ( n35640 , n35636 , n35639 );
buf ( n35641 , n35640 );
buf ( n35642 , n35641 );
nand ( n35643 , n23152 , n35642 );
nand ( n35644 , n35590 , n35616 , n35617 , n35643 );
buf ( n35645 , n35644 );
buf ( n35646 , n35645 );
buf ( n35647 , n275554 );
buf ( n35648 , n275554 );
or ( n35649 , n30256 , n26364 );
nand ( n35650 , n30318 , n26370 );
nand ( n35651 , n30361 , n26374 );
not ( n35652 , n14640 );
and ( n35653 , n33953 , n14714 );
not ( n35654 , n35653 );
or ( n35655 , n35652 , n35654 );
or ( n35656 , n35653 , n14640 );
nand ( n35657 , n35655 , n35656 );
not ( n35658 , n26390 );
and ( n35659 , n35657 , n35658 );
nand ( n35660 , n30374 , n32188 );
nand ( n35661 , n26395 , n24937 );
nand ( n35662 , n17542 , n14641 );
nand ( n35663 , n35660 , n35661 , n35662 );
nor ( n35664 , n35659 , n35663 );
and ( n35665 , n35650 , n35651 , n35664 );
nand ( n35666 , n35649 , n35665 );
buf ( n35667 , n35666 );
buf ( n35668 , n35667 );
not ( n35669 , n275925 );
buf ( n35670 , n35669 );
buf ( n35671 , n35670 );
buf ( n35672 , n275554 );
and ( n35673 , n23907 , n30506 );
not ( n35674 , n23907 );
not ( n35675 , n19478 );
buf ( n35676 , n19605 );
not ( n35677 , n35676 );
or ( n35678 , n35675 , n35677 );
or ( n35679 , n35676 , n19478 );
nand ( n35680 , n35678 , n35679 );
buf ( n35681 , n35680 );
and ( n35682 , n35674 , n35681 );
nor ( n35683 , n35673 , n35682 );
not ( n35684 , n35683 );
and ( n35685 , n35684 , n20987 );
not ( n35686 , n20340 );
nand ( n35687 , n20070 , n35686 );
not ( n35688 , n35687 );
not ( n35689 , n20337 );
or ( n35690 , n35688 , n35689 );
or ( n35691 , n35687 , n20337 );
nand ( n35692 , n35690 , n35691 );
buf ( n35693 , n35692 );
nand ( n35694 , n35693 , n21001 );
nand ( n35695 , n20400 , n20504 );
not ( n35696 , n35695 );
not ( n35697 , n20500 );
or ( n35698 , n35696 , n35697 );
buf ( n35699 , n20500 );
or ( n35700 , n35699 , n35695 );
nand ( n35701 , n35698 , n35700 );
buf ( n35702 , n35701 );
nand ( n35703 , n35702 , n19358 );
not ( n35704 , n20551 );
not ( n35705 , n20547 );
or ( n35706 , n35704 , n35705 );
or ( n35707 , n20547 , n20551 );
nand ( n35708 , n35706 , n35707 );
buf ( n35709 , n35708 );
and ( n35710 , n35709 , n19290 );
buf ( n35711 , n20550 );
buf ( n35712 , n35711 );
buf ( n35713 , n35712 );
buf ( n35714 , n35713 );
and ( n35715 , n19219 , n35714 );
nor ( n35716 , n35710 , n35715 );
nand ( n35717 , n35694 , n35703 , n35716 );
nor ( n35718 , n35685 , n35717 );
or ( n35719 , n35718 , n21030 );
nand ( n35720 , n21030 , n18339 );
nand ( n35721 , n35719 , n35720 );
buf ( n35722 , n35721 );
buf ( n35723 , n35722 );
not ( n35724 , n275929 );
buf ( n35725 , n35724 );
buf ( n35726 , n35725 );
not ( n35727 , n275929 );
buf ( n35728 , n35727 );
buf ( n35729 , n35728 );
buf ( n35730 , n27664 );
buf ( n35731 , n35730 );
or ( n35732 , n23835 , n20743 );
and ( n35733 , n23866 , n17405 );
nand ( n35734 , n17411 , n23881 );
nand ( n35735 , n20785 , n15557 );
nand ( n35736 , n17562 , n13959 );
and ( n35737 , n17532 , n17533 );
not ( n35738 , n17532 );
and ( n35739 , n35738 , n13949 );
nor ( n35740 , n35737 , n35739 );
nand ( n35741 , n35740 , n17545 );
nand ( n35742 , n35734 , n35735 , n35736 , n35741 );
nor ( n35743 , n35733 , n35742 );
nand ( n35744 , n23850 , n16970 );
and ( n35745 , n35743 , n35744 );
nand ( n35746 , n35732 , n35745 );
buf ( n35747 , n35746 );
buf ( n35748 , n35747 );
or ( n35749 , n32366 , n26365 );
nand ( n35750 , n32380 , n26370 );
nand ( n35751 , n32393 , n26374 );
and ( n35752 , n17510 , n13617 );
not ( n35753 , n17510 );
not ( n35754 , n13616 );
and ( n35755 , n35753 , n35754 );
nor ( n35756 , n35752 , n35755 );
nand ( n35757 , n31180 , n35756 );
nand ( n35758 , n32401 , n26393 );
nand ( n35759 , n26395 , n32405 );
nor ( n35760 , n14830 , n35754 );
not ( n35761 , n35760 );
and ( n35762 , n35758 , n35759 , n35761 );
and ( n35763 , n35750 , n35751 , n35757 , n35762 );
nand ( n35764 , n35749 , n35763 );
buf ( n35765 , n35764 );
buf ( n35766 , n35765 );
not ( n35767 , n275805 );
nand ( n35768 , n35767 , n275837 );
not ( n35769 , n35768 );
not ( n35770 , n275767 );
or ( n35771 , n35769 , n35770 );
or ( n35772 , n275767 , n35768 );
nand ( n35773 , n35771 , n35772 );
buf ( n35774 , n35773 );
buf ( n35775 , n35774 );
buf ( n35776 , n275554 );
buf ( n35777 , n275554 );
not ( n35778 , n275925 );
buf ( n35779 , n35778 );
buf ( n35780 , n35779 );
buf ( n35781 , n275554 );
not ( n35782 , n275550 );
buf ( n35783 , n35782 );
buf ( n35784 , n35783 );
not ( n35785 , n275929 );
buf ( n35786 , n35785 );
buf ( n35787 , n35786 );
not ( n35788 , n275550 );
buf ( n35789 , n35788 );
buf ( n35790 , n35789 );
not ( n35791 , n277355 );
or ( n35792 , n35791 , n9158 );
nand ( n35793 , n9369 , n9158 );
nand ( n35794 , n35792 , n35793 );
buf ( n35795 , n35794 );
buf ( n35796 , n35795 );
not ( n35797 , n275550 );
buf ( n35798 , n35797 );
buf ( n35799 , n35798 );
buf ( n35800 , n19496 );
not ( n35801 , n35800 );
not ( n35802 , n35801 );
and ( n35803 , n21039 , n35802 );
not ( n35804 , n21039 );
not ( n35805 , n19621 );
not ( n35806 , n19605 );
nand ( n35807 , n35806 , n19478 );
not ( n35808 , n35807 );
or ( n35809 , n35805 , n35808 );
or ( n35810 , n35807 , n19621 );
nand ( n35811 , n35809 , n35810 );
buf ( n35812 , n35811 );
and ( n35813 , n35804 , n35812 );
nor ( n35814 , n35803 , n35813 );
or ( n35815 , n35814 , n19216 );
nand ( n35816 , n20387 , n20506 );
not ( n35817 , n35816 );
not ( n35818 , n20400 );
not ( n35819 , n20500 );
or ( n35820 , n35818 , n35819 );
nand ( n35821 , n35820 , n20504 );
not ( n35822 , n35821 );
or ( n35823 , n35817 , n35822 );
or ( n35824 , n35821 , n35816 );
nand ( n35825 , n35823 , n35824 );
buf ( n35826 , n35825 );
and ( n35827 , n35826 , n19360 );
not ( n35828 , n19317 );
and ( n35829 , n19658 , n18408 );
not ( n35830 , n19658 );
and ( n35831 , n35830 , n19659 );
nor ( n35832 , n35829 , n35831 );
not ( n35833 , n35832 );
and ( n35834 , n35828 , n35833 );
buf ( n35835 , n20548 );
buf ( n35836 , n35835 );
buf ( n35837 , n35836 );
and ( n35838 , n33162 , n35837 );
nor ( n35839 , n35834 , n35838 );
not ( n35840 , n21600 );
not ( n35841 , n20551 );
nand ( n35842 , n35841 , n20547 );
not ( n35843 , n35842 );
or ( n35844 , n35840 , n35843 );
or ( n35845 , n35842 , n21600 );
nand ( n35846 , n35844 , n35845 );
buf ( n35847 , n35846 );
nand ( n35848 , n35847 , n29075 );
nand ( n35849 , n19387 , n18402 );
nand ( n35850 , n35839 , n35848 , n35849 );
nor ( n35851 , n35827 , n35850 );
nand ( n35852 , n19983 , n20344 );
not ( n35853 , n35852 );
not ( n35854 , n20070 );
not ( n35855 , n20337 );
or ( n35856 , n35854 , n35855 );
nand ( n35857 , n35856 , n35686 );
not ( n35858 , n35857 );
or ( n35859 , n35853 , n35858 );
or ( n35860 , n35857 , n35852 );
nand ( n35861 , n35859 , n35860 );
buf ( n35862 , n35861 );
not ( n35863 , n19353 );
nand ( n35864 , n35862 , n35863 );
and ( n35865 , n35851 , n35864 );
nand ( n35866 , n35815 , n35865 );
buf ( n35867 , n35866 );
buf ( n35868 , n35867 );
not ( n35869 , n275550 );
buf ( n35870 , n35869 );
buf ( n35871 , n35870 );
buf ( n35872 , n275554 );
not ( n35873 , n20846 );
and ( n35874 , n32271 , n35873 );
not ( n35875 , n20889 );
not ( n35876 , n32290 );
or ( n35877 , n35875 , n35876 );
and ( n35878 , n32309 , n20927 );
not ( n35879 , n17409 );
not ( n35880 , n32323 );
or ( n35881 , n35879 , n35880 );
nand ( n35882 , n20940 , n32327 );
nand ( n35883 , n35881 , n35882 );
nor ( n35884 , n35878 , n35883 );
nand ( n35885 , n35877 , n35884 );
nor ( n35886 , n35874 , n35885 );
or ( n35887 , n35886 , n21697 );
nand ( n35888 , n21696 , n13888 );
nand ( n35889 , n35887 , n35888 );
buf ( n35890 , n35889 );
buf ( n35891 , n35890 );
not ( n35892 , n275929 );
buf ( n35893 , n35892 );
buf ( n35894 , n35893 );
not ( n35895 , n275925 );
buf ( n35896 , n35895 );
buf ( n35897 , n35896 );
buf ( n35898 , n275554 );
nand ( n35899 , n34055 , n28408 );
not ( n35900 , n28429 );
nand ( n35901 , n34063 , n35900 );
and ( n35902 , n34073 , n29163 );
nor ( n35903 , n29172 , n12136 );
not ( n35904 , n12271 );
or ( n35905 , n28459 , n35904 );
nand ( n35906 , n20649 , n9306 );
nand ( n35907 , n35905 , n35906 );
nor ( n35908 , n35902 , n35903 , n35907 );
not ( n35909 , n28450 );
nand ( n35910 , n35909 , n11607 );
nand ( n35911 , n35899 , n35901 , n35908 , n35910 );
buf ( n35912 , n35911 );
buf ( n35913 , n35912 );
or ( n35914 , n35801 , n21774 );
nand ( n35915 , n21770 , n9517 );
nand ( n35916 , n35914 , n35915 );
buf ( n35917 , n35916 );
buf ( n35918 , n35917 );
not ( n35919 , n275929 );
buf ( n35920 , n35919 );
buf ( n35921 , n35920 );
buf ( n35922 , n275554 );
or ( n35923 , n22816 , n19216 );
nand ( n35924 , n22836 , n19360 );
nand ( n35925 , n22858 , n19354 );
not ( n35926 , n34284 );
not ( n35927 , n19318 );
or ( n35928 , n35926 , n35927 );
or ( n35929 , n19291 , n22865 );
nand ( n35930 , n35928 , n35929 );
nor ( n35931 , n32248 , n22872 );
not ( n35932 , n18878 );
nor ( n35933 , n35932 , n19388 );
nor ( n35934 , n35930 , n35931 , n35933 );
and ( n35935 , n35924 , n35925 , n35934 );
nand ( n35936 , n35923 , n35935 );
buf ( n35937 , n35936 );
buf ( n35938 , n35937 );
or ( n35939 , n35472 , n21030 );
nand ( n35940 , n21030 , n18474 );
nand ( n35941 , n35939 , n35940 );
buf ( n35942 , n35941 );
buf ( n35943 , n35942 );
or ( n35944 , n29410 , n19216 );
and ( n35945 , n29444 , n19360 );
not ( n35946 , n19317 );
and ( n35947 , n29474 , n19020 );
not ( n35948 , n29474 );
and ( n35949 , n35948 , n29475 );
nor ( n35950 , n35947 , n35949 );
not ( n35951 , n35950 );
and ( n35952 , n35946 , n35951 );
and ( n35953 , n33162 , n29459 );
nor ( n35954 , n35952 , n35953 );
nand ( n35955 , n29454 , n29075 );
nand ( n35956 , n33840 , n19010 );
nand ( n35957 , n35954 , n35955 , n35956 );
nor ( n35958 , n35945 , n35957 );
nand ( n35959 , n29427 , n33157 );
and ( n35960 , n35958 , n35959 );
nand ( n35961 , n35944 , n35960 );
buf ( n35962 , n35961 );
buf ( n35963 , n35962 );
buf ( n35964 , n21161 );
not ( n35965 , n35964 );
or ( n35966 , n35965 , n21774 );
nand ( n35967 , n21774 , n9562 );
nand ( n35968 , n35966 , n35967 );
buf ( n35969 , n35968 );
buf ( n35970 , n35969 );
not ( n35971 , n275550 );
buf ( n35972 , n35971 );
buf ( n35973 , n35972 );
or ( n35974 , n32228 , n27590 );
not ( n35975 , n22191 );
nand ( n35976 , n35975 , n11080 );
nand ( n35977 , n35974 , n35976 );
buf ( n35978 , n35977 );
buf ( n35979 , n35978 );
or ( n35980 , n32627 , n26365 );
nand ( n35981 , n32653 , n26370 );
nand ( n35982 , n32679 , n26374 );
not ( n35983 , n13794 );
and ( n35984 , n17531 , n35983 );
not ( n35985 , n17531 );
and ( n35986 , n35985 , n13795 );
nor ( n35987 , n35984 , n35986 );
nor ( n35988 , n26390 , n35987 );
nand ( n35989 , n32689 , n26393 );
nand ( n35990 , n26395 , n32694 );
nand ( n35991 , n17542 , n13795 );
nand ( n35992 , n35989 , n35990 , n35991 );
nor ( n35993 , n35988 , n35992 );
and ( n35994 , n35981 , n35982 , n35993 );
nand ( n35995 , n35980 , n35994 );
buf ( n35996 , n35995 );
buf ( n35997 , n35996 );
or ( n35998 , n33527 , n27589 );
not ( n35999 , n22191 );
nand ( n36000 , n35999 , n11134 );
nand ( n36001 , n35998 , n36000 );
buf ( n36002 , n36001 );
buf ( n36003 , n36002 );
buf ( n36004 , n275554 );
buf ( n36005 , n275554 );
not ( n36006 , n275550 );
buf ( n36007 , n36006 );
buf ( n36008 , n36007 );
buf ( n36009 , n275554 );
buf ( n36010 , n275554 );
buf ( n36011 , n275554 );
not ( n36012 , n275925 );
buf ( n36013 , n36012 );
buf ( n36014 , n36013 );
not ( n36015 , n275925 );
buf ( n36016 , n36015 );
buf ( n36017 , n36016 );
buf ( n36018 , n275554 );
buf ( n36019 , n275554 );
buf ( n36020 , n275554 );
buf ( n36021 , n275554 );
not ( n36022 , n275925 );
buf ( n36023 , n36022 );
buf ( n36024 , n36023 );
buf ( n36025 , n275554 );
buf ( n36026 , n275554 );
not ( n36027 , n20616 );
not ( n36028 , n20637 );
or ( n36029 , n36027 , n36028 );
nand ( n36030 , n36029 , n9102 );
nand ( n36031 , n11730 , n36030 );
and ( n36032 , n20585 , n36031 );
not ( n36033 , n20585 );
and ( n36034 , n36033 , n9101 );
or ( n36035 , n36032 , n36034 );
buf ( n36036 , n36035 );
not ( n36037 , n11550 );
not ( n36038 , n36037 );
or ( n36039 , n36036 , n36038 );
not ( n36040 , n11730 );
not ( n36041 , n36040 );
not ( n36042 , n36030 );
or ( n36043 , n36041 , n36042 );
nand ( n36044 , n20627 , n20616 );
nand ( n36045 , n36043 , n36044 );
not ( n36046 , n36045 );
not ( n36047 , n36046 );
and ( n36048 , n36047 , n275657 );
buf ( n36049 , n36037 );
buf ( n36050 , n11538 );
not ( n36051 , n36050 );
nor ( n36052 , n36049 , n36051 );
not ( n36053 , n36052 );
nand ( n36054 , n36049 , n36051 );
nand ( n36055 , n36053 , n36054 );
not ( n36056 , n36055 );
buf ( n36057 , n11577 );
not ( n36058 , n36057 );
buf ( n36059 , n11616 );
nor ( n36060 , n36058 , n36059 );
not ( n36061 , n36060 );
buf ( n36062 , n11639 );
not ( n36063 , n36062 );
not ( n36064 , n11655 );
buf ( n36065 , n36064 );
nand ( n36066 , n36063 , n36065 );
nand ( n36067 , n36061 , n36066 );
not ( n36068 , n36067 );
not ( n36069 , n36068 );
buf ( n36070 , n10881 );
not ( n36071 , n36070 );
buf ( n36072 , n10841 );
nor ( n36073 , n36071 , n36072 );
not ( n36074 , n36073 );
buf ( n36075 , n10907 );
not ( n36076 , n36075 );
not ( n36077 , n10924 );
buf ( n36078 , n36077 );
nand ( n36079 , n36076 , n36078 );
not ( n36080 , n36079 );
or ( n36081 , n36074 , n36080 );
not ( n36082 , n36078 );
nand ( n36083 , n36082 , n36075 );
nand ( n36084 , n36081 , n36083 );
buf ( n36085 , n10780 );
not ( n36086 , n36085 );
buf ( n36087 , n26407 );
nand ( n36088 , n36086 , n36087 );
buf ( n36089 , n10765 );
not ( n36090 , n36089 );
buf ( n36091 , n10718 );
nand ( n36092 , n36090 , n36091 );
and ( n36093 , n36088 , n36092 );
and ( n36094 , n36084 , n36093 );
not ( n36095 , n36088 );
not ( n36096 , n36089 );
nor ( n36097 , n36096 , n36091 );
not ( n36098 , n36097 );
or ( n36099 , n36095 , n36098 );
not ( n36100 , n36087 );
nand ( n36101 , n36100 , n36085 );
nand ( n36102 , n36099 , n36101 );
nor ( n36103 , n36094 , n36102 );
not ( n36104 , n36070 );
nand ( n36105 , n36104 , n36072 );
and ( n36106 , n36079 , n36105 );
buf ( n36107 , n11092 );
not ( n36108 , n36107 );
not ( n36109 , n276323 );
not ( n36110 , n36109 );
buf ( n36111 , n36110 );
nand ( n36112 , n36108 , n36111 );
not ( n36113 , n36112 );
buf ( n36114 , n10996 );
xor ( n36115 , n36114 , n20623 );
buf ( n36116 , n10966 );
not ( n36117 , n36116 );
and ( n36118 , n36115 , n36117 );
and ( n36119 , n36114 , n20623 );
or ( n36120 , n36118 , n36119 );
buf ( n36121 , n11130 );
not ( n36122 , n36121 );
buf ( n36123 , n11144 );
nand ( n36124 , n36122 , n36123 );
and ( n36125 , n36120 , n36124 );
not ( n36126 , n36125 );
or ( n36127 , n36113 , n36126 );
not ( n36128 , n36123 );
nand ( n36129 , n36128 , n36121 );
not ( n36130 , n36129 );
and ( n36131 , n36112 , n36130 );
not ( n36132 , n36107 );
nor ( n36133 , n36132 , n36111 );
nor ( n36134 , n36131 , n36133 );
nand ( n36135 , n36127 , n36134 );
nand ( n36136 , n36106 , n36093 , n36135 );
nand ( n36137 , n36103 , n36136 );
not ( n36138 , n36137 );
or ( n36139 , n36069 , n36138 );
and ( n36140 , n36058 , n36059 );
not ( n36141 , n36140 );
not ( n36142 , n36066 );
or ( n36143 , n36141 , n36142 );
not ( n36144 , n36065 );
nand ( n36145 , n36144 , n36062 );
nand ( n36146 , n36143 , n36145 );
not ( n36147 , n36146 );
nand ( n36148 , n36139 , n36147 );
not ( n36149 , n36148 );
or ( n36150 , n36056 , n36149 );
or ( n36151 , n36148 , n36055 );
nand ( n36152 , n36150 , n36151 );
buf ( n36153 , n36152 );
not ( n36154 , n36153 );
nor ( n36155 , n20581 , n20616 );
not ( n36156 , n36155 );
or ( n36157 , n36154 , n36156 );
not ( n36158 , n20637 );
nor ( n36159 , n36158 , n20616 );
buf ( n36160 , n11522 );
not ( n36161 , n36160 );
buf ( n36162 , n36037 );
nor ( n36163 , n36161 , n36162 );
not ( n36164 , n36163 );
not ( n36165 , n36160 );
nand ( n36166 , n36165 , n36162 );
nand ( n36167 , n36164 , n36166 );
not ( n36168 , n36167 );
buf ( n36169 , n11577 );
not ( n36170 , n36169 );
buf ( n36171 , n11602 );
nor ( n36172 , n36170 , n36171 );
not ( n36173 , n36172 );
buf ( n36174 , n11626 );
not ( n36175 , n36174 );
buf ( n36176 , n36064 );
nand ( n36177 , n36175 , n36176 );
nand ( n36178 , n36173 , n36177 );
not ( n36179 , n36178 );
not ( n36180 , n36179 );
buf ( n36181 , n10874 );
not ( n36182 , n36181 );
buf ( n36183 , n10841 );
nor ( n36184 , n36182 , n36183 );
not ( n36185 , n36184 );
buf ( n36186 , n10902 );
not ( n36187 , n36186 );
buf ( n36188 , n36077 );
nand ( n36189 , n36187 , n36188 );
not ( n36190 , n36189 );
or ( n36191 , n36185 , n36190 );
not ( n36192 , n36188 );
nand ( n36193 , n36192 , n36186 );
nand ( n36194 , n36191 , n36193 );
buf ( n36195 , n10800 );
not ( n36196 , n36195 );
buf ( n36197 , n26407 );
nand ( n36198 , n36196 , n36197 );
buf ( n36199 , n10753 );
not ( n36200 , n36199 );
buf ( n36201 , n10718 );
nand ( n36202 , n36200 , n36201 );
and ( n36203 , n36198 , n36202 );
nand ( n36204 , n36194 , n36203 );
not ( n36205 , n36199 );
nor ( n36206 , n36205 , n36201 );
and ( n36207 , n36206 , n36198 );
not ( n36208 , n36195 );
nor ( n36209 , n36208 , n36197 );
nor ( n36210 , n36207 , n36209 );
nand ( n36211 , n36204 , n36210 );
not ( n36212 , n36181 );
nand ( n36213 , n36212 , n36183 );
and ( n36214 , n36189 , n36213 );
buf ( n36215 , n11073 );
not ( n36216 , n36215 );
buf ( n36217 , n36110 );
nand ( n36218 , n36216 , n36217 );
not ( n36219 , n36218 );
buf ( n36220 , n10991 );
xor ( n36221 , n20633 , n36220 );
buf ( n36222 , n10966 );
not ( n36223 , n36222 );
and ( n36224 , n36221 , n36223 );
and ( n36225 , n20633 , n36220 );
or ( n36226 , n36224 , n36225 );
buf ( n36227 , n11127 );
not ( n36228 , n36227 );
buf ( n36229 , n11144 );
nand ( n36230 , n36228 , n36229 );
and ( n36231 , n36226 , n36230 );
not ( n36232 , n36231 );
or ( n36233 , n36219 , n36232 );
not ( n36234 , n36229 );
nand ( n36235 , n36234 , n36227 );
not ( n36236 , n36235 );
and ( n36237 , n36218 , n36236 );
not ( n36238 , n36215 );
nor ( n36239 , n36238 , n36217 );
nor ( n36240 , n36237 , n36239 );
nand ( n36241 , n36233 , n36240 );
and ( n36242 , n36214 , n36203 , n36241 );
or ( n36243 , n36211 , n36242 );
not ( n36244 , n36243 );
or ( n36245 , n36180 , n36244 );
and ( n36246 , n36170 , n36171 );
not ( n36247 , n36246 );
not ( n36248 , n36177 );
or ( n36249 , n36247 , n36248 );
not ( n36250 , n36176 );
nand ( n36251 , n36250 , n36174 );
nand ( n36252 , n36249 , n36251 );
not ( n36253 , n36252 );
nand ( n36254 , n36245 , n36253 );
not ( n36255 , n36254 );
or ( n36256 , n36168 , n36255 );
or ( n36257 , n36254 , n36167 );
nand ( n36258 , n36256 , n36257 );
buf ( n36259 , n36258 );
nand ( n36260 , n36159 , n36259 );
nand ( n36261 , n36157 , n36260 );
nor ( n36262 , n36048 , n36261 );
nand ( n36263 , n36039 , n36262 );
nand ( n36264 , n36263 , n20645 );
or ( n36265 , n36031 , n20644 );
nand ( n36266 , n36265 , n20657 );
and ( n36267 , n36266 , n20580 );
buf ( n36268 , n36037 );
not ( n36269 , n36268 );
buf ( n36270 , n11538 );
nand ( n36271 , n36269 , n36270 );
not ( n36272 , n36268 );
nor ( n36273 , n36272 , n36270 );
not ( n36274 , n36273 );
nand ( n36275 , n36271 , n36274 );
not ( n36276 , n36275 );
buf ( n36277 , n36064 );
not ( n36278 , n36277 );
buf ( n36279 , n11639 );
nand ( n36280 , n36278 , n36279 );
buf ( n36281 , n11577 );
buf ( n36282 , n11616 );
not ( n36283 , n36282 );
or ( n36284 , n36281 , n36283 );
and ( n36285 , n36280 , n36284 );
not ( n36286 , n36285 );
buf ( n36287 , n26407 );
not ( n36288 , n36287 );
buf ( n36289 , n10780 );
nand ( n36290 , n36288 , n36289 );
buf ( n36291 , n10718 );
not ( n36292 , n36291 );
buf ( n36293 , n10765 );
nand ( n36294 , n36292 , n36293 );
and ( n36295 , n36290 , n36294 );
not ( n36296 , n36295 );
buf ( n36297 , n11130 );
not ( n36298 , n36297 );
buf ( n36299 , n11144 );
nand ( n36300 , n36298 , n36299 );
not ( n36301 , n36300 );
buf ( n36302 , n36110 );
not ( n36303 , n36302 );
buf ( n36304 , n11092 );
nand ( n36305 , n36303 , n36304 );
nand ( n36306 , n36301 , n36305 );
not ( n36307 , n36304 );
nand ( n36308 , n36307 , n36302 );
nand ( n36309 , n36306 , n36308 );
not ( n36310 , n36305 );
buf ( n36311 , n10996 );
not ( n36312 , n36311 );
xor ( n36313 , n20601 , n36312 );
buf ( n36314 , n10966 );
and ( n36315 , n36313 , n36314 );
and ( n36316 , n20601 , n36312 );
or ( n36317 , n36315 , n36316 );
not ( n36318 , n36299 );
nand ( n36319 , n36318 , n36297 );
nand ( n36320 , n36317 , n36319 );
nor ( n36321 , n36310 , n36320 );
nor ( n36322 , n36309 , n36321 );
buf ( n36323 , n36077 );
not ( n36324 , n36323 );
buf ( n36325 , n10907 );
nand ( n36326 , n36324 , n36325 );
buf ( n36327 , n10841 );
not ( n36328 , n36327 );
buf ( n36329 , n10881 );
nand ( n36330 , n36328 , n36329 );
nand ( n36331 , n36326 , n36330 );
nor ( n36332 , n36322 , n36331 );
not ( n36333 , n36332 );
or ( n36334 , n36296 , n36333 );
not ( n36335 , n36327 );
nor ( n36336 , n36335 , n36329 );
not ( n36337 , n36336 );
not ( n36338 , n36326 );
or ( n36339 , n36337 , n36338 );
not ( n36340 , n36325 );
nand ( n36341 , n36340 , n36323 );
nand ( n36342 , n36339 , n36341 );
and ( n36343 , n36295 , n36342 );
not ( n36344 , n36291 );
nor ( n36345 , n36344 , n36293 );
not ( n36346 , n36345 );
not ( n36347 , n36290 );
or ( n36348 , n36346 , n36347 );
not ( n36349 , n36289 );
nand ( n36350 , n36349 , n36287 );
nand ( n36351 , n36348 , n36350 );
nor ( n36352 , n36343 , n36351 );
nand ( n36353 , n36334 , n36352 );
not ( n36354 , n36353 );
or ( n36355 , n36286 , n36354 );
and ( n36356 , n36281 , n36283 );
not ( n36357 , n36356 );
not ( n36358 , n36280 );
or ( n36359 , n36357 , n36358 );
not ( n36360 , n36279 );
nand ( n36361 , n36360 , n36277 );
nand ( n36362 , n36359 , n36361 );
not ( n36363 , n36362 );
nand ( n36364 , n36355 , n36363 );
not ( n36365 , n36364 );
or ( n36366 , n36276 , n36365 );
or ( n36367 , n36364 , n36275 );
nand ( n36368 , n36366 , n36367 );
buf ( n36369 , n36368 );
nand ( n36370 , n36267 , n36369 );
and ( n36371 , n36266 , n20588 );
buf ( n36372 , n36037 );
not ( n36373 , n36372 );
buf ( n36374 , n11522 );
nand ( n36375 , n36373 , n36374 );
not ( n36376 , n36372 );
nor ( n36377 , n36376 , n36374 );
not ( n36378 , n36377 );
nand ( n36379 , n36375 , n36378 );
not ( n36380 , n36379 );
buf ( n36381 , n36064 );
not ( n36382 , n36381 );
buf ( n36383 , n11626 );
nand ( n36384 , n36382 , n36383 );
buf ( n36385 , n11577 );
not ( n36386 , n36385 );
buf ( n36387 , n11602 );
nand ( n36388 , n36386 , n36387 );
and ( n36389 , n36384 , n36388 );
not ( n36390 , n36389 );
buf ( n36391 , n26407 );
not ( n36392 , n36391 );
buf ( n36393 , n10800 );
nand ( n36394 , n36392 , n36393 );
buf ( n36395 , n10718 );
not ( n36396 , n36395 );
buf ( n36397 , n10753 );
nand ( n36398 , n36396 , n36397 );
and ( n36399 , n36394 , n36398 );
not ( n36400 , n36399 );
buf ( n36401 , n36110 );
not ( n36402 , n36401 );
buf ( n36403 , n11073 );
nand ( n36404 , n36402 , n36403 );
buf ( n36405 , n11144 );
not ( n36406 , n36405 );
buf ( n36407 , n11127 );
nor ( n36408 , n36406 , n36407 );
nand ( n36409 , n36404 , n36408 );
not ( n36410 , n36403 );
nand ( n36411 , n36410 , n36401 );
nand ( n36412 , n36409 , n36411 );
not ( n36413 , n36404 );
buf ( n36414 , n10991 );
not ( n36415 , n36414 );
xor ( n36416 , n20593 , n36415 );
buf ( n36417 , n10966 );
and ( n36418 , n36416 , n36417 );
and ( n36419 , n20593 , n36415 );
or ( n36420 , n36418 , n36419 );
not ( n36421 , n36405 );
nand ( n36422 , n36421 , n36407 );
nand ( n36423 , n36420 , n36422 );
nor ( n36424 , n36413 , n36423 );
nor ( n36425 , n36412 , n36424 );
buf ( n36426 , n36077 );
not ( n36427 , n36426 );
buf ( n36428 , n10902 );
nand ( n36429 , n36427 , n36428 );
buf ( n36430 , n10841 );
not ( n36431 , n36430 );
buf ( n36432 , n10874 );
nand ( n36433 , n36431 , n36432 );
nand ( n36434 , n36429 , n36433 );
nor ( n36435 , n36425 , n36434 );
not ( n36436 , n36435 );
or ( n36437 , n36400 , n36436 );
not ( n36438 , n36430 );
nor ( n36439 , n36438 , n36432 );
not ( n36440 , n36439 );
not ( n36441 , n36429 );
or ( n36442 , n36440 , n36441 );
not ( n36443 , n36428 );
nand ( n36444 , n36443 , n36426 );
nand ( n36445 , n36442 , n36444 );
and ( n36446 , n36399 , n36445 );
not ( n36447 , n36395 );
nor ( n36448 , n36447 , n36397 );
not ( n36449 , n36448 );
not ( n36450 , n36394 );
or ( n36451 , n36449 , n36450 );
not ( n36452 , n36393 );
nand ( n36453 , n36452 , n36391 );
nand ( n36454 , n36451 , n36453 );
nor ( n36455 , n36446 , n36454 );
nand ( n36456 , n36437 , n36455 );
not ( n36457 , n36456 );
or ( n36458 , n36390 , n36457 );
not ( n36459 , n36387 );
nand ( n36460 , n36459 , n36385 );
not ( n36461 , n36460 );
nand ( n36462 , n36461 , n36384 );
not ( n36463 , n36383 );
nand ( n36464 , n36463 , n36381 );
nand ( n36465 , n36462 , n36464 );
not ( n36466 , n36465 );
nand ( n36467 , n36458 , n36466 );
not ( n36468 , n36467 );
or ( n36469 , n36380 , n36468 );
or ( n36470 , n36467 , n36379 );
nand ( n36471 , n36469 , n36470 );
buf ( n36472 , n36471 );
nand ( n36473 , n36371 , n36472 );
nor ( n36474 , n20657 , n20586 );
and ( n36475 , n36474 , n36037 );
or ( n36476 , n20654 , n275656 );
nand ( n36477 , n20649 , n9315 );
nand ( n36478 , n36476 , n36477 );
nor ( n36479 , n36475 , n36478 );
nand ( n36480 , n36264 , n36370 , n36473 , n36479 );
buf ( n36481 , n36480 );
buf ( n36482 , n36481 );
not ( n36483 , n11366 );
or ( n36484 , n36483 , n9158 );
not ( n36485 , n11343 );
or ( n36486 , n36485 , n9157 );
nand ( n36487 , n36484 , n36486 );
buf ( n36488 , n36487 );
buf ( n36489 , n36488 );
xor ( n36490 , n31683 , n31687 );
and ( n36491 , n36490 , n31693 );
and ( n36492 , n31683 , n31687 );
or ( n36493 , n36491 , n36492 );
buf ( n36494 , RI21a12910_76);
not ( n36495 , n36494 );
not ( n36496 , n36495 );
buf ( n36497 , n36496 );
buf ( n36498 , RI210bf3f0_290);
not ( n36499 , n36498 );
not ( n36500 , n36499 );
buf ( n36501 , n36500 );
xor ( n36502 , n36497 , n36501 );
buf ( n36503 , RI21078a40_505);
not ( n36504 , n36503 );
not ( n36505 , n36504 );
buf ( n36506 , n36505 );
not ( n36507 , n36506 );
xor ( n36508 , n36502 , n36507 );
xor ( n36509 , n36493 , n36508 );
or ( n36510 , n31712 , n31701 );
nand ( n36511 , n36510 , n31699 );
xor ( n36512 , n36509 , n36511 );
buf ( n36513 , n36512 );
buf ( n36514 , n36513 );
or ( n36515 , n34423 , n14908 );
and ( n36516 , n34499 , n20763 );
nand ( n36517 , n35653 , n17545 , n14641 );
nand ( n36518 , n20785 , n24939 );
nand ( n36519 , n32339 , n34510 );
nand ( n36520 , n17562 , n14654 );
nand ( n36521 , n36517 , n36518 , n36519 , n36520 );
nor ( n36522 , n36516 , n36521 );
nand ( n36523 , n34463 , n16970 );
nand ( n36524 , n36515 , n36522 , n36523 );
buf ( n36525 , n36524 );
buf ( n36526 , n36525 );
nand ( n36527 , n29702 , n31422 );
nand ( n36528 , n29747 , n31437 );
nand ( n36529 , n29764 , n31449 );
not ( n36530 , n32053 );
and ( n36531 , n36530 , n12355 );
not ( n36532 , n277961 );
or ( n36533 , n31453 , n36532 );
nand ( n36534 , n28236 , n277973 );
nand ( n36535 , n36533 , n36534 );
nor ( n36536 , n36531 , n36535 );
nand ( n36537 , n28242 , n12156 );
and ( n36538 , n36529 , n36536 , n36537 );
nand ( n36539 , n36527 , n36528 , n36538 );
buf ( n36540 , n36539 );
buf ( n36541 , n36540 );
not ( n36542 , n275929 );
buf ( n36543 , n36542 );
buf ( n36544 , n36543 );
buf ( n36545 , n275554 );
buf ( n36546 , n275554 );
buf ( n36547 , n275554 );
buf ( n36548 , n275554 );
not ( n36549 , n275929 );
buf ( n36550 , n36549 );
buf ( n36551 , n36550 );
buf ( n36552 , n275554 );
buf ( n36553 , n275554 );
or ( n36554 , n24448 , n21030 );
nand ( n36555 , n21030 , n18387 );
nand ( n36556 , n36554 , n36555 );
buf ( n36557 , n36556 );
buf ( n36558 , n36557 );
not ( n36559 , n24814 );
or ( n36560 , n36559 , n28252 );
nand ( n36561 , n29046 , n277336 );
nand ( n36562 , n36560 , n36561 );
buf ( n36563 , n36562 );
buf ( n36564 , n36563 );
buf ( n36565 , n275554 );
not ( n36566 , n275929 );
buf ( n36567 , n36566 );
buf ( n36568 , n36567 );
not ( n36569 , n11594 );
or ( n36570 , n36569 , n9158 );
not ( n36571 , n11577 );
or ( n36572 , n9157 , n36571 );
nand ( n36573 , n36570 , n36572 );
buf ( n36574 , n36573 );
buf ( n36575 , n36574 );
buf ( n36576 , n275554 );
and ( n36577 , n14830 , n13369 );
not ( n36578 , n14830 );
and ( n36579 , n36578 , n24935 );
or ( n36580 , n36577 , n36579 );
buf ( n36581 , n36580 );
buf ( n36582 , n36581 );
or ( n36583 , n35683 , n19216 );
nand ( n36584 , n35693 , n35150 );
nand ( n36585 , n35702 , n19360 );
and ( n36586 , n35709 , n29075 );
not ( n36587 , n18345 );
not ( n36588 , n19657 );
not ( n36589 , n36588 );
or ( n36590 , n36587 , n36589 );
or ( n36591 , n36588 , n18345 );
nand ( n36592 , n36590 , n36591 );
not ( n36593 , n36592 );
nor ( n36594 , n36593 , n19317 );
nor ( n36595 , n36586 , n36594 );
nand ( n36596 , n19221 , n35714 );
nand ( n36597 , n19387 , n18335 );
and ( n36598 , n36595 , n36596 , n36597 );
and ( n36599 , n36584 , n36585 , n36598 );
nand ( n36600 , n36583 , n36599 );
buf ( n36601 , n36600 );
buf ( n36602 , n36601 );
buf ( n36603 , n275554 );
not ( n36604 , n275929 );
buf ( n36605 , n36604 );
buf ( n36606 , n36605 );
or ( n36607 , n34672 , n20953 );
nand ( n36608 , n20950 , n13682 );
nand ( n36609 , n36607 , n36608 );
buf ( n36610 , n36609 );
buf ( n36611 , n36610 );
not ( n36612 , n275925 );
buf ( n36613 , n36612 );
buf ( n36614 , n36613 );
not ( n36615 , n24672 );
or ( n36616 , n36615 , n29044 );
nand ( n36617 , n28252 , n9496 );
nand ( n36618 , n36616 , n36617 );
buf ( n36619 , n36618 );
buf ( n36620 , n36619 );
and ( n36621 , n20711 , n14542 );
not ( n36622 , n20711 );
not ( n36623 , n34686 );
not ( n36624 , n34687 );
and ( n36625 , n36623 , n36624 );
not ( n36626 , n36623 );
and ( n36627 , n36626 , n34687 );
nor ( n36628 , n36625 , n36627 );
buf ( n36629 , n36628 );
and ( n36630 , n36622 , n36629 );
nor ( n36631 , n36621 , n36630 );
or ( n36632 , n36631 , n14908 );
xor ( n36633 , n17431 , n34728 );
buf ( n36634 , n36633 );
nand ( n36635 , n32339 , n36634 );
buf ( n36636 , n16753 );
buf ( n36637 , n36636 );
buf ( n36638 , n36637 );
nand ( n36639 , n20785 , n36638 );
not ( n36640 , n17299 );
nand ( n36641 , n17310 , n17314 );
not ( n36642 , n36641 );
or ( n36643 , n36640 , n36642 );
or ( n36644 , n36641 , n17299 );
nand ( n36645 , n36643 , n36644 );
buf ( n36646 , n36645 );
and ( n36647 , n17405 , n36646 );
not ( n36648 , n14549 );
nor ( n36649 , n17561 , n36648 );
nor ( n36650 , n36647 , n36649 );
not ( n36651 , n20765 );
not ( n36652 , n14544 );
not ( n36653 , n36652 );
and ( n36654 , n36651 , n36653 );
nand ( n36655 , n16803 , n16760 );
not ( n36656 , n36655 );
not ( n36657 , n16727 );
or ( n36658 , n36657 , n16724 );
nand ( n36659 , n36658 , n16707 );
not ( n36660 , n36659 );
or ( n36661 , n36656 , n36660 );
or ( n36662 , n36655 , n36659 );
nand ( n36663 , n36661 , n36662 );
buf ( n36664 , n36663 );
and ( n36665 , n36664 , n16968 );
nor ( n36666 , n36654 , n36665 );
and ( n36667 , n36635 , n36639 , n36650 , n36666 );
nand ( n36668 , n36632 , n36667 );
buf ( n36669 , n36668 );
buf ( n36670 , n36669 );
or ( n36671 , n275860 , n275684 );
not ( n36672 , n36671 );
or ( n36673 , n32738 , n275665 );
nand ( n36674 , n36673 , n275856 );
not ( n36675 , n36674 );
or ( n36676 , n36672 , n36675 );
or ( n36677 , n36674 , n36671 );
nand ( n36678 , n36676 , n36677 );
buf ( n36679 , n36678 );
buf ( n36680 , n36679 );
buf ( n36681 , n275554 );
not ( n36682 , n19156 );
or ( n36683 , n19143 , n36682 );
nand ( n36684 , n36683 , n19163 );
buf ( n36685 , n36684 );
buf ( n36686 , n36685 );
not ( n36687 , n275550 );
buf ( n36688 , n36687 );
buf ( n36689 , n36688 );
nand ( n36690 , n25064 , n25087 );
buf ( n36691 , n25337 );
not ( n36692 , n36691 );
buf ( n36693 , n25093 );
nor ( n36694 , n36692 , n36693 );
buf ( n36695 , n36694 );
buf ( n36696 , n36695 );
not ( n36697 , n36696 );
buf ( n36698 , n25264 );
buf ( n36699 , n25128 );
buf ( n36700 , n25103 );
not ( n36701 , n36700 );
buf ( n36702 , n36701 );
buf ( n36703 , n36702 );
and ( n36704 , n36698 , n36699 , n36703 );
buf ( n36705 , n36702 );
not ( n36706 , n36705 );
buf ( n36707 , n25329 );
not ( n36708 , n36707 );
or ( n36709 , n36706 , n36708 );
buf ( n36710 , n25309 );
nand ( n36711 , n36709 , n36710 );
buf ( n36712 , n36711 );
buf ( n36713 , n36712 );
nor ( n36714 , n36704 , n36713 );
buf ( n36715 , n36714 );
buf ( n36716 , n36715 );
not ( n36717 , n36716 );
or ( n36718 , n36697 , n36717 );
buf ( n36719 , n36715 );
buf ( n36720 , n36695 );
or ( n36721 , n36719 , n36720 );
nand ( n36722 , n36718 , n36721 );
buf ( n36723 , n36722 );
buf ( n36724 , n36723 );
not ( n36725 , n36724 );
nor ( n36726 , n36725 , n25389 );
nand ( n36727 , n25397 , n275668 );
buf ( n36728 , n25425 );
buf ( n36729 , n25660 );
nor ( n36730 , n36728 , n36729 );
buf ( n36731 , n36730 );
buf ( n36732 , n36731 );
not ( n36733 , n36732 );
buf ( n36734 , n25586 );
buf ( n36735 , n25453 );
buf ( n36736 , n25432 );
not ( n36737 , n36736 );
buf ( n36738 , n36737 );
buf ( n36739 , n36738 );
and ( n36740 , n36734 , n36735 , n36739 );
buf ( n36741 , n36738 );
not ( n36742 , n36741 );
buf ( n36743 , n25642 );
not ( n36744 , n36743 );
or ( n36745 , n36742 , n36744 );
buf ( n36746 , n25653 );
nand ( n36747 , n36745 , n36746 );
buf ( n36748 , n36747 );
buf ( n36749 , n36748 );
nor ( n36750 , n36740 , n36749 );
buf ( n36751 , n36750 );
buf ( n36752 , n36751 );
not ( n36753 , n36752 );
or ( n36754 , n36733 , n36753 );
buf ( n36755 , n36751 );
buf ( n36756 , n36731 );
or ( n36757 , n36755 , n36756 );
nand ( n36758 , n36754 , n36757 );
buf ( n36759 , n36758 );
buf ( n36760 , n36759 );
and ( n36761 , n25402 , n36760 );
not ( n36762 , n18749 );
nor ( n36763 , n19639 , n36762 );
nor ( n36764 , n36761 , n36763 );
buf ( n36765 , n25974 );
buf ( n36766 , n25741 );
and ( n36767 , n36765 , n36766 );
buf ( n36768 , n36767 );
buf ( n36769 , n36768 );
not ( n36770 , n36769 );
buf ( n36771 , n25902 );
buf ( n36772 , n25770 );
buf ( n36773 , n25748 );
and ( n36774 , n36771 , n36772 , n36773 );
buf ( n36775 , n25748 );
not ( n36776 , n36775 );
buf ( n36777 , n25956 );
not ( n36778 , n36777 );
or ( n36779 , n36776 , n36778 );
buf ( n36780 , n25964 );
nand ( n36781 , n36779 , n36780 );
buf ( n36782 , n36781 );
buf ( n36783 , n36782 );
nor ( n36784 , n36774 , n36783 );
buf ( n36785 , n36784 );
buf ( n36786 , n36785 );
not ( n36787 , n36786 );
or ( n36788 , n36770 , n36787 );
buf ( n36789 , n36785 );
buf ( n36790 , n36768 );
or ( n36791 , n36789 , n36790 );
nand ( n36792 , n36788 , n36791 );
buf ( n36793 , n36792 );
buf ( n36794 , n36793 );
nand ( n36795 , n25717 , n36794 );
nand ( n36796 , n36727 , n36764 , n36795 );
nor ( n36797 , n36726 , n36796 );
buf ( n36798 , n26278 );
not ( n36799 , n36798 );
buf ( n36800 , n26058 );
nor ( n36801 , n36799 , n36800 );
buf ( n36802 , n36801 );
buf ( n36803 , n36802 );
not ( n36804 , n36803 );
buf ( n36805 , n26212 );
buf ( n36806 , n26078 );
buf ( n36807 , n26050 );
and ( n36808 , n36805 , n36806 , n36807 );
buf ( n36809 , n26050 );
not ( n36810 , n36809 );
buf ( n36811 , n26270 );
not ( n36812 , n36811 );
or ( n36813 , n36810 , n36812 );
buf ( n36814 , n26253 );
nand ( n36815 , n36813 , n36814 );
buf ( n36816 , n36815 );
buf ( n36817 , n36816 );
nor ( n36818 , n36808 , n36817 );
buf ( n36819 , n36818 );
buf ( n36820 , n36819 );
not ( n36821 , n36820 );
or ( n36822 , n36804 , n36821 );
buf ( n36823 , n36819 );
buf ( n36824 , n36802 );
or ( n36825 , n36823 , n36824 );
nand ( n36826 , n36822 , n36825 );
buf ( n36827 , n36826 );
buf ( n36828 , n36827 );
nand ( n36829 , n26027 , n36828 );
nand ( n36830 , n36690 , n36797 , n36829 );
buf ( n36831 , n36830 );
buf ( n36832 , n36831 );
buf ( n36833 , n275554 );
not ( n36834 , n32154 );
and ( n36835 , n36834 , n23788 );
nand ( n36836 , n32164 , n20889 );
nand ( n36837 , n32174 , n24711 );
and ( n36838 , n32187 , n17409 );
and ( n36839 , n20940 , n32192 );
nor ( n36840 , n36838 , n36839 );
nand ( n36841 , n36836 , n36837 , n36840 );
nor ( n36842 , n36835 , n36841 );
or ( n36843 , n36842 , n20953 );
nand ( n36844 , n20950 , n13635 );
nand ( n36845 , n36843 , n36844 );
buf ( n36846 , n36845 );
buf ( n36847 , n36846 );
buf ( n36848 , n9157 );
buf ( n36849 , n36848 );
not ( n36850 , n275925 );
buf ( n36851 , n36850 );
buf ( n36852 , n36851 );
or ( n36853 , n24330 , n24452 );
nand ( n36854 , n28146 , n18930 );
nand ( n36855 , n36853 , n36854 );
buf ( n36856 , n36855 );
buf ( n36857 , n36856 );
not ( n36858 , n10958 );
not ( n36859 , n9157 );
or ( n36860 , n36858 , n36859 );
not ( n36861 , n36077 );
or ( n36862 , n9157 , n36861 );
nand ( n36863 , n36860 , n36862 );
buf ( n36864 , n36863 );
buf ( n36865 , n36864 );
not ( n36866 , n20713 );
or ( n36867 , n36866 , n29044 );
nand ( n36868 , n29046 , n9675 );
nand ( n36869 , n36867 , n36868 );
buf ( n36870 , n36869 );
buf ( n36871 , n36870 );
not ( n36872 , n275929 );
buf ( n36873 , n36872 );
buf ( n36874 , n36873 );
buf ( n36875 , n275554 );
not ( n36876 , n275925 );
buf ( n36877 , n36876 );
buf ( n36878 , n36877 );
not ( n36879 , n23403 );
or ( n36880 , n36879 , n20743 );
and ( n36881 , n23433 , n20763 );
nand ( n36882 , n32339 , n23442 );
nand ( n36883 , n20785 , n23447 );
nand ( n36884 , n17560 , n13757 );
and ( n36885 , n17522 , n17523 );
not ( n36886 , n17522 );
and ( n36887 , n36886 , n13746 );
nor ( n36888 , n36885 , n36887 );
nand ( n36889 , n17545 , n36888 );
nand ( n36890 , n36882 , n36883 , n36884 , n36889 );
nor ( n36891 , n36881 , n36890 );
nand ( n36892 , n23418 , n16970 );
and ( n36893 , n36891 , n36892 );
nand ( n36894 , n36880 , n36893 );
buf ( n36895 , n36894 );
buf ( n36896 , n36895 );
buf ( n36897 , n275554 );
not ( n36898 , n26423 );
or ( n36899 , n36898 , n29046 );
nand ( n36900 , n28252 , n9575 );
nand ( n36901 , n36899 , n36900 );
buf ( n36902 , n36901 );
buf ( n36903 , n36902 );
not ( n36904 , n275925 );
buf ( n36905 , n36904 );
buf ( n36906 , n36905 );
buf ( n36907 , n275554 );
buf ( n36908 , n275554 );
and ( n36909 , n14830 , n13226 );
not ( n36910 , n14830 );
and ( n36911 , n36910 , n15962 );
or ( n36912 , n36909 , n36911 );
buf ( n36913 , n36912 );
buf ( n36914 , n36913 );
not ( n36915 , n275550 );
buf ( n36916 , n36915 );
buf ( n36917 , n36916 );
not ( n36918 , n275929 );
buf ( n36919 , n36918 );
buf ( n36920 , n36919 );
buf ( n36921 , n275554 );
not ( n36922 , n34302 );
not ( n36923 , n29702 );
or ( n36924 , n36922 , n36923 );
and ( n36925 , n29747 , n35900 );
nand ( n36926 , n29764 , n34307 );
nand ( n36927 , n28451 , n277973 );
nand ( n36928 , n29171 , n12355 );
nand ( n36929 , n34311 , n12156 );
nand ( n36930 , n20649 , n9329 );
and ( n36931 , n36928 , n36929 , n36930 );
nand ( n36932 , n36926 , n36927 , n36931 );
nor ( n36933 , n36925 , n36932 );
nand ( n36934 , n36924 , n36933 );
buf ( n36935 , n36934 );
buf ( n36936 , n36935 );
buf ( n36937 , n275554 );
not ( n36938 , n275929 );
buf ( n36939 , n36938 );
buf ( n36940 , n36939 );
not ( n36941 , n275925 );
buf ( n36942 , n36941 );
buf ( n36943 , n36942 );
buf ( n36944 , n275554 );
not ( n36945 , n20820 );
or ( n36946 , n36945 , n29046 );
nand ( n36947 , n28252 , n9505 );
nand ( n36948 , n36946 , n36947 );
buf ( n36949 , n36948 );
buf ( n36950 , n36949 );
buf ( n36951 , n275554 );
not ( n36952 , n275925 );
buf ( n36953 , n36952 );
buf ( n36954 , n36953 );
buf ( n36955 , n275554 );
not ( n36956 , n275550 );
buf ( n36957 , n36956 );
buf ( n36958 , n36957 );
buf ( n36959 , n275554 );
not ( n36960 , n34302 );
not ( n36961 , n35012 );
or ( n36962 , n36960 , n36961 );
and ( n36963 , n35037 , n28430 );
nand ( n36964 , n35044 , n34307 );
nand ( n36965 , n28451 , n277625 );
and ( n36966 , n32755 , n12198 );
and ( n36967 , n34311 , n12365 );
and ( n36968 , n34313 , n9350 );
nor ( n36969 , n36966 , n36967 , n36968 );
nand ( n36970 , n36964 , n36965 , n36969 );
nor ( n36971 , n36963 , n36970 );
nand ( n36972 , n36962 , n36971 );
buf ( n36973 , n36972 );
buf ( n36974 , n36973 );
not ( n36975 , n30610 );
and ( n36976 , n36975 , n20987 );
not ( n36977 , n19358 );
not ( n36978 , n30649 );
or ( n36979 , n36977 , n36978 );
and ( n36980 , n30624 , n21001 );
or ( n36981 , n30636 , n19289 );
or ( n36982 , n24440 , n30629 );
nand ( n36983 , n36981 , n36982 );
nor ( n36984 , n36980 , n36983 );
nand ( n36985 , n36979 , n36984 );
nor ( n36986 , n36976 , n36985 );
or ( n36987 , n36986 , n24450 );
nand ( n36988 , n24450 , n18368 );
nand ( n36989 , n36987 , n36988 );
buf ( n36990 , n36989 );
buf ( n36991 , n36990 );
not ( n36992 , n11331 );
or ( n36993 , n36992 , n9158 );
not ( n36994 , n11302 );
or ( n36995 , n36994 , n9157 );
nand ( n36996 , n36993 , n36995 );
buf ( n36997 , n36996 );
buf ( n36998 , n36997 );
not ( n36999 , n25119 );
not ( n37000 , n22335 );
or ( n37001 , n36999 , n37000 );
nand ( n37002 , n19977 , n275557 );
nand ( n37003 , n37001 , n37002 );
buf ( n37004 , n37003 );
buf ( n37005 , n37004 );
buf ( n37006 , n275554 );
not ( n37007 , n275929 );
buf ( n37008 , n37007 );
buf ( n37009 , n37008 );
buf ( n37010 , n275554 );
not ( n37011 , n275550 );
buf ( n37012 , n37011 );
buf ( n37013 , n37012 );
buf ( n37014 , n275554 );
not ( n37015 , n34157 );
or ( n37016 , n37015 , n21774 );
nand ( n37017 , n21774 , n277460 );
nand ( n37018 , n37016 , n37017 );
buf ( n37019 , n37018 );
buf ( n37020 , n37019 );
buf ( n37021 , n275554 );
not ( n37022 , n275925 );
buf ( n37023 , n37022 );
buf ( n37024 , n37023 );
not ( n37025 , n275550 );
buf ( n37026 , n37025 );
buf ( n37027 , n37026 );
buf ( n37028 , n275554 );
not ( n37029 , n275929 );
buf ( n37030 , n37029 );
buf ( n37031 , n37030 );
not ( n37032 , n275925 );
buf ( n37033 , n37032 );
buf ( n37034 , n37033 );
not ( n37035 , n13976 );
or ( n37036 , n37035 , n29046 );
nand ( n37037 , n28252 , n9765 );
nand ( n37038 , n37036 , n37037 );
buf ( n37039 , n37038 );
buf ( n37040 , n37039 );
and ( n37041 , n22193 , n278013 );
not ( n37042 , n22193 );
not ( n37043 , n29599 );
buf ( n37044 , n29671 );
buf ( n37045 , n29649 );
nand ( n37046 , n37044 , n37045 );
buf ( n37047 , n37046 );
buf ( n37048 , n37047 );
not ( n37049 , n37048 );
buf ( n37050 , n27281 );
not ( n37051 , n37050 );
buf ( n37052 , n27479 );
not ( n37053 , n37052 );
or ( n37054 , n37051 , n37053 );
buf ( n37055 , n27276 );
nand ( n37056 , n37054 , n37055 );
buf ( n37057 , n37056 );
buf ( n37058 , n37057 );
not ( n37059 , n37058 );
or ( n37060 , n37049 , n37059 );
buf ( n37061 , n37057 );
buf ( n37062 , n37047 );
or ( n37063 , n37061 , n37062 );
nand ( n37064 , n37060 , n37063 );
buf ( n37065 , n37064 );
buf ( n37066 , n37065 );
not ( n37067 , n37066 );
or ( n37068 , n37043 , n37067 );
nand ( n37069 , n29723 , n29735 );
not ( n37070 , n37069 );
not ( n37071 , n27185 );
not ( n37072 , n29728 );
or ( n37073 , n37071 , n37072 );
nand ( n37074 , n37073 , n27187 );
not ( n37075 , n37074 );
or ( n37076 , n37070 , n37075 );
or ( n37077 , n37074 , n37069 );
nand ( n37078 , n37076 , n37077 );
buf ( n37079 , n37078 );
and ( n37080 , n37079 , n23655 );
not ( n37081 , n22052 );
xnor ( n37082 , n31441 , n29755 );
buf ( n37083 , n37082 );
not ( n37084 , n37083 );
or ( n37085 , n37081 , n37084 );
and ( n37086 , n22007 , n12288 );
and ( n37087 , n23679 , n12295 );
nor ( n37088 , n37086 , n37087 );
nand ( n37089 , n37085 , n37088 );
nor ( n37090 , n37080 , n37089 );
nand ( n37091 , n37068 , n37090 );
and ( n37092 , n37042 , n37091 );
or ( n37093 , n37041 , n37092 );
buf ( n37094 , n37093 );
buf ( n37095 , n37094 );
not ( n37096 , n275550 );
buf ( n37097 , n37096 );
buf ( n37098 , n37097 );
buf ( n37099 , n275554 );
not ( n37100 , n275550 );
buf ( n37101 , n37100 );
buf ( n37102 , n37101 );
not ( n37103 , n36631 );
not ( n37104 , n23789 );
and ( n37105 , n37103 , n37104 );
not ( n37106 , n20927 );
not ( n37107 , n36646 );
or ( n37108 , n37106 , n37107 );
and ( n37109 , n36664 , n20889 );
and ( n37110 , n36634 , n17409 );
and ( n37111 , n17499 , n36638 );
nor ( n37112 , n37110 , n37111 );
not ( n37113 , n37112 );
nor ( n37114 , n37109 , n37113 );
nand ( n37115 , n37108 , n37114 );
nor ( n37116 , n37105 , n37115 );
or ( n37117 , n37116 , n27647 );
nand ( n37118 , n21696 , n14554 );
nand ( n37119 , n37117 , n37118 );
buf ( n37120 , n37119 );
buf ( n37121 , n37120 );
not ( n37122 , n275550 );
buf ( n37123 , n37122 );
buf ( n37124 , n37123 );
not ( n37125 , n275925 );
buf ( n37126 , n37125 );
buf ( n37127 , n37126 );
nand ( n37128 , n25064 , n28957 );
buf ( n37129 , n28543 );
not ( n37130 , n37129 );
buf ( n37131 , n37130 );
buf ( n37132 , n37131 );
buf ( n37133 , n28586 );
nand ( n37134 , n37132 , n37133 );
buf ( n37135 , n37134 );
buf ( n37136 , n37135 );
not ( n37137 , n37136 );
buf ( n37138 , n35262 );
buf ( n37139 , n28523 );
not ( n37140 , n37139 );
buf ( n37141 , n37140 );
buf ( n37142 , n37141 );
or ( n37143 , n37138 , n37142 );
buf ( n37144 , n25131 );
buf ( n37145 , n28523 );
buf ( n37146 , n25264 );
nand ( n37147 , n37144 , n37145 , n37146 );
buf ( n37148 , n37147 );
buf ( n37149 , n37148 );
buf ( n37150 , n28573 );
nand ( n37151 , n37143 , n37149 , n37150 );
buf ( n37152 , n37151 );
buf ( n37153 , n37152 );
not ( n37154 , n37153 );
or ( n37155 , n37137 , n37154 );
buf ( n37156 , n37152 );
buf ( n37157 , n37135 );
or ( n37158 , n37156 , n37157 );
nand ( n37159 , n37155 , n37158 );
buf ( n37160 , n37159 );
buf ( n37161 , n37160 );
not ( n37162 , n37161 );
nor ( n37163 , n37162 , n25389 );
nand ( n37164 , n25397 , n31686 );
buf ( n37165 , n28691 );
not ( n37166 , n37165 );
buf ( n37167 , n37166 );
buf ( n37168 , n37167 );
buf ( n37169 , n28723 );
and ( n37170 , n37168 , n37169 );
buf ( n37171 , n37170 );
buf ( n37172 , n37171 );
not ( n37173 , n37172 );
buf ( n37174 , n25456 );
buf ( n37175 , n28667 );
buf ( n37176 , n25586 );
and ( n37177 , n37174 , n37175 , n37176 );
buf ( n37178 , n35297 );
buf ( n37179 , n28664 );
or ( n37180 , n37178 , n37179 );
buf ( n37181 , n28714 );
nand ( n37182 , n37180 , n37181 );
buf ( n37183 , n37182 );
buf ( n37184 , n37183 );
nor ( n37185 , n37177 , n37184 );
buf ( n37186 , n37185 );
buf ( n37187 , n37186 );
not ( n37188 , n37187 );
or ( n37189 , n37173 , n37188 );
buf ( n37190 , n37186 );
buf ( n37191 , n37171 );
or ( n37192 , n37190 , n37191 );
nand ( n37193 , n37189 , n37192 );
buf ( n37194 , n37193 );
buf ( n37195 , n37194 );
and ( n37196 , n25402 , n37195 );
nor ( n37197 , n19639 , n29481 );
nor ( n37198 , n37196 , n37197 );
buf ( n37199 , n28832 );
not ( n37200 , n37199 );
buf ( n37201 , n37200 );
buf ( n37202 , n37201 );
buf ( n37203 , n28864 );
and ( n37204 , n37202 , n37203 );
buf ( n37205 , n37204 );
buf ( n37206 , n37205 );
not ( n37207 , n37206 );
buf ( n37208 , n25773 );
buf ( n37209 , n28808 );
buf ( n37210 , n25902 );
and ( n37211 , n37208 , n37209 , n37210 );
buf ( n37212 , n35332 );
buf ( n37213 , n28805 );
or ( n37214 , n37212 , n37213 );
buf ( n37215 , n28855 );
nand ( n37216 , n37214 , n37215 );
buf ( n37217 , n37216 );
buf ( n37218 , n37217 );
nor ( n37219 , n37211 , n37218 );
buf ( n37220 , n37219 );
buf ( n37221 , n37220 );
not ( n37222 , n37221 );
or ( n37223 , n37207 , n37222 );
buf ( n37224 , n37220 );
buf ( n37225 , n37205 );
or ( n37226 , n37224 , n37225 );
nand ( n37227 , n37223 , n37226 );
buf ( n37228 , n37227 );
buf ( n37229 , n37228 );
nand ( n37230 , n28761 , n37229 );
nand ( n37231 , n37164 , n37198 , n37230 );
nor ( n37232 , n37163 , n37231 );
buf ( n37233 , n28964 );
not ( n37234 , n37233 );
buf ( n37235 , n37234 );
buf ( n37236 , n37235 );
buf ( n37237 , n29005 );
and ( n37238 , n37236 , n37237 );
buf ( n37239 , n37238 );
buf ( n37240 , n37239 );
not ( n37241 , n37240 );
buf ( n37242 , n26081 );
buf ( n37243 , n28947 );
buf ( n37244 , n26212 );
and ( n37245 , n37242 , n37243 , n37244 );
buf ( n37246 , n35367 );
buf ( n37247 , n28944 );
or ( n37248 , n37246 , n37247 );
buf ( n37249 , n28992 );
nand ( n37250 , n37248 , n37249 );
buf ( n37251 , n37250 );
buf ( n37252 , n37251 );
nor ( n37253 , n37245 , n37252 );
buf ( n37254 , n37253 );
buf ( n37255 , n37254 );
not ( n37256 , n37255 );
or ( n37257 , n37241 , n37256 );
buf ( n37258 , n37254 );
buf ( n37259 , n37239 );
or ( n37260 , n37258 , n37259 );
nand ( n37261 , n37257 , n37260 );
buf ( n37262 , n37261 );
buf ( n37263 , n37262 );
nand ( n37264 , n26027 , n37263 );
nand ( n37265 , n37128 , n37232 , n37264 );
buf ( n37266 , n37265 );
buf ( n37267 , n37266 );
not ( n37268 , n275925 );
buf ( n37269 , n37268 );
buf ( n37270 , n37269 );
not ( n37271 , n31467 );
and ( n37272 , n37271 , n36496 );
nor ( n37273 , n26386 , n17523 );
nor ( n37274 , n37272 , n37273 );
buf ( n37275 , n12799 );
nand ( n37276 , n22914 , n37275 );
buf ( n37277 , n37275 );
buf ( n37278 , n37277 );
buf ( n37279 , n37278 );
buf ( n37280 , n13750 );
buf ( n37281 , n37280 );
nor ( n37282 , n37279 , n37281 );
buf ( n37283 , n37282 );
buf ( n37284 , n37283 );
buf ( n37285 , n37278 );
buf ( n37286 , n37280 );
and ( n37287 , n37285 , n37286 );
buf ( n37288 , n37287 );
buf ( n37289 , n37288 );
nor ( n37290 , n37284 , n37289 );
buf ( n37291 , n37290 );
buf ( n37292 , n37291 );
not ( n37293 , n37292 );
buf ( n37294 , n23140 );
buf ( n37295 , n31484 );
buf ( n37296 , n31514 );
nor ( n37297 , n37295 , n37296 );
buf ( n37298 , n37297 );
buf ( n37299 , n37298 );
buf ( n37300 , n31506 );
nand ( n37301 , n37299 , n37300 );
buf ( n37302 , n37301 );
buf ( n37303 , n37302 );
not ( n37304 , n37303 );
buf ( n37305 , n37304 );
buf ( n37306 , n37305 );
buf ( n37307 , n34525 );
buf ( n37308 , n37307 );
buf ( n37309 , n37308 );
buf ( n37310 , n13774 );
buf ( n37311 , n37310 );
nor ( n37312 , n37309 , n37311 );
buf ( n37313 , n37312 );
buf ( n37314 , n37313 );
not ( n37315 , n37314 );
buf ( n37316 , n37315 );
buf ( n37317 , n37316 );
and ( n37318 , n37294 , n37306 , n37317 );
buf ( n37319 , n37298 );
buf ( n37320 , n31537 );
and ( n37321 , n37319 , n37320 );
buf ( n37322 , n31484 );
buf ( n37323 , n31544 );
or ( n37324 , n37322 , n37323 );
buf ( n37325 , n31478 );
nand ( n37326 , n37324 , n37325 );
buf ( n37327 , n37326 );
buf ( n37328 , n37327 );
nor ( n37329 , n37321 , n37328 );
buf ( n37330 , n37329 );
buf ( n37331 , n37330 );
buf ( n37332 , n37313 );
or ( n37333 , n37331 , n37332 );
buf ( n37334 , n37308 );
buf ( n37335 , n37310 );
nand ( n37336 , n37334 , n37335 );
buf ( n37337 , n37336 );
buf ( n37338 , n37337 );
nand ( n37339 , n37333 , n37338 );
buf ( n37340 , n37339 );
buf ( n37341 , n37340 );
nor ( n37342 , n37318 , n37341 );
buf ( n37343 , n37342 );
buf ( n37344 , n37343 );
not ( n37345 , n37344 );
or ( n37346 , n37293 , n37345 );
buf ( n37347 , n37343 );
buf ( n37348 , n37291 );
or ( n37349 , n37347 , n37348 );
nand ( n37350 , n37346 , n37349 );
buf ( n37351 , n37350 );
buf ( n37352 , n37351 );
nand ( n37353 , n22918 , n37352 );
buf ( n37354 , n37277 );
buf ( n37355 , n37354 );
buf ( n37356 , n13757 );
buf ( n37357 , n37356 );
nor ( n37358 , n37355 , n37357 );
buf ( n37359 , n37358 );
buf ( n37360 , n37359 );
buf ( n37361 , n37354 );
buf ( n37362 , n37356 );
and ( n37363 , n37361 , n37362 );
buf ( n37364 , n37363 );
buf ( n37365 , n37364 );
nor ( n37366 , n37360 , n37365 );
buf ( n37367 , n37366 );
buf ( n37368 , n37367 );
not ( n37369 , n37368 );
buf ( n37370 , n23365 );
buf ( n37371 , n31578 );
buf ( n37372 , n31606 );
nor ( n37373 , n37371 , n37372 );
buf ( n37374 , n37373 );
buf ( n37375 , n37374 );
buf ( n37376 , n31599 );
nand ( n37377 , n37375 , n37376 );
buf ( n37378 , n37377 );
buf ( n37379 , n37378 );
not ( n37380 , n37379 );
buf ( n37381 , n37380 );
buf ( n37382 , n37381 );
buf ( n37383 , n37307 );
buf ( n37384 , n37383 );
buf ( n37385 , n13779 );
buf ( n37386 , n37385 );
nor ( n37387 , n37384 , n37386 );
buf ( n37388 , n37387 );
buf ( n37389 , n37388 );
not ( n37390 , n37389 );
buf ( n37391 , n37390 );
buf ( n37392 , n37391 );
and ( n37393 , n37370 , n37382 , n37392 );
buf ( n37394 , n37374 );
buf ( n37395 , n31629 );
and ( n37396 , n37394 , n37395 );
buf ( n37397 , n31578 );
buf ( n37398 , n31636 );
or ( n37399 , n37397 , n37398 );
buf ( n37400 , n31572 );
nand ( n37401 , n37399 , n37400 );
buf ( n37402 , n37401 );
buf ( n37403 , n37402 );
nor ( n37404 , n37396 , n37403 );
buf ( n37405 , n37404 );
buf ( n37406 , n37405 );
buf ( n37407 , n37388 );
or ( n37408 , n37406 , n37407 );
buf ( n37409 , n37383 );
buf ( n37410 , n37385 );
nand ( n37411 , n37409 , n37410 );
buf ( n37412 , n37411 );
buf ( n37413 , n37412 );
nand ( n37414 , n37408 , n37413 );
buf ( n37415 , n37414 );
buf ( n37416 , n37415 );
nor ( n37417 , n37393 , n37416 );
buf ( n37418 , n37417 );
buf ( n37419 , n37418 );
not ( n37420 , n37419 );
or ( n37421 , n37369 , n37420 );
buf ( n37422 , n37418 );
buf ( n37423 , n37367 );
or ( n37424 , n37422 , n37423 );
nand ( n37425 , n37421 , n37424 );
buf ( n37426 , n37425 );
buf ( n37427 , n37426 );
nand ( n37428 , n23152 , n37427 );
nand ( n37429 , n37274 , n37276 , n37353 , n37428 );
buf ( n37430 , n37429 );
buf ( n37431 , n37430 );
not ( n37432 , n275550 );
buf ( n37433 , n37432 );
buf ( n37434 , n37433 );
and ( n37435 , n31306 , n35873 );
not ( n37436 , n20889 );
not ( n37437 , n31356 );
or ( n37438 , n37436 , n37437 );
and ( n37439 , n31320 , n20927 );
not ( n37440 , n17409 );
not ( n37441 , n31327 );
or ( n37442 , n37440 , n37441 );
nand ( n37443 , n20940 , n31332 );
nand ( n37444 , n37442 , n37443 );
nor ( n37445 , n37439 , n37444 );
nand ( n37446 , n37438 , n37445 );
nor ( n37447 , n37435 , n37446 );
or ( n37448 , n37447 , n27647 );
nand ( n37449 , n21696 , n13914 );
nand ( n37450 , n37448 , n37449 );
buf ( n37451 , n37450 );
buf ( n37452 , n37451 );
buf ( n37453 , n275554 );
not ( n37454 , n275929 );
buf ( n37455 , n37454 );
buf ( n37456 , n37455 );
buf ( n37457 , n275554 );
not ( n37458 , n275925 );
buf ( n37459 , n37458 );
buf ( n37460 , n37459 );
buf ( n37461 , n275554 );
or ( n37462 , n35069 , n27179 );
not ( n37463 , n27179 );
not ( n37464 , n277416 );
or ( n37465 , n37463 , n37464 );
nand ( n37466 , n37462 , n37465 );
buf ( n37467 , n37466 );
buf ( n37468 , n37467 );
not ( n37469 , n275550 );
buf ( n37470 , n37469 );
buf ( n37471 , n37470 );
not ( n37472 , n275550 );
buf ( n37473 , n37472 );
buf ( n37474 , n37473 );
not ( n37475 , n18189 );
not ( n37476 , n22335 );
or ( n37477 , n37475 , n37476 );
not ( n37478 , n29919 );
or ( n37479 , n37478 , n22335 );
nand ( n37480 , n37477 , n37479 );
buf ( n37481 , n37480 );
buf ( n37482 , n37481 );
buf ( n37483 , n275554 );
not ( n37484 , n31056 );
and ( n37485 , n37484 , n26638 );
not ( n37486 , n21001 );
not ( n37487 , n31122 );
or ( n37488 , n37486 , n37487 );
and ( n37489 , n31076 , n19358 );
not ( n37490 , n31098 );
not ( n37491 , n19219 );
or ( n37492 , n37490 , n37491 );
nand ( n37493 , n31094 , n19290 );
nand ( n37494 , n37492 , n37493 );
nor ( n37495 , n37489 , n37494 );
nand ( n37496 , n37488 , n37495 );
nor ( n37497 , n37485 , n37496 );
or ( n37498 , n37497 , n21030 );
nand ( n37499 , n21030 , n18825 );
nand ( n37500 , n37498 , n37499 );
buf ( n37501 , n37500 );
buf ( n37502 , n37501 );
not ( n37503 , n275929 );
buf ( n37504 , n37503 );
buf ( n37505 , n37504 );
not ( n37506 , n24050 );
or ( n37507 , n37506 , n22335 );
nand ( n37508 , n28818 , n22335 );
nand ( n37509 , n37507 , n37508 );
buf ( n37510 , n37509 );
buf ( n37511 , n37510 );
not ( n37512 , n275925 );
buf ( n37513 , n37512 );
buf ( n37514 , n37513 );
not ( n37515 , n16794 );
not ( n37516 , n23806 );
or ( n37517 , n37515 , n37516 );
buf ( n37518 , n22998 );
nand ( n37519 , n14830 , n37518 );
nand ( n37520 , n37517 , n37519 );
buf ( n37521 , n37520 );
buf ( n37522 , n37521 );
or ( n37523 , n23787 , n14909 );
and ( n37524 , n23759 , n17405 );
nand ( n37525 , n17411 , n23764 );
nand ( n37526 , n20785 , n23769 );
nand ( n37527 , n17562 , n13846 );
and ( n37528 , n17524 , n13856 );
not ( n37529 , n17524 );
not ( n37530 , n13855 );
and ( n37531 , n37529 , n37530 );
nor ( n37532 , n37528 , n37531 );
nand ( n37533 , n17545 , n37532 );
nand ( n37534 , n37525 , n37526 , n37527 , n37533 );
nor ( n37535 , n37524 , n37534 );
nand ( n37536 , n23729 , n16970 );
nand ( n37537 , n37523 , n37535 , n37536 );
buf ( n37538 , n37537 );
buf ( n37539 , n37538 );
buf ( n37540 , n275554 );
not ( n37541 , n275925 );
buf ( n37542 , n37541 );
buf ( n37543 , n37542 );
buf ( n37544 , n275554 );
buf ( n37545 , n275554 );
or ( n37546 , n33901 , n26364 );
nand ( n37547 , n33927 , n26370 );
nand ( n37548 , n33949 , n26374 );
not ( n37549 , n33958 );
not ( n37550 , n37549 );
not ( n37551 , n26390 );
and ( n37552 , n37550 , n37551 );
nand ( n37553 , n33968 , n32188 );
nand ( n37554 , n26395 , n24891 );
nand ( n37555 , n17542 , n14714 );
nand ( n37556 , n37553 , n37554 , n37555 );
nor ( n37557 , n37552 , n37556 );
and ( n37558 , n37547 , n37548 , n37557 );
nand ( n37559 , n37546 , n37558 );
buf ( n37560 , n37559 );
buf ( n37561 , n37560 );
and ( n37562 , n18208 , n35964 );
not ( n37563 , n18208 );
not ( n37564 , n23955 );
not ( n37565 , n37564 );
not ( n37566 , n21113 );
nor ( n37567 , n37566 , n21164 );
not ( n37568 , n37567 );
or ( n37569 , n37565 , n37568 );
or ( n37570 , n37567 , n37564 );
nand ( n37571 , n37569 , n37570 );
buf ( n37572 , n37571 );
and ( n37573 , n37563 , n37572 );
nor ( n37574 , n37562 , n37573 );
not ( n37575 , n37574 );
and ( n37576 , n37575 , n21174 );
not ( n37577 , n21001 );
not ( n37578 , n24175 );
nand ( n37579 , n37578 , n24196 );
not ( n37580 , n37579 );
not ( n37581 , n21363 );
nor ( n37582 , n37581 , n21469 );
not ( n37583 , n37582 );
nor ( n37584 , n37583 , n21417 );
not ( n37585 , n37584 );
not ( n37586 , n20337 );
or ( n37587 , n37585 , n37586 );
not ( n37588 , n37582 );
not ( n37589 , n21485 );
or ( n37590 , n37588 , n37589 );
not ( n37591 , n21491 );
not ( n37592 , n21362 );
and ( n37593 , n37591 , n37592 );
nor ( n37594 , n37593 , n21360 );
nand ( n37595 , n37590 , n37594 );
not ( n37596 , n37595 );
nand ( n37597 , n37587 , n37596 );
not ( n37598 , n37597 );
or ( n37599 , n37580 , n37598 );
or ( n37600 , n37597 , n37579 );
nand ( n37601 , n37599 , n37600 );
buf ( n37602 , n37601 );
not ( n37603 , n37602 );
or ( n37604 , n37577 , n37603 );
not ( n37605 , n24241 );
nand ( n37606 , n37605 , n24246 );
not ( n37607 , n37606 );
and ( n37608 , n21547 , n21515 );
not ( n37609 , n37608 );
nor ( n37610 , n37609 , n21563 );
not ( n37611 , n37610 );
not ( n37612 , n20500 );
or ( n37613 , n37611 , n37612 );
and ( n37614 , n37608 , n21576 );
not ( n37615 , n21515 );
not ( n37616 , n21585 );
or ( n37617 , n37615 , n37616 );
nand ( n37618 , n37617 , n21518 );
nor ( n37619 , n37614 , n37618 );
nand ( n37620 , n37613 , n37619 );
not ( n37621 , n37620 );
or ( n37622 , n37607 , n37621 );
or ( n37623 , n37620 , n37606 );
nand ( n37624 , n37622 , n37623 );
buf ( n37625 , n37624 );
and ( n37626 , n37625 , n19358 );
not ( n37627 , n19290 );
not ( n37628 , n24308 );
nand ( n37629 , n21611 , n21597 );
nor ( n37630 , n21605 , n37629 );
and ( n37631 , n37630 , n20547 );
not ( n37632 , n37631 );
or ( n37633 , n37628 , n37632 );
or ( n37634 , n37631 , n24308 );
nand ( n37635 , n37633 , n37634 );
buf ( n37636 , n37635 );
not ( n37637 , n37636 );
or ( n37638 , n37627 , n37637 );
buf ( n37639 , n24307 );
buf ( n37640 , n37639 );
buf ( n37641 , n37640 );
nand ( n37642 , n27619 , n37641 );
nand ( n37643 , n37638 , n37642 );
nor ( n37644 , n37626 , n37643 );
nand ( n37645 , n37604 , n37644 );
nor ( n37646 , n37576 , n37645 );
or ( n37647 , n37646 , n24450 );
nand ( n37648 , n24452 , n18692 );
nand ( n37649 , n37647 , n37648 );
buf ( n37650 , n37649 );
buf ( n37651 , n37650 );
not ( n37652 , n275929 );
buf ( n37653 , n37652 );
buf ( n37654 , n37653 );
or ( n37655 , n37646 , n21030 );
nand ( n37656 , n21030 , n18705 );
nand ( n37657 , n37655 , n37656 );
buf ( n37658 , n37657 );
buf ( n37659 , n37658 );
buf ( n37660 , n275554 );
not ( n37661 , n28304 );
and ( n37662 , n29153 , n37661 );
and ( n37663 , n29126 , n28328 );
nor ( n37664 , n37662 , n37663 );
not ( n37665 , n28218 );
and ( n37666 , n29138 , n37665 );
nor ( n37667 , n28241 , n12336 );
nor ( n37668 , n37666 , n37667 );
and ( n37669 , n31451 , n12264 );
not ( n37670 , n10752 );
or ( n37671 , n28233 , n37670 );
not ( n37672 , n10761 );
not ( n37673 , n37672 );
or ( n37674 , n28356 , n37673 );
nand ( n37675 , n37671 , n37674 );
nor ( n37676 , n37669 , n37675 );
nand ( n37677 , n37664 , n37668 , n37676 );
buf ( n37678 , n37677 );
buf ( n37679 , n37678 );
buf ( n37680 , n275554 );
not ( n37681 , n23088 );
not ( n37682 , n14830 );
or ( n37683 , n37681 , n37682 );
nand ( n37684 , n16321 , n23806 );
nand ( n37685 , n37683 , n37684 );
buf ( n37686 , n37685 );
buf ( n37687 , n37686 );
not ( n37688 , n275925 );
buf ( n37689 , n37688 );
buf ( n37690 , n37689 );
buf ( n37691 , n275554 );
not ( n37692 , n275550 );
buf ( n37693 , n37692 );
buf ( n37694 , n37693 );
buf ( n37695 , n275554 );
nand ( n37696 , n35012 , n31422 );
nand ( n37697 , n35037 , n31437 );
nand ( n37698 , n35044 , n31449 );
and ( n37699 , n32054 , n12198 );
not ( n37700 , n277625 );
not ( n37701 , n28357 );
or ( n37702 , n37700 , n37701 );
or ( n37703 , n32061 , n277614 );
nand ( n37704 , n37702 , n37703 );
nor ( n37705 , n37699 , n37704 );
nand ( n37706 , n31460 , n12365 );
and ( n37707 , n37698 , n37705 , n37706 );
nand ( n37708 , n37696 , n37697 , n37707 );
buf ( n37709 , n37708 );
buf ( n37710 , n37709 );
buf ( n37711 , n275554 );
not ( n37712 , n275550 );
buf ( n37713 , n37712 );
buf ( n37714 , n37713 );
not ( n37715 , n275550 );
buf ( n37716 , n37715 );
buf ( n37717 , n37716 );
not ( n37718 , n275929 );
buf ( n37719 , n37718 );
buf ( n37720 , n37719 );
not ( n37721 , n275550 );
buf ( n37722 , n37721 );
buf ( n37723 , n37722 );
buf ( n37724 , n275554 );
buf ( n37725 , n275554 );
buf ( n37726 , n275554 );
buf ( n37727 , n275554 );
and ( n37728 , n9158 , n9083 );
not ( n37729 , n9158 );
and ( n37730 , n37729 , n277531 );
or ( n37731 , n37728 , n37730 );
buf ( n37732 , n37731 );
buf ( n37733 , n37732 );
not ( n37734 , n275925 );
buf ( n37735 , n37734 );
buf ( n37736 , n37735 );
not ( n37737 , n275550 );
buf ( n37738 , n37737 );
buf ( n37739 , n37738 );
and ( n37740 , n37271 , n275648 );
nor ( n37741 , n14830 , n17512 );
nor ( n37742 , n37740 , n37741 );
nand ( n37743 , n22914 , n35488 );
buf ( n37744 , n23066 );
buf ( n37745 , n23109 );
and ( n37746 , n37744 , n37745 );
buf ( n37747 , n37746 );
buf ( n37748 , n37747 );
not ( n37749 , n37748 );
buf ( n37750 , n30540 );
buf ( n37751 , n23097 );
and ( n37752 , n37750 , n37751 );
buf ( n37753 , n23126 );
nor ( n37754 , n37752 , n37753 );
buf ( n37755 , n37754 );
buf ( n37756 , n37755 );
not ( n37757 , n37756 );
or ( n37758 , n37749 , n37757 );
buf ( n37759 , n37755 );
buf ( n37760 , n37747 );
or ( n37761 , n37759 , n37760 );
nand ( n37762 , n37758 , n37761 );
buf ( n37763 , n37762 );
buf ( n37764 , n37763 );
nand ( n37765 , n22918 , n37764 );
buf ( n37766 , n23294 );
buf ( n37767 , n23334 );
and ( n37768 , n37766 , n37767 );
buf ( n37769 , n37768 );
buf ( n37770 , n37769 );
not ( n37771 , n37770 );
buf ( n37772 , n30574 );
buf ( n37773 , n23322 );
and ( n37774 , n37772 , n37773 );
buf ( n37775 , n23351 );
nor ( n37776 , n37774 , n37775 );
buf ( n37777 , n37776 );
buf ( n37778 , n37777 );
not ( n37779 , n37778 );
or ( n37780 , n37771 , n37779 );
buf ( n37781 , n37777 );
buf ( n37782 , n37769 );
or ( n37783 , n37781 , n37782 );
nand ( n37784 , n37780 , n37783 );
buf ( n37785 , n37784 );
buf ( n37786 , n37785 );
nand ( n37787 , n23152 , n37786 );
nand ( n37788 , n37742 , n37743 , n37765 , n37787 );
buf ( n37789 , n37788 );
buf ( n37790 , n37789 );
nand ( n37791 , n34359 , n23603 );
nand ( n37792 , n34376 , n23655 );
and ( n37793 , n34383 , n29371 );
or ( n37794 , n22008 , n12352 );
or ( n37795 , n23680 , n34387 );
nand ( n37796 , n37794 , n37795 );
nor ( n37797 , n37793 , n37796 );
and ( n37798 , n37791 , n37792 , n37797 );
or ( n37799 , n37798 , n27179 );
nand ( n37800 , n23708 , n11256 );
nand ( n37801 , n37799 , n37800 );
buf ( n37802 , n37801 );
buf ( n37803 , n37802 );
not ( n37804 , n275550 );
buf ( n37805 , n37804 );
buf ( n37806 , n37805 );
and ( n37807 , n27589 , n10746 );
not ( n37808 , n27589 );
and ( n37809 , n37808 , n29155 );
or ( n37810 , n37807 , n37809 );
buf ( n37811 , n37810 );
buf ( n37812 , n37811 );
or ( n37813 , n23835 , n26365 );
nand ( n37814 , n23850 , n26370 );
nand ( n37815 , n23866 , n26374 );
not ( n37816 , n35740 );
nor ( n37817 , n37816 , n26390 );
nand ( n37818 , n23881 , n26393 );
nand ( n37819 , n26395 , n15557 );
nand ( n37820 , n17542 , n13949 );
nand ( n37821 , n37818 , n37819 , n37820 );
nor ( n37822 , n37817 , n37821 );
and ( n37823 , n37814 , n37815 , n37822 );
nand ( n37824 , n37813 , n37823 );
buf ( n37825 , n37824 );
buf ( n37826 , n37825 );
buf ( n37827 , n275554 );
buf ( n37828 , n275554 );
nand ( n37829 , n34811 , n29599 );
nand ( n37830 , n34837 , n30962 );
and ( n37831 , n34844 , n22052 );
or ( n37832 , n32722 , n12215 );
or ( n37833 , n22014 , n12166 );
nand ( n37834 , n37832 , n37833 );
nor ( n37835 , n37831 , n37834 );
and ( n37836 , n37829 , n37830 , n37835 );
or ( n37837 , n37836 , n27179 );
or ( n37838 , n37463 , n277560 );
nand ( n37839 , n37837 , n37838 );
buf ( n37840 , n37839 );
buf ( n37841 , n37840 );
not ( n37842 , n275550 );
buf ( n37843 , n37842 );
buf ( n37844 , n37843 );
not ( n37845 , n275929 );
buf ( n37846 , n37845 );
buf ( n37847 , n37846 );
or ( n37848 , n20985 , n19634 );
and ( n37849 , n34105 , n18324 );
nand ( n37850 , n20998 , n20353 );
nand ( n37851 , n19644 , n21022 );
nand ( n37852 , n21011 , n20515 );
nand ( n37853 , n19645 , n21018 );
nand ( n37854 , n37850 , n37851 , n37852 , n37853 );
nor ( n37855 , n37849 , n37854 );
nand ( n37856 , n37848 , n37855 );
buf ( n37857 , n37856 );
buf ( n37858 , n37857 );
buf ( n37859 , n275554 );
buf ( n37860 , n14599 );
and ( n37861 , n13373 , n37860 );
not ( n37862 , n13373 );
buf ( n37863 , n20829 );
and ( n37864 , n37863 , n20831 );
not ( n37865 , n37863 );
not ( n37866 , n20831 );
and ( n37867 , n37865 , n37866 );
nor ( n37868 , n37864 , n37867 );
buf ( n37869 , n37868 );
and ( n37870 , n37862 , n37869 );
nor ( n37871 , n37861 , n37870 );
or ( n37872 , n37871 , n14909 );
not ( n37873 , n16970 );
nand ( n37874 , n16498 , n16492 );
not ( n37875 , n37874 );
not ( n37876 , n16497 );
nor ( n37877 , n37876 , n16862 );
not ( n37878 , n37877 );
not ( n37879 , n32943 );
or ( n37880 , n37878 , n37879 );
not ( n37881 , n16497 );
not ( n37882 , n16874 );
or ( n37883 , n37881 , n37882 );
nand ( n37884 , n37883 , n16489 );
not ( n37885 , n37884 );
nand ( n37886 , n37880 , n37885 );
not ( n37887 , n37886 );
or ( n37888 , n37875 , n37887 );
or ( n37889 , n37886 , n37874 );
nand ( n37890 , n37888 , n37889 );
buf ( n37891 , n37890 );
not ( n37892 , n37891 );
or ( n37893 , n37873 , n37892 );
and ( n37894 , n17507 , n13574 );
not ( n37895 , n17507 );
not ( n37896 , n13573 );
and ( n37897 , n37895 , n37896 );
nor ( n37898 , n37894 , n37897 );
not ( n37899 , n37898 );
not ( n37900 , n17545 );
or ( n37901 , n37899 , n37900 );
not ( n37902 , n17417 );
not ( n37903 , n17415 );
and ( n37904 , n17433 , n37903 , n17421 );
not ( n37905 , n37904 );
or ( n37906 , n37902 , n37905 );
or ( n37907 , n37904 , n17417 );
nand ( n37908 , n37906 , n37907 );
buf ( n37909 , n37908 );
not ( n37910 , n37909 );
or ( n37911 , n17410 , n37910 );
nand ( n37912 , n37901 , n37911 );
buf ( n37913 , n17416 );
buf ( n37914 , n37913 );
buf ( n37915 , n37914 );
not ( n37916 , n37915 );
nor ( n37917 , n37916 , n17500 );
nor ( n37918 , n37912 , n37917 );
nand ( n37919 , n37893 , n37918 );
not ( n37920 , n17405 );
nor ( n37921 , n20896 , n17179 );
not ( n37922 , n37921 );
not ( n37923 , n32950 );
or ( n37924 , n37922 , n37923 );
not ( n37925 , n24698 );
not ( n37926 , n24702 );
or ( n37927 , n37925 , n37926 );
nand ( n37928 , n37927 , n24699 );
not ( n37929 , n37928 );
nand ( n37930 , n37924 , n37929 );
nand ( n37931 , n17159 , n17176 );
xnor ( n37932 , n37930 , n37931 );
buf ( n37933 , n37932 );
not ( n37934 , n37933 );
or ( n37935 , n37920 , n37934 );
nand ( n37936 , n17562 , n13571 );
nand ( n37937 , n37935 , n37936 );
nor ( n37938 , n37919 , n37937 );
nand ( n37939 , n37872 , n37938 );
buf ( n37940 , n37939 );
buf ( n37941 , n37940 );
not ( n37942 , n26551 );
or ( n37943 , n37942 , n21774 );
nand ( n37944 , n21770 , n9688 );
nand ( n37945 , n37943 , n37944 );
buf ( n37946 , n37945 );
buf ( n37947 , n37946 );
buf ( n37948 , n275554 );
buf ( n37949 , n275554 );
not ( n37950 , n275550 );
buf ( n37951 , n37950 );
buf ( n37952 , n37951 );
or ( n37953 , n31143 , n20742 );
nand ( n37954 , n31152 , n16970 );
nand ( n37955 , n31161 , n17405 );
not ( n37956 , n31169 );
not ( n37957 , n32339 );
or ( n37958 , n37956 , n37957 );
nand ( n37959 , n17545 , n31184 );
nand ( n37960 , n37958 , n37959 );
not ( n37961 , n31174 );
nor ( n37962 , n37961 , n17500 );
not ( n37963 , n13778 );
nor ( n37964 , n17561 , n37963 );
nor ( n37965 , n37960 , n37962 , n37964 );
and ( n37966 , n37954 , n37955 , n37965 );
nand ( n37967 , n37953 , n37966 );
buf ( n37968 , n37967 );
buf ( n37969 , n37968 );
not ( n37970 , n275925 );
buf ( n37971 , n37970 );
buf ( n37972 , n37971 );
not ( n37973 , n23774 );
or ( n37974 , n37973 , n29044 );
nand ( n37975 , n28252 , n9720 );
nand ( n37976 , n37974 , n37975 );
buf ( n37977 , n37976 );
buf ( n37978 , n37977 );
not ( n37979 , n275550 );
buf ( n37980 , n37979 );
buf ( n37981 , n37980 );
not ( n37982 , n275550 );
buf ( n37983 , n37982 );
buf ( n37984 , n37983 );
nand ( n37985 , n32811 , n33491 );
or ( n37986 , n37985 , n31448 );
and ( n37987 , n28350 , n277498 );
or ( n37988 , n28233 , n9396 );
nand ( n37989 , n37988 , n33500 );
nor ( n37990 , n37987 , n37989 );
nand ( n37991 , n37986 , n37990 );
buf ( n37992 , n37991 );
buf ( n37993 , n37992 );
buf ( n37994 , n275554 );
buf ( n37995 , n275554 );
not ( n37996 , n275550 );
buf ( n37997 , n37996 );
buf ( n37998 , n37997 );
not ( n37999 , n275550 );
buf ( n38000 , n37999 );
buf ( n38001 , n38000 );
buf ( n38002 , n275554 );
buf ( n38003 , n275554 );
not ( n38004 , n275929 );
buf ( n38005 , n38004 );
buf ( n38006 , n38005 );
not ( n38007 , n17965 );
not ( n38008 , n22335 );
or ( n38009 , n38007 , n38008 );
not ( n38010 , n27995 );
or ( n38011 , n38010 , n22335 );
nand ( n38012 , n38009 , n38011 );
buf ( n38013 , n38012 );
buf ( n38014 , n38013 );
not ( n38015 , n275929 );
buf ( n38016 , n38015 );
buf ( n38017 , n38016 );
buf ( n38018 , n275554 );
buf ( n38019 , n275554 );
buf ( n38020 , n275554 );
not ( n38021 , n275550 );
buf ( n38022 , n38021 );
buf ( n38023 , n38022 );
buf ( n38024 , n275554 );
not ( n38025 , n275549 );
not ( n38026 , n38025 );
buf ( n38027 , n38026 );
buf ( n38028 , n38027 );
buf ( n38029 , n275554 );
not ( n38030 , n275550 );
buf ( n38031 , n38030 );
buf ( n38032 , n38031 );
not ( n38033 , n27685 );
or ( n38034 , n38033 , n29046 );
nand ( n38035 , n28252 , n9531 );
nand ( n38036 , n38034 , n38035 );
buf ( n38037 , n38036 );
buf ( n38038 , n38037 );
buf ( n38039 , n275554 );
not ( n38040 , n275550 );
buf ( n38041 , n38040 );
buf ( n38042 , n38041 );
and ( n38043 , n26516 , n27810 );
not ( n38044 , n26516 );
not ( n38045 , n29857 );
not ( n38046 , n38045 );
not ( n38047 , n34165 );
or ( n38048 , n38046 , n38047 );
or ( n38049 , n38045 , n34165 );
nand ( n38050 , n38048 , n38049 );
buf ( n38051 , n38050 );
and ( n38052 , n38044 , n38051 );
nor ( n38053 , n38043 , n38052 );
or ( n38054 , n38053 , n19216 );
nand ( n38055 , n30024 , n30060 );
not ( n38056 , n38055 );
not ( n38057 , n30038 );
nand ( n38058 , n38057 , n30035 );
nor ( n38059 , n28014 , n38058 );
not ( n38060 , n38059 );
not ( n38061 , n30043 );
or ( n38062 , n38060 , n38061 );
not ( n38063 , n28037 );
not ( n38064 , n38058 );
and ( n38065 , n38063 , n38064 );
not ( n38066 , n30035 );
not ( n38067 , n30052 );
or ( n38068 , n38066 , n38067 );
nand ( n38069 , n38068 , n30057 );
nor ( n38070 , n38065 , n38069 );
nand ( n38071 , n38062 , n38070 );
not ( n38072 , n38071 );
or ( n38073 , n38056 , n38072 );
or ( n38074 , n38071 , n38055 );
nand ( n38075 , n38073 , n38074 );
buf ( n38076 , n38075 );
nand ( n38077 , n38076 , n33157 );
or ( n38078 , n30090 , n30120 );
not ( n38079 , n38078 );
nor ( n38080 , n35437 , n30099 );
not ( n38081 , n38080 );
nor ( n38082 , n38081 , n28079 );
not ( n38083 , n38082 );
not ( n38084 , n28092 );
or ( n38085 , n38083 , n38084 );
not ( n38086 , n38080 );
not ( n38087 , n28109 );
or ( n38088 , n38086 , n38087 );
not ( n38089 , n35434 );
not ( n38090 , n30113 );
or ( n38091 , n38089 , n38090 );
nand ( n38092 , n38091 , n30117 );
not ( n38093 , n38092 );
nand ( n38094 , n38088 , n38093 );
not ( n38095 , n38094 );
nand ( n38096 , n38085 , n38095 );
not ( n38097 , n38096 );
or ( n38098 , n38079 , n38097 );
or ( n38099 , n38096 , n38078 );
nand ( n38100 , n38098 , n38099 );
buf ( n38101 , n38100 );
nand ( n38102 , n38101 , n19360 );
not ( n38103 , n18507 );
and ( n38104 , n30148 , n38103 );
not ( n38105 , n30148 );
and ( n38106 , n38105 , n18508 );
nor ( n38107 , n38104 , n38106 );
not ( n38108 , n38107 );
nand ( n38109 , n38108 , n19318 );
not ( n38110 , n30163 );
not ( n38111 , n30158 );
nor ( n38112 , n27062 , n24300 , n28126 );
nor ( n38113 , n27059 , n28122 , n30162 );
nand ( n38114 , n38111 , n28125 , n38112 , n38113 );
nor ( n38115 , n28124 , n38114 );
not ( n38116 , n38115 );
or ( n38117 , n38110 , n38116 );
or ( n38118 , n38115 , n30163 );
nand ( n38119 , n38117 , n38118 );
buf ( n38120 , n38119 );
nand ( n38121 , n38120 , n29075 );
buf ( n38122 , n30076 );
buf ( n38123 , n38122 );
buf ( n38124 , n38123 );
buf ( n38125 , n38124 );
nand ( n38126 , n33162 , n38125 );
nand ( n38127 , n19387 , n18504 );
and ( n38128 , n38109 , n38121 , n38126 , n38127 );
and ( n38129 , n38077 , n38102 , n38128 );
nand ( n38130 , n38054 , n38129 );
buf ( n38131 , n38130 );
buf ( n38132 , n38131 );
and ( n38133 , n32940 , n21659 );
not ( n38134 , n20889 );
not ( n38135 , n32948 );
or ( n38136 , n38134 , n38135 );
and ( n38137 , n32955 , n20927 );
not ( n38138 , n17409 );
not ( n38139 , n32965 );
or ( n38140 , n38138 , n38139 );
not ( n38141 , n32958 );
or ( n38142 , n20939 , n38141 );
nand ( n38143 , n38140 , n38142 );
nor ( n38144 , n38137 , n38143 );
nand ( n38145 , n38136 , n38144 );
nor ( n38146 , n38133 , n38145 );
or ( n38147 , n38146 , n21697 );
nand ( n38148 , n21696 , n13649 );
nand ( n38149 , n38147 , n38148 );
buf ( n38150 , n38149 );
buf ( n38151 , n38150 );
not ( n38152 , n275929 );
buf ( n38153 , n38152 );
buf ( n38154 , n38153 );
or ( n38155 , n33544 , n21030 );
nand ( n38156 , n21030 , n18289 );
nand ( n38157 , n38155 , n38156 );
buf ( n38158 , n38157 );
buf ( n38159 , n38158 );
not ( n38160 , n275550 );
buf ( n38161 , n38160 );
buf ( n38162 , n38161 );
and ( n38163 , n37271 , n9413 );
nor ( n38164 , n38163 , n32316 );
nand ( n38165 , n22914 , n14880 );
buf ( n38166 , n14880 );
buf ( n38167 , n38166 );
buf ( n38168 , n38167 );
not ( n38169 , n38168 );
buf ( n38170 , n13888 );
buf ( n38171 , n38170 );
not ( n38172 , n38171 );
and ( n38173 , n38169 , n38172 );
buf ( n38174 , n38167 );
buf ( n38175 , n38170 );
and ( n38176 , n38174 , n38175 );
nor ( n38177 , n38173 , n38176 );
buf ( n38178 , n38177 );
buf ( n38179 , n38178 );
not ( n38180 , n38179 );
buf ( n38181 , n23140 );
buf ( n38182 , n37305 );
buf ( n38183 , n37283 );
buf ( n38184 , n37313 );
or ( n38185 , n38183 , n38184 );
buf ( n38186 , n38185 );
buf ( n38187 , n38186 );
buf ( n38188 , n12882 );
buf ( n38189 , n38188 );
buf ( n38190 , n38189 );
buf ( n38191 , n38190 );
buf ( n38192 , n13849 );
buf ( n38193 , n38192 );
nor ( n38194 , n38191 , n38193 );
buf ( n38195 , n38194 );
buf ( n38196 , n38195 );
nor ( n38197 , n38187 , n38196 );
buf ( n38198 , n38197 );
buf ( n38199 , n38198 );
and ( n38200 , n38181 , n38182 , n38199 );
buf ( n38201 , n37330 );
buf ( n38202 , n38198 );
not ( n38203 , n38202 );
buf ( n38204 , n38203 );
buf ( n38205 , n38204 );
or ( n38206 , n38201 , n38205 );
buf ( n38207 , n38195 );
buf ( n38208 , n37283 );
not ( n38209 , n38208 );
buf ( n38210 , n37337 );
not ( n38211 , n38210 );
and ( n38212 , n38209 , n38211 );
buf ( n38213 , n37288 );
nor ( n38214 , n38212 , n38213 );
buf ( n38215 , n38214 );
buf ( n38216 , n38215 );
or ( n38217 , n38207 , n38216 );
buf ( n38218 , n38190 );
buf ( n38219 , n38192 );
nand ( n38220 , n38218 , n38219 );
buf ( n38221 , n38220 );
buf ( n38222 , n38221 );
nand ( n38223 , n38206 , n38217 , n38222 );
buf ( n38224 , n38223 );
buf ( n38225 , n38224 );
nor ( n38226 , n38200 , n38225 );
buf ( n38227 , n38226 );
buf ( n38228 , n38227 );
not ( n38229 , n38228 );
or ( n38230 , n38180 , n38229 );
buf ( n38231 , n38227 );
buf ( n38232 , n38178 );
or ( n38233 , n38231 , n38232 );
nand ( n38234 , n38230 , n38233 );
buf ( n38235 , n38234 );
buf ( n38236 , n38235 );
nand ( n38237 , n22918 , n38236 );
buf ( n38238 , n38166 );
buf ( n38239 , n38238 );
not ( n38240 , n38239 );
buf ( n38241 , n13893 );
buf ( n38242 , n38241 );
not ( n38243 , n38242 );
and ( n38244 , n38240 , n38243 );
buf ( n38245 , n38238 );
buf ( n38246 , n38241 );
and ( n38247 , n38245 , n38246 );
nor ( n38248 , n38244 , n38247 );
buf ( n38249 , n38248 );
buf ( n38250 , n38249 );
not ( n38251 , n38250 );
buf ( n38252 , n23365 );
buf ( n38253 , n37381 );
buf ( n38254 , n37359 );
buf ( n38255 , n37388 );
or ( n38256 , n38254 , n38255 );
buf ( n38257 , n38256 );
buf ( n38258 , n38257 );
buf ( n38259 , n38189 );
buf ( n38260 , n38259 );
buf ( n38261 , n13846 );
buf ( n38262 , n38261 );
nor ( n38263 , n38260 , n38262 );
buf ( n38264 , n38263 );
buf ( n38265 , n38264 );
nor ( n38266 , n38258 , n38265 );
buf ( n38267 , n38266 );
buf ( n38268 , n38267 );
and ( n38269 , n38252 , n38253 , n38268 );
buf ( n38270 , n37405 );
buf ( n38271 , n38267 );
not ( n38272 , n38271 );
buf ( n38273 , n38272 );
buf ( n38274 , n38273 );
or ( n38275 , n38270 , n38274 );
buf ( n38276 , n38264 );
buf ( n38277 , n37359 );
not ( n38278 , n38277 );
buf ( n38279 , n37412 );
not ( n38280 , n38279 );
and ( n38281 , n38278 , n38280 );
buf ( n38282 , n37364 );
nor ( n38283 , n38281 , n38282 );
buf ( n38284 , n38283 );
buf ( n38285 , n38284 );
or ( n38286 , n38276 , n38285 );
buf ( n38287 , n38259 );
buf ( n38288 , n38261 );
nand ( n38289 , n38287 , n38288 );
buf ( n38290 , n38289 );
buf ( n38291 , n38290 );
nand ( n38292 , n38275 , n38286 , n38291 );
buf ( n38293 , n38292 );
buf ( n38294 , n38293 );
nor ( n38295 , n38269 , n38294 );
buf ( n38296 , n38295 );
buf ( n38297 , n38296 );
not ( n38298 , n38297 );
or ( n38299 , n38251 , n38298 );
buf ( n38300 , n38296 );
buf ( n38301 , n38249 );
or ( n38302 , n38300 , n38301 );
nand ( n38303 , n38299 , n38302 );
buf ( n38304 , n38303 );
buf ( n38305 , n38304 );
nand ( n38306 , n23152 , n38305 );
nand ( n38307 , n38164 , n38165 , n38237 , n38306 );
buf ( n38308 , n38307 );
buf ( n38309 , n38308 );
not ( n38310 , n275925 );
buf ( n38311 , n38310 );
buf ( n38312 , n38311 );
not ( n38313 , n275550 );
buf ( n38314 , n38313 );
buf ( n38315 , n38314 );
not ( n38316 , n275550 );
buf ( n38317 , n38316 );
buf ( n38318 , n38317 );
not ( n38319 , n275925 );
buf ( n38320 , n38319 );
buf ( n38321 , n38320 );
not ( n38322 , n275929 );
buf ( n38323 , n38322 );
buf ( n38324 , n38323 );
not ( n38325 , n275550 );
buf ( n38326 , n38325 );
buf ( n38327 , n38326 );
not ( n38328 , n32131 );
or ( n38329 , n38328 , n29044 );
nand ( n38330 , n29044 , n9548 );
nand ( n38331 , n38329 , n38330 );
buf ( n38332 , n38331 );
buf ( n38333 , n38332 );
or ( n38334 , n24494 , n26364 );
nand ( n38335 , n24574 , n26370 );
nand ( n38336 , n24607 , n26374 );
and ( n38337 , n33951 , n33952 );
not ( n38338 , n33951 );
and ( n38339 , n38338 , n14034 );
nor ( n38340 , n38337 , n38339 );
not ( n38341 , n38340 );
nor ( n38342 , n38341 , n26390 );
nand ( n38343 , n24617 , n32188 );
nand ( n38344 , n26395 , n24538 );
nand ( n38345 , n17542 , n14034 );
nand ( n38346 , n38343 , n38344 , n38345 );
nor ( n38347 , n38342 , n38346 );
and ( n38348 , n38335 , n38336 , n38347 );
nand ( n38349 , n38334 , n38348 );
buf ( n38350 , n38349 );
buf ( n38351 , n38350 );
or ( n38352 , n29517 , n19636 );
not ( n38353 , n30612 );
not ( n38354 , n38353 );
not ( n38355 , n29543 );
and ( n38356 , n38354 , n38355 );
and ( n38357 , n29579 , n20353 );
nor ( n38358 , n38356 , n38357 );
and ( n38359 , n29535 , n20515 );
not ( n38360 , n35321 );
nand ( n38361 , n29557 , n20560 );
nand ( n38362 , n19644 , n29548 );
nand ( n38363 , n38360 , n38361 , n38362 );
nor ( n38364 , n38359 , n38363 );
and ( n38365 , n38358 , n38364 );
nand ( n38366 , n38352 , n38365 );
buf ( n38367 , n38366 );
buf ( n38368 , n38367 );
not ( n38369 , n16012 );
or ( n38370 , n38369 , n23807 );
or ( n38371 , n17542 , n14890 );
nand ( n38372 , n38370 , n38371 );
buf ( n38373 , n38372 );
buf ( n38374 , n38373 );
buf ( n38375 , n275554 );
and ( n38376 , n33796 , n20987 );
not ( n38377 , n21001 );
not ( n38378 , n33805 );
or ( n38379 , n38377 , n38378 );
and ( n38380 , n33817 , n19358 );
not ( n38381 , n19290 );
not ( n38382 , n33826 );
or ( n38383 , n38381 , n38382 );
nand ( n38384 , n19219 , n33837 );
nand ( n38385 , n38383 , n38384 );
nor ( n38386 , n38380 , n38385 );
nand ( n38387 , n38379 , n38386 );
nor ( n38388 , n38376 , n38387 );
or ( n38389 , n38388 , n24452 );
nand ( n38390 , n24450 , n18953 );
nand ( n38391 , n38389 , n38390 );
buf ( n38392 , n38391 );
buf ( n38393 , n38392 );
or ( n38394 , n29464 , n24450 );
nand ( n38395 , n24452 , n19015 );
nand ( n38396 , n38394 , n38395 );
buf ( n38397 , n38396 );
buf ( n38398 , n38397 );
not ( n38399 , n15725 );
or ( n38400 , n38399 , n14830 );
nand ( n38401 , n14830 , n37275 );
nand ( n38402 , n38400 , n38401 );
buf ( n38403 , n38402 );
buf ( n38404 , n38403 );
or ( n38405 , n14806 , n26364 );
nand ( n38406 , n16954 , n26370 );
nand ( n38407 , n17401 , n26374 );
not ( n38408 , n17539 );
nor ( n38409 , n38408 , n26390 );
nand ( n38410 , n17496 , n32188 );
nand ( n38411 , n26395 , n15509 );
nand ( n38412 , n17542 , n14002 );
nand ( n38413 , n38410 , n38411 , n38412 );
nor ( n38414 , n38409 , n38413 );
and ( n38415 , n38406 , n38407 , n38414 );
nand ( n38416 , n38405 , n38415 );
buf ( n38417 , n38416 );
buf ( n38418 , n38417 );
nand ( n38419 , n25064 , n25119 );
buf ( n38420 , n25125 );
not ( n38421 , n38420 );
buf ( n38422 , n25316 );
nand ( n38423 , n38421 , n38422 );
buf ( n38424 , n38423 );
buf ( n38425 , n38424 );
not ( n38426 , n38425 );
buf ( n38427 , n25264 );
not ( n38428 , n38427 );
or ( n38429 , n38426 , n38428 );
buf ( n38430 , n25264 );
buf ( n38431 , n38424 );
or ( n38432 , n38430 , n38431 );
nand ( n38433 , n38429 , n38432 );
buf ( n38434 , n38433 );
buf ( n38435 , n38434 );
not ( n38436 , n38435 );
nor ( n38437 , n38436 , n25389 );
nand ( n38438 , n25397 , n275614 );
buf ( n38439 , n25450 );
not ( n38440 , n38439 );
buf ( n38441 , n25629 );
nand ( n38442 , n38440 , n38441 );
buf ( n38443 , n38442 );
buf ( n38444 , n38443 );
not ( n38445 , n38444 );
buf ( n38446 , n25586 );
not ( n38447 , n38446 );
or ( n38448 , n38445 , n38447 );
buf ( n38449 , n25586 );
buf ( n38450 , n38443 );
or ( n38451 , n38449 , n38450 );
nand ( n38452 , n38448 , n38451 );
buf ( n38453 , n38452 );
buf ( n38454 , n38453 );
and ( n38455 , n25402 , n38454 );
not ( n38456 , n18345 );
nor ( n38457 , n38456 , n19639 );
nor ( n38458 , n38455 , n38457 );
buf ( n38459 , n25767 );
not ( n38460 , n38459 );
buf ( n38461 , n25943 );
nand ( n38462 , n38460 , n38461 );
buf ( n38463 , n38462 );
buf ( n38464 , n38463 );
not ( n38465 , n38464 );
buf ( n38466 , n25902 );
not ( n38467 , n38466 );
or ( n38468 , n38465 , n38467 );
buf ( n38469 , n25902 );
buf ( n38470 , n38463 );
or ( n38471 , n38469 , n38470 );
nand ( n38472 , n38468 , n38471 );
buf ( n38473 , n38472 );
buf ( n38474 , n38473 );
nand ( n38475 , n28761 , n38474 );
nand ( n38476 , n38438 , n38458 , n38475 );
nor ( n38477 , n38437 , n38476 );
buf ( n38478 , n26075 );
not ( n38479 , n38478 );
buf ( n38480 , n26261 );
nand ( n38481 , n38479 , n38480 );
buf ( n38482 , n38481 );
buf ( n38483 , n38482 );
not ( n38484 , n38483 );
buf ( n38485 , n26212 );
not ( n38486 , n38485 );
or ( n38487 , n38484 , n38486 );
buf ( n38488 , n26212 );
buf ( n38489 , n38482 );
or ( n38490 , n38488 , n38489 );
nand ( n38491 , n38487 , n38490 );
buf ( n38492 , n38491 );
buf ( n38493 , n38492 );
nand ( n38494 , n26027 , n38493 );
nand ( n38495 , n38419 , n38477 , n38494 );
buf ( n38496 , n38495 );
buf ( n38497 , n38496 );
buf ( n38498 , n275554 );
not ( n38499 , n275550 );
buf ( n38500 , n38499 );
buf ( n38501 , n38500 );
not ( n38502 , n38053 );
and ( n38503 , n38502 , n26638 );
not ( n38504 , n21001 );
not ( n38505 , n38076 );
or ( n38506 , n38504 , n38505 );
and ( n38507 , n38101 , n19358 );
not ( n38508 , n38125 );
not ( n38509 , n27619 );
or ( n38510 , n38508 , n38509 );
nand ( n38511 , n38120 , n19290 );
nand ( n38512 , n38510 , n38511 );
nor ( n38513 , n38507 , n38512 );
nand ( n38514 , n38506 , n38513 );
nor ( n38515 , n38503 , n38514 );
or ( n38516 , n38515 , n35473 );
nand ( n38517 , n28146 , n18513 );
nand ( n38518 , n38516 , n38517 );
buf ( n38519 , n38518 );
buf ( n38520 , n38519 );
not ( n38521 , n275925 );
buf ( n38522 , n38521 );
buf ( n38523 , n38522 );
not ( n38524 , n32617 );
or ( n38525 , n38524 , n28252 );
nand ( n38526 , n28252 , n9692 );
nand ( n38527 , n38525 , n38526 );
buf ( n38528 , n38527 );
buf ( n38529 , n38528 );
not ( n38530 , n35814 );
and ( n38531 , n38530 , n23992 );
not ( n38532 , n21001 );
not ( n38533 , n35862 );
or ( n38534 , n38532 , n38533 );
and ( n38535 , n35826 , n19358 );
not ( n38536 , n19290 );
not ( n38537 , n35847 );
or ( n38538 , n38536 , n38537 );
nand ( n38539 , n19219 , n35837 );
nand ( n38540 , n38538 , n38539 );
nor ( n38541 , n38535 , n38540 );
nand ( n38542 , n38534 , n38541 );
nor ( n38543 , n38531 , n38542 );
or ( n38544 , n38543 , n21030 );
nand ( n38545 , n21030 , n18405 );
nand ( n38546 , n38544 , n38545 );
buf ( n38547 , n38546 );
buf ( n38548 , n38547 );
not ( n38549 , n275925 );
buf ( n38550 , n38549 );
buf ( n38551 , n38550 );
buf ( n38552 , n275554 );
buf ( n38553 , n275554 );
buf ( n38554 , n275554 );
buf ( n38555 , n275554 );
not ( n38556 , n275929 );
buf ( n38557 , n38556 );
buf ( n38558 , n38557 );
not ( n38559 , n27098 );
or ( n38560 , n38559 , n29046 );
nand ( n38561 , n29044 , n9566 );
nand ( n38562 , n38560 , n38561 );
buf ( n38563 , n38562 );
buf ( n38564 , n38563 );
not ( n38565 , n26626 );
not ( n38566 , n38565 );
not ( n38567 , n38566 );
or ( n38568 , n38567 , n21770 );
nand ( n38569 , n21774 , n9706 );
nand ( n38570 , n38568 , n38569 );
buf ( n38571 , n38570 );
buf ( n38572 , n38571 );
buf ( n38573 , n275554 );
not ( n38574 , n275798 );
nand ( n38575 , n38574 , n275839 );
not ( n38576 , n38575 );
not ( n38577 , n35767 );
not ( n38578 , n275767 );
or ( n38579 , n38577 , n38578 );
nand ( n38580 , n38579 , n275837 );
not ( n38581 , n38580 );
or ( n38582 , n38576 , n38581 );
or ( n38583 , n38580 , n38575 );
nand ( n38584 , n38582 , n38583 );
buf ( n38585 , n38584 );
buf ( n38586 , n38585 );
not ( n38587 , n277948 );
not ( n38588 , n27179 );
or ( n38589 , n38587 , n38588 );
not ( n38590 , n31734 );
or ( n38591 , n38590 , n27179 );
nand ( n38592 , n38589 , n38591 );
buf ( n38593 , n38592 );
buf ( n38594 , n38593 );
nand ( n38595 , n30448 , n28306 );
nand ( n38596 , n30472 , n28330 );
and ( n38597 , n28332 , n30488 );
and ( n38598 , n28350 , n12153 );
nor ( n38599 , n38597 , n38598 );
and ( n38600 , n28231 , n12207 );
or ( n38601 , n28354 , n11274 );
nand ( n38602 , n28357 , n11283 );
nand ( n38603 , n38601 , n38602 );
nor ( n38604 , n38600 , n38603 );
nand ( n38605 , n38595 , n38596 , n38599 , n38604 );
buf ( n38606 , n38605 );
buf ( n38607 , n38606 );
not ( n38608 , n16608 );
or ( n38609 , n38608 , n14830 );
nand ( n38610 , n31496 , n23807 );
nand ( n38611 , n38609 , n38610 );
buf ( n38612 , n38611 );
buf ( n38613 , n38612 );
not ( n38614 , n275550 );
buf ( n38615 , n38614 );
buf ( n38616 , n38615 );
buf ( n38617 , n275554 );
not ( n38618 , n275550 );
buf ( n38619 , n38618 );
buf ( n38620 , n38619 );
not ( n38621 , n24485 );
or ( n38622 , n38621 , n29046 );
nand ( n38623 , n28252 , n9740 );
nand ( n38624 , n38622 , n38623 );
buf ( n38625 , n38624 );
buf ( n38626 , n38625 );
not ( n38627 , n275929 );
buf ( n38628 , n38627 );
buf ( n38629 , n38628 );
not ( n38630 , n275550 );
buf ( n38631 , n38630 );
buf ( n38632 , n38631 );
buf ( n38633 , n275554 );
buf ( n38634 , n275554 );
not ( n38635 , n275929 );
buf ( n38636 , n38635 );
buf ( n38637 , n38636 );
buf ( n38638 , n275554 );
not ( n38639 , n275925 );
buf ( n38640 , n38639 );
buf ( n38641 , n38640 );
not ( n38642 , n275925 );
buf ( n38643 , n38642 );
buf ( n38644 , n38643 );
not ( n38645 , n275929 );
buf ( n38646 , n38645 );
buf ( n38647 , n38646 );
not ( n38648 , n18314 );
not ( n38649 , n24450 );
or ( n38650 , n38648 , n38649 );
or ( n38651 , n21026 , n24450 );
nand ( n38652 , n38650 , n38651 );
buf ( n38653 , n38652 );
buf ( n38654 , n38653 );
not ( n38655 , n26103 );
not ( n38656 , n22335 );
or ( n38657 , n38655 , n38656 );
nand ( n38658 , n20181 , n275557 );
nand ( n38659 , n38657 , n38658 );
buf ( n38660 , n38659 );
buf ( n38661 , n38660 );
not ( n38662 , n275929 );
buf ( n38663 , n38662 );
buf ( n38664 , n38663 );
not ( n38665 , n275929 );
buf ( n38666 , n38665 );
buf ( n38667 , n38666 );
not ( n38668 , n275925 );
buf ( n38669 , n38668 );
buf ( n38670 , n38669 );
not ( n38671 , n275929 );
buf ( n38672 , n38671 );
buf ( n38673 , n38672 );
or ( n38674 , n32699 , n23887 );
nand ( n38675 , n20951 , n13809 );
nand ( n38676 , n38674 , n38675 );
buf ( n38677 , n38676 );
buf ( n38678 , n38677 );
buf ( n38679 , n275554 );
not ( n38680 , n14841 );
not ( n38681 , n14896 );
and ( n38682 , n38680 , n38681 );
nor ( n38683 , n38682 , n14838 );
not ( n38684 , n24834 );
or ( n38685 , n38683 , n38684 );
nand ( n38686 , n38685 , n14830 );
buf ( n38687 , n38686 );
buf ( n38688 , n38687 );
buf ( n38689 , n275554 );
buf ( n38690 , n275554 );
buf ( n38691 , n275554 );
not ( n38692 , n275550 );
buf ( n38693 , n38692 );
buf ( n38694 , n38693 );
and ( n38695 , n23907 , n38566 );
not ( n38696 , n23907 );
not ( n38697 , n21140 );
nand ( n38698 , n38697 , n21163 , n21113 );
not ( n38699 , n38698 );
nand ( n38700 , n33060 , n23955 );
nor ( n38701 , n33067 , n38700 , n23980 );
nand ( n38702 , n38699 , n38701 , n19069 );
buf ( n38703 , n26628 );
xnor ( n38704 , n38702 , n38703 );
buf ( n38705 , n38704 );
and ( n38706 , n38696 , n38705 );
or ( n38707 , n38695 , n38706 );
and ( n38708 , n38707 , n27845 );
not ( n38709 , n21001 );
nand ( n38710 , n26911 , n26931 );
not ( n38711 , n38710 );
not ( n38712 , n26852 );
not ( n38713 , n24204 );
or ( n38714 , n38712 , n38713 );
not ( n38715 , n26928 );
nand ( n38716 , n38714 , n38715 );
not ( n38717 , n38716 );
or ( n38718 , n38711 , n38717 );
or ( n38719 , n38716 , n38710 );
nand ( n38720 , n38718 , n38719 );
buf ( n38721 , n38720 );
not ( n38722 , n38721 );
or ( n38723 , n38709 , n38722 );
nand ( n38724 , n31065 , n27036 );
not ( n38725 , n38724 );
not ( n38726 , n26990 );
not ( n38727 , n27020 );
or ( n38728 , n38726 , n38727 );
not ( n38729 , n27034 );
nand ( n38730 , n38728 , n38729 );
not ( n38731 , n38730 );
or ( n38732 , n38725 , n38731 );
or ( n38733 , n38730 , n38724 );
nand ( n38734 , n38732 , n38733 );
buf ( n38735 , n38734 );
and ( n38736 , n38735 , n19358 );
buf ( n38737 , n27069 );
buf ( n38738 , n38737 );
buf ( n38739 , n38738 );
not ( n38740 , n38739 );
not ( n38741 , n19219 );
or ( n38742 , n38740 , n38741 );
not ( n38743 , n27071 );
not ( n38744 , n27065 );
nand ( n38745 , n38744 , n24314 );
not ( n38746 , n38745 );
or ( n38747 , n38743 , n38746 );
or ( n38748 , n38745 , n27071 );
nand ( n38749 , n38747 , n38748 );
buf ( n38750 , n38749 );
nand ( n38751 , n38750 , n19290 );
nand ( n38752 , n38742 , n38751 );
nor ( n38753 , n38736 , n38752 );
nand ( n38754 , n38723 , n38753 );
nor ( n38755 , n38708 , n38754 );
or ( n38756 , n38755 , n28146 );
nand ( n38757 , n24450 , n18663 );
nand ( n38758 , n38756 , n38757 );
buf ( n38759 , n38758 );
buf ( n38760 , n38759 );
buf ( n38761 , n275554 );
buf ( n38762 , n275554 );
not ( n38763 , n16842 );
not ( n38764 , n23806 );
or ( n38765 , n38763 , n38764 );
nand ( n38766 , n14830 , n22969 );
nand ( n38767 , n38765 , n38766 );
buf ( n38768 , n38767 );
buf ( n38769 , n38768 );
not ( n38770 , n275929 );
buf ( n38771 , n38770 );
buf ( n38772 , n38771 );
buf ( n38773 , n275554 );
buf ( n38774 , n275554 );
and ( n38775 , n17562 , n14742 );
not ( n38776 , n17562 );
buf ( n38777 , n277460 );
buf ( n38778 , n38777 );
not ( n38779 , n38778 );
buf ( n38780 , n277495 );
buf ( n38781 , n38780 );
not ( n38782 , n38781 );
and ( n38783 , n38779 , n38782 );
buf ( n38784 , n38777 );
buf ( n38785 , n38780 );
and ( n38786 , n38784 , n38785 );
nor ( n38787 , n38783 , n38786 );
buf ( n38788 , n38787 );
buf ( n38789 , n38788 );
not ( n38790 , n38789 );
buf ( n38791 , n15387 );
buf ( n38792 , n15013 );
buf ( n38793 , n22226 );
buf ( n38794 , n24952 );
not ( n38795 , n38794 );
buf ( n38796 , n24995 );
nor ( n38797 , n38795 , n38796 );
buf ( n38798 , n38797 );
buf ( n38799 , n38798 );
and ( n38800 , n38793 , n38799 );
buf ( n38801 , n38800 );
buf ( n38802 , n38801 );
and ( n38803 , n38792 , n38802 );
buf ( n38804 , n38803 );
buf ( n38805 , n38804 );
and ( n38806 , n38791 , n38805 );
buf ( n38807 , n38801 );
not ( n38808 , n38807 );
buf ( n38809 , n15481 );
not ( n38810 , n38809 );
or ( n38811 , n38808 , n38810 );
buf ( n38812 , n22281 );
buf ( n38813 , n38798 );
and ( n38814 , n38812 , n38813 );
buf ( n38815 , n24979 );
buf ( n38816 , n24995 );
or ( n38817 , n38815 , n38816 );
buf ( n38818 , n25001 );
nand ( n38819 , n38817 , n38818 );
buf ( n38820 , n38819 );
buf ( n38821 , n38820 );
nor ( n38822 , n38814 , n38821 );
buf ( n38823 , n38822 );
buf ( n38824 , n38823 );
nand ( n38825 , n38811 , n38824 );
buf ( n38826 , n38825 );
buf ( n38827 , n38826 );
nor ( n38828 , n38806 , n38827 );
buf ( n38829 , n38828 );
buf ( n38830 , n38829 );
not ( n38831 , n38830 );
or ( n38832 , n38790 , n38831 );
buf ( n38833 , n38829 );
buf ( n38834 , n38788 );
or ( n38835 , n38833 , n38834 );
nand ( n38836 , n38832 , n38835 );
buf ( n38837 , n38836 );
buf ( n38838 , n38837 );
not ( n38839 , n38838 );
or ( n38840 , n38839 , n9432 );
nand ( n38841 , n277352 , n277460 );
nand ( n38842 , n38840 , n38841 );
and ( n38843 , n24834 , n38842 );
buf ( n38844 , n38843 );
not ( n38845 , n38844 );
nand ( n38846 , n23875 , n24897 , n24941 , n25024 );
nor ( n38847 , n30367 , n38846 );
not ( n38848 , n38847 );
or ( n38849 , n38845 , n38848 );
or ( n38850 , n38847 , n38844 );
nand ( n38851 , n38849 , n38850 );
buf ( n38852 , n38851 );
and ( n38853 , n38852 , n17409 );
and ( n38854 , n20940 , n38843 );
nor ( n38855 , n38853 , n38854 );
nand ( n38856 , n24837 , n38855 );
and ( n38857 , n38776 , n38856 );
or ( n38858 , n38775 , n38857 );
buf ( n38859 , n38858 );
buf ( n38860 , n38859 );
or ( n38861 , n33077 , n19216 );
and ( n38862 , n33099 , n19360 );
nand ( n38863 , n33116 , n29075 );
not ( n38864 , n19317 );
not ( n38865 , n33104 );
and ( n38866 , n38864 , n38865 );
and ( n38867 , n33162 , n33120 );
nor ( n38868 , n38866 , n38867 );
nand ( n38869 , n19387 , n18596 );
nand ( n38870 , n38863 , n38868 , n38869 );
nor ( n38871 , n38862 , n38870 );
nand ( n38872 , n33143 , n35863 );
and ( n38873 , n38871 , n38872 );
nand ( n38874 , n38861 , n38873 );
buf ( n38875 , n38874 );
buf ( n38876 , n38875 );
buf ( n38877 , n275554 );
not ( n38878 , n275925 );
buf ( n38879 , n38878 );
buf ( n38880 , n38879 );
not ( n38881 , n22936 );
not ( n38882 , n14830 );
or ( n38883 , n38881 , n38882 );
nand ( n38884 , n16384 , n27664 );
nand ( n38885 , n38883 , n38884 );
buf ( n38886 , n38885 );
buf ( n38887 , n38886 );
not ( n38888 , n10982 );
or ( n38889 , n9158 , n38888 );
buf ( n38890 , n10966 );
not ( n38891 , n38890 );
or ( n38892 , n9157 , n38891 );
nand ( n38893 , n38889 , n38892 );
buf ( n38894 , n38893 );
buf ( n38895 , n38894 );
not ( n38896 , n275929 );
buf ( n38897 , n38896 );
buf ( n38898 , n38897 );
or ( n38899 , n27696 , n20743 );
nand ( n38900 , n27711 , n16968 );
nand ( n38901 , n27724 , n20763 );
nand ( n38902 , n17411 , n27737 );
nand ( n38903 , n17502 , n27728 );
nand ( n38904 , n17562 , n13718 );
nand ( n38905 , n17545 , n32890 );
and ( n38906 , n38902 , n38903 , n38904 , n38905 );
and ( n38907 , n38900 , n38901 , n38906 );
nand ( n38908 , n38899 , n38907 );
buf ( n38909 , n38908 );
buf ( n38910 , n38909 );
not ( n38911 , n275925 );
buf ( n38912 , n38911 );
buf ( n38913 , n38912 );
not ( n38914 , n32992 );
not ( n38915 , n23789 );
and ( n38916 , n38914 , n38915 );
not ( n38917 , n20889 );
not ( n38918 , n33009 );
or ( n38919 , n38917 , n38918 );
and ( n38920 , n33026 , n20926 );
not ( n38921 , n17409 );
not ( n38922 , n33039 );
or ( n38923 , n38921 , n38922 );
nand ( n38924 , n20940 , n33044 );
nand ( n38925 , n38923 , n38924 );
nor ( n38926 , n38920 , n38925 );
nand ( n38927 , n38919 , n38926 );
nor ( n38928 , n38916 , n38927 );
or ( n38929 , n38928 , n21697 );
nand ( n38930 , n21696 , n13864 );
nand ( n38931 , n38929 , n38930 );
buf ( n38932 , n38931 );
buf ( n38933 , n38932 );
not ( n38934 , n275550 );
buf ( n38935 , n38934 );
buf ( n38936 , n38935 );
not ( n38937 , n24736 );
or ( n38938 , n38937 , n29044 );
nand ( n38939 , n29046 , n277457 );
nand ( n38940 , n38938 , n38939 );
buf ( n38941 , n38940 );
buf ( n38942 , n38941 );
not ( n38943 , n275925 );
buf ( n38944 , n38943 );
buf ( n38945 , n38944 );
buf ( n38946 , n275554 );
not ( n38947 , n16118 );
or ( n38948 , n38947 , n14830 );
or ( n38949 , n23806 , n14883 );
nand ( n38950 , n38948 , n38949 );
buf ( n38951 , n38950 );
buf ( n38952 , n38951 );
buf ( n38953 , n275554 );
not ( n38954 , n275925 );
buf ( n38955 , n38954 );
buf ( n38956 , n38955 );
buf ( n38957 , n275554 );
or ( n38958 , n36036 , n38891 );
and ( n38959 , n36047 , n275730 );
xor ( n38960 , n36114 , n20623 );
xor ( n38961 , n38960 , n36117 );
buf ( n38962 , n38961 );
not ( n38963 , n38962 );
not ( n38964 , n36155 );
or ( n38965 , n38963 , n38964 );
xor ( n38966 , n20633 , n36220 );
xor ( n38967 , n38966 , n36223 );
buf ( n38968 , n38967 );
nand ( n38969 , n36159 , n38968 );
nand ( n38970 , n38965 , n38969 );
nor ( n38971 , n38959 , n38970 );
nand ( n38972 , n38958 , n38971 );
nand ( n38973 , n38972 , n20645 );
xor ( n38974 , n20601 , n36312 );
xor ( n38975 , n38974 , n36314 );
buf ( n38976 , n38975 );
nand ( n38977 , n36267 , n38976 );
xor ( n38978 , n20593 , n36415 );
xor ( n38979 , n38978 , n36417 );
buf ( n38980 , n38979 );
nand ( n38981 , n36371 , n38980 );
and ( n38982 , n36474 , n38890 );
not ( n38983 , n11006 );
not ( n38984 , n34313 );
or ( n38985 , n38983 , n38984 );
or ( n38986 , n20654 , n275729 );
nand ( n38987 , n38985 , n38986 );
nor ( n38988 , n38982 , n38987 );
nand ( n38989 , n38973 , n38977 , n38981 , n38988 );
buf ( n38990 , n38989 );
buf ( n38991 , n38990 );
not ( n38992 , n16070 );
or ( n38993 , n38992 , n14830 );
nand ( n38994 , n14830 , n14885 );
nand ( n38995 , n38993 , n38994 );
buf ( n38996 , n38995 );
buf ( n38997 , n38996 );
or ( n38998 , n32785 , n21030 );
nand ( n38999 , n21030 , n19077 );
nand ( n39000 , n38998 , n38999 );
buf ( n39001 , n39000 );
buf ( n39002 , n39001 );
not ( n39003 , n275929 );
buf ( n39004 , n39003 );
buf ( n39005 , n39004 );
or ( n39006 , n25031 , n23887 );
not ( n39007 , n20951 );
or ( n39008 , n39007 , n14680 );
nand ( n39009 , n39006 , n39008 );
buf ( n39010 , n39009 );
buf ( n39011 , n39010 );
not ( n39012 , n18015 );
not ( n39013 , n22335 );
or ( n39014 , n39012 , n39013 );
not ( n39015 , n27884 );
or ( n39016 , n39015 , n22335 );
nand ( n39017 , n39014 , n39016 );
buf ( n39018 , n39017 );
buf ( n39019 , n39018 );
buf ( n39020 , n275554 );
not ( n39021 , n14806 );
and ( n39022 , n39021 , n23788 );
not ( n39023 , n20889 );
not ( n39024 , n16954 );
or ( n39025 , n39023 , n39024 );
and ( n39026 , n17401 , n20926 );
not ( n39027 , n15509 );
not ( n39028 , n20940 );
or ( n39029 , n39027 , n39028 );
nand ( n39030 , n17496 , n17409 );
nand ( n39031 , n39029 , n39030 );
nor ( n39032 , n39026 , n39031 );
nand ( n39033 , n39025 , n39032 );
nor ( n39034 , n39022 , n39033 );
or ( n39035 , n39034 , n21697 );
nand ( n39036 , n21696 , n13984 );
nand ( n39037 , n39035 , n39036 );
buf ( n39038 , n39037 );
buf ( n39039 , n39038 );
not ( n39040 , n19429 );
or ( n39041 , n39040 , n21774 );
nand ( n39042 , n21774 , n9509 );
nand ( n39043 , n39041 , n39042 );
buf ( n39044 , n39043 );
buf ( n39045 , n39044 );
buf ( n39046 , n275554 );
buf ( n39047 , n275554 );
not ( n39048 , n34302 );
not ( n39049 , n31420 );
or ( n39050 , n39048 , n39049 );
and ( n39051 , n31436 , n35900 );
nand ( n39052 , n31447 , n34307 );
nand ( n39053 , n28451 , n277941 );
nand ( n39054 , n29171 , n12294 );
nand ( n39055 , n34848 , n12357 );
nand ( n39056 , n20649 , n9327 );
and ( n39057 , n39054 , n39055 , n39056 );
nand ( n39058 , n39052 , n39053 , n39057 );
nor ( n39059 , n39051 , n39058 );
nand ( n39060 , n39050 , n39059 );
buf ( n39061 , n39060 );
buf ( n39062 , n39061 );
buf ( n39063 , n275554 );
or ( n39064 , n36631 , n26364 );
nand ( n39065 , n26389 , n26386 );
and ( n39066 , n39065 , n14545 );
nand ( n39067 , n36664 , n26367 );
nand ( n39068 , n36646 , n26374 );
nand ( n39069 , n26395 , n36638 );
nand ( n39070 , n32188 , n36634 );
nand ( n39071 , n39067 , n39068 , n39069 , n39070 );
nor ( n39072 , n39066 , n39071 );
nand ( n39073 , n39064 , n39072 );
buf ( n39074 , n39073 );
buf ( n39075 , n39074 );
not ( n39076 , n275550 );
buf ( n39077 , n39076 );
buf ( n39078 , n39077 );
buf ( n39079 , n275554 );
not ( n39080 , n33901 );
and ( n39081 , n39080 , n23788 );
not ( n39082 , n20889 );
not ( n39083 , n33927 );
or ( n39084 , n39082 , n39083 );
and ( n39085 , n33949 , n20926 );
nand ( n39086 , n33968 , n17409 );
nand ( n39087 , n20940 , n24891 );
nand ( n39088 , n39086 , n39087 );
nor ( n39089 , n39085 , n39088 );
nand ( n39090 , n39084 , n39089 );
nor ( n39091 , n39081 , n39090 );
or ( n39092 , n39091 , n23887 );
nand ( n39093 , n20953 , n14711 );
nand ( n39094 , n39092 , n39093 );
buf ( n39095 , n39094 );
buf ( n39096 , n39095 );
not ( n39097 , n275929 );
buf ( n39098 , n39097 );
buf ( n39099 , n39098 );
buf ( n39100 , n275554 );
not ( n39101 , n275925 );
buf ( n39102 , n39101 );
buf ( n39103 , n39102 );
or ( n39104 , n29377 , n27179 );
nand ( n39105 , n23708 , n11639 );
nand ( n39106 , n39104 , n39105 );
buf ( n39107 , n39106 );
buf ( n39108 , n39107 );
not ( n39109 , n16705 );
or ( n39110 , n39109 , n20961 );
not ( n39111 , n9435 );
or ( n39112 , n28247 , n39111 );
nand ( n39113 , n39110 , n39112 );
buf ( n39114 , n39113 );
buf ( n39115 , n39114 );
buf ( n39116 , n275554 );
not ( n39117 , n11120 );
or ( n39118 , n9158 , n39117 );
not ( n39119 , n36110 );
or ( n39120 , n9157 , n39119 );
nand ( n39121 , n39118 , n39120 );
buf ( n39122 , n39121 );
buf ( n39123 , n39122 );
and ( n39124 , n31468 , n275585 );
nor ( n39125 , n39124 , n34930 );
nand ( n39126 , n22914 , n31508 );
buf ( n39127 , n31517 );
buf ( n39128 , n31544 );
and ( n39129 , n39127 , n39128 );
buf ( n39130 , n39129 );
buf ( n39131 , n39130 );
not ( n39132 , n39131 );
buf ( n39133 , n23137 );
buf ( n39134 , n31506 );
and ( n39135 , n39133 , n39134 );
buf ( n39136 , n31493 );
buf ( n39137 , n30540 );
buf ( n39138 , n31506 );
and ( n39139 , n39136 , n39137 , n39138 );
buf ( n39140 , n39139 );
buf ( n39141 , n39140 );
buf ( n39142 , n31537 );
nor ( n39143 , n39135 , n39141 , n39142 );
buf ( n39144 , n39143 );
buf ( n39145 , n39144 );
not ( n39146 , n39145 );
or ( n39147 , n39132 , n39146 );
buf ( n39148 , n39144 );
buf ( n39149 , n39130 );
or ( n39150 , n39148 , n39149 );
nand ( n39151 , n39147 , n39150 );
buf ( n39152 , n39151 );
buf ( n39153 , n39152 );
nand ( n39154 , n22918 , n39153 );
buf ( n39155 , n31609 );
buf ( n39156 , n31636 );
and ( n39157 , n39155 , n39156 );
buf ( n39158 , n39157 );
buf ( n39159 , n39158 );
not ( n39160 , n39159 );
buf ( n39161 , n23362 );
buf ( n39162 , n31599 );
and ( n39163 , n39161 , n39162 );
buf ( n39164 , n31587 );
buf ( n39165 , n30574 );
buf ( n39166 , n31599 );
and ( n39167 , n39164 , n39165 , n39166 );
buf ( n39168 , n39167 );
buf ( n39169 , n39168 );
buf ( n39170 , n31629 );
nor ( n39171 , n39163 , n39169 , n39170 );
buf ( n39172 , n39171 );
buf ( n39173 , n39172 );
not ( n39174 , n39173 );
or ( n39175 , n39160 , n39174 );
buf ( n39176 , n39172 );
buf ( n39177 , n39158 );
or ( n39178 , n39176 , n39177 );
nand ( n39179 , n39175 , n39178 );
buf ( n39180 , n39179 );
buf ( n39181 , n39180 );
nand ( n39182 , n23152 , n39181 );
nand ( n39183 , n39125 , n39126 , n39154 , n39182 );
buf ( n39184 , n39183 );
buf ( n39185 , n39184 );
not ( n39186 , n35134 );
and ( n39187 , n39186 , n20987 );
not ( n39188 , n19358 );
not ( n39189 , n35145 );
or ( n39190 , n39188 , n39189 );
and ( n39191 , n35166 , n21001 );
or ( n39192 , n35183 , n19289 );
or ( n39193 , n22867 , n35189 );
nand ( n39194 , n39192 , n39193 );
nor ( n39195 , n39191 , n39194 );
nand ( n39196 , n39190 , n39195 );
nor ( n39197 , n39187 , n39196 );
or ( n39198 , n39197 , n24452 );
nand ( n39199 , n28146 , n18903 );
nand ( n39200 , n39198 , n39199 );
buf ( n39201 , n39200 );
buf ( n39202 , n39201 );
or ( n39203 , n37447 , n20951 );
nand ( n39204 , n20953 , n13924 );
nand ( n39205 , n39203 , n39204 );
buf ( n39206 , n39205 );
buf ( n39207 , n39206 );
not ( n39208 , n14560 );
not ( n39209 , n20950 );
or ( n39210 , n39208 , n39209 );
or ( n39211 , n37116 , n23887 );
nand ( n39212 , n39210 , n39211 );
buf ( n39213 , n39212 );
buf ( n39214 , n39213 );
not ( n39215 , n275550 );
buf ( n39216 , n39215 );
buf ( n39217 , n39216 );
or ( n39218 , n34035 , n21030 );
nand ( n39219 , n21030 , n18870 );
nand ( n39220 , n39218 , n39219 );
buf ( n39221 , n39220 );
buf ( n39222 , n39221 );
and ( n39223 , n9158 , n9123 );
not ( n39224 , n9158 );
and ( n39225 , n39224 , n277796 );
or ( n39226 , n39223 , n39225 );
buf ( n39227 , n39226 );
buf ( n39228 , n39227 );
buf ( n39229 , n275554 );
and ( n39230 , n9158 , n275946 );
not ( n39231 , n9158 );
and ( n39232 , n39231 , n11060 );
or ( n39233 , n39230 , n39232 );
buf ( n39234 , n39233 );
buf ( n39235 , n39234 );
buf ( n39236 , n19619 );
and ( n39237 , n18208 , n39236 );
not ( n39238 , n18208 );
buf ( n39239 , n21137 );
not ( n39240 , n39239 );
and ( n39241 , n19475 , n19621 );
nand ( n39242 , n19606 , n39241 );
not ( n39243 , n39242 );
or ( n39244 , n39240 , n39243 );
or ( n39245 , n39242 , n39239 );
nand ( n39246 , n39244 , n39245 );
buf ( n39247 , n39246 );
and ( n39248 , n39238 , n39247 );
nor ( n39249 , n39237 , n39248 );
or ( n39250 , n39249 , n19216 );
not ( n39251 , n21414 );
nand ( n39252 , n39251 , n21482 );
not ( n39253 , n39252 );
nor ( n39254 , n20072 , n19940 );
not ( n39255 , n39254 );
not ( n39256 , n20337 );
or ( n39257 , n39255 , n39256 );
not ( n39258 , n19941 );
not ( n39259 , n20345 );
or ( n39260 , n39258 , n39259 );
nand ( n39261 , n39260 , n19942 );
not ( n39262 , n39261 );
nand ( n39263 , n39257 , n39262 );
not ( n39264 , n39263 );
or ( n39265 , n39253 , n39264 );
or ( n39266 , n39263 , n39252 );
nand ( n39267 , n39265 , n39266 );
buf ( n39268 , n39267 );
and ( n39269 , n39268 , n33157 );
nand ( n39270 , n21560 , n21574 );
not ( n39271 , n39270 );
nor ( n39272 , n20401 , n20370 );
not ( n39273 , n39272 );
not ( n39274 , n20500 );
or ( n39275 , n39273 , n39274 );
or ( n39276 , n20508 , n20370 );
nand ( n39277 , n39276 , n20372 );
not ( n39278 , n39277 );
nand ( n39279 , n39275 , n39278 );
not ( n39280 , n39279 );
or ( n39281 , n39271 , n39280 );
or ( n39282 , n39279 , n39270 );
nand ( n39283 , n39281 , n39282 );
buf ( n39284 , n39283 );
and ( n39285 , n39284 , n19360 );
not ( n39286 , n19317 );
and ( n39287 , n29473 , n36762 );
not ( n39288 , n29473 );
and ( n39289 , n39288 , n18750 );
nor ( n39290 , n39287 , n39289 );
not ( n39291 , n39290 );
and ( n39292 , n39286 , n39291 );
buf ( n39293 , n21601 );
buf ( n39294 , n39293 );
and ( n39295 , n19221 , n39294 );
nor ( n39296 , n39292 , n39295 );
not ( n39297 , n21603 );
and ( n39298 , n20552 , n20521 );
nand ( n39299 , n20547 , n39298 );
not ( n39300 , n39299 );
or ( n39301 , n39297 , n39300 );
or ( n39302 , n39299 , n21603 );
nand ( n39303 , n39301 , n39302 );
buf ( n39304 , n39303 );
nand ( n39305 , n39304 , n29075 );
nand ( n39306 , n33840 , n18744 );
nand ( n39307 , n39296 , n39305 , n39306 );
nor ( n39308 , n39269 , n39285 , n39307 );
nand ( n39309 , n39250 , n39308 );
buf ( n39310 , n39309 );
buf ( n39311 , n39310 );
and ( n39312 , n23907 , n38566 );
not ( n39313 , n23907 );
and ( n39314 , n39313 , n38705 );
nor ( n39315 , n39312 , n39314 );
or ( n39316 , n39315 , n19216 );
and ( n39317 , n38735 , n19360 );
nand ( n39318 , n38750 , n29075 );
and ( n39319 , n33162 , n38739 );
and ( n39320 , n30138 , n30139 );
not ( n39321 , n30138 );
and ( n39322 , n39321 , n18668 );
nor ( n39323 , n39320 , n39322 );
not ( n39324 , n39323 );
nor ( n39325 , n39324 , n19317 );
nor ( n39326 , n39319 , n39325 );
nand ( n39327 , n19387 , n18680 );
nand ( n39328 , n39318 , n39326 , n39327 );
nor ( n39329 , n39317 , n39328 );
nand ( n39330 , n38721 , n35863 );
and ( n39331 , n39329 , n39330 );
nand ( n39332 , n39316 , n39331 );
buf ( n39333 , n39332 );
buf ( n39334 , n39333 );
and ( n39335 , n27179 , n277848 );
not ( n39336 , n27179 );
not ( n39337 , n29599 );
buf ( n39338 , n30837 );
buf ( n39339 , n30888 );
nand ( n39340 , n39338 , n39339 );
buf ( n39341 , n39340 );
buf ( n39342 , n39341 );
not ( n39343 , n39342 );
buf ( n39344 , n30830 );
buf ( n39345 , n39344 );
not ( n39346 , n39345 );
buf ( n39347 , n30823 );
nor ( n39348 , n39346 , n39347 );
buf ( n39349 , n39348 );
buf ( n39350 , n39349 );
not ( n39351 , n39350 );
buf ( n39352 , n27479 );
not ( n39353 , n39352 );
or ( n39354 , n39351 , n39353 );
buf ( n39355 , n39344 );
not ( n39356 , n39355 );
buf ( n39357 , n30869 );
buf ( n39358 , n39357 );
not ( n39359 , n39358 );
or ( n39360 , n39356 , n39359 );
buf ( n39361 , n30878 );
nand ( n39362 , n39360 , n39361 );
buf ( n39363 , n39362 );
buf ( n39364 , n39363 );
not ( n39365 , n39364 );
buf ( n39366 , n39365 );
buf ( n39367 , n39366 );
nand ( n39368 , n39354 , n39367 );
buf ( n39369 , n39368 );
buf ( n39370 , n39369 );
not ( n39371 , n39370 );
or ( n39372 , n39343 , n39371 );
buf ( n39373 , n39369 );
buf ( n39374 , n39341 );
or ( n39375 , n39373 , n39374 );
nand ( n39376 , n39372 , n39375 );
buf ( n39377 , n39376 );
buf ( n39378 , n39377 );
not ( n39379 , n39378 );
or ( n39380 , n39337 , n39379 );
nand ( n39381 , n30925 , n30953 );
not ( n39382 , n39381 );
not ( n39383 , n30921 );
nor ( n39384 , n39383 , n30932 );
not ( n39385 , n39384 );
not ( n39386 , n29728 );
or ( n39387 , n39385 , n39386 );
not ( n39388 , n30921 );
buf ( n39389 , n30945 );
not ( n39390 , n39389 );
or ( n39391 , n39388 , n39390 );
nand ( n39392 , n39391 , n30949 );
not ( n39393 , n39392 );
nand ( n39394 , n39387 , n39393 );
not ( n39395 , n39394 );
or ( n39396 , n39382 , n39395 );
or ( n39397 , n39394 , n39381 );
nand ( n39398 , n39396 , n39397 );
buf ( n39399 , n39398 );
and ( n39400 , n39399 , n23655 );
not ( n39401 , n23673 );
not ( n39402 , n30976 );
and ( n39403 , n29758 , n29750 );
not ( n39404 , n39403 );
or ( n39405 , n39402 , n39404 );
buf ( n39406 , n30972 );
nand ( n39407 , n39405 , n39406 );
not ( n39408 , n30979 );
nor ( n39409 , n39408 , n30972 );
nand ( n39410 , n31442 , n39409 );
nand ( n39411 , n39407 , n39410 );
buf ( n39412 , n39411 );
not ( n39413 , n39412 );
or ( n39414 , n39401 , n39413 );
and ( n39415 , n27520 , n12247 );
and ( n39416 , n22013 , n12182 );
nor ( n39417 , n39415 , n39416 );
nand ( n39418 , n39414 , n39417 );
nor ( n39419 , n39400 , n39418 );
nand ( n39420 , n39380 , n39419 );
and ( n39421 , n39336 , n39420 );
or ( n39422 , n39335 , n39421 );
buf ( n39423 , n39422 );
buf ( n39424 , n39423 );
not ( n39425 , n28436 );
buf ( n39426 , n28220 );
and ( n39427 , n39426 , n27495 );
not ( n39428 , n39426 );
not ( n39429 , n27495 );
and ( n39430 , n39428 , n39429 );
nor ( n39431 , n39427 , n39430 );
buf ( n39432 , n39431 );
not ( n39433 , n39432 );
or ( n39434 , n39425 , n39433 );
nand ( n39435 , n39434 , n9155 );
not ( n39436 , n22117 );
not ( n39437 , n39436 );
not ( n39438 , n22118 );
not ( n39439 , n39438 );
or ( n39440 , n39437 , n39439 );
buf ( n39441 , n22119 );
nand ( n39442 , n39440 , n39441 );
buf ( n39443 , n39442 );
nor ( n39444 , n39443 , n32812 );
buf ( n39445 , n21901 );
not ( n39446 , n39445 );
buf ( n39447 , n39446 );
buf ( n39448 , n39447 );
not ( n39449 , n39448 );
buf ( n39450 , n21903 );
not ( n39451 , n39450 );
or ( n39452 , n39449 , n39451 );
buf ( n39453 , n21903 );
not ( n39454 , n39453 );
buf ( n39455 , n39454 );
buf ( n39456 , n39455 );
buf ( n39457 , n21901 );
nand ( n39458 , n39456 , n39457 );
buf ( n39459 , n39458 );
buf ( n39460 , n39459 );
nand ( n39461 , n39452 , n39460 );
buf ( n39462 , n39461 );
buf ( n39463 , n39462 );
not ( n39464 , n32812 );
or ( n39465 , n39463 , n39464 );
nand ( n39466 , n39465 , n32815 );
or ( n39467 , n39444 , n39466 );
nand ( n39468 , n39467 , n9146 );
not ( n39469 , n39443 );
and ( n39470 , n11731 , n12687 , n12096 );
nand ( n39471 , n39469 , n39470 );
nand ( n39472 , n39468 , n39471 );
not ( n39473 , n11741 );
and ( n39474 , n39472 , n39473 );
or ( n39475 , n39443 , n32813 );
or ( n39476 , n39463 , n9136 );
nand ( n39477 , n39475 , n39476 );
nand ( n39478 , n39477 , n12108 );
nand ( n39479 , n12687 , n12101 );
or ( n39480 , n39463 , n39479 );
nand ( n39481 , n11732 , n11741 );
nand ( n39482 , n39480 , n39481 );
and ( n39483 , n20581 , n11060 );
not ( n39484 , n20581 );
and ( n39485 , n39484 , n275946 );
nor ( n39486 , n39483 , n39485 );
and ( n39487 , n39486 , n12688 );
nor ( n39488 , n39482 , n39487 );
nand ( n39489 , n39478 , n39488 );
nor ( n39490 , n39474 , n39489 );
nand ( n39491 , n39435 , n39490 );
or ( n39492 , n39491 , n35975 );
not ( n39493 , n11024 );
or ( n39494 , n22191 , n39493 );
nand ( n39495 , n39492 , n39494 );
buf ( n39496 , n39495 );
buf ( n39497 , n39496 );
buf ( n39498 , n275554 );
not ( n39499 , n275550 );
buf ( n39500 , n39499 );
buf ( n39501 , n39500 );
not ( n39502 , n275550 );
buf ( n39503 , n39502 );
buf ( n39504 , n39503 );
buf ( n39505 , n275554 );
buf ( n39506 , n275554 );
not ( n39507 , n278003 );
or ( n39508 , n39507 , n9158 );
or ( n39509 , n9144 , n9157 );
nand ( n39510 , n39508 , n39509 );
buf ( n39511 , n39510 );
buf ( n39512 , n39511 );
not ( n39513 , n275929 );
buf ( n39514 , n39513 );
buf ( n39515 , n39514 );
not ( n39516 , n275925 );
buf ( n39517 , n39516 );
buf ( n39518 , n39517 );
not ( n39519 , n275903 );
nor ( n39520 , n39519 , n275900 );
not ( n39521 , n39520 );
not ( n39522 , n275862 );
not ( n39523 , n39522 );
or ( n39524 , n39521 , n39523 );
or ( n39525 , n39522 , n39520 );
nand ( n39526 , n39524 , n39525 );
buf ( n39527 , n39526 );
buf ( n39528 , n39527 );
buf ( n39529 , n275554 );
not ( n39530 , n275929 );
buf ( n39531 , n39530 );
buf ( n39532 , n39531 );
not ( n39533 , n275929 );
buf ( n39534 , n39533 );
buf ( n39535 , n39534 );
buf ( n39536 , n275554 );
not ( n39537 , n275550 );
buf ( n39538 , n39537 );
buf ( n39539 , n39538 );
buf ( n39540 , n275554 );
buf ( n39541 , n275554 );
not ( n39542 , n33980 );
or ( n39543 , n21769 , n39542 );
not ( n39544 , n21769 );
not ( n39545 , n9469 );
or ( n39546 , n39544 , n39545 );
nand ( n39547 , n39543 , n39546 );
buf ( n39548 , n39547 );
buf ( n39549 , n39548 );
buf ( n39550 , n275554 );
buf ( n39551 , RI21a12898_77);
not ( n39552 , n39551 );
not ( n39553 , n39552 );
buf ( n39554 , n39553 );
buf ( n39555 , RI210beb80_291);
not ( n39556 , n39555 );
not ( n39557 , n39556 );
buf ( n39558 , n39557 );
xor ( n39559 , n39554 , n39558 );
buf ( n39560 , RI21077f78_506);
not ( n39561 , n39560 );
not ( n39562 , n39561 );
buf ( n39563 , n39562 );
not ( n39564 , n39563 );
xor ( n39565 , n39559 , n39564 );
xor ( n39566 , n36497 , n36501 );
and ( n39567 , n39566 , n36507 );
and ( n39568 , n36497 , n36501 );
or ( n39569 , n39567 , n39568 );
and ( n39570 , n39565 , n39569 );
not ( n39571 , n39570 );
or ( n39572 , n39565 , n39569 );
nand ( n39573 , n39571 , n39572 );
not ( n39574 , n39573 );
xor ( n39575 , n36493 , n36508 );
and ( n39576 , n39575 , n36511 );
and ( n39577 , n36493 , n36508 );
or ( n39578 , n39576 , n39577 );
not ( n39579 , n39578 );
or ( n39580 , n39574 , n39579 );
or ( n39581 , n39578 , n39573 );
nand ( n39582 , n39580 , n39581 );
buf ( n39583 , n39582 );
buf ( n39584 , n39583 );
buf ( n39585 , n275554 );
and ( n39586 , n21998 , n12686 );
nor ( n39587 , n39586 , n9100 );
buf ( n39588 , n9183 );
or ( n39589 , n39587 , n39588 );
nand ( n39590 , n39589 , n9411 );
nand ( n39591 , n39590 , n9158 );
buf ( n39592 , n39591 );
buf ( n39593 , n39592 );
buf ( n39594 , n275554 );
or ( n39595 , n33797 , n29866 );
and ( n39596 , n33817 , n20515 );
not ( n39597 , n37197 );
nand ( n39598 , n33826 , n29492 );
nand ( n39599 , n20563 , n33837 );
nand ( n39600 , n39597 , n39598 , n39599 );
nor ( n39601 , n39596 , n39600 );
nand ( n39602 , n33805 , n20353 );
not ( n39603 , n33832 );
nand ( n39604 , n39603 , n19648 );
and ( n39605 , n39601 , n39602 , n39604 );
nand ( n39606 , n39595 , n39605 );
buf ( n39607 , n39606 );
buf ( n39608 , n39607 );
or ( n39609 , n36842 , n21696 );
nand ( n39610 , n21697 , n13629 );
nand ( n39611 , n39609 , n39610 );
buf ( n39612 , n39611 );
buf ( n39613 , n39612 );
not ( n39614 , n22335 );
not ( n39615 , n25097 );
or ( n39616 , n39614 , n39615 );
not ( n39617 , n19887 );
or ( n39618 , n39617 , n22335 );
nand ( n39619 , n39616 , n39618 );
buf ( n39620 , n39619 );
buf ( n39621 , n39620 );
not ( n39622 , n22961 );
not ( n39623 , n14830 );
or ( n39624 , n39622 , n39623 );
nand ( n39625 , n16479 , n27664 );
nand ( n39626 , n39624 , n39625 );
buf ( n39627 , n39626 );
buf ( n39628 , n39627 );
not ( n39629 , n275925 );
buf ( n39630 , n39629 );
buf ( n39631 , n39630 );
not ( n39632 , n275550 );
buf ( n39633 , n39632 );
buf ( n39634 , n39633 );
not ( n39635 , n22944 );
not ( n39636 , n14830 );
or ( n39637 , n39635 , n39636 );
nand ( n39638 , n16435 , n27664 );
nand ( n39639 , n39637 , n39638 );
buf ( n39640 , n39639 );
buf ( n39641 , n39640 );
not ( n39642 , n275550 );
buf ( n39643 , n39642 );
buf ( n39644 , n39643 );
or ( n39645 , n34634 , n26364 );
nand ( n39646 , n34648 , n26370 );
nand ( n39647 , n34656 , n26374 );
and ( n39648 , n17504 , n13677 );
not ( n39649 , n17504 );
and ( n39650 , n39649 , n35588 );
nor ( n39651 , n39648 , n39650 );
nand ( n39652 , n31180 , n39651 );
and ( n39653 , n26395 , n34668 );
not ( n39654 , n32188 );
not ( n39655 , n34664 );
or ( n39656 , n39654 , n39655 );
not ( n39657 , n35589 );
nand ( n39658 , n39656 , n39657 );
nor ( n39659 , n39653 , n39658 );
and ( n39660 , n39646 , n39647 , n39652 , n39659 );
nand ( n39661 , n39645 , n39660 );
buf ( n39662 , n39661 );
buf ( n39663 , n39662 );
not ( n39664 , n26893 );
or ( n39665 , n39664 , n22335 );
or ( n39666 , n275557 , n19204 );
nand ( n39667 , n39665 , n39666 );
buf ( n39668 , n39667 );
buf ( n39669 , n39668 );
buf ( n39670 , n275554 );
buf ( n39671 , n275554 );
buf ( n39672 , n275554 );
not ( n39673 , n33077 );
and ( n39674 , n39673 , n23992 );
not ( n39675 , n21001 );
not ( n39676 , n33143 );
or ( n39677 , n39675 , n39676 );
and ( n39678 , n33099 , n19358 );
not ( n39679 , n19290 );
not ( n39680 , n33116 );
or ( n39681 , n39679 , n39680 );
nand ( n39682 , n19219 , n33120 );
nand ( n39683 , n39681 , n39682 );
nor ( n39684 , n39678 , n39683 );
nand ( n39685 , n39677 , n39684 );
nor ( n39686 , n39674 , n39685 );
or ( n39687 , n39686 , n21030 );
nand ( n39688 , n21030 , n18600 );
nand ( n39689 , n39687 , n39688 );
buf ( n39690 , n39689 );
buf ( n39691 , n39690 );
not ( n39692 , n275550 );
buf ( n39693 , n39692 );
buf ( n39694 , n39693 );
buf ( n39695 , n275554 );
not ( n39696 , n278051 );
or ( n39697 , n39696 , n9158 );
buf ( n39698 , n278032 );
not ( n39699 , n39698 );
or ( n39700 , n9157 , n39699 );
nand ( n39701 , n39697 , n39700 );
buf ( n39702 , n39701 );
buf ( n39703 , n39702 );
buf ( n39704 , n275554 );
buf ( n39705 , n275554 );
not ( n39706 , n34151 );
or ( n39707 , n39706 , n21774 );
nand ( n39708 , n21774 , n277340 );
nand ( n39709 , n39707 , n39708 );
buf ( n39710 , n39709 );
buf ( n39711 , n39710 );
not ( n39712 , n275925 );
buf ( n39713 , n39712 );
buf ( n39714 , n39713 );
not ( n39715 , n275929 );
buf ( n39716 , n39715 );
buf ( n39717 , n39716 );
buf ( n39718 , n275554 );
buf ( n39719 , n275554 );
buf ( n39720 , n275554 );
buf ( n39721 , RI210cdf40_249);
buf ( n39722 , n39721 );
not ( n39723 , n39722 );
buf ( n39724 , RI2107db58_464);
buf ( n39725 , n39724 );
not ( n39726 , n39725 );
or ( n39727 , n39723 , n39726 );
not ( n39728 , n39725 );
not ( n39729 , n39722 );
and ( n39730 , n39728 , n39729 );
buf ( n39731 , RI21069950_647);
buf ( n39732 , n39731 );
nor ( n39733 , n39730 , n39732 );
nand ( n39734 , n39727 , n39733 );
buf ( n39735 , n39734 );
buf ( n39736 , n39735 );
not ( n39737 , n34302 );
not ( n39738 , n39378 );
or ( n39739 , n39737 , n39738 );
and ( n39740 , n39399 , n35900 );
nand ( n39741 , n39412 , n34307 );
nand ( n39742 , n28451 , n277868 );
nand ( n39743 , n32755 , n12247 );
and ( n39744 , n34311 , n12182 );
and ( n39745 , n34313 , n9336 );
nor ( n39746 , n39744 , n39745 );
and ( n39747 , n39743 , n39746 );
nand ( n39748 , n39741 , n39742 , n39747 );
nor ( n39749 , n39740 , n39748 );
nand ( n39750 , n39739 , n39749 );
buf ( n39751 , n39750 );
buf ( n39752 , n39751 );
not ( n39753 , n275929 );
buf ( n39754 , n39753 );
buf ( n39755 , n39754 );
not ( n39756 , n275925 );
buf ( n39757 , n39756 );
buf ( n39758 , n39757 );
or ( n39759 , n27843 , n29866 );
nand ( n39760 , n28049 , n20353 );
nand ( n39761 , n28120 , n30132 );
not ( n39762 , n19649 );
not ( n39763 , n18652 );
and ( n39764 , n30145 , n39763 );
not ( n39765 , n30145 );
and ( n39766 , n39765 , n18653 );
nor ( n39767 , n39764 , n39766 );
not ( n39768 , n39767 );
and ( n39769 , n39762 , n39768 );
nand ( n39770 , n28140 , n31095 );
nand ( n39771 , n29494 , n27885 );
nand ( n39772 , n30179 , n18653 );
nand ( n39773 , n39770 , n39771 , n39772 );
nor ( n39774 , n39769 , n39773 );
and ( n39775 , n39760 , n39761 , n39774 );
nand ( n39776 , n39759 , n39775 );
buf ( n39777 , n39776 );
buf ( n39778 , n39777 );
or ( n39779 , n33994 , n32073 );
not ( n39780 , n19651 );
not ( n39781 , n18862 );
and ( n39782 , n39780 , n39781 );
nand ( n39783 , n34008 , n20353 );
nand ( n39784 , n34018 , n20515 );
and ( n39785 , n29492 , n34024 );
nor ( n39786 , n19639 , n30615 );
nor ( n39787 , n39785 , n39786 );
nand ( n39788 , n20563 , n34029 );
nand ( n39789 , n39783 , n39784 , n39787 , n39788 );
nor ( n39790 , n39782 , n39789 );
nand ( n39791 , n39779 , n39790 );
buf ( n39792 , n39791 );
buf ( n39793 , n39792 );
buf ( n39794 , n275554 );
buf ( n39795 , n275554 );
buf ( n39796 , n275554 );
buf ( n39797 , n275554 );
not ( n39798 , n275925 );
buf ( n39799 , n39798 );
buf ( n39800 , n39799 );
nand ( n39801 , n28186 , n27586 );
nand ( n39802 , n28196 , n27561 );
and ( n39803 , n39801 , n39802 );
nand ( n39804 , n28219 , n27576 );
and ( n39805 , n28231 , n12189 );
not ( n39806 , n10873 );
or ( n39807 , n28233 , n39806 );
nand ( n39808 , n28236 , n29169 );
nand ( n39809 , n39807 , n39808 );
nor ( n39810 , n39805 , n39809 );
nand ( n39811 , n31459 , n12233 );
nand ( n39812 , n39803 , n39804 , n39810 , n39811 );
buf ( n39813 , n39812 );
buf ( n39814 , n39813 );
not ( n39815 , n275929 );
buf ( n39816 , n39815 );
buf ( n39817 , n39816 );
not ( n39818 , n275929 );
buf ( n39819 , n39818 );
buf ( n39820 , n39819 );
not ( n39821 , n275929 );
buf ( n39822 , n39821 );
buf ( n39823 , n39822 );
not ( n39824 , n275929 );
buf ( n39825 , n39824 );
buf ( n39826 , n39825 );
not ( n39827 , n275550 );
buf ( n39828 , n39827 );
buf ( n39829 , n39828 );
and ( n39830 , n22335 , n28957 );
not ( n39831 , n22335 );
and ( n39832 , n39831 , n24086 );
or ( n39833 , n39830 , n39832 );
buf ( n39834 , n39833 );
buf ( n39835 , n39834 );
not ( n39836 , n275550 );
buf ( n39837 , n39836 );
buf ( n39838 , n39837 );
buf ( n39839 , n275554 );
and ( n39840 , n31719 , n277860 );
not ( n39841 , n31719 );
and ( n39842 , n39841 , n39420 );
or ( n39843 , n39840 , n39842 );
buf ( n39844 , n39843 );
buf ( n39845 , n39844 );
and ( n39846 , n9158 , n9041 );
not ( n39847 , n9158 );
and ( n39848 , n39847 , n277607 );
or ( n39849 , n39846 , n39848 );
buf ( n39850 , n39849 );
buf ( n39851 , n39850 );
buf ( n39852 , n275554 );
not ( n39853 , n275925 );
buf ( n39854 , n39853 );
buf ( n39855 , n39854 );
or ( n39856 , n36879 , n26365 );
nand ( n39857 , n23418 , n26370 );
nand ( n39858 , n23433 , n26374 );
not ( n39859 , n36888 );
nor ( n39860 , n39859 , n26390 );
not ( n39861 , n37273 );
nand ( n39862 , n23442 , n32188 );
nand ( n39863 , n26395 , n23447 );
nand ( n39864 , n39861 , n39862 , n39863 );
nor ( n39865 , n39860 , n39864 );
and ( n39866 , n39857 , n39858 , n39865 );
nand ( n39867 , n39856 , n39866 );
buf ( n39868 , n39867 );
buf ( n39869 , n39868 );
buf ( n39870 , n275554 );
nand ( n39871 , n25064 , n26103 );
buf ( n39872 , n25161 );
not ( n39873 , n39872 );
buf ( n39874 , n25239 );
nand ( n39875 , n39873 , n39874 );
buf ( n39876 , n39875 );
buf ( n39877 , n39876 );
not ( n39878 , n39877 );
buf ( n39879 , n25221 );
not ( n39880 , n39879 );
buf ( n39881 , n39880 );
buf ( n39882 , n39881 );
buf ( n39883 , n25170 );
or ( n39884 , n39882 , n39883 );
buf ( n39885 , n25233 );
nand ( n39886 , n39884 , n39885 );
buf ( n39887 , n39886 );
buf ( n39888 , n39887 );
not ( n39889 , n39888 );
or ( n39890 , n39878 , n39889 );
buf ( n39891 , n39887 );
buf ( n39892 , n39876 );
or ( n39893 , n39891 , n39892 );
nand ( n39894 , n39890 , n39893 );
buf ( n39895 , n39894 );
buf ( n39896 , n39895 );
not ( n39897 , n39896 );
nor ( n39898 , n39897 , n25389 );
nand ( n39899 , n25397 , n275773 );
buf ( n39900 , n25484 );
not ( n39901 , n39900 );
buf ( n39902 , n25560 );
nand ( n39903 , n39901 , n39902 );
buf ( n39904 , n39903 );
buf ( n39905 , n39904 );
not ( n39906 , n39905 );
buf ( n39907 , n31226 );
buf ( n39908 , n25491 );
or ( n39909 , n39907 , n39908 );
buf ( n39910 , n25554 );
nand ( n39911 , n39909 , n39910 );
buf ( n39912 , n39911 );
buf ( n39913 , n39912 );
not ( n39914 , n39913 );
or ( n39915 , n39906 , n39914 );
buf ( n39916 , n39912 );
buf ( n39917 , n39904 );
or ( n39918 , n39916 , n39917 );
nand ( n39919 , n39915 , n39918 );
buf ( n39920 , n39919 );
buf ( n39921 , n39920 );
and ( n39922 , n25402 , n39921 );
not ( n39923 , n18391 );
nor ( n39924 , n39923 , n19639 );
nor ( n39925 , n39922 , n39924 );
buf ( n39926 , n25800 );
not ( n39927 , n39926 );
buf ( n39928 , n25876 );
nand ( n39929 , n39927 , n39928 );
buf ( n39930 , n39929 );
buf ( n39931 , n39930 );
not ( n39932 , n39931 );
buf ( n39933 , n31247 );
buf ( n39934 , n25807 );
or ( n39935 , n39933 , n39934 );
buf ( n39936 , n25870 );
nand ( n39937 , n39935 , n39936 );
buf ( n39938 , n39937 );
buf ( n39939 , n39938 );
not ( n39940 , n39939 );
or ( n39941 , n39932 , n39940 );
buf ( n39942 , n39938 );
buf ( n39943 , n39930 );
or ( n39944 , n39942 , n39943 );
nand ( n39945 , n39941 , n39944 );
buf ( n39946 , n39945 );
buf ( n39947 , n39946 );
nand ( n39948 , n28761 , n39947 );
nand ( n39949 , n39899 , n39925 , n39948 );
nor ( n39950 , n39898 , n39949 );
buf ( n39951 , n26109 );
not ( n39952 , n39951 );
buf ( n39953 , n26186 );
nand ( n39954 , n39952 , n39953 );
buf ( n39955 , n39954 );
buf ( n39956 , n39955 );
not ( n39957 , n39956 );
buf ( n39958 , n31269 );
buf ( n39959 , n26116 );
or ( n39960 , n39958 , n39959 );
buf ( n39961 , n26180 );
nand ( n39962 , n39960 , n39961 );
buf ( n39963 , n39962 );
buf ( n39964 , n39963 );
not ( n39965 , n39964 );
or ( n39966 , n39957 , n39965 );
buf ( n39967 , n39963 );
buf ( n39968 , n39955 );
or ( n39969 , n39967 , n39968 );
nand ( n39970 , n39966 , n39969 );
buf ( n39971 , n39970 );
buf ( n39972 , n39971 );
nand ( n39973 , n26027 , n39972 );
nand ( n39974 , n39871 , n39950 , n39973 );
buf ( n39975 , n39974 );
buf ( n39976 , n39975 );
not ( n39977 , n275550 );
buf ( n39978 , n39977 );
buf ( n39979 , n39978 );
and ( n39980 , n22193 , n278062 );
not ( n39981 , n22193 );
and ( n39982 , n39981 , n27526 );
nor ( n39983 , n39980 , n39982 );
buf ( n39984 , n39983 );
buf ( n39985 , n39984 );
not ( n39986 , n11490 );
or ( n39987 , n36036 , n39986 );
and ( n39988 , n36045 , n275672 );
buf ( n39989 , n11490 );
buf ( n39990 , n11467 );
not ( n39991 , n39990 );
nand ( n39992 , n39989 , n39991 );
not ( n39993 , n39992 );
nor ( n39994 , n39989 , n39991 );
nor ( n39995 , n39993 , n39994 );
not ( n39996 , n39995 );
and ( n39997 , n36137 , n36068 , n36054 );
nand ( n39998 , n36146 , n36054 );
nand ( n39999 , n39998 , n36053 );
nor ( n40000 , n39997 , n39999 );
not ( n40001 , n40000 );
or ( n40002 , n39996 , n40001 );
or ( n40003 , n40000 , n39995 );
nand ( n40004 , n40002 , n40003 );
buf ( n40005 , n40004 );
not ( n40006 , n40005 );
not ( n40007 , n36155 );
or ( n40008 , n40006 , n40007 );
buf ( n40009 , n11490 );
buf ( n40010 , n11474 );
not ( n40011 , n40010 );
nand ( n40012 , n40009 , n40011 );
not ( n40013 , n40012 );
nor ( n40014 , n40009 , n40011 );
nor ( n40015 , n40013 , n40014 );
not ( n40016 , n40015 );
and ( n40017 , n36243 , n36179 , n36166 );
nand ( n40018 , n36252 , n36166 );
nand ( n40019 , n40018 , n36164 );
nor ( n40020 , n40017 , n40019 );
not ( n40021 , n40020 );
or ( n40022 , n40016 , n40021 );
or ( n40023 , n40020 , n40015 );
nand ( n40024 , n40022 , n40023 );
buf ( n40025 , n40024 );
nand ( n40026 , n36159 , n40025 );
nand ( n40027 , n40008 , n40026 );
nor ( n40028 , n39988 , n40027 );
nand ( n40029 , n39987 , n40028 );
nand ( n40030 , n40029 , n20645 );
buf ( n40031 , n11490 );
not ( n40032 , n40031 );
buf ( n40033 , n11467 );
nand ( n40034 , n40032 , n40033 );
not ( n40035 , n40034 );
not ( n40036 , n40031 );
nor ( n40037 , n40036 , n40033 );
nor ( n40038 , n40035 , n40037 );
not ( n40039 , n40038 );
and ( n40040 , n36353 , n36285 , n36271 );
not ( n40041 , n36271 );
or ( n40042 , n36363 , n40041 );
nand ( n40043 , n40042 , n36274 );
nor ( n40044 , n40040 , n40043 );
not ( n40045 , n40044 );
or ( n40046 , n40039 , n40045 );
or ( n40047 , n40044 , n40038 );
nand ( n40048 , n40046 , n40047 );
buf ( n40049 , n40048 );
nand ( n40050 , n36267 , n40049 );
buf ( n40051 , n11490 );
not ( n40052 , n40051 );
buf ( n40053 , n11474 );
nand ( n40054 , n40052 , n40053 );
not ( n40055 , n40054 );
not ( n40056 , n40051 );
nor ( n40057 , n40056 , n40053 );
nor ( n40058 , n40055 , n40057 );
not ( n40059 , n40058 );
and ( n40060 , n36456 , n36389 , n36375 );
not ( n40061 , n36375 );
or ( n40062 , n36466 , n40061 );
nand ( n40063 , n40062 , n36378 );
nor ( n40064 , n40060 , n40063 );
not ( n40065 , n40064 );
or ( n40066 , n40059 , n40065 );
or ( n40067 , n40064 , n40058 );
nand ( n40068 , n40066 , n40067 );
buf ( n40069 , n40068 );
nand ( n40070 , n36371 , n40069 );
and ( n40071 , n36474 , n11490 );
or ( n40072 , n20654 , n275671 );
nand ( n40073 , n20649 , n9310 );
nand ( n40074 , n40072 , n40073 );
nor ( n40075 , n40071 , n40074 );
nand ( n40076 , n40030 , n40050 , n40070 , n40075 );
buf ( n40077 , n40076 );
buf ( n40078 , n40077 );
buf ( n40079 , n275554 );
and ( n40080 , n21990 , n28408 );
or ( n40081 , n29172 , n12340 );
or ( n40082 , n28459 , n12128 );
nand ( n40083 , n20649 , n9277 );
nand ( n40084 , n40081 , n40082 , n40083 );
nor ( n40085 , n40080 , n40084 );
nand ( n40086 , n22049 , n29163 );
nand ( n40087 , n32751 , n22141 );
not ( n40088 , n28450 );
not ( n40089 , n10788 );
nand ( n40090 , n40088 , n40089 );
nand ( n40091 , n40085 , n40086 , n40087 , n40090 );
buf ( n40092 , n40091 );
buf ( n40093 , n40092 );
not ( n40094 , n275550 );
buf ( n40095 , n40094 );
buf ( n40096 , n40095 );
not ( n40097 , n275550 );
buf ( n40098 , n40097 );
buf ( n40099 , n40098 );
buf ( n40100 , n275554 );
not ( n40101 , n11159 );
or ( n40102 , n9158 , n40101 );
not ( n40103 , n11144 );
or ( n40104 , n9157 , n40103 );
nand ( n40105 , n40102 , n40104 );
buf ( n40106 , n40105 );
buf ( n40107 , n40106 );
buf ( n40108 , n275554 );
not ( n40109 , n35552 );
not ( n40110 , n275744 );
not ( n40111 , n40110 );
and ( n40112 , n40109 , n40111 );
and ( n40113 , n17542 , n14761 );
nor ( n40114 , n40112 , n40113 );
xor ( n40115 , n23235 , n23236 );
buf ( n40116 , n40115 );
buf ( n40117 , n40116 );
nand ( n40118 , n23152 , n40117 );
xor ( n40119 , n23006 , n23007 );
buf ( n40120 , n40119 );
buf ( n40121 , n40120 );
nand ( n40122 , n22918 , n40121 );
nand ( n40123 , n22914 , n29258 );
nand ( n40124 , n40114 , n40118 , n40122 , n40123 );
buf ( n40125 , n40124 );
buf ( n40126 , n40125 );
buf ( n40127 , n275554 );
not ( n40128 , n275550 );
buf ( n40129 , n40128 );
buf ( n40130 , n40129 );
not ( n40131 , n275925 );
buf ( n40132 , n40131 );
buf ( n40133 , n40132 );
not ( n40134 , n275925 );
buf ( n40135 , n40134 );
buf ( n40136 , n40135 );
buf ( n40137 , n275554 );
not ( n40138 , n275925 );
buf ( n40139 , n40138 );
buf ( n40140 , n40139 );
buf ( n40141 , n275554 );
buf ( n40142 , n275554 );
buf ( n40143 , n275554 );
not ( n40144 , n27783 );
or ( n40145 , n40144 , n21774 );
nand ( n40146 , n21774 , n9769 );
nand ( n40147 , n40145 , n40146 );
buf ( n40148 , n40147 );
buf ( n40149 , n40148 );
not ( n40150 , n275550 );
buf ( n40151 , n40150 );
buf ( n40152 , n40151 );
and ( n40153 , n19143 , n19201 );
nor ( n40154 , n40153 , n19140 );
or ( n40155 , n40154 , n25394 );
nand ( n40156 , n40155 , n19639 );
buf ( n40157 , n40156 );
buf ( n40158 , n40157 );
not ( n40159 , n275550 );
buf ( n40160 , n40159 );
buf ( n40161 , n40160 );
not ( n40162 , n275929 );
buf ( n40163 , n40162 );
buf ( n40164 , n40163 );
not ( n40165 , n275550 );
buf ( n40166 , n40165 );
buf ( n40167 , n40166 );
buf ( n40168 , n275554 );
not ( n40169 , n275929 );
buf ( n40170 , n40169 );
buf ( n40171 , n40170 );
or ( n40172 , n34739 , n21697 );
nand ( n40173 , n21697 , n13549 );
nand ( n40174 , n40172 , n40173 );
buf ( n40175 , n40174 );
buf ( n40176 , n40175 );
nand ( n40177 , n29346 , n28408 );
nand ( n40178 , n29359 , n28430 );
nand ( n40179 , n29369 , n28440 );
nand ( n40180 , n28451 , n32608 );
and ( n40181 , n28455 , n32605 );
or ( n40182 , n28459 , n12131 );
nand ( n40183 , n20649 , n9295 );
nand ( n40184 , n40182 , n40183 );
nor ( n40185 , n40181 , n40184 );
and ( n40186 , n40179 , n40180 , n40185 );
nand ( n40187 , n40177 , n40178 , n40186 );
buf ( n40188 , n40187 );
buf ( n40189 , n40188 );
or ( n40190 , n26636 , n32074 );
and ( n40191 , n27046 , n20515 );
and ( n40192 , n30141 , n18552 );
not ( n40193 , n30141 );
not ( n40194 , n18551 );
and ( n40195 , n40193 , n40194 );
nor ( n40196 , n40192 , n40195 );
not ( n40197 , n40196 );
not ( n40198 , n19650 );
or ( n40199 , n40197 , n40198 );
nand ( n40200 , n27079 , n31095 );
nand ( n40201 , n20563 , n27050 );
nand ( n40202 , n30179 , n18552 );
and ( n40203 , n40200 , n40201 , n40202 );
nand ( n40204 , n40199 , n40203 );
nor ( n40205 , n40191 , n40204 );
nand ( n40206 , n26944 , n20353 );
and ( n40207 , n40205 , n40206 );
nand ( n40208 , n40190 , n40207 );
buf ( n40209 , n40208 );
buf ( n40210 , n40209 );
not ( n40211 , n275550 );
buf ( n40212 , n40211 );
buf ( n40213 , n40212 );
buf ( n40214 , n275554 );
not ( n40215 , n275929 );
buf ( n40216 , n40215 );
buf ( n40217 , n40216 );
buf ( n40218 , n275554 );
not ( n40219 , n39432 );
or ( n40220 , n40219 , n28437 );
nand ( n40221 , n29234 , n11034 );
and ( n40222 , n28407 , n39463 );
and ( n40223 , n39443 , n28427 );
not ( n40224 , n28449 );
and ( n40225 , n40224 , n12316 );
nor ( n40226 , n40222 , n40223 , n40225 );
nand ( n40227 , n40220 , n40221 , n40226 );
buf ( n40228 , n40227 );
buf ( n40229 , n40228 );
not ( n40230 , n275550 );
buf ( n40231 , n40230 );
buf ( n40232 , n40231 );
not ( n40233 , n275929 );
buf ( n40234 , n40233 );
buf ( n40235 , n40234 );
not ( n40236 , n275929 );
buf ( n40237 , n40236 );
buf ( n40238 , n40237 );
and ( n40239 , n31468 , n275629 );
nor ( n40240 , n14830 , n37896 );
nor ( n40241 , n40239 , n40240 );
nand ( n40242 , n22914 , n22936 );
buf ( n40243 , n22956 );
not ( n40244 , n40243 );
buf ( n40245 , n22942 );
nor ( n40246 , n40244 , n40245 );
buf ( n40247 , n40246 );
buf ( n40248 , n40247 );
not ( n40249 , n40248 );
buf ( n40250 , n22996 );
buf ( n40251 , n23043 );
buf ( n40252 , n23054 );
not ( n40253 , n40252 );
buf ( n40254 , n40253 );
buf ( n40255 , n40254 );
and ( n40256 , n40250 , n40251 , n40255 );
buf ( n40257 , n40254 );
not ( n40258 , n40257 );
buf ( n40259 , n22984 );
not ( n40260 , n40259 );
or ( n40261 , n40258 , n40260 );
buf ( n40262 , n22950 );
nand ( n40263 , n40261 , n40262 );
buf ( n40264 , n40263 );
buf ( n40265 , n40264 );
nor ( n40266 , n40256 , n40265 );
buf ( n40267 , n40266 );
buf ( n40268 , n40267 );
not ( n40269 , n40268 );
or ( n40270 , n40249 , n40269 );
buf ( n40271 , n40267 );
buf ( n40272 , n40247 );
or ( n40273 , n40271 , n40272 );
nand ( n40274 , n40270 , n40273 );
buf ( n40275 , n40274 );
buf ( n40276 , n40275 );
nand ( n40277 , n22918 , n40276 );
buf ( n40278 , n23188 );
not ( n40279 , n40278 );
buf ( n40280 , n23175 );
nor ( n40281 , n40279 , n40280 );
buf ( n40282 , n40281 );
buf ( n40283 , n40282 );
not ( n40284 , n40283 );
buf ( n40285 , n23226 );
buf ( n40286 , n23272 );
buf ( n40287 , n23283 );
not ( n40288 , n40287 );
buf ( n40289 , n40288 );
buf ( n40290 , n40289 );
and ( n40291 , n40285 , n40286 , n40290 );
buf ( n40292 , n40289 );
not ( n40293 , n40292 );
buf ( n40294 , n23214 );
not ( n40295 , n40294 );
or ( n40296 , n40293 , n40295 );
buf ( n40297 , n23182 );
nand ( n40298 , n40296 , n40297 );
buf ( n40299 , n40298 );
buf ( n40300 , n40299 );
nor ( n40301 , n40291 , n40300 );
buf ( n40302 , n40301 );
buf ( n40303 , n40302 );
not ( n40304 , n40303 );
or ( n40305 , n40284 , n40304 );
buf ( n40306 , n40302 );
buf ( n40307 , n40282 );
or ( n40308 , n40306 , n40307 );
nand ( n40309 , n40305 , n40308 );
buf ( n40310 , n40309 );
buf ( n40311 , n40310 );
nand ( n40312 , n23152 , n40311 );
nand ( n40313 , n40241 , n40242 , n40277 , n40312 );
buf ( n40314 , n40313 );
buf ( n40315 , n40314 );
or ( n40316 , n33272 , n19216 );
and ( n40317 , n33236 , n19360 );
nand ( n40318 , n33245 , n29075 );
not ( n40319 , n19317 );
and ( n40320 , n30135 , n18614 );
not ( n40321 , n30135 );
and ( n40322 , n40321 , n30136 );
nor ( n40323 , n40320 , n40322 );
not ( n40324 , n40323 );
and ( n40325 , n40319 , n40324 );
and ( n40326 , n19221 , n33250 );
nor ( n40327 , n40325 , n40326 );
nand ( n40328 , n33840 , n18625 );
nand ( n40329 , n40318 , n40327 , n40328 );
nor ( n40330 , n40317 , n40329 );
nand ( n40331 , n33222 , n35863 );
nand ( n40332 , n40316 , n40330 , n40331 );
buf ( n40333 , n40332 );
buf ( n40334 , n40333 );
buf ( n40335 , n275554 );
or ( n40336 , n39034 , n23887 );
nand ( n40337 , n20953 , n13996 );
nand ( n40338 , n40336 , n40337 );
buf ( n40339 , n40338 );
buf ( n40340 , n40339 );
buf ( n40341 , n275554 );
not ( n40342 , n275550 );
buf ( n40343 , n40342 );
buf ( n40344 , n40343 );
and ( n40345 , n26516 , n33297 );
not ( n40346 , n26516 );
buf ( n40347 , n27814 );
not ( n40348 , n40347 );
nand ( n40349 , n26632 , n26553 );
not ( n40350 , n40349 );
or ( n40351 , n40348 , n40350 );
or ( n40352 , n40349 , n40347 );
nand ( n40353 , n40351 , n40352 );
buf ( n40354 , n40353 );
and ( n40355 , n40346 , n40354 );
nor ( n40356 , n40345 , n40355 );
not ( n40357 , n40356 );
and ( n40358 , n40357 , n26638 );
not ( n40359 , n21001 );
not ( n40360 , n28010 );
nand ( n40361 , n40360 , n28029 );
not ( n40362 , n40361 );
not ( n40363 , n26733 );
nor ( n40364 , n40363 , n26912 );
not ( n40365 , n40364 );
nor ( n40366 , n40365 , n26853 );
not ( n40367 , n40366 );
not ( n40368 , n26915 );
or ( n40369 , n40367 , n40368 );
not ( n40370 , n40364 );
not ( n40371 , n26928 );
or ( n40372 , n40370 , n40371 );
and ( n40373 , n26935 , n26733 );
not ( n40374 , n26734 );
nor ( n40375 , n40373 , n40374 );
nand ( n40376 , n40372 , n40375 );
not ( n40377 , n40376 );
nand ( n40378 , n40369 , n40377 );
not ( n40379 , n40378 );
or ( n40380 , n40362 , n40379 );
or ( n40381 , n40378 , n40361 );
nand ( n40382 , n40380 , n40381 );
buf ( n40383 , n40382 );
not ( n40384 , n40383 );
or ( n40385 , n40359 , n40384 );
not ( n40386 , n28075 );
nand ( n40387 , n40386 , n28098 );
not ( n40388 , n40387 );
nor ( n40389 , n27014 , n26959 );
not ( n40390 , n40389 );
nor ( n40391 , n40390 , n26991 );
not ( n40392 , n40391 );
not ( n40393 , n27020 );
or ( n40394 , n40392 , n40393 );
and ( n40395 , n40389 , n27034 );
not ( n40396 , n26960 );
not ( n40397 , n27039 );
or ( n40398 , n40396 , n40397 );
nand ( n40399 , n40398 , n26961 );
nor ( n40400 , n40395 , n40399 );
nand ( n40401 , n40394 , n40400 );
not ( n40402 , n40401 );
or ( n40403 , n40388 , n40402 );
or ( n40404 , n40401 , n40387 );
nand ( n40405 , n40403 , n40404 );
buf ( n40406 , n40405 );
and ( n40407 , n40406 , n19358 );
buf ( n40408 , n28129 );
buf ( n40409 , n40408 );
not ( n40410 , n40409 );
not ( n40411 , n19219 );
or ( n40412 , n40410 , n40411 );
not ( n40413 , n28131 );
nand ( n40414 , n35459 , n27055 );
nor ( n40415 , n27065 , n40414 );
nand ( n40416 , n24314 , n40415 );
not ( n40417 , n40416 );
or ( n40418 , n40413 , n40417 );
or ( n40419 , n40416 , n28131 );
nand ( n40420 , n40418 , n40419 );
buf ( n40421 , n40420 );
nand ( n40422 , n40421 , n19290 );
nand ( n40423 , n40412 , n40422 );
nor ( n40424 , n40407 , n40423 );
nand ( n40425 , n40385 , n40424 );
nor ( n40426 , n40358 , n40425 );
or ( n40427 , n40426 , n28146 );
nand ( n40428 , n24450 , n18530 );
nand ( n40429 , n40427 , n40428 );
buf ( n40430 , n40429 );
buf ( n40431 , n40430 );
buf ( n40432 , n275554 );
not ( n40433 , n275929 );
buf ( n40434 , n40433 );
buf ( n40435 , n40434 );
buf ( n40436 , n275554 );
not ( n40437 , n275550 );
buf ( n40438 , n40437 );
buf ( n40439 , n40438 );
or ( n40440 , n33196 , n28146 );
nand ( n40441 , n28146 , n18435 );
nand ( n40442 , n40440 , n40441 );
buf ( n40443 , n40442 );
buf ( n40444 , n40443 );
not ( n40445 , n275929 );
buf ( n40446 , n40445 );
buf ( n40447 , n40446 );
buf ( n40448 , n275554 );
not ( n40449 , n29395 );
or ( n40450 , n40449 , n21770 );
nand ( n40451 , n21774 , n9535 );
nand ( n40452 , n40450 , n40451 );
buf ( n40453 , n40452 );
buf ( n40454 , n40453 );
not ( n40455 , n34302 );
not ( n40456 , n37066 );
or ( n40457 , n40455 , n40456 );
and ( n40458 , n37079 , n35900 );
nand ( n40459 , n37083 , n34307 );
nand ( n40460 , n28451 , n278022 );
and ( n40461 , n32755 , n12288 );
or ( n40462 , n32757 , n12296 );
nand ( n40463 , n20649 , n9323 );
nand ( n40464 , n40462 , n40463 );
nor ( n40465 , n40461 , n40464 );
nand ( n40466 , n40459 , n40460 , n40465 );
nor ( n40467 , n40458 , n40466 );
nand ( n40468 , n40457 , n40467 );
buf ( n40469 , n40468 );
buf ( n40470 , n40469 );
nand ( n40471 , n30713 , n28306 );
nand ( n40472 , n30732 , n33875 );
and ( n40473 , n28332 , n30741 );
and ( n40474 , n28350 , n11953 );
nor ( n40475 , n40473 , n40474 );
and ( n40476 , n32054 , n12255 );
or ( n40477 , n28354 , n11473 );
not ( n40478 , n11464 );
nand ( n40479 , n28357 , n40478 );
nand ( n40480 , n40477 , n40479 );
nor ( n40481 , n40476 , n40480 );
nand ( n40482 , n40471 , n40472 , n40475 , n40481 );
buf ( n40483 , n40482 );
buf ( n40484 , n40483 );
nand ( n40485 , n28303 , n23603 );
nand ( n40486 , n28326 , n23655 );
and ( n40487 , n28348 , n29371 );
or ( n40488 , n23675 , n12244 );
or ( n40489 , n23680 , n12360 );
nand ( n40490 , n40488 , n40489 );
nor ( n40491 , n40487 , n40490 );
and ( n40492 , n40485 , n40486 , n40491 );
or ( n40493 , n40492 , n27179 );
nand ( n40494 , n23708 , n11415 );
nand ( n40495 , n40493 , n40494 );
buf ( n40496 , n40495 );
buf ( n40497 , n40496 );
or ( n40498 , n25031 , n21696 );
not ( n40499 , n27647 );
or ( n40500 , n40499 , n14671 );
nand ( n40501 , n40498 , n40500 );
buf ( n40502 , n40501 );
buf ( n40503 , n40502 );
not ( n40504 , n275929 );
buf ( n40505 , n40504 );
buf ( n40506 , n40505 );
buf ( n40507 , n275554 );
not ( n40508 , n275550 );
buf ( n40509 , n40508 );
buf ( n40510 , n40509 );
nand ( n40511 , n27265 , n33875 );
nand ( n40512 , n27488 , n28306 );
and ( n40513 , n28332 , n27518 );
and ( n40514 , n28242 , n12290 );
nor ( n40515 , n40513 , n40514 );
not ( n40516 , n12174 );
and ( n40517 , n28231 , n40516 );
or ( n40518 , n31453 , n278058 );
nand ( n40519 , n28236 , n10624 );
nand ( n40520 , n40518 , n40519 );
nor ( n40521 , n40517 , n40520 );
nand ( n40522 , n40511 , n40512 , n40515 , n40521 );
buf ( n40523 , n40522 );
buf ( n40524 , n40523 );
not ( n40525 , n275550 );
buf ( n40526 , n40525 );
buf ( n40527 , n40526 );
or ( n40528 , n37574 , n19216 );
and ( n40529 , n37625 , n19360 );
not ( n40530 , n19317 );
and ( n40531 , n29479 , n25713 );
not ( n40532 , n29479 );
and ( n40533 , n40532 , n18697 );
nor ( n40534 , n40531 , n40533 );
not ( n40535 , n40534 );
and ( n40536 , n40530 , n40535 );
and ( n40537 , n19221 , n37641 );
nor ( n40538 , n40536 , n40537 );
nand ( n40539 , n37636 , n29075 );
nand ( n40540 , n19387 , n18701 );
nand ( n40541 , n40538 , n40539 , n40540 );
nor ( n40542 , n40529 , n40541 );
nand ( n40543 , n37602 , n19354 );
and ( n40544 , n40542 , n40543 );
nand ( n40545 , n40528 , n40544 );
buf ( n40546 , n40545 );
buf ( n40547 , n40546 );
not ( n40548 , n275929 );
buf ( n40549 , n40548 );
buf ( n40550 , n40549 );
buf ( n40551 , n275554 );
nand ( n40552 , n28186 , n29216 );
nand ( n40553 , n28196 , n29205 );
and ( n40554 , n40552 , n40553 );
nand ( n40555 , n28219 , n29231 );
and ( n40556 , n28231 , n12142 );
not ( n40557 , n11126 );
or ( n40558 , n28233 , n40557 );
nand ( n40559 , n28236 , n11137 );
nand ( n40560 , n40558 , n40559 );
nor ( n40561 , n40556 , n40560 );
nand ( n40562 , n28242 , n12280 );
nand ( n40563 , n40554 , n40555 , n40561 , n40562 );
buf ( n40564 , n40563 );
buf ( n40565 , n40564 );
buf ( n40566 , n275554 );
not ( n40567 , n275925 );
buf ( n40568 , n40567 );
buf ( n40569 , n40568 );
not ( n40570 , n11514 );
or ( n40571 , n40570 , n9158 );
or ( n40572 , n39986 , n9157 );
nand ( n40573 , n40571 , n40572 );
buf ( n40574 , n40573 );
buf ( n40575 , n40574 );
not ( n40576 , n35072 );
or ( n40577 , n37836 , n40576 );
or ( n40578 , n22192 , n277568 );
nand ( n40579 , n40577 , n40578 );
buf ( n40580 , n40579 );
buf ( n40581 , n40580 );
or ( n40582 , n32627 , n20743 );
and ( n40583 , n32679 , n20763 );
not ( n40584 , n35987 );
not ( n40585 , n20765 );
and ( n40586 , n40584 , n40585 );
and ( n40587 , n17411 , n32689 );
nor ( n40588 , n40586 , n40587 );
nand ( n40589 , n20785 , n32694 );
nand ( n40590 , n17560 , n13806 );
nand ( n40591 , n40588 , n40589 , n40590 );
nor ( n40592 , n40583 , n40591 );
nand ( n40593 , n32653 , n16968 );
and ( n40594 , n40592 , n40593 );
nand ( n40595 , n40582 , n40594 );
buf ( n40596 , n40595 );
buf ( n40597 , n40596 );
not ( n40598 , n275929 );
buf ( n40599 , n40598 );
buf ( n40600 , n40599 );
buf ( n40601 , n275554 );
buf ( n40602 , n275554 );
buf ( n40603 , n275554 );
not ( n40604 , n275550 );
buf ( n40605 , n40604 );
buf ( n40606 , n40605 );
buf ( n40607 , n275554 );
not ( n40608 , n275929 );
buf ( n40609 , n40608 );
buf ( n40610 , n40609 );
buf ( n40611 , n275554 );
not ( n40612 , n275550 );
buf ( n40613 , n40612 );
buf ( n40614 , n40613 );
or ( n40615 , n35718 , n24450 );
nand ( n40616 , n24450 , n18350 );
nand ( n40617 , n40615 , n40616 );
buf ( n40618 , n40617 );
buf ( n40619 , n40618 );
not ( n40620 , n20673 );
not ( n40621 , n14895 );
and ( n40622 , n40620 , n40621 );
not ( n40623 , n20687 );
not ( n40624 , n24711 );
or ( n40625 , n40623 , n40624 );
nand ( n40626 , n20939 , n17408 );
and ( n40627 , n40626 , n20680 );
and ( n40628 , n20697 , n20889 );
nor ( n40629 , n40627 , n40628 );
nand ( n40630 , n40625 , n40629 );
nor ( n40631 , n40622 , n40630 );
or ( n40632 , n40631 , n21696 );
nand ( n40633 , n21696 , n14770 );
nand ( n40634 , n40632 , n40633 );
buf ( n40635 , n40634 );
buf ( n40636 , n40635 );
buf ( n40637 , n275554 );
not ( n40638 , n275929 );
buf ( n40639 , n40638 );
buf ( n40640 , n40639 );
or ( n40641 , n30668 , n21030 );
nand ( n40642 , n21030 , n18982 );
nand ( n40643 , n40641 , n40642 );
buf ( n40644 , n40643 );
buf ( n40645 , n40644 );
nand ( n40646 , n33596 , n31422 );
nand ( n40647 , n33611 , n31437 );
nand ( n40648 , n33621 , n31449 );
and ( n40649 , n28231 , n12302 );
not ( n40650 , n277672 );
not ( n40651 , n28357 );
or ( n40652 , n40650 , n40651 );
or ( n40653 , n32061 , n277662 );
nand ( n40654 , n40652 , n40653 );
nor ( n40655 , n40649 , n40654 );
nand ( n40656 , n31460 , n277696 );
and ( n40657 , n40648 , n40655 , n40656 );
nand ( n40658 , n40646 , n40647 , n40657 );
buf ( n40659 , n40658 );
buf ( n40660 , n40659 );
not ( n40661 , n39469 );
and ( n40662 , n28328 , n40661 );
or ( n40663 , n28233 , n11039 );
nand ( n40664 , n28236 , n11034 );
nand ( n40665 , n40663 , n40664 );
nor ( n40666 , n40662 , n40665 );
not ( n40667 , n40219 );
nand ( n40668 , n37665 , n40667 );
nand ( n40669 , n37661 , n39463 );
nand ( n40670 , n31459 , n12316 );
nand ( n40671 , n40666 , n40668 , n40669 , n40670 );
buf ( n40672 , n40671 );
buf ( n40673 , n40672 );
not ( n40674 , n11613 );
not ( n40675 , n31719 );
or ( n40676 , n40674 , n40675 );
nand ( n40677 , n34055 , n27489 );
nand ( n40678 , n34063 , n27266 );
and ( n40679 , n34073 , n22052 );
or ( n40680 , n22008 , n12136 );
or ( n40681 , n23680 , n35904 );
nand ( n40682 , n40680 , n40681 );
nor ( n40683 , n40679 , n40682 );
and ( n40684 , n40677 , n40678 , n40683 );
or ( n40685 , n40684 , n29379 );
nand ( n40686 , n40676 , n40685 );
buf ( n40687 , n40686 );
buf ( n40688 , n40687 );
not ( n40689 , n275925 );
buf ( n40690 , n40689 );
buf ( n40691 , n40690 );
not ( n40692 , n275929 );
buf ( n40693 , n40692 );
buf ( n40694 , n40693 );
not ( n40695 , n275925 );
buf ( n40696 , n40695 );
buf ( n40697 , n40696 );
and ( n40698 , n14830 , n38188 );
not ( n40699 , n14830 );
and ( n40700 , n40699 , n15610 );
or ( n40701 , n40698 , n40700 );
buf ( n40702 , n40701 );
buf ( n40703 , n40702 );
or ( n40704 , n22877 , n24452 );
nand ( n40705 , n24450 , n18891 );
nand ( n40706 , n40704 , n40705 );
buf ( n40707 , n40706 );
buf ( n40708 , n40707 );
or ( n40709 , n34517 , n21697 );
nand ( n40710 , n34674 , n14658 );
nand ( n40711 , n40709 , n40710 );
buf ( n40712 , n40711 );
buf ( n40713 , n40712 );
buf ( n40714 , n33407 );
buf ( n40715 , n33455 );
nand ( n40716 , n40714 , n40715 );
buf ( n40717 , n40716 );
buf ( n40718 , n40717 );
not ( n40719 , n40718 );
buf ( n40720 , n33400 );
not ( n40721 , n40720 );
buf ( n40722 , n31838 );
nor ( n40723 , n40721 , n40722 );
buf ( n40724 , n40723 );
buf ( n40725 , n40724 );
not ( n40726 , n40725 );
buf ( n40727 , n27479 );
not ( n40728 , n40727 );
or ( n40729 , n40726 , n40728 );
buf ( n40730 , n33400 );
not ( n40731 , n40730 );
buf ( n40732 , n31922 );
not ( n40733 , n40732 );
or ( n40734 , n40731 , n40733 );
buf ( n40735 , n33448 );
not ( n40736 , n40735 );
buf ( n40737 , n40736 );
buf ( n40738 , n40737 );
nand ( n40739 , n40734 , n40738 );
buf ( n40740 , n40739 );
buf ( n40741 , n40740 );
not ( n40742 , n40741 );
buf ( n40743 , n40742 );
buf ( n40744 , n40743 );
nand ( n40745 , n40729 , n40744 );
buf ( n40746 , n40745 );
buf ( n40747 , n40746 );
not ( n40748 , n40747 );
or ( n40749 , n40719 , n40748 );
buf ( n40750 , n40746 );
buf ( n40751 , n40717 );
or ( n40752 , n40750 , n40751 );
nand ( n40753 , n40749 , n40752 );
buf ( n40754 , n40753 );
buf ( n40755 , n40754 );
nand ( n40756 , n40755 , n31422 );
nand ( n40757 , n33336 , n33360 );
not ( n40758 , n40757 );
and ( n40759 , n31978 , n33332 );
not ( n40760 , n40759 );
not ( n40761 , n27260 );
or ( n40762 , n40760 , n40761 );
not ( n40763 , n33332 );
not ( n40764 , n32011 );
or ( n40765 , n40763 , n40764 );
not ( n40766 , n33356 );
nand ( n40767 , n40765 , n40766 );
not ( n40768 , n40767 );
nand ( n40769 , n40762 , n40768 );
not ( n40770 , n40769 );
or ( n40771 , n40758 , n40770 );
or ( n40772 , n40769 , n40757 );
nand ( n40773 , n40771 , n40772 );
buf ( n40774 , n40773 );
nand ( n40775 , n40774 , n31437 );
not ( n40776 , n32790 );
not ( n40777 , n40776 );
not ( n40778 , n34839 );
nand ( n40779 , n32045 , n32032 );
nor ( n40780 , n40778 , n40779 );
not ( n40781 , n40780 );
or ( n40782 , n40777 , n40781 );
or ( n40783 , n40780 , n40776 );
nand ( n40784 , n40782 , n40783 );
buf ( n40785 , n40784 );
nand ( n40786 , n40785 , n28332 );
buf ( n40787 , n12168 );
and ( n40788 , n32054 , n40787 );
not ( n40789 , n277362 );
not ( n40790 , n28357 );
or ( n40791 , n40789 , n40790 );
or ( n40792 , n32061 , n277368 );
nand ( n40793 , n40791 , n40792 );
nor ( n40794 , n40788 , n40793 );
nand ( n40795 , n31460 , n277411 );
and ( n40796 , n40786 , n40794 , n40795 );
nand ( n40797 , n40756 , n40775 , n40796 );
buf ( n40798 , n40797 );
buf ( n40799 , n40798 );
buf ( n40800 , n275554 );
not ( n40801 , n11674 );
or ( n40802 , n40801 , n9158 );
not ( n40803 , n36064 );
or ( n40804 , n40803 , n9157 );
nand ( n40805 , n40802 , n40804 );
buf ( n40806 , n40805 );
buf ( n40807 , n40806 );
buf ( n40808 , n275554 );
not ( n40809 , n35975 );
not ( n40810 , n277355 );
not ( n40811 , n32813 );
or ( n40812 , n40810 , n40811 );
nand ( n40813 , n40812 , n32832 );
nand ( n40814 , n40809 , n40813 );
or ( n40815 , n32828 , n40814 );
not ( n40816 , n40809 );
nand ( n40817 , n40816 , n9262 );
nand ( n40818 , n40815 , n40817 );
buf ( n40819 , n40818 );
buf ( n40820 , n40819 );
buf ( n40821 , n275554 );
not ( n40822 , n275842 );
nor ( n40823 , n40822 , n275833 );
not ( n40824 , n40823 );
not ( n40825 , n275807 );
nor ( n40826 , n40825 , n275840 );
not ( n40827 , n40826 );
or ( n40828 , n40824 , n40827 );
or ( n40829 , n40826 , n40823 );
nand ( n40830 , n40828 , n40829 );
buf ( n40831 , n40830 );
buf ( n40832 , n40831 );
or ( n40833 , n35412 , n19216 );
nand ( n40834 , n35431 , n33157 );
nand ( n40835 , n35453 , n19360 );
nand ( n40836 , n35467 , n29075 );
and ( n40837 , n30146 , n30147 );
not ( n40838 , n30146 );
and ( n40839 , n40838 , n18487 );
nor ( n40840 , n40837 , n40839 );
nand ( n40841 , n40840 , n19318 );
nand ( n40842 , n33162 , n30019 );
nand ( n40843 , n19387 , n18478 );
and ( n40844 , n40836 , n40841 , n40842 , n40843 );
and ( n40845 , n40834 , n40835 , n40844 );
nand ( n40846 , n40833 , n40845 );
buf ( n40847 , n40846 );
buf ( n40848 , n40847 );
not ( n40849 , n275925 );
buf ( n40850 , n40849 );
buf ( n40851 , n40850 );
buf ( n40852 , n275554 );
not ( n40853 , n275929 );
buf ( n40854 , n40853 );
buf ( n40855 , n40854 );
not ( n40856 , n275925 );
buf ( n40857 , n40856 );
buf ( n40858 , n40857 );
buf ( n40859 , n275554 );
not ( n40860 , n275550 );
buf ( n40861 , n40860 );
buf ( n40862 , n40861 );
buf ( n40863 , n275554 );
not ( n40864 , n275550 );
buf ( n40865 , n40864 );
buf ( n40866 , n40865 );
buf ( n40867 , n275554 );
not ( n40868 , n275929 );
buf ( n40869 , n40868 );
buf ( n40870 , n40869 );
not ( n40871 , n275929 );
buf ( n40872 , n40871 );
buf ( n40873 , n40872 );
not ( n40874 , n275925 );
buf ( n40875 , n40874 );
buf ( n40876 , n40875 );
or ( n40877 , n24683 , n14909 );
and ( n40878 , n17505 , n17506 );
not ( n40879 , n17505 );
and ( n40880 , n40879 , n13593 );
nor ( n40881 , n40878 , n40880 );
not ( n40882 , n40881 );
not ( n40883 , n17545 );
or ( n40884 , n40882 , n40883 );
not ( n40885 , n24720 );
or ( n40886 , n17410 , n40885 );
nand ( n40887 , n40884 , n40886 );
not ( n40888 , n24724 );
nor ( n40889 , n40888 , n17500 );
nor ( n40890 , n40887 , n40889 );
and ( n40891 , n24696 , n16968 );
not ( n40892 , n13584 );
nor ( n40893 , n17561 , n40892 );
nor ( n40894 , n40891 , n40893 );
nand ( n40895 , n24710 , n17405 );
and ( n40896 , n40890 , n40894 , n40895 );
nand ( n40897 , n40877 , n40896 );
buf ( n40898 , n40897 );
buf ( n40899 , n40898 );
not ( n40900 , n275925 );
buf ( n40901 , n40900 );
buf ( n40902 , n40901 );
buf ( n40903 , n275554 );
not ( n40904 , n275925 );
buf ( n40905 , n40904 );
buf ( n40906 , n40905 );
not ( n40907 , n18309 );
or ( n40908 , n21769 , n40907 );
not ( n40909 , n9439 );
or ( n40910 , n21772 , n40909 );
nand ( n40911 , n40908 , n40910 );
buf ( n40912 , n40911 );
buf ( n40913 , n40912 );
not ( n40914 , n275925 );
buf ( n40915 , n40914 );
buf ( n40916 , n40915 );
not ( n40917 , n275550 );
buf ( n40918 , n40917 );
buf ( n40919 , n40918 );
buf ( n40920 , n275554 );
not ( n40921 , n275929 );
buf ( n40922 , n40921 );
buf ( n40923 , n40922 );
not ( n40924 , n35121 );
or ( n40925 , n40924 , n21770 );
nand ( n40926 , n21774 , n9500 );
nand ( n40927 , n40925 , n40926 );
buf ( n40928 , n40927 );
buf ( n40929 , n40928 );
not ( n40930 , n33715 );
not ( n40931 , n29825 );
nand ( n40932 , n40931 , n34122 );
not ( n40933 , n40932 );
not ( n40934 , n40933 );
or ( n40935 , n40930 , n40934 );
buf ( n40936 , n34155 );
nand ( n40937 , n40935 , n40936 );
nor ( n40938 , n40932 , n34155 );
nand ( n40939 , n40938 , n33715 );
nand ( n40940 , n40937 , n40939 );
buf ( n40941 , n40940 );
and ( n40942 , n40941 , n34172 );
not ( n40943 , n29856 );
nor ( n40944 , n40943 , n33056 );
nor ( n40945 , n40942 , n40944 );
not ( n40946 , n40945 );
and ( n40947 , n40946 , n23992 );
not ( n40948 , n21001 );
buf ( n40949 , n34248 );
not ( n40950 , n40949 );
buf ( n40951 , n18463 );
buf ( n40952 , n40951 );
buf ( n40953 , n40952 );
not ( n40954 , n40953 );
or ( n40955 , n40950 , n40954 );
or ( n40956 , n40953 , n40949 );
nand ( n40957 , n40955 , n40956 );
not ( n40958 , n40957 );
and ( n40959 , n29966 , n29969 );
not ( n40960 , n40959 );
or ( n40961 , n40958 , n40960 );
or ( n40962 , n40959 , n40957 );
nand ( n40963 , n40961 , n40962 );
not ( n40964 , n40963 );
nand ( n40965 , n30039 , n29971 );
nor ( n40966 , n40965 , n28014 );
not ( n40967 , n40966 );
not ( n40968 , n30043 );
or ( n40969 , n40967 , n40968 );
not ( n40970 , n40965 );
and ( n40971 , n28036 , n40970 );
not ( n40972 , n29971 );
not ( n40973 , n30063 );
or ( n40974 , n40972 , n40973 );
nand ( n40975 , n40974 , n29972 );
nor ( n40976 , n40971 , n40975 );
nand ( n40977 , n40969 , n40976 );
not ( n40978 , n40977 );
or ( n40979 , n40964 , n40978 );
or ( n40980 , n40977 , n40963 );
nand ( n40981 , n40979 , n40980 );
buf ( n40982 , n40981 );
not ( n40983 , n40982 );
or ( n40984 , n40948 , n40983 );
buf ( n40985 , n34248 );
not ( n40986 , n40985 );
buf ( n40987 , n40952 );
not ( n40988 , n40987 );
not ( n40989 , n40988 );
or ( n40990 , n40986 , n40989 );
or ( n40991 , n40988 , n40985 );
nand ( n40992 , n40990 , n40991 );
not ( n40993 , n40992 );
and ( n40994 , n30073 , n30074 );
not ( n40995 , n40994 );
or ( n40996 , n40993 , n40995 );
or ( n40997 , n40994 , n40992 );
nand ( n40998 , n40996 , n40997 );
not ( n40999 , n40998 );
nand ( n41000 , n30102 , n30081 );
nor ( n41001 , n41000 , n28079 );
not ( n41002 , n41001 );
not ( n41003 , n28092 );
or ( n41004 , n41002 , n41003 );
not ( n41005 , n33731 );
not ( n41006 , n41000 );
and ( n41007 , n41005 , n41006 );
not ( n41008 , n30081 );
not ( n41009 , n30122 );
or ( n41010 , n41008 , n41009 );
nand ( n41011 , n41010 , n30082 );
nor ( n41012 , n41007 , n41011 );
nand ( n41013 , n41004 , n41012 );
not ( n41014 , n41013 );
or ( n41015 , n40999 , n41014 );
or ( n41016 , n41013 , n40998 );
nand ( n41017 , n41015 , n41016 );
buf ( n41018 , n41017 );
and ( n41019 , n41018 , n19358 );
not ( n41020 , n19290 );
not ( n41021 , n34251 );
nor ( n41022 , n30166 , n30156 );
nand ( n41023 , n30160 , n41022 );
nor ( n41024 , n28124 , n41023 );
not ( n41025 , n41024 );
or ( n41026 , n41021 , n41025 );
or ( n41027 , n41024 , n34251 );
nand ( n41028 , n41026 , n41027 );
buf ( n41029 , n41028 );
not ( n41030 , n41029 );
or ( n41031 , n41020 , n41030 );
not ( n41032 , n34249 );
buf ( n41033 , n41032 );
buf ( n41034 , n41033 );
nand ( n41035 , n19219 , n41034 );
nand ( n41036 , n41031 , n41035 );
nor ( n41037 , n41019 , n41036 );
nand ( n41038 , n40984 , n41037 );
nor ( n41039 , n40947 , n41038 );
or ( n41040 , n41039 , n21030 );
nand ( n41041 , n21030 , n18450 );
nand ( n41042 , n41040 , n41041 );
buf ( n41043 , n41042 );
buf ( n41044 , n41043 );
not ( n41045 , n275929 );
buf ( n41046 , n41045 );
buf ( n41047 , n41046 );
not ( n41048 , n275925 );
buf ( n41049 , n41048 );
buf ( n41050 , n41049 );
not ( n41051 , n275550 );
buf ( n41052 , n41051 );
buf ( n41053 , n41052 );
not ( n41054 , n275550 );
buf ( n41055 , n41054 );
buf ( n41056 , n41055 );
buf ( n41057 , n275554 );
buf ( n41058 , n275554 );
buf ( n41059 , n275554 );
not ( n41060 , n9158 );
not ( n41061 , n9061 );
or ( n41062 , n41060 , n41061 );
not ( n41063 , n277410 );
or ( n41064 , n41063 , n9158 );
nand ( n41065 , n41062 , n41064 );
buf ( n41066 , n41065 );
buf ( n41067 , n41066 );
buf ( n41068 , n275554 );
not ( n41069 , n39249 );
and ( n41070 , n41069 , n21174 );
not ( n41071 , n21001 );
not ( n41072 , n39268 );
or ( n41073 , n41071 , n41072 );
and ( n41074 , n39284 , n19358 );
not ( n41075 , n19290 );
not ( n41076 , n39304 );
or ( n41077 , n41075 , n41076 );
nand ( n41078 , n27619 , n39294 );
nand ( n41079 , n41077 , n41078 );
nor ( n41080 , n41074 , n41079 );
nand ( n41081 , n41073 , n41080 );
nor ( n41082 , n41070 , n41081 );
or ( n41083 , n41082 , n21030 );
nand ( n41084 , n21030 , n18747 );
nand ( n41085 , n41083 , n41084 );
buf ( n41086 , n41085 );
buf ( n41087 , n41086 );
buf ( n41088 , n275554 );
buf ( n41089 , n275554 );
and ( n41090 , n37271 , n275783 );
not ( n41091 , n32968 );
nand ( n41092 , n41091 , n29263 );
nor ( n41093 , n41090 , n41092 );
nand ( n41094 , n22914 , n22969 );
buf ( n41095 , n22975 );
not ( n41096 , n41095 );
buf ( n41097 , n22993 );
nor ( n41098 , n41096 , n41097 );
buf ( n41099 , n41098 );
buf ( n41100 , n41099 );
not ( n41101 , n41100 );
buf ( n41102 , n35600 );
not ( n41103 , n41102 );
or ( n41104 , n41101 , n41103 );
buf ( n41105 , n35600 );
buf ( n41106 , n41099 );
or ( n41107 , n41105 , n41106 );
nand ( n41108 , n41104 , n41107 );
buf ( n41109 , n41108 );
buf ( n41110 , n41109 );
nand ( n41111 , n22918 , n41110 );
buf ( n41112 , n23205 );
not ( n41113 , n41112 );
buf ( n41114 , n23223 );
nor ( n41115 , n41113 , n41114 );
buf ( n41116 , n41115 );
buf ( n41117 , n41116 );
not ( n41118 , n41117 );
buf ( n41119 , n35627 );
not ( n41120 , n41119 );
or ( n41121 , n41118 , n41120 );
buf ( n41122 , n35627 );
buf ( n41123 , n41116 );
or ( n41124 , n41122 , n41123 );
nand ( n41125 , n41121 , n41124 );
buf ( n41126 , n41125 );
buf ( n41127 , n41126 );
nand ( n41128 , n23152 , n41127 );
nand ( n41129 , n41093 , n41094 , n41111 , n41128 );
buf ( n41130 , n41129 );
buf ( n41131 , n41130 );
buf ( n41132 , n275554 );
or ( n41133 , n19102 , n19634 );
and ( n41134 , n34105 , n19088 );
and ( n41135 , n20353 , n19347 );
and ( n41136 , n19645 , n19311 );
nor ( n41137 , n41135 , n41136 );
nand ( n41138 , n19644 , n19286 );
nand ( n41139 , n20515 , n19372 );
nand ( n41140 , n41137 , n41138 , n41139 );
nor ( n41141 , n41134 , n41140 );
nand ( n41142 , n41133 , n41141 );
buf ( n41143 , n41142 );
buf ( n41144 , n41143 );
buf ( n41145 , n275554 );
or ( n41146 , n39091 , n21697 );
nand ( n41147 , n27647 , n14705 );
nand ( n41148 , n41146 , n41147 );
buf ( n41149 , n41148 );
buf ( n41150 , n41149 );
buf ( n41151 , n275554 );
not ( n41152 , n22335 );
not ( n41153 , n25087 );
or ( n41154 , n41152 , n41153 );
not ( n41155 , n21403 );
or ( n41156 , n41155 , n22335 );
nand ( n41157 , n41154 , n41156 );
buf ( n41158 , n41157 );
buf ( n41159 , n41158 );
buf ( n41160 , n275554 );
and ( n41161 , n19387 , n19047 );
not ( n41162 , n19387 );
and ( n41163 , n41162 , n34263 );
or ( n41164 , n41161 , n41163 );
buf ( n41165 , n41164 );
buf ( n41166 , n41165 );
or ( n41167 , n27112 , n26364 );
nand ( n41168 , n27131 , n26370 );
nand ( n41169 , n27149 , n26374 );
nand ( n41170 , n32176 , n35232 );
nand ( n41171 , n27157 , n26393 );
nand ( n41172 , n26395 , n27161 );
not ( n41173 , n33636 );
and ( n41174 , n41171 , n41172 , n41173 );
and ( n41175 , n41168 , n41169 , n41170 , n41174 );
nand ( n41176 , n41167 , n41175 );
buf ( n41177 , n41176 );
buf ( n41178 , n41177 );
not ( n41179 , n275925 );
buf ( n41180 , n41179 );
buf ( n41181 , n41180 );
not ( n41182 , n275925 );
buf ( n41183 , n41182 );
buf ( n41184 , n41183 );
buf ( n41185 , n275554 );
not ( n41186 , n275550 );
buf ( n41187 , n41186 );
buf ( n41188 , n41187 );
not ( n41189 , n275550 );
buf ( n41190 , n41189 );
buf ( n41191 , n41190 );
not ( n41192 , n275925 );
buf ( n41193 , n41192 );
buf ( n41194 , n41193 );
or ( n41195 , n35134 , n32073 );
and ( n41196 , n35166 , n20353 );
or ( n41197 , n20562 , n35189 );
or ( n41198 , n20559 , n35183 );
nor ( n41199 , n19639 , n19655 );
not ( n41200 , n41199 );
nand ( n41201 , n41197 , n41198 , n41200 );
nor ( n41202 , n41196 , n41201 );
nand ( n41203 , n35145 , n20515 );
nand ( n41204 , n19650 , n35173 );
and ( n41205 , n41202 , n41203 , n41204 );
nand ( n41206 , n41195 , n41205 );
buf ( n41207 , n41206 );
buf ( n41208 , n41207 );
not ( n41209 , n275929 );
buf ( n41210 , n41209 );
buf ( n41211 , n41210 );
not ( n41212 , n29820 );
or ( n41213 , n41212 , n21774 );
nand ( n41214 , n21770 , n9779 );
nand ( n41215 , n41213 , n41214 );
buf ( n41216 , n41215 );
buf ( n41217 , n41216 );
buf ( n41218 , n275554 );
and ( n41219 , n24450 , n19050 );
not ( n41220 , n24450 );
and ( n41221 , n41220 , n34263 );
or ( n41222 , n41219 , n41221 );
buf ( n41223 , n41222 );
buf ( n41224 , n41223 );
not ( n41225 , n275929 );
buf ( n41226 , n41225 );
buf ( n41227 , n41226 );
and ( n41228 , n22335 , n25067 );
not ( n41229 , n22335 );
and ( n41230 , n41229 , n24153 );
or ( n41231 , n41228 , n41230 );
buf ( n41232 , n41231 );
buf ( n41233 , n41232 );
buf ( n41234 , n275554 );
buf ( n41235 , n275554 );
buf ( n41236 , n275554 );
not ( n41237 , n13358 );
not ( n41238 , n27665 );
or ( n41239 , n41237 , n41238 );
not ( n41240 , n24889 );
or ( n41241 , n41240 , n27665 );
nand ( n41242 , n41239 , n41241 );
buf ( n41243 , n41242 );
buf ( n41244 , n41243 );
not ( n41245 , n275929 );
buf ( n41246 , n41245 );
buf ( n41247 , n41246 );
buf ( n41248 , n275554 );
not ( n41249 , n275925 );
buf ( n41250 , n41249 );
buf ( n41251 , n41250 );
not ( n41252 , n275925 );
buf ( n41253 , n41252 );
buf ( n41254 , n41253 );
or ( n41255 , n26438 , n20743 );
nand ( n41256 , n26462 , n16970 );
nand ( n41257 , n26483 , n17405 );
nand ( n41258 , n32339 , n26493 );
nand ( n41259 , n20785 , n26498 );
nand ( n41260 , n17562 , n13695 );
and ( n41261 , n17516 , n13699 );
not ( n41262 , n17516 );
not ( n41263 , n13698 );
and ( n41264 , n41262 , n41263 );
nor ( n41265 , n41261 , n41264 );
nand ( n41266 , n17545 , n41265 );
and ( n41267 , n41258 , n41259 , n41260 , n41266 );
and ( n41268 , n41256 , n41257 , n41267 );
nand ( n41269 , n41255 , n41268 );
buf ( n41270 , n41269 );
buf ( n41271 , n41270 );
buf ( n41272 , n275554 );
buf ( n41273 , n275554 );
buf ( n41274 , n275554 );
not ( n41275 , n275929 );
buf ( n41276 , n41275 );
buf ( n41277 , n41276 );
buf ( n41278 , n275554 );
and ( n41279 , n23706 , n277658 );
not ( n41280 , n23706 );
and ( n41281 , n41280 , n33629 );
or ( n41282 , n41279 , n41281 );
buf ( n41283 , n41282 );
buf ( n41284 , n41283 );
buf ( n41285 , n275554 );
buf ( n41286 , n275554 );
buf ( n41287 , n275554 );
buf ( n41288 , n275554 );
not ( n41289 , n275925 );
buf ( n41290 , n41289 );
buf ( n41291 , n41290 );
or ( n41292 , n41039 , n24452 );
nand ( n41293 , n24450 , n18461 );
nand ( n41294 , n41292 , n41293 );
buf ( n41295 , n41294 );
buf ( n41296 , n41295 );
buf ( n41297 , n275554 );
not ( n41298 , n275925 );
buf ( n41299 , n41298 );
buf ( n41300 , n41299 );
or ( n41301 , n24494 , n14909 );
nand ( n41302 , n24574 , n16970 );
and ( n41303 , n24607 , n17405 );
nand ( n41304 , n17411 , n24617 );
nand ( n41305 , n20785 , n24538 );
nand ( n41306 , n38340 , n17545 );
nand ( n41307 , n17562 , n14029 );
nand ( n41308 , n41304 , n41305 , n41306 , n41307 );
nor ( n41309 , n41303 , n41308 );
and ( n41310 , n41302 , n41309 );
nand ( n41311 , n41301 , n41310 );
buf ( n41312 , n41311 );
buf ( n41313 , n41312 );
not ( n41314 , n275550 );
buf ( n41315 , n41314 );
buf ( n41316 , n41315 );
buf ( n41317 , n275554 );
buf ( n41318 , n275554 );
not ( n41319 , n275550 );
buf ( n41320 , n41319 );
buf ( n41321 , n41320 );
not ( n41322 , n275925 );
buf ( n41323 , n41322 );
buf ( n41324 , n41323 );
not ( n41325 , n275550 );
buf ( n41326 , n41325 );
buf ( n41327 , n41326 );
not ( n41328 , n27832 );
or ( n41329 , n41328 , n21774 );
nand ( n41330 , n21774 , n9761 );
nand ( n41331 , n41329 , n41330 );
buf ( n41332 , n41331 );
buf ( n41333 , n41332 );
buf ( n41334 , n275554 );
buf ( n41335 , n275554 );
not ( n41336 , n9419 );
not ( n41337 , n9426 );
or ( n41338 , n41336 , n41337 );
not ( n41339 , n9426 );
not ( n41340 , n9419 );
and ( n41341 , n41339 , n41340 );
buf ( n41342 , RI210699c8_646);
buf ( n41343 , n41342 );
nor ( n41344 , n41341 , n41343 );
nand ( n41345 , n41338 , n41344 );
buf ( n41346 , n41345 );
buf ( n41347 , n41346 );
not ( n41348 , n34302 );
not ( n41349 , n40755 );
or ( n41350 , n41348 , n41349 );
and ( n41351 , n40774 , n28430 );
nand ( n41352 , n40785 , n34307 );
nand ( n41353 , n28451 , n277362 );
and ( n41354 , n32755 , n40787 );
and ( n41355 , n34848 , n277411 );
and ( n41356 , n34313 , n9364 );
nor ( n41357 , n41354 , n41355 , n41356 );
nand ( n41358 , n41352 , n41353 , n41357 );
nor ( n41359 , n41351 , n41358 );
nand ( n41360 , n41350 , n41359 );
buf ( n41361 , n41360 );
buf ( n41362 , n41361 );
not ( n41363 , n275929 );
buf ( n41364 , n41363 );
buf ( n41365 , n41364 );
buf ( n41366 , n275554 );
buf ( n41367 , n275554 );
not ( n41368 , n275550 );
buf ( n41369 , n41368 );
buf ( n41370 , n41369 );
not ( n41371 , n275925 );
buf ( n41372 , n41371 );
buf ( n41373 , n41372 );
not ( n41374 , n275925 );
buf ( n41375 , n41374 );
buf ( n41376 , n41375 );
buf ( n41377 , n275554 );
not ( n41378 , n275925 );
buf ( n41379 , n41378 );
buf ( n41380 , n41379 );
not ( n41381 , n275929 );
buf ( n41382 , n41381 );
buf ( n41383 , n41382 );
buf ( n41384 , n275554 );
not ( n41385 , n34245 );
nand ( n41386 , n30160 , n30167 , n34252 );
nor ( n41387 , n28124 , n41386 );
not ( n41388 , n41387 );
or ( n41389 , n41385 , n41388 );
or ( n41390 , n41387 , n34245 );
nand ( n41391 , n41389 , n41390 );
buf ( n41392 , n41391 );
and ( n41393 , n41392 , n19290 );
and ( n41394 , n19219 , n34244 );
nor ( n41395 , n41393 , n41394 );
and ( n41396 , n34174 , n41395 );
or ( n41397 , n41396 , n28146 );
or ( n41398 , n33546 , n18841 );
nand ( n41399 , n41397 , n41398 );
buf ( n41400 , n41399 );
buf ( n41401 , n41400 );
and ( n41402 , n31468 , n275596 );
nor ( n41403 , n41402 , n35760 );
nand ( n41404 , n22914 , n35108 );
buf ( n41405 , n23086 );
not ( n41406 , n41405 );
buf ( n41407 , n23123 );
nand ( n41408 , n41406 , n41407 );
buf ( n41409 , n41408 );
buf ( n41410 , n41409 );
not ( n41411 , n41410 );
buf ( n41412 , n30540 );
not ( n41413 , n41412 );
buf ( n41414 , n41413 );
buf ( n41415 , n41414 );
buf ( n41416 , n23094 );
or ( n41417 , n41415 , n41416 );
buf ( n41418 , n23117 );
nand ( n41419 , n41417 , n41418 );
buf ( n41420 , n41419 );
buf ( n41421 , n41420 );
not ( n41422 , n41421 );
or ( n41423 , n41411 , n41422 );
buf ( n41424 , n41420 );
buf ( n41425 , n41409 );
or ( n41426 , n41424 , n41425 );
nand ( n41427 , n41423 , n41426 );
buf ( n41428 , n41427 );
buf ( n41429 , n41428 );
nand ( n41430 , n22918 , n41429 );
buf ( n41431 , n23312 );
not ( n41432 , n41431 );
buf ( n41433 , n23348 );
nand ( n41434 , n41432 , n41433 );
buf ( n41435 , n41434 );
buf ( n41436 , n41435 );
not ( n41437 , n41436 );
buf ( n41438 , n30574 );
not ( n41439 , n41438 );
buf ( n41440 , n41439 );
buf ( n41441 , n41440 );
buf ( n41442 , n23319 );
or ( n41443 , n41441 , n41442 );
buf ( n41444 , n23342 );
nand ( n41445 , n41443 , n41444 );
buf ( n41446 , n41445 );
buf ( n41447 , n41446 );
not ( n41448 , n41447 );
or ( n41449 , n41437 , n41448 );
buf ( n41450 , n41446 );
buf ( n41451 , n41435 );
or ( n41452 , n41450 , n41451 );
nand ( n41453 , n41449 , n41452 );
buf ( n41454 , n41453 );
buf ( n41455 , n41454 );
nand ( n41456 , n23152 , n41455 );
nand ( n41457 , n41403 , n41404 , n41430 , n41456 );
buf ( n41458 , n41457 );
buf ( n41459 , n41458 );
not ( n41460 , n275925 );
buf ( n41461 , n41460 );
buf ( n41462 , n41461 );
not ( n41463 , n275925 );
buf ( n41464 , n41463 );
buf ( n41465 , n41464 );
not ( n41466 , n277452 );
or ( n41467 , n41466 , n9158 );
nand ( n41468 , n9228 , n9158 );
nand ( n41469 , n41467 , n41468 );
buf ( n41470 , n41469 );
buf ( n41471 , n41470 );
or ( n41472 , n30610 , n19216 );
and ( n41473 , n30624 , n19354 );
not ( n41474 , n30628 );
not ( n41475 , n33162 );
or ( n41476 , n41474 , n41475 );
not ( n41477 , n19291 );
not ( n41478 , n30636 );
and ( n41479 , n41477 , n41478 );
and ( n41480 , n19318 , n30617 );
nor ( n41481 , n41479 , n41480 );
nand ( n41482 , n41476 , n41481 );
nor ( n41483 , n41473 , n41482 );
nand ( n41484 , n30649 , n19360 );
nand ( n41485 , n19387 , n18356 );
and ( n41486 , n41483 , n41484 , n41485 );
nand ( n41487 , n41472 , n41486 );
buf ( n41488 , n41487 );
buf ( n41489 , n41488 );
nand ( n41490 , n25064 , n28818 );
buf ( n41491 , n28533 );
buf ( n41492 , n28593 );
nor ( n41493 , n41491 , n41492 );
buf ( n41494 , n41493 );
buf ( n41495 , n41494 );
not ( n41496 , n41495 );
buf ( n41497 , n28514 );
buf ( n41498 , n28523 );
buf ( n41499 , n37131 );
and ( n41500 , n41497 , n41498 , n41499 );
buf ( n41501 , n28573 );
buf ( n41502 , n28543 );
or ( n41503 , n41501 , n41502 );
buf ( n41504 , n28586 );
nand ( n41505 , n41503 , n41504 );
buf ( n41506 , n41505 );
buf ( n41507 , n41506 );
nor ( n41508 , n41500 , n41507 );
buf ( n41509 , n41508 );
buf ( n41510 , n41509 );
not ( n41511 , n41510 );
or ( n41512 , n41496 , n41511 );
buf ( n41513 , n41509 );
buf ( n41514 , n41494 );
or ( n41515 , n41513 , n41514 );
nand ( n41516 , n41512 , n41515 );
buf ( n41517 , n41516 );
buf ( n41518 , n41517 );
not ( n41519 , n41518 );
nor ( n41520 , n41519 , n25389 );
nand ( n41521 , n25397 , n36500 );
buf ( n41522 , n28729 );
not ( n41523 , n41522 );
buf ( n41524 , n28684 );
nor ( n41525 , n41523 , n41524 );
buf ( n41526 , n41525 );
buf ( n41527 , n41526 );
not ( n41528 , n41527 );
buf ( n41529 , n28655 );
buf ( n41530 , n28667 );
buf ( n41531 , n37167 );
and ( n41532 , n41529 , n41530 , n41531 );
buf ( n41533 , n28714 );
buf ( n41534 , n28691 );
or ( n41535 , n41533 , n41534 );
buf ( n41536 , n28723 );
nand ( n41537 , n41535 , n41536 );
buf ( n41538 , n41537 );
buf ( n41539 , n41538 );
nor ( n41540 , n41532 , n41539 );
buf ( n41541 , n41540 );
buf ( n41542 , n41541 );
not ( n41543 , n41542 );
or ( n41544 , n41528 , n41543 );
buf ( n41545 , n41541 );
buf ( n41546 , n41526 );
or ( n41547 , n41545 , n41546 );
nand ( n41548 , n41544 , n41547 );
buf ( n41549 , n41548 );
buf ( n41550 , n41549 );
and ( n41551 , n25402 , n41550 );
nor ( n41552 , n41551 , n29496 );
buf ( n41553 , n28870 );
not ( n41554 , n41553 );
buf ( n41555 , n28824 );
nor ( n41556 , n41554 , n41555 );
buf ( n41557 , n41556 );
buf ( n41558 , n41557 );
not ( n41559 , n41558 );
buf ( n41560 , n28796 );
buf ( n41561 , n28808 );
buf ( n41562 , n37201 );
and ( n41563 , n41560 , n41561 , n41562 );
buf ( n41564 , n28855 );
buf ( n41565 , n28832 );
or ( n41566 , n41564 , n41565 );
buf ( n41567 , n28864 );
nand ( n41568 , n41566 , n41567 );
buf ( n41569 , n41568 );
buf ( n41570 , n41569 );
nor ( n41571 , n41563 , n41570 );
buf ( n41572 , n41571 );
buf ( n41573 , n41572 );
not ( n41574 , n41573 );
or ( n41575 , n41559 , n41574 );
buf ( n41576 , n41572 );
buf ( n41577 , n41557 );
or ( n41578 , n41576 , n41577 );
nand ( n41579 , n41575 , n41578 );
buf ( n41580 , n41579 );
buf ( n41581 , n41580 );
nand ( n41582 , n28761 , n41581 );
nand ( n41583 , n41521 , n41552 , n41582 );
nor ( n41584 , n41520 , n41583 );
buf ( n41585 , n28955 );
buf ( n41586 , n29012 );
nor ( n41587 , n41585 , n41586 );
buf ( n41588 , n41587 );
buf ( n41589 , n41588 );
not ( n41590 , n41589 );
buf ( n41591 , n28935 );
buf ( n41592 , n28947 );
buf ( n41593 , n37235 );
and ( n41594 , n41591 , n41592 , n41593 );
buf ( n41595 , n28992 );
buf ( n41596 , n28964 );
or ( n41597 , n41595 , n41596 );
buf ( n41598 , n29005 );
nand ( n41599 , n41597 , n41598 );
buf ( n41600 , n41599 );
buf ( n41601 , n41600 );
nor ( n41602 , n41594 , n41601 );
buf ( n41603 , n41602 );
buf ( n41604 , n41603 );
not ( n41605 , n41604 );
or ( n41606 , n41590 , n41605 );
buf ( n41607 , n41603 );
buf ( n41608 , n41588 );
or ( n41609 , n41607 , n41608 );
nand ( n41610 , n41606 , n41609 );
buf ( n41611 , n41610 );
buf ( n41612 , n41611 );
nand ( n41613 , n26027 , n41612 );
nand ( n41614 , n41490 , n41584 , n41613 );
buf ( n41615 , n41614 );
buf ( n41616 , n41615 );
or ( n41617 , n30495 , n31719 );
or ( n41618 , n35071 , n11268 );
nand ( n41619 , n41617 , n41618 );
buf ( n41620 , n41619 );
buf ( n41621 , n41620 );
or ( n41622 , n36036 , n40103 );
and ( n41623 , n36045 , n275711 );
not ( n41624 , n36120 );
nand ( n41625 , n36124 , n36129 );
not ( n41626 , n41625 );
or ( n41627 , n41624 , n41626 );
or ( n41628 , n41625 , n36120 );
nand ( n41629 , n41627 , n41628 );
buf ( n41630 , n41629 );
not ( n41631 , n41630 );
not ( n41632 , n36155 );
or ( n41633 , n41631 , n41632 );
not ( n41634 , n36159 );
not ( n41635 , n41634 );
not ( n41636 , n36226 );
nand ( n41637 , n36230 , n36235 );
not ( n41638 , n41637 );
or ( n41639 , n41636 , n41638 );
or ( n41640 , n41637 , n36226 );
nand ( n41641 , n41639 , n41640 );
buf ( n41642 , n41641 );
nand ( n41643 , n41635 , n41642 );
nand ( n41644 , n41633 , n41643 );
nor ( n41645 , n41623 , n41644 );
nand ( n41646 , n41622 , n41645 );
nand ( n41647 , n41646 , n20645 );
not ( n41648 , n36317 );
nand ( n41649 , n36319 , n36300 );
not ( n41650 , n41649 );
or ( n41651 , n41648 , n41650 );
or ( n41652 , n41649 , n36317 );
nand ( n41653 , n41651 , n41652 );
buf ( n41654 , n41653 );
nand ( n41655 , n36267 , n41654 );
not ( n41656 , n36420 );
not ( n41657 , n36408 );
nand ( n41658 , n36422 , n41657 );
not ( n41659 , n41658 );
or ( n41660 , n41656 , n41659 );
or ( n41661 , n41658 , n36420 );
nand ( n41662 , n41660 , n41661 );
buf ( n41663 , n41662 );
nand ( n41664 , n36371 , n41663 );
and ( n41665 , n36474 , n11144 );
not ( n41666 , n11137 );
not ( n41667 , n34313 );
or ( n41668 , n41666 , n41667 );
or ( n41669 , n20654 , n275710 );
nand ( n41670 , n41668 , n41669 );
nor ( n41671 , n41665 , n41670 );
nand ( n41672 , n41647 , n41655 , n41664 , n41671 );
buf ( n41673 , n41672 );
buf ( n41674 , n41673 );
not ( n41675 , n275929 );
buf ( n41676 , n41675 );
buf ( n41677 , n41676 );
not ( n41678 , n275929 );
buf ( n41679 , n41678 );
buf ( n41680 , n41679 );
buf ( n41681 , n275554 );
buf ( n41682 , n25639 );
buf ( n41683 , n25442 );
nand ( n41684 , n41682 , n41683 );
buf ( n41685 , n41684 );
buf ( n41686 , n41685 );
not ( n41687 , n41686 );
buf ( n41688 , n25586 );
not ( n41689 , n41688 );
buf ( n41690 , n41689 );
buf ( n41691 , n41690 );
buf ( n41692 , n25450 );
or ( n41693 , n41691 , n41692 );
buf ( n41694 , n25629 );
nand ( n41695 , n41693 , n41694 );
buf ( n41696 , n41695 );
buf ( n41697 , n41696 );
not ( n41698 , n41697 );
or ( n41699 , n41687 , n41698 );
buf ( n41700 , n41696 );
buf ( n41701 , n41685 );
or ( n41702 , n41700 , n41701 );
nand ( n41703 , n41699 , n41702 );
buf ( n41704 , n41703 );
buf ( n41705 , n41704 );
and ( n41706 , n25402 , n41705 );
nor ( n41707 , n19639 , n19659 );
nor ( n41708 , n41706 , n41707 );
nand ( n41709 , n25397 , n275600 );
buf ( n41710 , n25953 );
buf ( n41711 , n25759 );
nand ( n41712 , n41710 , n41711 );
buf ( n41713 , n41712 );
buf ( n41714 , n41713 );
not ( n41715 , n41714 );
buf ( n41716 , n25902 );
not ( n41717 , n41716 );
buf ( n41718 , n41717 );
buf ( n41719 , n41718 );
buf ( n41720 , n25767 );
or ( n41721 , n41719 , n41720 );
buf ( n41722 , n25943 );
nand ( n41723 , n41721 , n41722 );
buf ( n41724 , n41723 );
buf ( n41725 , n41724 );
not ( n41726 , n41725 );
or ( n41727 , n41715 , n41726 );
buf ( n41728 , n41724 );
buf ( n41729 , n41713 );
or ( n41730 , n41728 , n41729 );
nand ( n41731 , n41727 , n41730 );
buf ( n41732 , n41731 );
buf ( n41733 , n41732 );
nand ( n41734 , n28761 , n41733 );
nand ( n41735 , n41708 , n41709 , n41734 );
buf ( n41736 , n25115 );
buf ( n41737 , n25326 );
nand ( n41738 , n41736 , n41737 );
buf ( n41739 , n41738 );
buf ( n41740 , n41739 );
not ( n41741 , n41740 );
buf ( n41742 , n25264 );
not ( n41743 , n41742 );
buf ( n41744 , n41743 );
buf ( n41745 , n41744 );
buf ( n41746 , n25125 );
or ( n41747 , n41745 , n41746 );
buf ( n41748 , n25316 );
nand ( n41749 , n41747 , n41748 );
buf ( n41750 , n41749 );
buf ( n41751 , n41750 );
not ( n41752 , n41751 );
or ( n41753 , n41741 , n41752 );
buf ( n41754 , n41750 );
buf ( n41755 , n41739 );
or ( n41756 , n41754 , n41755 );
nand ( n41757 , n41753 , n41756 );
buf ( n41758 , n41757 );
buf ( n41759 , n41758 );
not ( n41760 , n41759 );
nor ( n41761 , n41760 , n25389 );
nor ( n41762 , n41735 , n41761 );
buf ( n41763 , n25753 );
nand ( n41764 , n25064 , n41763 );
buf ( n41765 , n26068 );
not ( n41766 , n41765 );
buf ( n41767 , n26267 );
nand ( n41768 , n41766 , n41767 );
buf ( n41769 , n41768 );
buf ( n41770 , n41769 );
not ( n41771 , n41770 );
buf ( n41772 , n26212 );
not ( n41773 , n41772 );
buf ( n41774 , n41773 );
buf ( n41775 , n41774 );
buf ( n41776 , n26075 );
or ( n41777 , n41775 , n41776 );
buf ( n41778 , n26261 );
nand ( n41779 , n41777 , n41778 );
buf ( n41780 , n41779 );
buf ( n41781 , n41780 );
not ( n41782 , n41781 );
or ( n41783 , n41771 , n41782 );
buf ( n41784 , n41780 );
buf ( n41785 , n41769 );
or ( n41786 , n41784 , n41785 );
nand ( n41787 , n41783 , n41786 );
buf ( n41788 , n41787 );
buf ( n41789 , n41788 );
nand ( n41790 , n26027 , n41789 );
nand ( n41791 , n41762 , n41764 , n41790 );
buf ( n41792 , n41791 );
buf ( n41793 , n41792 );
not ( n41794 , n275929 );
buf ( n41795 , n41794 );
buf ( n41796 , n41795 );
buf ( n41797 , n275554 );
buf ( n41798 , n275554 );
not ( n41799 , n275925 );
buf ( n41800 , n41799 );
buf ( n41801 , n41800 );
or ( n41802 , n29410 , n19636 );
not ( n41803 , n38353 );
not ( n41804 , n35950 );
and ( n41805 , n41803 , n41804 );
and ( n41806 , n29427 , n20353 );
nor ( n41807 , n41805 , n41806 );
and ( n41808 , n29444 , n20515 );
nor ( n41809 , n19639 , n29475 );
not ( n41810 , n41809 );
nand ( n41811 , n29454 , n20560 );
nand ( n41812 , n19644 , n29459 );
nand ( n41813 , n41810 , n41811 , n41812 );
nor ( n41814 , n41808 , n41813 );
and ( n41815 , n41807 , n41814 );
nand ( n41816 , n41802 , n41815 );
buf ( n41817 , n41816 );
buf ( n41818 , n41817 );
not ( n41819 , n275550 );
buf ( n41820 , n41819 );
buf ( n41821 , n41820 );
or ( n41822 , n23684 , n31719 );
or ( n41823 , n35071 , n11526 );
nand ( n41824 , n41822 , n41823 );
buf ( n41825 , n41824 );
buf ( n41826 , n41825 );
not ( n41827 , n275893 );
nand ( n41828 , n41827 , n275905 );
not ( n41829 , n41828 );
or ( n41830 , n39522 , n275900 );
nand ( n41831 , n41830 , n275903 );
not ( n41832 , n41831 );
or ( n41833 , n41829 , n41832 );
or ( n41834 , n41831 , n41828 );
nand ( n41835 , n41833 , n41834 );
buf ( n41836 , n41835 );
buf ( n41837 , n41836 );
not ( n41838 , n275929 );
buf ( n41839 , n41838 );
buf ( n41840 , n41839 );
buf ( n41841 , n275554 );
buf ( n41842 , n275554 );
or ( n41843 , n20947 , n27647 );
nand ( n41844 , n34674 , n13474 );
nand ( n41845 , n41843 , n41844 );
buf ( n41846 , n41845 );
buf ( n41847 , n41846 );
not ( n41848 , n275929 );
buf ( n41849 , n41848 );
buf ( n41850 , n41849 );
not ( n41851 , n275925 );
buf ( n41852 , n41851 );
buf ( n41853 , n41852 );
not ( n41854 , n275925 );
buf ( n41855 , n41854 );
buf ( n41856 , n41855 );
or ( n41857 , n38755 , n21030 );
nand ( n41858 , n21030 , n18674 );
nand ( n41859 , n41857 , n41858 );
buf ( n41860 , n41859 );
buf ( n41861 , n41860 );
not ( n41862 , n275550 );
buf ( n41863 , n41862 );
buf ( n41864 , n41863 );
buf ( n41865 , n275554 );
buf ( n41866 , n275554 );
buf ( n41867 , n275554 );
buf ( n41868 , n275554 );
buf ( n41869 , n275554 );
not ( n41870 , n275929 );
buf ( n41871 , n41870 );
buf ( n41872 , n41871 );
buf ( n41873 , n275554 );
not ( n41874 , n275925 );
buf ( n41875 , n41874 );
buf ( n41876 , n41875 );
or ( n41877 , n36036 , n9144 );
and ( n41878 , n36047 , n9423 );
buf ( n41879 , n9137 );
buf ( n41880 , n41879 );
buf ( n41881 , n277957 );
xnor ( n41882 , n41880 , n41881 );
not ( n41883 , n41882 );
nand ( n41884 , n36106 , n36135 );
not ( n41885 , n36084 );
not ( n41886 , n36102 );
and ( n41887 , n41884 , n41885 , n41886 );
nor ( n41888 , n41887 , n36067 );
not ( n41889 , n41888 );
nand ( n41890 , n39992 , n36054 );
nor ( n41891 , n36102 , n36093 );
nor ( n41892 , n41890 , n41891 );
not ( n41893 , n41892 );
or ( n41894 , n41889 , n41893 );
not ( n41895 , n36146 );
not ( n41896 , n41890 );
not ( n41897 , n41896 );
or ( n41898 , n41895 , n41897 );
and ( n41899 , n36052 , n39992 );
nor ( n41900 , n41899 , n39994 );
nand ( n41901 , n41898 , n41900 );
not ( n41902 , n41901 );
nand ( n41903 , n41894 , n41902 );
buf ( n41904 , n11290 );
not ( n41905 , n41904 );
buf ( n41906 , n11302 );
nand ( n41907 , n41905 , n41906 );
buf ( n41908 , n11256 );
not ( n41909 , n41908 );
buf ( n41910 , n11202 );
nand ( n41911 , n41909 , n41910 );
and ( n41912 , n41907 , n41911 );
buf ( n41913 , n11372 );
not ( n41914 , n41913 );
buf ( n41915 , n11343 );
nand ( n41916 , n41914 , n41915 );
buf ( n41917 , n11432 );
buf ( n41918 , n11415 );
not ( n41919 , n41918 );
nand ( n41920 , n41917 , n41919 );
and ( n41921 , n41916 , n41920 );
and ( n41922 , n41912 , n41921 );
buf ( n41923 , n278066 );
not ( n41924 , n41923 );
not ( n41925 , n10630 );
buf ( n41926 , n41925 );
nand ( n41927 , n41924 , n41926 );
not ( n41928 , n41927 );
buf ( n41929 , n278032 );
not ( n41930 , n41929 );
buf ( n41931 , n278010 );
nor ( n41932 , n41930 , n41931 );
nor ( n41933 , n41928 , n41932 );
buf ( n41934 , n277948 );
not ( n41935 , n41934 );
buf ( n41936 , n277906 );
nand ( n41937 , n41935 , n41936 );
and ( n41938 , n41933 , n41937 );
and ( n41939 , n41903 , n41922 , n41938 );
not ( n41940 , n41938 );
not ( n41941 , n41920 );
not ( n41942 , n41915 );
nand ( n41943 , n41942 , n41913 );
or ( n41944 , n41941 , n41943 );
or ( n41945 , n41917 , n41919 );
nand ( n41946 , n41944 , n41945 );
not ( n41947 , n41946 );
not ( n41948 , n41912 );
or ( n41949 , n41947 , n41948 );
not ( n41950 , n41908 );
nor ( n41951 , n41950 , n41910 );
and ( n41952 , n41907 , n41951 );
not ( n41953 , n41904 );
nor ( n41954 , n41953 , n41906 );
nor ( n41955 , n41952 , n41954 );
nand ( n41956 , n41949 , n41955 );
not ( n41957 , n41956 );
or ( n41958 , n41940 , n41957 );
not ( n41959 , n41926 );
nand ( n41960 , n41959 , n41923 );
or ( n41961 , n41932 , n41960 );
not ( n41962 , n41929 );
nand ( n41963 , n41962 , n41931 );
nand ( n41964 , n41961 , n41963 );
and ( n41965 , n41964 , n41937 );
not ( n41966 , n41934 );
nor ( n41967 , n41966 , n41936 );
nor ( n41968 , n41965 , n41967 );
nand ( n41969 , n41958 , n41968 );
nor ( n41970 , n41939 , n41969 );
not ( n41971 , n41970 );
or ( n41972 , n41883 , n41971 );
or ( n41973 , n41970 , n41882 );
nand ( n41974 , n41972 , n41973 );
buf ( n41975 , n41974 );
not ( n41976 , n41975 );
not ( n41977 , n36155 );
or ( n41978 , n41976 , n41977 );
buf ( n41979 , n41879 );
buf ( n41980 , n277962 );
xnor ( n41981 , n41979 , n41980 );
not ( n41982 , n41981 );
nand ( n41983 , n36214 , n36241 );
not ( n41984 , n36194 );
and ( n41985 , n41983 , n41984 , n36210 );
nor ( n41986 , n41985 , n36178 );
not ( n41987 , n41986 );
and ( n41988 , n40012 , n36166 );
not ( n41989 , n41988 );
not ( n41990 , n36210 );
nor ( n41991 , n41990 , n36203 );
nor ( n41992 , n41989 , n41991 );
not ( n41993 , n41992 );
or ( n41994 , n41987 , n41993 );
not ( n41995 , n36252 );
not ( n41996 , n41988 );
or ( n41997 , n41995 , n41996 );
and ( n41998 , n36163 , n40012 );
nor ( n41999 , n41998 , n40014 );
nand ( n42000 , n41997 , n41999 );
not ( n42001 , n42000 );
nand ( n42002 , n41994 , n42001 );
buf ( n42003 , n11275 );
not ( n42004 , n42003 );
buf ( n42005 , n11302 );
nand ( n42006 , n42004 , n42005 );
buf ( n42007 , n11252 );
not ( n42008 , n42007 );
buf ( n42009 , n11202 );
nand ( n42010 , n42008 , n42009 );
and ( n42011 , n42006 , n42010 );
buf ( n42012 , n11378 );
not ( n42013 , n42012 );
buf ( n42014 , n11343 );
nand ( n42015 , n42013 , n42014 );
buf ( n42016 , n11432 );
buf ( n42017 , n11411 );
not ( n42018 , n42017 );
nand ( n42019 , n42016 , n42018 );
and ( n42020 , n42015 , n42019 );
and ( n42021 , n42011 , n42020 );
buf ( n42022 , n278059 );
not ( n42023 , n42022 );
buf ( n42024 , n41925 );
nand ( n42025 , n42023 , n42024 );
not ( n42026 , n42025 );
buf ( n42027 , n278032 );
not ( n42028 , n42027 );
buf ( n42029 , n278016 );
nor ( n42030 , n42028 , n42029 );
nor ( n42031 , n42026 , n42030 );
buf ( n42032 , n277934 );
not ( n42033 , n42032 );
buf ( n42034 , n277906 );
nand ( n42035 , n42033 , n42034 );
and ( n42036 , n42031 , n42035 );
and ( n42037 , n42002 , n42021 , n42036 );
not ( n42038 , n42036 );
not ( n42039 , n42019 );
not ( n42040 , n42012 );
nor ( n42041 , n42040 , n42014 );
not ( n42042 , n42041 );
or ( n42043 , n42039 , n42042 );
or ( n42044 , n42016 , n42018 );
nand ( n42045 , n42043 , n42044 );
not ( n42046 , n42045 );
not ( n42047 , n42011 );
or ( n42048 , n42046 , n42047 );
not ( n42049 , n42007 );
nor ( n42050 , n42049 , n42009 );
and ( n42051 , n42006 , n42050 );
not ( n42052 , n42003 );
nor ( n42053 , n42052 , n42005 );
nor ( n42054 , n42051 , n42053 );
nand ( n42055 , n42048 , n42054 );
not ( n42056 , n42055 );
or ( n42057 , n42038 , n42056 );
not ( n42058 , n42024 );
nand ( n42059 , n42058 , n42022 );
or ( n42060 , n42030 , n42059 );
not ( n42061 , n42027 );
nand ( n42062 , n42061 , n42029 );
nand ( n42063 , n42060 , n42062 );
and ( n42064 , n42063 , n42035 );
not ( n42065 , n42032 );
nor ( n42066 , n42065 , n42034 );
nor ( n42067 , n42064 , n42066 );
nand ( n42068 , n42057 , n42067 );
nor ( n42069 , n42037 , n42068 );
not ( n42070 , n42069 );
or ( n42071 , n41982 , n42070 );
or ( n42072 , n42069 , n41981 );
nand ( n42073 , n42071 , n42072 );
buf ( n42074 , n42073 );
nand ( n42075 , n41635 , n42074 );
nand ( n42076 , n41978 , n42075 );
nor ( n42077 , n41878 , n42076 );
nand ( n42078 , n41877 , n42077 );
nand ( n42079 , n42078 , n20645 );
buf ( n42080 , n41879 );
buf ( n42081 , n42080 );
buf ( n42082 , n277957 );
xnor ( n42083 , n42081 , n42082 );
not ( n42084 , n42083 );
and ( n42085 , n40034 , n36271 );
nand ( n42086 , n42085 , n36362 );
and ( n42087 , n36273 , n40034 );
nor ( n42088 , n42087 , n40037 );
nand ( n42089 , n42086 , n42088 );
not ( n42090 , n42089 );
or ( n42091 , n36295 , n36351 );
or ( n42092 , n36332 , n36351 , n36342 );
and ( n42093 , n36285 , n42092 );
nand ( n42094 , n42091 , n42093 , n42085 );
nand ( n42095 , n42090 , n42094 );
buf ( n42096 , n11343 );
not ( n42097 , n42096 );
buf ( n42098 , n11372 );
nand ( n42099 , n42097 , n42098 );
buf ( n42100 , n11432 );
not ( n42101 , n42100 );
buf ( n42102 , n11415 );
nand ( n42103 , n42101 , n42102 );
nand ( n42104 , n42099 , n42103 );
not ( n42105 , n42104 );
not ( n42106 , n42105 );
buf ( n42107 , n11290 );
not ( n42108 , n42107 );
buf ( n42109 , n11302 );
nor ( n42110 , n42108 , n42109 );
buf ( n42111 , n11256 );
not ( n42112 , n42111 );
buf ( n42113 , n11202 );
nor ( n42114 , n42112 , n42113 );
or ( n42115 , n42110 , n42114 );
nor ( n42116 , n42106 , n42115 );
buf ( n42117 , n41925 );
buf ( n42118 , n42117 );
not ( n42119 , n42118 );
buf ( n42120 , n278066 );
nand ( n42121 , n42119 , n42120 );
not ( n42122 , n42121 );
buf ( n42123 , n278010 );
not ( n42124 , n42123 );
buf ( n42125 , n39698 );
nor ( n42126 , n42124 , n42125 );
nor ( n42127 , n42122 , n42126 );
buf ( n42128 , n277906 );
not ( n42129 , n42128 );
buf ( n42130 , n277948 );
nand ( n42131 , n42129 , n42130 );
and ( n42132 , n42127 , n42131 );
and ( n42133 , n42095 , n42116 , n42132 );
not ( n42134 , n42132 );
nor ( n42135 , n42097 , n42098 );
and ( n42136 , n42135 , n42103 );
not ( n42137 , n42100 );
nor ( n42138 , n42137 , n42102 );
nor ( n42139 , n42136 , n42138 );
or ( n42140 , n42115 , n42139 );
not ( n42141 , n42111 );
nand ( n42142 , n42141 , n42113 );
or ( n42143 , n42110 , n42142 );
not ( n42144 , n42107 );
nand ( n42145 , n42144 , n42109 );
nand ( n42146 , n42140 , n42143 , n42145 );
not ( n42147 , n42146 );
or ( n42148 , n42134 , n42147 );
not ( n42149 , n42120 );
nand ( n42150 , n42149 , n42118 );
or ( n42151 , n42126 , n42150 );
not ( n42152 , n42123 );
nand ( n42153 , n42152 , n42125 );
nand ( n42154 , n42151 , n42153 );
and ( n42155 , n42154 , n42131 );
not ( n42156 , n42128 );
nor ( n42157 , n42156 , n42130 );
nor ( n42158 , n42155 , n42157 );
nand ( n42159 , n42148 , n42158 );
nor ( n42160 , n42133 , n42159 );
not ( n42161 , n42160 );
or ( n42162 , n42084 , n42161 );
or ( n42163 , n42160 , n42083 );
nand ( n42164 , n42162 , n42163 );
buf ( n42165 , n42164 );
nand ( n42166 , n36267 , n42165 );
buf ( n42167 , n42080 );
buf ( n42168 , n277962 );
xnor ( n42169 , n42167 , n42168 );
not ( n42170 , n42169 );
and ( n42171 , n40054 , n36375 );
nand ( n42172 , n42171 , n36465 );
and ( n42173 , n36377 , n40054 );
nor ( n42174 , n42173 , n40057 );
nand ( n42175 , n42172 , n42174 );
not ( n42176 , n42175 );
or ( n42177 , n36399 , n36454 );
or ( n42178 , n36435 , n36454 , n36445 );
and ( n42179 , n36389 , n42178 );
nand ( n42180 , n42177 , n42179 , n42171 );
nand ( n42181 , n42176 , n42180 );
buf ( n42182 , n11343 );
not ( n42183 , n42182 );
buf ( n42184 , n11378 );
nand ( n42185 , n42183 , n42184 );
buf ( n42186 , n11432 );
not ( n42187 , n42186 );
buf ( n42188 , n11411 );
nand ( n42189 , n42187 , n42188 );
nand ( n42190 , n42185 , n42189 );
not ( n42191 , n42190 );
not ( n42192 , n42191 );
buf ( n42193 , n11275 );
not ( n42194 , n42193 );
buf ( n42195 , n11302 );
nor ( n42196 , n42194 , n42195 );
buf ( n42197 , n11252 );
not ( n42198 , n42197 );
buf ( n42199 , n11202 );
nor ( n42200 , n42198 , n42199 );
or ( n42201 , n42196 , n42200 );
nor ( n42202 , n42192 , n42201 );
buf ( n42203 , n42117 );
not ( n42204 , n42203 );
buf ( n42205 , n278059 );
nand ( n42206 , n42204 , n42205 );
not ( n42207 , n42206 );
buf ( n42208 , n278016 );
not ( n42209 , n42208 );
buf ( n42210 , n39698 );
nor ( n42211 , n42209 , n42210 );
nor ( n42212 , n42207 , n42211 );
buf ( n42213 , n277906 );
not ( n42214 , n42213 );
buf ( n42215 , n277934 );
nand ( n42216 , n42214 , n42215 );
and ( n42217 , n42212 , n42216 );
and ( n42218 , n42181 , n42202 , n42217 );
not ( n42219 , n42217 );
nor ( n42220 , n42183 , n42184 );
and ( n42221 , n42220 , n42189 );
not ( n42222 , n42186 );
nor ( n42223 , n42222 , n42188 );
nor ( n42224 , n42221 , n42223 );
or ( n42225 , n42201 , n42224 );
not ( n42226 , n42197 );
nand ( n42227 , n42226 , n42199 );
or ( n42228 , n42196 , n42227 );
not ( n42229 , n42193 );
nand ( n42230 , n42229 , n42195 );
nand ( n42231 , n42225 , n42228 , n42230 );
not ( n42232 , n42231 );
or ( n42233 , n42219 , n42232 );
not ( n42234 , n42205 );
nand ( n42235 , n42234 , n42203 );
or ( n42236 , n42211 , n42235 );
not ( n42237 , n42208 );
nand ( n42238 , n42237 , n42210 );
nand ( n42239 , n42236 , n42238 );
and ( n42240 , n42239 , n42216 );
not ( n42241 , n42213 );
nor ( n42242 , n42241 , n42215 );
nor ( n42243 , n42240 , n42242 );
nand ( n42244 , n42233 , n42243 );
nor ( n42245 , n42218 , n42244 );
not ( n42246 , n42245 );
or ( n42247 , n42170 , n42246 );
or ( n42248 , n42245 , n42169 );
nand ( n42249 , n42247 , n42248 );
buf ( n42250 , n42249 );
nand ( n42251 , n36371 , n42250 );
and ( n42252 , n36474 , n9137 );
or ( n42253 , n20654 , n9422 );
nand ( n42254 , n42253 , n36930 );
nor ( n42255 , n42252 , n42254 );
nand ( n42256 , n42079 , n42166 , n42251 , n42255 );
buf ( n42257 , n42256 );
buf ( n42258 , n42257 );
not ( n42259 , n275550 );
buf ( n42260 , n42259 );
buf ( n42261 , n42260 );
not ( n42262 , n22335 );
not ( n42263 , n25276 );
or ( n42264 , n42262 , n42263 );
not ( n42265 , n21446 );
or ( n42266 , n42265 , n22335 );
nand ( n42267 , n42264 , n42266 );
buf ( n42268 , n42267 );
buf ( n42269 , n42268 );
buf ( n42270 , n275554 );
not ( n42271 , n23401 );
or ( n42272 , n42271 , n29046 );
nand ( n42273 , n29044 , n9728 );
nand ( n42274 , n42272 , n42273 );
buf ( n42275 , n42274 );
buf ( n42276 , n42275 );
not ( n42277 , n275929 );
buf ( n42278 , n42277 );
buf ( n42279 , n42278 );
buf ( n42280 , n275554 );
buf ( n42281 , n275554 );
not ( n42282 , n275929 );
buf ( n42283 , n42282 );
buf ( n42284 , n42283 );
buf ( n42285 , n275554 );
buf ( n42286 , n275554 );
not ( n42287 , n275925 );
buf ( n42288 , n42287 );
buf ( n42289 , n42288 );
or ( n42290 , n40426 , n21030 );
nand ( n42291 , n21030 , n18543 );
nand ( n42292 , n42290 , n42291 );
buf ( n42293 , n42292 );
buf ( n42294 , n42293 );
not ( n42295 , n26231 );
and ( n42296 , n22335 , n42295 );
not ( n42297 , n22335 );
and ( n42298 , n42297 , n21301 );
or ( n42299 , n42296 , n42298 );
buf ( n42300 , n42299 );
buf ( n42301 , n42300 );
and ( n42302 , n39578 , n39572 );
nor ( n42303 , n42302 , n39570 );
buf ( n42304 , n9416 );
not ( n42305 , n42304 );
buf ( n42306 , n9413 );
not ( n42307 , n42306 );
buf ( n42308 , n9423 );
not ( n42309 , n42308 );
and ( n42310 , n42307 , n42309 );
and ( n42311 , n42308 , n42306 );
nor ( n42312 , n42310 , n42311 );
not ( n42313 , n42312 );
or ( n42314 , n42305 , n42313 );
or ( n42315 , n42312 , n42304 );
nand ( n42316 , n42314 , n42315 );
not ( n42317 , n42316 );
xor ( n42318 , n39554 , n39558 );
and ( n42319 , n42318 , n39564 );
and ( n42320 , n39554 , n39558 );
or ( n42321 , n42319 , n42320 );
not ( n42322 , n42321 );
and ( n42323 , n42317 , n42322 );
and ( n42324 , n42316 , n42321 );
nor ( n42325 , n42323 , n42324 );
xnor ( n42326 , n42303 , n42325 );
buf ( n42327 , n42326 );
buf ( n42328 , n42327 );
buf ( n42329 , n275554 );
or ( n42330 , n33272 , n32073 );
and ( n42331 , n33236 , n20515 );
or ( n42332 , n19649 , n40323 );
nand ( n42333 , n33245 , n29492 );
nand ( n42334 , n20563 , n33250 );
nand ( n42335 , n275557 , n18614 );
nand ( n42336 , n42332 , n42333 , n42334 , n42335 );
nor ( n42337 , n42331 , n42336 );
nand ( n42338 , n33222 , n20353 );
nand ( n42339 , n42330 , n42337 , n42338 );
buf ( n42340 , n42339 );
buf ( n42341 , n42340 );
not ( n42342 , n275550 );
buf ( n42343 , n42342 );
buf ( n42344 , n42343 );
nand ( n42345 , n25064 , n42295 );
buf ( n42346 , n25297 );
buf ( n42347 , n25364 );
and ( n42348 , n42346 , n42347 );
buf ( n42349 , n42348 );
buf ( n42350 , n42349 );
not ( n42351 , n42350 );
buf ( n42352 , n25340 );
buf ( n42353 , n25285 );
and ( n42354 , n42352 , n42353 );
buf ( n42355 , n25131 );
buf ( n42356 , n25264 );
buf ( n42357 , n25285 );
and ( n42358 , n42355 , n42356 , n42357 );
buf ( n42359 , n42358 );
buf ( n42360 , n42359 );
buf ( n42361 , n25357 );
nor ( n42362 , n42354 , n42360 , n42361 );
buf ( n42363 , n42362 );
buf ( n42364 , n42363 );
not ( n42365 , n42364 );
or ( n42366 , n42351 , n42365 );
buf ( n42367 , n42363 );
buf ( n42368 , n42349 );
or ( n42369 , n42367 , n42368 );
nand ( n42370 , n42366 , n42369 );
buf ( n42371 , n42370 );
buf ( n42372 , n42371 );
not ( n42373 , n42372 );
nor ( n42374 , n42373 , n25389 );
nand ( n42375 , n25397 , n275576 );
buf ( n42376 , n25615 );
buf ( n42377 , n25693 );
nor ( n42378 , n42376 , n42377 );
buf ( n42379 , n42378 );
buf ( n42380 , n42379 );
not ( n42381 , n42380 );
buf ( n42382 , n25456 );
buf ( n42383 , n25586 );
buf ( n42384 , n25606 );
and ( n42385 , n42382 , n42383 , n42384 );
buf ( n42386 , n25666 );
buf ( n42387 , n25606 );
and ( n42388 , n42386 , n42387 );
buf ( n42389 , n25683 );
nor ( n42390 , n42388 , n42389 );
buf ( n42391 , n42390 );
buf ( n42392 , n42391 );
not ( n42393 , n42392 );
buf ( n42394 , n42393 );
buf ( n42395 , n42394 );
nor ( n42396 , n42385 , n42395 );
buf ( n42397 , n42396 );
buf ( n42398 , n42397 );
not ( n42399 , n42398 );
or ( n42400 , n42381 , n42399 );
buf ( n42401 , n42397 );
buf ( n42402 , n42379 );
or ( n42403 , n42401 , n42402 );
nand ( n42404 , n42400 , n42403 );
buf ( n42405 , n42404 );
buf ( n42406 , n42405 );
and ( n42407 , n25402 , n42406 );
nor ( n42408 , n42407 , n32086 );
buf ( n42409 , n25928 );
buf ( n42410 , n26004 );
nor ( n42411 , n42409 , n42410 );
buf ( n42412 , n42411 );
buf ( n42413 , n42412 );
not ( n42414 , n42413 );
buf ( n42415 , n25773 );
buf ( n42416 , n25902 );
buf ( n42417 , n25920 );
and ( n42418 , n42415 , n42416 , n42417 );
buf ( n42419 , n25977 );
buf ( n42420 , n25920 );
and ( n42421 , n42419 , n42420 );
buf ( n42422 , n25994 );
nor ( n42423 , n42421 , n42422 );
buf ( n42424 , n42423 );
buf ( n42425 , n42424 );
not ( n42426 , n42425 );
buf ( n42427 , n42426 );
buf ( n42428 , n42427 );
nor ( n42429 , n42418 , n42428 );
buf ( n42430 , n42429 );
buf ( n42431 , n42430 );
not ( n42432 , n42431 );
or ( n42433 , n42414 , n42432 );
buf ( n42434 , n42430 );
buf ( n42435 , n42412 );
or ( n42436 , n42434 , n42435 );
nand ( n42437 , n42433 , n42436 );
buf ( n42438 , n42437 );
buf ( n42439 , n42438 );
nand ( n42440 , n28761 , n42439 );
nand ( n42441 , n42375 , n42408 , n42440 );
nor ( n42442 , n42374 , n42441 );
buf ( n42443 , n26241 );
buf ( n42444 , n26305 );
and ( n42445 , n42443 , n42444 );
buf ( n42446 , n42445 );
buf ( n42447 , n42446 );
not ( n42448 , n42447 );
buf ( n42449 , n26281 );
buf ( n42450 , n26229 );
and ( n42451 , n42449 , n42450 );
buf ( n42452 , n26081 );
buf ( n42453 , n26212 );
buf ( n42454 , n26229 );
and ( n42455 , n42452 , n42453 , n42454 );
buf ( n42456 , n42455 );
buf ( n42457 , n42456 );
buf ( n42458 , n26298 );
nor ( n42459 , n42451 , n42457 , n42458 );
buf ( n42460 , n42459 );
buf ( n42461 , n42460 );
not ( n42462 , n42461 );
or ( n42463 , n42448 , n42462 );
buf ( n42464 , n42460 );
buf ( n42465 , n42446 );
or ( n42466 , n42464 , n42465 );
nand ( n42467 , n42463 , n42466 );
buf ( n42468 , n42467 );
buf ( n42469 , n42468 );
nand ( n42470 , n26027 , n42469 );
nand ( n42471 , n42345 , n42442 , n42470 );
buf ( n42472 , n42471 );
buf ( n42473 , n42472 );
buf ( n42474 , n275554 );
not ( n42475 , n275550 );
buf ( n42476 , n42475 );
buf ( n42477 , n42476 );
not ( n42478 , n15777 );
or ( n42479 , n42478 , n14830 );
or ( n42480 , n23806 , n14903 );
nand ( n42481 , n42479 , n42480 );
buf ( n42482 , n42481 );
buf ( n42483 , n42482 );
not ( n42484 , n275925 );
buf ( n42485 , n42484 );
buf ( n42486 , n42485 );
not ( n42487 , n29856 );
or ( n42488 , n42487 , n21774 );
nand ( n42489 , n21774 , n9787 );
nand ( n42490 , n42488 , n42489 );
buf ( n42491 , n42490 );
buf ( n42492 , n42491 );
not ( n42493 , n275550 );
buf ( n42494 , n42493 );
buf ( n42495 , n42494 );
not ( n42496 , n275925 );
buf ( n42497 , n42496 );
buf ( n42498 , n42497 );
buf ( n42499 , n275554 );
not ( n42500 , n275925 );
buf ( n42501 , n42500 );
buf ( n42502 , n42501 );
buf ( n42503 , n275554 );
buf ( n42504 , n275554 );
buf ( n42505 , n275554 );
buf ( n42506 , n275554 );
buf ( n42507 , n275554 );
buf ( n42508 , n275554 );
or ( n42509 , n36036 , n36485 );
and ( n42510 , n36045 , n275887 );
nand ( n42511 , n41943 , n41916 );
not ( n42512 , n42511 );
not ( n42513 , n41903 );
or ( n42514 , n42512 , n42513 );
or ( n42515 , n41903 , n42511 );
nand ( n42516 , n42514 , n42515 );
buf ( n42517 , n42516 );
not ( n42518 , n42517 );
not ( n42519 , n36155 );
or ( n42520 , n42518 , n42519 );
not ( n42521 , n42041 );
nand ( n42522 , n42521 , n42015 );
not ( n42523 , n42522 );
not ( n42524 , n42002 );
or ( n42525 , n42523 , n42524 );
or ( n42526 , n42002 , n42522 );
nand ( n42527 , n42525 , n42526 );
buf ( n42528 , n42527 );
nand ( n42529 , n41635 , n42528 );
nand ( n42530 , n42520 , n42529 );
nor ( n42531 , n42510 , n42530 );
nand ( n42532 , n42509 , n42531 );
nand ( n42533 , n42532 , n20645 );
not ( n42534 , n42135 );
nand ( n42535 , n42099 , n42534 );
not ( n42536 , n42535 );
not ( n42537 , n42095 );
or ( n42538 , n42536 , n42537 );
or ( n42539 , n42095 , n42535 );
nand ( n42540 , n42538 , n42539 );
buf ( n42541 , n42540 );
nand ( n42542 , n36267 , n42541 );
not ( n42543 , n42220 );
nand ( n42544 , n42185 , n42543 );
not ( n42545 , n42544 );
not ( n42546 , n42181 );
or ( n42547 , n42545 , n42546 );
or ( n42548 , n42181 , n42544 );
nand ( n42549 , n42547 , n42548 );
buf ( n42550 , n42549 );
nand ( n42551 , n36371 , n42550 );
and ( n42552 , n36474 , n11343 );
or ( n42553 , n20654 , n275886 );
nand ( n42554 , n42553 , n28461 );
nor ( n42555 , n42552 , n42554 );
nand ( n42556 , n42533 , n42542 , n42551 , n42555 );
buf ( n42557 , n42556 );
buf ( n42558 , n42557 );
not ( n42559 , n275550 );
buf ( n42560 , n42559 );
buf ( n42561 , n42560 );
and ( n42562 , n29126 , n32751 );
not ( n42563 , n12264 );
not ( n42564 , n29171 );
or ( n42565 , n42563 , n42564 );
and ( n42566 , n28458 , n10740 );
nand ( n42567 , n20649 , n9291 );
not ( n42568 , n42567 );
nor ( n42569 , n42566 , n42568 );
nand ( n42570 , n42565 , n42569 );
nor ( n42571 , n42562 , n42570 );
nand ( n42572 , n29138 , n29163 );
nand ( n42573 , n29153 , n28408 );
not ( n42574 , n28450 );
nand ( n42575 , n42574 , n37672 );
nand ( n42576 , n42571 , n42572 , n42573 , n42575 );
buf ( n42577 , n42576 );
buf ( n42578 , n42577 );
buf ( n42579 , n275554 );
buf ( n42580 , n275554 );
buf ( n42581 , n275554 );
buf ( n42582 , n275554 );
not ( n42583 , n275929 );
buf ( n42584 , n42583 );
buf ( n42585 , n42584 );
or ( n42586 , n39315 , n19634 );
and ( n42587 , n29471 , n38735 );
not ( n42588 , n39323 );
not ( n42589 , n30612 );
or ( n42590 , n42588 , n42589 );
nand ( n42591 , n38750 , n29492 );
nand ( n42592 , n20563 , n38739 );
nand ( n42593 , n30179 , n18668 );
and ( n42594 , n42591 , n42592 , n42593 );
nand ( n42595 , n42590 , n42594 );
nor ( n42596 , n42587 , n42595 );
nand ( n42597 , n38721 , n20353 );
and ( n42598 , n42596 , n42597 );
nand ( n42599 , n42586 , n42598 );
buf ( n42600 , n42599 );
buf ( n42601 , n42600 );
not ( n42602 , n275925 );
buf ( n42603 , n42602 );
buf ( n42604 , n42603 );
not ( n42605 , n27810 );
or ( n42606 , n42605 , n21774 );
nand ( n42607 , n21774 , n9752 );
nand ( n42608 , n42606 , n42607 );
buf ( n42609 , n42608 );
buf ( n42610 , n42609 );
buf ( n42611 , n275554 );
or ( n42612 , n39197 , n21030 );
nand ( n42613 , n21030 , n18912 );
nand ( n42614 , n42612 , n42613 );
buf ( n42615 , n42614 );
buf ( n42616 , n42615 );
not ( n42617 , n22335 );
not ( n42618 , n25267 );
or ( n42619 , n42617 , n42618 );
not ( n42620 , n21351 );
or ( n42621 , n42620 , n22335 );
nand ( n42622 , n42619 , n42621 );
buf ( n42623 , n42622 );
buf ( n42624 , n42623 );
and ( n42625 , n23706 , n277833 );
not ( n42626 , n23706 );
not ( n42627 , n29599 );
buf ( n42628 , n39344 );
buf ( n42629 , n30878 );
nand ( n42630 , n42628 , n42629 );
buf ( n42631 , n42630 );
buf ( n42632 , n42631 );
not ( n42633 , n42632 );
buf ( n42634 , n30820 );
not ( n42635 , n42634 );
buf ( n42636 , n27479 );
not ( n42637 , n42636 );
or ( n42638 , n42635 , n42637 );
buf ( n42639 , n39357 );
not ( n42640 , n42639 );
buf ( n42641 , n42640 );
buf ( n42642 , n42641 );
nand ( n42643 , n42638 , n42642 );
buf ( n42644 , n42643 );
buf ( n42645 , n42644 );
not ( n42646 , n42645 );
or ( n42647 , n42633 , n42646 );
buf ( n42648 , n42644 );
buf ( n42649 , n42631 );
or ( n42650 , n42648 , n42649 );
nand ( n42651 , n42647 , n42650 );
buf ( n42652 , n42651 );
buf ( n42653 , n42652 );
not ( n42654 , n42653 );
or ( n42655 , n42627 , n42654 );
nand ( n42656 , n30921 , n30949 );
not ( n42657 , n42656 );
not ( n42658 , n30931 );
not ( n42659 , n29728 );
or ( n42660 , n42658 , n42659 );
not ( n42661 , n39389 );
nand ( n42662 , n42660 , n42661 );
not ( n42663 , n42662 );
or ( n42664 , n42657 , n42663 );
or ( n42665 , n42662 , n42656 );
nand ( n42666 , n42664 , n42665 );
buf ( n42667 , n42666 );
and ( n42668 , n42667 , n30962 );
not ( n42669 , n23673 );
not ( n42670 , n30977 );
not ( n42671 , n39403 );
or ( n42672 , n42670 , n42671 );
buf ( n42673 , n39403 );
or ( n42674 , n42673 , n30977 );
nand ( n42675 , n42672 , n42674 );
buf ( n42676 , n42675 );
not ( n42677 , n42676 );
or ( n42678 , n42669 , n42677 );
and ( n42679 , n27520 , n11826 );
and ( n42680 , n22013 , n12248 );
nor ( n42681 , n42679 , n42680 );
nand ( n42682 , n42678 , n42681 );
nor ( n42683 , n42668 , n42682 );
nand ( n42684 , n42655 , n42683 );
and ( n42685 , n42626 , n42684 );
or ( n42686 , n42625 , n42685 );
buf ( n42687 , n42686 );
buf ( n42688 , n42687 );
buf ( n42689 , n275554 );
buf ( n42690 , n275554 );
or ( n42691 , n33994 , n19216 );
nand ( n42692 , n34008 , n35150 );
nor ( n42693 , n32248 , n34030 );
not ( n42694 , n34024 );
not ( n42695 , n29075 );
or ( n42696 , n42694 , n42695 );
nand ( n42697 , n19318 , n30615 );
nand ( n42698 , n42696 , n42697 );
nor ( n42699 , n42693 , n42698 );
nand ( n42700 , n34018 , n19360 );
nand ( n42701 , n19387 , n18866 );
and ( n42702 , n42692 , n42699 , n42700 , n42701 );
nand ( n42703 , n42691 , n42702 );
buf ( n42704 , n42703 );
buf ( n42705 , n42704 );
nand ( n42706 , n25063 , n17586 );
xor ( n42707 , n25182 , n25185 );
buf ( n42708 , n42707 );
buf ( n42709 , n42708 );
and ( n42710 , n34544 , n42709 );
not ( n42711 , n275750 );
not ( n42712 , n25396 );
or ( n42713 , n42711 , n42712 );
xor ( n42714 , n25503 , n25504 );
buf ( n42715 , n42714 );
buf ( n42716 , n42715 );
and ( n42717 , n25402 , n42716 );
xor ( n42718 , n25819 , n25820 );
buf ( n42719 , n42718 );
buf ( n42720 , n42719 );
not ( n42721 , n42720 );
not ( n42722 , n28761 );
or ( n42723 , n42721 , n42722 );
nand ( n42724 , n275557 , n18283 );
nand ( n42725 , n42723 , n42724 );
nor ( n42726 , n42717 , n42725 );
nand ( n42727 , n42713 , n42726 );
nor ( n42728 , n42710 , n42727 );
xor ( n42729 , n26128 , n26130 );
buf ( n42730 , n42729 );
buf ( n42731 , n42730 );
nand ( n42732 , n26027 , n42731 );
nand ( n42733 , n42706 , n42728 , n42732 );
buf ( n42734 , n42733 );
buf ( n42735 , n42734 );
buf ( n42736 , n275554 );
buf ( n42737 , n275554 );
buf ( n42738 , n275554 );
not ( n42739 , n275925 );
buf ( n42740 , n42739 );
buf ( n42741 , n42740 );
or ( n42742 , n41082 , n28146 );
nand ( n42743 , n24452 , n18754 );
nand ( n42744 , n42742 , n42743 );
buf ( n42745 , n42744 );
buf ( n42746 , n42745 );
and ( n42747 , n31719 , n277707 );
not ( n42748 , n31719 );
not ( n42749 , n29599 );
buf ( n42750 , n31891 );
buf ( n42751 , n31907 );
nand ( n42752 , n42750 , n42751 );
buf ( n42753 , n42752 );
buf ( n42754 , n42753 );
not ( n42755 , n42754 );
buf ( n42756 , n30798 );
not ( n42757 , n42756 );
buf ( n42758 , n30840 );
nor ( n42759 , n42757 , n42758 );
buf ( n42760 , n42759 );
buf ( n42761 , n42760 );
not ( n42762 , n42761 );
buf ( n42763 , n30823 );
nor ( n42764 , n42762 , n42763 );
buf ( n42765 , n42764 );
buf ( n42766 , n42765 );
not ( n42767 , n42766 );
buf ( n42768 , n27479 );
not ( n42769 , n42768 );
or ( n42770 , n42767 , n42769 );
buf ( n42771 , n42760 );
buf ( n42772 , n39357 );
and ( n42773 , n42771 , n42772 );
buf ( n42774 , n30798 );
not ( n42775 , n42774 );
buf ( n42776 , n30891 );
not ( n42777 , n42776 );
or ( n42778 , n42775 , n42777 );
buf ( n42779 , n30806 );
nand ( n42780 , n42778 , n42779 );
buf ( n42781 , n42780 );
buf ( n42782 , n42781 );
nor ( n42783 , n42773 , n42782 );
buf ( n42784 , n42783 );
buf ( n42785 , n42784 );
nand ( n42786 , n42770 , n42785 );
buf ( n42787 , n42786 );
buf ( n42788 , n42787 );
not ( n42789 , n42788 );
or ( n42790 , n42755 , n42789 );
buf ( n42791 , n42787 );
buf ( n42792 , n42753 );
or ( n42793 , n42791 , n42792 );
nand ( n42794 , n42790 , n42793 );
buf ( n42795 , n42794 );
buf ( n42796 , n42795 );
not ( n42797 , n42796 );
or ( n42798 , n42749 , n42797 );
nand ( n42799 , n31975 , n32006 );
not ( n42800 , n42799 );
nor ( n42801 , n30926 , n30913 );
not ( n42802 , n42801 );
nor ( n42803 , n42802 , n30932 );
not ( n42804 , n42803 );
not ( n42805 , n29728 );
or ( n42806 , n42804 , n42805 );
not ( n42807 , n42801 );
not ( n42808 , n39389 );
or ( n42809 , n42807 , n42808 );
and ( n42810 , n30954 , n30912 );
nor ( n42811 , n42810 , n30915 );
nand ( n42812 , n42809 , n42811 );
not ( n42813 , n42812 );
nand ( n42814 , n42806 , n42813 );
not ( n42815 , n42814 );
or ( n42816 , n42800 , n42815 );
or ( n42817 , n42814 , n42799 );
nand ( n42818 , n42816 , n42817 );
buf ( n42819 , n42818 );
and ( n42820 , n42819 , n23655 );
not ( n42821 , n23673 );
not ( n42822 , n32035 );
not ( n42823 , n42822 );
nor ( n42824 , n30982 , n30966 );
not ( n42825 , n42824 );
or ( n42826 , n42823 , n42825 );
or ( n42827 , n42824 , n42822 );
nand ( n42828 , n42826 , n42827 );
buf ( n42829 , n42828 );
not ( n42830 , n42829 );
or ( n42831 , n42821 , n42830 );
and ( n42832 , n27520 , n12371 );
and ( n42833 , n22013 , n12304 );
nor ( n42834 , n42832 , n42833 );
nand ( n42835 , n42831 , n42834 );
nor ( n42836 , n42820 , n42835 );
nand ( n42837 , n42798 , n42836 );
and ( n42838 , n42748 , n42837 );
or ( n42839 , n42747 , n42838 );
buf ( n42840 , n42839 );
buf ( n42841 , n42840 );
not ( n42842 , n275550 );
buf ( n42843 , n42842 );
buf ( n42844 , n42843 );
not ( n42845 , n275925 );
buf ( n42846 , n42845 );
buf ( n42847 , n42846 );
buf ( n42848 , n275554 );
not ( n42849 , n275550 );
buf ( n42850 , n42849 );
buf ( n42851 , n42850 );
buf ( n42852 , n275554 );
not ( n42853 , n21990 );
not ( n42854 , n42853 );
not ( n42855 , n28304 );
and ( n42856 , n42854 , n42855 );
and ( n42857 , n22141 , n28328 );
nor ( n42858 , n42856 , n42857 );
and ( n42859 , n22049 , n37665 );
nor ( n42860 , n28241 , n12128 );
nor ( n42861 , n42859 , n42860 );
and ( n42862 , n31451 , n12337 );
not ( n42863 , n10799 );
or ( n42864 , n28233 , n42863 );
not ( n42865 , n40089 );
or ( n42866 , n28356 , n42865 );
nand ( n42867 , n42864 , n42866 );
nor ( n42868 , n42862 , n42867 );
nand ( n42869 , n42858 , n42861 , n42868 );
buf ( n42870 , n42869 );
buf ( n42871 , n42870 );
and ( n42872 , n28196 , n31767 );
and ( n42873 , n28186 , n31780 );
nor ( n42874 , n42872 , n42873 );
not ( n42875 , n12282 );
and ( n42876 , n31451 , n42875 );
or ( n42877 , n28233 , n11072 );
nand ( n42878 , n28357 , n31784 );
nand ( n42879 , n42877 , n42878 );
nor ( n42880 , n42876 , n42879 );
nand ( n42881 , n28219 , n31744 );
nand ( n42882 , n31459 , n12192 );
nand ( n42883 , n42874 , n42880 , n42881 , n42882 );
buf ( n42884 , n42883 );
buf ( n42885 , n42884 );
not ( n42886 , n275550 );
buf ( n42887 , n42886 );
buf ( n42888 , n42887 );
not ( n42889 , n275925 );
buf ( n42890 , n42889 );
buf ( n42891 , n42890 );
not ( n42892 , n275925 );
buf ( n42893 , n42892 );
buf ( n42894 , n42893 );
not ( n42895 , n275929 );
buf ( n42896 , n42895 );
buf ( n42897 , n42896 );
or ( n42898 , n19143 , n19167 );
nand ( n42899 , n42898 , n19631 );
buf ( n42900 , n42899 );
buf ( n42901 , n42900 );
not ( n42902 , n29795 );
or ( n42903 , n42902 , n21774 );
nand ( n42904 , n21774 , n9744 );
nand ( n42905 , n42903 , n42904 );
buf ( n42906 , n42905 );
buf ( n42907 , n42906 );
not ( n42908 , n275550 );
buf ( n42909 , n42908 );
buf ( n42910 , n42909 );
buf ( n42911 , n275554 );
not ( n42912 , n275929 );
buf ( n42913 , n42912 );
buf ( n42914 , n42913 );
buf ( n42915 , n275554 );
not ( n42916 , n16201 );
or ( n42917 , n42916 , n14830 );
nand ( n42918 , n23069 , n23807 );
nand ( n42919 , n42917 , n42918 );
buf ( n42920 , n42919 );
buf ( n42921 , n42920 );
buf ( n42922 , n275554 );
buf ( n42923 , n29057 );
not ( n42924 , n42923 );
not ( n42925 , n14759 );
nand ( n42926 , n42925 , n24813 );
buf ( n42927 , n42926 );
not ( n42928 , n42927 );
not ( n42929 , n42928 );
not ( n42930 , n42929 );
or ( n42931 , n42924 , n42930 );
not ( n42932 , n42928 );
buf ( n42933 , n16332 );
buf ( n42934 , n16766 );
buf ( n42935 , n16440 );
buf ( n42936 , n16763 );
buf ( n42937 , n42936 );
and ( n42938 , n42933 , n42934 , n42935 , n42937 );
not ( n42939 , n42938 );
not ( n42940 , n16815 );
buf ( n42941 , n42940 );
buf ( n42942 , n16485 );
nand ( n42943 , n42941 , n42942 );
nor ( n42944 , n42939 , n42943 );
buf ( n42945 , n42944 );
buf ( n42946 , n16212 );
buf ( n42947 , n16151 );
and ( n42948 , n42946 , n42947 );
not ( n42949 , n42948 );
buf ( n42950 , n16296 );
buf ( n42951 , n17202 );
nand ( n42952 , n42950 , n42951 );
nor ( n42953 , n42949 , n42952 );
buf ( n42954 , n16650 );
buf ( n42955 , n16614 );
and ( n42956 , n42954 , n42955 );
nand ( n42957 , n42945 , n42953 , n42956 );
buf ( n42958 , n16509 );
not ( n42959 , n42958 );
and ( n42960 , n42957 , n42959 );
not ( n42961 , n42957 );
and ( n42962 , n42961 , n42958 );
nor ( n42963 , n42960 , n42962 );
buf ( n42964 , n42963 );
not ( n42965 , n42964 );
or ( n42966 , n42932 , n42965 );
nand ( n42967 , n42931 , n42966 );
buf ( n42968 , n42967 );
not ( n42969 , n34927 );
buf ( n42970 , n42969 );
not ( n42971 , n42970 );
nor ( n42972 , n42968 , n42971 );
buf ( n42973 , n31140 );
not ( n42974 , n42973 );
buf ( n42975 , n42927 );
not ( n42976 , n42975 );
or ( n42977 , n42974 , n42976 );
buf ( n42978 , n15839 );
buf ( n42979 , n42978 );
not ( n42980 , n42979 );
and ( n42981 , n42944 , n42953 );
not ( n42982 , n42956 );
nor ( n42983 , n42982 , n42959 );
nand ( n42984 , n42981 , n42983 );
not ( n42985 , n42984 );
or ( n42986 , n42980 , n42985 );
or ( n42987 , n42984 , n42979 );
nand ( n42988 , n42986 , n42987 );
buf ( n42989 , n42988 );
not ( n42990 , n42989 );
or ( n42991 , n42932 , n42990 );
nand ( n42992 , n42977 , n42991 );
buf ( n42993 , n42992 );
buf ( n42994 , n17450 );
buf ( n42995 , n42994 );
buf ( n42996 , n42995 );
buf ( n42997 , n42996 );
not ( n42998 , n42997 );
nor ( n42999 , n42993 , n42998 );
nor ( n43000 , n42972 , n42999 );
buf ( n43001 , n34092 );
not ( n43002 , n43001 );
not ( n43003 , n42975 );
or ( n43004 , n43002 , n43003 );
buf ( n43005 , n42927 );
nand ( n43006 , n42945 , n42953 , n42954 );
buf ( n43007 , n42955 );
not ( n43008 , n43007 );
and ( n43009 , n43006 , n43008 );
not ( n43010 , n43006 );
and ( n43011 , n43010 , n43007 );
nor ( n43012 , n43009 , n43011 );
buf ( n43013 , n43012 );
not ( n43014 , n43013 );
or ( n43015 , n43005 , n43014 );
nand ( n43016 , n43004 , n43015 );
buf ( n43017 , n43016 );
buf ( n43018 , n26497 );
not ( n43019 , n43018 );
nor ( n43020 , n43017 , n43019 );
not ( n43021 , n26423 );
not ( n43022 , n43021 );
not ( n43023 , n43022 );
not ( n43024 , n42927 );
not ( n43025 , n43024 );
not ( n43026 , n43025 );
or ( n43027 , n43023 , n43026 );
buf ( n43028 , n42927 );
xor ( n43029 , n42981 , n42954 );
buf ( n43030 , n43029 );
not ( n43031 , n43030 );
or ( n43032 , n43028 , n43031 );
nand ( n43033 , n43027 , n43032 );
buf ( n43034 , n43033 );
buf ( n43035 , n27728 );
not ( n43036 , n43035 );
nor ( n43037 , n43034 , n43036 );
nor ( n43038 , n43020 , n43037 );
nand ( n43039 , n43000 , n43038 );
not ( n43040 , n27685 );
not ( n43041 , n43040 );
not ( n43042 , n43041 );
not ( n43043 , n42975 );
or ( n43044 , n43042 , n43043 );
not ( n43045 , n42946 );
nor ( n43046 , n42952 , n43045 );
nand ( n43047 , n42945 , n43046 );
not ( n43048 , n42947 );
and ( n43049 , n43047 , n43048 );
not ( n43050 , n43047 );
and ( n43051 , n43050 , n42947 );
nor ( n43052 , n43049 , n43051 );
buf ( n43053 , n43052 );
not ( n43054 , n43053 );
or ( n43055 , n43005 , n43054 );
nand ( n43056 , n43044 , n43055 );
buf ( n43057 , n43056 );
buf ( n43058 , n27161 );
not ( n43059 , n43058 );
nor ( n43060 , n43057 , n43059 );
not ( n43061 , n42952 );
nand ( n43062 , n43061 , n42945 );
and ( n43063 , n43062 , n43045 );
not ( n43064 , n43062 );
and ( n43065 , n43064 , n42946 );
nor ( n43066 , n43063 , n43065 );
buf ( n43067 , n43066 );
not ( n43068 , n43067 );
or ( n43069 , n43028 , n43068 );
not ( n43070 , n27098 );
not ( n43071 , n43070 );
nand ( n43072 , n43025 , n43071 );
nand ( n43073 , n43069 , n43072 );
buf ( n43074 , n43073 );
buf ( n43075 , n20943 );
not ( n43076 , n43075 );
nor ( n43077 , n43074 , n43076 );
nor ( n43078 , n43060 , n43077 );
buf ( n43079 , n32353 );
not ( n43080 , n43079 );
not ( n43081 , n43005 );
or ( n43082 , n43080 , n43081 );
xor ( n43083 , n42950 , n42945 );
buf ( n43084 , n43083 );
not ( n43085 , n43084 );
or ( n43086 , n43028 , n43085 );
nand ( n43087 , n43082 , n43086 );
buf ( n43088 , n43087 );
buf ( n43089 , n32192 );
not ( n43090 , n43089 );
nand ( n43091 , n43088 , n43090 );
buf ( n43092 , n32405 );
not ( n43093 , n43092 );
not ( n43094 , n20820 );
not ( n43095 , n43094 );
not ( n43096 , n43095 );
not ( n43097 , n43024 );
not ( n43098 , n43097 );
or ( n43099 , n43096 , n43098 );
nand ( n43100 , n42945 , n42950 );
not ( n43101 , n42951 );
and ( n43102 , n43100 , n43101 );
not ( n43103 , n43100 );
and ( n43104 , n43103 , n42951 );
nor ( n43105 , n43102 , n43104 );
buf ( n43106 , n43105 );
not ( n43107 , n43106 );
or ( n43108 , n42932 , n43107 );
nand ( n43109 , n43099 , n43108 );
buf ( n43110 , n43109 );
nand ( n43111 , n43093 , n43110 );
and ( n43112 , n43091 , n43111 );
not ( n43113 , n43092 );
nor ( n43114 , n43113 , n43110 );
nor ( n43115 , n43112 , n43114 );
and ( n43116 , n43078 , n43115 );
nand ( n43117 , n43074 , n43076 );
or ( n43118 , n43060 , n43117 );
nand ( n43119 , n43057 , n43059 );
nand ( n43120 , n43118 , n43119 );
nor ( n43121 , n43116 , n43120 );
or ( n43122 , n43039 , n43121 );
nand ( n43123 , n43034 , n43036 );
or ( n43124 , n43020 , n43123 );
nand ( n43125 , n43017 , n43019 );
nand ( n43126 , n43124 , n43125 );
and ( n43127 , n43000 , n43126 );
nand ( n43128 , n42968 , n42971 );
or ( n43129 , n42999 , n43128 );
nand ( n43130 , n42993 , n42998 );
nand ( n43131 , n43129 , n43130 );
nor ( n43132 , n43127 , n43131 );
nand ( n43133 , n43122 , n43132 );
not ( n43134 , n43133 );
buf ( n43135 , n28249 );
buf ( n43136 , n43135 );
not ( n43137 , n43136 );
not ( n43138 , n42932 );
or ( n43139 , n43137 , n43138 );
not ( n43140 , n42975 );
not ( n43141 , n43140 );
buf ( n43142 , n42934 );
not ( n43143 , n43142 );
not ( n43144 , n42937 );
and ( n43145 , n43143 , n43144 );
nand ( n43146 , n43142 , n42937 );
not ( n43147 , n43146 );
nor ( n43148 , n43145 , n43147 );
buf ( n43149 , n43148 );
not ( n43150 , n43149 );
or ( n43151 , n43141 , n43150 );
nand ( n43152 , n43139 , n43151 );
buf ( n43153 , n43152 );
not ( n43154 , n34722 );
buf ( n43155 , n43154 );
not ( n43156 , n43155 );
nor ( n43157 , n43153 , n43156 );
buf ( n43158 , n20679 );
not ( n43159 , n43158 );
buf ( n43160 , n16705 );
buf ( n43161 , n43160 );
buf ( n43162 , n43161 );
buf ( n43163 , n43162 );
nor ( n43164 , n43159 , n43163 );
buf ( n43165 , n14542 );
not ( n43166 , n43165 );
buf ( n43167 , n21685 );
and ( n43168 , n43166 , n43167 );
or ( n43169 , n43164 , n43168 );
or ( n43170 , n43166 , n43167 );
nand ( n43171 , n43169 , n43170 );
buf ( n43172 , n14564 );
buf ( n43173 , n43172 );
buf ( n43174 , n43173 );
not ( n43175 , n43174 );
buf ( n43176 , n36638 );
nand ( n43177 , n43175 , n43176 );
and ( n43178 , n43171 , n43177 );
not ( n43179 , n43176 );
and ( n43180 , n43174 , n43179 );
nor ( n43181 , n43178 , n43180 );
or ( n43182 , n43157 , n43181 );
nand ( n43183 , n43153 , n43156 );
nand ( n43184 , n43182 , n43183 );
not ( n43185 , n42927 );
not ( n43186 , n43185 );
buf ( n43187 , n42941 );
nand ( n43188 , n43147 , n43187 );
xnor ( n43189 , n43188 , n42942 );
buf ( n43190 , n43189 );
not ( n43191 , n43190 );
or ( n43192 , n43186 , n43191 );
not ( n43193 , n43024 );
buf ( n43194 , n24672 );
buf ( n43195 , n43194 );
nand ( n43196 , n43193 , n43195 );
nand ( n43197 , n43192 , n43196 );
buf ( n43198 , n43197 );
buf ( n43199 , n34668 );
not ( n43200 , n43199 );
nor ( n43201 , n43198 , n43200 );
buf ( n43202 , n34623 );
buf ( n43203 , n43202 );
not ( n43204 , n43203 );
not ( n43205 , n42975 );
or ( n43206 , n43204 , n43205 );
not ( n43207 , n43187 );
not ( n43208 , n43146 );
or ( n43209 , n43207 , n43208 );
or ( n43210 , n43146 , n43187 );
nand ( n43211 , n43209 , n43210 );
buf ( n43212 , n43211 );
not ( n43213 , n43212 );
or ( n43214 , n43028 , n43213 );
nand ( n43215 , n43206 , n43214 );
buf ( n43216 , n43215 );
buf ( n43217 , n32958 );
not ( n43218 , n43217 );
nor ( n43219 , n43216 , n43218 );
nor ( n43220 , n43201 , n43219 );
buf ( n43221 , n32131 );
buf ( n43222 , n43221 );
not ( n43223 , n43222 );
not ( n43224 , n42975 );
or ( n43225 , n43223 , n43224 );
not ( n43226 , n42943 );
nand ( n43227 , n43226 , n43147 , n42935 );
xnor ( n43228 , n43227 , n42933 );
buf ( n43229 , n43228 );
not ( n43230 , n43229 );
or ( n43231 , n43028 , n43230 );
nand ( n43232 , n43225 , n43231 );
buf ( n43233 , n43232 );
buf ( n43234 , n37915 );
not ( n43235 , n43234 );
nor ( n43236 , n43233 , n43235 );
buf ( n43237 , n37860 );
buf ( n43238 , n43237 );
not ( n43239 , n43238 );
not ( n43240 , n43097 );
or ( n43241 , n43239 , n43240 );
nor ( n43242 , n43146 , n42943 );
xor ( n43243 , n43242 , n42935 );
buf ( n43244 , n43243 );
not ( n43245 , n43244 );
or ( n43246 , n43186 , n43245 );
nand ( n43247 , n43241 , n43246 );
buf ( n43248 , n43247 );
buf ( n43249 , n24724 );
not ( n43250 , n43249 );
nor ( n43251 , n43248 , n43250 );
nor ( n43252 , n43236 , n43251 );
nand ( n43253 , n43184 , n43220 , n43252 );
not ( n43254 , n43253 );
nand ( n43255 , n43216 , n43218 );
nand ( n43256 , n43198 , n43200 );
and ( n43257 , n43255 , n43256 );
nor ( n43258 , n43257 , n43201 );
and ( n43259 , n43252 , n43258 );
nand ( n43260 , n43248 , n43250 );
or ( n43261 , n43236 , n43260 );
nand ( n43262 , n43233 , n43235 );
nand ( n43263 , n43261 , n43262 );
nor ( n43264 , n43259 , n43263 );
not ( n43265 , n43264 );
or ( n43266 , n43254 , n43265 );
nor ( n43267 , n43088 , n43090 );
nor ( n43268 , n43114 , n43267 );
nand ( n43269 , n43078 , n43268 );
nor ( n43270 , n43039 , n43269 );
nand ( n43271 , n43266 , n43270 );
nand ( n43272 , n43134 , n43271 );
buf ( n43273 , n24937 );
not ( n43274 , n43273 );
not ( n43275 , n24767 );
not ( n43276 , n43275 );
not ( n43277 , n43276 );
not ( n43278 , n43025 );
or ( n43279 , n43277 , n43278 );
nor ( n43280 , n42943 , n42952 );
and ( n43281 , n42978 , n42958 );
nand ( n43282 , n43280 , n42948 , n43281 );
nand ( n43283 , n42956 , n42938 );
nor ( n43284 , n43282 , n43283 );
buf ( n43285 , n43284 );
not ( n43286 , n17070 );
buf ( n43287 , n43286 );
buf ( n43288 , n15733 );
buf ( n43289 , n17011 );
buf ( n43290 , n16016 );
nand ( n43291 , n43287 , n43288 , n43289 , n43290 );
not ( n43292 , n43291 );
buf ( n43293 , n15621 );
buf ( n43294 , n43293 );
buf ( n43295 , n15800 );
buf ( n43296 , n43295 );
nand ( n43297 , n43294 , n43296 );
buf ( n43298 , n15966 );
buf ( n43299 , n16027 );
nand ( n43300 , n43298 , n43299 );
nor ( n43301 , n43297 , n43300 );
nand ( n43302 , n43292 , n43301 );
not ( n43303 , n43302 );
buf ( n43304 , n16975 );
buf ( n43305 , n15512 );
and ( n43306 , n43304 , n43305 );
buf ( n43307 , n30271 );
not ( n43308 , n43307 );
buf ( n43309 , n24541 );
buf ( n43310 , n43309 );
not ( n43311 , n43310 );
nor ( n43312 , n43308 , n43311 );
and ( n43313 , n43306 , n43312 );
nand ( n43314 , n43285 , n43303 , n43313 );
buf ( n43315 , n30322 );
not ( n43316 , n43315 );
xor ( n43317 , n43314 , n43316 );
buf ( n43318 , n43317 );
not ( n43319 , n43318 );
or ( n43320 , n43005 , n43319 );
nand ( n43321 , n43279 , n43320 );
buf ( n43322 , n43321 );
not ( n43323 , n43322 );
not ( n43324 , n43323 );
or ( n43325 , n43274 , n43324 );
nand ( n43326 , n43313 , n43315 );
nor ( n43327 , n43326 , n43302 );
nand ( n43328 , n43327 , n43285 );
buf ( n43329 , n34431 );
not ( n43330 , n43329 );
and ( n43331 , n43328 , n43330 );
not ( n43332 , n43328 );
and ( n43333 , n43332 , n43329 );
nor ( n43334 , n43331 , n43333 );
buf ( n43335 , n43334 );
not ( n43336 , n43335 );
or ( n43337 , n42929 , n43336 );
not ( n43338 , n24790 );
not ( n43339 , n43338 );
nand ( n43340 , n43097 , n43339 );
nand ( n43341 , n43337 , n43340 );
buf ( n43342 , n43341 );
not ( n43343 , n43342 );
buf ( n43344 , n24939 );
nand ( n43345 , n43343 , n43344 );
nand ( n43346 , n43325 , n43345 );
buf ( n43347 , n25020 );
not ( n43348 , n43347 );
nand ( n43349 , n43315 , n43329 );
not ( n43350 , n43349 );
nand ( n43351 , n43350 , n43313 );
nor ( n43352 , n43351 , n43302 );
nand ( n43353 , n43352 , n43285 );
buf ( n43354 , n14683 );
buf ( n43355 , n43354 );
and ( n43356 , n43353 , n43355 );
not ( n43357 , n43353 );
not ( n43358 , n43355 );
and ( n43359 , n43357 , n43358 );
nor ( n43360 , n43356 , n43359 );
buf ( n43361 , n43360 );
not ( n43362 , n43361 );
or ( n43363 , n42975 , n43362 );
nand ( n43364 , n43193 , n24813 );
nand ( n43365 , n43363 , n43364 );
buf ( n43366 , n43365 );
not ( n43367 , n43366 );
not ( n43368 , n43367 );
or ( n43369 , n43348 , n43368 );
buf ( n43370 , n14747 );
not ( n43371 , n43370 );
and ( n43372 , n43371 , n43355 );
not ( n43373 , n43371 );
and ( n43374 , n43373 , n43358 );
nor ( n43375 , n43372 , n43374 );
not ( n43376 , n43375 );
nor ( n43377 , n43349 , n43355 );
and ( n43378 , n43303 , n43313 , n43377 );
nand ( n43379 , n43285 , n43378 );
not ( n43380 , n43379 );
or ( n43381 , n43376 , n43380 );
or ( n43382 , n43379 , n43375 );
nand ( n43383 , n43381 , n43382 );
buf ( n43384 , n43383 );
not ( n43385 , n43384 );
not ( n43386 , n43140 );
or ( n43387 , n43385 , n43386 );
not ( n43388 , n14759 );
nand ( n43389 , n43387 , n43388 );
buf ( n43390 , n43389 );
buf ( n43391 , n38843 );
not ( n43392 , n43391 );
nand ( n43393 , n43390 , n43392 );
nand ( n43394 , n43369 , n43393 );
nor ( n43395 , n43346 , n43394 );
not ( n43396 , n24485 );
not ( n43397 , n43193 );
or ( n43398 , n43396 , n43397 );
not ( n43399 , n43306 );
nor ( n43400 , n43399 , n43311 );
nand ( n43401 , n43285 , n43303 , n43400 );
buf ( n43402 , n43307 );
not ( n43403 , n43402 );
and ( n43404 , n43401 , n43403 );
not ( n43405 , n43401 );
and ( n43406 , n43405 , n43402 );
nor ( n43407 , n43404 , n43406 );
buf ( n43408 , n43407 );
not ( n43409 , n43408 );
or ( n43410 , n43005 , n43409 );
nand ( n43411 , n43398 , n43410 );
buf ( n43412 , n43411 );
buf ( n43413 , n24891 );
not ( n43414 , n43413 );
nor ( n43415 , n43412 , n43414 );
nor ( n43416 , n43302 , n43399 );
nand ( n43417 , n43285 , n43416 );
and ( n43418 , n43417 , n43311 );
not ( n43419 , n43417 );
and ( n43420 , n43419 , n43310 );
nor ( n43421 , n43418 , n43420 );
buf ( n43422 , n43421 );
not ( n43423 , n43422 );
or ( n43424 , n43186 , n43423 );
nand ( n43425 , n42975 , n14057 );
nand ( n43426 , n43424 , n43425 );
buf ( n43427 , n43426 );
buf ( n43428 , n24538 );
not ( n43429 , n43428 );
nor ( n43430 , n43427 , n43429 );
nor ( n43431 , n43415 , n43430 );
not ( n43432 , n43431 );
not ( n43433 , n42975 );
not ( n43434 , n14796 );
or ( n43435 , n43433 , n43434 );
nand ( n43436 , n43285 , n43303 , n43304 );
not ( n43437 , n43305 );
and ( n43438 , n43436 , n43437 );
not ( n43439 , n43436 );
and ( n43440 , n43439 , n43305 );
nor ( n43441 , n43438 , n43440 );
buf ( n43442 , n43441 );
not ( n43443 , n43442 );
or ( n43444 , n42975 , n43443 );
nand ( n43445 , n43435 , n43444 );
buf ( n43446 , n43445 );
buf ( n43447 , n15509 );
not ( n43448 , n43447 );
nor ( n43449 , n43446 , n43448 );
not ( n43450 , n43449 );
not ( n43451 , n13976 );
not ( n43452 , n43451 );
not ( n43453 , n43452 );
not ( n43454 , n43005 );
or ( n43455 , n43453 , n43454 );
nand ( n43456 , n43285 , n43303 );
not ( n43457 , n43304 );
and ( n43458 , n43456 , n43457 );
not ( n43459 , n43456 );
and ( n43460 , n43459 , n43304 );
nor ( n43461 , n43458 , n43460 );
buf ( n43462 , n43461 );
not ( n43463 , n43462 );
or ( n43464 , n43028 , n43463 );
nand ( n43465 , n43455 , n43464 );
buf ( n43466 , n43465 );
not ( n43467 , n43466 );
buf ( n43468 , n15557 );
nand ( n43469 , n43467 , n43468 );
nand ( n43470 , n43450 , n43469 );
nor ( n43471 , n43432 , n43470 );
nand ( n43472 , n43395 , n43471 );
not ( n43473 , n23822 );
not ( n43474 , n43473 );
not ( n43475 , n43474 );
not ( n43476 , n43025 );
or ( n43477 , n43475 , n43476 );
not ( n43478 , n43297 );
buf ( n43479 , n43288 );
and ( n43480 , n43479 , n43289 );
nand ( n43481 , n43478 , n43480 );
and ( n43482 , n43299 , n43287 );
nand ( n43483 , n43482 , n43290 );
nor ( n43484 , n43481 , n43483 );
nand ( n43485 , n43285 , n43484 );
not ( n43486 , n43298 );
and ( n43487 , n43485 , n43486 );
not ( n43488 , n43485 );
and ( n43489 , n43488 , n43298 );
nor ( n43490 , n43487 , n43489 );
buf ( n43491 , n43490 );
not ( n43492 , n43491 );
or ( n43493 , n43028 , n43492 );
nand ( n43494 , n43477 , n43493 );
buf ( n43495 , n43494 );
buf ( n43496 , n32694 );
not ( n43497 , n43496 );
nor ( n43498 , n43495 , n43497 );
buf ( n43499 , n32617 );
not ( n43500 , n43499 );
not ( n43501 , n43186 );
or ( n43502 , n43500 , n43501 );
not ( n43503 , n43482 );
nor ( n43504 , n43503 , n43481 );
nand ( n43505 , n43285 , n43504 );
not ( n43506 , n43290 );
and ( n43507 , n43505 , n43506 );
not ( n43508 , n43505 );
and ( n43509 , n43508 , n43290 );
nor ( n43510 , n43507 , n43509 );
buf ( n43511 , n43510 );
not ( n43512 , n43511 );
or ( n43513 , n43186 , n43512 );
nand ( n43514 , n43502 , n43513 );
buf ( n43515 , n43514 );
not ( n43516 , n33043 );
buf ( n43517 , n43516 );
not ( n43518 , n43517 );
nor ( n43519 , n43515 , n43518 );
nor ( n43520 , n43498 , n43519 );
not ( n43521 , n43287 );
nor ( n43522 , n43481 , n43521 );
nand ( n43523 , n43285 , n43522 );
not ( n43524 , n43299 );
and ( n43525 , n43523 , n43524 );
not ( n43526 , n43523 );
and ( n43527 , n43526 , n43299 );
nor ( n43528 , n43525 , n43527 );
buf ( n43529 , n43528 );
not ( n43530 , n43529 );
or ( n43531 , n43005 , n43530 );
not ( n43532 , n32980 );
not ( n43533 , n43532 );
nand ( n43534 , n42929 , n43533 );
nand ( n43535 , n43531 , n43534 );
buf ( n43536 , n43535 );
buf ( n43537 , n20788 );
not ( n43538 , n43537 );
nor ( n43539 , n43536 , n43538 );
not ( n43540 , n31331 );
buf ( n43541 , n43540 );
not ( n43542 , n43541 );
buf ( n43543 , n20713 );
not ( n43544 , n43543 );
not ( n43545 , n43097 );
or ( n43546 , n43544 , n43545 );
not ( n43547 , n43481 );
nand ( n43548 , n43547 , n43285 );
and ( n43549 , n43548 , n43521 );
not ( n43550 , n43548 );
and ( n43551 , n43550 , n43287 );
nor ( n43552 , n43549 , n43551 );
buf ( n43553 , n43552 );
not ( n43554 , n43553 );
or ( n43555 , n43005 , n43554 );
nand ( n43556 , n43546 , n43555 );
buf ( n43557 , n43556 );
nor ( n43558 , n43542 , n43557 );
nor ( n43559 , n43539 , n43558 );
nand ( n43560 , n43520 , n43559 );
not ( n43561 , n43560 );
buf ( n43562 , n31303 );
not ( n43563 , n43562 );
or ( n43564 , n43185 , n43563 );
not ( n43565 , n43289 );
nor ( n43566 , n43297 , n43565 );
nand ( n43567 , n43285 , n43566 );
xnor ( n43568 , n43567 , n43479 );
buf ( n43569 , n43568 );
nand ( n43570 , n43024 , n43569 );
nand ( n43571 , n43564 , n43570 );
buf ( n43572 , n43571 );
buf ( n43573 , n32326 );
not ( n43574 , n43573 );
nor ( n43575 , n43572 , n43574 );
buf ( n43576 , n29042 );
not ( n43577 , n43576 );
not ( n43578 , n42975 );
or ( n43579 , n43577 , n43578 );
not ( n43580 , n43297 );
nand ( n43581 , n43580 , n43285 );
and ( n43582 , n43581 , n43565 );
not ( n43583 , n43581 );
and ( n43584 , n43583 , n43289 );
nor ( n43585 , n43582 , n43584 );
buf ( n43586 , n43585 );
not ( n43587 , n43586 );
or ( n43588 , n42975 , n43587 );
nand ( n43589 , n43579 , n43588 );
buf ( n43590 , n43589 );
buf ( n43591 , n23769 );
not ( n43592 , n43591 );
nor ( n43593 , n43590 , n43592 );
nor ( n43594 , n43575 , n43593 );
not ( n43595 , n43594 );
buf ( n43596 , n31174 );
not ( n43597 , n43596 );
buf ( n43598 , n23401 );
not ( n43599 , n43598 );
not ( n43600 , n43186 );
or ( n43601 , n43599 , n43600 );
buf ( n43602 , n43296 );
not ( n43603 , n43602 );
not ( n43604 , n43285 );
not ( n43605 , n43604 );
or ( n43606 , n43603 , n43605 );
or ( n43607 , n43604 , n43602 );
nand ( n43608 , n43606 , n43607 );
buf ( n43609 , n43608 );
not ( n43610 , n43609 );
or ( n43611 , n43028 , n43610 );
nand ( n43612 , n43601 , n43611 );
buf ( n43613 , n43612 );
not ( n43614 , n43613 );
not ( n43615 , n43614 );
or ( n43616 , n43597 , n43615 );
not ( n43617 , n23774 );
not ( n43618 , n43617 );
not ( n43619 , n43618 );
not ( n43620 , n43193 );
or ( n43621 , n43619 , n43620 );
nand ( n43622 , n43285 , n43602 );
buf ( n43623 , n43294 );
not ( n43624 , n43623 );
and ( n43625 , n43622 , n43624 );
not ( n43626 , n43622 );
and ( n43627 , n43626 , n43623 );
nor ( n43628 , n43625 , n43627 );
buf ( n43629 , n43628 );
not ( n43630 , n43629 );
or ( n43631 , n42929 , n43630 );
nand ( n43632 , n43621 , n43631 );
buf ( n43633 , n43632 );
buf ( n43634 , n23446 );
not ( n43635 , n43634 );
nor ( n43636 , n43633 , n43635 );
not ( n43637 , n43636 );
nand ( n43638 , n43616 , n43637 );
nor ( n43639 , n43595 , n43638 );
nand ( n43640 , n43561 , n43639 );
nor ( n43641 , n43472 , n43640 );
and ( n43642 , n43272 , n43641 );
not ( n43643 , n43596 );
nand ( n43644 , n43643 , n43613 );
nand ( n43645 , n43633 , n43635 );
and ( n43646 , n43644 , n43645 );
nor ( n43647 , n43646 , n43636 );
and ( n43648 , n43594 , n43647 );
nand ( n43649 , n43590 , n43592 );
or ( n43650 , n43575 , n43649 );
nand ( n43651 , n43572 , n43574 );
nand ( n43652 , n43650 , n43651 );
nor ( n43653 , n43648 , n43652 );
not ( n43654 , n43653 );
not ( n43655 , n43560 );
and ( n43656 , n43654 , n43655 );
not ( n43657 , n43520 );
not ( n43658 , n43541 );
nand ( n43659 , n43658 , n43557 );
or ( n43660 , n43539 , n43659 );
nand ( n43661 , n43536 , n43538 );
nand ( n43662 , n43660 , n43661 );
not ( n43663 , n43662 );
or ( n43664 , n43657 , n43663 );
not ( n43665 , n43498 );
nand ( n43666 , n43515 , n43518 );
not ( n43667 , n43666 );
and ( n43668 , n43665 , n43667 );
and ( n43669 , n43495 , n43497 );
nor ( n43670 , n43668 , n43669 );
nand ( n43671 , n43664 , n43670 );
nor ( n43672 , n43656 , n43671 );
or ( n43673 , n43672 , n43472 );
not ( n43674 , n43431 );
not ( n43675 , n43468 );
nand ( n43676 , n43675 , n43466 );
or ( n43677 , n43449 , n43676 );
nand ( n43678 , n43446 , n43448 );
nand ( n43679 , n43677 , n43678 );
not ( n43680 , n43679 );
or ( n43681 , n43674 , n43680 );
not ( n43682 , n43415 );
nand ( n43683 , n43427 , n43429 );
not ( n43684 , n43683 );
and ( n43685 , n43682 , n43684 );
and ( n43686 , n43412 , n43414 );
nor ( n43687 , n43685 , n43686 );
nand ( n43688 , n43681 , n43687 );
and ( n43689 , n43688 , n43395 );
not ( n43690 , n43322 );
nor ( n43691 , n43690 , n43273 );
and ( n43692 , n43345 , n43691 );
not ( n43693 , n43342 );
nor ( n43694 , n43693 , n43344 );
nor ( n43695 , n43692 , n43694 );
or ( n43696 , n43695 , n43394 );
not ( n43697 , n43366 );
nor ( n43698 , n43697 , n43347 );
and ( n43699 , n43698 , n43393 );
nor ( n43700 , n43390 , n43392 );
nor ( n43701 , n43699 , n43700 );
nand ( n43702 , n43696 , n43701 );
nor ( n43703 , n43689 , n43702 );
nand ( n43704 , n43673 , n43703 );
nor ( n43705 , n43642 , n43704 );
buf ( n43706 , n43705 );
and ( n43707 , n17540 , n43706 );
not ( n43708 , n17540 );
not ( n43709 , n43706 );
and ( n43710 , n43708 , n43709 );
nor ( n43711 , n43707 , n43710 );
not ( n43712 , n14886 );
and ( n43713 , n43711 , n43712 );
buf ( n43714 , n16151 );
not ( n43715 , n43714 );
buf ( n43716 , n27159 );
nor ( n43717 , n43715 , n43716 );
not ( n43718 , n43717 );
buf ( n43719 , n16650 );
not ( n43720 , n43719 );
buf ( n43721 , n27726 );
nor ( n43722 , n43720 , n43721 );
not ( n43723 , n43721 );
nor ( n43724 , n43723 , n43719 );
or ( n43725 , n43722 , n43724 );
not ( n43726 , n43725 );
or ( n43727 , n43718 , n43726 );
or ( n43728 , n43725 , n43717 );
nand ( n43729 , n43727 , n43728 );
not ( n43730 , n43722 );
buf ( n43731 , n16614 );
not ( n43732 , n43731 );
buf ( n43733 , n26495 );
nor ( n43734 , n43732 , n43733 );
not ( n43735 , n43733 );
nor ( n43736 , n43735 , n43731 );
or ( n43737 , n43734 , n43736 );
not ( n43738 , n43737 );
or ( n43739 , n43730 , n43738 );
or ( n43740 , n43737 , n43722 );
nand ( n43741 , n43739 , n43740 );
not ( n43742 , n43734 );
buf ( n43743 , n16509 );
not ( n43744 , n43743 );
buf ( n43745 , n34924 );
nor ( n43746 , n43744 , n43745 );
not ( n43747 , n43745 );
nor ( n43748 , n43747 , n43743 );
or ( n43749 , n43746 , n43748 );
not ( n43750 , n43749 );
or ( n43751 , n43742 , n43750 );
or ( n43752 , n43749 , n43734 );
nand ( n43753 , n43751 , n43752 );
buf ( n43754 , n43293 );
not ( n43755 , n43754 );
buf ( n43756 , n23445 );
nor ( n43757 , n43755 , n43756 );
not ( n43758 , n43757 );
buf ( n43759 , n17011 );
not ( n43760 , n43759 );
buf ( n43761 , n23767 );
nor ( n43762 , n43760 , n43761 );
not ( n43763 , n43761 );
nor ( n43764 , n43763 , n43759 );
or ( n43765 , n43762 , n43764 );
not ( n43766 , n43765 );
or ( n43767 , n43758 , n43766 );
or ( n43768 , n43765 , n43757 );
nand ( n43769 , n43767 , n43768 );
nand ( n43770 , n43729 , n43741 , n43753 , n43769 );
not ( n43771 , n43746 );
buf ( n43772 , n15839 );
not ( n43773 , n43772 );
buf ( n43774 , n42994 );
nor ( n43775 , n43773 , n43774 );
not ( n43776 , n43774 );
nor ( n43777 , n43776 , n43772 );
or ( n43778 , n43775 , n43777 );
not ( n43779 , n43778 );
or ( n43780 , n43771 , n43779 );
or ( n43781 , n43778 , n43746 );
nand ( n43782 , n43780 , n43781 );
not ( n43783 , n43775 );
buf ( n43784 , n43295 );
not ( n43785 , n43784 );
buf ( n43786 , n31171 );
nor ( n43787 , n43785 , n43786 );
not ( n43788 , n43786 );
nor ( n43789 , n43788 , n43784 );
or ( n43790 , n43787 , n43789 );
not ( n43791 , n43790 );
or ( n43792 , n43783 , n43791 );
or ( n43793 , n43790 , n43775 );
nand ( n43794 , n43792 , n43793 );
not ( n43795 , n43787 );
not ( n43796 , n43756 );
nor ( n43797 , n43796 , n43754 );
or ( n43798 , n43757 , n43797 );
not ( n43799 , n43798 );
or ( n43800 , n43795 , n43799 );
or ( n43801 , n43798 , n43787 );
nand ( n43802 , n43800 , n43801 );
buf ( n43803 , n14747 );
buf ( n43804 , n38843 );
xor ( n43805 , n43803 , n43804 );
not ( n43806 , n43805 );
buf ( n43807 , n43354 );
not ( n43808 , n43807 );
buf ( n43809 , n25020 );
or ( n43810 , n43808 , n43809 );
not ( n43811 , n43810 );
and ( n43812 , n43806 , n43811 );
and ( n43813 , n43805 , n43810 );
nor ( n43814 , n43812 , n43813 );
nand ( n43815 , n43782 , n43794 , n43802 , n43814 );
nor ( n43816 , n43770 , n43815 );
not ( n43817 , n43762 );
buf ( n43818 , n15733 );
not ( n43819 , n43818 );
buf ( n43820 , n32325 );
nor ( n43821 , n43819 , n43820 );
not ( n43822 , n43820 );
nor ( n43823 , n43822 , n43818 );
or ( n43824 , n43821 , n43823 );
not ( n43825 , n43824 );
or ( n43826 , n43817 , n43825 );
or ( n43827 , n43824 , n43762 );
nand ( n43828 , n43826 , n43827 );
not ( n43829 , n43821 );
buf ( n43830 , n43286 );
buf ( n43831 , n43830 );
not ( n43832 , n43831 );
buf ( n43833 , n31329 );
nor ( n43834 , n43832 , n43833 );
not ( n43835 , n43833 );
nor ( n43836 , n43835 , n43831 );
or ( n43837 , n43834 , n43836 );
not ( n43838 , n43837 );
or ( n43839 , n43829 , n43838 );
or ( n43840 , n43837 , n43821 );
nand ( n43841 , n43839 , n43840 );
not ( n43842 , n43834 );
buf ( n43843 , n16027 );
not ( n43844 , n43843 );
buf ( n43845 , n20786 );
nor ( n43846 , n43844 , n43845 );
not ( n43847 , n43846 );
not ( n43848 , n43843 );
nand ( n43849 , n43848 , n43845 );
nand ( n43850 , n43847 , n43849 );
not ( n43851 , n43850 );
or ( n43852 , n43842 , n43851 );
or ( n43853 , n43850 , n43834 );
nand ( n43854 , n43852 , n43853 );
not ( n43855 , n43846 );
buf ( n43856 , n16016 );
not ( n43857 , n43856 );
buf ( n43858 , n33041 );
nor ( n43859 , n43857 , n43858 );
not ( n43860 , n43859 );
not ( n43861 , n43856 );
nand ( n43862 , n43861 , n43858 );
nand ( n43863 , n43860 , n43862 );
not ( n43864 , n43863 );
or ( n43865 , n43855 , n43864 );
or ( n43866 , n43863 , n43846 );
nand ( n43867 , n43865 , n43866 );
nand ( n43868 , n43828 , n43841 , n43854 , n43867 );
not ( n43869 , n43859 );
buf ( n43870 , n15966 );
not ( n43871 , n43870 );
buf ( n43872 , n32692 );
nor ( n43873 , n43871 , n43872 );
not ( n43874 , n43872 );
nor ( n43875 , n43874 , n43870 );
or ( n43876 , n43873 , n43875 );
not ( n43877 , n43876 );
or ( n43878 , n43869 , n43877 );
or ( n43879 , n43876 , n43859 );
nand ( n43880 , n43878 , n43879 );
buf ( n43881 , n15561 );
not ( n43882 , n43881 );
buf ( n43883 , n15557 );
nor ( n43884 , n43882 , n43883 );
not ( n43885 , n43884 );
buf ( n43886 , n15509 );
not ( n43887 , n43886 );
buf ( n43888 , n15513 );
not ( n43889 , n43888 );
not ( n43890 , n43889 );
or ( n43891 , n43887 , n43890 );
nor ( n43892 , n43889 , n43886 );
not ( n43893 , n43892 );
nand ( n43894 , n43891 , n43893 );
not ( n43895 , n43894 );
or ( n43896 , n43885 , n43895 );
or ( n43897 , n43894 , n43884 );
nand ( n43898 , n43896 , n43897 );
not ( n43899 , n43892 );
buf ( n43900 , n24538 );
not ( n43901 , n43900 );
buf ( n43902 , n43309 );
not ( n43903 , n43902 );
not ( n43904 , n43903 );
or ( n43905 , n43901 , n43904 );
nor ( n43906 , n43903 , n43900 );
not ( n43907 , n43906 );
nand ( n43908 , n43905 , n43907 );
not ( n43909 , n43908 );
or ( n43910 , n43899 , n43909 );
or ( n43911 , n43908 , n43892 );
nand ( n43912 , n43910 , n43911 );
not ( n43913 , n43906 );
buf ( n43914 , n24891 );
not ( n43915 , n43914 );
buf ( n43916 , n30326 );
not ( n43917 , n43916 );
not ( n43918 , n43917 );
or ( n43919 , n43915 , n43918 );
nor ( n43920 , n43917 , n43914 );
not ( n43921 , n43920 );
nand ( n43922 , n43919 , n43921 );
not ( n43923 , n43922 );
or ( n43924 , n43913 , n43923 );
or ( n43925 , n43922 , n43906 );
nand ( n43926 , n43924 , n43925 );
nand ( n43927 , n43880 , n43898 , n43912 , n43926 );
nor ( n43928 , n43868 , n43927 );
not ( n43929 , n43920 );
buf ( n43930 , n30322 );
not ( n43931 , n43930 );
buf ( n43932 , n24937 );
nor ( n43933 , n43931 , n43932 );
not ( n43934 , n43933 );
not ( n43935 , n43930 );
nand ( n43936 , n43935 , n43932 );
nand ( n43937 , n43934 , n43936 );
not ( n43938 , n43937 );
or ( n43939 , n43929 , n43938 );
or ( n43940 , n43937 , n43920 );
nand ( n43941 , n43939 , n43940 );
not ( n43942 , n43933 );
buf ( n43943 , n34432 );
not ( n43944 , n43943 );
buf ( n43945 , n24939 );
nor ( n43946 , n43944 , n43945 );
not ( n43947 , n43945 );
nor ( n43948 , n43947 , n43943 );
or ( n43949 , n43946 , n43948 );
not ( n43950 , n43949 );
or ( n43951 , n43942 , n43950 );
or ( n43952 , n43949 , n43933 );
nand ( n43953 , n43951 , n43952 );
buf ( n43954 , n42940 );
buf ( n43955 , n43954 );
not ( n43956 , n43955 );
buf ( n43957 , n32957 );
nor ( n43958 , n43956 , n43957 );
not ( n43959 , n43958 );
buf ( n43960 , n16485 );
not ( n43961 , n43960 );
buf ( n43962 , n34666 );
nor ( n43963 , n43961 , n43962 );
not ( n43964 , n43962 );
nor ( n43965 , n43964 , n43960 );
or ( n43966 , n43963 , n43965 );
not ( n43967 , n43966 );
or ( n43968 , n43959 , n43967 );
or ( n43969 , n43966 , n43958 );
nand ( n43970 , n43968 , n43969 );
nand ( n43971 , n43941 , n43953 , n43970 );
not ( n43972 , n43883 );
not ( n43973 , n43882 );
or ( n43974 , n43972 , n43973 );
not ( n43975 , n43884 );
nand ( n43976 , n43974 , n43975 );
not ( n43977 , n43976 );
not ( n43978 , n43873 );
and ( n43979 , n43977 , n43978 );
and ( n43980 , n43976 , n43873 );
nor ( n43981 , n43979 , n43980 );
not ( n43982 , n43808 );
not ( n43983 , n43809 );
or ( n43984 , n43982 , n43983 );
nand ( n43985 , n43984 , n43810 );
not ( n43986 , n43985 );
not ( n43987 , n43946 );
and ( n43988 , n43986 , n43987 );
and ( n43989 , n43985 , n43946 );
nor ( n43990 , n43988 , n43989 );
nor ( n43991 , n43971 , n43981 , n43990 );
buf ( n43992 , n17202 );
not ( n43993 , n43992 );
buf ( n43994 , n32403 );
nor ( n43995 , n43993 , n43994 );
not ( n43996 , n43995 );
buf ( n43997 , n16212 );
not ( n43998 , n43997 );
buf ( n43999 , n20941 );
nor ( n44000 , n43998 , n43999 );
not ( n44001 , n43999 );
nor ( n44002 , n44001 , n43997 );
or ( n44003 , n44000 , n44002 );
not ( n44004 , n44003 );
or ( n44005 , n43996 , n44004 );
or ( n44006 , n44003 , n43995 );
nand ( n44007 , n44005 , n44006 );
not ( n44008 , n43963 );
buf ( n44009 , n16440 );
not ( n44010 , n44009 );
buf ( n44011 , n24722 );
nor ( n44012 , n44010 , n44011 );
not ( n44013 , n44011 );
nor ( n44014 , n44013 , n44009 );
or ( n44015 , n44012 , n44014 );
not ( n44016 , n44015 );
or ( n44017 , n44008 , n44016 );
or ( n44018 , n44015 , n43963 );
nand ( n44019 , n44017 , n44018 );
not ( n44020 , n44000 );
not ( n44021 , n43717 );
not ( n44022 , n43714 );
nand ( n44023 , n44022 , n43716 );
nand ( n44024 , n44021 , n44023 );
not ( n44025 , n44024 );
or ( n44026 , n44020 , n44025 );
or ( n44027 , n44024 , n44000 );
nand ( n44028 , n44026 , n44027 );
buf ( n44029 , n16766 );
buf ( n44030 , n42936 );
xnor ( n44031 , n44029 , n44030 );
not ( n44032 , n34721 );
buf ( n44033 , n44032 );
and ( n44034 , n44031 , n44033 );
nor ( n44035 , n44031 , n44033 );
buf ( n44036 , n36637 );
buf ( n44037 , n43173 );
xnor ( n44038 , n44036 , n44037 );
buf ( n44039 , n20679 );
not ( n44040 , n44039 );
buf ( n44041 , n43162 );
not ( n44042 , n44041 );
or ( n44043 , n44040 , n44042 );
or ( n44044 , n44041 , n44039 );
nand ( n44045 , n44043 , n44044 );
buf ( n44046 , n21685 );
buf ( n44047 , n14542 );
xnor ( n44048 , n44046 , n44047 );
nand ( n44049 , n44038 , n44045 , n44048 );
nor ( n44050 , n44034 , n44035 , n44049 );
nand ( n44051 , n44007 , n44019 , n44028 , n44050 );
not ( n44052 , n44030 );
nor ( n44053 , n44052 , n44033 );
not ( n44054 , n44053 );
not ( n44055 , n43957 );
nor ( n44056 , n44055 , n43955 );
or ( n44057 , n43958 , n44056 );
not ( n44058 , n44057 );
or ( n44059 , n44054 , n44058 );
or ( n44060 , n44057 , n44053 );
nand ( n44061 , n44059 , n44060 );
buf ( n44062 , n16332 );
not ( n44063 , n44062 );
buf ( n44064 , n37913 );
nor ( n44065 , n44063 , n44064 );
not ( n44066 , n44065 );
buf ( n44067 , n16296 );
not ( n44068 , n44067 );
buf ( n44069 , n32190 );
nor ( n44070 , n44068 , n44069 );
not ( n44071 , n44070 );
not ( n44072 , n44067 );
nand ( n44073 , n44072 , n44069 );
nand ( n44074 , n44071 , n44073 );
not ( n44075 , n44074 );
or ( n44076 , n44066 , n44075 );
or ( n44077 , n44074 , n44065 );
nand ( n44078 , n44076 , n44077 );
not ( n44079 , n44012 );
not ( n44080 , n44065 );
not ( n44081 , n44062 );
nand ( n44082 , n44081 , n44064 );
nand ( n44083 , n44080 , n44082 );
not ( n44084 , n44083 );
or ( n44085 , n44079 , n44084 );
or ( n44086 , n44083 , n44012 );
nand ( n44087 , n44085 , n44086 );
not ( n44088 , n44070 );
not ( n44089 , n43995 );
not ( n44090 , n43992 );
nand ( n44091 , n44090 , n43994 );
nand ( n44092 , n44089 , n44091 );
not ( n44093 , n44092 );
or ( n44094 , n44088 , n44093 );
or ( n44095 , n44092 , n44070 );
nand ( n44096 , n44094 , n44095 );
nand ( n44097 , n44061 , n44078 , n44087 , n44096 );
nor ( n44098 , n44051 , n44097 );
and ( n44099 , n43816 , n43928 , n43991 , n44098 );
buf ( n44100 , n44099 );
nor ( n44101 , n44100 , n43712 , n14905 );
nor ( n44102 , n43713 , n44101 );
nor ( n44103 , n22898 , n14900 );
not ( n44104 , n44103 );
or ( n44105 , n44102 , n44104 );
not ( n44106 , n43712 );
buf ( n44107 , n25020 );
not ( n44108 , n44107 );
not ( n44109 , n44108 );
buf ( n44110 , n24815 );
not ( n44111 , n44110 );
or ( n44112 , n44109 , n44111 );
buf ( n44113 , n24737 );
not ( n44114 , n44113 );
buf ( n44115 , n38843 );
nand ( n44116 , n44114 , n44115 );
nand ( n44117 , n44112 , n44116 );
buf ( n44118 , n24937 );
not ( n44119 , n44118 );
not ( n44120 , n44119 );
not ( n44121 , n43275 );
buf ( n44122 , n44121 );
not ( n44123 , n44122 );
or ( n44124 , n44120 , n44123 );
not ( n44125 , n43338 );
buf ( n44126 , n44125 );
buf ( n44127 , n24939 );
not ( n44128 , n44127 );
nand ( n44129 , n44126 , n44128 );
nand ( n44130 , n44124 , n44129 );
nor ( n44131 , n44117 , n44130 );
buf ( n44132 , n24538 );
not ( n44133 , n44132 );
not ( n44134 , n44133 );
buf ( n44135 , n14057 );
buf ( n44136 , n44135 );
not ( n44137 , n44136 );
or ( n44138 , n44134 , n44137 );
buf ( n44139 , n24485 );
buf ( n44140 , n44139 );
buf ( n44141 , n24891 );
not ( n44142 , n44141 );
nand ( n44143 , n44140 , n44142 );
nand ( n44144 , n44138 , n44143 );
buf ( n44145 , n15557 );
not ( n44146 , n44145 );
not ( n44147 , n44146 );
not ( n44148 , n43451 );
buf ( n44149 , n44148 );
not ( n44150 , n44149 );
or ( n44151 , n44147 , n44150 );
buf ( n44152 , n14796 );
buf ( n44153 , n15509 );
not ( n44154 , n44153 );
nand ( n44155 , n44152 , n44154 );
nand ( n44156 , n44151 , n44155 );
nor ( n44157 , n44144 , n44156 );
nand ( n44158 , n44131 , n44157 );
buf ( n44159 , n34925 );
not ( n44160 , n44159 );
not ( n44161 , n44160 );
buf ( n44162 , n42923 );
not ( n44163 , n44162 );
or ( n44164 , n44161 , n44163 );
buf ( n44165 , n42995 );
not ( n44166 , n44165 );
buf ( n44167 , n42973 );
nand ( n44168 , n44166 , n44167 );
nand ( n44169 , n44164 , n44168 );
buf ( n44170 , n27727 );
not ( n44171 , n44170 );
not ( n44172 , n44171 );
not ( n44173 , n43021 );
buf ( n44174 , n44173 );
not ( n44175 , n44174 );
or ( n44176 , n44172 , n44175 );
buf ( n44177 , n26496 );
not ( n44178 , n44177 );
buf ( n44179 , n43001 );
nand ( n44180 , n44178 , n44179 );
nand ( n44181 , n44176 , n44180 );
nor ( n44182 , n44169 , n44181 );
buf ( n44183 , n20942 );
not ( n44184 , n44183 );
not ( n44185 , n44184 );
not ( n44186 , n43070 );
buf ( n44187 , n44186 );
not ( n44188 , n44187 );
or ( n44189 , n44185 , n44188 );
buf ( n44190 , n27160 );
not ( n44191 , n44190 );
not ( n44192 , n43040 );
buf ( n44193 , n44192 );
nand ( n44194 , n44191 , n44193 );
nand ( n44195 , n44189 , n44194 );
buf ( n44196 , n32191 );
not ( n44197 , n44196 );
not ( n44198 , n44197 );
buf ( n44199 , n43079 );
not ( n44200 , n44199 );
or ( n44201 , n44198 , n44200 );
buf ( n44202 , n32404 );
not ( n44203 , n44202 );
not ( n44204 , n43094 );
buf ( n44205 , n44204 );
nand ( n44206 , n44203 , n44205 );
nand ( n44207 , n44201 , n44206 );
nor ( n44208 , n44195 , n44207 );
buf ( n44209 , n37914 );
not ( n44210 , n44209 );
buf ( n44211 , n43221 );
nand ( n44212 , n44210 , n44211 );
buf ( n44213 , n24722 );
not ( n44214 , n44213 );
buf ( n44215 , n43237 );
nand ( n44216 , n44214 , n44215 );
and ( n44217 , n44212 , n44216 );
not ( n44218 , n44217 );
buf ( n44219 , n34719 );
not ( n44220 , n44219 );
buf ( n44221 , n43135 );
nand ( n44222 , n44220 , n44221 );
buf ( n44223 , n43160 );
not ( n44224 , n44223 );
buf ( n44225 , n20678 );
nor ( n44226 , n44224 , n44225 );
buf ( n44227 , n14542 );
buf ( n44228 , n21683 );
not ( n44229 , n44228 );
and ( n44230 , n44227 , n44229 );
or ( n44231 , n44226 , n44230 );
or ( n44232 , n44227 , n44229 );
nand ( n44233 , n44231 , n44232 );
buf ( n44234 , n36636 );
not ( n44235 , n44234 );
buf ( n44236 , n43172 );
nand ( n44237 , n44235 , n44236 );
nand ( n44238 , n44222 , n44233 , n44237 );
not ( n44239 , n44234 );
nor ( n44240 , n44239 , n44236 );
nand ( n44241 , n44222 , n44240 );
not ( n44242 , n44221 );
nand ( n44243 , n44242 , n44219 );
nand ( n44244 , n44238 , n44241 , n44243 );
buf ( n44245 , n34667 );
not ( n44246 , n44245 );
buf ( n44247 , n43194 );
nand ( n44248 , n44246 , n44247 );
buf ( n44249 , n32957 );
not ( n44250 , n44249 );
buf ( n44251 , n43202 );
nand ( n44252 , n44250 , n44251 );
and ( n44253 , n44244 , n44248 , n44252 );
not ( n44254 , n44253 );
or ( n44255 , n44218 , n44254 );
not ( n44256 , n44249 );
nor ( n44257 , n44256 , n44251 );
not ( n44258 , n44257 );
not ( n44259 , n44248 );
or ( n44260 , n44258 , n44259 );
not ( n44261 , n44247 );
nand ( n44262 , n44261 , n44245 );
nand ( n44263 , n44260 , n44262 );
and ( n44264 , n44217 , n44263 );
not ( n44265 , n44213 );
nor ( n44266 , n44265 , n44215 );
not ( n44267 , n44266 );
not ( n44268 , n44212 );
or ( n44269 , n44267 , n44268 );
not ( n44270 , n44211 );
nand ( n44271 , n44270 , n44209 );
nand ( n44272 , n44269 , n44271 );
nor ( n44273 , n44264 , n44272 );
nand ( n44274 , n44255 , n44273 );
and ( n44275 , n44182 , n44208 , n44274 );
not ( n44276 , n44182 );
nor ( n44277 , n44199 , n44197 );
not ( n44278 , n44277 );
not ( n44279 , n44206 );
or ( n44280 , n44278 , n44279 );
not ( n44281 , n44205 );
nand ( n44282 , n44281 , n44202 );
nand ( n44283 , n44280 , n44282 );
not ( n44284 , n44283 );
not ( n44285 , n44195 );
not ( n44286 , n44285 );
or ( n44287 , n44284 , n44286 );
nor ( n44288 , n44187 , n44184 );
and ( n44289 , n44194 , n44288 );
not ( n44290 , n44193 );
and ( n44291 , n44290 , n44190 );
nor ( n44292 , n44289 , n44291 );
nand ( n44293 , n44287 , n44292 );
not ( n44294 , n44293 );
or ( n44295 , n44276 , n44294 );
not ( n44296 , n44169 );
nor ( n44297 , n44174 , n44171 );
not ( n44298 , n44297 );
not ( n44299 , n44180 );
or ( n44300 , n44298 , n44299 );
not ( n44301 , n44179 );
nand ( n44302 , n44301 , n44177 );
nand ( n44303 , n44300 , n44302 );
and ( n44304 , n44296 , n44303 );
nor ( n44305 , n44162 , n44160 );
not ( n44306 , n44305 );
not ( n44307 , n44168 );
or ( n44308 , n44306 , n44307 );
not ( n44309 , n44167 );
nand ( n44310 , n44309 , n44165 );
nand ( n44311 , n44308 , n44310 );
nor ( n44312 , n44304 , n44311 );
nand ( n44313 , n44295 , n44312 );
nor ( n44314 , n44275 , n44313 );
buf ( n44315 , n33042 );
not ( n44316 , n44315 );
not ( n44317 , n44316 );
buf ( n44318 , n43499 );
not ( n44319 , n44318 );
or ( n44320 , n44317 , n44319 );
buf ( n44321 , n43474 );
buf ( n44322 , n32693 );
not ( n44323 , n44322 );
nand ( n44324 , n44321 , n44323 );
nand ( n44325 , n44320 , n44324 );
buf ( n44326 , n31330 );
not ( n44327 , n44326 );
not ( n44328 , n44327 );
buf ( n44329 , n43543 );
not ( n44330 , n44329 );
or ( n44331 , n44328 , n44330 );
buf ( n44332 , n43533 );
buf ( n44333 , n20787 );
not ( n44334 , n44333 );
nand ( n44335 , n44332 , n44334 );
nand ( n44336 , n44331 , n44335 );
nor ( n44337 , n44325 , n44336 );
buf ( n44338 , n23768 );
buf ( n44339 , n44338 );
not ( n44340 , n44339 );
not ( n44341 , n44340 );
not ( n44342 , n43576 );
not ( n44343 , n44342 );
buf ( n44344 , n44343 );
not ( n44345 , n44344 );
or ( n44346 , n44341 , n44345 );
buf ( n44347 , n43562 );
buf ( n44348 , n32326 );
not ( n44349 , n44348 );
nand ( n44350 , n44347 , n44349 );
nand ( n44351 , n44346 , n44350 );
buf ( n44352 , n31172 );
not ( n44353 , n44352 );
not ( n44354 , n44353 );
buf ( n44355 , n43598 );
not ( n44356 , n44355 );
or ( n44357 , n44354 , n44356 );
not ( n44358 , n43617 );
buf ( n44359 , n44358 );
buf ( n44360 , n23446 );
not ( n44361 , n44360 );
nand ( n44362 , n44359 , n44361 );
nand ( n44363 , n44357 , n44362 );
nor ( n44364 , n44351 , n44363 );
nand ( n44365 , n44337 , n44364 );
nor ( n44366 , n44158 , n44314 , n44365 );
nor ( n44367 , n44359 , n44361 );
nor ( n44368 , n44355 , n44353 );
or ( n44369 , n44367 , n44368 );
nand ( n44370 , n44369 , n44362 );
or ( n44371 , n44351 , n44370 );
nor ( n44372 , n44344 , n44340 );
and ( n44373 , n44350 , n44372 );
nor ( n44374 , n44347 , n44349 );
nor ( n44375 , n44373 , n44374 );
nand ( n44376 , n44371 , n44375 );
and ( n44377 , n44376 , n44337 );
nor ( n44378 , n44329 , n44327 );
and ( n44379 , n44335 , n44378 );
nor ( n44380 , n44332 , n44334 );
nor ( n44381 , n44379 , n44380 );
or ( n44382 , n44381 , n44325 );
nor ( n44383 , n44318 , n44316 );
and ( n44384 , n44324 , n44383 );
nor ( n44385 , n44321 , n44323 );
nor ( n44386 , n44384 , n44385 );
nand ( n44387 , n44382 , n44386 );
nor ( n44388 , n44377 , n44387 );
or ( n44389 , n44158 , n44388 );
nor ( n44390 , n44152 , n44154 );
nor ( n44391 , n44149 , n44146 );
or ( n44392 , n44390 , n44391 );
nand ( n44393 , n44392 , n44155 );
or ( n44394 , n44144 , n44393 );
nor ( n44395 , n44136 , n44133 );
and ( n44396 , n44143 , n44395 );
nor ( n44397 , n44140 , n44142 );
nor ( n44398 , n44396 , n44397 );
nand ( n44399 , n44394 , n44398 );
and ( n44400 , n44131 , n44399 );
nor ( n44401 , n44122 , n44119 );
and ( n44402 , n44129 , n44401 );
nor ( n44403 , n44126 , n44128 );
nor ( n44404 , n44402 , n44403 );
or ( n44405 , n44117 , n44404 );
nor ( n44406 , n44110 , n44108 );
and ( n44407 , n44116 , n44406 );
not ( n44408 , n44113 );
nor ( n44409 , n44408 , n44115 );
nor ( n44410 , n44407 , n44409 );
nand ( n44411 , n44405 , n44410 );
nor ( n44412 , n44400 , n44411 );
nand ( n44413 , n44389 , n44412 );
nor ( n44414 , n44366 , n44413 );
buf ( n44415 , n44414 );
not ( n44416 , n44415 );
or ( n44417 , n44106 , n44416 );
buf ( n44418 , n25020 );
not ( n44419 , n44418 );
buf ( n44420 , n24815 );
not ( n44421 , n44420 );
not ( n44422 , n44421 );
or ( n44423 , n44419 , n44422 );
buf ( n44424 , n38843 );
not ( n44425 , n44424 );
buf ( n44426 , n24737 );
nand ( n44427 , n44425 , n44426 );
nand ( n44428 , n44423 , n44427 );
not ( n44429 , n44428 );
not ( n44430 , n43338 );
buf ( n44431 , n44430 );
buf ( n44432 , n24939 );
not ( n44433 , n44432 );
nor ( n44434 , n44431 , n44433 );
buf ( n44435 , n24937 );
not ( n44436 , n44435 );
buf ( n44437 , n44121 );
nor ( n44438 , n44436 , n44437 );
nor ( n44439 , n44434 , n44438 );
nand ( n44440 , n44429 , n44439 );
buf ( n44441 , n24891 );
not ( n44442 , n44441 );
buf ( n44443 , n44139 );
nor ( n44444 , n44442 , n44443 );
buf ( n44445 , n24538 );
not ( n44446 , n44445 );
buf ( n44447 , n44135 );
nor ( n44448 , n44446 , n44447 );
nor ( n44449 , n44444 , n44448 );
buf ( n44450 , n14796 );
buf ( n44451 , n15509 );
not ( n44452 , n44451 );
nor ( n44453 , n44450 , n44452 );
buf ( n44454 , n44148 );
buf ( n44455 , n15557 );
not ( n44456 , n44455 );
nor ( n44457 , n44454 , n44456 );
nor ( n44458 , n44453 , n44457 );
nand ( n44459 , n44449 , n44458 );
nor ( n44460 , n44440 , n44459 );
not ( n44461 , n44460 );
buf ( n44462 , n42973 );
not ( n44463 , n44462 );
buf ( n44464 , n42996 );
nand ( n44465 , n44463 , n44464 );
buf ( n44466 , n42923 );
not ( n44467 , n44466 );
buf ( n44468 , n34926 );
nand ( n44469 , n44467 , n44468 );
nand ( n44470 , n44465 , n44469 );
buf ( n44471 , n43001 );
not ( n44472 , n44471 );
buf ( n44473 , n26497 );
nand ( n44474 , n44472 , n44473 );
not ( n44475 , n43021 );
buf ( n44476 , n44475 );
not ( n44477 , n44476 );
buf ( n44478 , n27727 );
nand ( n44479 , n44477 , n44478 );
nand ( n44480 , n44474 , n44479 );
nor ( n44481 , n44470 , n44480 );
buf ( n44482 , n27160 );
not ( n44483 , n44482 );
buf ( n44484 , n43041 );
nor ( n44485 , n44483 , n44484 );
buf ( n44486 , n20942 );
not ( n44487 , n44486 );
buf ( n44488 , n43071 );
nor ( n44489 , n44487 , n44488 );
nor ( n44490 , n44485 , n44489 );
not ( n44491 , n44490 );
buf ( n44492 , n32191 );
not ( n44493 , n44492 );
buf ( n44494 , n43079 );
not ( n44495 , n44494 );
not ( n44496 , n44495 );
or ( n44497 , n44493 , n44496 );
buf ( n44498 , n43095 );
buf ( n44499 , n32404 );
not ( n44500 , n44499 );
nor ( n44501 , n44498 , n44500 );
not ( n44502 , n44501 );
nand ( n44503 , n44497 , n44502 );
nor ( n44504 , n44491 , n44503 );
buf ( n44505 , n37914 );
not ( n44506 , n44505 );
buf ( n44507 , n43222 );
nor ( n44508 , n44506 , n44507 );
buf ( n44509 , n24723 );
not ( n44510 , n44509 );
buf ( n44511 , n43237 );
nor ( n44512 , n44510 , n44511 );
nor ( n44513 , n44508 , n44512 );
buf ( n44514 , n43194 );
buf ( n44515 , n34667 );
not ( n44516 , n44515 );
nor ( n44517 , n44514 , n44516 );
buf ( n44518 , n32957 );
not ( n44519 , n44518 );
buf ( n44520 , n43202 );
nor ( n44521 , n44519 , n44520 );
nor ( n44522 , n44517 , n44521 );
buf ( n44523 , n43135 );
not ( n44524 , n44523 );
buf ( n44525 , n34720 );
nand ( n44526 , n44524 , n44525 );
buf ( n44527 , n20678 );
not ( n44528 , n44527 );
buf ( n44529 , n43161 );
nor ( n44530 , n44528 , n44529 );
buf ( n44531 , n14542 );
not ( n44532 , n44531 );
buf ( n44533 , n21684 );
and ( n44534 , n44532 , n44533 );
or ( n44535 , n44530 , n44534 );
or ( n44536 , n44532 , n44533 );
nand ( n44537 , n44535 , n44536 );
buf ( n44538 , n43172 );
not ( n44539 , n44538 );
buf ( n44540 , n36637 );
nand ( n44541 , n44539 , n44540 );
nand ( n44542 , n44526 , n44537 , n44541 );
not ( n44543 , n44538 );
nor ( n44544 , n44543 , n44540 );
nand ( n44545 , n44526 , n44544 );
not ( n44546 , n44525 );
nand ( n44547 , n44546 , n44523 );
nand ( n44548 , n44542 , n44545 , n44547 );
nand ( n44549 , n44513 , n44522 , n44548 );
not ( n44550 , n44518 );
nand ( n44551 , n44550 , n44520 );
or ( n44552 , n44517 , n44551 );
nand ( n44553 , n44514 , n44516 );
nand ( n44554 , n44552 , n44553 );
nand ( n44555 , n44513 , n44554 );
not ( n44556 , n44508 );
not ( n44557 , n44511 );
nor ( n44558 , n44557 , n44509 );
and ( n44559 , n44556 , n44558 );
not ( n44560 , n44507 );
nor ( n44561 , n44560 , n44505 );
nor ( n44562 , n44559 , n44561 );
nand ( n44563 , n44549 , n44555 , n44562 );
and ( n44564 , n44481 , n44504 , n44563 );
not ( n44565 , n44481 );
not ( n44566 , n44490 );
not ( n44567 , n44492 );
nand ( n44568 , n44567 , n44494 );
or ( n44569 , n44501 , n44568 );
nand ( n44570 , n44498 , n44500 );
nand ( n44571 , n44569 , n44570 );
not ( n44572 , n44571 );
or ( n44573 , n44566 , n44572 );
not ( n44574 , n44485 );
not ( n44575 , n44488 );
nor ( n44576 , n44575 , n44486 );
and ( n44577 , n44574 , n44576 );
not ( n44578 , n44484 );
nor ( n44579 , n44578 , n44482 );
nor ( n44580 , n44577 , n44579 );
nand ( n44581 , n44573 , n44580 );
not ( n44582 , n44581 );
or ( n44583 , n44565 , n44582 );
not ( n44584 , n44470 );
not ( n44585 , n44474 );
not ( n44586 , n44478 );
nand ( n44587 , n44586 , n44476 );
or ( n44588 , n44585 , n44587 );
not ( n44589 , n44473 );
nand ( n44590 , n44589 , n44471 );
nand ( n44591 , n44588 , n44590 );
and ( n44592 , n44584 , n44591 );
not ( n44593 , n44465 );
not ( n44594 , n44468 );
nand ( n44595 , n44594 , n44466 );
or ( n44596 , n44593 , n44595 );
not ( n44597 , n44464 );
nand ( n44598 , n44597 , n44462 );
nand ( n44599 , n44596 , n44598 );
nor ( n44600 , n44592 , n44599 );
nand ( n44601 , n44583 , n44600 );
nor ( n44602 , n44564 , n44601 );
not ( n44603 , n43473 );
buf ( n44604 , n44603 );
buf ( n44605 , n32693 );
not ( n44606 , n44605 );
nor ( n44607 , n44604 , n44606 );
buf ( n44608 , n43499 );
buf ( n44609 , n33042 );
not ( n44610 , n44609 );
nor ( n44611 , n44608 , n44610 );
nor ( n44612 , n44607 , n44611 );
not ( n44613 , n43532 );
buf ( n44614 , n44613 );
buf ( n44615 , n20787 );
not ( n44616 , n44615 );
nor ( n44617 , n44614 , n44616 );
buf ( n44618 , n43543 );
buf ( n44619 , n31330 );
not ( n44620 , n44619 );
nor ( n44621 , n44618 , n44620 );
nor ( n44622 , n44617 , n44621 );
nand ( n44623 , n44612 , n44622 );
not ( n44624 , n44623 );
buf ( n44625 , n43562 );
buf ( n44626 , n32326 );
not ( n44627 , n44626 );
nor ( n44628 , n44625 , n44627 );
not ( n44629 , n44342 );
buf ( n44630 , n44629 );
buf ( n44631 , n44338 );
not ( n44632 , n44631 );
nor ( n44633 , n44630 , n44632 );
nor ( n44634 , n44628 , n44633 );
not ( n44635 , n44634 );
not ( n44636 , n31173 );
buf ( n44637 , n44636 );
not ( n44638 , n44637 );
buf ( n44639 , n43598 );
not ( n44640 , n44639 );
not ( n44641 , n44640 );
or ( n44642 , n44638 , n44641 );
buf ( n44643 , n44358 );
buf ( n44644 , n23446 );
not ( n44645 , n44644 );
nor ( n44646 , n44643 , n44645 );
not ( n44647 , n44646 );
nand ( n44648 , n44642 , n44647 );
nor ( n44649 , n44635 , n44648 );
nand ( n44650 , n44624 , n44649 );
nor ( n44651 , n44461 , n44602 , n44650 );
nand ( n44652 , n44643 , n44645 );
not ( n44653 , n44637 );
nand ( n44654 , n44653 , n44639 );
and ( n44655 , n44652 , n44654 );
nor ( n44656 , n44655 , n44646 );
and ( n44657 , n44634 , n44656 );
nand ( n44658 , n44630 , n44632 );
or ( n44659 , n44628 , n44658 );
nand ( n44660 , n44625 , n44627 );
nand ( n44661 , n44659 , n44660 );
nor ( n44662 , n44657 , n44661 );
or ( n44663 , n44662 , n44623 );
nand ( n44664 , n44618 , n44620 );
or ( n44665 , n44617 , n44664 );
nand ( n44666 , n44614 , n44616 );
nand ( n44667 , n44665 , n44666 );
and ( n44668 , n44667 , n44612 );
nand ( n44669 , n44608 , n44610 );
or ( n44670 , n44607 , n44669 );
nand ( n44671 , n44604 , n44606 );
nand ( n44672 , n44670 , n44671 );
nor ( n44673 , n44668 , n44672 );
nand ( n44674 , n44663 , n44673 );
not ( n44675 , n44674 );
not ( n44676 , n44460 );
or ( n44677 , n44675 , n44676 );
not ( n44678 , n44440 );
nand ( n44679 , n44450 , n44452 );
nand ( n44680 , n44454 , n44456 );
and ( n44681 , n44679 , n44680 );
nor ( n44682 , n44681 , n44453 );
not ( n44683 , n44682 );
not ( n44684 , n44449 );
or ( n44685 , n44683 , n44684 );
not ( n44686 , n44444 );
not ( n44687 , n44447 );
nor ( n44688 , n44687 , n44445 );
and ( n44689 , n44686 , n44688 );
not ( n44690 , n44443 );
nor ( n44691 , n44690 , n44441 );
nor ( n44692 , n44689 , n44691 );
nand ( n44693 , n44685 , n44692 );
and ( n44694 , n44678 , n44693 );
not ( n44695 , n44434 );
not ( n44696 , n44437 );
nor ( n44697 , n44696 , n44435 );
and ( n44698 , n44695 , n44697 );
not ( n44699 , n44431 );
nor ( n44700 , n44699 , n44432 );
nor ( n44701 , n44698 , n44700 );
or ( n44702 , n44428 , n44701 );
nor ( n44703 , n44421 , n44418 );
and ( n44704 , n44427 , n44703 );
not ( n44705 , n44424 );
nor ( n44706 , n44705 , n44426 );
nor ( n44707 , n44704 , n44706 );
nand ( n44708 , n44702 , n44707 );
nor ( n44709 , n44694 , n44708 );
nand ( n44710 , n44677 , n44709 );
nor ( n44711 , n44651 , n44710 );
buf ( n44712 , n44711 );
or ( n44713 , n44712 , n43712 );
nand ( n44714 , n44417 , n44713 );
or ( n44715 , n44714 , n26359 );
nand ( n44716 , n44714 , n17543 );
nand ( n44717 , n14894 , n14847 );
nand ( n44718 , n44715 , n44716 , n44717 );
and ( n44719 , n44718 , n14838 );
nand ( n44720 , n44100 , n14886 , n44103 , n14905 );
not ( n44721 , n22899 );
not ( n44722 , n23151 );
not ( n44723 , n14907 );
or ( n44724 , n44722 , n44723 );
nand ( n44725 , n44724 , n22898 );
not ( n44726 , n44725 );
or ( n44727 , n44721 , n44726 );
nand ( n44728 , n44727 , n14847 );
nand ( n44729 , n44720 , n44728 );
nor ( n44730 , n44719 , n44729 );
nand ( n44731 , n44105 , n44730 );
buf ( n44732 , n44731 );
buf ( n44733 , n44732 );
buf ( n44734 , n275554 );
not ( n44735 , n275925 );
buf ( n44736 , n44735 );
buf ( n44737 , n44736 );
buf ( n44738 , n275554 );
or ( n44739 , n27843 , n19216 );
buf ( n44740 , n35150 );
nand ( n44741 , n28049 , n44740 );
nand ( n44742 , n28120 , n19360 );
nand ( n44743 , n28140 , n29075 );
not ( n44744 , n39767 );
not ( n44745 , n19317 );
and ( n44746 , n44744 , n44745 );
and ( n44747 , n33162 , n27885 );
nor ( n44748 , n44746 , n44747 );
nand ( n44749 , n19387 , n18638 );
and ( n44750 , n44743 , n44748 , n44749 );
and ( n44751 , n44741 , n44742 , n44750 );
nand ( n44752 , n44739 , n44751 );
buf ( n44753 , n44752 );
buf ( n44754 , n44753 );
buf ( n44755 , n275554 );
not ( n44756 , n275929 );
buf ( n44757 , n44756 );
buf ( n44758 , n44757 );
or ( n44759 , n35814 , n32074 );
not ( n44760 , n38353 );
not ( n44761 , n35832 );
and ( n44762 , n44760 , n44761 );
and ( n44763 , n35862 , n20353 );
nor ( n44764 , n44762 , n44763 );
and ( n44765 , n35826 , n20515 );
not ( n44766 , n41707 );
nand ( n44767 , n35847 , n31095 );
nand ( n44768 , n19644 , n35837 );
nand ( n44769 , n44766 , n44767 , n44768 );
nor ( n44770 , n44765 , n44769 );
and ( n44771 , n44764 , n44770 );
nand ( n44772 , n44759 , n44771 );
buf ( n44773 , n44772 );
buf ( n44774 , n44773 );
buf ( n44775 , n275554 );
buf ( n44776 , n275554 );
nand ( n44777 , n25064 , n18071 );
buf ( n44778 , n25205 );
buf ( n44779 , n25212 );
nand ( n44780 , n44778 , n44779 );
buf ( n44781 , n44780 );
buf ( n44782 , n44781 );
not ( n44783 , n44782 );
buf ( n44784 , n25180 );
not ( n44785 , n44784 );
buf ( n44786 , n25218 );
nand ( n44787 , n44785 , n44786 );
buf ( n44788 , n44787 );
buf ( n44789 , n44788 );
not ( n44790 , n44789 );
or ( n44791 , n44783 , n44790 );
buf ( n44792 , n44788 );
buf ( n44793 , n44781 );
or ( n44794 , n44792 , n44793 );
nand ( n44795 , n44791 , n44794 );
buf ( n44796 , n44795 );
buf ( n44797 , n44796 );
not ( n44798 , n44797 );
nor ( n44799 , n44798 , n25389 );
nand ( n44800 , n25397 , n275689 );
buf ( n44801 , n25524 );
buf ( n44802 , n25531 );
nand ( n44803 , n44801 , n44802 );
buf ( n44804 , n44803 );
buf ( n44805 , n44804 );
not ( n44806 , n44805 );
buf ( n44807 , n25501 );
not ( n44808 , n44807 );
buf ( n44809 , n25537 );
nand ( n44810 , n44808 , n44809 );
buf ( n44811 , n44810 );
buf ( n44812 , n44811 );
not ( n44813 , n44812 );
or ( n44814 , n44806 , n44813 );
buf ( n44815 , n44811 );
buf ( n44816 , n44804 );
or ( n44817 , n44815 , n44816 );
nand ( n44818 , n44814 , n44817 );
buf ( n44819 , n44818 );
buf ( n44820 , n44819 );
and ( n44821 , n25402 , n44820 );
nor ( n44822 , n44821 , n39786 );
buf ( n44823 , n25840 );
buf ( n44824 , n25847 );
nand ( n44825 , n44823 , n44824 );
buf ( n44826 , n44825 );
buf ( n44827 , n44826 );
not ( n44828 , n44827 );
buf ( n44829 , n25817 );
not ( n44830 , n44829 );
buf ( n44831 , n25853 );
nand ( n44832 , n44830 , n44831 );
buf ( n44833 , n44832 );
buf ( n44834 , n44833 );
not ( n44835 , n44834 );
or ( n44836 , n44828 , n44835 );
buf ( n44837 , n44833 );
buf ( n44838 , n44826 );
or ( n44839 , n44837 , n44838 );
nand ( n44840 , n44836 , n44839 );
buf ( n44841 , n44840 );
buf ( n44842 , n44841 );
nand ( n44843 , n28761 , n44842 );
nand ( n44844 , n44800 , n44822 , n44843 );
nor ( n44845 , n44799 , n44844 );
buf ( n44846 , n26126 );
not ( n44847 , n44846 );
buf ( n44848 , n26163 );
nand ( n44849 , n44847 , n44848 );
buf ( n44850 , n44849 );
buf ( n44851 , n44850 );
not ( n44852 , n44851 );
buf ( n44853 , n26150 );
buf ( n44854 , n26157 );
nand ( n44855 , n44853 , n44854 );
buf ( n44856 , n44855 );
buf ( n44857 , n44856 );
not ( n44858 , n44857 );
or ( n44859 , n44852 , n44858 );
buf ( n44860 , n44850 );
buf ( n44861 , n44856 );
or ( n44862 , n44860 , n44861 );
nand ( n44863 , n44859 , n44862 );
buf ( n44864 , n44863 );
buf ( n44865 , n44864 );
nand ( n44866 , n26027 , n44865 );
nand ( n44867 , n44777 , n44845 , n44866 );
buf ( n44868 , n44867 );
buf ( n44869 , n44868 );
or ( n44870 , n32914 , n21697 );
nand ( n44871 , n34674 , n13818 );
nand ( n44872 , n44870 , n44871 );
buf ( n44873 , n44872 );
buf ( n44874 , n44873 );
not ( n44875 , n33256 );
or ( n44876 , n44875 , n21774 );
nand ( n44877 , n21774 , n9724 );
nand ( n44878 , n44876 , n44877 );
buf ( n44879 , n44878 );
buf ( n44880 , n44879 );
not ( n44881 , n10737 );
not ( n44882 , n9157 );
or ( n44883 , n44881 , n44882 );
not ( n44884 , n10718 );
or ( n44885 , n9157 , n44884 );
nand ( n44886 , n44883 , n44885 );
buf ( n44887 , n44886 );
buf ( n44888 , n44887 );
not ( n44889 , n37871 );
not ( n44890 , n23789 );
and ( n44891 , n44889 , n44890 );
nand ( n44892 , n37891 , n20889 );
nand ( n44893 , n37933 , n24711 );
and ( n44894 , n37909 , n17409 );
and ( n44895 , n20940 , n37915 );
nor ( n44896 , n44894 , n44895 );
nand ( n44897 , n44892 , n44893 , n44896 );
nor ( n44898 , n44891 , n44897 );
or ( n44899 , n44898 , n20950 );
nand ( n44900 , n20950 , n13578 );
nand ( n44901 , n44899 , n44900 );
buf ( n44902 , n44901 );
buf ( n44903 , n44902 );
not ( n44904 , n275550 );
buf ( n44905 , n44904 );
buf ( n44906 , n44905 );
and ( n44907 , n20711 , n29057 );
not ( n44908 , n20711 );
not ( n44909 , n14228 );
not ( n44910 , n44909 );
not ( n44911 , n34859 );
nor ( n44912 , n34861 , n44911 );
not ( n44913 , n44912 );
or ( n44914 , n44910 , n44913 );
or ( n44915 , n44912 , n44909 );
nand ( n44916 , n44914 , n44915 );
buf ( n44917 , n44916 );
and ( n44918 , n44908 , n44917 );
nor ( n44919 , n44907 , n44918 );
or ( n44920 , n44919 , n26364 );
nand ( n44921 , n16881 , n16886 );
not ( n44922 , n44921 );
nand ( n44923 , n16668 , n34871 );
nor ( n44924 , n44923 , n26445 );
not ( n44925 , n44924 );
not ( n44926 , n20875 );
or ( n44927 , n44925 , n44926 );
not ( n44928 , n26451 );
not ( n44929 , n44923 );
and ( n44930 , n44928 , n44929 );
or ( n44931 , n34880 , n16618 );
nand ( n44932 , n44931 , n34872 );
nor ( n44933 , n44930 , n44932 );
nand ( n44934 , n44927 , n44933 );
not ( n44935 , n44934 );
or ( n44936 , n44922 , n44935 );
or ( n44937 , n44934 , n44921 );
nand ( n44938 , n44936 , n44937 );
buf ( n44939 , n44938 );
nand ( n44940 , n44939 , n26370 );
not ( n44941 , n17133 );
nand ( n44942 , n44941 , n17356 );
not ( n44943 , n44942 );
nand ( n44944 , n17121 , n34889 );
nor ( n44945 , n44944 , n17229 );
not ( n44946 , n44945 );
not ( n44947 , n20913 );
or ( n44948 , n44946 , n44947 );
not ( n44949 , n26473 );
not ( n44950 , n44944 );
and ( n44951 , n44949 , n44950 );
not ( n44952 , n34889 );
not ( n44953 , n17352 );
or ( n44954 , n44952 , n44953 );
nand ( n44955 , n44954 , n17354 );
nor ( n44956 , n44951 , n44955 );
nand ( n44957 , n44948 , n44956 );
not ( n44958 , n44957 );
or ( n44959 , n44943 , n44958 );
or ( n44960 , n44957 , n44942 );
nand ( n44961 , n44959 , n44960 );
buf ( n44962 , n44961 );
nand ( n44963 , n44962 , n26374 );
and ( n44964 , n17519 , n17520 );
not ( n44965 , n17519 );
and ( n44966 , n44965 , n13491 );
nor ( n44967 , n44964 , n44966 );
nand ( n44968 , n32176 , n44967 );
not ( n44969 , n17451 );
not ( n44970 , n34916 );
and ( n44971 , n44970 , n26486 , n17458 );
not ( n44972 , n44971 );
or ( n44973 , n44969 , n44972 );
or ( n44974 , n44971 , n17451 );
nand ( n44975 , n44973 , n44974 );
buf ( n44976 , n44975 );
nand ( n44977 , n44976 , n26393 );
buf ( n44978 , n42996 );
nand ( n44979 , n26395 , n44978 );
not ( n44980 , n31470 );
and ( n44981 , n44977 , n44979 , n44980 );
and ( n44982 , n44940 , n44963 , n44968 , n44981 );
nand ( n44983 , n44920 , n44982 );
buf ( n44984 , n44983 );
buf ( n44985 , n44984 );
and ( n44986 , n31719 , n277618 );
not ( n44987 , n31719 );
and ( n44988 , n44987 , n35052 );
or ( n44989 , n44986 , n44988 );
buf ( n44990 , n44989 );
buf ( n44991 , n44990 );
buf ( n44992 , n275554 );
buf ( n44993 , n275554 );
not ( n44994 , n11238 );
or ( n44995 , n44994 , n9158 );
not ( n44996 , n11202 );
or ( n44997 , n44996 , n9157 );
nand ( n44998 , n44995 , n44997 );
buf ( n44999 , n44998 );
buf ( n45000 , n44999 );
nand ( n45001 , n42796 , n31422 );
nand ( n45002 , n42819 , n28330 );
nand ( n45003 , n42829 , n31449 );
and ( n45004 , n36530 , n12371 );
not ( n45005 , n277715 );
not ( n45006 , n28357 );
or ( n45007 , n45005 , n45006 );
or ( n45008 , n32061 , n277703 );
nand ( n45009 , n45007 , n45008 );
nor ( n45010 , n45004 , n45009 );
nand ( n45011 , n31460 , n12304 );
and ( n45012 , n45003 , n45010 , n45011 );
nand ( n45013 , n45001 , n45002 , n45012 );
buf ( n45014 , n45013 );
buf ( n45015 , n45014 );
not ( n45016 , n275929 );
buf ( n45017 , n45016 );
buf ( n45018 , n45017 );
buf ( n45019 , n275554 );
buf ( n45020 , n275554 );
buf ( n45021 , n275554 );
or ( n45022 , n38388 , n21030 );
nand ( n45023 , n21030 , n18963 );
nand ( n45024 , n45022 , n45023 );
buf ( n45025 , n45024 );
buf ( n45026 , n45025 );
buf ( n45027 , n275554 );
not ( n45028 , n275550 );
buf ( n45029 , n45028 );
buf ( n45030 , n45029 );
and ( n45031 , n14830 , n13099 );
not ( n45032 , n14830 );
and ( n45033 , n45032 , n16692 );
or ( n45034 , n45031 , n45033 );
buf ( n45035 , n45034 );
buf ( n45036 , n45035 );
not ( n45037 , n275929 );
buf ( n45038 , n45037 );
buf ( n45039 , n45038 );
buf ( n45040 , n275554 );
and ( n45041 , n31142 , n23788 );
nand ( n45042 , n31152 , n20889 );
nand ( n45043 , n31161 , n20926 );
and ( n45044 , n31169 , n17409 );
and ( n45045 , n20940 , n31174 );
nor ( n45046 , n45044 , n45045 );
nand ( n45047 , n45042 , n45043 , n45046 );
nor ( n45048 , n45041 , n45047 );
or ( n45049 , n45048 , n20950 );
nand ( n45050 , n20950 , n13783 );
nand ( n45051 , n45049 , n45050 );
buf ( n45052 , n45051 );
buf ( n45053 , n45052 );
buf ( n45054 , n275554 );
buf ( n45055 , n275554 );
not ( n45056 , n24767 );
or ( n45057 , n45056 , n29044 );
nand ( n45058 , n29046 , n9783 );
nand ( n45059 , n45057 , n45058 );
buf ( n45060 , n45059 );
buf ( n45061 , n45060 );
or ( n45062 , n40684 , n23708 );
nand ( n45063 , n27641 , n11616 );
nand ( n45064 , n45062 , n45063 );
buf ( n45065 , n45064 );
buf ( n45066 , n45065 );
buf ( n45067 , n275554 );
buf ( n45068 , n275554 );
not ( n45069 , n275925 );
buf ( n45070 , n45069 );
buf ( n45071 , n45070 );
buf ( n45072 , n275554 );
not ( n45073 , n275929 );
buf ( n45074 , n45073 );
buf ( n45075 , n45074 );
not ( n45076 , n34623 );
or ( n45077 , n45076 , n29046 );
nand ( n45078 , n29044 , n9488 );
nand ( n45079 , n45077 , n45078 );
buf ( n45080 , n45079 );
buf ( n45081 , n45080 );
buf ( n45082 , n275554 );
buf ( n45083 , n275554 );
not ( n45084 , n275826 );
nand ( n45085 , n45084 , n275844 );
not ( n45086 , n45085 );
or ( n45087 , n40826 , n275833 );
nand ( n45088 , n45087 , n275842 );
not ( n45089 , n45088 );
or ( n45090 , n45086 , n45089 );
or ( n45091 , n45088 , n45085 );
nand ( n45092 , n45090 , n45091 );
buf ( n45093 , n45092 );
buf ( n45094 , n45093 );
buf ( n45095 , n275554 );
buf ( n45096 , n275554 );
buf ( n45097 , n275554 );
not ( n45098 , n38025 );
buf ( n45099 , n45098 );
buf ( n45100 , n45099 );
not ( n45101 , n278010 );
not ( n45102 , n27179 );
or ( n45103 , n45101 , n45102 );
not ( n45104 , n37091 );
or ( n45105 , n45104 , n27179 );
nand ( n45106 , n45103 , n45105 );
buf ( n45107 , n45106 );
buf ( n45108 , n45107 );
buf ( n45109 , n275554 );
buf ( n45110 , n275554 );
not ( n45111 , n275925 );
buf ( n45112 , n45111 );
buf ( n45113 , n45112 );
not ( n45114 , n275929 );
buf ( n45115 , n45114 );
buf ( n45116 , n45115 );
and ( n45117 , n20950 , n14745 );
not ( n45118 , n20950 );
and ( n45119 , n45118 , n38856 );
or ( n45120 , n45117 , n45119 );
buf ( n45121 , n45120 );
buf ( n45122 , n45121 );
buf ( n45123 , n275554 );
not ( n45124 , n275550 );
buf ( n45125 , n45124 );
buf ( n45126 , n45125 );
or ( n45127 , n37798 , n22193 );
or ( n45128 , n29380 , n11259 );
nand ( n45129 , n45127 , n45128 );
buf ( n45130 , n45129 );
buf ( n45131 , n45130 );
buf ( n45132 , n275554 );
buf ( n45133 , n275554 );
not ( n45134 , n275550 );
buf ( n45135 , n45134 );
buf ( n45136 , n45135 );
and ( n45137 , n14830 , n13339 );
not ( n45138 , n14830 );
and ( n45139 , n45138 , n38842 );
or ( n45140 , n45137 , n45139 );
buf ( n45141 , n45140 );
buf ( n45142 , n45141 );
not ( n45143 , n21769 );
buf ( n45144 , n45143 );
buf ( n45145 , n45144 );
not ( n45146 , n275929 );
buf ( n45147 , n45146 );
buf ( n45148 , n45147 );
or ( n45149 , n30748 , n31719 );
or ( n45150 , n35071 , n11477 );
nand ( n45151 , n45149 , n45150 );
buf ( n45152 , n45151 );
buf ( n45153 , n45152 );
not ( n45154 , n20142 );
not ( n45155 , n275557 );
or ( n45156 , n45154 , n45155 );
nand ( n45157 , n22335 , n25164 );
nand ( n45158 , n45156 , n45157 );
buf ( n45159 , n45158 );
buf ( n45160 , n45159 );
not ( n45161 , n31303 );
or ( n45162 , n45161 , n29044 );
nand ( n45163 , n29046 , n9702 );
nand ( n45164 , n45162 , n45163 );
buf ( n45165 , n45164 );
buf ( n45166 , n45165 );
not ( n45167 , n34302 );
not ( n45168 , n42653 );
or ( n45169 , n45167 , n45168 );
and ( n45170 , n42667 , n35900 );
nand ( n45171 , n42676 , n34307 );
nand ( n45172 , n28451 , n277839 );
nand ( n45173 , n32755 , n11826 );
and ( n45174 , n34311 , n12248 );
and ( n45175 , n34313 , n9333 );
nor ( n45176 , n45174 , n45175 );
and ( n45177 , n45173 , n45176 );
nand ( n45178 , n45171 , n45172 , n45177 );
nor ( n45179 , n45170 , n45178 );
nand ( n45180 , n45169 , n45179 );
buf ( n45181 , n45180 );
buf ( n45182 , n45181 );
or ( n45183 , n34869 , n20743 );
nand ( n45184 , n34887 , n16970 );
nand ( n45185 , n34906 , n17405 );
nand ( n45186 , n32339 , n34922 );
nand ( n45187 , n17502 , n34928 );
nand ( n45188 , n17562 , n13522 );
nand ( n45189 , n17545 , n34912 );
and ( n45190 , n45186 , n45187 , n45188 , n45189 );
and ( n45191 , n45184 , n45185 , n45190 );
nand ( n45192 , n45183 , n45191 );
buf ( n45193 , n45192 );
buf ( n45194 , n45193 );
or ( n45195 , n34634 , n14909 );
not ( n45196 , n16970 );
not ( n45197 , n34648 );
or ( n45198 , n45196 , n45197 );
not ( n45199 , n39651 );
not ( n45200 , n17545 );
or ( n45201 , n45199 , n45200 );
not ( n45202 , n34664 );
or ( n45203 , n17410 , n45202 );
nand ( n45204 , n45201 , n45203 );
not ( n45205 , n34668 );
nor ( n45206 , n45205 , n17501 );
nor ( n45207 , n45204 , n45206 );
nand ( n45208 , n45198 , n45207 );
not ( n45209 , n17405 );
not ( n45210 , n34656 );
or ( n45211 , n45209 , n45210 );
nand ( n45212 , n17562 , n13670 );
nand ( n45213 , n45211 , n45212 );
nor ( n45214 , n45208 , n45213 );
nand ( n45215 , n45195 , n45214 );
buf ( n45216 , n45215 );
buf ( n45217 , n45216 );
buf ( n45218 , n275554 );
buf ( n45219 , n275554 );
nand ( n45220 , n25064 , n18131 );
xor ( n45221 , n25188 , n25189 );
xor ( n45222 , n45221 , n25191 );
buf ( n45223 , n45222 );
buf ( n45224 , n45223 );
and ( n45225 , n34544 , n45224 );
not ( n45226 , n275725 );
not ( n45227 , n25396 );
or ( n45228 , n45226 , n45227 );
xor ( n45229 , n25507 , n25508 );
xor ( n45230 , n45229 , n25510 );
buf ( n45231 , n45230 );
buf ( n45232 , n45231 );
and ( n45233 , n25402 , n45232 );
xor ( n45234 , n25823 , n25824 );
xor ( n45235 , n45234 , n25826 );
buf ( n45236 , n45235 );
buf ( n45237 , n45236 );
not ( n45238 , n45237 );
not ( n45239 , n28761 );
or ( n45240 , n45238 , n45239 );
nand ( n45241 , n275557 , n19088 );
nand ( n45242 , n45240 , n45241 );
nor ( n45243 , n45233 , n45242 );
nand ( n45244 , n45228 , n45243 );
nor ( n45245 , n45225 , n45244 );
xor ( n45246 , n26133 , n26134 );
xor ( n45247 , n45246 , n26136 );
buf ( n45248 , n45247 );
buf ( n45249 , n45248 );
nand ( n45250 , n26027 , n45249 );
nand ( n45251 , n45220 , n45245 , n45250 );
buf ( n45252 , n45251 );
buf ( n45253 , n45252 );
buf ( n45254 , n275554 );
not ( n45255 , n275550 );
buf ( n45256 , n45255 );
buf ( n45257 , n45256 );
not ( n45258 , n31041 );
or ( n45259 , n45258 , n21770 );
nand ( n45260 , n21774 , n9679 );
nand ( n45261 , n45259 , n45260 );
buf ( n45262 , n45261 );
buf ( n45263 , n45262 );
buf ( n45264 , n275554 );
not ( n45265 , n275550 );
buf ( n45266 , n45265 );
buf ( n45267 , n45266 );
not ( n45268 , n275929 );
buf ( n45269 , n45268 );
buf ( n45270 , n45269 );
buf ( n45271 , n275554 );
buf ( n45272 , n275554 );
not ( n45273 , n275925 );
buf ( n45274 , n45273 );
buf ( n45275 , n45274 );
not ( n45276 , n275925 );
buf ( n45277 , n45276 );
buf ( n45278 , n45277 );
buf ( n45279 , n275554 );
buf ( n45280 , n275554 );
not ( n45281 , n22052 );
not ( n45282 , n27505 );
nor ( n45283 , n27569 , n27571 );
not ( n45284 , n45283 );
or ( n45285 , n45282 , n45284 );
or ( n45286 , n45283 , n27505 );
nand ( n45287 , n45285 , n45286 );
buf ( n45288 , n45287 );
not ( n45289 , n45288 );
or ( n45290 , n45281 , n45289 );
nand ( n45291 , n22084 , n22088 );
not ( n45292 , n45291 );
not ( n45293 , n27578 );
not ( n45294 , n22128 );
or ( n45295 , n45293 , n45294 );
nand ( n45296 , n45295 , n27579 );
not ( n45297 , n45296 );
or ( n45298 , n45292 , n45297 );
or ( n45299 , n45296 , n45291 );
nand ( n45300 , n45298 , n45299 );
buf ( n45301 , n45300 );
nand ( n45302 , n45301 , n22057 );
nand ( n45303 , n45290 , n45302 );
not ( n45304 , n23603 );
buf ( n45305 , n21940 );
buf ( n45306 , n21839 );
nand ( n45307 , n45305 , n45306 );
buf ( n45308 , n45307 );
buf ( n45309 , n45308 );
not ( n45310 , n45309 );
buf ( n45311 , n21945 );
not ( n45312 , n45311 );
buf ( n45313 , n21938 );
not ( n45314 , n45313 );
or ( n45315 , n45312 , n45314 );
buf ( n45316 , n27535 );
nand ( n45317 , n45315 , n45316 );
buf ( n45318 , n45317 );
buf ( n45319 , n45318 );
not ( n45320 , n45319 );
or ( n45321 , n45310 , n45320 );
buf ( n45322 , n45318 );
buf ( n45323 , n45308 );
or ( n45324 , n45322 , n45323 );
nand ( n45325 , n45321 , n45324 );
buf ( n45326 , n45325 );
buf ( n45327 , n45326 );
not ( n45328 , n45327 );
or ( n45329 , n45304 , n45328 );
not ( n45330 , n32722 );
not ( n45331 , n12261 );
and ( n45332 , n45330 , n45331 );
and ( n45333 , n23679 , n11848 );
nor ( n45334 , n45332 , n45333 );
nand ( n45335 , n45329 , n45334 );
nor ( n45336 , n45303 , n45335 );
or ( n45337 , n45336 , n22193 );
or ( n45338 , n22192 , n10910 );
nand ( n45339 , n45337 , n45338 );
buf ( n45340 , n45339 );
buf ( n45341 , n45340 );
or ( n45342 , n26438 , n26364 );
nand ( n45343 , n26462 , n26370 );
nand ( n45344 , n26483 , n26374 );
nand ( n45345 , n32176 , n41265 );
nand ( n45346 , n26493 , n26393 );
nand ( n45347 , n26395 , n26498 );
nor ( n45348 , n14830 , n41263 );
not ( n45349 , n45348 );
and ( n45350 , n45346 , n45347 , n45349 );
and ( n45351 , n45343 , n45344 , n45345 , n45350 );
nand ( n45352 , n45342 , n45351 );
buf ( n45353 , n45352 );
buf ( n45354 , n45353 );
buf ( n45355 , n275554 );
not ( n45356 , n275550 );
buf ( n45357 , n45356 );
buf ( n45358 , n45357 );
buf ( n45359 , n275554 );
not ( n45360 , n275929 );
buf ( n45361 , n45360 );
buf ( n45362 , n45361 );
not ( n45363 , n275929 );
buf ( n45364 , n45363 );
buf ( n45365 , n45364 );
not ( n45366 , n275925 );
buf ( n45367 , n45366 );
buf ( n45368 , n45367 );
or ( n45369 , n45048 , n21696 );
nand ( n45370 , n27647 , n13774 );
nand ( n45371 , n45369 , n45370 );
buf ( n45372 , n45371 );
buf ( n45373 , n45372 );
not ( n45374 , n275925 );
buf ( n45375 , n45374 );
buf ( n45376 , n45375 );
buf ( n45377 , n275554 );
or ( n45378 , n35412 , n29866 );
nand ( n45379 , n35431 , n20353 );
nand ( n45380 , n35453 , n30132 );
not ( n45381 , n34104 );
not ( n45382 , n40840 );
not ( n45383 , n45382 );
and ( n45384 , n45381 , n45383 );
nand ( n45385 , n35467 , n20560 );
nand ( n45386 , n29494 , n30019 );
nand ( n45387 , n30179 , n18487 );
nand ( n45388 , n45385 , n45386 , n45387 );
nor ( n45389 , n45384 , n45388 );
and ( n45390 , n45379 , n45380 , n45389 );
nand ( n45391 , n45378 , n45390 );
buf ( n45392 , n45391 );
buf ( n45393 , n45392 );
not ( n45394 , n275550 );
buf ( n45395 , n45394 );
buf ( n45396 , n45395 );
not ( n45397 , n275550 );
buf ( n45398 , n45397 );
buf ( n45399 , n45398 );
not ( n45400 , n16550 );
or ( n45401 , n45400 , n14830 );
nand ( n45402 , n31508 , n23807 );
nand ( n45403 , n45401 , n45402 );
buf ( n45404 , n45403 );
buf ( n45405 , n45404 );
not ( n45406 , n27265 );
not ( n45407 , n35900 );
or ( n45408 , n45406 , n45407 );
nand ( n45409 , n27488 , n28408 );
nand ( n45410 , n27518 , n34307 );
nand ( n45411 , n28451 , n10624 );
nand ( n45412 , n29171 , n40516 );
nand ( n45413 , n34311 , n12290 );
nand ( n45414 , n20649 , n9312 );
and ( n45415 , n45412 , n45413 , n45414 );
and ( n45416 , n45410 , n45411 , n45415 );
nand ( n45417 , n45408 , n45409 , n45416 );
buf ( n45418 , n45417 );
buf ( n45419 , n45418 );
buf ( n45420 , n275554 );
buf ( n45421 , n275554 );
not ( n45422 , n275925 );
buf ( n45423 , n45422 );
buf ( n45424 , n45423 );
not ( n45425 , n275550 );
buf ( n45426 , n45425 );
buf ( n45427 , n45426 );
not ( n45428 , n275929 );
buf ( n45429 , n45428 );
buf ( n45430 , n45429 );
not ( n45431 , n275925 );
buf ( n45432 , n45431 );
buf ( n45433 , n45432 );
or ( n45434 , n20985 , n19216 );
nand ( n45435 , n20998 , n19354 );
not ( n45436 , n19291 );
not ( n45437 , n21018 );
not ( n45438 , n45437 );
and ( n45439 , n45436 , n45438 );
and ( n45440 , n19318 , n18324 );
nor ( n45441 , n45439 , n45440 );
nand ( n45442 , n21011 , n19360 );
nand ( n45443 , n19221 , n21022 );
nand ( n45444 , n45435 , n45441 , n45442 , n45443 );
not ( n45445 , n18327 );
nor ( n45446 , n45445 , n19388 );
nor ( n45447 , n45444 , n45446 );
nand ( n45448 , n45434 , n45447 );
buf ( n45449 , n45448 );
buf ( n45450 , n45449 );
not ( n45451 , n275550 );
buf ( n45452 , n45451 );
buf ( n45453 , n45452 );
not ( n45454 , n275929 );
buf ( n45455 , n45454 );
buf ( n45456 , n45455 );
buf ( n45457 , n275554 );
not ( n45458 , n275925 );
buf ( n45459 , n45458 );
buf ( n45460 , n45459 );
not ( n45461 , n275929 );
buf ( n45462 , n45461 );
buf ( n45463 , n45462 );
buf ( n45464 , n275554 );
not ( n45465 , n275925 );
buf ( n45466 , n45465 );
buf ( n45467 , n45466 );
buf ( n45468 , n275554 );
not ( n45469 , n275550 );
buf ( n45470 , n45469 );
buf ( n45471 , n45470 );
or ( n45472 , n24683 , n26364 );
nand ( n45473 , n24696 , n26370 );
nand ( n45474 , n24710 , n26374 );
nand ( n45475 , n35658 , n40881 );
and ( n45476 , n26395 , n24724 );
not ( n45477 , n32188 );
not ( n45478 , n24720 );
or ( n45479 , n45477 , n45478 );
nor ( n45480 , n14830 , n17506 );
not ( n45481 , n45480 );
nand ( n45482 , n45479 , n45481 );
nor ( n45483 , n45476 , n45482 );
nand ( n45484 , n45473 , n45474 , n45475 , n45483 );
not ( n45485 , n45484 );
nand ( n45486 , n45472 , n45485 );
buf ( n45487 , n45486 );
buf ( n45488 , n45487 );
and ( n45489 , n22335 , n18201 );
not ( n45490 , n22335 );
and ( n45491 , n45490 , n29963 );
or ( n45492 , n45489 , n45491 );
buf ( n45493 , n45492 );
buf ( n45494 , n45493 );
buf ( n45495 , n275554 );
not ( n45496 , n26083 );
not ( n45497 , n22335 );
or ( n45498 , n45496 , n45497 );
nand ( n45499 , n20064 , n275557 );
nand ( n45500 , n45498 , n45499 );
buf ( n45501 , n45500 );
buf ( n45502 , n45501 );
not ( n45503 , n275550 );
buf ( n45504 , n45503 );
buf ( n45505 , n45504 );
and ( n45506 , n275745 , n275741 );
not ( n45507 , n275745 );
and ( n45508 , n45507 , n275742 );
nor ( n45509 , n45506 , n45508 );
xor ( n45510 , n45509 , n275751 );
buf ( n45511 , n45510 );
buf ( n45512 , n45511 );
not ( n45513 , n14795 );
or ( n45514 , n45513 , n29046 );
nand ( n45515 , n29044 , n9757 );
nand ( n45516 , n45514 , n45515 );
buf ( n45517 , n45516 );
buf ( n45518 , n45517 );
nand ( n45519 , n23602 , n28408 );
nand ( n45520 , n23654 , n32751 );
nand ( n45521 , n23671 , n29163 );
nand ( n45522 , n28451 , n33882 );
and ( n45523 , n32755 , n23676 );
or ( n45524 , n32757 , n12258 );
nand ( n45525 , n45524 , n36477 );
nor ( n45526 , n45523 , n45525 );
and ( n45527 , n45521 , n45522 , n45526 );
nand ( n45528 , n45519 , n45520 , n45527 );
buf ( n45529 , n45528 );
buf ( n45530 , n45529 );
or ( n45531 , n20673 , n26363 );
nand ( n45532 , n39065 , n14761 );
not ( n45533 , n26385 );
and ( n45534 , n45533 , n20680 );
and ( n45535 , n26367 , n20697 );
and ( n45536 , n26374 , n20687 );
nor ( n45537 , n45534 , n45535 , n45536 );
nand ( n45538 , n45531 , n45532 , n45537 );
buf ( n45539 , n45538 );
buf ( n45540 , n45539 );
not ( n45541 , n275925 );
buf ( n45542 , n45541 );
buf ( n45543 , n45542 );
or ( n45544 , n38543 , n28146 );
nand ( n45545 , n24452 , n18412 );
nand ( n45546 , n45544 , n45545 );
buf ( n45547 , n45546 );
buf ( n45548 , n45547 );
not ( n45549 , n11570 );
or ( n45550 , n45549 , n9158 );
or ( n45551 , n36038 , n9157 );
nand ( n45552 , n45550 , n45551 );
buf ( n45553 , n45552 );
buf ( n45554 , n45553 );
not ( n45555 , n275925 );
buf ( n45556 , n45555 );
buf ( n45557 , n45556 );
or ( n45558 , n22146 , n22158 );
nand ( n45559 , n45558 , n23685 );
buf ( n45560 , n45559 );
buf ( n45561 , n45560 );
not ( n45562 , n275550 );
buf ( n45563 , n45562 );
buf ( n45564 , n45563 );
not ( n45565 , n275550 );
buf ( n45566 , n45565 );
buf ( n45567 , n45566 );
not ( n45568 , n275929 );
buf ( n45569 , n45568 );
buf ( n45570 , n45569 );
buf ( n45571 , n275554 );
and ( n45572 , n22904 , n275864 );
nor ( n45573 , n45572 , n45348 );
nand ( n45574 , n22914 , n31496 );
buf ( n45575 , n31502 );
not ( n45576 , n45575 );
buf ( n45577 , n31534 );
nand ( n45578 , n45576 , n45577 );
buf ( n45579 , n45578 );
buf ( n45580 , n45579 );
not ( n45581 , n45580 );
buf ( n45582 , n23137 );
not ( n45583 , n45582 );
buf ( n45584 , n45583 );
buf ( n45585 , n45584 );
buf ( n45586 , n22924 );
or ( n45587 , n45585 , n45586 );
buf ( n45588 , n22924 );
not ( n45589 , n45588 );
buf ( n45590 , n31493 );
buf ( n45591 , n30540 );
nand ( n45592 , n45589 , n45590 , n45591 );
buf ( n45593 , n45592 );
buf ( n45594 , n45593 );
buf ( n45595 , n22930 );
nand ( n45596 , n45587 , n45594 , n45595 );
buf ( n45597 , n45596 );
buf ( n45598 , n45597 );
not ( n45599 , n45598 );
or ( n45600 , n45581 , n45599 );
buf ( n45601 , n45597 );
buf ( n45602 , n45579 );
or ( n45603 , n45601 , n45602 );
nand ( n45604 , n45600 , n45603 );
buf ( n45605 , n45604 );
buf ( n45606 , n45605 );
nand ( n45607 , n22918 , n45606 );
buf ( n45608 , n31595 );
not ( n45609 , n45608 );
buf ( n45610 , n31626 );
nand ( n45611 , n45609 , n45610 );
buf ( n45612 , n45611 );
buf ( n45613 , n45612 );
not ( n45614 , n45613 );
buf ( n45615 , n23362 );
not ( n45616 , n45615 );
buf ( n45617 , n45616 );
buf ( n45618 , n45617 );
buf ( n45619 , n23158 );
or ( n45620 , n45618 , n45619 );
buf ( n45621 , n23158 );
not ( n45622 , n45621 );
buf ( n45623 , n31587 );
buf ( n45624 , n30574 );
nand ( n45625 , n45622 , n45623 , n45624 );
buf ( n45626 , n45625 );
buf ( n45627 , n45626 );
buf ( n45628 , n23164 );
nand ( n45629 , n45620 , n45627 , n45628 );
buf ( n45630 , n45629 );
buf ( n45631 , n45630 );
not ( n45632 , n45631 );
or ( n45633 , n45614 , n45632 );
buf ( n45634 , n45630 );
buf ( n45635 , n45612 );
or ( n45636 , n45634 , n45635 );
nand ( n45637 , n45633 , n45636 );
buf ( n45638 , n45637 );
buf ( n45639 , n45638 );
nand ( n45640 , n23152 , n45639 );
nand ( n45641 , n45573 , n45574 , n45607 , n45640 );
buf ( n45642 , n45641 );
buf ( n45643 , n45642 );
not ( n45644 , n275929 );
buf ( n45645 , n45644 );
buf ( n45646 , n45645 );
not ( n45647 , n275925 );
buf ( n45648 , n45647 );
buf ( n45649 , n45648 );
not ( n45650 , n24452 );
not ( n45651 , n18715 );
or ( n45652 , n45650 , n45651 );
or ( n45653 , n21629 , n28146 );
nand ( n45654 , n45652 , n45653 );
buf ( n45655 , n45654 );
buf ( n45656 , n45655 );
not ( n45657 , n275929 );
buf ( n45658 , n45657 );
buf ( n45659 , n45658 );
buf ( n45660 , n275554 );
not ( n45661 , n21080 );
or ( n45662 , n45661 , n21774 );
nand ( n45663 , n21774 , n9544 );
nand ( n45664 , n45662 , n45663 );
buf ( n45665 , n45664 );
buf ( n45666 , n45665 );
and ( n45667 , n9158 , n9072 );
not ( n45668 , n9158 );
and ( n45669 , n45668 , n277747 );
or ( n45670 , n45667 , n45669 );
buf ( n45671 , n45670 );
buf ( n45672 , n45671 );
buf ( n45673 , n275554 );
buf ( n45674 , n275554 );
or ( n45675 , n36036 , n40803 );
not ( n45676 , n36046 );
and ( n45677 , n45676 , n275605 );
nand ( n45678 , n36066 , n36145 );
not ( n45679 , n45678 );
not ( n45680 , n36137 );
or ( n45681 , n45680 , n36060 );
not ( n45682 , n36140 );
nand ( n45683 , n45681 , n45682 );
not ( n45684 , n45683 );
or ( n45685 , n45679 , n45684 );
or ( n45686 , n45683 , n45678 );
nand ( n45687 , n45685 , n45686 );
buf ( n45688 , n45687 );
not ( n45689 , n45688 );
not ( n45690 , n36155 );
or ( n45691 , n45689 , n45690 );
nand ( n45692 , n36177 , n36251 );
not ( n45693 , n45692 );
not ( n45694 , n36243 );
or ( n45695 , n45694 , n36172 );
not ( n45696 , n36246 );
nand ( n45697 , n45695 , n45696 );
not ( n45698 , n45697 );
or ( n45699 , n45693 , n45698 );
or ( n45700 , n45697 , n45692 );
nand ( n45701 , n45699 , n45700 );
buf ( n45702 , n45701 );
nand ( n45703 , n41635 , n45702 );
nand ( n45704 , n45691 , n45703 );
nor ( n45705 , n45677 , n45704 );
nand ( n45706 , n45675 , n45705 );
nand ( n45707 , n45706 , n20645 );
nand ( n45708 , n36280 , n36361 );
not ( n45709 , n45708 );
not ( n45710 , n36353 );
not ( n45711 , n36284 );
or ( n45712 , n45710 , n45711 );
not ( n45713 , n36356 );
nand ( n45714 , n45712 , n45713 );
not ( n45715 , n45714 );
or ( n45716 , n45709 , n45715 );
or ( n45717 , n45714 , n45708 );
nand ( n45718 , n45716 , n45717 );
buf ( n45719 , n45718 );
nand ( n45720 , n36267 , n45719 );
nand ( n45721 , n36384 , n36464 );
not ( n45722 , n45721 );
not ( n45723 , n36456 );
not ( n45724 , n36388 );
or ( n45725 , n45723 , n45724 );
nand ( n45726 , n45725 , n36460 );
not ( n45727 , n45726 );
or ( n45728 , n45722 , n45727 );
or ( n45729 , n45726 , n45721 );
nand ( n45730 , n45728 , n45729 );
buf ( n45731 , n45730 );
nand ( n45732 , n36371 , n45731 );
and ( n45733 , n36474 , n36064 );
or ( n45734 , n20654 , n275604 );
nand ( n45735 , n45734 , n40183 );
nor ( n45736 , n45733 , n45735 );
nand ( n45737 , n45707 , n45720 , n45732 , n45736 );
buf ( n45738 , n45737 );
buf ( n45739 , n45738 );
not ( n45740 , n275925 );
buf ( n45741 , n45740 );
buf ( n45742 , n45741 );
or ( n45743 , n40492 , n31719 );
or ( n45744 , n35071 , n11418 );
nand ( n45745 , n45743 , n45744 );
buf ( n45746 , n45745 );
buf ( n45747 , n45746 );
or ( n45748 , n32728 , n31719 );
or ( n45749 , n35071 , n11382 );
nand ( n45750 , n45748 , n45749 );
buf ( n45751 , n45750 );
buf ( n45752 , n45751 );
and ( n45753 , n37271 , n31682 );
nor ( n45754 , n45753 , n31177 );
buf ( n45755 , n37316 );
buf ( n45756 , n37337 );
and ( n45757 , n45755 , n45756 );
buf ( n45758 , n45757 );
buf ( n45759 , n45758 );
not ( n45760 , n45759 );
buf ( n45761 , n31493 );
buf ( n45762 , n37305 );
buf ( n45763 , n30540 );
and ( n45764 , n45761 , n45762 , n45763 );
buf ( n45765 , n45584 );
buf ( n45766 , n37302 );
or ( n45767 , n45765 , n45766 );
buf ( n45768 , n37330 );
nand ( n45769 , n45767 , n45768 );
buf ( n45770 , n45769 );
buf ( n45771 , n45770 );
nor ( n45772 , n45764 , n45771 );
buf ( n45773 , n45772 );
buf ( n45774 , n45773 );
not ( n45775 , n45774 );
or ( n45776 , n45760 , n45775 );
buf ( n45777 , n45773 );
buf ( n45778 , n45758 );
or ( n45779 , n45777 , n45778 );
nand ( n45780 , n45776 , n45779 );
buf ( n45781 , n45780 );
buf ( n45782 , n45781 );
nand ( n45783 , n22918 , n45782 );
nand ( n45784 , n22914 , n34525 );
buf ( n45785 , n37391 );
buf ( n45786 , n37412 );
and ( n45787 , n45785 , n45786 );
buf ( n45788 , n45787 );
buf ( n45789 , n45788 );
not ( n45790 , n45789 );
buf ( n45791 , n31587 );
buf ( n45792 , n37381 );
buf ( n45793 , n30574 );
and ( n45794 , n45791 , n45792 , n45793 );
buf ( n45795 , n45617 );
buf ( n45796 , n37378 );
or ( n45797 , n45795 , n45796 );
buf ( n45798 , n37405 );
nand ( n45799 , n45797 , n45798 );
buf ( n45800 , n45799 );
buf ( n45801 , n45800 );
nor ( n45802 , n45794 , n45801 );
buf ( n45803 , n45802 );
buf ( n45804 , n45803 );
not ( n45805 , n45804 );
or ( n45806 , n45790 , n45805 );
buf ( n45807 , n45803 );
buf ( n45808 , n45788 );
or ( n45809 , n45807 , n45808 );
nand ( n45810 , n45806 , n45809 );
buf ( n45811 , n45810 );
buf ( n45812 , n45811 );
nand ( n45813 , n23152 , n45812 );
nand ( n45814 , n45754 , n45783 , n45784 , n45813 );
buf ( n45815 , n45814 );
buf ( n45816 , n45815 );
buf ( n45817 , n275554 );
buf ( n45818 , n275554 );
not ( n45819 , n275550 );
buf ( n45820 , n45819 );
buf ( n45821 , n45820 );
buf ( n45822 , n275554 );
buf ( n45823 , n275554 );
buf ( n45824 , n275554 );
buf ( n45825 , n275554 );
and ( n45826 , n9158 , n9117 );
not ( n45827 , n9158 );
and ( n45828 , n45827 , n277820 );
or ( n45829 , n45826 , n45828 );
buf ( n45830 , n45829 );
buf ( n45831 , n45830 );
buf ( n45832 , n275554 );
buf ( n45833 , n275554 );
or ( n45834 , n38515 , n21030 );
nand ( n45835 , n21030 , n18497 );
nand ( n45836 , n45834 , n45835 );
buf ( n45837 , n45836 );
buf ( n45838 , n45837 );
not ( n45839 , n275929 );
buf ( n45840 , n45839 );
buf ( n45841 , n45840 );
buf ( n45842 , n275554 );
not ( n45843 , n275550 );
buf ( n45844 , n45843 );
buf ( n45845 , n45844 );
not ( n45846 , n275550 );
buf ( n45847 , n45846 );
buf ( n45848 , n45847 );
not ( n45849 , n275925 );
buf ( n45850 , n45849 );
buf ( n45851 , n45850 );
buf ( n45852 , n275554 );
buf ( n45853 , n275554 );
buf ( n45854 , n275554 );
or ( n45855 , n44898 , n21696 );
nand ( n45856 , n21696 , n13568 );
nand ( n45857 , n45855 , n45856 );
buf ( n45858 , n45857 );
buf ( n45859 , n45858 );
buf ( n45860 , n275554 );
buf ( n45861 , n275554 );
or ( n45862 , n36036 , n39119 );
and ( n45863 , n45676 , n275693 );
not ( n45864 , n36125 );
nand ( n45865 , n45864 , n36129 );
not ( n45866 , n45865 );
not ( n45867 , n36133 );
nand ( n45868 , n45867 , n36112 );
not ( n45869 , n45868 );
or ( n45870 , n45866 , n45869 );
or ( n45871 , n45868 , n45865 );
nand ( n45872 , n45870 , n45871 );
buf ( n45873 , n45872 );
not ( n45874 , n45873 );
not ( n45875 , n36155 );
or ( n45876 , n45874 , n45875 );
not ( n45877 , n36231 );
nand ( n45878 , n45877 , n36235 );
not ( n45879 , n45878 );
not ( n45880 , n36239 );
nand ( n45881 , n45880 , n36218 );
not ( n45882 , n45881 );
or ( n45883 , n45879 , n45882 );
or ( n45884 , n45881 , n45878 );
nand ( n45885 , n45883 , n45884 );
buf ( n45886 , n45885 );
nand ( n45887 , n36159 , n45886 );
nand ( n45888 , n45876 , n45887 );
nor ( n45889 , n45863 , n45888 );
nand ( n45890 , n45862 , n45889 );
nand ( n45891 , n45890 , n20645 );
nand ( n45892 , n36320 , n36300 );
not ( n45893 , n45892 );
not ( n45894 , n36310 );
nand ( n45895 , n45894 , n36308 );
not ( n45896 , n45895 );
or ( n45897 , n45893 , n45896 );
or ( n45898 , n45895 , n45892 );
nand ( n45899 , n45897 , n45898 );
buf ( n45900 , n45899 );
nand ( n45901 , n36267 , n45900 );
nand ( n45902 , n36423 , n41657 );
not ( n45903 , n45902 );
not ( n45904 , n36413 );
nand ( n45905 , n45904 , n36411 );
not ( n45906 , n45905 );
or ( n45907 , n45903 , n45906 );
or ( n45908 , n45905 , n45902 );
nand ( n45909 , n45907 , n45908 );
buf ( n45910 , n45909 );
nand ( n45911 , n36371 , n45910 );
and ( n45912 , n36474 , n36110 );
or ( n45913 , n20654 , n275692 );
nand ( n45914 , n45913 , n31787 );
nor ( n45915 , n45912 , n45914 );
nand ( n45916 , n45891 , n45901 , n45911 , n45915 );
buf ( n45917 , n45916 );
buf ( n45918 , n45917 );
buf ( n45919 , n275554 );
or ( n45920 , n32272 , n20743 );
and ( n45921 , n20763 , n32309 );
not ( n45922 , n20765 );
not ( n45923 , n32314 );
and ( n45924 , n45922 , n45923 );
and ( n45925 , n17411 , n32323 );
nor ( n45926 , n45924 , n45925 );
nand ( n45927 , n17502 , n32327 );
nand ( n45928 , n17560 , n13893 );
nand ( n45929 , n45926 , n45927 , n45928 );
nor ( n45930 , n45921 , n45929 );
nand ( n45931 , n32290 , n16970 );
and ( n45932 , n45930 , n45931 );
nand ( n45933 , n45920 , n45932 );
buf ( n45934 , n45933 );
buf ( n45935 , n45934 );
buf ( n45936 , n30506 );
buf ( n45937 , n45936 );
not ( n45938 , n45937 );
not ( n45939 , n19066 );
nand ( n45940 , n45939 , n34151 );
buf ( n45941 , n45940 );
not ( n45942 , n45941 );
or ( n45943 , n45938 , n45942 );
not ( n45944 , n19066 );
nand ( n45945 , n45944 , n34151 );
buf ( n45946 , n45945 );
buf ( n45947 , n45946 );
buf ( n45948 , n19992 );
not ( n45949 , n45948 );
buf ( n45950 , n20114 );
buf ( n45951 , n20428 );
nand ( n45952 , n45950 , n45951 );
not ( n45953 , n45952 );
buf ( n45954 , n20109 );
buf ( n45955 , n45954 );
buf ( n45956 , n18919 );
buf ( n45957 , n45956 );
nand ( n45958 , n45955 , n45957 );
buf ( n45959 , n45958 );
not ( n45960 , n45959 );
buf ( n45961 , n20207 );
nand ( n45962 , n45953 , n45960 , n45961 );
not ( n45963 , n45962 );
or ( n45964 , n45949 , n45963 );
or ( n45965 , n45962 , n45948 );
nand ( n45966 , n45964 , n45965 );
buf ( n45967 , n45966 );
not ( n45968 , n45967 );
or ( n45969 , n45947 , n45968 );
nand ( n45970 , n45943 , n45969 );
buf ( n45971 , n45970 );
buf ( n45972 , n22871 );
not ( n45973 , n45972 );
nor ( n45974 , n45971 , n45973 );
not ( n45975 , n45946 );
not ( n45976 , n45975 );
nor ( n45977 , n45952 , n45959 );
xor ( n45978 , n45977 , n45961 );
buf ( n45979 , n45978 );
not ( n45980 , n45979 );
or ( n45981 , n45976 , n45980 );
buf ( n45982 , n22800 );
buf ( n45983 , n45982 );
nand ( n45984 , n45941 , n45983 );
nand ( n45985 , n45981 , n45984 );
buf ( n45986 , n45985 );
buf ( n45987 , n35188 );
not ( n45988 , n45987 );
nor ( n45989 , n45986 , n45988 );
nor ( n45990 , n45974 , n45989 );
not ( n45991 , n45975 );
not ( n45992 , n45951 );
nand ( n45993 , n45960 , n45950 );
not ( n45994 , n45993 );
or ( n45995 , n45992 , n45994 );
or ( n45996 , n45993 , n45951 );
nand ( n45997 , n45995 , n45996 );
buf ( n45998 , n45997 );
not ( n45999 , n45998 );
or ( n46000 , n45991 , n45999 );
not ( n46001 , n45940 );
not ( n46002 , n46001 );
buf ( n46003 , n35121 );
buf ( n46004 , n46003 );
nand ( n46005 , n46002 , n46004 );
nand ( n46006 , n46000 , n46005 );
buf ( n46007 , n46006 );
buf ( n46008 , n24442 );
not ( n46009 , n46008 );
nor ( n46010 , n46007 , n46009 );
not ( n46011 , n45950 );
not ( n46012 , n45959 );
or ( n46013 , n46011 , n46012 );
or ( n46014 , n45959 , n45950 );
nand ( n46015 , n46013 , n46014 );
buf ( n46016 , n46015 );
not ( n46017 , n46016 );
or ( n46018 , n45991 , n46017 );
buf ( n46019 , n24386 );
buf ( n46020 , n46019 );
nand ( n46021 , n45941 , n46020 );
nand ( n46022 , n46018 , n46021 );
buf ( n46023 , n46022 );
buf ( n46024 , n30628 );
not ( n46025 , n46024 );
nor ( n46026 , n46023 , n46025 );
nor ( n46027 , n46010 , n46026 );
not ( n46028 , n45946 );
not ( n46029 , n46028 );
not ( n46030 , n45955 );
not ( n46031 , n45957 );
and ( n46032 , n46030 , n46031 );
nor ( n46033 , n46032 , n45960 );
buf ( n46034 , n46033 );
not ( n46035 , n46034 );
or ( n46036 , n46029 , n46035 );
buf ( n46037 , n30599 );
buf ( n46038 , n46037 );
nand ( n46039 , n46002 , n46038 );
nand ( n46040 , n46036 , n46039 );
buf ( n46041 , n46040 );
buf ( n46042 , n34029 );
not ( n46043 , n46042 );
nor ( n46044 , n46041 , n46043 );
buf ( n46045 , n24645 );
not ( n46046 , n46045 );
buf ( n46047 , n18309 );
nor ( n46048 , n46046 , n46047 );
buf ( n46049 , n19092 );
not ( n46050 , n46049 );
buf ( n46051 , n19286 );
and ( n46052 , n46050 , n46051 );
or ( n46053 , n46048 , n46052 );
or ( n46054 , n46050 , n46051 );
nand ( n46055 , n46053 , n46054 );
buf ( n46056 , n33980 );
buf ( n46057 , n46056 );
not ( n46058 , n46057 );
buf ( n46059 , n21022 );
nand ( n46060 , n46058 , n46059 );
and ( n46061 , n46055 , n46060 );
not ( n46062 , n46059 );
and ( n46063 , n46057 , n46062 );
nor ( n46064 , n46061 , n46063 );
or ( n46065 , n46044 , n46064 );
nand ( n46066 , n46041 , n46043 );
nand ( n46067 , n46065 , n46066 );
nand ( n46068 , n45990 , n46027 , n46067 );
not ( n46069 , n46024 );
nand ( n46070 , n46069 , n46023 );
not ( n46071 , n46008 );
nand ( n46072 , n46071 , n46007 );
and ( n46073 , n46070 , n46072 );
nor ( n46074 , n46073 , n46010 );
nand ( n46075 , n46074 , n45990 );
not ( n46076 , n45974 );
and ( n46077 , n45986 , n45988 );
and ( n46078 , n46076 , n46077 );
and ( n46079 , n45971 , n45973 );
nor ( n46080 , n46078 , n46079 );
nand ( n46081 , n46068 , n46075 , n46080 );
not ( n46082 , n46081 );
not ( n46083 , n46028 );
not ( n46084 , n45952 );
nand ( n46085 , n45961 , n45948 );
nor ( n46086 , n45958 , n46085 );
buf ( n46087 , n46086 );
nand ( n46088 , n46084 , n46087 );
buf ( n46089 , n21366 );
buf ( n46090 , n19668 );
and ( n46091 , n46089 , n46090 );
buf ( n46092 , n19937 );
buf ( n46093 , n19952 );
buf ( n46094 , n46093 );
nand ( n46095 , n46092 , n46094 );
not ( n46096 , n46095 );
nand ( n46097 , n46091 , n46096 );
nor ( n46098 , n46088 , n46097 );
buf ( n46099 , n21356 );
buf ( n46100 , n46099 );
buf ( n46101 , n21418 );
buf ( n46102 , n46101 );
nand ( n46103 , n46100 , n46102 );
buf ( n46104 , n21307 );
buf ( n46105 , n46104 );
not ( n46106 , n46105 );
nor ( n46107 , n46103 , n46106 );
nand ( n46108 , n46098 , n46107 );
buf ( n46109 , n24158 );
buf ( n46110 , n46109 );
not ( n46111 , n46110 );
and ( n46112 , n46108 , n46111 );
not ( n46113 , n46108 );
and ( n46114 , n46113 , n46110 );
nor ( n46115 , n46112 , n46114 );
buf ( n46116 , n46115 );
not ( n46117 , n46116 );
or ( n46118 , n46083 , n46117 );
buf ( n46119 , n33794 );
buf ( n46120 , n46119 );
nand ( n46121 , n45941 , n46120 );
nand ( n46122 , n46118 , n46121 );
buf ( n46123 , n46122 );
buf ( n46124 , n37641 );
not ( n46125 , n46124 );
nor ( n46126 , n46123 , n46125 );
buf ( n46127 , n21624 );
not ( n46128 , n46127 );
not ( n46129 , n46088 );
nor ( n46130 , n46097 , n46103 );
nand ( n46131 , n46129 , n46130 );
and ( n46132 , n46131 , n46106 );
not ( n46133 , n46131 );
and ( n46134 , n46133 , n46105 );
nor ( n46135 , n46132 , n46134 );
buf ( n46136 , n46135 );
not ( n46137 , n46136 );
or ( n46138 , n46029 , n46137 );
buf ( n46139 , n35964 );
buf ( n46140 , n46139 );
nand ( n46141 , n45947 , n46140 );
nand ( n46142 , n46138 , n46141 );
buf ( n46143 , n46142 );
nor ( n46144 , n46128 , n46143 );
nor ( n46145 , n46126 , n46144 );
buf ( n46146 , n46100 );
not ( n46147 , n46146 );
not ( n46148 , n46088 );
not ( n46149 , n46102 );
nor ( n46150 , n46097 , n46149 );
nand ( n46151 , n46148 , n46150 );
not ( n46152 , n46151 );
or ( n46153 , n46147 , n46152 );
or ( n46154 , n46151 , n46146 );
nand ( n46155 , n46153 , n46154 );
buf ( n46156 , n46155 );
not ( n46157 , n46156 );
or ( n46158 , n46083 , n46157 );
buf ( n46159 , n21080 );
buf ( n46160 , n46159 );
nand ( n46161 , n45941 , n46160 );
nand ( n46162 , n46158 , n46161 );
buf ( n46163 , n46162 );
buf ( n46164 , n29548 );
not ( n46165 , n46164 );
nor ( n46166 , n46163 , n46165 );
buf ( n46167 , n29459 );
not ( n46168 , n46167 );
and ( n46169 , n46098 , n46102 );
not ( n46170 , n46098 );
and ( n46171 , n46170 , n46149 );
nor ( n46172 , n46169 , n46171 );
buf ( n46173 , n46172 );
not ( n46174 , n46173 );
or ( n46175 , n46083 , n46174 );
buf ( n46176 , n29506 );
buf ( n46177 , n46176 );
nand ( n46178 , n46002 , n46177 );
nand ( n46179 , n46175 , n46178 );
buf ( n46180 , n46179 );
nor ( n46181 , n46168 , n46180 );
nor ( n46182 , n46166 , n46181 );
nand ( n46183 , n46145 , n46182 );
not ( n46184 , n46088 );
not ( n46185 , n46090 );
nor ( n46186 , n46095 , n46185 );
nand ( n46187 , n46184 , n46186 );
buf ( n46188 , n46089 );
xnor ( n46189 , n46187 , n46188 );
buf ( n46190 , n46189 );
not ( n46191 , n46190 );
or ( n46192 , n45941 , n46191 );
not ( n46193 , n46001 );
buf ( n46194 , n29394 );
not ( n46195 , n46194 );
buf ( n46196 , n46195 );
nand ( n46197 , n46193 , n46196 );
nand ( n46198 , n46192 , n46197 );
buf ( n46199 , n46198 );
buf ( n46200 , n39294 );
not ( n46201 , n46200 );
nor ( n46202 , n46199 , n46201 );
buf ( n46203 , n39236 );
buf ( n46204 , n46203 );
not ( n46205 , n46204 );
not ( n46206 , n45941 );
or ( n46207 , n46205 , n46206 );
buf ( n46208 , n46088 );
not ( n46209 , n46208 );
nand ( n46210 , n46209 , n46096 );
and ( n46211 , n46210 , n46185 );
not ( n46212 , n46210 );
and ( n46213 , n46212 , n46090 );
nor ( n46214 , n46211 , n46213 );
buf ( n46215 , n46214 );
not ( n46216 , n46215 );
or ( n46217 , n45941 , n46216 );
nand ( n46218 , n46207 , n46217 );
buf ( n46219 , n46218 );
buf ( n46220 , n20566 );
not ( n46221 , n46220 );
nor ( n46222 , n46219 , n46221 );
nor ( n46223 , n46202 , n46222 );
buf ( n46224 , n19429 );
buf ( n46225 , n46224 );
not ( n46226 , n46225 );
not ( n46227 , n46002 );
or ( n46228 , n46226 , n46227 );
buf ( n46229 , n45946 );
nand ( n46230 , n46184 , n46094 );
xnor ( n46231 , n46230 , n46092 );
buf ( n46232 , n46231 );
not ( n46233 , n46232 );
or ( n46234 , n46229 , n46233 );
nand ( n46235 , n46228 , n46234 );
buf ( n46236 , n46235 );
buf ( n46237 , n35837 );
not ( n46238 , n46237 );
nor ( n46239 , n46236 , n46238 );
and ( n46240 , n46094 , n46209 );
not ( n46241 , n46094 );
and ( n46242 , n46241 , n46208 );
nor ( n46243 , n46240 , n46242 );
buf ( n46244 , n46243 );
not ( n46245 , n46244 );
or ( n46246 , n45976 , n46245 );
buf ( n46247 , n35800 );
buf ( n46248 , n46247 );
nand ( n46249 , n45947 , n46248 );
nand ( n46250 , n46246 , n46249 );
buf ( n46251 , n46250 );
buf ( n46252 , n35714 );
not ( n46253 , n46252 );
nor ( n46254 , n46251 , n46253 );
nor ( n46255 , n46239 , n46254 );
nand ( n46256 , n46223 , n46255 );
nor ( n46257 , n46183 , n46256 );
not ( n46258 , n46257 );
or ( n46259 , n46082 , n46258 );
not ( n46260 , n46183 );
not ( n46261 , n46223 );
not ( n46262 , n46237 );
nand ( n46263 , n46262 , n46236 );
not ( n46264 , n46263 );
nand ( n46265 , n46251 , n46253 );
not ( n46266 , n46265 );
or ( n46267 , n46264 , n46266 );
not ( n46268 , n46239 );
nand ( n46269 , n46267 , n46268 );
or ( n46270 , n46261 , n46269 );
not ( n46271 , n46220 );
nand ( n46272 , n46271 , n46219 );
or ( n46273 , n46202 , n46272 );
nand ( n46274 , n46199 , n46201 );
nand ( n46275 , n46273 , n46274 );
not ( n46276 , n46275 );
nand ( n46277 , n46270 , n46276 );
and ( n46278 , n46260 , n46277 );
not ( n46279 , n46145 );
not ( n46280 , n46167 );
nand ( n46281 , n46280 , n46180 );
or ( n46282 , n46166 , n46281 );
nand ( n46283 , n46163 , n46165 );
nand ( n46284 , n46282 , n46283 );
not ( n46285 , n46284 );
or ( n46286 , n46279 , n46285 );
not ( n46287 , n46126 );
not ( n46288 , n46127 );
nand ( n46289 , n46288 , n46143 );
not ( n46290 , n46289 );
and ( n46291 , n46287 , n46290 );
and ( n46292 , n46123 , n46125 );
nor ( n46293 , n46291 , n46292 );
nand ( n46294 , n46286 , n46293 );
nor ( n46295 , n46278 , n46294 );
nand ( n46296 , n46259 , n46295 );
buf ( n46297 , n30177 );
not ( n46298 , n46297 );
not ( n46299 , n29856 );
not ( n46300 , n46001 );
not ( n46301 , n46300 );
or ( n46302 , n46299 , n46301 );
nand ( n46303 , n46110 , n46105 );
nor ( n46304 , n46103 , n46303 );
nor ( n46305 , n45952 , n46095 );
nand ( n46306 , n46304 , n46086 , n46305 , n46091 );
not ( n46307 , n46306 );
buf ( n46308 , n24055 );
buf ( n46309 , n46308 );
buf ( n46310 , n24091 );
buf ( n46311 , n46310 );
nand ( n46312 , n46309 , n46311 );
buf ( n46313 , n28000 );
buf ( n46314 , n46313 );
buf ( n46315 , n26691 );
buf ( n46316 , n46315 );
nand ( n46317 , n46314 , n46316 );
nor ( n46318 , n46312 , n46317 );
buf ( n46319 , n26796 );
buf ( n46320 , n46319 );
buf ( n46321 , n26860 );
buf ( n46322 , n46321 );
nand ( n46323 , n46320 , n46322 );
buf ( n46324 , n26683 );
buf ( n46325 , n46324 );
buf ( n46326 , n26788 );
buf ( n46327 , n46326 );
nand ( n46328 , n46325 , n46327 );
nor ( n46329 , n46323 , n46328 );
nand ( n46330 , n46318 , n46329 );
buf ( n46331 , n28055 );
buf ( n46332 , n46331 );
buf ( n46333 , n28052 );
buf ( n46334 , n46333 );
nand ( n46335 , n46332 , n46334 );
buf ( n46336 , n30086 );
buf ( n46337 , n46336 );
buf ( n46338 , n30078 );
nand ( n46339 , n46337 , n46338 );
nor ( n46340 , n46335 , n46339 );
not ( n46341 , n46340 );
nor ( n46342 , n46330 , n46341 );
nand ( n46343 , n46307 , n46342 );
buf ( n46344 , n29967 );
not ( n46345 , n46344 );
and ( n46346 , n46343 , n46345 );
not ( n46347 , n46343 );
and ( n46348 , n46347 , n46344 );
nor ( n46349 , n46346 , n46348 );
buf ( n46350 , n46349 );
not ( n46351 , n46350 );
or ( n46352 , n46229 , n46351 );
nand ( n46353 , n46302 , n46352 );
buf ( n46354 , n46353 );
not ( n46355 , n46354 );
not ( n46356 , n46355 );
or ( n46357 , n46298 , n46356 );
not ( n46358 , n29820 );
and ( n46359 , n46300 , n46358 );
not ( n46360 , n46300 );
and ( n46361 , n46340 , n46344 );
not ( n46362 , n46330 );
nand ( n46363 , n46307 , n46361 , n46362 );
buf ( n46364 , n40952 );
not ( n46365 , n46364 );
and ( n46366 , n46363 , n46365 );
not ( n46367 , n46363 );
and ( n46368 , n46367 , n46364 );
nor ( n46369 , n46366 , n46368 );
buf ( n46370 , n46369 );
not ( n46371 , n46370 );
and ( n46372 , n46360 , n46371 );
nor ( n46373 , n46359 , n46372 );
buf ( n46374 , n46373 );
not ( n46375 , n46374 );
buf ( n46376 , n41034 );
nand ( n46377 , n46375 , n46376 );
nand ( n46378 , n46357 , n46377 );
buf ( n46379 , n34244 );
not ( n46380 , n46379 );
nand ( n46381 , n46344 , n46364 );
nor ( n46382 , n46341 , n46381 );
nand ( n46383 , n46307 , n46382 , n46362 );
buf ( n46384 , n18848 );
buf ( n46385 , n46384 );
and ( n46386 , n46383 , n46385 );
not ( n46387 , n46383 );
not ( n46388 , n46385 );
and ( n46389 , n46387 , n46388 );
nor ( n46390 , n46386 , n46389 );
buf ( n46391 , n46390 );
not ( n46392 , n46391 );
or ( n46393 , n45941 , n46392 );
buf ( n46394 , n34151 );
nand ( n46395 , n46002 , n46394 );
nand ( n46396 , n46393 , n46395 );
buf ( n46397 , n46396 );
not ( n46398 , n46397 );
not ( n46399 , n46398 );
or ( n46400 , n46380 , n46399 );
buf ( n46401 , n19054 );
buf ( n46402 , n46401 );
not ( n46403 , n46402 );
and ( n46404 , n46403 , n46388 );
not ( n46405 , n46403 );
and ( n46406 , n46405 , n46385 );
nor ( n46407 , n46404 , n46406 );
not ( n46408 , n46407 );
nor ( n46409 , n46381 , n46385 );
and ( n46410 , n46340 , n46409 );
nand ( n46411 , n46410 , n46362 );
nor ( n46412 , n46306 , n46411 );
not ( n46413 , n46412 );
or ( n46414 , n46408 , n46413 );
or ( n46415 , n46412 , n46407 );
nand ( n46416 , n46414 , n46415 );
buf ( n46417 , n46416 );
not ( n46418 , n46417 );
not ( n46419 , n45975 );
or ( n46420 , n46418 , n46419 );
nand ( n46421 , n46420 , n45939 );
buf ( n46422 , n46421 );
buf ( n46423 , n34241 );
not ( n46424 , n46423 );
nand ( n46425 , n46422 , n46424 );
nand ( n46426 , n46400 , n46425 );
nor ( n46427 , n46378 , n46426 );
not ( n46428 , n29795 );
not ( n46429 , n46428 );
not ( n46430 , n46429 );
not ( n46431 , n45941 );
or ( n46432 , n46430 , n46431 );
not ( n46433 , n46337 );
nor ( n46434 , n46335 , n46433 );
nand ( n46435 , n46307 , n46362 , n46434 );
not ( n46436 , n46338 );
and ( n46437 , n46435 , n46436 );
not ( n46438 , n46435 );
and ( n46439 , n46438 , n46338 );
nor ( n46440 , n46437 , n46439 );
buf ( n46441 , n46440 );
not ( n46442 , n46441 );
or ( n46443 , n46083 , n46442 );
nand ( n46444 , n46432 , n46443 );
buf ( n46445 , n46444 );
buf ( n46446 , n38125 );
not ( n46447 , n46446 );
nor ( n46448 , n46445 , n46447 );
buf ( n46449 , n27810 );
not ( n46450 , n46449 );
not ( n46451 , n45947 );
or ( n46452 , n46450 , n46451 );
nor ( n46453 , n46330 , n46335 );
nand ( n46454 , n46307 , n46453 );
xor ( n46455 , n46454 , n46433 );
buf ( n46456 , n46455 );
not ( n46457 , n46456 );
or ( n46458 , n46029 , n46457 );
nand ( n46459 , n46452 , n46458 );
buf ( n46460 , n46459 );
buf ( n46461 , n30019 );
not ( n46462 , n46461 );
nor ( n46463 , n46460 , n46462 );
nor ( n46464 , n46448 , n46463 );
buf ( n46465 , n27832 );
not ( n46466 , n46465 );
not ( n46467 , n45941 );
or ( n46468 , n46466 , n46467 );
not ( n46469 , n46332 );
nor ( n46470 , n46330 , n46469 );
nand ( n46471 , n46307 , n46470 );
not ( n46472 , n46334 );
and ( n46473 , n46471 , n46472 );
not ( n46474 , n46471 );
and ( n46475 , n46474 , n46334 );
nor ( n46476 , n46473 , n46475 );
buf ( n46477 , n46476 );
not ( n46478 , n46477 );
or ( n46479 , n46029 , n46478 );
nand ( n46480 , n46468 , n46479 );
buf ( n46481 , n46480 );
buf ( n46482 , n27885 );
not ( n46483 , n46482 );
nor ( n46484 , n46481 , n46483 );
buf ( n46485 , n27783 );
not ( n46486 , n46485 );
not ( n46487 , n45941 );
or ( n46488 , n46486 , n46487 );
nand ( n46489 , n46307 , n46362 );
and ( n46490 , n46489 , n46469 );
not ( n46491 , n46489 );
and ( n46492 , n46491 , n46332 );
nor ( n46493 , n46490 , n46492 );
buf ( n46494 , n46493 );
not ( n46495 , n46494 );
or ( n46496 , n45976 , n46495 );
nand ( n46497 , n46488 , n46496 );
buf ( n46498 , n46497 );
buf ( n46499 , n27932 );
not ( n46500 , n46499 );
nor ( n46501 , n46498 , n46500 );
nor ( n46502 , n46484 , n46501 );
and ( n46503 , n46464 , n46502 );
nand ( n46504 , n46427 , n46503 );
not ( n46505 , n26551 );
not ( n46506 , n46505 );
buf ( n46507 , n46506 );
not ( n46508 , n46507 );
not ( n46509 , n45941 );
or ( n46510 , n46508 , n46509 );
not ( n46511 , n46312 );
not ( n46512 , n46327 );
not ( n46513 , n46320 );
nor ( n46514 , n46512 , n46513 );
nand ( n46515 , n46511 , n46514 );
and ( n46516 , n46322 , n46316 );
nand ( n46517 , n46516 , n46325 );
nor ( n46518 , n46515 , n46517 );
nand ( n46519 , n46518 , n46307 );
buf ( n46520 , n46314 );
not ( n46521 , n46520 );
and ( n46522 , n46519 , n46521 );
not ( n46523 , n46519 );
and ( n46524 , n46523 , n46520 );
nor ( n46525 , n46522 , n46524 );
buf ( n46526 , n46525 );
not ( n46527 , n46526 );
or ( n46528 , n46229 , n46527 );
nand ( n46529 , n46510 , n46528 );
buf ( n46530 , n46529 );
buf ( n46531 , n40409 );
not ( n46532 , n46531 );
nor ( n46533 , n46530 , n46532 );
buf ( n46534 , n27050 );
not ( n46535 , n46534 );
not ( n46536 , n33296 );
buf ( n46537 , n46536 );
not ( n46538 , n46537 );
not ( n46539 , n46002 );
or ( n46540 , n46538 , n46539 );
not ( n46541 , n46516 );
nor ( n46542 , n46541 , n46515 );
nand ( n46543 , n46307 , n46542 );
not ( n46544 , n46325 );
and ( n46545 , n46543 , n46544 );
not ( n46546 , n46543 );
and ( n46547 , n46546 , n46325 );
nor ( n46548 , n46545 , n46547 );
buf ( n46549 , n46548 );
not ( n46550 , n46549 );
or ( n46551 , n45947 , n46550 );
nand ( n46552 , n46540 , n46551 );
buf ( n46553 , n46552 );
nor ( n46554 , n46535 , n46553 );
nor ( n46555 , n46533 , n46554 );
not ( n46556 , n21759 );
buf ( n46557 , n46556 );
not ( n46558 , n46557 );
not ( n46559 , n46002 );
or ( n46560 , n46558 , n46559 );
not ( n46561 , n46322 );
nor ( n46562 , n46515 , n46561 );
nand ( n46563 , n46307 , n46562 );
not ( n46564 , n46316 );
and ( n46565 , n46563 , n46564 );
not ( n46566 , n46563 );
and ( n46567 , n46566 , n46316 );
nor ( n46568 , n46565 , n46567 );
buf ( n46569 , n46568 );
not ( n46570 , n46569 );
or ( n46571 , n45947 , n46570 );
nand ( n46572 , n46560 , n46571 );
buf ( n46573 , n46572 );
buf ( n46574 , n31098 );
not ( n46575 , n46574 );
nor ( n46576 , n46573 , n46575 );
buf ( n46577 , n38739 );
not ( n46578 , n46577 );
not ( n46579 , n46515 );
nand ( n46580 , n46579 , n46307 );
and ( n46581 , n46580 , n46561 );
not ( n46582 , n46580 );
and ( n46583 , n46582 , n46322 );
nor ( n46584 , n46581 , n46583 );
buf ( n46585 , n46584 );
not ( n46586 , n46585 );
or ( n46587 , n45947 , n46586 );
buf ( n46588 , n31040 );
not ( n46589 , n46588 );
nand ( n46590 , n46300 , n46589 );
nand ( n46591 , n46587 , n46590 );
buf ( n46592 , n46591 );
nor ( n46593 , n46578 , n46592 );
nor ( n46594 , n46576 , n46593 );
and ( n46595 , n46555 , n46594 );
not ( n46596 , n33249 );
buf ( n46597 , n46596 );
not ( n46598 , n46597 );
nand ( n46599 , n46307 , n46511 );
and ( n46600 , n46599 , n46513 );
not ( n46601 , n46599 );
not ( n46602 , n46513 );
and ( n46603 , n46601 , n46602 );
nor ( n46604 , n46600 , n46603 );
buf ( n46605 , n46604 );
not ( n46606 , n46605 );
or ( n46607 , n45991 , n46606 );
not ( n46608 , n29110 );
not ( n46609 , n46608 );
nand ( n46610 , n45941 , n46609 );
nand ( n46611 , n46607 , n46610 );
buf ( n46612 , n46611 );
not ( n46613 , n46612 );
not ( n46614 , n46613 );
or ( n46615 , n46598 , n46614 );
nor ( n46616 , n46312 , n46513 );
nand ( n46617 , n46307 , n46616 );
and ( n46618 , n46617 , n46512 );
not ( n46619 , n46617 );
and ( n46620 , n46619 , n46327 );
nor ( n46621 , n46618 , n46620 );
buf ( n46622 , n46621 );
not ( n46623 , n46622 );
or ( n46624 , n45941 , n46623 );
not ( n46625 , n38565 );
not ( n46626 , n46625 );
not ( n46627 , n46626 );
nand ( n46628 , n46300 , n46627 );
nand ( n46629 , n46624 , n46628 );
buf ( n46630 , n46629 );
not ( n46631 , n46630 );
buf ( n46632 , n33120 );
nand ( n46633 , n46631 , n46632 );
nand ( n46634 , n46615 , n46633 );
buf ( n46635 , n33837 );
not ( n46636 , n46635 );
buf ( n46637 , n46311 );
not ( n46638 , n46637 );
not ( n46639 , n46306 );
or ( n46640 , n46638 , n46639 );
or ( n46641 , n46306 , n46637 );
nand ( n46642 , n46640 , n46641 );
buf ( n46643 , n46642 );
not ( n46644 , n46643 );
or ( n46645 , n45976 , n46644 );
buf ( n46646 , n23930 );
buf ( n46647 , n46646 );
nand ( n46648 , n45947 , n46647 );
nand ( n46649 , n46645 , n46648 );
buf ( n46650 , n46649 );
not ( n46651 , n46650 );
not ( n46652 , n46651 );
or ( n46653 , n46636 , n46652 );
nand ( n46654 , n46307 , n46637 );
buf ( n46655 , n46309 );
not ( n46656 , n46655 );
xor ( n46657 , n46654 , n46656 );
buf ( n46658 , n46657 );
not ( n46659 , n46658 );
or ( n46660 , n46229 , n46659 );
buf ( n46661 , n33255 );
not ( n46662 , n46661 );
nand ( n46663 , n45941 , n46662 );
nand ( n46664 , n46660 , n46663 );
buf ( n46665 , n46664 );
not ( n46666 , n46665 );
buf ( n46667 , n24325 );
nand ( n46668 , n46666 , n46667 );
nand ( n46669 , n46653 , n46668 );
nor ( n46670 , n46634 , n46669 );
nand ( n46671 , n46595 , n46670 );
nor ( n46672 , n46504 , n46671 );
and ( n46673 , n46296 , n46672 );
not ( n46674 , n46667 );
nand ( n46675 , n46674 , n46665 );
not ( n46676 , n46675 );
not ( n46677 , n46635 );
nand ( n46678 , n46677 , n46650 );
not ( n46679 , n46678 );
or ( n46680 , n46676 , n46679 );
nand ( n46681 , n46680 , n46668 );
or ( n46682 , n46634 , n46681 );
not ( n46683 , n46632 );
nor ( n46684 , n46630 , n46683 );
not ( n46685 , n46597 );
nand ( n46686 , n46685 , n46612 );
or ( n46687 , n46684 , n46686 );
nand ( n46688 , n46630 , n46683 );
nand ( n46689 , n46687 , n46688 );
not ( n46690 , n46689 );
nand ( n46691 , n46682 , n46690 );
and ( n46692 , n46595 , n46691 );
not ( n46693 , n46555 );
not ( n46694 , n46577 );
nand ( n46695 , n46694 , n46592 );
or ( n46696 , n46576 , n46695 );
nand ( n46697 , n46573 , n46575 );
nand ( n46698 , n46696 , n46697 );
not ( n46699 , n46698 );
or ( n46700 , n46693 , n46699 );
not ( n46701 , n46533 );
not ( n46702 , n46534 );
nand ( n46703 , n46702 , n46553 );
not ( n46704 , n46703 );
and ( n46705 , n46701 , n46704 );
and ( n46706 , n46530 , n46532 );
nor ( n46707 , n46705 , n46706 );
nand ( n46708 , n46700 , n46707 );
nor ( n46709 , n46692 , n46708 );
or ( n46710 , n46709 , n46504 );
not ( n46711 , n46464 );
not ( n46712 , n46499 );
nand ( n46713 , n46712 , n46498 );
or ( n46714 , n46713 , n46484 );
nand ( n46715 , n46481 , n46483 );
nand ( n46716 , n46714 , n46715 );
not ( n46717 , n46716 );
or ( n46718 , n46711 , n46717 );
not ( n46719 , n46448 );
nand ( n46720 , n46460 , n46462 );
not ( n46721 , n46720 );
and ( n46722 , n46719 , n46721 );
and ( n46723 , n46445 , n46447 );
nor ( n46724 , n46722 , n46723 );
nand ( n46725 , n46718 , n46724 );
and ( n46726 , n46725 , n46427 );
not ( n46727 , n46354 );
nor ( n46728 , n46727 , n46297 );
and ( n46729 , n46377 , n46728 );
not ( n46730 , n46374 );
nor ( n46731 , n46730 , n46376 );
nor ( n46732 , n46729 , n46731 );
or ( n46733 , n46732 , n46426 );
not ( n46734 , n46397 );
nor ( n46735 , n46734 , n46379 );
and ( n46736 , n46735 , n46425 );
nor ( n46737 , n46422 , n46424 );
nor ( n46738 , n46736 , n46737 );
nand ( n46739 , n46733 , n46738 );
nor ( n46740 , n46726 , n46739 );
nand ( n46741 , n46710 , n46740 );
nor ( n46742 , n46673 , n46741 );
buf ( n46743 , n46742 );
not ( n46744 , n46743 );
not ( n46745 , n19212 );
nand ( n46746 , n46745 , n19206 , n19140 );
not ( n46747 , n46746 );
and ( n46748 , n46744 , n46747 );
and ( n46749 , n19206 , n19140 , n19212 );
and ( n46750 , n46743 , n46749 );
nor ( n46751 , n46748 , n46750 );
nand ( n46752 , n19380 , n19639 );
or ( n46753 , n46751 , n46752 );
or ( n46754 , n19195 , n19146 );
nor ( n46755 , n46754 , n46746 );
and ( n46756 , n46743 , n46755 );
not ( n46757 , n46754 );
not ( n46758 , n46749 );
not ( n46759 , n46758 );
and ( n46760 , n46757 , n46759 );
buf ( n46761 , n41032 );
not ( n46762 , n46761 );
buf ( n46763 , n29820 );
nor ( n46764 , n46762 , n46763 );
buf ( n46765 , n29856 );
buf ( n46766 , n30176 );
not ( n46767 , n46766 );
nor ( n46768 , n46765 , n46767 );
nor ( n46769 , n46764 , n46768 );
not ( n46770 , n46769 );
buf ( n46771 , n34244 );
not ( n46772 , n46771 );
buf ( n46773 , n34152 );
not ( n46774 , n46773 );
not ( n46775 , n46774 );
or ( n46776 , n46772 , n46775 );
buf ( n46777 , n34158 );
buf ( n46778 , n34241 );
not ( n46779 , n46778 );
nand ( n46780 , n46777 , n46779 );
nand ( n46781 , n46776 , n46780 );
nor ( n46782 , n46770 , n46781 );
buf ( n46783 , n38123 );
not ( n46784 , n46783 );
buf ( n46785 , n29795 );
nor ( n46786 , n46784 , n46785 );
buf ( n46787 , n30019 );
not ( n46788 , n46787 );
buf ( n46789 , n27810 );
nor ( n46790 , n46788 , n46789 );
nor ( n46791 , n46786 , n46790 );
buf ( n46792 , n27885 );
not ( n46793 , n46792 );
buf ( n46794 , n27832 );
nor ( n46795 , n46793 , n46794 );
buf ( n46796 , n27932 );
not ( n46797 , n46796 );
buf ( n46798 , n27783 );
nor ( n46799 , n46797 , n46798 );
nor ( n46800 , n46795 , n46799 );
and ( n46801 , n46791 , n46800 );
nand ( n46802 , n46782 , n46801 );
buf ( n46803 , n24324 );
not ( n46804 , n46803 );
not ( n46805 , n46661 );
buf ( n46806 , n46805 );
nand ( n46807 , n46804 , n46806 );
buf ( n46808 , n33836 );
not ( n46809 , n46808 );
buf ( n46810 , n46646 );
nand ( n46811 , n46809 , n46810 );
and ( n46812 , n46807 , n46811 );
not ( n46813 , n46803 );
nor ( n46814 , n46813 , n46806 );
nor ( n46815 , n46812 , n46814 );
not ( n46816 , n46815 );
buf ( n46817 , n33119 );
not ( n46818 , n46817 );
buf ( n46819 , n46625 );
nor ( n46820 , n46818 , n46819 );
buf ( n46821 , n33248 );
not ( n46822 , n46821 );
not ( n46823 , n46608 );
buf ( n46824 , n46823 );
nor ( n46825 , n46822 , n46824 );
nor ( n46826 , n46820 , n46825 );
not ( n46827 , n46826 );
or ( n46828 , n46816 , n46827 );
not ( n46829 , n46820 );
not ( n46830 , n46824 );
nor ( n46831 , n46830 , n46821 );
and ( n46832 , n46829 , n46831 );
not ( n46833 , n46819 );
nor ( n46834 , n46833 , n46817 );
nor ( n46835 , n46832 , n46834 );
nand ( n46836 , n46828 , n46835 );
buf ( n46837 , n40408 );
not ( n46838 , n46837 );
not ( n46839 , n46505 );
buf ( n46840 , n46839 );
nor ( n46841 , n46838 , n46840 );
buf ( n46842 , n27049 );
not ( n46843 , n46842 );
buf ( n46844 , n46536 );
nor ( n46845 , n46843 , n46844 );
nor ( n46846 , n46841 , n46845 );
buf ( n46847 , n31097 );
not ( n46848 , n46847 );
buf ( n46849 , n46556 );
nor ( n46850 , n46848 , n46849 );
buf ( n46851 , n38737 );
not ( n46852 , n46851 );
not ( n46853 , n46588 );
buf ( n46854 , n46853 );
nor ( n46855 , n46852 , n46854 );
nor ( n46856 , n46850 , n46855 );
nand ( n46857 , n46846 , n46856 );
not ( n46858 , n46857 );
and ( n46859 , n46836 , n46858 );
not ( n46860 , n46846 );
not ( n46861 , n46851 );
nand ( n46862 , n46861 , n46854 );
or ( n46863 , n46850 , n46862 );
not ( n46864 , n46849 );
or ( n46865 , n46864 , n46847 );
nand ( n46866 , n46863 , n46865 );
not ( n46867 , n46866 );
or ( n46868 , n46860 , n46867 );
not ( n46869 , n46841 );
not ( n46870 , n46844 );
nor ( n46871 , n46870 , n46842 );
and ( n46872 , n46869 , n46871 );
not ( n46873 , n46840 );
nor ( n46874 , n46873 , n46837 );
nor ( n46875 , n46872 , n46874 );
nand ( n46876 , n46868 , n46875 );
nor ( n46877 , n46859 , n46876 );
or ( n46878 , n46802 , n46877 );
not ( n46879 , n46792 );
nand ( n46880 , n46879 , n46794 );
not ( n46881 , n46796 );
nand ( n46882 , n46881 , n46798 );
and ( n46883 , n46880 , n46882 );
nor ( n46884 , n46883 , n46795 );
not ( n46885 , n46884 );
not ( n46886 , n46791 );
or ( n46887 , n46885 , n46886 );
not ( n46888 , n46786 );
not ( n46889 , n46789 );
nor ( n46890 , n46889 , n46787 );
and ( n46891 , n46888 , n46890 );
not ( n46892 , n46785 );
nor ( n46893 , n46892 , n46783 );
nor ( n46894 , n46891 , n46893 );
nand ( n46895 , n46887 , n46894 );
and ( n46896 , n46782 , n46895 );
not ( n46897 , n46764 );
not ( n46898 , n46765 );
nor ( n46899 , n46898 , n46766 );
and ( n46900 , n46897 , n46899 );
not ( n46901 , n46763 );
nor ( n46902 , n46901 , n46761 );
nor ( n46903 , n46900 , n46902 );
or ( n46904 , n46781 , n46903 );
not ( n46905 , n46773 );
nor ( n46906 , n46905 , n46771 );
and ( n46907 , n46780 , n46906 );
nor ( n46908 , n46777 , n46779 );
nor ( n46909 , n46907 , n46908 );
nand ( n46910 , n46904 , n46909 );
nor ( n46911 , n46896 , n46910 );
nand ( n46912 , n46878 , n46911 );
buf ( n46913 , n33794 );
buf ( n46914 , n37640 );
not ( n46915 , n46914 );
nor ( n46916 , n46913 , n46915 );
buf ( n46917 , n21622 );
not ( n46918 , n46917 );
buf ( n46919 , n35964 );
nor ( n46920 , n46918 , n46919 );
nor ( n46921 , n46916 , n46920 );
buf ( n46922 , n46159 );
buf ( n46923 , n29547 );
not ( n46924 , n46923 );
nor ( n46925 , n46922 , n46924 );
buf ( n46926 , n29458 );
not ( n46927 , n46926 );
buf ( n46928 , n46176 );
nor ( n46929 , n46927 , n46928 );
nor ( n46930 , n46925 , n46929 );
and ( n46931 , n46921 , n46930 );
buf ( n46932 , n39293 );
not ( n46933 , n46932 );
not ( n46934 , n46194 );
buf ( n46935 , n46934 );
nor ( n46936 , n46933 , n46935 );
buf ( n46937 , n20565 );
not ( n46938 , n46937 );
buf ( n46939 , n39236 );
nor ( n46940 , n46938 , n46939 );
nor ( n46941 , n46936 , n46940 );
not ( n46942 , n46941 );
buf ( n46943 , n35712 );
not ( n46944 , n46943 );
buf ( n46945 , n46247 );
not ( n46946 , n46945 );
not ( n46947 , n46946 );
or ( n46948 , n46944 , n46947 );
buf ( n46949 , n46224 );
buf ( n46950 , n35836 );
not ( n46951 , n46950 );
nor ( n46952 , n46949 , n46951 );
not ( n46953 , n46952 );
nand ( n46954 , n46948 , n46953 );
nor ( n46955 , n46942 , n46954 );
buf ( n46956 , n22869 );
not ( n46957 , n46956 );
buf ( n46958 , n45936 );
nor ( n46959 , n46957 , n46958 );
buf ( n46960 , n35187 );
not ( n46961 , n46960 );
buf ( n46962 , n45982 );
nor ( n46963 , n46961 , n46962 );
nor ( n46964 , n46959 , n46963 );
buf ( n46965 , n46003 );
buf ( n46966 , n24441 );
not ( n46967 , n46966 );
nor ( n46968 , n46965 , n46967 );
buf ( n46969 , n30627 );
not ( n46970 , n46969 );
buf ( n46971 , n46019 );
nor ( n46972 , n46970 , n46971 );
nor ( n46973 , n46968 , n46972 );
buf ( n46974 , n46037 );
not ( n46975 , n46974 );
buf ( n46976 , n34028 );
nand ( n46977 , n46975 , n46976 );
buf ( n46978 , n24644 );
not ( n46979 , n46978 );
buf ( n46980 , n18309 );
nor ( n46981 , n46979 , n46980 );
buf ( n46982 , n19284 );
not ( n46983 , n46982 );
buf ( n46984 , n19092 );
nor ( n46985 , n46983 , n46984 );
or ( n46986 , n46981 , n46985 );
not ( n46987 , n46984 );
or ( n46988 , n46987 , n46982 );
nand ( n46989 , n46986 , n46988 );
buf ( n46990 , n46056 );
not ( n46991 , n46990 );
buf ( n46992 , n21021 );
nand ( n46993 , n46991 , n46992 );
nand ( n46994 , n46977 , n46989 , n46993 );
not ( n46995 , n46990 );
nor ( n46996 , n46995 , n46992 );
nand ( n46997 , n46977 , n46996 );
not ( n46998 , n46976 );
nand ( n46999 , n46998 , n46974 );
nand ( n47000 , n46994 , n46997 , n46999 );
nand ( n47001 , n46964 , n46973 , n47000 );
not ( n47002 , n46969 );
nand ( n47003 , n47002 , n46971 );
or ( n47004 , n46968 , n47003 );
nand ( n47005 , n46965 , n46967 );
nand ( n47006 , n47004 , n47005 );
nand ( n47007 , n46964 , n47006 );
not ( n47008 , n46959 );
not ( n47009 , n46962 );
nor ( n47010 , n47009 , n46960 );
and ( n47011 , n47008 , n47010 );
not ( n47012 , n46958 );
nor ( n47013 , n47012 , n46956 );
nor ( n47014 , n47011 , n47013 );
nand ( n47015 , n47001 , n47007 , n47014 );
nand ( n47016 , n46931 , n46955 , n47015 );
not ( n47017 , n46941 );
not ( n47018 , n46943 );
nand ( n47019 , n47018 , n46945 );
or ( n47020 , n46952 , n47019 );
not ( n47021 , n46949 );
or ( n47022 , n47021 , n46950 );
nand ( n47023 , n47020 , n47022 );
not ( n47024 , n47023 );
or ( n47025 , n47017 , n47024 );
not ( n47026 , n46936 );
not ( n47027 , n46939 );
nor ( n47028 , n47027 , n46937 );
and ( n47029 , n47026 , n47028 );
not ( n47030 , n46935 );
nor ( n47031 , n47030 , n46932 );
nor ( n47032 , n47029 , n47031 );
nand ( n47033 , n47025 , n47032 );
nand ( n47034 , n47033 , n46931 );
not ( n47035 , n46926 );
nand ( n47036 , n47035 , n46928 );
or ( n47037 , n46925 , n47036 );
nand ( n47038 , n46922 , n46924 );
nand ( n47039 , n47037 , n47038 );
and ( n47040 , n47039 , n46921 );
not ( n47041 , n46917 );
nand ( n47042 , n47041 , n46919 );
or ( n47043 , n46916 , n47042 );
nand ( n47044 , n46913 , n46915 );
nand ( n47045 , n47043 , n47044 );
nor ( n47046 , n47040 , n47045 );
nand ( n47047 , n47016 , n47034 , n47046 );
not ( n47048 , n46808 );
nor ( n47049 , n47048 , n46810 );
nor ( n47050 , n46814 , n47049 );
nand ( n47051 , n46826 , n47050 );
nor ( n47052 , n46857 , n47051 );
and ( n47053 , n47047 , n46782 , n47052 , n46801 );
nor ( n47054 , n46912 , n47053 );
buf ( n47055 , n47054 );
nor ( n47056 , n19315 , n19141 );
not ( n47057 , n47056 );
or ( n47058 , n47055 , n47057 );
nor ( n47059 , n19213 , n19141 );
nand ( n47060 , n47055 , n47059 );
buf ( n47061 , n29967 );
not ( n47062 , n47061 );
buf ( n47063 , n29964 );
nor ( n47064 , n47062 , n47063 );
not ( n47065 , n47064 );
buf ( n47066 , n34247 );
not ( n47067 , n47066 );
buf ( n47068 , n40951 );
not ( n47069 , n47068 );
not ( n47070 , n47069 );
or ( n47071 , n47067 , n47070 );
not ( n47072 , n47066 );
nand ( n47073 , n47072 , n47068 );
nand ( n47074 , n47071 , n47073 );
not ( n47075 , n47074 );
or ( n47076 , n47065 , n47075 );
or ( n47077 , n47074 , n47064 );
nand ( n47078 , n47076 , n47077 );
buf ( n47079 , n19668 );
not ( n47080 , n47079 );
buf ( n47081 , n20564 );
nor ( n47082 , n47080 , n47081 );
not ( n47083 , n47082 );
buf ( n47084 , n21601 );
not ( n47085 , n47084 );
buf ( n47086 , n21366 );
nand ( n47087 , n47085 , n47086 );
not ( n47088 , n47086 );
nand ( n47089 , n47088 , n47084 );
nand ( n47090 , n47087 , n47089 );
not ( n47091 , n47090 );
or ( n47092 , n47083 , n47091 );
or ( n47093 , n47090 , n47082 );
nand ( n47094 , n47092 , n47093 );
buf ( n47095 , n20428 );
not ( n47096 , n47095 );
buf ( n47097 , n20531 );
nor ( n47098 , n47096 , n47097 );
not ( n47099 , n47098 );
buf ( n47100 , n35186 );
not ( n47101 , n47100 );
buf ( n47102 , n20207 );
nand ( n47103 , n47101 , n47102 );
not ( n47104 , n47102 );
nand ( n47105 , n47104 , n47100 );
nand ( n47106 , n47103 , n47105 );
not ( n47107 , n47106 );
or ( n47108 , n47099 , n47107 );
or ( n47109 , n47106 , n47098 );
nand ( n47110 , n47108 , n47109 );
buf ( n47111 , n45956 );
buf ( n47112 , n45954 );
not ( n47113 , n47112 );
and ( n47114 , n47111 , n47113 );
not ( n47115 , n47111 );
and ( n47116 , n47115 , n47112 );
nor ( n47117 , n47114 , n47116 );
not ( n47118 , n47117 );
buf ( n47119 , n34027 );
not ( n47120 , n47119 );
and ( n47121 , n47118 , n47120 );
and ( n47122 , n47117 , n47119 );
nor ( n47123 , n47121 , n47122 );
buf ( n47124 , n24644 );
not ( n47125 , n47124 );
buf ( n47126 , n18309 );
not ( n47127 , n47126 );
or ( n47128 , n47125 , n47127 );
or ( n47129 , n47126 , n47124 );
nand ( n47130 , n47128 , n47129 );
buf ( n47131 , n21020 );
buf ( n47132 , n46056 );
xnor ( n47133 , n47131 , n47132 );
buf ( n47134 , n19285 );
buf ( n47135 , n19092 );
xnor ( n47136 , n47134 , n47135 );
and ( n47137 , n47123 , n47130 , n47133 , n47136 );
nand ( n47138 , n47078 , n47094 , n47110 , n47137 );
nor ( n47139 , n47113 , n47119 );
not ( n47140 , n47139 );
buf ( n47141 , n20114 );
not ( n47142 , n47141 );
buf ( n47143 , n30626 );
nor ( n47144 , n47142 , n47143 );
not ( n47145 , n47143 );
nor ( n47146 , n47145 , n47141 );
or ( n47147 , n47144 , n47146 );
not ( n47148 , n47147 );
or ( n47149 , n47140 , n47148 );
or ( n47150 , n47147 , n47139 );
nand ( n47151 , n47149 , n47150 );
not ( n47152 , n47144 );
not ( n47153 , n47097 );
nor ( n47154 , n47153 , n47095 );
or ( n47155 , n47098 , n47154 );
not ( n47156 , n47155 );
or ( n47157 , n47152 , n47156 );
or ( n47158 , n47155 , n47144 );
nand ( n47159 , n47157 , n47158 );
buf ( n47160 , n46093 );
not ( n47161 , n47160 );
buf ( n47162 , n35711 );
nor ( n47163 , n47161 , n47162 );
not ( n47164 , n47163 );
buf ( n47165 , n19937 );
buf ( n47166 , n47165 );
not ( n47167 , n47166 );
buf ( n47168 , n35835 );
nor ( n47169 , n47167 , n47168 );
not ( n47170 , n47168 );
nor ( n47171 , n47170 , n47166 );
or ( n47172 , n47169 , n47171 );
not ( n47173 , n47172 );
or ( n47174 , n47164 , n47173 );
or ( n47175 , n47172 , n47163 );
nand ( n47176 , n47174 , n47175 );
not ( n47177 , n47073 );
not ( n47178 , n47177 );
buf ( n47179 , n46384 );
not ( n47180 , n47179 );
buf ( n47181 , n34244 );
nor ( n47182 , n47180 , n47181 );
and ( n47183 , n47180 , n47181 );
or ( n47184 , n47182 , n47183 );
not ( n47185 , n47184 );
or ( n47186 , n47178 , n47185 );
or ( n47187 , n47184 , n47177 );
nand ( n47188 , n47186 , n47187 );
nand ( n47189 , n47151 , n47159 , n47176 , n47188 );
nor ( n47190 , n47138 , n47189 );
not ( n47191 , n47064 );
not ( n47192 , n47061 );
nand ( n47193 , n47192 , n47063 );
nand ( n47194 , n47191 , n47193 );
buf ( n47195 , n38122 );
not ( n47196 , n47195 );
buf ( n47197 , n30078 );
nand ( n47198 , n47196 , n47197 );
xnor ( n47199 , n47194 , n47198 );
not ( n47200 , n47162 );
nor ( n47201 , n47200 , n47160 );
or ( n47202 , n47163 , n47201 );
buf ( n47203 , n19992 );
not ( n47204 , n47203 );
buf ( n47205 , n22868 );
nor ( n47206 , n47204 , n47205 );
and ( n47207 , n47202 , n47206 );
nor ( n47208 , n47202 , n47206 );
nor ( n47209 , n47207 , n47208 );
not ( n47210 , n47205 );
nor ( n47211 , n47210 , n47203 );
or ( n47212 , n47206 , n47211 );
not ( n47213 , n47103 );
and ( n47214 , n47212 , n47213 );
nor ( n47215 , n47212 , n47213 );
nor ( n47216 , n47214 , n47215 );
nor ( n47217 , n47199 , n47209 , n47216 );
not ( n47218 , n47169 );
not ( n47219 , n47082 );
not ( n47220 , n47079 );
nand ( n47221 , n47220 , n47081 );
nand ( n47222 , n47219 , n47221 );
not ( n47223 , n47222 );
or ( n47224 , n47218 , n47223 );
or ( n47225 , n47222 , n47169 );
nand ( n47226 , n47224 , n47225 );
buf ( n47227 , n30019 );
not ( n47228 , n47227 );
buf ( n47229 , n46336 );
nand ( n47230 , n47228 , n47229 );
not ( n47231 , n47230 );
not ( n47232 , n47231 );
not ( n47233 , n47197 );
nand ( n47234 , n47233 , n47195 );
nand ( n47235 , n47198 , n47234 );
not ( n47236 , n47235 );
or ( n47237 , n47232 , n47236 );
or ( n47238 , n47235 , n47231 );
nand ( n47239 , n47237 , n47238 );
nand ( n47240 , n47190 , n47217 , n47226 , n47239 );
buf ( n47241 , n46321 );
buf ( n47242 , n27069 );
not ( n47243 , n47242 );
and ( n47244 , n47241 , n47243 );
not ( n47245 , n47242 );
nor ( n47246 , n47245 , n47241 );
or ( n47247 , n47244 , n47246 );
not ( n47248 , n47247 );
buf ( n47249 , n33118 );
not ( n47250 , n47249 );
buf ( n47251 , n46326 );
nand ( n47252 , n47250 , n47251 );
not ( n47253 , n47252 );
and ( n47254 , n47248 , n47253 );
and ( n47255 , n47247 , n47252 );
nor ( n47256 , n47254 , n47255 );
buf ( n47257 , n46315 );
not ( n47258 , n47257 );
buf ( n47259 , n27066 );
nor ( n47260 , n47258 , n47259 );
not ( n47261 , n47260 );
buf ( n47262 , n46324 );
buf ( n47263 , n27048 );
not ( n47264 , n47263 );
and ( n47265 , n47262 , n47264 );
nor ( n47266 , n47262 , n47264 );
or ( n47267 , n47265 , n47266 );
not ( n47268 , n47267 );
or ( n47269 , n47261 , n47268 );
or ( n47270 , n47267 , n47260 );
nand ( n47271 , n47269 , n47270 );
buf ( n47272 , n46099 );
not ( n47273 , n47272 );
buf ( n47274 , n29546 );
nor ( n47275 , n47273 , n47274 );
not ( n47276 , n47275 );
buf ( n47277 , n46104 );
not ( n47278 , n47277 );
buf ( n47279 , n21621 );
nor ( n47280 , n47278 , n47279 );
not ( n47281 , n47279 );
nor ( n47282 , n47281 , n47277 );
or ( n47283 , n47280 , n47282 );
not ( n47284 , n47283 );
or ( n47285 , n47276 , n47284 );
or ( n47286 , n47283 , n47275 );
nand ( n47287 , n47285 , n47286 );
not ( n47288 , n47280 );
buf ( n47289 , n46109 );
not ( n47290 , n47289 );
buf ( n47291 , n37639 );
nor ( n47292 , n47290 , n47291 );
not ( n47293 , n47291 );
nor ( n47294 , n47293 , n47289 );
or ( n47295 , n47292 , n47294 );
not ( n47296 , n47295 );
or ( n47297 , n47288 , n47296 );
or ( n47298 , n47295 , n47280 );
nand ( n47299 , n47297 , n47298 );
nand ( n47300 , n47256 , n47271 , n47287 , n47299 );
buf ( n47301 , n27058 );
not ( n47302 , n47301 );
buf ( n47303 , n46319 );
nand ( n47304 , n47302 , n47303 );
not ( n47305 , n47304 );
not ( n47306 , n47305 );
not ( n47307 , n47251 );
nand ( n47308 , n47307 , n47249 );
nand ( n47309 , n47252 , n47308 );
not ( n47310 , n47309 );
or ( n47311 , n47306 , n47310 );
or ( n47312 , n47309 , n47305 );
nand ( n47313 , n47311 , n47312 );
buf ( n47314 , n27932 );
not ( n47315 , n47314 );
buf ( n47316 , n46331 );
nand ( n47317 , n47315 , n47316 );
not ( n47318 , n47317 );
not ( n47319 , n47318 );
buf ( n47320 , n27885 );
not ( n47321 , n47320 );
buf ( n47322 , n46333 );
nand ( n47323 , n47321 , n47322 );
not ( n47324 , n47322 );
nand ( n47325 , n47324 , n47320 );
nand ( n47326 , n47323 , n47325 );
not ( n47327 , n47326 );
or ( n47328 , n47319 , n47327 );
or ( n47329 , n47326 , n47318 );
nand ( n47330 , n47328 , n47329 );
buf ( n47331 , n46313 );
buf ( n47332 , n28129 );
not ( n47333 , n47332 );
and ( n47334 , n47331 , n47333 );
not ( n47335 , n47334 );
not ( n47336 , n47316 );
nand ( n47337 , n47336 , n47314 );
nand ( n47338 , n47317 , n47337 );
not ( n47339 , n47338 );
or ( n47340 , n47335 , n47339 );
or ( n47341 , n47338 , n47334 );
nand ( n47342 , n47340 , n47341 );
not ( n47343 , n47323 );
not ( n47344 , n47343 );
not ( n47345 , n47229 );
nand ( n47346 , n47345 , n47227 );
nand ( n47347 , n47230 , n47346 );
not ( n47348 , n47347 );
or ( n47349 , n47344 , n47348 );
or ( n47350 , n47347 , n47343 );
nand ( n47351 , n47349 , n47350 );
nand ( n47352 , n47313 , n47330 , n47342 , n47351 );
nor ( n47353 , n47300 , n47352 );
not ( n47354 , n47244 );
not ( n47355 , n47259 );
nor ( n47356 , n47355 , n47257 );
or ( n47357 , n47260 , n47356 );
not ( n47358 , n47357 );
or ( n47359 , n47354 , n47358 );
or ( n47360 , n47357 , n47244 );
nand ( n47361 , n47359 , n47360 );
not ( n47362 , n47265 );
nor ( n47363 , n47331 , n47333 );
or ( n47364 , n47334 , n47363 );
not ( n47365 , n47364 );
or ( n47366 , n47362 , n47365 );
or ( n47367 , n47364 , n47265 );
nand ( n47368 , n47366 , n47367 );
buf ( n47369 , n24323 );
not ( n47370 , n47369 );
buf ( n47371 , n46308 );
nand ( n47372 , n47370 , n47371 );
not ( n47373 , n47372 );
not ( n47374 , n47373 );
not ( n47375 , n47303 );
nand ( n47376 , n47375 , n47301 );
nand ( n47377 , n47304 , n47376 );
not ( n47378 , n47377 );
or ( n47379 , n47374 , n47378 );
or ( n47380 , n47377 , n47373 );
nand ( n47381 , n47379 , n47380 );
not ( n47382 , n47292 );
buf ( n47383 , n33835 );
not ( n47384 , n47383 );
buf ( n47385 , n46310 );
nand ( n47386 , n47384 , n47385 );
not ( n47387 , n47385 );
nand ( n47388 , n47387 , n47383 );
nand ( n47389 , n47386 , n47388 );
not ( n47390 , n47389 );
or ( n47391 , n47382 , n47390 );
or ( n47392 , n47389 , n47292 );
nand ( n47393 , n47391 , n47392 );
nand ( n47394 , n47361 , n47368 , n47381 , n47393 );
not ( n47395 , n47087 );
not ( n47396 , n47395 );
buf ( n47397 , n46101 );
not ( n47398 , n47397 );
buf ( n47399 , n29457 );
nor ( n47400 , n47398 , n47399 );
not ( n47401 , n47399 );
nor ( n47402 , n47401 , n47397 );
or ( n47403 , n47400 , n47402 );
not ( n47404 , n47403 );
or ( n47405 , n47396 , n47404 );
or ( n47406 , n47403 , n47395 );
nand ( n47407 , n47405 , n47406 );
not ( n47408 , n47400 );
not ( n47409 , n47274 );
nor ( n47410 , n47409 , n47272 );
or ( n47411 , n47275 , n47410 );
not ( n47412 , n47411 );
or ( n47413 , n47408 , n47412 );
or ( n47414 , n47411 , n47400 );
nand ( n47415 , n47413 , n47414 );
not ( n47416 , n47386 );
not ( n47417 , n47416 );
not ( n47418 , n47371 );
nand ( n47419 , n47418 , n47369 );
nand ( n47420 , n47372 , n47419 );
not ( n47421 , n47420 );
or ( n47422 , n47417 , n47421 );
or ( n47423 , n47420 , n47416 );
nand ( n47424 , n47422 , n47423 );
not ( n47425 , n47182 );
buf ( n47426 , n46401 );
buf ( n47427 , n34241 );
xor ( n47428 , n47426 , n47427 );
not ( n47429 , n47428 );
or ( n47430 , n47425 , n47429 );
or ( n47431 , n47428 , n47182 );
nand ( n47432 , n47430 , n47431 );
nand ( n47433 , n47407 , n47415 , n47424 , n47432 );
nor ( n47434 , n47394 , n47433 );
nand ( n47435 , n47353 , n47434 );
nor ( n47436 , n47240 , n47435 );
buf ( n47437 , n47436 );
nand ( n47438 , n47437 , n46749 );
nand ( n47439 , n47058 , n47060 , n47438 );
nor ( n47440 , n19380 , n30179 );
and ( n47441 , n47439 , n47440 );
nor ( n47442 , n46760 , n47441 );
buf ( n47443 , n21623 );
not ( n47444 , n47443 );
not ( n47445 , n47444 );
buf ( n47446 , n46139 );
not ( n47447 , n47446 );
or ( n47448 , n47445 , n47447 );
buf ( n47449 , n46119 );
buf ( n47450 , n37640 );
not ( n47451 , n47450 );
nand ( n47452 , n47449 , n47451 );
nand ( n47453 , n47448 , n47452 );
buf ( n47454 , n29458 );
not ( n47455 , n47454 );
not ( n47456 , n47455 );
buf ( n47457 , n46176 );
not ( n47458 , n47457 );
or ( n47459 , n47456 , n47458 );
buf ( n47460 , n46159 );
buf ( n47461 , n29547 );
not ( n47462 , n47461 );
nand ( n47463 , n47460 , n47462 );
nand ( n47464 , n47459 , n47463 );
nor ( n47465 , n47453 , n47464 );
buf ( n47466 , n35836 );
not ( n47467 , n47466 );
buf ( n47468 , n46224 );
nand ( n47469 , n47467 , n47468 );
buf ( n47470 , n46247 );
buf ( n47471 , n35713 );
not ( n47472 , n47471 );
nor ( n47473 , n47470 , n47472 );
and ( n47474 , n47469 , n47473 );
not ( n47475 , n47466 );
nor ( n47476 , n47475 , n47468 );
nor ( n47477 , n47474 , n47476 );
buf ( n47478 , n20565 );
not ( n47479 , n47478 );
not ( n47480 , n47479 );
buf ( n47481 , n46203 );
not ( n47482 , n47481 );
or ( n47483 , n47480 , n47482 );
buf ( n47484 , n39293 );
not ( n47485 , n47484 );
buf ( n47486 , n46195 );
nand ( n47487 , n47485 , n47486 );
nand ( n47488 , n47483 , n47487 );
or ( n47489 , n47477 , n47488 );
nor ( n47490 , n47481 , n47479 );
and ( n47491 , n47487 , n47490 );
not ( n47492 , n47484 );
nor ( n47493 , n47492 , n47486 );
nor ( n47494 , n47491 , n47493 );
nand ( n47495 , n47489 , n47494 );
and ( n47496 , n47465 , n47495 );
nor ( n47497 , n47457 , n47455 );
and ( n47498 , n47463 , n47497 );
nor ( n47499 , n47460 , n47462 );
nor ( n47500 , n47498 , n47499 );
or ( n47501 , n47500 , n47453 );
nor ( n47502 , n47446 , n47444 );
and ( n47503 , n47452 , n47502 );
nor ( n47504 , n47449 , n47451 );
nor ( n47505 , n47503 , n47504 );
nand ( n47506 , n47501 , n47505 );
nor ( n47507 , n47496 , n47506 );
not ( n47508 , n47472 );
not ( n47509 , n47470 );
or ( n47510 , n47508 , n47509 );
nand ( n47511 , n47510 , n47469 );
nor ( n47512 , n47488 , n47511 );
buf ( n47513 , n22870 );
not ( n47514 , n47513 );
buf ( n47515 , n45936 );
nand ( n47516 , n47514 , n47515 );
buf ( n47517 , n35187 );
not ( n47518 , n47517 );
buf ( n47519 , n45982 );
nand ( n47520 , n47518 , n47519 );
and ( n47521 , n47516 , n47520 );
not ( n47522 , n47521 );
buf ( n47523 , n34028 );
not ( n47524 , n47523 );
buf ( n47525 , n46037 );
nand ( n47526 , n47524 , n47525 );
buf ( n47527 , n18309 );
not ( n47528 , n47527 );
buf ( n47529 , n24644 );
nor ( n47530 , n47528 , n47529 );
buf ( n47531 , n19092 );
buf ( n47532 , n19284 );
not ( n47533 , n47532 );
and ( n47534 , n47531 , n47533 );
or ( n47535 , n47530 , n47534 );
or ( n47536 , n47531 , n47533 );
nand ( n47537 , n47535 , n47536 );
buf ( n47538 , n21020 );
not ( n47539 , n47538 );
buf ( n47540 , n46056 );
nand ( n47541 , n47539 , n47540 );
and ( n47542 , n47526 , n47537 , n47541 );
not ( n47543 , n47538 );
nor ( n47544 , n47543 , n47540 );
not ( n47545 , n47544 );
not ( n47546 , n47526 );
or ( n47547 , n47545 , n47546 );
not ( n47548 , n47525 );
nand ( n47549 , n47548 , n47523 );
nand ( n47550 , n47547 , n47549 );
nor ( n47551 , n47542 , n47550 );
buf ( n47552 , n30627 );
not ( n47553 , n47552 );
not ( n47554 , n47553 );
buf ( n47555 , n46019 );
not ( n47556 , n47555 );
or ( n47557 , n47554 , n47556 );
buf ( n47558 , n24441 );
not ( n47559 , n47558 );
buf ( n47560 , n46003 );
nand ( n47561 , n47559 , n47560 );
nand ( n47562 , n47557 , n47561 );
nor ( n47563 , n47551 , n47562 );
not ( n47564 , n47563 );
or ( n47565 , n47522 , n47564 );
nor ( n47566 , n47555 , n47553 );
not ( n47567 , n47566 );
not ( n47568 , n47561 );
or ( n47569 , n47567 , n47568 );
not ( n47570 , n47560 );
nand ( n47571 , n47570 , n47558 );
nand ( n47572 , n47569 , n47571 );
and ( n47573 , n47521 , n47572 );
not ( n47574 , n47517 );
nor ( n47575 , n47574 , n47519 );
not ( n47576 , n47575 );
not ( n47577 , n47516 );
or ( n47578 , n47576 , n47577 );
not ( n47579 , n47515 );
nand ( n47580 , n47579 , n47513 );
nand ( n47581 , n47578 , n47580 );
nor ( n47582 , n47573 , n47581 );
nand ( n47583 , n47565 , n47582 );
nand ( n47584 , n47465 , n47512 , n47583 );
nand ( n47585 , n47507 , n47584 );
buf ( n47586 , n27049 );
not ( n47587 , n47586 );
not ( n47588 , n47587 );
buf ( n47589 , n46536 );
not ( n47590 , n47589 );
or ( n47591 , n47588 , n47590 );
buf ( n47592 , n40408 );
not ( n47593 , n47592 );
buf ( n47594 , n46506 );
nand ( n47595 , n47593 , n47594 );
nand ( n47596 , n47591 , n47595 );
buf ( n47597 , n38738 );
not ( n47598 , n47597 );
not ( n47599 , n47598 );
buf ( n47600 , n46589 );
not ( n47601 , n47600 );
or ( n47602 , n47599 , n47601 );
buf ( n47603 , n46557 );
buf ( n47604 , n31097 );
not ( n47605 , n47604 );
nand ( n47606 , n47603 , n47605 );
nand ( n47607 , n47602 , n47606 );
nor ( n47608 , n47596 , n47607 );
not ( n47609 , n47608 );
buf ( n47610 , n33248 );
not ( n47611 , n47610 );
not ( n47612 , n47611 );
buf ( n47613 , n46609 );
not ( n47614 , n47613 );
or ( n47615 , n47612 , n47614 );
not ( n47616 , n46626 );
buf ( n47617 , n47616 );
buf ( n47618 , n33119 );
not ( n47619 , n47618 );
nand ( n47620 , n47617 , n47619 );
nand ( n47621 , n47615 , n47620 );
not ( n47622 , n47621 );
buf ( n47623 , n46662 );
buf ( n47624 , n24324 );
not ( n47625 , n47624 );
nand ( n47626 , n47623 , n47625 );
buf ( n47627 , n46646 );
buf ( n47628 , n33836 );
not ( n47629 , n47628 );
nand ( n47630 , n47627 , n47629 );
and ( n47631 , n47626 , n47630 );
nand ( n47632 , n47622 , n47631 );
nor ( n47633 , n47609 , n47632 );
buf ( n47634 , n34244 );
not ( n47635 , n47634 );
not ( n47636 , n47635 );
not ( n47637 , n34153 );
buf ( n47638 , n47637 );
not ( n47639 , n47638 );
or ( n47640 , n47636 , n47639 );
buf ( n47641 , n34158 );
not ( n47642 , n47641 );
buf ( n47643 , n34241 );
nand ( n47644 , n47642 , n47643 );
nand ( n47645 , n47640 , n47644 );
buf ( n47646 , n30176 );
not ( n47647 , n47646 );
not ( n47648 , n47647 );
buf ( n47649 , n29856 );
not ( n47650 , n47649 );
or ( n47651 , n47648 , n47650 );
buf ( n47652 , n29820 );
buf ( n47653 , n41033 );
not ( n47654 , n47653 );
nand ( n47655 , n47652 , n47654 );
nand ( n47656 , n47651 , n47655 );
nor ( n47657 , n47645 , n47656 );
buf ( n47658 , n30019 );
not ( n47659 , n47658 );
not ( n47660 , n47659 );
buf ( n47661 , n46449 );
not ( n47662 , n47661 );
or ( n47663 , n47660 , n47662 );
not ( n47664 , n46428 );
buf ( n47665 , n47664 );
buf ( n47666 , n38124 );
not ( n47667 , n47666 );
nand ( n47668 , n47665 , n47667 );
nand ( n47669 , n47663 , n47668 );
buf ( n47670 , n27932 );
not ( n47671 , n47670 );
not ( n47672 , n47671 );
buf ( n47673 , n46485 );
not ( n47674 , n47673 );
or ( n47675 , n47672 , n47674 );
buf ( n47676 , n46465 );
buf ( n47677 , n27885 );
not ( n47678 , n47677 );
nand ( n47679 , n47676 , n47678 );
nand ( n47680 , n47675 , n47679 );
nor ( n47681 , n47669 , n47680 );
nand ( n47682 , n47585 , n47633 , n47657 , n47681 );
nor ( n47683 , n47623 , n47625 );
nor ( n47684 , n47627 , n47629 );
or ( n47685 , n47683 , n47684 );
nand ( n47686 , n47685 , n47626 );
or ( n47687 , n47621 , n47686 );
nor ( n47688 , n47613 , n47611 );
and ( n47689 , n47620 , n47688 );
nor ( n47690 , n47617 , n47619 );
nor ( n47691 , n47689 , n47690 );
nand ( n47692 , n47687 , n47691 );
nand ( n47693 , n47692 , n47608 );
not ( n47694 , n47596 );
nor ( n47695 , n47600 , n47598 );
not ( n47696 , n47695 );
not ( n47697 , n47606 );
or ( n47698 , n47696 , n47697 );
not ( n47699 , n47603 );
nand ( n47700 , n47699 , n47604 );
nand ( n47701 , n47698 , n47700 );
and ( n47702 , n47694 , n47701 );
nor ( n47703 , n47589 , n47587 );
not ( n47704 , n47703 );
not ( n47705 , n47595 );
or ( n47706 , n47704 , n47705 );
not ( n47707 , n47594 );
nand ( n47708 , n47707 , n47592 );
nand ( n47709 , n47706 , n47708 );
nor ( n47710 , n47702 , n47709 );
nand ( n47711 , n47693 , n47710 );
nand ( n47712 , n47711 , n47657 , n47681 );
nor ( n47713 , n47676 , n47678 );
nor ( n47714 , n47673 , n47671 );
or ( n47715 , n47713 , n47714 );
nand ( n47716 , n47715 , n47679 );
or ( n47717 , n47669 , n47716 );
nor ( n47718 , n47661 , n47659 );
and ( n47719 , n47668 , n47718 );
nor ( n47720 , n47665 , n47667 );
nor ( n47721 , n47719 , n47720 );
nand ( n47722 , n47717 , n47721 );
and ( n47723 , n47657 , n47722 );
nor ( n47724 , n47649 , n47647 );
and ( n47725 , n47655 , n47724 );
nor ( n47726 , n47652 , n47654 );
nor ( n47727 , n47725 , n47726 );
or ( n47728 , n47645 , n47727 );
nor ( n47729 , n47638 , n47635 );
and ( n47730 , n47644 , n47729 );
not ( n47731 , n47641 );
nor ( n47732 , n47731 , n47643 );
nor ( n47733 , n47730 , n47732 );
nand ( n47734 , n47728 , n47733 );
nor ( n47735 , n47723 , n47734 );
and ( n47736 , n47682 , n47712 , n47735 );
buf ( n47737 , n47736 );
or ( n47738 , n47737 , n46752 );
nand ( n47739 , n47738 , n46754 );
and ( n47740 , n47739 , n47059 );
not ( n47741 , n47737 );
not ( n47742 , n46752 );
nand ( n47743 , n47742 , n47056 );
nor ( n47744 , n47741 , n47743 );
nor ( n47745 , n47740 , n47744 );
not ( n47746 , n47437 );
not ( n47747 , n47440 );
nor ( n47748 , n47747 , n46746 );
and ( n47749 , n47746 , n47748 );
not ( n47750 , n25388 );
not ( n47751 , n19214 );
or ( n47752 , n47750 , n47751 );
nand ( n47753 , n47752 , n25045 );
and ( n47754 , n47753 , n25048 );
nor ( n47755 , n47754 , n19146 );
not ( n47756 , n47748 );
not ( n47757 , n47056 );
and ( n47758 , n47756 , n47757 );
nor ( n47759 , n47758 , n46754 );
nor ( n47760 , n47749 , n47755 , n47759 );
nand ( n47761 , n47442 , n47745 , n47760 );
nor ( n47762 , n46756 , n47761 );
nand ( n47763 , n46753 , n47762 );
buf ( n47764 , n47763 );
buf ( n47765 , n47764 );
not ( n47766 , n275550 );
buf ( n47767 , n47766 );
buf ( n47768 , n47767 );
or ( n47769 , n36036 , n23381 );
and ( n47770 , n36045 , n39562 );
not ( n47771 , n41937 );
nor ( n47772 , n47771 , n41967 );
not ( n47773 , n47772 );
and ( n47774 , n41903 , n41922 , n41933 );
not ( n47775 , n41933 );
not ( n47776 , n41956 );
or ( n47777 , n47775 , n47776 );
not ( n47778 , n41964 );
nand ( n47779 , n47777 , n47778 );
nor ( n47780 , n47774 , n47779 );
not ( n47781 , n47780 );
or ( n47782 , n47773 , n47781 );
or ( n47783 , n47780 , n47772 );
nand ( n47784 , n47782 , n47783 );
buf ( n47785 , n47784 );
not ( n47786 , n47785 );
not ( n47787 , n36155 );
or ( n47788 , n47786 , n47787 );
not ( n47789 , n42035 );
nor ( n47790 , n47789 , n42066 );
not ( n47791 , n47790 );
and ( n47792 , n42002 , n42021 , n42031 );
not ( n47793 , n42031 );
not ( n47794 , n42055 );
or ( n47795 , n47793 , n47794 );
not ( n47796 , n42063 );
nand ( n47797 , n47795 , n47796 );
nor ( n47798 , n47792 , n47797 );
not ( n47799 , n47798 );
or ( n47800 , n47791 , n47799 );
or ( n47801 , n47798 , n47790 );
nand ( n47802 , n47800 , n47801 );
buf ( n47803 , n47802 );
nand ( n47804 , n36159 , n47803 );
nand ( n47805 , n47788 , n47804 );
nor ( n47806 , n47770 , n47805 );
nand ( n47807 , n47769 , n47806 );
nand ( n47808 , n47807 , n20645 );
not ( n47809 , n42131 );
nor ( n47810 , n47809 , n42157 );
not ( n47811 , n47810 );
and ( n47812 , n42095 , n42116 , n42127 );
not ( n47813 , n42127 );
not ( n47814 , n42146 );
or ( n47815 , n47813 , n47814 );
not ( n47816 , n42154 );
nand ( n47817 , n47815 , n47816 );
nor ( n47818 , n47812 , n47817 );
not ( n47819 , n47818 );
or ( n47820 , n47811 , n47819 );
or ( n47821 , n47818 , n47810 );
nand ( n47822 , n47820 , n47821 );
buf ( n47823 , n47822 );
nand ( n47824 , n36267 , n47823 );
not ( n47825 , n42216 );
nor ( n47826 , n47825 , n42242 );
not ( n47827 , n47826 );
and ( n47828 , n42181 , n42202 , n42212 );
not ( n47829 , n42212 );
not ( n47830 , n42231 );
or ( n47831 , n47829 , n47830 );
not ( n47832 , n42239 );
nand ( n47833 , n47831 , n47832 );
nor ( n47834 , n47828 , n47833 );
not ( n47835 , n47834 );
or ( n47836 , n47827 , n47835 );
or ( n47837 , n47834 , n47826 );
nand ( n47838 , n47836 , n47837 );
buf ( n47839 , n47838 );
nand ( n47840 , n36371 , n47839 );
and ( n47841 , n36474 , n277906 );
or ( n47842 , n20654 , n39561 );
nand ( n47843 , n47842 , n39056 );
nor ( n47844 , n47841 , n47843 );
nand ( n47845 , n47808 , n47824 , n47840 , n47844 );
buf ( n47846 , n47845 );
buf ( n47847 , n47846 );
not ( n47848 , n275925 );
buf ( n47849 , n47848 );
buf ( n47850 , n47849 );
not ( n47851 , n275925 );
buf ( n47852 , n47851 );
buf ( n47853 , n47852 );
buf ( n47854 , n275554 );
or ( n47855 , n33723 , n19216 );
and ( n47856 , n33737 , n19360 );
nand ( n47857 , n33754 , n29075 );
and ( n47858 , n33162 , n27932 );
nor ( n47859 , n33743 , n19317 );
nor ( n47860 , n47858 , n47859 );
nand ( n47861 , n19387 , n18800 );
nand ( n47862 , n47857 , n47860 , n47861 );
nor ( n47863 , n47856 , n47862 );
nand ( n47864 , n33773 , n35150 );
and ( n47865 , n47863 , n47864 );
nand ( n47866 , n47855 , n47865 );
buf ( n47867 , n47866 );
buf ( n47868 , n47867 );
not ( n47869 , n275929 );
buf ( n47870 , n47869 );
buf ( n47871 , n47870 );
or ( n47872 , n21657 , n26364 );
and ( n47873 , n39065 , n14528 );
and ( n47874 , n21678 , n26367 );
and ( n47875 , n26384 , n21681 );
nor ( n47876 , n47874 , n47875 );
nand ( n47877 , n26395 , n21685 );
nand ( n47878 , n26374 , n21668 );
nand ( n47879 , n47876 , n47877 , n47878 );
nor ( n47880 , n47873 , n47879 );
nand ( n47881 , n47872 , n47880 );
buf ( n47882 , n47881 );
buf ( n47883 , n47882 );
or ( n47884 , n27165 , n21696 );
nand ( n47885 , n34674 , n13452 );
nand ( n47886 , n47884 , n47885 );
buf ( n47887 , n47886 );
buf ( n47888 , n47887 );
not ( n47889 , n275929 );
buf ( n47890 , n47889 );
buf ( n47891 , n47890 );
not ( n47892 , n27641 );
nand ( n47893 , n47892 , n40813 );
or ( n47894 , n32828 , n47893 );
buf ( n47895 , n9254 );
nand ( n47896 , n27641 , n47895 );
nand ( n47897 , n47894 , n47896 );
buf ( n47898 , n47897 );
buf ( n47899 , n47898 );
buf ( n47900 , n275554 );
buf ( n47901 , n275554 );
not ( n47902 , n275929 );
buf ( n47903 , n47902 );
buf ( n47904 , n47903 );
not ( n47905 , n275929 );
buf ( n47906 , n47905 );
buf ( n47907 , n47906 );
not ( n47908 , n275550 );
buf ( n47909 , n47908 );
buf ( n47910 , n47909 );
or ( n47911 , n30256 , n14909 );
nand ( n47912 , n30318 , n16970 );
and ( n47913 , n30361 , n17405 );
nand ( n47914 , n35657 , n17545 );
nand ( n47915 , n32339 , n30374 );
nand ( n47916 , n17502 , n24937 );
nand ( n47917 , n17562 , n14631 );
nand ( n47918 , n47914 , n47915 , n47916 , n47917 );
nor ( n47919 , n47913 , n47918 );
and ( n47920 , n47912 , n47919 );
nand ( n47921 , n47911 , n47920 );
buf ( n47922 , n47921 );
buf ( n47923 , n47922 );
or ( n47924 , n32992 , n20743 );
and ( n47925 , n33026 , n17405 );
not ( n47926 , n33032 );
not ( n47927 , n20765 );
and ( n47928 , n47926 , n47927 );
and ( n47929 , n32339 , n33039 );
nor ( n47930 , n47928 , n47929 );
nand ( n47931 , n20785 , n33044 );
nand ( n47932 , n17562 , n13870 );
nand ( n47933 , n47930 , n47931 , n47932 );
nor ( n47934 , n47925 , n47933 );
nand ( n47935 , n33009 , n16970 );
and ( n47936 , n47934 , n47935 );
nand ( n47937 , n47924 , n47936 );
buf ( n47938 , n47937 );
buf ( n47939 , n47938 );
buf ( n47940 , n275554 );
not ( n47941 , n275550 );
buf ( n47942 , n47941 );
buf ( n47943 , n47942 );
buf ( n47944 , n275554 );
not ( n47945 , n275925 );
buf ( n47946 , n47945 );
buf ( n47947 , n47946 );
buf ( n47948 , n275554 );
buf ( n47949 , n275554 );
buf ( n47950 , n275554 );
nand ( n47951 , n22192 , n32833 );
or ( n47952 , n32828 , n47951 );
nand ( n47953 , n40816 , n9387 );
nand ( n47954 , n47952 , n47953 );
buf ( n47955 , n47954 );
buf ( n47956 , n47955 );
buf ( n47957 , n275554 );
not ( n47958 , n275929 );
buf ( n47959 , n47958 );
buf ( n47960 , n47959 );
not ( n47961 , n275929 );
buf ( n47962 , n47961 );
buf ( n47963 , n47962 );
or ( n47964 , n36036 , n26418 );
and ( n47965 , n45676 , n275873 );
not ( n47966 , n41945 );
nor ( n47967 , n47966 , n41941 );
not ( n47968 , n47967 );
and ( n47969 , n41896 , n36068 );
and ( n47970 , n47969 , n36137 , n41916 );
not ( n47971 , n41916 );
or ( n47972 , n41902 , n47971 );
nand ( n47973 , n47972 , n41943 );
nor ( n47974 , n47970 , n47973 );
not ( n47975 , n47974 );
or ( n47976 , n47968 , n47975 );
or ( n47977 , n47974 , n47967 );
nand ( n47978 , n47976 , n47977 );
buf ( n47979 , n47978 );
not ( n47980 , n47979 );
not ( n47981 , n36155 );
or ( n47982 , n47980 , n47981 );
and ( n47983 , n42044 , n42019 );
not ( n47984 , n47983 );
and ( n47985 , n41988 , n36179 );
and ( n47986 , n47985 , n36243 , n42015 );
not ( n47987 , n42015 );
or ( n47988 , n42001 , n47987 );
nand ( n47989 , n47988 , n42521 );
nor ( n47990 , n47986 , n47989 );
not ( n47991 , n47990 );
or ( n47992 , n47984 , n47991 );
or ( n47993 , n47990 , n47983 );
nand ( n47994 , n47992 , n47993 );
buf ( n47995 , n47994 );
nand ( n47996 , n36159 , n47995 );
nand ( n47997 , n47982 , n47996 );
nor ( n47998 , n47965 , n47997 );
nand ( n47999 , n47964 , n47998 );
nand ( n48000 , n47999 , n20645 );
not ( n48001 , n42103 );
nor ( n48002 , n48001 , n42138 );
not ( n48003 , n48002 );
and ( n48004 , n42085 , n36285 );
and ( n48005 , n48004 , n36353 , n42099 );
nand ( n48006 , n42089 , n42099 );
nand ( n48007 , n48006 , n42534 );
nor ( n48008 , n48005 , n48007 );
not ( n48009 , n48008 );
or ( n48010 , n48003 , n48009 );
or ( n48011 , n48008 , n48002 );
nand ( n48012 , n48010 , n48011 );
buf ( n48013 , n48012 );
nand ( n48014 , n36267 , n48013 );
not ( n48015 , n42189 );
nor ( n48016 , n48015 , n42223 );
not ( n48017 , n48016 );
and ( n48018 , n42171 , n36389 );
and ( n48019 , n48018 , n36456 , n42185 );
nand ( n48020 , n42175 , n42185 );
nand ( n48021 , n48020 , n42543 );
nor ( n48022 , n48019 , n48021 );
not ( n48023 , n48022 );
or ( n48024 , n48017 , n48023 );
or ( n48025 , n48022 , n48016 );
nand ( n48026 , n48024 , n48025 );
buf ( n48027 , n48026 );
nand ( n48028 , n36371 , n48027 );
and ( n48029 , n36474 , n11432 );
or ( n48030 , n20654 , n275872 );
nand ( n48031 , n48030 , n32759 );
nor ( n48032 , n48029 , n48031 );
nand ( n48033 , n48000 , n48014 , n48028 , n48032 );
buf ( n48034 , n48033 );
buf ( n48035 , n48034 );
not ( n48036 , n275929 );
buf ( n48037 , n48036 );
buf ( n48038 , n48037 );
not ( n48039 , n275929 );
buf ( n48040 , n48039 );
buf ( n48041 , n48040 );
buf ( n48042 , n275554 );
not ( n48043 , n14542 );
or ( n48044 , n48043 , n20961 );
not ( n48045 , n9444 );
or ( n48046 , n28247 , n48045 );
nand ( n48047 , n48044 , n48046 );
buf ( n48048 , n48047 );
buf ( n48049 , n48048 );
not ( n48050 , n275929 );
buf ( n48051 , n48050 );
buf ( n48052 , n48051 );
not ( n48053 , n275925 );
buf ( n48054 , n48053 );
buf ( n48055 , n48054 );
and ( n48056 , n21030 , n18642 );
not ( n48057 , n21030 );
and ( n48058 , n48057 , n28145 );
nor ( n48059 , n48056 , n48058 );
buf ( n48060 , n48059 );
buf ( n48061 , n48060 );
or ( n48062 , n44919 , n20743 );
nand ( n48063 , n44939 , n16970 );
nand ( n48064 , n44962 , n17405 );
nand ( n48065 , n17411 , n44976 );
nand ( n48066 , n20785 , n44978 );
nand ( n48067 , n17562 , n13495 );
nand ( n48068 , n17545 , n44967 );
and ( n48069 , n48065 , n48066 , n48067 , n48068 );
and ( n48070 , n48063 , n48064 , n48069 );
nand ( n48071 , n48062 , n48070 );
buf ( n48072 , n48071 );
buf ( n48073 , n48072 );
or ( n48074 , n31056 , n19216 );
and ( n48075 , n31076 , n19360 );
nand ( n48076 , n31094 , n29075 );
and ( n48077 , n33162 , n31098 );
not ( n48078 , n31083 );
nor ( n48079 , n48078 , n29537 );
nor ( n48080 , n48077 , n48079 );
nand ( n48081 , n19387 , n18830 );
nand ( n48082 , n48076 , n48080 , n48081 );
nor ( n48083 , n48075 , n48082 );
nand ( n48084 , n31122 , n44740 );
and ( n48085 , n48083 , n48084 );
nand ( n48086 , n48074 , n48085 );
buf ( n48087 , n48086 );
buf ( n48088 , n48087 );
nand ( n48089 , n25064 , n25097 );
buf ( n48090 , n36702 );
buf ( n48091 , n25309 );
and ( n48092 , n48090 , n48091 );
buf ( n48093 , n48092 );
buf ( n48094 , n48093 );
not ( n48095 , n48094 );
buf ( n48096 , n25264 );
buf ( n48097 , n25128 );
and ( n48098 , n48096 , n48097 );
buf ( n48099 , n25329 );
nor ( n48100 , n48098 , n48099 );
buf ( n48101 , n48100 );
buf ( n48102 , n48101 );
not ( n48103 , n48102 );
or ( n48104 , n48095 , n48103 );
buf ( n48105 , n48101 );
buf ( n48106 , n48093 );
or ( n48107 , n48105 , n48106 );
nand ( n48108 , n48104 , n48107 );
buf ( n48109 , n48108 );
buf ( n48110 , n48109 );
not ( n48111 , n48110 );
nor ( n48112 , n48111 , n25389 );
nand ( n48113 , n25397 , n275652 );
buf ( n48114 , n36738 );
buf ( n48115 , n25653 );
and ( n48116 , n48114 , n48115 );
buf ( n48117 , n48116 );
buf ( n48118 , n48117 );
not ( n48119 , n48118 );
buf ( n48120 , n25586 );
buf ( n48121 , n25453 );
and ( n48122 , n48120 , n48121 );
buf ( n48123 , n25642 );
nor ( n48124 , n48122 , n48123 );
buf ( n48125 , n48124 );
buf ( n48126 , n48125 );
not ( n48127 , n48126 );
or ( n48128 , n48119 , n48127 );
buf ( n48129 , n48125 );
buf ( n48130 , n48117 );
or ( n48131 , n48129 , n48130 );
nand ( n48132 , n48128 , n48131 );
buf ( n48133 , n48132 );
buf ( n48134 , n48133 );
and ( n48135 , n25402 , n48134 );
nor ( n48136 , n48135 , n20517 );
buf ( n48137 , n25748 );
buf ( n48138 , n25964 );
and ( n48139 , n48137 , n48138 );
buf ( n48140 , n48139 );
buf ( n48141 , n48140 );
not ( n48142 , n48141 );
buf ( n48143 , n25902 );
buf ( n48144 , n25770 );
and ( n48145 , n48143 , n48144 );
buf ( n48146 , n25956 );
nor ( n48147 , n48145 , n48146 );
buf ( n48148 , n48147 );
buf ( n48149 , n48148 );
not ( n48150 , n48149 );
or ( n48151 , n48142 , n48150 );
buf ( n48152 , n48148 );
buf ( n48153 , n48140 );
or ( n48154 , n48152 , n48153 );
nand ( n48155 , n48151 , n48154 );
buf ( n48156 , n48155 );
buf ( n48157 , n48156 );
nand ( n48158 , n25717 , n48157 );
nand ( n48159 , n48113 , n48136 , n48158 );
nor ( n48160 , n48112 , n48159 );
buf ( n48161 , n26050 );
buf ( n48162 , n26253 );
and ( n48163 , n48161 , n48162 );
buf ( n48164 , n48163 );
buf ( n48165 , n48164 );
not ( n48166 , n48165 );
buf ( n48167 , n26212 );
buf ( n48168 , n26078 );
and ( n48169 , n48167 , n48168 );
buf ( n48170 , n26270 );
nor ( n48171 , n48169 , n48170 );
buf ( n48172 , n48171 );
buf ( n48173 , n48172 );
not ( n48174 , n48173 );
or ( n48175 , n48166 , n48174 );
buf ( n48176 , n48172 );
buf ( n48177 , n48164 );
or ( n48178 , n48176 , n48177 );
nand ( n48179 , n48175 , n48178 );
buf ( n48180 , n48179 );
buf ( n48181 , n48180 );
nand ( n48182 , n26027 , n48181 );
nand ( n48183 , n48089 , n48160 , n48182 );
buf ( n48184 , n48183 );
buf ( n48185 , n48184 );
not ( n48186 , n275929 );
buf ( n48187 , n48186 );
buf ( n48188 , n48187 );
not ( n48189 , n26679 );
or ( n48190 , n48189 , n22335 );
or ( n48191 , n275557 , n19191 );
nand ( n48192 , n48190 , n48191 );
buf ( n48193 , n48192 );
buf ( n48194 , n48193 );
or ( n48195 , n39686 , n28146 );
nand ( n48196 , n24450 , n18587 );
nand ( n48197 , n48195 , n48196 );
buf ( n48198 , n48197 );
buf ( n48199 , n48198 );
not ( n48200 , n275550 );
buf ( n48201 , n48200 );
buf ( n48202 , n48201 );
not ( n48203 , n275550 );
buf ( n48204 , n48203 );
buf ( n48205 , n48204 );
buf ( n48206 , n275554 );
buf ( n48207 , n275554 );
buf ( n48208 , n275554 );
buf ( n48209 , n275554 );
buf ( n48210 , n275554 );
not ( n48211 , n39588 );
and ( n48212 , n9100 , n48211 , n9158 );
buf ( n48213 , n48212 );
buf ( n48214 , n48213 );
nor ( n48215 , n275916 , n275914 );
not ( n48216 , n48215 );
not ( n48217 , n275907 );
or ( n48218 , n48216 , n48217 );
or ( n48219 , n275907 , n48215 );
nand ( n48220 , n48218 , n48219 );
buf ( n48221 , n48220 );
buf ( n48222 , n48221 );
not ( n48223 , n275925 );
buf ( n48224 , n48223 );
buf ( n48225 , n48224 );
not ( n48226 , n275929 );
buf ( n48227 , n48226 );
buf ( n48228 , n48227 );
not ( n48229 , n275925 );
buf ( n48230 , n48229 );
buf ( n48231 , n48230 );
not ( n48232 , n275925 );
buf ( n48233 , n48232 );
buf ( n48234 , n48233 );
not ( n48235 , n275929 );
buf ( n48236 , n48235 );
buf ( n48237 , n48236 );
not ( n48238 , n275550 );
buf ( n48239 , n48238 );
buf ( n48240 , n48239 );
not ( n48241 , n275925 );
buf ( n48242 , n48241 );
buf ( n48243 , n48242 );
not ( n48244 , n34302 );
not ( n48245 , n31962 );
or ( n48246 , n48244 , n48245 );
and ( n48247 , n32029 , n28430 );
nand ( n48248 , n32051 , n34307 );
nand ( n48249 , n28451 , n32057 );
and ( n48250 , n32755 , n32055 );
and ( n48251 , n34848 , n277533 );
and ( n48252 , n34313 , n9355 );
nor ( n48253 , n48250 , n48251 , n48252 );
nand ( n48254 , n48248 , n48249 , n48253 );
nor ( n48255 , n48247 , n48254 );
nand ( n48256 , n48246 , n48255 );
buf ( n48257 , n48256 );
buf ( n48258 , n48257 );
not ( n48259 , n275925 );
buf ( n48260 , n48259 );
buf ( n48261 , n48260 );
not ( n48262 , n33794 );
or ( n48263 , n48262 , n21774 );
nand ( n48264 , n21774 , n9527 );
nand ( n48265 , n48263 , n48264 );
buf ( n48266 , n48265 );
buf ( n48267 , n48266 );
not ( n48268 , n275550 );
buf ( n48269 , n48268 );
buf ( n48270 , n48269 );
not ( n48271 , n275925 );
buf ( n48272 , n48271 );
buf ( n48273 , n48272 );
not ( n48274 , n275929 );
buf ( n48275 , n48274 );
buf ( n48276 , n48275 );
not ( n48277 , n275550 );
buf ( n48278 , n48277 );
buf ( n48279 , n48278 );
nand ( n48280 , n25064 , n25276 );
buf ( n48281 , n25282 );
not ( n48282 , n48281 );
buf ( n48283 , n25348 );
nand ( n48284 , n48282 , n48283 );
buf ( n48285 , n48284 );
buf ( n48286 , n48285 );
not ( n48287 , n48286 );
buf ( n48288 , n28514 );
not ( n48289 , n48288 );
or ( n48290 , n48287 , n48289 );
buf ( n48291 , n28514 );
buf ( n48292 , n48285 );
or ( n48293 , n48291 , n48292 );
nand ( n48294 , n48290 , n48293 );
buf ( n48295 , n48294 );
buf ( n48296 , n48295 );
not ( n48297 , n48296 );
nor ( n48298 , n48297 , n25389 );
nand ( n48299 , n25397 , n275882 );
buf ( n48300 , n25603 );
not ( n48301 , n48300 );
buf ( n48302 , n25674 );
nand ( n48303 , n48301 , n48302 );
buf ( n48304 , n48303 );
buf ( n48305 , n48304 );
not ( n48306 , n48305 );
buf ( n48307 , n28655 );
not ( n48308 , n48307 );
or ( n48309 , n48306 , n48308 );
buf ( n48310 , n28655 );
buf ( n48311 , n48304 );
or ( n48312 , n48310 , n48311 );
nand ( n48313 , n48309 , n48312 );
buf ( n48314 , n48313 );
buf ( n48315 , n48314 );
and ( n48316 , n25402 , n48315 );
nor ( n48317 , n48316 , n41809 );
buf ( n48318 , n25917 );
not ( n48319 , n48318 );
buf ( n48320 , n25985 );
nand ( n48321 , n48319 , n48320 );
buf ( n48322 , n48321 );
buf ( n48323 , n48322 );
not ( n48324 , n48323 );
buf ( n48325 , n28796 );
not ( n48326 , n48325 );
or ( n48327 , n48324 , n48326 );
buf ( n48328 , n28796 );
buf ( n48329 , n48322 );
or ( n48330 , n48328 , n48329 );
nand ( n48331 , n48327 , n48330 );
buf ( n48332 , n48331 );
buf ( n48333 , n48332 );
nand ( n48334 , n25717 , n48333 );
nand ( n48335 , n48299 , n48317 , n48334 );
nor ( n48336 , n48298 , n48335 );
buf ( n48337 , n26226 );
not ( n48338 , n48337 );
buf ( n48339 , n26289 );
nand ( n48340 , n48338 , n48339 );
buf ( n48341 , n48340 );
buf ( n48342 , n48341 );
not ( n48343 , n48342 );
buf ( n48344 , n28935 );
not ( n48345 , n48344 );
or ( n48346 , n48343 , n48345 );
buf ( n48347 , n28935 );
buf ( n48348 , n48341 );
or ( n48349 , n48347 , n48348 );
nand ( n48350 , n48346 , n48349 );
buf ( n48351 , n48350 );
buf ( n48352 , n48351 );
nand ( n48353 , n26027 , n48352 );
nand ( n48354 , n48280 , n48336 , n48353 );
buf ( n48355 , n48354 );
buf ( n48356 , n48355 );
nand ( n48357 , n30906 , n31422 );
nand ( n48358 , n30961 , n31437 );
nand ( n48359 , n30988 , n31449 );
and ( n48360 , n36530 , n12185 );
not ( n48361 , n277771 );
not ( n48362 , n28357 );
or ( n48363 , n48361 , n48362 );
or ( n48364 , n32061 , n277762 );
nand ( n48365 , n48363 , n48364 );
nor ( n48366 , n48360 , n48365 );
nand ( n48367 , n31460 , n12370 );
and ( n48368 , n48359 , n48366 , n48367 );
nand ( n48369 , n48357 , n48358 , n48368 );
buf ( n48370 , n48369 );
buf ( n48371 , n48370 );
buf ( n48372 , n275554 );
or ( n48373 , n35683 , n19636 );
nand ( n48374 , n35693 , n20353 );
nand ( n48375 , n35702 , n20515 );
nand ( n48376 , n19648 , n36592 );
nand ( n48377 , n35709 , n19645 );
nand ( n48378 , n19644 , n35714 );
not ( n48379 , n38457 );
and ( n48380 , n48377 , n48378 , n48379 );
and ( n48381 , n48374 , n48375 , n48376 , n48380 );
nand ( n48382 , n48373 , n48381 );
buf ( n48383 , n48382 );
buf ( n48384 , n48383 );
or ( n48385 , n35212 , n28146 );
nand ( n48386 , n24450 , n18794 );
nand ( n48387 , n48385 , n48386 );
buf ( n48388 , n48387 );
buf ( n48389 , n48388 );
buf ( n48390 , n275554 );
or ( n48391 , n23696 , n12108 , n11729 );
not ( n48392 , n23687 );
and ( n48393 , n12097 , n11729 );
and ( n48394 , n12108 , n9136 );
nor ( n48395 , n48393 , n48394 );
or ( n48396 , n48392 , n48395 );
nand ( n48397 , n48391 , n48396 );
nand ( n48398 , n48397 , n28436 , n11732 );
or ( n48399 , n37985 , n48398 );
not ( n48400 , n48397 );
and ( n48401 , n48400 , n32819 , n9271 );
not ( n48402 , n22146 );
or ( n48403 , n48402 , n12679 , n11729 );
nand ( n48404 , n48403 , n23696 );
and ( n48405 , n12679 , n277356 );
not ( n48406 , n12679 );
and ( n48407 , n48406 , n9367 );
nor ( n48408 , n48405 , n48407 );
nor ( n48409 , n48408 , n11729 );
and ( n48410 , n48404 , n48409 );
not ( n48411 , n48404 );
and ( n48412 , n48411 , n9271 );
nor ( n48413 , n48410 , n48412 );
nor ( n48414 , n48413 , n32819 );
nor ( n48415 , n48401 , n48414 );
nand ( n48416 , n48399 , n48415 );
buf ( n48417 , n48416 );
buf ( n48418 , n48417 );
not ( n48419 , n275925 );
buf ( n48420 , n48419 );
buf ( n48421 , n48420 );
buf ( n48422 , n275554 );
not ( n48423 , n275929 );
buf ( n48424 , n48423 );
buf ( n48425 , n48424 );
buf ( n48426 , n275554 );
buf ( n48427 , n275554 );
and ( n48428 , n20950 , n14765 );
not ( n48429 , n20950 );
and ( n48430 , n48429 , n40631 );
nor ( n48431 , n48428 , n48430 );
buf ( n48432 , n48431 );
buf ( n48433 , n48432 );
buf ( n48434 , n275554 );
buf ( n48435 , n275554 );
buf ( n48436 , n275554 );
buf ( n48437 , n275554 );
not ( n48438 , n275925 );
buf ( n48439 , n48438 );
buf ( n48440 , n48439 );
not ( n48441 , n275929 );
buf ( n48442 , n48441 );
buf ( n48443 , n48442 );
or ( n48444 , n39249 , n19636 );
not ( n48445 , n38353 );
not ( n48446 , n39290 );
and ( n48447 , n48445 , n48446 );
and ( n48448 , n39268 , n20353 );
nor ( n48449 , n48447 , n48448 );
and ( n48450 , n39284 , n20515 );
not ( n48451 , n36763 );
nand ( n48452 , n39304 , n20560 );
nand ( n48453 , n19644 , n39294 );
nand ( n48454 , n48451 , n48452 , n48453 );
nor ( n48455 , n48450 , n48454 );
and ( n48456 , n48449 , n48455 );
nand ( n48457 , n48444 , n48456 );
buf ( n48458 , n48457 );
buf ( n48459 , n48458 );
not ( n48460 , n275925 );
buf ( n48461 , n48460 );
buf ( n48462 , n48461 );
not ( n48463 , n275929 );
buf ( n48464 , n48463 );
buf ( n48465 , n48464 );
not ( n48466 , n275925 );
buf ( n48467 , n48466 );
buf ( n48468 , n48467 );
or ( n48469 , n39491 , n27640 );
nand ( n48470 , n27640 , n11018 );
nand ( n48471 , n48469 , n48470 );
buf ( n48472 , n48471 );
buf ( n48473 , n48472 );
not ( n48474 , n275925 );
buf ( n48475 , n48474 );
buf ( n48476 , n48475 );
buf ( n48477 , n275554 );
buf ( n48478 , n275554 );
nand ( n48479 , n28398 , n28306 );
nand ( n48480 , n28426 , n33875 );
and ( n48481 , n28332 , n28433 );
and ( n48482 , n28242 , n12220 );
nor ( n48483 , n48481 , n48482 );
and ( n48484 , n28231 , n28456 );
or ( n48485 , n28354 , n11377 );
nand ( n48486 , n28236 , n11392 );
nand ( n48487 , n48485 , n48486 );
nor ( n48488 , n48484 , n48487 );
nand ( n48489 , n48479 , n48480 , n48483 , n48488 );
buf ( n48490 , n48489 );
buf ( n48491 , n48490 );
not ( n48492 , n275925 );
buf ( n48493 , n48492 );
buf ( n48494 , n48493 );
or ( n48495 , n40356 , n19216 );
and ( n48496 , n40406 , n19360 );
nand ( n48497 , n40421 , n29075 );
and ( n48498 , n33162 , n40409 );
and ( n48499 , n30142 , n18525 );
not ( n48500 , n30142 );
and ( n48501 , n48500 , n30143 );
nor ( n48502 , n48499 , n48501 );
nor ( n48503 , n48502 , n29537 );
nor ( n48504 , n48498 , n48503 );
nand ( n48505 , n19387 , n18536 );
nand ( n48506 , n48497 , n48504 , n48505 );
nor ( n48507 , n48496 , n48506 );
nand ( n48508 , n40383 , n44740 );
and ( n48509 , n48507 , n48508 );
nand ( n48510 , n48495 , n48509 );
buf ( n48511 , n48510 );
buf ( n48512 , n48511 );
or ( n48513 , n31307 , n26365 );
nand ( n48514 , n31356 , n26370 );
nand ( n48515 , n31320 , n26374 );
not ( n48516 , n31339 );
nor ( n48517 , n48516 , n26390 );
nand ( n48518 , n31327 , n26393 );
nand ( n48519 , n26395 , n31332 );
nand ( n48520 , n17542 , n13910 );
nand ( n48521 , n48518 , n48519 , n48520 );
nor ( n48522 , n48517 , n48521 );
and ( n48523 , n48514 , n48515 , n48522 );
nand ( n48524 , n48513 , n48523 );
buf ( n48525 , n48524 );
buf ( n48526 , n48525 );
or ( n48527 , n23886 , n21696 );
nand ( n48528 , n21697 , n13945 );
nand ( n48529 , n48527 , n48528 );
buf ( n48530 , n48529 );
buf ( n48531 , n48530 );
not ( n48532 , n275929 );
buf ( n48533 , n48532 );
buf ( n48534 , n48533 );
or ( n48535 , n32941 , n14908 );
not ( n48536 , n17501 );
not ( n48537 , n38141 );
and ( n48538 , n48536 , n48537 );
and ( n48539 , n32948 , n16968 );
nor ( n48540 , n48538 , n48539 );
not ( n48541 , n20765 );
not ( n48542 , n32974 );
and ( n48543 , n48541 , n48542 );
and ( n48544 , n17411 , n32965 );
nor ( n48545 , n48543 , n48544 );
and ( n48546 , n17405 , n32955 );
not ( n48547 , n13644 );
nor ( n48548 , n17561 , n48547 );
nor ( n48549 , n48546 , n48548 );
and ( n48550 , n48540 , n48545 , n48549 );
nand ( n48551 , n48535 , n48550 );
buf ( n48552 , n48551 );
buf ( n48553 , n48552 );
not ( n48554 , n275929 );
buf ( n48555 , n48554 );
buf ( n48556 , n48555 );
or ( n48557 , n38928 , n23887 );
nand ( n48558 , n20951 , n13875 );
nand ( n48559 , n48557 , n48558 );
buf ( n48560 , n48559 );
buf ( n48561 , n48560 );
buf ( n48562 , n275554 );
buf ( n48563 , n275554 );
and ( n48564 , n27179 , n277551 );
not ( n48565 , n27179 );
and ( n48566 , n48565 , n32123 );
or ( n48567 , n48564 , n48566 );
buf ( n48568 , n48567 );
buf ( n48569 , n48568 );
not ( n48570 , n34302 );
not ( n48571 , n33596 );
or ( n48572 , n48570 , n48571 );
and ( n48573 , n33611 , n28430 );
nand ( n48574 , n33621 , n34307 );
nand ( n48575 , n28451 , n277672 );
and ( n48576 , n32755 , n12302 );
and ( n48577 , n34311 , n277696 );
and ( n48578 , n34313 , n9345 );
nor ( n48579 , n48576 , n48577 , n48578 );
nand ( n48580 , n48574 , n48575 , n48579 );
nor ( n48581 , n48573 , n48580 );
nand ( n48582 , n48572 , n48581 );
buf ( n48583 , n48582 );
buf ( n48584 , n48583 );
or ( n48585 , n26636 , n19216 );
and ( n48586 , n27046 , n19360 );
nand ( n48587 , n27079 , n29075 );
and ( n48588 , n33162 , n27050 );
and ( n48589 , n19318 , n40196 );
nor ( n48590 , n48588 , n48589 );
nand ( n48591 , n19387 , n18563 );
nand ( n48592 , n48587 , n48590 , n48591 );
nor ( n48593 , n48586 , n48592 );
nand ( n48594 , n26944 , n35150 );
and ( n48595 , n48593 , n48594 );
nand ( n48596 , n48585 , n48595 );
buf ( n48597 , n48596 );
buf ( n48598 , n48597 );
or ( n48599 , n37574 , n32074 );
not ( n48600 , n19649 );
not ( n48601 , n40534 );
and ( n48602 , n48600 , n48601 );
and ( n48603 , n37602 , n20353 );
nor ( n48604 , n48602 , n48603 );
and ( n48605 , n37625 , n20515 );
not ( n48606 , n25714 );
nand ( n48607 , n37636 , n20560 );
nand ( n48608 , n29494 , n37641 );
nand ( n48609 , n48606 , n48607 , n48608 );
nor ( n48610 , n48605 , n48609 );
and ( n48611 , n48604 , n48610 );
nand ( n48612 , n48599 , n48611 );
buf ( n48613 , n48612 );
buf ( n48614 , n48613 );
not ( n48615 , n275925 );
buf ( n48616 , n48615 );
buf ( n48617 , n48616 );
buf ( n48618 , n275554 );
not ( n48619 , n275550 );
buf ( n48620 , n48619 );
buf ( n48621 , n48620 );
buf ( n48622 , n275554 );
not ( n48623 , n275550 );
buf ( n48624 , n48623 );
buf ( n48625 , n48624 );
buf ( n48626 , n275554 );
buf ( n48627 , n275554 );
not ( n48628 , n275929 );
buf ( n48629 , n48628 );
buf ( n48630 , n48629 );
not ( n48631 , n275929 );
buf ( n48632 , n48631 );
buf ( n48633 , n48632 );
buf ( n48634 , n275554 );
not ( n48635 , n275550 );
buf ( n48636 , n48635 );
buf ( n48637 , n48636 );
not ( n48638 , n275925 );
buf ( n48639 , n48638 );
buf ( n48640 , n48639 );
or ( n48641 , n23989 , n19216 );
and ( n48642 , n24296 , n19360 );
nand ( n48643 , n24320 , n29075 );
not ( n48644 , n19317 );
not ( n48645 , n29487 );
and ( n48646 , n48644 , n48645 );
and ( n48647 , n33162 , n24325 );
nor ( n48648 , n48646 , n48647 );
nand ( n48649 , n19387 , n18945 );
nand ( n48650 , n48643 , n48648 , n48649 );
nor ( n48651 , n48642 , n48650 );
nand ( n48652 , n24213 , n35863 );
nand ( n48653 , n48641 , n48651 , n48652 );
buf ( n48654 , n48653 );
buf ( n48655 , n48654 );
or ( n48656 , n21172 , n19216 );
and ( n48657 , n21592 , n19360 );
not ( n48658 , n19317 );
not ( n48659 , n32080 );
and ( n48660 , n48658 , n48659 );
and ( n48661 , n19221 , n21624 );
nor ( n48662 , n48660 , n48661 );
nand ( n48663 , n21618 , n29075 );
nand ( n48664 , n19387 , n18731 );
nand ( n48665 , n48662 , n48663 , n48664 );
nor ( n48666 , n48657 , n48665 );
nand ( n48667 , n21499 , n19354 );
and ( n48668 , n48666 , n48667 );
nand ( n48669 , n48656 , n48668 );
buf ( n48670 , n48669 );
buf ( n48671 , n48670 );
buf ( n48672 , n275554 );
buf ( n48673 , n275554 );
not ( n48674 , n275925 );
buf ( n48675 , n48674 );
buf ( n48676 , n48675 );
not ( n48677 , n275929 );
buf ( n48678 , n48677 );
buf ( n48679 , n48678 );
buf ( n48680 , n275554 );
buf ( n48681 , n275554 );
or ( n48682 , n34696 , n26364 );
not ( n48683 , n26390 );
not ( n48684 , n13555 );
and ( n48685 , n48683 , n48684 );
nand ( n48686 , n34706 , n26370 );
nand ( n48687 , n34717 , n26374 );
nand ( n48688 , n26395 , n34723 );
and ( n48689 , n26393 , n34734 );
nor ( n48690 , n14830 , n32972 );
nor ( n48691 , n48689 , n48690 );
nand ( n48692 , n48686 , n48687 , n48688 , n48691 );
nor ( n48693 , n48685 , n48692 );
nand ( n48694 , n48682 , n48693 );
buf ( n48695 , n48694 );
buf ( n48696 , n48695 );
not ( n48697 , n18115 );
not ( n48698 , n22335 );
or ( n48699 , n48697 , n48698 );
not ( n48700 , n20292 );
or ( n48701 , n22335 , n48700 );
nand ( n48702 , n48699 , n48701 );
buf ( n48703 , n48702 );
buf ( n48704 , n48703 );
not ( n48705 , n275925 );
buf ( n48706 , n48705 );
buf ( n48707 , n48706 );
not ( n48708 , n275929 );
buf ( n48709 , n48708 );
buf ( n48710 , n48709 );
buf ( n48711 , n275554 );
not ( n48712 , n13278 );
not ( n48713 , n27665 );
or ( n48714 , n48712 , n48713 );
not ( n48715 , n24536 );
or ( n48716 , n48715 , n27665 );
nand ( n48717 , n48714 , n48716 );
buf ( n48718 , n48717 );
buf ( n48719 , n48718 );
buf ( n48720 , n275554 );
not ( n48721 , n275929 );
buf ( n48722 , n48721 );
buf ( n48723 , n48722 );
not ( n48724 , n275929 );
buf ( n48725 , n48724 );
buf ( n48726 , n48725 );
buf ( n48727 , n275554 );
or ( n48728 , n37497 , n28146 );
nand ( n48729 , n24450 , n18814 );
nand ( n48730 , n48728 , n48729 );
buf ( n48731 , n48730 );
buf ( n48732 , n48731 );
buf ( n48733 , n275554 );
not ( n48734 , n275925 );
buf ( n48735 , n48734 );
buf ( n48736 , n48735 );
not ( n48737 , n23759 );
not ( n48738 , n48737 );
not ( n48739 , n26373 );
and ( n48740 , n48738 , n48739 );
and ( n48741 , n23729 , n26370 );
nor ( n48742 , n48740 , n48741 );
or ( n48743 , n23787 , n26364 );
nor ( n48744 , n26386 , n37530 );
not ( n48745 , n48744 );
nand ( n48746 , n23764 , n32188 );
not ( n48747 , n26390 );
nand ( n48748 , n48747 , n37532 );
nand ( n48749 , n26395 , n23769 );
nand ( n48750 , n48745 , n48746 , n48748 , n48749 );
not ( n48751 , n48750 );
nand ( n48752 , n48742 , n48743 , n48751 );
buf ( n48753 , n48752 );
buf ( n48754 , n48753 );
not ( n48755 , n275929 );
buf ( n48756 , n48755 );
buf ( n48757 , n48756 );
buf ( n48758 , n275554 );
not ( n48759 , n275929 );
buf ( n48760 , n48759 );
buf ( n48761 , n48760 );
not ( n48762 , n275929 );
buf ( n48763 , n48762 );
buf ( n48764 , n48763 );
nand ( n48765 , n25064 , n26091 );
buf ( n48766 , n32428 );
buf ( n48767 , n25249 );
and ( n48768 , n48766 , n48767 );
buf ( n48769 , n48768 );
buf ( n48770 , n48769 );
not ( n48771 , n48770 );
buf ( n48772 , n25224 );
buf ( n48773 , n25242 );
nor ( n48774 , n48772 , n48773 );
buf ( n48775 , n48774 );
buf ( n48776 , n48775 );
not ( n48777 , n48776 );
or ( n48778 , n48771 , n48777 );
buf ( n48779 , n48775 );
buf ( n48780 , n48769 );
or ( n48781 , n48779 , n48780 );
nand ( n48782 , n48778 , n48781 );
buf ( n48783 , n48782 );
buf ( n48784 , n48783 );
not ( n48785 , n48784 );
nor ( n48786 , n48785 , n25389 );
nand ( n48787 , n25397 , n275812 );
buf ( n48788 , n32465 );
buf ( n48789 , n25571 );
nand ( n48790 , n48788 , n48789 );
buf ( n48791 , n48790 );
buf ( n48792 , n48791 );
not ( n48793 , n48792 );
buf ( n48794 , n32475 );
not ( n48795 , n48794 );
buf ( n48796 , n25543 );
nand ( n48797 , n48795 , n48796 );
buf ( n48798 , n48797 );
buf ( n48799 , n48798 );
not ( n48800 , n48799 );
or ( n48801 , n48793 , n48800 );
buf ( n48802 , n48798 );
buf ( n48803 , n48791 );
or ( n48804 , n48802 , n48803 );
nand ( n48805 , n48801 , n48804 );
buf ( n48806 , n48805 );
buf ( n48807 , n48806 );
and ( n48808 , n25402 , n48807 );
nor ( n48809 , n48808 , n41199 );
buf ( n48810 , n32509 );
buf ( n48811 , n25887 );
nand ( n48812 , n48810 , n48811 );
buf ( n48813 , n48812 );
buf ( n48814 , n48813 );
not ( n48815 , n48814 );
buf ( n48816 , n32519 );
not ( n48817 , n48816 );
buf ( n48818 , n25859 );
nand ( n48819 , n48817 , n48818 );
buf ( n48820 , n48819 );
buf ( n48821 , n48820 );
not ( n48822 , n48821 );
or ( n48823 , n48815 , n48822 );
buf ( n48824 , n48820 );
buf ( n48825 , n48813 );
or ( n48826 , n48824 , n48825 );
nand ( n48827 , n48823 , n48826 );
buf ( n48828 , n48827 );
buf ( n48829 , n48828 );
nand ( n48830 , n25717 , n48829 );
nand ( n48831 , n48787 , n48809 , n48830 );
nor ( n48832 , n48786 , n48831 );
buf ( n48833 , n26197 );
buf ( n48834 , n32552 );
nand ( n48835 , n48833 , n48834 );
buf ( n48836 , n48835 );
buf ( n48837 , n48836 );
not ( n48838 , n48837 );
buf ( n48839 , n26189 );
not ( n48840 , n48839 );
buf ( n48841 , n26169 );
nand ( n48842 , n48840 , n48841 );
buf ( n48843 , n48842 );
buf ( n48844 , n48843 );
not ( n48845 , n48844 );
or ( n48846 , n48838 , n48845 );
buf ( n48847 , n48843 );
buf ( n48848 , n48836 );
or ( n48849 , n48847 , n48848 );
nand ( n48850 , n48846 , n48849 );
buf ( n48851 , n48850 );
buf ( n48852 , n48851 );
nand ( n48853 , n26027 , n48852 );
nand ( n48854 , n48765 , n48832 , n48853 );
buf ( n48855 , n48854 );
buf ( n48856 , n48855 );
buf ( n48857 , n275554 );
and ( n48858 , n22193 , n277830 );
not ( n48859 , n22193 );
and ( n48860 , n48859 , n42684 );
or ( n48861 , n48858 , n48860 );
buf ( n48862 , n48861 );
buf ( n48863 , n48862 );
not ( n48864 , n275925 );
buf ( n48865 , n48864 );
buf ( n48866 , n48865 );
buf ( n48867 , n275554 );
buf ( n48868 , n275554 );
not ( n48869 , n275929 );
buf ( n48870 , n48869 );
buf ( n48871 , n48870 );
and ( n48872 , n31468 , n275698 );
nor ( n48873 , n48872 , n48690 );
nand ( n48874 , n22914 , n37518 );
buf ( n48875 , n23004 );
not ( n48876 , n48875 );
buf ( n48877 , n23040 );
nand ( n48878 , n48876 , n48877 );
buf ( n48879 , n48878 );
buf ( n48880 , n48879 );
not ( n48881 , n48880 );
buf ( n48882 , n23027 );
buf ( n48883 , n23034 );
nand ( n48884 , n48882 , n48883 );
buf ( n48885 , n48884 );
buf ( n48886 , n48885 );
not ( n48887 , n48886 );
or ( n48888 , n48881 , n48887 );
buf ( n48889 , n48879 );
buf ( n48890 , n48885 );
or ( n48891 , n48889 , n48890 );
nand ( n48892 , n48888 , n48891 );
buf ( n48893 , n48892 );
buf ( n48894 , n48893 );
nand ( n48895 , n22918 , n48894 );
buf ( n48896 , n23233 );
not ( n48897 , n48896 );
buf ( n48898 , n23269 );
nand ( n48899 , n48897 , n48898 );
buf ( n48900 , n48899 );
buf ( n48901 , n48900 );
not ( n48902 , n48901 );
buf ( n48903 , n23256 );
buf ( n48904 , n23263 );
nand ( n48905 , n48903 , n48904 );
buf ( n48906 , n48905 );
buf ( n48907 , n48906 );
not ( n48908 , n48907 );
or ( n48909 , n48902 , n48908 );
buf ( n48910 , n48900 );
buf ( n48911 , n48906 );
or ( n48912 , n48910 , n48911 );
nand ( n48913 , n48909 , n48912 );
buf ( n48914 , n48913 );
buf ( n48915 , n48914 );
nand ( n48916 , n23152 , n48915 );
nand ( n48917 , n48873 , n48874 , n48895 , n48916 );
buf ( n48918 , n48917 );
buf ( n48919 , n48918 );
not ( n48920 , n44919 );
and ( n48921 , n48920 , n20847 );
nand ( n48922 , n44939 , n20889 );
nand ( n48923 , n44962 , n20927 );
and ( n48924 , n44976 , n17409 );
and ( n48925 , n20940 , n44978 );
nor ( n48926 , n48924 , n48925 );
nand ( n48927 , n48922 , n48923 , n48926 );
nor ( n48928 , n48921 , n48927 );
or ( n48929 , n48928 , n20950 );
nand ( n48930 , n20953 , n13506 );
nand ( n48931 , n48929 , n48930 );
buf ( n48932 , n48931 );
buf ( n48933 , n48932 );
not ( n48934 , n275929 );
buf ( n48935 , n48934 );
buf ( n48936 , n48935 );
not ( n48937 , n275550 );
buf ( n48938 , n48937 );
buf ( n48939 , n48938 );
not ( n48940 , n275925 );
buf ( n48941 , n48940 );
buf ( n48942 , n48941 );
buf ( n48943 , n275554 );
buf ( n48944 , n275554 );
not ( n48945 , n22800 );
or ( n48946 , n48945 , n21770 );
nand ( n48947 , n21774 , n9587 );
nand ( n48948 , n48946 , n48947 );
buf ( n48949 , n48948 );
buf ( n48950 , n48949 );
not ( n48951 , n275644 );
nand ( n48952 , n48951 , n275850 );
not ( n48953 , n48952 );
not ( n48954 , n24348 );
not ( n48955 , n48954 );
or ( n48956 , n48953 , n48955 );
or ( n48957 , n48954 , n48952 );
nand ( n48958 , n48956 , n48957 );
buf ( n48959 , n48958 );
buf ( n48960 , n48959 );
buf ( n48961 , n275554 );
or ( n48962 , n36036 , n39699 );
and ( n48963 , n36047 , n36505 );
not ( n48964 , n41963 );
nor ( n48965 , n48964 , n41932 );
not ( n48966 , n48965 );
and ( n48967 , n41903 , n41922 , n41927 );
not ( n48968 , n41927 );
not ( n48969 , n41956 );
or ( n48970 , n48968 , n48969 );
nand ( n48971 , n48970 , n41960 );
nor ( n48972 , n48967 , n48971 );
not ( n48973 , n48972 );
or ( n48974 , n48966 , n48973 );
or ( n48975 , n48972 , n48965 );
nand ( n48976 , n48974 , n48975 );
buf ( n48977 , n48976 );
not ( n48978 , n48977 );
not ( n48979 , n36155 );
or ( n48980 , n48978 , n48979 );
not ( n48981 , n42062 );
nor ( n48982 , n48981 , n42030 );
not ( n48983 , n48982 );
and ( n48984 , n42002 , n42021 , n42025 );
not ( n48985 , n42025 );
not ( n48986 , n42055 );
or ( n48987 , n48985 , n48986 );
nand ( n48988 , n48987 , n42059 );
nor ( n48989 , n48984 , n48988 );
not ( n48990 , n48989 );
or ( n48991 , n48983 , n48990 );
or ( n48992 , n48989 , n48982 );
nand ( n48993 , n48991 , n48992 );
buf ( n48994 , n48993 );
nand ( n48995 , n36159 , n48994 );
nand ( n48996 , n48980 , n48995 );
nor ( n48997 , n48963 , n48996 );
nand ( n48998 , n48962 , n48997 );
nand ( n48999 , n48998 , n20645 );
not ( n49000 , n42153 );
nor ( n49001 , n49000 , n42126 );
not ( n49002 , n49001 );
and ( n49003 , n42095 , n42116 , n42121 );
not ( n49004 , n42121 );
not ( n49005 , n42146 );
or ( n49006 , n49004 , n49005 );
nand ( n49007 , n49006 , n42150 );
nor ( n49008 , n49003 , n49007 );
not ( n49009 , n49008 );
or ( n49010 , n49002 , n49009 );
or ( n49011 , n49008 , n49001 );
nand ( n49012 , n49010 , n49011 );
buf ( n49013 , n49012 );
nand ( n49014 , n36267 , n49013 );
not ( n49015 , n42238 );
nor ( n49016 , n49015 , n42211 );
not ( n49017 , n49016 );
and ( n49018 , n42181 , n42202 , n42206 );
not ( n49019 , n42206 );
not ( n49020 , n42231 );
or ( n49021 , n49019 , n49020 );
nand ( n49022 , n49021 , n42235 );
nor ( n49023 , n49018 , n49022 );
not ( n49024 , n49023 );
or ( n49025 , n49017 , n49024 );
or ( n49026 , n49023 , n49016 );
nand ( n49027 , n49025 , n49026 );
buf ( n49028 , n49027 );
nand ( n49029 , n36371 , n49028 );
and ( n49030 , n36474 , n39698 );
or ( n49031 , n20654 , n36504 );
nand ( n49032 , n49031 , n40463 );
nor ( n49033 , n49030 , n49032 );
nand ( n49034 , n48999 , n49014 , n49029 , n49033 );
buf ( n49035 , n49034 );
buf ( n49036 , n49035 );
not ( n49037 , n275925 );
buf ( n49038 , n49037 );
buf ( n49039 , n49038 );
buf ( n49040 , n275554 );
or ( n49041 , n36036 , n36571 );
and ( n49042 , n36047 , n275619 );
not ( n49043 , n36060 );
nand ( n49044 , n49043 , n45682 );
not ( n49045 , n49044 );
not ( n49046 , n36137 );
or ( n49047 , n49045 , n49046 );
or ( n49048 , n36137 , n49044 );
nand ( n49049 , n49047 , n49048 );
buf ( n49050 , n49049 );
not ( n49051 , n49050 );
not ( n49052 , n36155 );
or ( n49053 , n49051 , n49052 );
not ( n49054 , n36172 );
nand ( n49055 , n49054 , n45696 );
not ( n49056 , n49055 );
not ( n49057 , n36243 );
or ( n49058 , n49056 , n49057 );
or ( n49059 , n36243 , n49055 );
nand ( n49060 , n49058 , n49059 );
buf ( n49061 , n49060 );
nand ( n49062 , n36159 , n49061 );
nand ( n49063 , n49053 , n49062 );
nor ( n49064 , n49042 , n49063 );
nand ( n49065 , n49041 , n49064 );
nand ( n49066 , n49065 , n20645 );
not ( n49067 , n45711 );
nand ( n49068 , n49067 , n45713 );
not ( n49069 , n49068 );
not ( n49070 , n36353 );
or ( n49071 , n49069 , n49070 );
or ( n49072 , n36353 , n49068 );
nand ( n49073 , n49071 , n49072 );
buf ( n49074 , n49073 );
nand ( n49075 , n36267 , n49074 );
not ( n49076 , n45724 );
nand ( n49077 , n49076 , n36460 );
not ( n49078 , n49077 );
not ( n49079 , n36456 );
or ( n49080 , n49078 , n49079 );
or ( n49081 , n36456 , n49077 );
nand ( n49082 , n49080 , n49081 );
buf ( n49083 , n49082 );
nand ( n49084 , n36371 , n49083 );
and ( n49085 , n36474 , n11577 );
or ( n49086 , n20654 , n275618 );
nand ( n49087 , n49086 , n35906 );
nor ( n49088 , n49085 , n49087 );
nand ( n49089 , n49066 , n49075 , n49084 , n49088 );
buf ( n49090 , n49089 );
buf ( n49091 , n49090 );
not ( n49092 , n275925 );
buf ( n49093 , n49092 );
buf ( n49094 , n49093 );
not ( n49095 , n275925 );
buf ( n49096 , n49095 );
buf ( n49097 , n49096 );
not ( n49098 , n275925 );
buf ( n49099 , n49098 );
buf ( n49100 , n49099 );
not ( n49101 , n275550 );
buf ( n49102 , n49101 );
buf ( n49103 , n49102 );
not ( n49104 , n275929 );
buf ( n49105 , n49104 );
buf ( n49106 , n49105 );
not ( n49107 , n275929 );
buf ( n49108 , n49107 );
buf ( n49109 , n49108 );
buf ( n49110 , n275554 );
or ( n49111 , n30379 , n23887 );
nand ( n49112 , n20953 , n14645 );
nand ( n49113 , n49111 , n49112 );
buf ( n49114 , n49113 );
buf ( n49115 , n49114 );
not ( n49116 , n275550 );
buf ( n49117 , n49116 );
buf ( n49118 , n49117 );
buf ( n49119 , n275554 );
not ( n49120 , n275925 );
buf ( n49121 , n49120 );
buf ( n49122 , n49121 );
buf ( n49123 , n275554 );
buf ( n49124 , n275554 );
not ( n49125 , n275929 );
buf ( n49126 , n49125 );
buf ( n49127 , n49126 );
not ( n49128 , n275929 );
buf ( n49129 , n49128 );
buf ( n49130 , n49129 );
or ( n49131 , n36036 , n44996 );
and ( n49132 , n45676 , n275580 );
not ( n49133 , n41911 );
nor ( n49134 , n49133 , n41951 );
not ( n49135 , n49134 );
and ( n49136 , n47969 , n36137 , n41921 );
not ( n49137 , n41921 );
or ( n49138 , n41902 , n49137 );
not ( n49139 , n41946 );
nand ( n49140 , n49138 , n49139 );
nor ( n49141 , n49136 , n49140 );
not ( n49142 , n49141 );
or ( n49143 , n49135 , n49142 );
or ( n49144 , n49141 , n49134 );
nand ( n49145 , n49143 , n49144 );
buf ( n49146 , n49145 );
not ( n49147 , n49146 );
not ( n49148 , n36155 );
or ( n49149 , n49147 , n49148 );
not ( n49150 , n42010 );
nor ( n49151 , n49150 , n42050 );
not ( n49152 , n49151 );
and ( n49153 , n47985 , n36243 , n42020 );
not ( n49154 , n42020 );
or ( n49155 , n42001 , n49154 );
not ( n49156 , n42045 );
nand ( n49157 , n49155 , n49156 );
nor ( n49158 , n49153 , n49157 );
not ( n49159 , n49158 );
or ( n49160 , n49152 , n49159 );
or ( n49161 , n49158 , n49151 );
nand ( n49162 , n49160 , n49161 );
buf ( n49163 , n49162 );
nand ( n49164 , n36159 , n49163 );
nand ( n49165 , n49149 , n49164 );
nor ( n49166 , n49132 , n49165 );
nand ( n49167 , n49131 , n49166 );
nand ( n49168 , n49167 , n20645 );
not ( n49169 , n42142 );
nor ( n49170 , n49169 , n42114 );
not ( n49171 , n49170 );
and ( n49172 , n48004 , n36353 , n42105 );
nand ( n49173 , n42089 , n42105 );
nand ( n49174 , n49173 , n42139 );
nor ( n49175 , n49172 , n49174 );
not ( n49176 , n49175 );
or ( n49177 , n49171 , n49176 );
or ( n49178 , n49175 , n49170 );
nand ( n49179 , n49177 , n49178 );
buf ( n49180 , n49179 );
nand ( n49181 , n36267 , n49180 );
not ( n49182 , n42227 );
nor ( n49183 , n49182 , n42200 );
not ( n49184 , n49183 );
and ( n49185 , n48018 , n36456 , n42191 );
nand ( n49186 , n42175 , n42191 );
nand ( n49187 , n49186 , n42224 );
nor ( n49188 , n49185 , n49187 );
not ( n49189 , n49188 );
or ( n49190 , n49184 , n49189 );
or ( n49191 , n49188 , n49183 );
nand ( n49192 , n49190 , n49191 );
buf ( n49193 , n49192 );
nand ( n49194 , n36371 , n49193 );
and ( n49195 , n36474 , n11202 );
or ( n49196 , n20654 , n275579 );
nand ( n49197 , n49196 , n34389 );
nor ( n49198 , n49195 , n49197 );
nand ( n49199 , n49168 , n49181 , n49194 , n49198 );
buf ( n49200 , n49199 );
buf ( n49201 , n49200 );
not ( n49202 , n275925 );
buf ( n49203 , n49202 );
buf ( n49204 , n49203 );
buf ( n49205 , n275554 );
not ( n49206 , n39236 );
or ( n49207 , n49206 , n21770 );
nand ( n49208 , n21774 , n9570 );
nand ( n49209 , n49207 , n49208 );
buf ( n49210 , n49209 );
buf ( n49211 , n49210 );
nand ( n49212 , n25064 , n32873 );
buf ( n49213 , n28602 );
not ( n49214 , n49213 );
buf ( n49215 , n28556 );
nor ( n49216 , n49214 , n49215 );
buf ( n49217 , n49216 );
buf ( n49218 , n49217 );
not ( n49219 , n49218 );
buf ( n49220 , n28514 );
buf ( n49221 , n28523 );
buf ( n49222 , n28546 );
not ( n49223 , n49222 );
buf ( n49224 , n49223 );
buf ( n49225 , n49224 );
and ( n49226 , n49220 , n49221 , n49225 );
buf ( n49227 , n28573 );
buf ( n49228 , n28546 );
or ( n49229 , n49227 , n49228 );
buf ( n49230 , n28596 );
nand ( n49231 , n49229 , n49230 );
buf ( n49232 , n49231 );
buf ( n49233 , n49232 );
nor ( n49234 , n49226 , n49233 );
buf ( n49235 , n49234 );
buf ( n49236 , n49235 );
not ( n49237 , n49236 );
or ( n49238 , n49219 , n49237 );
buf ( n49239 , n49235 );
buf ( n49240 , n49217 );
or ( n49241 , n49239 , n49240 );
nand ( n49242 , n49238 , n49241 );
buf ( n49243 , n49242 );
buf ( n49244 , n49243 );
and ( n49245 , n34544 , n49244 );
not ( n49246 , n39557 );
not ( n49247 , n25396 );
or ( n49248 , n49246 , n49247 );
buf ( n49249 , n28741 );
not ( n49250 , n49249 );
buf ( n49251 , n28675 );
nor ( n49252 , n49250 , n49251 );
buf ( n49253 , n49252 );
buf ( n49254 , n49253 );
not ( n49255 , n49254 );
buf ( n49256 , n28655 );
buf ( n49257 , n28667 );
buf ( n49258 , n28694 );
and ( n49259 , n49256 , n49257 , n49258 );
buf ( n49260 , n28732 );
not ( n49261 , n49260 );
buf ( n49262 , n28714 );
not ( n49263 , n49262 );
buf ( n49264 , n28694 );
nand ( n49265 , n49263 , n49264 );
buf ( n49266 , n49265 );
buf ( n49267 , n49266 );
nand ( n49268 , n49261 , n49267 );
buf ( n49269 , n49268 );
buf ( n49270 , n49269 );
nor ( n49271 , n49259 , n49270 );
buf ( n49272 , n49271 );
buf ( n49273 , n49272 );
not ( n49274 , n49273 );
or ( n49275 , n49255 , n49274 );
buf ( n49276 , n49272 );
buf ( n49277 , n49253 );
or ( n49278 , n49276 , n49277 );
nand ( n49279 , n49275 , n49278 );
buf ( n49280 , n49279 );
buf ( n49281 , n49280 );
and ( n49282 , n25402 , n49281 );
buf ( n49283 , n28882 );
not ( n49284 , n49283 );
buf ( n49285 , n28815 );
nor ( n49286 , n49284 , n49285 );
buf ( n49287 , n49286 );
buf ( n49288 , n49287 );
not ( n49289 , n49288 );
buf ( n49290 , n28796 );
buf ( n49291 , n28808 );
buf ( n49292 , n28835 );
and ( n49293 , n49290 , n49291 , n49292 );
buf ( n49294 , n28873 );
not ( n49295 , n49294 );
buf ( n49296 , n28855 );
not ( n49297 , n49296 );
buf ( n49298 , n28835 );
nand ( n49299 , n49297 , n49298 );
buf ( n49300 , n49299 );
buf ( n49301 , n49300 );
nand ( n49302 , n49295 , n49301 );
buf ( n49303 , n49302 );
buf ( n49304 , n49303 );
nor ( n49305 , n49293 , n49304 );
buf ( n49306 , n49305 );
buf ( n49307 , n49306 );
not ( n49308 , n49307 );
or ( n49309 , n49289 , n49308 );
buf ( n49310 , n49306 );
buf ( n49311 , n49287 );
or ( n49312 , n49310 , n49311 );
nand ( n49313 , n49309 , n49312 );
buf ( n49314 , n49313 );
buf ( n49315 , n49314 );
not ( n49316 , n49315 );
not ( n49317 , n28761 );
or ( n49318 , n49316 , n49317 );
nand ( n49319 , n49318 , n42335 );
nor ( n49320 , n49282 , n49319 );
nand ( n49321 , n49248 , n49320 );
nor ( n49322 , n49245 , n49321 );
buf ( n49323 , n29021 );
not ( n49324 , n49323 );
buf ( n49325 , n28975 );
nor ( n49326 , n49324 , n49325 );
buf ( n49327 , n49326 );
buf ( n49328 , n49327 );
not ( n49329 , n49328 );
buf ( n49330 , n28935 );
buf ( n49331 , n28947 );
buf ( n49332 , n28967 );
not ( n49333 , n49332 );
buf ( n49334 , n49333 );
buf ( n49335 , n49334 );
and ( n49336 , n49330 , n49331 , n49335 );
buf ( n49337 , n28992 );
buf ( n49338 , n28967 );
or ( n49339 , n49337 , n49338 );
buf ( n49340 , n29015 );
nand ( n49341 , n49339 , n49340 );
buf ( n49342 , n49341 );
buf ( n49343 , n49342 );
nor ( n49344 , n49336 , n49343 );
buf ( n49345 , n49344 );
buf ( n49346 , n49345 );
not ( n49347 , n49346 );
or ( n49348 , n49329 , n49347 );
buf ( n49349 , n49345 );
buf ( n49350 , n49327 );
or ( n49351 , n49349 , n49350 );
nand ( n49352 , n49348 , n49351 );
buf ( n49353 , n49352 );
buf ( n49354 , n49353 );
nand ( n49355 , n26027 , n49354 );
nand ( n49356 , n49212 , n49322 , n49355 );
buf ( n49357 , n49356 );
buf ( n49358 , n49357 );
buf ( n49359 , n275554 );
nand ( n49360 , n34811 , n31422 );
nand ( n49361 , n34837 , n28330 );
nand ( n49362 , n34844 , n31449 );
and ( n49363 , n32054 , n277554 );
not ( n49364 , n277573 );
not ( n49365 , n28357 );
or ( n49366 , n49364 , n49365 );
or ( n49367 , n32061 , n277564 );
nand ( n49368 , n49366 , n49367 );
nor ( n49369 , n49363 , n49368 );
nand ( n49370 , n31460 , n277609 );
and ( n49371 , n49362 , n49369 , n49370 );
nand ( n49372 , n49360 , n49361 , n49371 );
buf ( n49373 , n49372 );
buf ( n49374 , n49373 );
not ( n49375 , n275550 );
buf ( n49376 , n49375 );
buf ( n49377 , n49376 );
not ( n49378 , n10841 );
or ( n49379 , n36036 , n49378 );
and ( n49380 , n45676 , n275792 );
not ( n49381 , n36073 );
nand ( n49382 , n49381 , n36105 );
not ( n49383 , n49382 );
not ( n49384 , n36135 );
or ( n49385 , n49383 , n49384 );
or ( n49386 , n36135 , n49382 );
nand ( n49387 , n49385 , n49386 );
buf ( n49388 , n49387 );
not ( n49389 , n49388 );
not ( n49390 , n36155 );
or ( n49391 , n49389 , n49390 );
not ( n49392 , n36184 );
nand ( n49393 , n49392 , n36213 );
not ( n49394 , n49393 );
not ( n49395 , n36241 );
or ( n49396 , n49394 , n49395 );
or ( n49397 , n36241 , n49393 );
nand ( n49398 , n49396 , n49397 );
buf ( n49399 , n49398 );
nand ( n49400 , n41635 , n49399 );
nand ( n49401 , n49391 , n49400 );
nor ( n49402 , n49380 , n49401 );
nand ( n49403 , n49379 , n49402 );
nand ( n49404 , n49403 , n20645 );
not ( n49405 , n36336 );
nand ( n49406 , n49405 , n36330 );
not ( n49407 , n49406 );
not ( n49408 , n36322 );
not ( n49409 , n49408 );
or ( n49410 , n49407 , n49409 );
or ( n49411 , n49408 , n49406 );
nand ( n49412 , n49410 , n49411 );
buf ( n49413 , n49412 );
nand ( n49414 , n36267 , n49413 );
not ( n49415 , n36439 );
nand ( n49416 , n49415 , n36433 );
not ( n49417 , n49416 );
not ( n49418 , n36425 );
not ( n49419 , n49418 );
or ( n49420 , n49417 , n49419 );
or ( n49421 , n49418 , n49416 );
nand ( n49422 , n49420 , n49421 );
buf ( n49423 , n49422 );
nand ( n49424 , n36371 , n49423 );
and ( n49425 , n36474 , n10841 );
or ( n49426 , n20654 , n275791 );
nand ( n49427 , n49426 , n29177 );
nor ( n49428 , n49425 , n49427 );
nand ( n49429 , n49404 , n49414 , n49424 , n49428 );
buf ( n49430 , n49429 );
buf ( n49431 , n49430 );
not ( n49432 , n275925 );
buf ( n49433 , n49432 );
buf ( n49434 , n49433 );
not ( n49435 , n275925 );
buf ( n49436 , n49435 );
buf ( n49437 , n49436 );
not ( n49438 , n275929 );
buf ( n49439 , n49438 );
buf ( n49440 , n49439 );
not ( n49441 , n275925 );
buf ( n49442 , n49441 );
buf ( n49443 , n49442 );
nand ( n49444 , n39378 , n31422 );
nand ( n49445 , n39399 , n28330 );
nand ( n49446 , n39412 , n31449 );
and ( n49447 , n36530 , n12247 );
not ( n49448 , n277868 );
not ( n49449 , n28357 );
or ( n49450 , n49448 , n49449 );
or ( n49451 , n32061 , n277853 );
nand ( n49452 , n49450 , n49451 );
nor ( n49453 , n49447 , n49452 );
nand ( n49454 , n31460 , n12182 );
and ( n49455 , n49446 , n49453 , n49454 );
nand ( n49456 , n49444 , n49445 , n49455 );
buf ( n49457 , n49456 );
buf ( n49458 , n49457 );
xor ( n49459 , n275742 , n275753 );
xor ( n49460 , n49459 , n275756 );
buf ( n49461 , n49460 );
buf ( n49462 , n49461 );
not ( n49463 , n275929 );
buf ( n49464 , n49463 );
buf ( n49465 , n49464 );
buf ( n49466 , n275554 );
buf ( n49467 , n275554 );
buf ( n49468 , n275554 );
not ( n49469 , n275925 );
buf ( n49470 , n49469 );
buf ( n49471 , n49470 );
buf ( n49472 , n275554 );
or ( n49473 , n32366 , n20743 );
nand ( n49474 , n32380 , n16968 );
nand ( n49475 , n32393 , n20763 );
nand ( n49476 , n17411 , n32401 );
nand ( n49477 , n17502 , n32405 );
nand ( n49478 , n17560 , n13611 );
nand ( n49479 , n17545 , n35756 );
and ( n49480 , n49476 , n49477 , n49478 , n49479 );
and ( n49481 , n49474 , n49475 , n49480 );
nand ( n49482 , n49473 , n49481 );
buf ( n49483 , n49482 );
buf ( n49484 , n49483 );
buf ( n49485 , n275554 );
not ( n49486 , n275929 );
buf ( n49487 , n49486 );
buf ( n49488 , n49487 );
or ( n49489 , n27742 , n27647 );
nand ( n49490 , n21696 , n13724 );
nand ( n49491 , n49489 , n49490 );
buf ( n49492 , n49491 );
buf ( n49493 , n49492 );
not ( n49494 , n275929 );
buf ( n49495 , n49494 );
buf ( n49496 , n49495 );
not ( n49497 , n275929 );
buf ( n49498 , n49497 );
buf ( n49499 , n49498 );
not ( n49500 , n275550 );
buf ( n49501 , n49500 );
buf ( n49502 , n49501 );
not ( n49503 , n31140 );
or ( n49504 , n49503 , n29046 );
nand ( n49505 , n28252 , n9523 );
nand ( n49506 , n49504 , n49505 );
buf ( n49507 , n49506 );
buf ( n49508 , n49507 );
not ( n49509 , n37860 );
or ( n49510 , n49509 , n28252 );
nand ( n49511 , n28252 , n9583 );
nand ( n49512 , n49510 , n49511 );
buf ( n49513 , n49512 );
buf ( n49514 , n49513 );
buf ( n49515 , n275554 );
buf ( n49516 , n275554 );
or ( n49517 , n23452 , n21697 );
nand ( n49518 , n21696 , n13750 );
nand ( n49519 , n49517 , n49518 );
buf ( n49520 , n49519 );
buf ( n49521 , n49520 );
buf ( n49522 , n275554 );
buf ( n49523 , n275554 );
not ( n49524 , n275929 );
buf ( n49525 , n49524 );
buf ( n49526 , n49525 );
not ( n49527 , n275550 );
buf ( n49528 , n49527 );
buf ( n49529 , n49528 );
or ( n49530 , n40356 , n32074 );
and ( n49531 , n40406 , n20515 );
not ( n49532 , n48502 );
not ( n49533 , n49532 );
not ( n49534 , n30612 );
or ( n49535 , n49533 , n49534 );
nand ( n49536 , n40421 , n31095 );
nand ( n49537 , n20563 , n40409 );
nand ( n49538 , n30179 , n18525 );
and ( n49539 , n49536 , n49537 , n49538 );
nand ( n49540 , n49535 , n49539 );
nor ( n49541 , n49531 , n49540 );
nand ( n49542 , n40383 , n20353 );
and ( n49543 , n49541 , n49542 );
nand ( n49544 , n49530 , n49543 );
buf ( n49545 , n49544 );
buf ( n49546 , n49545 );
not ( n49547 , n275925 );
buf ( n49548 , n49547 );
buf ( n49549 , n49548 );
nand ( n49550 , n40755 , n29599 );
nand ( n49551 , n40774 , n30962 );
and ( n49552 , n40785 , n22052 );
and ( n49553 , n27520 , n40787 );
and ( n49554 , n22013 , n277411 );
nor ( n49555 , n49553 , n49554 );
not ( n49556 , n49555 );
nor ( n49557 , n49552 , n49556 );
and ( n49558 , n49550 , n49551 , n49557 );
or ( n49559 , n49558 , n27179 );
not ( n49560 , n277376 );
or ( n49561 , n37463 , n49560 );
nand ( n49562 , n49559 , n49561 );
buf ( n49563 , n49562 );
buf ( n49564 , n49563 );
not ( n49565 , n275550 );
buf ( n49566 , n49565 );
buf ( n49567 , n49566 );
buf ( n49568 , n275554 );
not ( n49569 , n32980 );
or ( n49570 , n49569 , n28252 );
nand ( n49571 , n29046 , n9667 );
nand ( n49572 , n49570 , n49571 );
buf ( n49573 , n49572 );
buf ( n49574 , n49573 );
and ( n49575 , n31719 , n277966 );
not ( n49576 , n31719 );
and ( n49577 , n49576 , n29773 );
or ( n49578 , n49575 , n49577 );
buf ( n49579 , n49578 );
buf ( n49580 , n49579 );
not ( n49581 , n21772 );
not ( n49582 , n30599 );
or ( n49583 , n49581 , n49582 );
nand ( n49584 , n21773 , n9462 );
nand ( n49585 , n49583 , n49584 );
buf ( n49586 , n49585 );
buf ( n49587 , n49586 );
or ( n49588 , n32354 , n29044 );
nand ( n49589 , n29044 , n9513 );
nand ( n49590 , n49588 , n49589 );
buf ( n49591 , n49590 );
buf ( n49592 , n49591 );
buf ( n49593 , n275554 );
not ( n49594 , n22335 );
not ( n49595 , n41763 );
or ( n49596 , n49594 , n49595 );
not ( n49597 , n19927 );
or ( n49598 , n49597 , n22335 );
nand ( n49599 , n49596 , n49598 );
buf ( n49600 , n49599 );
buf ( n49601 , n49600 );
not ( n49602 , n275925 );
buf ( n49603 , n49602 );
buf ( n49604 , n49603 );
and ( n49605 , n37271 , n39553 );
nor ( n49606 , n49605 , n48744 );
nand ( n49607 , n22914 , n38188 );
buf ( n49608 , n38221 );
not ( n49609 , n49608 );
buf ( n49610 , n38195 );
nor ( n49611 , n49609 , n49610 );
buf ( n49612 , n49611 );
buf ( n49613 , n49612 );
not ( n49614 , n49613 );
buf ( n49615 , n23140 );
buf ( n49616 , n37305 );
buf ( n49617 , n38186 );
not ( n49618 , n49617 );
buf ( n49619 , n49618 );
buf ( n49620 , n49619 );
and ( n49621 , n49615 , n49616 , n49620 );
buf ( n49622 , n37330 );
buf ( n49623 , n38186 );
or ( n49624 , n49622 , n49623 );
buf ( n49625 , n38215 );
nand ( n49626 , n49624 , n49625 );
buf ( n49627 , n49626 );
buf ( n49628 , n49627 );
nor ( n49629 , n49621 , n49628 );
buf ( n49630 , n49629 );
buf ( n49631 , n49630 );
not ( n49632 , n49631 );
or ( n49633 , n49614 , n49632 );
buf ( n49634 , n49630 );
buf ( n49635 , n49612 );
or ( n49636 , n49634 , n49635 );
nand ( n49637 , n49633 , n49636 );
buf ( n49638 , n49637 );
buf ( n49639 , n49638 );
nand ( n49640 , n22918 , n49639 );
buf ( n49641 , n38290 );
not ( n49642 , n49641 );
buf ( n49643 , n38264 );
nor ( n49644 , n49642 , n49643 );
buf ( n49645 , n49644 );
buf ( n49646 , n49645 );
not ( n49647 , n49646 );
buf ( n49648 , n23365 );
buf ( n49649 , n37381 );
buf ( n49650 , n38257 );
not ( n49651 , n49650 );
buf ( n49652 , n49651 );
buf ( n49653 , n49652 );
and ( n49654 , n49648 , n49649 , n49653 );
buf ( n49655 , n37405 );
buf ( n49656 , n38257 );
or ( n49657 , n49655 , n49656 );
buf ( n49658 , n38284 );
nand ( n49659 , n49657 , n49658 );
buf ( n49660 , n49659 );
buf ( n49661 , n49660 );
nor ( n49662 , n49654 , n49661 );
buf ( n49663 , n49662 );
buf ( n49664 , n49663 );
not ( n49665 , n49664 );
or ( n49666 , n49647 , n49665 );
buf ( n49667 , n49663 );
buf ( n49668 , n49645 );
or ( n49669 , n49667 , n49668 );
nand ( n49670 , n49666 , n49669 );
buf ( n49671 , n49670 );
buf ( n49672 , n49671 );
nand ( n49673 , n23152 , n49672 );
nand ( n49674 , n49606 , n49607 , n49640 , n49673 );
buf ( n49675 , n49674 );
buf ( n49676 , n49675 );
and ( n49677 , n20961 , n9466 );
not ( n49678 , n20961 );
and ( n49679 , n49678 , n14564 );
or ( n49680 , n49677 , n49679 );
buf ( n49681 , n49680 );
buf ( n49682 , n49681 );
buf ( n49683 , n275554 );
buf ( n49684 , n275554 );
buf ( n49685 , n275554 );
not ( n49686 , n10907 );
not ( n49687 , n23708 );
or ( n49688 , n49686 , n49687 );
or ( n49689 , n45336 , n23705 );
nand ( n49690 , n49688 , n49689 );
buf ( n49691 , n49690 );
buf ( n49692 , n49691 );
and ( n49693 , n45327 , n28408 );
or ( n49694 , n28454 , n12261 );
or ( n49695 , n32757 , n12266 );
nand ( n49696 , n20649 , n9281 );
nand ( n49697 , n49694 , n49695 , n49696 );
nor ( n49698 , n49693 , n49697 );
nand ( n49699 , n45288 , n29163 );
nand ( n49700 , n45301 , n32751 );
not ( n49701 , n28450 );
nand ( n49702 , n49701 , n10917 );
nand ( n49703 , n49698 , n49699 , n49700 , n49702 );
buf ( n49704 , n49703 );
buf ( n49705 , n49704 );
not ( n49706 , n275929 );
buf ( n49707 , n49706 );
buf ( n49708 , n49707 );
or ( n49709 , n34696 , n14908 );
nand ( n49710 , n32339 , n34734 );
nand ( n49711 , n20785 , n34723 );
not ( n49712 , n17561 );
not ( n49713 , n13545 );
not ( n49714 , n49713 );
and ( n49715 , n49712 , n49714 );
and ( n49716 , n17405 , n34717 );
nor ( n49717 , n49715 , n49716 );
and ( n49718 , n34706 , n16968 );
nor ( n49719 , n20765 , n13555 );
nor ( n49720 , n49718 , n49719 );
and ( n49721 , n49710 , n49711 , n49717 , n49720 );
nand ( n49722 , n49709 , n49721 );
buf ( n49723 , n49722 );
buf ( n49724 , n49723 );
buf ( n49725 , n275554 );
buf ( n49726 , n275554 );
buf ( n49727 , n275554 );
buf ( n49728 , n275554 );
buf ( n49729 , n275554 );
not ( n49730 , n275925 );
buf ( n49731 , n49730 );
buf ( n49732 , n49731 );
nand ( n49733 , n42653 , n31422 );
nand ( n49734 , n42667 , n31437 );
nand ( n49735 , n42676 , n31449 );
and ( n49736 , n36530 , n11826 );
not ( n49737 , n277839 );
not ( n49738 , n28236 );
or ( n49739 , n49737 , n49738 );
or ( n49740 , n31453 , n277826 );
nand ( n49741 , n49739 , n49740 );
nor ( n49742 , n49736 , n49741 );
nand ( n49743 , n31460 , n12248 );
and ( n49744 , n49735 , n49742 , n49743 );
nand ( n49745 , n49733 , n49734 , n49744 );
buf ( n49746 , n49745 );
buf ( n49747 , n49746 );
buf ( n49748 , n275554 );
not ( n49749 , n275925 );
buf ( n49750 , n49749 );
buf ( n49751 , n49750 );
not ( n49752 , n23822 );
or ( n49753 , n49752 , n28252 );
nand ( n49754 , n28252 , n9684 );
nand ( n49755 , n49753 , n49754 );
buf ( n49756 , n49755 );
buf ( n49757 , n49756 );
buf ( n49758 , n275554 );
buf ( n49759 , n275554 );
not ( n49760 , n275925 );
buf ( n49761 , n49760 );
buf ( n49762 , n49761 );
not ( n49763 , n275925 );
buf ( n49764 , n49763 );
buf ( n49765 , n49764 );
buf ( n49766 , n275554 );
buf ( n49767 , n275554 );
not ( n49768 , n41925 );
or ( n49769 , n36036 , n49768 );
and ( n49770 , n36047 , n31691 );
and ( n49771 , n41960 , n41927 );
not ( n49772 , n49771 );
and ( n49773 , n41922 , n47969 , n36137 );
not ( n49774 , n41956 );
nand ( n49775 , n41922 , n41901 );
nand ( n49776 , n49774 , n49775 );
nor ( n49777 , n49773 , n49776 );
not ( n49778 , n49777 );
or ( n49779 , n49772 , n49778 );
or ( n49780 , n49777 , n49771 );
nand ( n49781 , n49779 , n49780 );
buf ( n49782 , n49781 );
not ( n49783 , n49782 );
not ( n49784 , n36155 );
or ( n49785 , n49783 , n49784 );
and ( n49786 , n42059 , n42025 );
not ( n49787 , n49786 );
and ( n49788 , n42021 , n47985 , n36243 );
not ( n49789 , n42000 );
not ( n49790 , n42021 );
or ( n49791 , n49789 , n49790 );
not ( n49792 , n42055 );
nand ( n49793 , n49791 , n49792 );
nor ( n49794 , n49788 , n49793 );
not ( n49795 , n49794 );
or ( n49796 , n49787 , n49795 );
or ( n49797 , n49794 , n49786 );
nand ( n49798 , n49796 , n49797 );
buf ( n49799 , n49798 );
nand ( n49800 , n36159 , n49799 );
nand ( n49801 , n49785 , n49800 );
nor ( n49802 , n49770 , n49801 );
nand ( n49803 , n49769 , n49802 );
nand ( n49804 , n49803 , n20645 );
and ( n49805 , n42121 , n42150 );
not ( n49806 , n49805 );
and ( n49807 , n42116 , n48004 , n36353 );
not ( n49808 , n42146 );
nand ( n49809 , n42116 , n42089 );
nand ( n49810 , n49808 , n49809 );
nor ( n49811 , n49807 , n49810 );
not ( n49812 , n49811 );
or ( n49813 , n49806 , n49812 );
or ( n49814 , n49811 , n49805 );
nand ( n49815 , n49813 , n49814 );
buf ( n49816 , n49815 );
nand ( n49817 , n36267 , n49816 );
and ( n49818 , n42206 , n42235 );
not ( n49819 , n49818 );
and ( n49820 , n42202 , n48018 , n36456 );
not ( n49821 , n42231 );
nand ( n49822 , n42202 , n42175 );
nand ( n49823 , n49821 , n49822 );
nor ( n49824 , n49820 , n49823 );
not ( n49825 , n49824 );
or ( n49826 , n49819 , n49825 );
or ( n49827 , n49824 , n49818 );
nand ( n49828 , n49826 , n49827 );
buf ( n49829 , n49828 );
nand ( n49830 , n36371 , n49829 );
and ( n49831 , n36474 , n41925 );
or ( n49832 , n20654 , n31690 );
nand ( n49833 , n49832 , n45414 );
nor ( n49834 , n49831 , n49833 );
nand ( n49835 , n49804 , n49817 , n49830 , n49834 );
buf ( n49836 , n49835 );
buf ( n49837 , n49836 );
and ( n49838 , n21696 , n14739 );
not ( n49839 , n21696 );
and ( n49840 , n49839 , n38856 );
or ( n49841 , n49838 , n49840 );
buf ( n49842 , n49841 );
buf ( n49843 , n49842 );
not ( n49844 , n275929 );
buf ( n49845 , n49844 );
buf ( n49846 , n49845 );
or ( n49847 , n36036 , n36994 );
and ( n49848 , n36047 , n275566 );
not ( n49849 , n41907 );
nor ( n49850 , n49849 , n41954 );
not ( n49851 , n49850 );
nand ( n49852 , n41921 , n41911 );
not ( n49853 , n49852 );
and ( n49854 , n47969 , n36137 , n49853 );
or ( n49855 , n41902 , n49852 );
and ( n49856 , n41946 , n41911 );
nor ( n49857 , n49856 , n41951 );
nand ( n49858 , n49855 , n49857 );
nor ( n49859 , n49854 , n49858 );
not ( n49860 , n49859 );
or ( n49861 , n49851 , n49860 );
or ( n49862 , n49859 , n49850 );
nand ( n49863 , n49861 , n49862 );
buf ( n49864 , n49863 );
not ( n49865 , n49864 );
not ( n49866 , n36155 );
or ( n49867 , n49865 , n49866 );
not ( n49868 , n42006 );
nor ( n49869 , n49868 , n42053 );
not ( n49870 , n49869 );
nand ( n49871 , n42020 , n42010 );
not ( n49872 , n49871 );
and ( n49873 , n47985 , n36243 , n49872 );
or ( n49874 , n42001 , n49871 );
and ( n49875 , n42045 , n42010 );
nor ( n49876 , n49875 , n42050 );
nand ( n49877 , n49874 , n49876 );
nor ( n49878 , n49873 , n49877 );
not ( n49879 , n49878 );
or ( n49880 , n49870 , n49879 );
or ( n49881 , n49878 , n49869 );
nand ( n49882 , n49880 , n49881 );
buf ( n49883 , n49882 );
nand ( n49884 , n36159 , n49883 );
nand ( n49885 , n49867 , n49884 );
nor ( n49886 , n49848 , n49885 );
nand ( n49887 , n49847 , n49886 );
nand ( n49888 , n49887 , n20645 );
not ( n49889 , n42145 );
nor ( n49890 , n49889 , n42110 );
not ( n49891 , n49890 );
nor ( n49892 , n42104 , n42114 );
and ( n49893 , n48004 , n36353 , n49892 );
or ( n49894 , n42139 , n42114 );
nand ( n49895 , n42089 , n49892 );
nand ( n49896 , n49894 , n49895 , n42142 );
nor ( n49897 , n49893 , n49896 );
not ( n49898 , n49897 );
or ( n49899 , n49891 , n49898 );
or ( n49900 , n49897 , n49890 );
nand ( n49901 , n49899 , n49900 );
buf ( n49902 , n49901 );
nand ( n49903 , n36267 , n49902 );
not ( n49904 , n42230 );
nor ( n49905 , n49904 , n42196 );
not ( n49906 , n49905 );
nor ( n49907 , n42190 , n42200 );
and ( n49908 , n48018 , n36456 , n49907 );
or ( n49909 , n42224 , n42200 );
nand ( n49910 , n42175 , n49907 );
nand ( n49911 , n49909 , n49910 , n42227 );
nor ( n49912 , n49908 , n49911 );
not ( n49913 , n49912 );
or ( n49914 , n49906 , n49913 );
or ( n49915 , n49912 , n49905 );
nand ( n49916 , n49914 , n49915 );
buf ( n49917 , n49916 );
nand ( n49918 , n36371 , n49917 );
and ( n49919 , n36474 , n11302 );
or ( n49920 , n20654 , n275565 );
nand ( n49921 , n49920 , n35101 );
nor ( n49922 , n49919 , n49921 );
nand ( n49923 , n49888 , n49903 , n49918 , n49922 );
buf ( n49924 , n49923 );
buf ( n49925 , n49924 );
not ( n49926 , n275929 );
buf ( n49927 , n49926 );
buf ( n49928 , n49927 );
not ( n49929 , n275550 );
buf ( n49930 , n49929 );
buf ( n49931 , n49930 );
or ( n49932 , n27624 , n28146 );
nand ( n49933 , n24452 , n18770 );
nand ( n49934 , n49932 , n49933 );
buf ( n49935 , n49934 );
buf ( n49936 , n49935 );
or ( n49937 , n36986 , n21030 );
nand ( n49938 , n21030 , n18364 );
nand ( n49939 , n49937 , n49938 );
buf ( n49940 , n49939 );
buf ( n49941 , n49940 );
not ( n49942 , n275550 );
buf ( n49943 , n49942 );
buf ( n49944 , n49943 );
nand ( n49945 , n37066 , n28306 );
nand ( n49946 , n37079 , n31437 );
nand ( n49947 , n37083 , n31449 );
and ( n49948 , n31451 , n12288 );
not ( n49949 , n278015 );
or ( n49950 , n28354 , n49949 );
nand ( n49951 , n28236 , n278022 );
nand ( n49952 , n49950 , n49951 );
nor ( n49953 , n49948 , n49952 );
nand ( n49954 , n31460 , n12295 );
and ( n49955 , n49947 , n49953 , n49954 );
nand ( n49956 , n49945 , n49946 , n49955 );
buf ( n49957 , n49956 );
buf ( n49958 , n49957 );
buf ( n49959 , n275554 );
or ( n49960 , n32409 , n20953 );
nand ( n49961 , n20953 , n13620 );
nand ( n49962 , n49960 , n49961 );
buf ( n49963 , n49962 );
buf ( n49964 , n49963 );
not ( n49965 , n275550 );
buf ( n49966 , n49965 );
buf ( n49967 , n49966 );
buf ( n49968 , n275554 );
and ( n49969 , n27664 , n16718 );
not ( n49970 , n27664 );
and ( n49971 , n49970 , n29258 );
or ( n49972 , n49969 , n49971 );
buf ( n49973 , n49972 );
buf ( n49974 , n49973 );
or ( n49975 , n22143 , n23708 );
nand ( n49976 , n27641 , n10780 );
nand ( n49977 , n49975 , n49976 );
buf ( n49978 , n49977 );
buf ( n49979 , n49978 );
not ( n49980 , n10858 );
or ( n49981 , n9158 , n49980 );
or ( n49982 , n9157 , n49378 );
nand ( n49983 , n49981 , n49982 );
buf ( n49984 , n49983 );
buf ( n49985 , n49984 );
buf ( n49986 , n275554 );
or ( n49987 , n49558 , n40576 );
not ( n49988 , n277381 );
or ( n49989 , n22192 , n49988 );
nand ( n49990 , n49987 , n49989 );
buf ( n49991 , n49990 );
buf ( n49992 , n49991 );
not ( n49993 , n34302 );
not ( n49994 , n42796 );
or ( n49995 , n49993 , n49994 );
and ( n49996 , n42819 , n35900 );
nand ( n49997 , n42829 , n34307 );
nand ( n49998 , n28451 , n277715 );
nand ( n49999 , n29171 , n12371 );
and ( n50000 , n34311 , n12304 );
and ( n50001 , n34313 , n9341 );
nor ( n50002 , n50000 , n50001 );
and ( n50003 , n49999 , n50002 );
nand ( n50004 , n49997 , n49998 , n50003 );
nor ( n50005 , n49996 , n50004 );
nand ( n50006 , n49995 , n50005 );
buf ( n50007 , n50006 );
buf ( n50008 , n50007 );
buf ( n50009 , n275554 );
buf ( n50010 , n275554 );
buf ( n50011 , n275554 );
not ( n50012 , n275550 );
buf ( n50013 , n50012 );
buf ( n50014 , n50013 );
buf ( n50015 , n275554 );
or ( n50016 , n41396 , n21030 );
or ( n50017 , n21029 , n18837 );
nand ( n50018 , n50016 , n50017 );
buf ( n50019 , n50018 );
buf ( n50020 , n50019 );
buf ( n50021 , n275554 );
buf ( n50022 , n275554 );
buf ( n50023 , n275554 );
and ( n50024 , n31468 , n275821 );
nor ( n50025 , n50024 , n45480 );
nand ( n50026 , n22914 , n22944 );
buf ( n50027 , n22950 );
buf ( n50028 , n40254 );
nand ( n50029 , n50027 , n50028 );
buf ( n50030 , n50029 );
buf ( n50031 , n50030 );
not ( n50032 , n50031 );
buf ( n50033 , n22984 );
not ( n50034 , n50033 );
buf ( n50035 , n23046 );
nand ( n50036 , n50034 , n50035 );
buf ( n50037 , n50036 );
buf ( n50038 , n50037 );
not ( n50039 , n50038 );
or ( n50040 , n50032 , n50039 );
buf ( n50041 , n50037 );
buf ( n50042 , n50030 );
or ( n50043 , n50041 , n50042 );
nand ( n50044 , n50040 , n50043 );
buf ( n50045 , n50044 );
buf ( n50046 , n50045 );
nand ( n50047 , n22918 , n50046 );
buf ( n50048 , n23182 );
buf ( n50049 , n40289 );
nand ( n50050 , n50048 , n50049 );
buf ( n50051 , n50050 );
buf ( n50052 , n50051 );
not ( n50053 , n50052 );
buf ( n50054 , n23214 );
not ( n50055 , n50054 );
buf ( n50056 , n23275 );
nand ( n50057 , n50055 , n50056 );
buf ( n50058 , n50057 );
buf ( n50059 , n50058 );
not ( n50060 , n50059 );
or ( n50061 , n50053 , n50060 );
buf ( n50062 , n50058 );
buf ( n50063 , n50051 );
or ( n50064 , n50062 , n50063 );
nand ( n50065 , n50061 , n50064 );
buf ( n50066 , n50065 );
buf ( n50067 , n50066 );
nand ( n50068 , n23152 , n50067 );
nand ( n50069 , n50025 , n50026 , n50047 , n50068 );
buf ( n50070 , n50069 );
buf ( n50071 , n50070 );
buf ( n50072 , n275554 );
buf ( n50073 , n275554 );
not ( n50074 , n275929 );
buf ( n50075 , n50074 );
buf ( n50076 , n50075 );
not ( n50077 , n275550 );
buf ( n50078 , n50077 );
buf ( n50079 , n50078 );
not ( n50080 , n275550 );
buf ( n50081 , n50080 );
buf ( n50082 , n50081 );
not ( n50083 , n275925 );
buf ( n50084 , n50083 );
buf ( n50085 , n50084 );
buf ( n50086 , n275554 );
not ( n50087 , n275929 );
buf ( n50088 , n50087 );
buf ( n50089 , n50088 );
not ( n50090 , n275550 );
buf ( n50091 , n50090 );
buf ( n50092 , n50091 );
and ( n50093 , n22335 , n18038 );
not ( n50094 , n22335 );
and ( n50095 , n50094 , n30017 );
or ( n50096 , n50093 , n50095 );
buf ( n50097 , n50096 );
buf ( n50098 , n50097 );
or ( n50099 , n36036 , n26408 );
and ( n50100 , n45676 , n275638 );
and ( n50101 , n36088 , n36101 );
not ( n50102 , n50101 );
and ( n50103 , n36106 , n36135 , n36092 );
not ( n50104 , n36083 );
or ( n50105 , n50104 , n36073 );
nand ( n50106 , n50105 , n36079 );
not ( n50107 , n50106 );
nand ( n50108 , n50107 , n36092 );
not ( n50109 , n36097 );
nand ( n50110 , n50108 , n50109 );
nor ( n50111 , n50103 , n50110 );
not ( n50112 , n50111 );
or ( n50113 , n50102 , n50112 );
or ( n50114 , n50111 , n50101 );
nand ( n50115 , n50113 , n50114 );
buf ( n50116 , n50115 );
not ( n50117 , n50116 );
not ( n50118 , n36155 );
or ( n50119 , n50117 , n50118 );
not ( n50120 , n36198 );
nor ( n50121 , n50120 , n36209 );
not ( n50122 , n50121 );
and ( n50123 , n36214 , n36241 , n36202 );
not ( n50124 , n36193 );
or ( n50125 , n50124 , n36184 );
nand ( n50126 , n50125 , n36189 );
not ( n50127 , n50126 );
nand ( n50128 , n50127 , n36202 );
not ( n50129 , n36206 );
nand ( n50130 , n50128 , n50129 );
nor ( n50131 , n50123 , n50130 );
not ( n50132 , n50131 );
or ( n50133 , n50122 , n50132 );
or ( n50134 , n50131 , n50121 );
nand ( n50135 , n50133 , n50134 );
buf ( n50136 , n50135 );
nand ( n50137 , n41635 , n50136 );
nand ( n50138 , n50119 , n50137 );
nor ( n50139 , n50100 , n50138 );
nand ( n50140 , n50099 , n50139 );
nand ( n50141 , n50140 , n20645 );
and ( n50142 , n36350 , n36290 );
not ( n50143 , n50142 );
and ( n50144 , n36342 , n36294 );
not ( n50145 , n36294 );
nor ( n50146 , n36322 , n36331 , n50145 );
nor ( n50147 , n50144 , n50146 , n36345 );
not ( n50148 , n50147 );
or ( n50149 , n50143 , n50148 );
or ( n50150 , n50147 , n50142 );
nand ( n50151 , n50149 , n50150 );
buf ( n50152 , n50151 );
nand ( n50153 , n36267 , n50152 );
and ( n50154 , n36453 , n36394 );
not ( n50155 , n50154 );
and ( n50156 , n36445 , n36398 );
not ( n50157 , n36398 );
nor ( n50158 , n36425 , n36434 , n50157 );
nor ( n50159 , n50156 , n50158 , n36448 );
not ( n50160 , n50159 );
or ( n50161 , n50155 , n50160 );
or ( n50162 , n50159 , n50154 );
nand ( n50163 , n50161 , n50162 );
buf ( n50164 , n50163 );
nand ( n50165 , n36371 , n50164 );
and ( n50166 , n36474 , n26407 );
or ( n50167 , n20654 , n275637 );
nand ( n50168 , n50167 , n40083 );
nor ( n50169 , n50166 , n50168 );
nand ( n50170 , n50141 , n50153 , n50165 , n50169 );
buf ( n50171 , n50170 );
buf ( n50172 , n50171 );
not ( n50173 , n45327 );
not ( n50174 , n50173 );
not ( n50175 , n28304 );
and ( n50176 , n50174 , n50175 );
and ( n50177 , n45301 , n28328 );
nor ( n50178 , n50176 , n50177 );
and ( n50179 , n45288 , n37665 );
nor ( n50180 , n28241 , n12266 );
nor ( n50181 , n50179 , n50180 );
and ( n50182 , n31451 , n12236 );
not ( n50183 , n10917 );
not ( n50184 , n28236 );
or ( n50185 , n50183 , n50184 );
not ( n50186 , n10902 );
or ( n50187 , n31453 , n50186 );
nand ( n50188 , n50185 , n50187 );
nor ( n50189 , n50182 , n50188 );
nand ( n50190 , n50178 , n50181 , n50189 );
buf ( n50191 , n50190 );
buf ( n50192 , n50191 );
not ( n50193 , n275925 );
buf ( n50194 , n50193 );
buf ( n50195 , n50194 );
or ( n50196 , n24400 , n19634 );
and ( n50197 , n24429 , n20353 );
or ( n50198 , n20562 , n24443 );
or ( n50199 , n20559 , n24438 );
not ( n50200 , n39924 );
nand ( n50201 , n50198 , n50199 , n50200 );
nor ( n50202 , n50197 , n50201 );
nand ( n50203 , n24415 , n20515 );
nand ( n50204 , n19650 , n32242 );
and ( n50205 , n50202 , n50203 , n50204 );
nand ( n50206 , n50196 , n50205 );
buf ( n50207 , n50206 );
buf ( n50208 , n50207 );
nand ( n50209 , n30713 , n28408 );
nand ( n50210 , n30732 , n32751 );
nand ( n50211 , n30741 , n29163 );
nand ( n50212 , n28451 , n40478 );
and ( n50213 , n32755 , n12255 );
or ( n50214 , n32757 , n12240 );
nand ( n50215 , n50214 , n40073 );
nor ( n50216 , n50213 , n50215 );
and ( n50217 , n50211 , n50212 , n50216 );
nand ( n50218 , n50209 , n50210 , n50217 );
buf ( n50219 , n50218 );
buf ( n50220 , n50219 );
or ( n50221 , n48928 , n27647 );
nand ( n50222 , n34674 , n13501 );
nand ( n50223 , n50221 , n50222 );
buf ( n50224 , n50223 );
buf ( n50225 , n50224 );
not ( n50226 , n275929 );
buf ( n50227 , n50226 );
buf ( n50228 , n50227 );
not ( n50229 , n275550 );
buf ( n50230 , n50229 );
buf ( n50231 , n50230 );
buf ( n50232 , n275554 );
buf ( n50233 , n275554 );
or ( n50234 , n36036 , n36861 );
and ( n50235 , n45676 , n275778 );
and ( n50236 , n36079 , n36083 );
not ( n50237 , n50236 );
and ( n50238 , n36135 , n36105 );
nor ( n50239 , n50238 , n36073 );
not ( n50240 , n50239 );
or ( n50241 , n50237 , n50240 );
or ( n50242 , n50239 , n50236 );
nand ( n50243 , n50241 , n50242 );
buf ( n50244 , n50243 );
not ( n50245 , n50244 );
not ( n50246 , n36155 );
or ( n50247 , n50245 , n50246 );
and ( n50248 , n36189 , n36193 );
not ( n50249 , n50248 );
and ( n50250 , n36241 , n36213 );
nor ( n50251 , n50250 , n36184 );
not ( n50252 , n50251 );
or ( n50253 , n50249 , n50252 );
or ( n50254 , n50251 , n50248 );
nand ( n50255 , n50253 , n50254 );
buf ( n50256 , n50255 );
nand ( n50257 , n41635 , n50256 );
nand ( n50258 , n50247 , n50257 );
nor ( n50259 , n50235 , n50258 );
nand ( n50260 , n50234 , n50259 );
nand ( n50261 , n50260 , n20645 );
and ( n50262 , n36341 , n36326 );
not ( n50263 , n50262 );
and ( n50264 , n49408 , n36330 );
nor ( n50265 , n50264 , n36336 );
not ( n50266 , n50265 );
or ( n50267 , n50263 , n50266 );
or ( n50268 , n50265 , n50262 );
nand ( n50269 , n50267 , n50268 );
buf ( n50270 , n50269 );
nand ( n50271 , n36267 , n50270 );
and ( n50272 , n36444 , n36429 );
not ( n50273 , n50272 );
and ( n50274 , n49418 , n36433 );
nor ( n50275 , n50274 , n36439 );
not ( n50276 , n50275 );
or ( n50277 , n50273 , n50276 );
or ( n50278 , n50275 , n50272 );
nand ( n50279 , n50277 , n50278 );
buf ( n50280 , n50279 );
nand ( n50281 , n36371 , n50280 );
and ( n50282 , n36474 , n36077 );
or ( n50283 , n20654 , n275777 );
nand ( n50284 , n50283 , n49696 );
nor ( n50285 , n50282 , n50284 );
nand ( n50286 , n50261 , n50271 , n50281 , n50285 );
buf ( n50287 , n50286 );
buf ( n50288 , n50287 );
buf ( n50289 , n275554 );
not ( n50290 , n275550 );
buf ( n50291 , n50290 );
buf ( n50292 , n50291 );
buf ( n50293 , n275554 );
or ( n50294 , n38146 , n20950 );
nand ( n50295 , n20950 , n13657 );
nand ( n50296 , n50294 , n50295 );
buf ( n50297 , n50296 );
buf ( n50298 , n50297 );
and ( n50299 , n9158 , n41925 );
not ( n50300 , n9158 );
and ( n50301 , n50300 , n10644 );
or ( n50302 , n50299 , n50301 );
buf ( n50303 , n50302 );
buf ( n50304 , n50303 );
not ( n50305 , n275929 );
buf ( n50306 , n50305 );
buf ( n50307 , n50306 );
buf ( n50308 , n275554 );
or ( n50309 , n38053 , n29866 );
nand ( n50310 , n38076 , n20353 );
nand ( n50311 , n38101 , n30132 );
not ( n50312 , n34104 );
not ( n50313 , n38107 );
and ( n50314 , n50312 , n50313 );
nand ( n50315 , n38120 , n31095 );
nand ( n50316 , n29494 , n38125 );
nand ( n50317 , n30179 , n18508 );
nand ( n50318 , n50315 , n50316 , n50317 );
nor ( n50319 , n50314 , n50318 );
and ( n50320 , n50310 , n50311 , n50319 );
nand ( n50321 , n50309 , n50320 );
buf ( n50322 , n50321 );
buf ( n50323 , n50322 );
buf ( n50324 , n275554 );
buf ( n50325 , n275554 );
buf ( n50326 , n275554 );
or ( n50327 , n26502 , n27647 );
nand ( n50328 , n34674 , n13689 );
nand ( n50329 , n50327 , n50328 );
buf ( n50330 , n50329 );
buf ( n50331 , n50330 );
not ( n50332 , n275929 );
buf ( n50333 , n50332 );
buf ( n50334 , n50333 );
or ( n50335 , n40945 , n19216 );
and ( n50336 , n41018 , n19360 );
nand ( n50337 , n30149 , n19318 , n18440 );
nand ( n50338 , n41029 , n29075 );
nand ( n50339 , n33162 , n41034 );
nand ( n50340 , n19387 , n18457 );
nand ( n50341 , n50337 , n50338 , n50339 , n50340 );
nor ( n50342 , n50336 , n50341 );
nand ( n50343 , n40982 , n35150 );
nand ( n50344 , n50335 , n50342 , n50343 );
buf ( n50345 , n50344 );
buf ( n50346 , n50345 );
buf ( n50347 , n275554 );
and ( n50348 , n23706 , n277710 );
not ( n50349 , n23706 );
and ( n50350 , n50349 , n42837 );
or ( n50351 , n50348 , n50350 );
buf ( n50352 , n50351 );
buf ( n50353 , n50352 );
not ( n50354 , n275929 );
buf ( n50355 , n50354 );
buf ( n50356 , n50355 );
buf ( n50357 , n275554 );
buf ( n50358 , n275554 );
not ( n50359 , n17991 );
not ( n50360 , n22335 );
or ( n50361 , n50359 , n50360 );
not ( n50362 , n27930 );
or ( n50363 , n50362 , n22335 );
nand ( n50364 , n50361 , n50363 );
buf ( n50365 , n50364 );
buf ( n50366 , n50365 );
not ( n50367 , n275550 );
buf ( n50368 , n50367 );
buf ( n50369 , n50368 );
not ( n50370 , n275929 );
buf ( n50371 , n50370 );
buf ( n50372 , n50371 );
buf ( n50373 , n275554 );
or ( n50374 , n41396 , n19387 );
or ( n50375 , n19388 , n18845 );
nand ( n50376 , n50374 , n50375 );
buf ( n50377 , n50376 );
buf ( n50378 , n50377 );
not ( n50379 , n275925 );
buf ( n50380 , n50379 );
buf ( n50381 , n50380 );
not ( n50382 , n24790 );
or ( n50383 , n50382 , n29046 );
nand ( n50384 , n28252 , n9775 );
nand ( n50385 , n50383 , n50384 );
buf ( n50386 , n50385 );
buf ( n50387 , n50386 );
not ( n50388 , n275550 );
buf ( n50389 , n50388 );
buf ( n50390 , n50389 );
buf ( n50391 , n275554 );
buf ( n50392 , n275554 );
not ( n50393 , n275925 );
buf ( n50394 , n50393 );
buf ( n50395 , n50394 );
or ( n50396 , n36036 , n44884 );
and ( n50397 , n45676 , n275816 );
nand ( n50398 , n50109 , n36092 );
not ( n50399 , n50398 );
nand ( n50400 , n41884 , n50106 );
not ( n50401 , n50400 );
or ( n50402 , n50399 , n50401 );
or ( n50403 , n50400 , n50398 );
nand ( n50404 , n50402 , n50403 );
buf ( n50405 , n50404 );
not ( n50406 , n50405 );
not ( n50407 , n36155 );
or ( n50408 , n50406 , n50407 );
nand ( n50409 , n50129 , n36202 );
not ( n50410 , n50409 );
nand ( n50411 , n41983 , n50126 );
not ( n50412 , n50411 );
or ( n50413 , n50410 , n50412 );
or ( n50414 , n50411 , n50409 );
nand ( n50415 , n50413 , n50414 );
buf ( n50416 , n50415 );
nand ( n50417 , n41635 , n50416 );
nand ( n50418 , n50408 , n50417 );
nor ( n50419 , n50397 , n50418 );
nand ( n50420 , n50396 , n50419 );
nand ( n50421 , n50420 , n20645 );
nor ( n50422 , n50145 , n36345 );
not ( n50423 , n50422 );
nor ( n50424 , n36332 , n36342 );
not ( n50425 , n50424 );
or ( n50426 , n50423 , n50425 );
or ( n50427 , n50424 , n50422 );
nand ( n50428 , n50426 , n50427 );
buf ( n50429 , n50428 );
nand ( n50430 , n36267 , n50429 );
nor ( n50431 , n50157 , n36448 );
not ( n50432 , n50431 );
nor ( n50433 , n36435 , n36445 );
not ( n50434 , n50433 );
or ( n50435 , n50432 , n50434 );
or ( n50436 , n50433 , n50431 );
nand ( n50437 , n50435 , n50436 );
buf ( n50438 , n50437 );
nand ( n50439 , n36371 , n50438 );
and ( n50440 , n36474 , n10718 );
or ( n50441 , n20654 , n275815 );
nand ( n50442 , n50441 , n42567 );
nor ( n50443 , n50440 , n50442 );
nand ( n50444 , n50421 , n50430 , n50439 , n50443 );
buf ( n50445 , n50444 );
buf ( n50446 , n50445 );
not ( n50447 , n275925 );
buf ( n50448 , n50447 );
buf ( n50449 , n50448 );
buf ( n50450 , n275554 );
not ( n50451 , n34869 );
and ( n50452 , n50451 , n26440 );
nand ( n50453 , n34887 , n20889 );
nand ( n50454 , n34906 , n20927 );
and ( n50455 , n34922 , n17409 );
and ( n50456 , n20940 , n34928 );
nor ( n50457 , n50455 , n50456 );
nand ( n50458 , n50453 , n50454 , n50457 );
nor ( n50459 , n50452 , n50458 );
or ( n50460 , n50459 , n21696 );
nand ( n50461 , n34674 , n13517 );
nand ( n50462 , n50460 , n50461 );
buf ( n50463 , n50462 );
buf ( n50464 , n50463 );
buf ( n50465 , n275554 );
not ( n50466 , n275929 );
buf ( n50467 , n50466 );
buf ( n50468 , n50467 );
buf ( n50469 , n275554 );
not ( n50470 , n26782 );
or ( n50471 , n50470 , n22335 );
or ( n50472 , n275557 , n19183 );
nand ( n50473 , n50471 , n50472 );
buf ( n50474 , n50473 );
buf ( n50475 , n50474 );
not ( n50476 , n275550 );
buf ( n50477 , n50476 );
buf ( n50478 , n50477 );
not ( n50479 , n275550 );
buf ( n50480 , n50479 );
buf ( n50481 , n50480 );
buf ( n50482 , n275554 );
not ( n50483 , n275925 );
buf ( n50484 , n50483 );
buf ( n50485 , n50484 );
not ( n50486 , n275929 );
buf ( n50487 , n50486 );
buf ( n50488 , n50487 );
not ( n50489 , n19092 );
or ( n50490 , n21769 , n50489 );
not ( n50491 , n9448 );
or ( n50492 , n39544 , n50491 );
nand ( n50493 , n50490 , n50492 );
buf ( n50494 , n50493 );
buf ( n50495 , n50494 );
not ( n50496 , n275550 );
buf ( n50497 , n50496 );
buf ( n50498 , n50497 );
or ( n50499 , n50459 , n20951 );
nand ( n50500 , n20953 , n13531 );
nand ( n50501 , n50499 , n50500 );
buf ( n50502 , n50501 );
buf ( n50503 , n50502 );
buf ( n50504 , n275554 );
or ( n50505 , n35886 , n20951 );
nand ( n50506 , n20950 , n13902 );
nand ( n50507 , n50505 , n50506 );
buf ( n50508 , n50507 );
buf ( n50509 , n50508 );
not ( n50510 , n275550 );
buf ( n50511 , n50510 );
buf ( n50512 , n50511 );
buf ( n50513 , n275554 );
buf ( n50514 , n275554 );
not ( n50515 , n20103 );
not ( n50516 , n275557 );
or ( n50517 , n50515 , n50516 );
nand ( n50518 , n22335 , n18071 );
nand ( n50519 , n50517 , n50518 );
buf ( n50520 , n50519 );
buf ( n50521 , n50520 );
or ( n50522 , n20844 , n26364 );
nand ( n50523 , n20885 , n26370 );
nand ( n50524 , n20924 , n26374 );
nand ( n50525 , n32176 , n24366 );
nand ( n50526 , n20937 , n26393 );
nand ( n50527 , n26395 , n20943 );
not ( n50528 , n37741 );
and ( n50529 , n50526 , n50527 , n50528 );
and ( n50530 , n50523 , n50524 , n50525 , n50529 );
nand ( n50531 , n50522 , n50530 );
buf ( n50532 , n50531 );
buf ( n50533 , n50532 );
buf ( n50534 , n275554 );
or ( n50535 , n37871 , n26364 );
nand ( n50536 , n37891 , n26370 );
nand ( n50537 , n37933 , n26374 );
nand ( n50538 , n35658 , n37898 );
and ( n50539 , n26395 , n37915 );
not ( n50540 , n32188 );
not ( n50541 , n37909 );
or ( n50542 , n50540 , n50541 );
not ( n50543 , n40240 );
nand ( n50544 , n50542 , n50543 );
nor ( n50545 , n50539 , n50544 );
and ( n50546 , n50536 , n50537 , n50538 , n50545 );
nand ( n50547 , n50535 , n50546 );
buf ( n50548 , n50547 );
buf ( n50549 , n50548 );
buf ( n50550 , n275554 );
and ( C0 , n275561 , n275560 );
endmodule

