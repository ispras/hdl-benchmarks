// IWLS benchmark module "decod" printed on Wed May 29 16:32:29 2002
module decod(a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u);
input
  a,
  b,
  c,
  d,
  e;
output
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r,
  s,
  t,
  u;
wire
  o0,
  \[7] ,
  \[8] ,
  \[9] ,
  \[10] ,
  \[0] ,
  \[11] ,
  \[1] ,
  \[12] ,
  \[2] ,
  \[13] ,
  \[3] ,
  \[14] ,
  \[4] ,
  \[15] ,
  \[5] ,
  n0,
  \[6] ;
assign
  o0 = e & a,
  \[7]  = o0 & (~b & (~c & ~d)),
  \[8]  = n0 & (b & (c & d)),
  \[9]  = n0 & (b & (c & ~d)),
  \[10]  = n0 & (b & (~c & d)),
  \[0]  = o0 & (b & (c & d)),
  \[11]  = n0 & (b & (~c & ~d)),
  \[1]  = o0 & (b & (c & ~d)),
  \[12]  = n0 & (~b & (c & d)),
  f = \[0] ,
  g = \[1] ,
  h = \[2] ,
  i = \[3] ,
  j = \[4] ,
  k = \[5] ,
  l = \[6] ,
  m = \[7] ,
  n = \[8] ,
  o = \[9] ,
  p = \[10] ,
  q = \[11] ,
  r = \[12] ,
  s = \[13] ,
  t = \[14] ,
  \[2]  = o0 & (b & (~c & d)),
  \[13]  = n0 & (~b & (c & ~d)),
  u = \[15] ,
  \[3]  = o0 & (b & (~c & ~d)),
  \[14]  = n0 & (~b & (~c & d)),
  \[4]  = o0 & (~b & (c & d)),
  \[15]  = n0 & (~b & (~c & ~d)),
  \[5]  = o0 & (~b & (c & ~d)),
  n0 = e & ~a,
  \[6]  = o0 & (~b & (~c & d));
endmodule

