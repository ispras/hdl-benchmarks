module logical_xor_1_1(a, b, c);
  input a;
  input b;
  output c;
  assign c = a ^^ b;
endmodule
