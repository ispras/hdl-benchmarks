// IWLS benchmark module "comp" printed on Wed May 29 16:31:29 2002
module comp(a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, \x , y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0);
input
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r,
  s,
  t,
  u,
  v,
  w,
  \x ,
  y,
  z,
  a0,
  b0,
  c0,
  d0,
  e0,
  f0;
output
  g0,
  h0,
  i0;
wire
  m0,
  \[15] ,
  \[16] ,
  o0,
  o1,
  o2,
  \[17] ,
  \[18] ,
  q0,
  s0,
  \[0] ,
  \[1] ,
  b2,
  b3,
  \[2] ,
  c1,
  d1,
  w0,
  e1,
  x0,
  f1,
  \[10] ,
  \[9] ,
  \[11] ,
  \[12] ;
assign
  m0 = (f0 & ~p) | \[15] ,
  \[15]  = (e0 & ~o) | \[9] ,
  \[16]  = (a0 & ~k) | \[10] ,
  o0 = (~d1 & (b0 & ~l)) | (\[16]  & ~d1),
  o1 = c0 & ~m,
  o2 = u & ~e,
  \[17]  = (w & ~g) | \[11] ,
  \[18]  = (s & ~c) | \[12] ,
  q0 = (\x  & ~h) | \[17] ,
  s0 = (t & ~d) | \[18] ,
  \[0]  = ~\[1]  & ~\[2] ,
  \[1]  = ~o0 & (~d1 & (~m0 & (~c1 & (~x0 & ~w0)))),
  b2 = y & ~i,
  b3 = q & ~a,
  \[2]  = (~o0 & (c1 & (~x0 & ~w0))) | ((d1 & (~x0 & ~w0)) | ((e1 & ~x0) | f1)),
  c1 = (~\[15]  & (~f0 & p)) | ((~\[9]  & (~e0 & o)) | ((~o1 & (~d0 & n)) | (~c0 & m))),
  d1 = (~\[16]  & (~b0 & l)) | ((~\[10]  & (~a0 & k)) | ((~b2 & (~z & j)) | (~y & i))),
  w0 = q0 | e1,
  e1 = (~\[17]  & (~\x  & h)) | ((~\[11]  & (~w & g)) | ((~o2 & (~v & f)) | (~u & e))),
  x0 = s0 | f1,
  f1 = (~\[18]  & (~t & d)) | ((~\[12]  & (~s & c)) | ((~b3 & (~r & b)) | (~q & a))),
  g0 = \[0] ,
  h0 = \[1] ,
  \[10]  = (z & ~j) | b2,
  i0 = \[2] ,
  \[9]  = (d0 & ~n) | o1,
  \[11]  = (v & ~f) | o2,
  \[12]  = (r & ~b) | b3;
endmodule

