module s9234_1_bench(
  blif_clk_net,
  blif_reset_net,
  g89,
  g94,
  g98,
  g102,
  g107,
  g301,
  g306,
  g310,
  g314,
  g319,
  g557,
  g558,
  g559,
  g560,
  g561,
  g562,
  g563,
  g564,
  g705,
  g639,
  g567,
  g45,
  g42,
  g39,
  g702,
  g32,
  g38,
  g46,
  g36,
  g47,
  g40,
  g37,
  g41,
  g22,
  g44,
  g23,
  g2584,
  g3222,
  g3600,
  g4307,
  g4321,
  g4422,
  g4809,
  g5137,
  g5468,
  g5469,
  g5692,
  g6282,
  g6284,
  g6360,
  g6362,
  g6364,
  g6366,
  g6368,
  g6370,
  g6372,
  g6374,
  g6728,
  g1290,
  g4121,
  g4108,
  g4106,
  g4103,
  g1293,
  g4099,
  g4102,
  g4109,
  g4100,
  g4112,
  g4105,
  g4101,
  g4110,
  g4104,
  g4107,
  g4098);
input blif_clk_net;
input blif_reset_net;
input g89;
input g94;
input g98;
input g102;
input g107;
input g301;
input g306;
input g310;
input g314;
input g319;
input g557;
input g558;
input g559;
input g560;
input g561;
input g562;
input g563;
input g564;
input g705;
input g639;
input g567;
input g45;
input g42;
input g39;
input g702;
input g32;
input g38;
input g46;
input g36;
input g47;
input g40;
input g37;
input g41;
input g22;
input g44;
input g23;
output g2584;
output g3222;
output g3600;
output g4307;
output g4321;
output g4422;
output g4809;
output g5137;
output g5468;
output g5469;
output g5692;
output g6282;
output g6284;
output g6360;
output g6362;
output g6364;
output g6366;
output g6368;
output g6370;
output g6372;
output g6374;
output g6728;
output g1290;
output g4121;
output g4108;
output g4106;
output g4103;
output g1293;
output g4099;
output g4102;
output g4109;
output g4100;
output g4112;
output g4105;
output g4101;
output g4110;
output g4104;
output g4107;
output g4098;
reg g678;
reg g332;
reg g123;
reg g207;
reg g695;
reg g461;
reg g18;
reg g292;
reg g331;
reg g689;
reg g24;
reg g465;
reg g84;
reg g291;
reg g676;
reg g622;
reg g117;
reg g278;
reg g128;
reg g598;
reg g554;
reg g496;
reg g179;
reg g48;
reg g590;
reg g551;
reg g682;
reg g11;
reg g606;
reg g188;
reg g646;
reg g327;
reg g361;
reg g289;
reg g398;
reg g684;
reg g619;
reg g208;
reg g248;
reg g390;
reg g625;
reg g681;
reg g437;
reg g276;
reg g3;
reg g323;
reg g224;
reg g685;
reg g43;
reg g157;
reg g282;
reg g697;
reg g206;
reg g449;
reg g118;
reg g528;
reg g284;
reg g426;
reg g634;
reg g669;
reg g520;
reg g281;
reg g175;
reg g15;
reg g631;
reg g69;
reg g693;
reg g337;
reg g457;
reg g486;
reg g471;
reg g328;
reg g285;
reg g418;
reg g402;
reg g297;
reg g212;
reg g410;
reg g430;
reg g33;
reg g662;
reg g453;
reg g269;
reg g574;
reg g441;
reg g664;
reg g349;
reg g211;
reg g586;
reg g571;
reg g29;
reg g326;
reg g698;
reg g654;
reg g293;
reg g690;
reg g445;
reg g374;
reg g6;
reg g687;
reg g357;
reg g386;
reg g504;
reg g665;
reg g166;
reg g541;
reg g74;
reg g338;
reg g696;
reg g516;
reg g536;
reg g683;
reg g353;
reg g545;
reg g254;
reg g341;
reg g290;
reg g2;
reg g287;
reg g336;
reg g345;
reg g628;
reg g679;
reg g28;
reg g688;
reg g283;
reg g613;
reg g10;
reg g14;
reg g680;
reg g143;
reg g672;
reg g667;
reg g366;
reg g279;
reg g492;
reg g170;
reg g686;
reg g288;
reg g638;
reg g602;
reg g642;
reg g280;
reg g663;
reg g610;
reg g148;
reg g209;
reg g675;
reg g478;
reg g122;
reg g54;
reg g594;
reg g286;
reg g489;
reg g616;
reg g79;
reg g218;
reg g242;
reg g578;
reg g184;
reg g119;
reg g668;
reg g139;
reg g422;
reg g210;
reg g394;
reg g230;
reg g25;
reg g204;
reg g658;
reg g650;
reg g378;
reg g508;
reg g548;
reg g370;
reg g406;
reg g236;
reg g500;
reg g205;
reg g197;
reg g666;
reg g114;
reg g524;
reg g260;
reg g111;
reg g131;
reg g7;
reg g19;
reg g677;
reg g582;
reg g485;
reg g699;
reg g193;
reg g135;
reg g382;
reg g414;
reg g434;
reg g266;
reg g49;
reg g152;
reg g692;
reg g277;
reg g127;
reg g161;
reg g512;
reg g532;
reg g64;
reg g694;
reg g691;
reg g1;
reg g59;
wire g2171;
wire I2596;
wire g3491;
wire g3610;
wire I8764;
wire g4355;
wire g6579;
wire I3711;
wire g4610;
wire g3892;
wire g3277;
wire g4396;
wire g4866;
wire g6365;
wire g3783;
wire g3603;
wire g4111;
wire I5793;
wire g2887;
wire I5743;
wire g6136;
wire g1276;
wire g3885;
wire I8494;
wire g1946;
wire g6034;
wire g3034;
wire g4847;
wire I9085;
wire g2776;
wire I4667;
wire g6542;
wire g6426;
wire I7463;
wire g5729;
wire g6561;
wire I4452;
wire I7963;
wire g2039;
wire g5788;
wire g6293;
wire g6577;
wire g5711;
wire I4678;
wire I5517;
wire I8872;
wire I6923;
wire g5925;
wire g5805;
wire g5216;
wire g1110;
wire I7333;
wire I8491;
wire g5025;
wire I2753;
wire g5119;
wire g2098;
wire g5099;
wire I5526;
wire I2479;
wire I4961;
wire g4342;
wire g4623;
wire g3150;
wire g5445;
wire g5778;
wire I2442;
wire g3864;
wire g4432;
wire g736;
wire g3761;
wire I2299;
wire g4157;
wire g5680;
wire g4835;
wire g4136;
wire g1628;
wire g6544;
wire I4173;
wire g4276;
wire I3556;
wire I2150;
wire g2535;
wire g6419;
wire I4526;
wire I3298;
wire g3554;
wire I8335;
wire I5195;
wire g6358;
wire g2416;
wire I2738;
wire I8821;
wire I2845;
wire g6261;
wire g1387;
wire g3366;
wire I8564;
wire g3638;
wire g4236;
wire g2859;
wire g3534;
wire I9031;
wire I8393;
wire g5498;
wire I7039;
wire g1589;
wire g5874;
wire I8209;
wire g4401;
wire I7571;
wire g6890;
wire g940;
wire I6371;
wire g2135;
wire g3670;
wire g3922;
wire g6114;
wire g4454;
wire g1822;
wire g6847;
wire g6818;
wire g5491;
wire g1063;
wire g4830;
wire g6015;
wire I5433;
wire I7692;
wire g1206;
wire I3894;
wire g5726;
wire g6853;
wire I7906;
wire g2177;
wire g4150;
wire g3029;
wire I6660;
wire g1925;
wire g6827;
wire I5603;
wire g835;
wire g4811;
wire g5673;
wire I9116;
wire I5023;
wire g5329;
wire I8196;
wire g5295;
wire g6743;
wire I2449;
wire g6101;
wire I7481;
wire g3067;
wire g3748;
wire g1841;
wire I9128;
wire g4854;
wire I7987;
wire g1829;
wire g6279;
wire g6605;
wire I9179;
wire I3019;
wire g5318;
wire g6879;
wire I6318;
wire g6837;
wire g6594;
wire g6494;
wire g3598;
wire I8713;
wire g6155;
wire I6895;
wire g1369;
wire I5233;
wire I8202;
wire g5602;
wire I2521;
wire I3137;
wire I7509;
wire g2087;
wire g893;
wire g6923;
wire I8370;
wire I2716;
wire g6333;
wire g2709;
wire g2315;
wire g6108;
wire I2420;
wire g809;
wire g5694;
wire g6142;
wire g5135;
wire I8110;
wire g3755;
wire I8285;
wire g2018;
wire g5363;
wire I2073;
wire g3848;
wire g3128;
wire g1567;
wire I6386;
wire g6587;
wire g1784;
wire g3931;
wire g3200;
wire g5185;
wire g4459;
wire g6549;
wire g4717;
wire I6093;
wire g6523;
wire g3342;
wire I2179;
wire I3534;
wire g4068;
wire g4127;
wire g4526;
wire g1813;
wire g4144;
wire g1366;
wire g5947;
wire g5946;
wire g1982;
wire I7433;
wire g3619;
wire g1344;
wire g5935;
wire g2780;
wire g6086;
wire g4619;
wire I3434;
wire I9011;
wire I6456;
wire I3056;
wire g2941;
wire I3855;
wire g4644;
wire I8653;
wire g3990;
wire I8626;
wire g2727;
wire g2340;
wire I2343;
wire I2499;
wire g3851;
wire g2307;
wire g3333;
wire g4756;
wire g6556;
wire g3936;
wire g3154;
wire I4684;
wire g4114;
wire g3646;
wire I5944;
wire g1192;
wire g3013;
wire g1665;
wire g3701;
wire I2728;
wire g4634;
wire I8378;
wire g5478;
wire g4839;
wire I6311;
wire g6822;
wire g2767;
wire g6401;
wire I8056;
wire I3358;
wire I3620;
wire g1922;
wire I7593;
wire I5783;
wire I4008;
wire I4246;
wire g5958;
wire g4699;
wire g5512;
wire I5708;
wire g4461;
wire I2284;
wire g4168;
wire g6488;
wire g4720;
wire g6150;
wire I2608;
wire I7143;
wire g5489;
wire g6269;
wire g3869;
wire I3068;
wire g3109;
wire I8800;
wire I3028;
wire g2688;
wire g4178;
wire I8837;
wire I8369;
wire g1853;
wire g3768;
wire I5702;
wire I4646;
wire g965;
wire I3244;
wire I4204;
wire g3382;
wire I5505;
wire g5141;
wire g2157;
wire g1695;
wire g2954;
wire g5541;
wire I8089;
wire g5198;
wire g3912;
wire g6691;
wire g3973;
wire I6543;
wire I7440;
wire I1980;
wire g2356;
wire g5269;
wire g4600;
wire g6065;
wire I4340;
wire g5629;
wire g6536;
wire g6055;
wire g4266;
wire g3778;
wire g4702;
wire g1861;
wire g2078;
wire I8946;
wire I3485;
wire I6177;
wire g2915;
wire g4120;
wire g5373;
wire g1847;
wire I5427;
wire g3958;
wire g3807;
wire g6900;
wire g5074;
wire g6147;
wire g2112;
wire g6093;
wire g4603;
wire g6185;
wire I8066;
wire g2733;
wire I6612;
wire g2876;
wire I2023;
wire g5565;
wire I5720;
wire g932;
wire g1675;
wire I2278;
wire I5460;
wire I4166;
wire g6371;
wire I2508;
wire I2324;
wire g4777;
wire g5047;
wire I8500;
wire I2825;
wire I6819;
wire I3340;
wire g6654;
wire g4249;
wire I8997;
wire g3991;
wire g3465;
wire g2030;
wire g4637;
wire g5916;
wire g2025;
wire g2265;
wire g1887;
wire g4285;
wire I2961;
wire I7002;
wire g5274;
wire I5648;
wire g2796;
wire g5536;
wire I6963;
wire I5400;
wire g5159;
wire g5210;
wire I5644;
wire I3699;
wire g3053;
wire g1960;
wire g4468;
wire I7197;
wire I2880;
wire g1637;
wire g3571;
wire g4803;
wire g5142;
wire g6416;
wire g3094;
wire g3463;
wire g6239;
wire g4333;
wire g4508;
wire I5768;
wire I3071;
wire g4812;
wire I3740;
wire g1219;
wire g3377;
wire I5442;
wire I6143;
wire I3328;
wire I4252;
wire g1043;
wire g6176;
wire g6909;
wire I7313;
wire I2290;
wire I6475;
wire I3954;
wire g3772;
wire g4267;
wire I5865;
wire g2419;
wire g3144;
wire I2134;
wire g3651;
wire I2013;
wire g1899;
wire g6884;
wire g2712;
wire I8476;
wire I2143;
wire g1641;
wire g3779;
wire g3329;
wire g1703;
wire I2221;
wire I4623;
wire g4628;
wire g4566;
wire I8730;
wire g4698;
wire g3834;
wire g1319;
wire I7170;
wire g1123;
wire I8273;
wire g4732;
wire I7871;
wire I2399;
wire I2199;
wire g6327;
wire g5894;
wire I5837;
wire g5601;
wire g2719;
wire I8809;
wire I6391;
wire g3697;
wire g6434;
wire g4002;
wire I5214;
wire g5527;
wire g4661;
wire I2109;
wire I5071;
wire I5209;
wire I9098;
wire I8512;
wire g6252;
wire g4435;
wire g5948;
wire g4824;
wire g2864;
wire g2781;
wire g2961;
wire I8659;
wire g6569;
wire g4387;
wire g5624;
wire I7097;
wire I2334;
wire g2771;
wire I5019;
wire I5301;
wire g5054;
wire g3028;
wire g6301;
wire g5996;
wire g5191;
wire g1518;
wire g5160;
wire I1947;
wire g4900;
wire g4219;
wire I8897;
wire g4790;
wire g2766;
wire g3517;
wire g1327;
wire g1334;
wire I2340;
wire g709;
wire I3112;
wire g5454;
wire I8432;
wire g5177;
wire g4170;
wire g2253;
wire g3375;
wire g2975;
wire g3082;
wire I6403;
wire I6063;
wire g3874;
wire I7521;
wire g2515;
wire I4809;
wire I8620;
wire g5676;
wire g6899;
wire I2349;
wire g4382;
wire I8650;
wire g2850;
wire I2601;
wire g5010;
wire I2663;
wire g1236;
wire g6767;
wire g6670;
wire I5068;
wire g6465;
wire g4225;
wire g4565;
wire g4188;
wire g4853;
wire g5251;
wire I6420;
wire g3661;
wire I3999;
wire g2588;
wire I3990;
wire I6661;
wire I2611;
wire g1583;
wire g6420;
wire g4678;
wire g4222;
wire g5630;
wire g3631;
wire g3726;
wire g2494;
wire I7478;
wire g3457;
wire g4404;
wire I7254;
wire g5687;
wire I6346;
wire g5582;
wire I7230;
wire g3829;
wire g1046;
wire g850;
wire I3031;
wire g4607;
wire g6260;
wire I3468;
wire g3871;
wire I8834;
wire g5554;
wire I4009;
wire I7570;
wire g6679;
wire g6456;
wire I8576;
wire g1575;
wire g3593;
wire g2440;
wire g3966;
wire I8255;
wire g3177;
wire I8074;
wire I3540;
wire I6659;
wire g2959;
wire g4873;
wire g6444;
wire I6579;
wire I8961;
wire g6376;
wire I4445;
wire g4596;
wire g897;
wire I8441;
wire g4613;
wire g6771;
wire I6362;
wire g3302;
wire g5797;
wire I3641;
wire I3779;
wire g2091;
wire I7058;
wire g6429;
wire g5085;
wire g5515;
wire I8727;
wire g1160;
wire I7802;
wire I2653;
wire g6553;
wire g3986;
wire g2343;
wire I3691;
wire g4048;
wire g5617;
wire g1880;
wire I3516;
wire g5435;
wire g3299;
wire I8180;
wire g6601;
wire g4840;
wire g4446;
wire g5486;
wire g1116;
wire I5532;
wire I2943;
wire g2647;
wire I8524;
wire I8423;
wire I7972;
wire g3684;
wire I5382;
wire I8479;
wire g1684;
wire g945;
wire g6937;
wire g1233;
wire g5358;
wire g1439;
wire g5138;
wire I7223;
wire g3118;
wire I2998;
wire g5242;
wire g4585;
wire g862;
wire g4180;
wire g1484;
wire I5760;
wire I6417;
wire g3290;
wire I4123;
wire g4502;
wire g6308;
wire I9170;
wire g6044;
wire g2541;
wire I8913;
wire g3658;
wire g1998;
wire g3228;
wire g3903;
wire g5864;
wire g3859;
wire g6616;
wire I7167;
wire g2906;
wire g1076;
wire g3671;
wire g2754;
wire I5686;
wire I1825;
wire g3782;
wire I2630;
wire I8860;
wire I8079;
wire g3076;
wire I2428;
wire I1874;
wire I3816;
wire I3109;
wire g5395;
wire g5553;
wire g3535;
wire I3927;
wire I8975;
wire I8165;
wire g5937;
wire g2720;
wire g5450;
wire g2243;
wire I7372;
wire g3367;
wire g5492;
wire g2608;
wire g6812;
wire I6549;
wire I4334;
wire g5310;
wire I7686;
wire g6102;
wire g2179;
wire I4159;
wire g6402;
wire g6828;
wire g4723;
wire I4273;
wire I9119;
wire g4054;
wire I2627;
wire I2721;
wire g1821;
wire I3575;
wire g2158;
wire g6848;
wire I6473;
wire g929;
wire g1581;
wire I9092;
wire g2104;
wire I8195;
wire g6817;
wire g3195;
wire g3840;
wire g3480;
wire g4044;
wire I7173;
wire g6094;
wire g4451;
wire g5499;
wire I6733;
wire g3821;
wire g3923;
wire g6535;
wire I8656;
wire g4213;
wire g6924;
wire g3289;
wire I6956;
wire g1842;
wire I5630;
wire g6070;
wire g3276;
wire g4730;
wire g3459;
wire g3902;
wire g3291;
wire g1108;
wire g2631;
wire I7153;
wire g3972;
wire I5328;
wire g1820;
wire g894;
wire g2800;
wire g4137;
wire g4494;
wire g3743;
wire I3313;
wire g6541;
wire g3611;
wire g6135;
wire g6543;
wire I7267;
wire g1711;
wire g5303;
wire I5309;
wire I8203;
wire g1891;
wire g4611;
wire g3490;
wire g5693;
wire I5385;
wire g4155;
wire g2568;
wire g3886;
wire g849;
wire I6933;
wire g2891;
wire g4156;
wire I8309;
wire I6340;
wire g4356;
wire I3528;
wire I3833;
wire g3379;
wire g6427;
wire I6072;
wire I3569;
wire g1498;
wire I7548;
wire g6248;
wire g2607;
wire I5622;
wire g4343;
wire g6500;
wire g5250;
wire g6697;
wire I2542;
wire I2408;
wire g5875;
wire g3833;
wire g5777;
wire g2663;
wire g4657;
wire I6995;
wire g749;
wire g6896;
wire I5177;
wire I8573;
wire I3629;
wire g5682;
wire g6271;
wire I3965;
wire g4395;
wire I6615;
wire I2620;
wire I5109;
wire g3685;
wire g2213;
wire g4134;
wire g6614;
wire I3614;
wire g5087;
wire g3343;
wire I3419;
wire I8150;
wire I4347;
wire g1052;
wire g5446;
wire g5351;
wire g6309;
wire I9185;
wire g5049;
wire I5705;
wire g2858;
wire g1059;
wire g1720;
wire g760;
wire I5264;
wire g3984;
wire I5654;
wire g4057;
wire g1833;
wire g4115;
wire g1696;
wire g3332;
wire g5477;
wire g3095;
wire I2391;
wire I7576;
wire g5062;
wire g3437;
wire g4460;
wire g6268;
wire I8147;
wire g5936;
wire I2683;
wire g1594;
wire I4205;
wire I4223;
wire g5149;
wire g2059;
wire g4160;
wire I6170;
wire g5540;
wire g5888;
wire I2067;
wire g3911;
wire g4932;
wire g3760;
wire I2014;
wire g6770;
wire I4288;
wire I6706;
wire g1772;
wire I4195;
wire g5277;
wire I6444;
wire g1762;
wire g3767;
wire I3471;
wire I3013;
wire I7562;
wire g6748;
wire g6125;
wire g2701;
wire I7587;
wire I7336;
wire g2839;
wire g4179;
wire g5197;
wire g5217;
wire g3180;
wire I3395;
wire g2357;
wire g2136;
wire g6373;
wire g2111;
wire g5326;
wire g2015;
wire g6690;
wire g4218;
wire g4374;
wire I4031;
wire g4601;
wire g3792;
wire g3383;
wire I5784;
wire g4703;
wire I7796;
wire I3047;
wire g6512;
wire g5451;
wire I8888;
wire g6738;
wire g5379;
wire g4778;
wire I7081;
wire I3596;
wire g6066;
wire g5372;
wire g4669;
wire g1220;
wire I2676;
wire g4247;
wire g6334;
wire g4865;
wire g3901;
wire I2358;
wire g3963;
wire g6588;
wire g2079;
wire g1848;
wire g2585;
wire g3327;
wire I7698;
wire g3883;
wire g2053;
wire g4221;
wire g3683;
wire g1620;
wire g1609;
wire g6524;
wire g1555;
wire g6744;
wire g2550;
wire g6941;
wire g6077;
wire I2898;
wire g4716;
wire g6363;
wire g4248;
wire g3649;
wire g3127;
wire g5387;
wire I8638;
wire g5660;
wire I3669;
wire g6685;
wire I8665;
wire g2306;
wire g710;
wire I6561;
wire I2072;
wire g4527;
wire I2877;
wire g6035;
wire I7104;
wire I2893;
wire g4145;
wire g3891;
wire g5231;
wire I2682;
wire I5081;
wire g2672;
wire g2134;
wire g4708;
wire g5186;
wire g4309;
wire I8818;
wire g2509;
wire I8857;
wire g5995;
wire g5782;
wire g6493;
wire g4126;
wire g1690;
wire I9233;
wire g1854;
wire g3203;
wire I3934;
wire g1988;
wire g4237;
wire I5484;
wire g2726;
wire I8707;
wire g2675;
wire g1111;
wire I2617;
wire g2252;
wire g4667;
wire g5943;
wire g3626;
wire g6310;
wire I8420;
wire I6114;
wire I4939;
wire g3930;
wire g6530;
wire I6534;
wire g1797;
wire g1398;
wire g5069;
wire g6507;
wire I2498;
wire g4226;
wire I9208;
wire g5330;
wire I5882;
wire g6156;
wire g6141;
wire I8379;
wire g2043;
wire I4935;
wire g6236;
wire I9038;
wire I5548;
wire g1459;
wire I8159;
wire I8411;
wire g6322;
wire I7556;
wire g4597;
wire g1642;
wire g1274;
wire g2882;
wire I8044;
wire g3704;
wire g1335;
wire I2537;
wire I2675;
wire g4047;
wire g3238;
wire I6685;
wire g5234;
wire g2370;
wire g5863;
wire g2554;
wire g6417;
wire g6698;
wire g5924;
wire g3326;
wire I5659;
wire I5252;
wire I8541;
wire g3376;
wire I6187;
wire I3083;
wire g1122;
wire I2053;
wire g4457;
wire I5952;
wire g6144;
wire I9101;
wire g5574;
wire g6669;
wire g2953;
wire g1519;
wire I8177;
wire I8544;
wire g1283;
wire I3653;
wire I3617;
wire g5202;
wire g2042;
wire g2295;
wire g3921;
wire g6799;
wire g1593;
wire g6435;
wire I8246;
wire I7583;
wire I5208;
wire I6299;
wire I2916;
wire g1117;
wire g6572;
wire g1318;
wire I3647;
wire g1655;
wire g5485;
wire g1759;
wire g6492;
wire I8582;
wire g2212;
wire g6048;
wire g5531;
wire g5048;
wire I2785;
wire g4670;
wire g4513;
wire I8290;
wire I1995;
wire I5692;
wire g6883;
wire I8916;
wire g6302;
wire g4388;
wire g6706;
wire g4660;
wire g6803;
wire I3952;
wire g5524;
wire I4516;
wire g6511;
wire I6126;
wire I5249;
wire g1654;
wire g2625;
wire I3843;
wire g5178;
wire I7646;
wire I3093;
wire g6655;
wire I7091;
wire g4206;
wire g3858;
wire g6710;
wire I3074;
wire g6754;
wire g4842;
wire I6775;
wire I5481;
wire g6117;
wire I5647;
wire I9137;
wire g1426;
wire g5166;
wire g4161;
wire g2024;
wire g5228;
wire g6660;
wire I6962;
wire g4636;
wire g2740;
wire I3502;
wire g2734;
wire g899;
wire g6747;
wire g1664;
wire g5537;
wire I3441;
wire g2066;
wire g5821;
wire g6421;
wire g6930;
wire g5143;
wire g5211;
wire g6314;
wire g3052;
wire g950;
wire I3158;
wire g5120;
wire g3192;
wire I6102;
wire I7535;
wire g1769;
wire I5403;
wire I6099;
wire g4948;
wire g4764;
wire g4559;
wire g830;
wire I8467;
wire g6085;
wire g6720;
wire I2122;
wire I8881;
wire I6084;
wire g719;
wire I2207;
wire g4805;
wire g5436;
wire I3361;
wire g6130;
wire g4503;
wire g3223;
wire g6554;
wire I7342;
wire g1161;
wire I8279;
wire g3672;
wire g5245;
wire I4444;
wire g3650;
wire g6450;
wire I6414;
wire g6841;
wire g1702;
wire g5218;
wire g3616;
wire g6915;
wire g3301;
wire g4769;
wire g4035;
wire I9021;
wire g5804;
wire g6617;
wire g1292;
wire g5787;
wire I5520;
wire I6105;
wire g2936;
wire g3054;
wire I6231;
wire g6167;
wire I5412;
wire I7549;
wire g3985;
wire g2933;
wire g3161;
wire g3176;
wire g898;
wire g6173;
wire I2883;
wire g4189;
wire g1683;
wire g948;
wire g6736;
wire g4181;
wire g834;
wire g4240;
wire g3229;
wire g6701;
wire g5883;
wire g939;
wire g4662;
wire g2907;
wire g2875;
wire g6255;
wire g861;
wire g6792;
wire g6600;
wire g4798;
wire I7971;
wire I5116;
wire g5170;
wire g4800;
wire I7073;
wire g6768;
wire g4789;
wire I6816;
wire g5053;
wire g5854;
wire g2174;
wire g1411;
wire g3499;
wire I3346;
wire g2819;
wire g3729;
wire I7224;
wire g4436;
wire g4509;
wire g3601;
wire g5623;
wire I2835;
wire g3845;
wire I3776;
wire g2656;
wire g2137;
wire g6838;
wire g5562;
wire I6525;
wire I6033;
wire g3992;
wire g3374;
wire g1001;
wire g4403;
wire I4229;
wire I4267;
wire g5209;
wire g4443;
wire g1282;
wire I3697;
wire g3315;
wire g1729;
wire g3629;
wire I7065;
wire g6162;
wire g1852;
wire g1402;
wire I6008;
wire g4429;
wire g6604;
wire I8030;
wire I4940;
wire g3453;
wire I7098;
wire I5938;
wire I5236;
wire g3873;
wire I8894;
wire I7683;
wire g1546;
wire I2989;
wire g4804;
wire g3089;
wire g2164;
wire g5281;
wire I3222;
wire I5316;
wire g1574;
wire g6622;
wire g4545;
wire I4240;
wire g6109;
wire I3493;
wire g1573;
wire g2125;
wire I2791;
wire g4472;
wire g6628;
wire g6319;
wire I3788;
wire g4564;
wire g5424;
wire I5668;
wire I2958;
wire g6739;
wire g5433;
wire g1191;
wire I3893;
wire g4328;
wire g4606;
wire I6054;
wire g5406;
wire g3854;
wire g3828;
wire g3669;
wire g5429;
wire I1938;
wire I6321;
wire g3288;
wire g5583;
wire g3143;
wire g1045;
wire I8417;
wire I3741;
wire g1584;
wire g3458;
wire g4053;
wire I4366;
wire g3773;
wire g3660;
wire g2682;
wire I2004;
wire g3884;
wire I5594;
wire g6940;
wire g6099;
wire I6452;
wire g5051;
wire I5189;
wire g5183;
wire g4712;
wire g4715;
wire I5609;
wire g4758;
wire g6140;
wire g3757;
wire g1978;
wire g6568;
wire I5782;
wire I2473;
wire I4784;
wire g2586;
wire g6529;
wire g3529;
wire g2705;
wire g3718;
wire g5992;
wire g4363;
wire g6157;
wire I5084;
wire g6335;
wire I6630;
wire I1969;
wire I6649;
wire g928;
wire I3874;
wire g2671;
wire g6454;
wire g6294;
wire g6250;
wire g4129;
wire g2551;
wire g3084;
wire g4116;
wire I6531;
wire I7543;
wire g2923;
wire g5068;
wire g1556;
wire g5752;
wire g6431;
wire g6849;
wire g3090;
wire g6300;
wire g6745;
wire g4658;
wire I2373;
wire g2577;
wire g5994;
wire g5151;
wire I2405;
wire g2524;
wire I8138;
wire I2811;
wire I9082;
wire g3933;
wire g3728;
wire g4786;
wire I7550;
wire g4238;
wire I1871;
wire I1924;
wire I6567;
wire g3357;
wire g1743;
wire I1856;
wire g2089;
wire g4173;
wire I2172;
wire g5696;
wire g6558;
wire g1774;
wire g5376;
wire g5443;
wire I2922;
wire I4964;
wire I2062;
wire I4402;
wire I2899;
wire g3075;
wire I3935;
wire g6731;
wire g6406;
wire g1831;
wire I8235;
wire g5147;
wire I6976;
wire g6298;
wire g6864;
wire g5552;
wire g3680;
wire I7707;
wire I4315;
wire g1249;
wire g3354;
wire g6534;
wire g2769;
wire g5230;
wire g2744;
wire I3099;
wire g2913;
wire I7209;
wire g4583;
wire I6582;
wire I6182;
wire g6589;
wire g4772;
wire I5790;
wire g5949;
wire g1529;
wire I8535;
wire I5436;
wire g4631;
wire I6809;
wire g1481;
wire g4722;
wire g5668;
wire g4967;
wire g3541;
wire I2074;
wire g3019;
wire g1595;
wire g3820;
wire I8755;
wire g6593;
wire I4802;
wire g2230;
wire g1721;
wire g5476;
wire g4246;
wire g6230;
wire g6259;
wire g2835;
wire g5955;
wire I4919;
wire g6340;
wire g3690;
wire g3286;
wire I7261;
wire I8681;
wire g2692;
wire g5791;
wire I3906;
wire I8552;
wire g5563;
wire I2749;
wire g4608;
wire I1978;
wire g5632;
wire g4560;
wire g3209;
wire I8093;
wire I8360;
wire g6902;
wire I6740;
wire g1845;
wire g1710;
wire g6263;
wire g4394;
wire g996;
wire I5308;
wire g5681;
wire g3785;
wire I9164;
wire g1514;
wire g4933;
wire g3275;
wire g6684;
wire I5451;
wire I2979;
wire g1826;
wire g4292;
wire g3928;
wire I7577;
wire I2910;
wire g6351;
wire g2865;
wire g3612;
wire g4135;
wire g5449;
wire I4324;
wire g3320;
wire g1359;
wire I4258;
wire g6074;
wire I2681;
wire g1267;
wire I3206;
wire I5948;
wire I2244;
wire g3862;
wire g3364;
wire g5386;
wire I2417;
wire I7838;
wire I3723;
wire g5546;
wire g6878;
wire g4045;
wire g5309;
wire g2160;
wire g3311;
wire I8907;
wire g3841;
wire g2787;
wire I3942;
wire g4162;
wire I3007;
wire g4871;
wire g821;
wire I4537;
wire g5227;
wire I5320;
wire g6505;
wire I2724;
wire g4378;
wire I8300;
wire g4493;
wire g4340;
wire I1841;
wire g6281;
wire I8778;
wire g5776;
wire I9014;
wire I4510;
wire g6229;
wire g5439;
wire g3368;
wire g5418;
wire g5915;
wire g2602;
wire I4410;
wire I5037;
wire I4955;
wire g2106;
wire g6032;
wire I3478;
wire g3031;
wire g2155;
wire I6437;
wire g2612;
wire I7232;
wire g4549;
wire g1060;
wire g5246;
wire g2687;
wire I2992;
wire I3659;
wire g3186;
wire g4524;
wire I6992;
wire g3532;
wire g4186;
wire g5117;
wire g2119;
wire g2244;
wire g4314;
wire g2805;
wire I5753;
wire g3983;
wire I5756;
wire I9110;
wire g3703;
wire I2382;
wire I4040;
wire I8863;
wire g5327;
wire g4625;
wire g1918;
wire g1560;
wire g4837;
wire I7514;
wire g2653;
wire I4151;
wire I2119;
wire g1773;
wire I7042;
wire g4832;
wire I3400;
wire g2956;
wire I7358;
wire g6796;
wire g4385;
wire I6334;
wire g3867;
wire I9173;
wire g3893;
wire I4471;
wire g2853;
wire g1706;
wire g4210;
wire I6474;
wire g5452;
wire g6276;
wire I2890;
wire g1578;
wire I6186;
wire g4372;
wire I7069;
wire g3742;
wire g4004;
wire g3538;
wire g6118;
wire g3608;
wire g6829;
wire g5675;
wire g798;
wire g1460;
wire g5530;
wire g1288;
wire I7150;
wire g6124;
wire g5774;
wire g3340;
wire g2752;
wire g2609;
wire g3777;
wire g3969;
wire g2175;
wire I9095;
wire g5140;
wire g1734;
wire g4700;
wire g3489;
wire g6741;
wire g3190;
wire I3457;
wire g6830;
wire I8488;
wire g1679;
wire I8724;
wire g4380;
wire g6483;
wire I9158;
wire g3633;
wire I5359;
wire g5045;
wire g6931;
wire g6839;
wire g3733;
wire g4428;
wire g5649;
wire g2802;
wire g2758;
wire I4321;
wire g3232;
wire g1940;
wire g5331;
wire g4220;
wire g3663;
wire g5857;
wire g4488;
wire g1838;
wire g5356;
wire g4851;
wire g5012;
wire g1321;
wire g1931;
wire I6078;
wire I3698;
wire g3876;
wire g3498;
wire I3413;
wire g1011;
wire I7536;
wire g5256;
wire I8884;
wire g2118;
wire g5165;
wire g6189;
wire g4456;
wire I6812;
wire I4261;
wire g1332;
wire g2791;
wire g5505;
wire g2497;
wire I6051;
wire g5741;
wire g938;
wire g6704;
wire g4914;
wire I4243;
wire I5091;
wire g4531;
wire g3191;
wire g5584;
wire g1577;
wire g4406;
wire g6133;
wire g6913;
wire I3050;
wire g2268;
wire I5430;
wire g1190;
wire g4598;
wire g3504;
wire g6439;
wire I4351;
wire I5424;
wire I2805;
wire g4371;
wire g4227;
wire g4819;
wire g5407;
wire g4701;
wire g3341;
wire g4536;
wire g2826;
wire g3488;
wire I5197;
wire I1988;
wire g6844;
wire g6893;
wire g5391;
wire I7099;
wire g2934;
wire g6618;
wire g5061;
wire g5923;
wire I7245;
wire g4195;
wire g3421;
wire I8521;
wire g2275;
wire I2385;
wire I3678;
wire I3268;
wire g1328;
wire I8081;
wire g6057;
wire g6729;
wire I5418;
wire g6571;
wire g5910;
wire g6504;
wire I7528;
wire g1682;
wire g2818;
wire g6447;
wire I3399;
wire g6321;
wire g2813;
wire g1928;
wire I3755;
wire I5243;
wire g5233;
wire g1291;
wire g5637;
wire g2916;
wire g1969;
wire g3751;
wire g6486;
wire I6283;
wire I3864;
wire I6783;
wire I4468;
wire g1138;
wire g4471;
wire g4349;
wire g2446;
wire I8806;
wire I6485;
wire g3644;
wire g3609;
wire g1935;
wire I7029;
wire g3522;
wire g3929;
wire g1410;
wire I6377;
wire I8591;
wire g3857;
wire g5171;
wire I5998;
wire I7237;
wire g3837;
wire g1088;
wire I9131;
wire g5880;
wire g3905;
wire g3989;
wire I3505;
wire g3434;
wire I5637;
wire g2908;
wire g3710;
wire g2293;
wire g5308;
wire g3842;
wire g4353;
wire g4046;
wire g6824;
wire g1250;
wire g2544;
wire I9028;
wire g4845;
wire I9035;
wire I5394;
wire g4511;
wire g2892;
wire I3059;
wire g5112;
wire g1395;
wire g4017;
wire g3971;
wire g2096;
wire g6491;
wire I3846;
wire I2485;
wire g5813;
wire g2743;
wire I3970;
wire g2166;
wire g4265;
wire g4430;
wire I7113;
wire g2008;
wire g5670;
wire I7640;
wire g2073;
wire I2700;
wire I3717;
wire g6313;
wire I9052;
wire I4371;
wire I4437;
wire g4763;
wire I7355;
wire I6289;
wire I6269;
wire g3451;
wire I7541;
wire I4743;
wire g2323;
wire g1905;
wire g3030;
wire g4500;
wire g3309;
wire I6096;
wire I5406;
wire I2707;
wire I7193;
wire g5603;
wire I2797;
wire g4043;
wire I6406;
wire g4399;
wire g6650;
wire I6081;
wire g930;
wire I4212;
wire g5077;
wire g6621;
wire I3800;
wire I8264;
wire I2982;
wire I5933;
wire I5537;
wire g2834;
wire g1586;
wire I8644;
wire g1659;
wire g6243;
wire g6240;
wire I6315;
wire g2995;
wire g6693;
wire g6468;
wire I9122;
wire I3148;
wire I4501;
wire I8594;
wire g2067;
wire g2196;
wire g4609;
wire g3815;
wire g1375;
wire I3456;
wire g6673;
wire I4433;
wire g848;
wire I5454;
wire I5153;
wire g2555;
wire g6842;
wire I7808;
wire I7210;
wire g4205;
wire g2845;
wire g1534;
wire I6666;
wire I8171;
wire g3001;
wire g4561;
wire I5056;
wire I5876;
wire g6514;
wire I5926;
wire I5696;
wire I2776;
wire g3236;
wire g5201;
wire g6151;
wire g3756;
wire g6361;
wire I2854;
wire g2721;
wire g2505;
wire g3502;
wire g1733;
wire I6570;
wire g1039;
wire g6644;
wire I8153;
wire g6886;
wire g4941;
wire g6084;
wire I2015;
wire g2001;
wire g4949;
wire g5059;
wire I6918;
wire g2413;
wire g5381;
wire I2674;
wire I3961;
wire g2897;
wire I5094;
wire I6964;
wire g2924;
wire g3022;
wire I8276;
wire g5434;
wire I6763;
wire I3247;
wire g6705;
wire g5193;
wire g1275;
wire I4495;
wire g3117;
wire g2084;
wire I4920;
wire g4783;
wire I3037;
wire g6436;
wire g2777;
wire g5575;
wire g6345;
wire g2460;
wire g5695;
wire g3355;
wire g4492;
wire I5633;
wire g6014;
wire g3239;
wire g5260;
wire g6659;
wire I2218;
wire g5892;
wire g2296;
wire g2866;
wire g2484;
wire g6329;
wire g5628;
wire I9074;
wire g4501;
wire I2287;
wire I6792;
wire I6305;
wire g1115;
wire g4512;
wire I7596;
wire I8875;
wire g1317;
wire g6287;
wire g1407;
wire g2405;
wire g4825;
wire g6715;
wire g4622;
wire g5052;
wire g3136;
wire g5908;
wire g4010;
wire g1222;
wire g5444;
wire g4706;
wire g2768;
wire g6521;
wire g5148;
wire g4874;
wire I1917;
wire g3040;
wire I2970;
wire g3618;
wire g4584;
wire g3259;
wire g3540;
wire g6299;
wire g5179;
wire g4239;
wire g5350;
wire g5475;
wire I3331;
wire I6750;
wire g3212;
wire g5375;
wire g3769;
wire I7490;
wire I8426;
wire g6258;
wire g2138;
wire I4203;
wire g847;
wire I2293;
wire I8082;
wire g3215;
wire g4630;
wire g3007;
wire g3298;
wire g5545;
wire g5374;
wire g5956;
wire g5199;
wire I2973;
wire I7856;
wire g5812;
wire g1557;
wire g6623;
wire I8696;
wire g5357;
wire g3208;
wire g6262;
wire I3488;
wire g3681;
wire I8368;
wire I3044;
wire g6231;
wire g5780;
wire g3914;
wire g2330;
wire g6123;
wire g6592;
wire g5568;
wire I8629;
wire g6336;
wire g4228;
wire I3086;
wire g4491;
wire g3913;
wire g3678;
wire g6179;
wire g6798;
wire g1724;
wire g6692;
wire I3708;
wire I6540;
wire I6692;
wire g1094;
wire g5219;
wire g6056;
wire g6489;
wire I8674;
wire I3560;
wire g3114;
wire g5164;
wire I3804;
wire I6723;
wire g6687;
wire g6901;
wire g2728;
wire g1846;
wire g4826;
wire I7346;
wire I1961;
wire g4757;
wire g5050;
wire g2086;
wire I9077;
wire g5184;
wire g3321;
wire g5794;
wire g4863;
wire I8632;
wire g3861;
wire g2670;
wire g4128;
wire g3939;
wire g6746;
wire I2763;
wire g2981;
wire g5304;
wire g4354;
wire g1979;
wire g1330;
wire g6107;
wire g4117;
wire I4681;
wire g1957;
wire I8693;
wire I5597;
wire I2457;
wire g1894;
wire g6158;
wire I5333;
wire I2306;
wire g5521;
wire g4759;
wire I2788;
wire g1345;
wire g4848;
wire I2108;
wire g6330;
wire g4714;
wire g6295;
wire g921;
wire g2650;
wire g4379;
wire g4677;
wire g5488;
wire g3622;
wire g5152;
wire g3932;
wire g3384;
wire I3152;
wire g4617;
wire g1358;
wire g6533;
wire g4123;
wire I4414;
wire g4169;
wire g6312;
wire g4797;
wire g2618;
wire g3356;
wire g2525;
wire g2242;
wire g5993;
wire I8444;
wire g5714;
wire g4059;
wire g4752;
wire I8229;
wire I3225;
wire g5060;
wire I5910;
wire g5824;
wire I1853;
wire g2695;
wire g3334;
wire g4187;
wire I2091;
wire g6657;
wire g4277;
wire g2320;
wire I2940;
wire g6357;
wire g3630;
wire g3852;
wire I4420;
wire g6645;
wire I3352;
wire g3628;
wire g4624;
wire I6015;
wire I7439;
wire g5576;
wire g1832;
wire I1832;
wire g2408;
wire g3187;
wire I3284;
wire g5667;
wire g6892;
wire g2060;
wire I5618;
wire g3770;
wire I2870;
wire I7542;
wire g5457;
wire g5265;
wire I8462;
wire I8258;
wire g4001;
wire I2593;
wire g2686;
wire I8940;
wire g6400;
wire g3806;
wire I3411;
wire I9065;
wire g5018;
wire g2659;
wire I5767;
wire g2870;
wire I5006;
wire g4599;
wire g3512;
wire I7534;
wire I2491;
wire I2967;
wire g6316;
wire g4151;
wire g1477;
wire g5551;
wire g4684;
wire g6555;
wire g2753;
wire I6185;
wire g3539;
wire I6434;
wire g4386;
wire g5292;
wire I1979;
wire g2178;
wire I9051;
wire g6115;
wire I2635;
wire g4838;
wire I3105;
wire g4146;
wire g6926;
wire I6789;
wire g6280;
wire g4373;
wire g2333;
wire g5698;
wire I6390;
wire g3533;
wire g6877;
wire g6480;
wire g3957;
wire g5939;
wire I3764;
wire g927;
wire g2955;
wire I9152;
wire g4736;
wire g6795;
wire g1205;
wire I3916;
wire g6277;
wire I6801;
wire g3287;
wire g6148;
wire g3433;
wire g5950;
wire g2367;
wire g2944;
wire g4393;
wire g4433;
wire g3847;
wire g2312;
wire g1783;
wire I8891;
wire g1627;
wire g6033;
wire g1656;
wire g6519;
wire g6100;
wire I4593;
wire I6495;
wire g5872;
wire g4132;
wire I6036;
wire g4643;
wire I8201;
wire I5307;
wire I2986;
wire g4760;
wire g2410;
wire I4331;
wire g1351;
wire g5518;
wire I6942;
wire g6567;
wire g5773;
wire I4941;
wire g3613;
wire g2105;
wire I2245;
wire g5622;
wire g6110;
wire I4398;
wire I1844;
wire I7578;
wire I4424;
wire g3365;
wire g6352;
wire I4211;
wire g2172;
wire I3161;
wire g5775;
wire g6076;
wire g1875;
wire I7966;
wire g1814;
wire I4358;
wire I7116;
wire g4341;
wire g3312;
wire I6087;
wire g5497;
wire I3004;
wire g2113;
wire I5169;
wire I3425;
wire g1030;
wire I4455;
wire I8614;
wire g3023;
wire I4226;
wire I6677;
wire I2735;
wire g5226;
wire g3014;
wire I5053;
wire g6506;
wire I6949;
wire I8779;
wire g6562;
wire g1528;
wire I1994;
wire g2156;
wire g3369;
wire g5684;
wire I2574;
wire g3162;
wire g6699;
wire g5067;
wire I2037;
wire g4158;
wire g3267;
wire I3644;
wire I3933;
wire g4946;
wire I4507;
wire I5615;
wire g4740;
wire g1966;
wire I4587;
wire g5247;
wire I8647;
wire I7799;
wire g4080;
wire I7055;
wire I5078;
wire g3300;
wire g4308;
wire I8588;
wire g6499;
wire g5953;
wire I6023;
wire g1643;
wire g2090;
wire I7487;
wire g5638;
wire g3750;
wire g2664;
wire g4434;
wire g6925;
wire g1480;
wire I6874;
wire I5388;
wire I8189;
wire g3926;
wire I5487;
wire g6446;
wire g3682;
wire g4445;
wire I2315;
wire I4150;
wire g4334;
wire g6619;
wire g5533;
wire g952;
wire g5604;
wire g2409;
wire g6160;
wire g6075;
wire g6914;
wire g2867;
wire g3336;
wire g5621;
wire g946;
wire I7238;
wire g2294;
wire I7441;
wire I5508;
wire g6730;
wire g1934;
wire g6307;
wire I5242;
wire g5895;
wire g2026;
wire g4579;
wire I5545;
wire g3659;
wire g6253;
wire g3904;
wire g900;
wire g3836;
wire I4276;
wire g1678;
wire I8220;
wire I3140;
wire g4915;
wire g1782;
wire g1329;
wire g3970;
wire g5467;
wire g2931;
wire I3258;
wire I3513;
wire g2889;
wire g1825;
wire g6910;
wire g6437;
wire g3771;
wire I6253;
wire g2827;
wire g1394;
wire g6809;
wire g1273;
wire g2117;
wire g5011;
wire g6821;
wire I4300;
wire g4058;
wire g4679;
wire I6057;
wire g6716;
wire g3881;
wire I2995;
wire I5119;
wire g4550;
wire g4537;
wire I5493;
wire g2803;
wire g3784;
wire g1943;
wire I8570;
wire g5136;
wire I3316;
wire g1326;
wire g6876;
wire g6742;
wire I5591;
wire g5889;
wire g4453;
wire I7811;
wire I6400;
wire g4364;
wire I7689;
wire g5364;
wire g4427;
wire I3212;
wire g6898;
wire g6441;
wire g6481;
wire g6457;
wire g5945;
wire g1576;
wire I5196;
wire g5662;
wire g6703;
wire g3965;
wire g4515;
wire g2790;
wire I3675;
wire g6126;
wire g6599;
wire g4802;
wire I2696;
wire g3662;
wire g2461;
wire g6620;
wire g2254;
wire g6451;
wire I2949;
wire g5431;
wire g937;
wire g804;
wire g3656;
wire I7501;
wire g3732;
wire g4405;
wire g1638;
wire g2267;
wire g3093;
wire I5351;
wire g3233;
wire g6212;
wire g4489;
wire g5951;
wire g5618;
wire g3505;
wire g4042;
wire I6132;
wire I3465;
wire g4639;
wire I3455;
wire g4779;
wire g3647;
wire I2346;
wire I5065;
wire g2921;
wire g4507;
wire g2713;
wire g2085;
wire g2214;
wire g1917;
wire I6701;
wire I7246;
wire g6609;
wire g2962;
wire g6152;
wire g6885;
wire g5066;
wire g4020;
wire g6405;
wire g2884;
wire g3679;
wire I6349;
wire g3135;
wire I3662;
wire g6634;
wire g6708;
wire g5200;
wire I3235;
wire I8984;
wire g5487;
wire I4921;
wire g2619;
wire g3237;
wire g4731;
wire g5157;
wire g5084;
wire g6415;
wire g2044;
wire I7264;
wire g6083;
wire I3398;
wire g6346;
wire g3328;
wire g4616;
wire g6513;
wire I4023;
wire g6651;
wire g3835;
wire g5504;
wire g2241;
wire I7190;
wire g5380;
wire g1333;
wire I3364;
wire g5627;
wire g4784;
wire g4685;
wire g3896;
wire g6286;
wire g1289;
wire g5232;
wire I5302;
wire g5909;
wire g6938;
wire g5192;
wire g1038;
wire I5043;
wire g5261;
wire g6789;
wire g1470;
wire I8243;
wire I4545;
wire I2507;
wire g6656;
wire I7007;
wire g1316;
wire I1865;
wire I3337;
wire I2952;
wire I8295;
wire g4510;
wire g4194;
wire I4217;
wire g4823;
wire g5865;
wire g2485;
wire I3858;
wire g4567;
wire g2009;
wire I9041;
wire g4140;
wire g5111;
wire g1221;
wire g3335;
wire g3452;
wire g3002;
wire I5188;
wire g6241;
wire g2145;
wire g3466;
wire g2437;
wire g4284;
wire g6766;
wire g6490;
wire I2527;
wire g2165;
wire I7187;
wire I2741;
wire I2131;
wire I8518;
wire I3271;
wire g5441;
wire I4050;
wire g2068;
wire g1857;
wire g5098;
wire g3875;
wire g3352;
wire g5158;
wire I7161;
wire g931;
wire g6082;
wire I3971;
wire g3464;
wire g3982;
wire g2099;
wire I6766;
wire g5975;
wire g6089;
wire I4986;
wire g1535;
wire g6777;
wire g3816;
wire I6798;
wire g1044;
wire g3960;
wire g4744;
wire g6797;
wire g4852;
wire g2391;
wire g1950;
wire I3720;
wire g2430;
wire g2950;
wire g2759;
wire g5172;
wire I8958;
wire g3759;
wire g6238;
wire I6292;
wire I3376;
wire g2842;
wire g6790;
wire I8854;
wire I7352;
wire I7339;
wire g3359;
wire g3046;
wire g985;
wire g3104;
wire I8267;
wire g5912;
wire I8120;
wire I3794;
wire I3379;
wire I3525;
wire g6713;
wire g4816;
wire g5360;
wire I8774;
wire I5568;
wire g2095;
wire I8981;
wire g5570;
wire g4021;
wire g1331;
wire g5672;
wire g3338;
wire g3322;
wire g6712;
wire g3182;
wire g6686;
wire g5605;
wire g3085;
wire I5716;
wire I2464;
wire g6646;
wire g2860;
wire g4929;
wire g4397;
wire I3215;
wire g6888;
wire g4849;
wire I2552;
wire g2920;
wire I3096;
wire I3169;
wire g3234;
wire I8249;
wire I3752;
wire g1883;
wire g3995;
wire I3188;
wire g2215;
wire I3823;
wire g5248;
wire g2256;
wire I8119;
wire I2364;
wire g6695;
wire g2997;
wire g5110;
wire g4633;
wire g6825;
wire g1036;
wire g4289;
wire I8240;
wire I7176;
wire I5761;
wire g913;
wire g2434;
wire g6461;
wire I8515;
wire g3133;
wire I8815;
wire g2029;
wire g6788;
wire g1564;
wire I5987;
wire I8678;
wire I2897;
wire I6004;
wire I8456;
wire g1423;
wire g3999;
wire I2821;
wire I3080;
wire I3382;
wire g6522;
wire g3371;
wire I3367;
wire I6867;
wire g5593;
wire I3294;
wire I7978;
wire g858;
wire g4904;
wire g1348;
wire g2061;
wire g6305;
wire I2330;
wire g5500;
wire g4051;
wire g5173;
wire g2538;
wire g3980;
wire g3575;
wire I4903;
wire I8473;
wire I8531;
wire I4382;
wire I7679;
wire I1932;
wire I2904;
wire g5890;
wire g6707;
wire I8156;
wire g1660;
wire g4793;
wire g1645;
wire I4546;
wire g1175;
wire g4656;
wire g4202;
wire I8107;
wire g6516;
wire I2703;
wire g3643;
wire I4182;
wire g3123;
wire g6469;
wire I5640;
wire g5708;
wire g4683;
wire g1474;
wire I8394;
wire g4147;
wire I9182;
wire I5439;
wire g1502;
wire g4464;
wire I8453;
wire g1047;
wire g4229;
wire g5224;
wire I3729;
wire g6170;
wire g6116;
wire g6153;
wire g6424;
wire I5360;
wire g5560;
wire I4757;
wire g3049;
wire I4019;
wire g5264;
wire I9230;
wire g3196;
wire g1731;
wire g5723;
wire g6242;
wire g5122;
wire g1650;
wire g5599;
wire I2671;
wire I3304;
wire g1671;
wire g5509;
wire I3334;
wire g5503;
wire g6324;
wire g6068;
wire g6449;
wire g4426;
wire g3625;
wire g873;
wire I8386;
wire I3848;
wire g3882;
wire g6440;
wire g1937;
wire g3503;
wire g865;
wire g3699;
wire g5873;
wire g5678;
wire I6410;
wire g2233;
wire g6933;
wire I2828;
wire g3907;
wire I5496;
wire g6127;
wire I6558;
wire g3956;
wire I3370;
wire g1570;
wire I4255;
wire g3283;
wire I8183;
wire I5890;
wire g2793;
wire g854;
wire g1416;
wire g5094;
wire g4788;
wire g3242;
wire I4220;
wire I3126;
wire g5241;
wire g3460;
wire g4514;
wire g3962;
wire g5661;
wire I2867;
wire g5860;
wire g1749;
wire I5027;
wire g5432;
wire I5293;
wire I2614;
wire g5801;
wire g6574;
wire I7239;
wire g4299;
wire g1837;
wire g1836;
wire g3665;
wire I8270;
wire g5139;
wire g1788;
wire g2968;
wire g6040;
wire g3813;
wire g4592;
wire g2599;
wire g6311;
wire I8211;
wire g4517;
wire g2973;
wire I8597;
wire g4532;
wire g3838;
wire I3876;
wire I2029;
wire I2712;
wire g4947;
wire g4250;
wire g4666;
wire I7600;
wire g4877;
wire g4322;
wire g2644;
wire g6802;
wire I3638;
wire g4521;
wire I8579;
wire I5851;
wire g4808;
wire g6408;
wire g5044;
wire I3989;
wire g6288;
wire g5220;
wire I3770;
wire g3545;
wire I9008;
wire g5017;
wire g6438;
wire I9044;
wire I3301;
wire I5536;
wire I5499;
wire g2594;
wire g3654;
wire g3199;
wire I8002;
wire g846;
wire I3065;
wire g1559;
wire g6624;
wire g4857;
wire I8527;
wire I8910;
wire g5392;
wire g6315;
wire g5886;
wire g2565;
wire I4210;
wire g5014;
wire g3940;
wire g2518;
wire g4719;
wire I7563;
wire I8878;
wire g6342;
wire I3412;
wire I2057;
wire g3484;
wire g5090;
wire g5550;
wire g5482;
wire I5502;
wire g6784;
wire g3230;
wire I4160;
wire I3155;
wire I2768;
wire g5569;
wire g3942;
wire g2932;
wire g2909;
wire g4447;
wire g3967;
wire I2814;
wire I3608;
wire g4038;
wire I5226;
wire I9050;
wire g1725;
wire g944;
wire g3520;
wire g4039;
wire g6443;
wire g3224;
wire g4766;
wire g1543;
wire g5428;
wire g1681;
wire g1323;
wire g6911;
wire g949;
wire g6165;
wire I5472;
wire I8034;
wire g4040;
wire I4498;
wire g3978;
wire g6582;
wire g1513;
wire g4133;
wire g6265;
wire g6432;
wire g4739;
wire g6904;
wire g5917;
wire I3883;
wire g4113;
wire g3063;
wire g2820;
wire I2604;
wire I3733;
wire g1858;
wire g5466;
wire g2634;
wire I5899;
wire g1624;
wire g4339;
wire I5626;
wire g1608;
wire g6359;
wire I3915;
wire g3898;
wire I3923;
wire I6930;
wire g6560;
wire g5116;
wire g4588;
wire g1037;
wire I6045;
wire g5952;
wire I1970;
wire I2929;
wire I2688;
wire g2176;
wire I6697;
wire I3288;
wire g1890;
wire g4141;
wire g3167;
wire g1670;
wire g5878;
wire I8168;
wire g3787;
wire g2890;
wire I2731;
wire I3240;
wire I7475;
wire g4050;
wire g3981;
wire g3790;
wire g6598;
wire g6875;
wire I9059;
wire g3855;
wire g3284;
wire g1542;
wire g1056;
wire I3496;
wire g1633;
wire g6625;
wire g3330;
wire I5457;
wire g3483;
wire I8773;
wire g3955;
wire g1253;
wire g1588;
wire I9107;
wire g3745;
wire I4161;
wire g6341;
wire g2108;
wire I7529;
wire g5740;
wire I1927;
wire g2010;
wire I2296;
wire I5857;
wire g6840;
wire g6608;
wire g5299;
wire g872;
wire g4183;
wire g6566;
wire g2583;
wire g1761;
wire g2922;
wire I6576;
wire I7960;
wire I7996;
wire I8843;
wire I6327;
wire g1113;
wire g5095;
wire g5677;
wire I5030;
wire g4346;
wire g6274;
wire I2301;
wire I5409;
wire g3325;
wire g2836;
wire I7035;
wire g2902;
wire g6247;
wire I6337;
wire g926;
wire I8358;
wire g2958;
wire I7564;
wire g4834;
wire g1791;
wire I3909;
wire g3906;
wire g1461;
wire g3889;
wire g2364;
wire I8103;
wire g5378;
wire g1975;
wire g5182;
wire g5731;
wire g6816;
wire g3558;
wire I8136;
wire I6672;
wire g2746;
wire g2390;
wire g3589;
wire g6128;
wire g2581;
wire g6283;
wire I8118;
wire I7119;
wire I6042;
wire g3353;
wire g2678;
wire g2603;
wire g6640;
wire g3530;
wire g4490;
wire g3479;
wire g3037;
wire g4499;
wire I3811;
wire g2940;
wire g3246;
wire g6794;
wire g2032;
wire g4686;
wire g3865;
wire g4850;
wire I4474;
wire I7270;
wire g6052;
wire g3860;
wire g5495;
wire g3849;
wire g5697;
wire g5324;
wire I3635;
wire g6832;
wire g6498;
wire I5059;
wire g4272;
wire g5577;
wire g4525;
wire I2275;
wire g2883;
wire I6607;
wire g4152;
wire I3408;
wire g1419;
wire g5065;
wire g2706;
wire g2004;
wire I2643;
wire g2575;
wire g4638;
wire g4118;
wire g3074;
wire g6527;
wire g5189;
wire I5600;
wire g2806;
wire g4041;
wire g3802;
wire g5818;
wire g1563;
wire g1422;
wire g4671;
wire I8567;
wire g2056;
wire I5217;
wire g1315;
wire g3693;
wire g5922;
wire I4234;
wire g6091;
wire g3158;
wire I9161;
wire I4303;
wire I3687;
wire I5187;
wire g4827;
wire g4640;
wire I2185;
wire I2955;
wire g3362;
wire g3642;
wire I5343;
wire I2528;
wire g5442;
wire g6296;
wire I4522;
wire I4233;
wire I8414;
wire I3546;
wire g6774;
wire g3878;
wire g1661;
wire g2757;
wire I4312;
wire I8687;
wire g6846;
wire I7208;
wire I6247;
wire I8503;
wire g1006;
wire g6778;
wire g3758;
wire g2945;
wire g6137;
wire I4783;
wire I6448;
wire g6347;
wire g6289;
wire I3274;
wire g6895;
wire g2311;
wire g1337;
wire g4232;
wire I6745;
wire g6583;
wire g6485;
wire g6412;
wire I5562;
wire I4777;
wire g6385;
wire g6591;
wire g845;
wire g3308;
wire g6182;
wire g3705;
wire g5954;
wire g6414;
wire g5314;
wire g6332;
wire g3346;
wire g1954;
wire g4022;
wire g3207;
wire g3775;
wire g1644;
wire g3844;
wire I4791;
wire I8447;
wire I3537;
wire I7110;
wire g3763;
wire g5155;
wire I6937;
wire I3310;
wire I2802;
wire g4713;
wire g784;
wire I8345;
wire g3183;
wire g5145;
wire g4707;
wire g4362;
wire g5659;
wire I2544;
wire g4410;
wire g6232;
wire I8994;
wire g5559;
wire I5551;
wire g1550;
wire g6145;
wire g3258;
wire g3935;
wire g4465;
wire g791;
wire g5664;
wire g6122;
wire g4164;
wire g5388;
wire g3723;
wire g3358;
wire I8061;
wire I5674;
wire g4861;
wire g3486;
wire g6132;
wire g5163;
wire g5474;
wire g901;
wire g3171;
wire g3296;
wire g5779;
wire g2324;
wire I5223;
wire g4578;
wire g3799;
wire g5852;
wire I2204;
wire g3425;
wire I5736;
wire g3927;
wire I4483;
wire g6397;
wire g6689;
wire g5440;
wire g6733;
wire g4034;
wire g4377;
wire I5731;
wire g6758;
wire g1255;
wire g1209;
wire g6531;
wire g2316;
wire I8349;
wire I2080;
wire g3719;
wire g3615;
wire g5212;
wire g4645;
wire g4193;
wire I6621;
wire I8282;
wire I5490;
wire g3796;
wire I3767;
wire I5904;
wire I7522;
wire g908;
wire I1958;
wire g4245;
wire g3537;
wire g4653;
wire I4547;
wire g1378;
wire g2339;
wire g6306;
wire g2872;
wire g4498;
wire I6769;
wire g6709;
wire g878;
wire g743;
wire g3996;
wire g4015;
wire g3519;
wire I3349;
wire g2506;
wire I6302;
wire g2350;
wire I2864;
wire g6580;
wire g3360;
wire g6154;
wire g4794;
wire I2935;
wire g2255;
wire g6081;
wire g4191;
wire I4528;
wire I2578;
wire I9155;
wire I5204;
wire g6474;
wire I8603;
wire g5578;
wire g5064;
wire I6111;
wire I8450;
wire I2237;
wire g5174;
wire I2658;
wire g1174;
wire I7216;
wire g5866;
wire g4655;
wire I6194;
wire g1287;
wire I9057;
wire g6826;
wire I7451;
wire g1802;
wire g3780;
wire g6348;
wire I5893;
wire I2907;
wire g6482;
wire g6318;
wire g1672;
wire g3564;
wire g4993;
wire g5598;
wire g6611;
wire g4463;
wire g6683;
wire g6337;
wire g1473;
wire I2394;
wire I4184;
wire g4691;
wire g3691;
wire g3776;
wire I7484;
wire I4170;
wire g4148;
wire g1735;
wire I8395;
wire I5848;
wire g4541;
wire I7318;
wire I3077;
wire g1793;
wire g5700;
wire g3041;
wire I1935;
wire g6912;
wire g4262;
wire I6175;
wire g5121;
wire g1636;
wire g6515;
wire g6442;
wire I4309;
wire I6343;
wire I2842;
wire g2007;
wire g6880;
wire I5923;
wire g2807;
wire g3373;
wire g3057;
wire g6425;
wire g5561;
wire g4003;
wire g6088;
wire g4504;
wire g951;
wire g5437;
wire I4671;
wire I3519;
wire g5671;
wire g6854;
wire g910;
wire I3847;
wire g4762;
wire I8210;
wire g1270;
wire g3797;
wire g4928;
wire g5481;
wire I3946;
wire g2861;
wire g2021;
wire g3086;
wire I2779;
wire I3578;
wire I2424;
wire I3090;
wire I8966;
wire g6724;
wire I3749;
wire g4687;
wire g3450;
wire I5868;
wire I4980;
wire g6073;
wire g3988;
wire g3337;
wire g4785;
wire I4504;
wire g1533;
wire g6750;
wire I2388;
wire g6927;
wire g2996;
wire I6090;
wire I6001;
wire g5751;
wire g4632;
wire I9104;
wire g6647;
wire g6787;
wire g3877;
wire g706;
wire g5903;
wire I5535;
wire I4010;
wire I1953;
wire g5566;
wire g5169;
wire g3677;
wire I6885;
wire I5445;
wire g4172;
wire g6850;
wire g6694;
wire g1647;
wire g4286;
wire g2946;
wire g6576;
wire I8329;
wire I5825;
wire I8040;
wire g5382;
wire I3826;
wire I3531;
wire g2903;
wire I4318;
wire g3350;
wire I8129;
wire g3814;
wire I8716;
wire g4486;
wire g2814;
wire g6407;
wire g2467;
wire I3445;
wire I6552;
wire g5887;
wire g1742;
wire I2021;
wire g5571;
wire g6166;
wire I7077;
wire g3424;
wire g3521;
wire g6039;
wire I5415;
wire I3251;
wire g5118;
wire g4568;
wire g6906;
wire I5244;
wire I3840;
wire g4270;
wire I4362;
wire g1232;
wire g4185;
wire g2877;
wire g6783;
wire g4440;
wire I4152;
wire g6665;
wire g3140;
wire g6188;
wire g838;
wire I8803;
wire g6834;
wire g3657;
wire g6801;
wire g4872;
wire I5478;
wire g5162;
wire g4858;
wire g3752;
wire g2914;
wire I1838;
wire g2986;
wire I6324;
wire g3528;
wire g1558;
wire g5410;
wire g5817;
wire I6743;
wire g5532;
wire g3868;
wire I3599;
wire g1994;
wire I8080;
wire g3511;
wire g2804;
wire I7981;
wire I5871;
wire g4582;
wire g2291;
wire I2584;
wire g6105;
wire g4577;
wire g4771;
wire g5398;
wire g4801;
wire g6251;
wire g943;
wire g3941;
wire I7497;
wire g5225;
wire g6487;
wire I8831;
wire g3113;
wire g4086;
wire I4249;
wire g2731;
wire I4391;
wire g2234;
wire g1680;
wire g6732;
wire g1541;
wire g716;
wire I8070;
wire g3968;
wire I5270;
wire g2121;
wire g6843;
wire g3688;
wire g6448;
wire g2347;
wire g1049;
wire g3282;
wire I5879;
wire I7434;
wire g2896;
wire g4765;
wire g3597;
wire I6772;
wire g2716;
wire I8113;
wire I3830;
wire g4516;
wire g5508;
wire g3870;
wire g4425;
wire I2817;
wire g5620;
wire g3271;
wire I5606;
wire g3231;
wire I3871;
wire g5742;
wire g3698;
wire g5502;
wire g3247;
wire I6069;
wire I5124;
wire I2169;
wire g4590;
wire I6026;
wire I2795;
wire I5463;
wire g5705;
wire g5808;
wire I2246;
wire g3850;
wire I7704;
wire I7506;
wire I8972;
wire g5091;
wire g6323;
wire g1279;
wire g2745;
wire g6573;
wire g3319;
wire g3664;
wire g4530;
wire g3635;
wire I2234;
wire g3500;
wire I3861;
wire g2967;
wire g6134;
wire g2849;
wire I7061;
wire I1877;
wire I7244;
wire g5249;
wire g5800;
wire g2643;
wire g2792;
wire g4593;
wire g5479;
wire g3235;
wire g4533;
wire g6919;
wire g4351;
wire I7969;
wire g1775;
wire g6430;
wire I4519;
wire g1689;
wire I2175;
wire g4520;
wire g5402;
wire g2422;
wire I3134;
wire g3147;
wire g4163;
wire g1789;
wire g6557;
wire I5300;
wire g4627;
wire I3572;
wire I2300;
wire g2772;
wire g6275;
wire g5683;
wire g1815;
wire g3744;
wire g2974;
wire g4950;
wire g6584;
wire g4348;
wire g3934;
wire g1114;
wire I8470;
wire g6503;
wire g1790;
wire g1585;
wire I6392;
wire g3887;
wire g923;
wire I8699;
wire g5323;
wire g6106;
wire I2379;
wire g6326;
wire g5663;
wire g1732;
wire g6793;
wire g4936;
wire I7231;
wire g1919;
wire g4251;
wire g2582;
wire I9058;
wire I3001;
wire g1760;
wire g3557;
wire g6637;
wire g6272;
wire I5269;
wire I8538;
wire I2767;
wire g4831;
wire g4780;
wire g1716;
wire g4727;
wire g3977;
wire g4487;
wire I2272;
wire g5496;
wire g5046;
wire I6537;
wire I6952;
wire I3785;
wire g3689;
wire I5040;
wire g3531;
wire g6727;
wire I7517;
wire g2957;
wire I4282;
wire g909;
wire g4589;
wire I7608;
wire g6920;
wire g6613;
wire g6658;
wire g1824;
wire I3726;
wire g6051;
wire I4477;
wire I3773;
wire g5213;
wire g2035;
wire g1320;
wire g2336;
wire I2370;
wire I6244;
wire g3225;
wire I2140;
wire g6932;
wire I2526;
wire I7637;
wire g2107;
wire g1418;
wire g5415;
wire g3604;
wire g4184;
wire g5567;
wire g5325;
wire g866;
wire I2476;
wire g1539;
wire g3170;
wire g6433;
wire g6559;
wire g3897;
wire g1756;
wire g6565;
wire I5523;
wire I7295;
wire g3099;
wire g4383;
wire g5879;
wire g5115;
wire I2919;
wire I3914;
wire g5399;
wire g3166;
wire I3232;
wire g4718;
wire g3064;
wire g839;
wire g4293;
wire g5458;
wire I6927;
wire g2097;
wire I5929;
wire g5465;
wire g2698;
wire I2445;
wire g2576;
wire I9002;
wire g4159;
wire g855;
wire g3747;
wire g6266;
wire I8991;
wire I9113;
wire g2622;
wire g2691;
wire g6264;
wire g1499;
wire g5921;
wire g3363;
wire g3285;
wire g5686;
wire g3544;
wire g2100;
wire g3954;
wire I3127;
wire g3880;
wire g4522;
wire g5558;
wire I1880;
wire I4297;
wire g1055;
wire g4400;
wire g4569;
wire g5307;
wire g6894;
wire g1878;
wire I5294;
wire g5669;
wire g3310;
wire g2276;
wire I3474;
wire g5940;
wire I2668;
wire I3681;
wire g5273;
wire I2003;
wire g6939;
wire g2170;
wire g5918;
wire g4614;
wire g4230;
wire I2162;
wire g3487;
wire g2895;
wire g2195;
wire g1042;
wire g5377;
wire g4654;
wire g1808;
wire I4706;
wire g3297;
wire g3527;
wire g4894;
wire I5469;
wire I3190;
wire g4370;
wire g5291;
wire g1997;
wire g4138;
wire g1336;
wire g3791;
wire g6233;
wire g6688;
wire g6497;
wire I3168;
wire g5278;
wire g6131;
wire g1972;
wire I3522;
wire I7701;
wire g4864;
wire I6546;
wire I1835;
wire g1363;
wire g6097;
wire g4233;
wire I8969;
wire g4131;
wire I8348;
wire g6121;
wire g4192;
wire g4244;
wire g3124;
wire g6823;
wire I3202;
wire g5383;
wire g4352;
wire I2090;
wire I4480;
wire g3781;
wire g4122;
wire I3391;
wire g4704;
wire g5146;
wire I2128;
wire g5473;
wire g6193;
wire I2543;
wire g754;
wire I8866;
wire I4183;
wire I4343;
wire g4391;
wire g5900;
wire g6062;
wire g6545;
wire I6359;
wire g6903;
wire g4347;
wire g2919;
wire I4794;
wire I2946;
wire g3762;
wire g4646;
wire g1776;
wire I9064;
wire I8668;
wire g5876;
wire g4119;
wire I8752;
wire I2060;
wire g4774;
wire g6740;
wire I8623;
wire I2355;
wire g5544;
wire g6092;
wire g3387;
wire g2822;
wire g774;
wire g3307;
wire I8600;
wire g2868;
wire g3073;
wire g6338;
wire g6590;
wire g6714;
wire g3632;
wire g4846;
wire I2041;
wire g3692;
wire g3803;
wire I7555;
wire g714;
wire g5634;
wire g3323;
wire I9140;
wire g5893;
wire I5885;
wire I8117;
wire I4513;
wire I2623;
wire g4870;
wire I2281;
wire g4455;
wire g2088;
wire I3325;
wire g1384;
wire g6297;
wire I9143;
wire g5355;
wire g6159;
wire g5447;
wire g3157;
wire g3083;
wire I1952;
wire I3388;
wire I8585;
wire g4672;
wire I5843;
wire g2443;
wire g4692;
wire I5556;
wire I5514;
wire g1691;
wire g5150;
wire g4828;
wire I7590;
wire I7311;
wire g5156;
wire I8137;
wire I8828;
wire I3115;
wire g5370;
wire I8635;
wire g6069;
wire g6773;
wire g6908;
wire g3645;
wire g2092;
wire g3786;
wire g6413;
wire I4821;
wire g4149;
wire g889;
wire I5840;
wire g5631;
wire g6528;
wire I6756;
wire I7829;
wire g1830;
wire I6959;
wire I3428;
wire g6455;
wire I2361;
wire I2453;
wire I7466;
wire I3481;
wire g5315;
wire g6525;
wire I1963;
wire g4910;
wire g6723;
wire I2193;
wire I2756;
wire I4059;
wire I5376;
wire g1324;
wire g3478;
wire g5082;
wire g1632;
wire g6445;
wire g2640;
wire I5907;
wire g1755;
wire g4437;
wire g6936;
wire g3846;
wire g6257;
wire g4688;
wire g6921;
wire g4252;
wire g4563;
wire g6249;
wire I8641;
wire g1472;
wire g6806;
wire I8217;
wire I2047;
wire g1834;
wire I6488;
wire g1294;
wire g3501;
wire g1084;
wire g3181;
wire g1688;
wire g3648;
wire I7634;
wire I3593;
wire I6139;
wire g6510;
wire I6028;
wire g4813;
wire g5600;
wire g1177;
wire g1391;
wire g5626;
wire g1551;
wire g4591;
wire I5228;
wire g4534;
wire I8186;
wire g3627;
wire g3462;
wire I3509;
wire g4519;
wire g6496;
wire g2795;
wire I9024;
wire I4688;
wire I6989;
wire g1908;
wire g5016;
wire g4741;
wire I6573;
wire I3761;
wire I4489;
wire I3499;
wire I5542;
wire g3240;
wire I7999;
wire g5092;
wire I1962;
wire g3344;
wire g6700;
wire g5403;
wire g3146;
wire g2966;
wire g5385;
wire g6851;
wire I4762;
wire g6897;
wire g5438;
wire g2817;
wire I3739;
wire g5944;
wire g6237;
wire g6080;
wire g5359;
wire g5352;
wire g4345;
wire I2887;
wire g1648;
wire g4130;
wire I3602;
wire g6508;
wire g5507;
wire I6986;
wire I8127;
wire g6317;
wire g3653;
wire g1692;
wire g4271;
wire g6615;
wire I2228;
wire I3902;
wire g4806;
wire g6907;
wire I8812;
wire g2591;
wire g942;
wire g3518;
wire g6163;
wire g4036;
wire g3667;
wire g1070;
wire g3617;
wire I2692;
wire I8385;
wire g2904;
wire g2470;
wire g1763;
wire I7284;
wire I2796;
wire g3853;
wire I9125;
wire I3550;
wire I7225;
wire I5766;
wire I5475;
wire g5480;
wire g2041;
wire I7604;
wire g4768;
wire g5884;
wire g6603;
wire g6800;
wire g6087;
wire g2905;
wire g5423;
wire g2062;
wire g1726;
wire I2337;
wire g1295;
wire I3543;
wire g4319;
wire I2231;
wire g3096;
wire g5161;
wire g5096;
wire g947;
wire g1549;
wire g852;
wire g4452;
wire g6734;
wire I7892;
wire g3304;
wire I6066;
wire g4694;
wire g5214;
wire g6737;
wire g6782;
wire g1911;
wire g6036;
wire g5114;
wire I3178;
wire I2182;
wire g2231;
wire g6820;
wire g4375;
wire g1963;
wire g3788;
wire g5311;
wire I8840;
wire g4829;
wire g5816;
wire g6917;
wire I2913;
wire I2766;
wire I6108;
wire g2738;
wire I4279;
wire g2264;
wire g4855;
wire g4032;
wire I7472;
wire g4424;
wire g3317;
wire g5572;
wire g1686;
wire I7312;
wire g895;
wire g5042;
wire g4441;
wire g851;
wire g1582;
wire I2352;
wire g2874;
wire g2120;
wire g4761;
wire g4868;
wire I3581;
wire I3255;
wire I3746;
wire g1352;
wire g2846;
wire g5899;
wire g1173;
wire g3605;
wire g3831;
wire g815;
wire g5579;
wire g2346;
wire g1417;
wire I2581;
wire g5535;
wire I8988;
wire g1157;
wire g6078;
wire g5237;
wire g3567;
wire I2082;
wire g5538;
wire g1603;
wire g5904;
wire I5448;
wire I7527;
wire g856;
wire I6250;
wire g3440;
wire g3890;
wire g5362;
wire I5259;
wire g1118;
wire g5897;
wire g4190;
wire g6648;
wire g3441;
wire I3953;
wire I8548;
wire I6118;
wire g1953;
wire g6244;
wire g4357;
wire g2284;
wire g6143;
wire g6303;
wire I9005;
wire g1819;
wire g1985;
wire I6464;
wire g3132;
wire I4375;
wire g6696;
wire g5869;
wire g6453;
wire g6575;
wire g2292;
wire I5612;
wire g5781;
wire I2848;
wire g6367;
wire g3060;
wire I5759;
wire g844;
wire g6652;
wire g6291;
wire I4133;
wire I5103;
wire I3373;
wire g5587;
wire g6786;
wire g4444;
wire I2318;
wire g2435;
wire g4776;
wire I6599;
wire I3462;
wire g3900;
wire I8359;
wire g3997;
wire g5168;
wire g4844;
wire g6928;
wire g6596;
wire I3452;
wire g4580;
wire g5580;
wire I2566;
wire I8174;
wire g4626;
wire g2821;
wire g918;
wire I1971;
wire I2745;
wire I5271;
wire g5648;
wire g5086;
wire I3278;
wire I5207;
wire g1673;
wire g6855;
wire g5190;
wire g3731;
wire I7012;
wire I3034;
wire g2327;
wire g1897;
wire g4177;
wire I9149;
wire g2760;
wire I4486;
wire I4327;
wire I2934;
wire g4016;
wire g6835;
wire g2755;
wire g6518;
wire g2871;
wire g6467;
wire I6507;
wire I2860;
wire g2862;
wire g6717;
wire g6473;
wire g5597;
wire g1285;
wire g4389;
wire g5369;
wire g3641;
wire I2050;
wire I7569;
wire g4014;
wire g4302;
wire g4735;
wire g6047;
wire I6625;
wire I6646;
wire g4280;
wire I5723;
wire g5646;
wire g3987;
wire g3351;
wire g6682;
wire g837;
wire g4745;
wire g1741;
wire g5411;
wire I3322;
wire I6680;
wire g1639;
wire g6881;
wire g1450;
wire g4074;
wire I3584;
wire g3378;
wire I7832;
wire g5615;
wire g2764;
wire g2103;
wire I6355;
wire I6308;
wire I1862;
wire I5777;
wire g4439;
wire g4369;
wire g3636;
wire g5124;
wire g3724;
wire g5590;
wire g2732;
wire g2893;
wire g1540;
wire I2022;
wire I3446;
wire g1204;
wire g4791;
wire I5148;
wire g1653;
wire g5901;
wire I7217;
wire g4528;
wire I1986;
wire I3782;
wire g6597;
wire g3173;
wire g5877;
wire g3380;
wire g3156;
wire I8332;
wire g3306;
wire g6290;
wire I7258;
wire g3765;
wire g3070;
wire g4523;
wire g6422;
wire I6753;
wire g6452;
wire g1805;
wire g5448;
wire g5556;
wire g6410;
wire I8684;
wire I5913;
wire I8194;
wire g4384;
wire I3319;
wire g5353;
wire I9236;
wire I8429;
wire I6352;
wire I7469;
wire I6330;
wire I7835;
wire I7852;
wire g4320;
wire g2163;
wire g2808;
wire g6095;
wire I6048;
wire g5920;
wire g6661;
wire g6267;
wire I6972;
wire g843;
wire g6585;
wire g3454;
wire g5175;
wire g4668;
wire g3100;
wire g4673;
wire g6520;
wire g1770;
wire g4142;
wire g6098;
wire g2840;
wire g5180;
wire I8671;
wire g1017;
wire I1951;
wire g4281;
wire g4360;
wire g5685;
wire g3964;
wire g6538;
wire I3684;
wire g3725;
wire g4125;
wire I2190;
wire I6759;
wire I8367;
wire I7859;
wire I6441;
wire g922;
wire g6722;
wire g5187;
wire g5557;
wire I5896;
wire I8978;
wire I4066;
wire I8261;
wire g1415;
wire g4651;
wire g3016;
wire g5784;
wire g3673;
wire g1739;
wire g3959;
wire g715;
wire g1936;
wire g5730;
wire g4641;
wire I6587;
wire I8509;
wire g4367;
wire I3758;
wire g6735;
wire g6353;
wire g2949;
wire g6526;
wire I2312;
wire g2838;
wire g1781;
wire I2005;
wire g2782;
wire I2137;
wire I4462;
wire g6548;
wire g3510;
wire g2947;
wire g2667;
wire g5862;
wire g4241;
wire g2788;
wire I2839;
wire g3279;
wire g2831;
wire g2927;
wire I8347;
wire g6916;
wire g6120;
wire g3294;
wire g6234;
wire g5013;
wire I3291;
wire g1339;
wire g4544;
wire I3983;
wire g4647;
wire g6791;
wire g4416;
wire I4291;
wire I6499;
wire I6500;
wire g2952;
wire I3040;
wire g1747;
wire I2159;
wire I8376;
wire g6394;
wire g4705;
wire I4198;
wire g3766;
wire g5701;
wire I6528;
wire g5484;
wire g3292;
wire g1203;
wire g4390;
wire g5543;
wire I7979;
wire g6478;
wire g1552;
wire g1257;
wire g5255;
wire I2061;
wire g4711;
wire g2436;
wire g1381;
wire g1991;
wire g2628;
wire g5270;
wire g2263;
wire g1143;
wire I2215;
wire g3103;
wire I5258;
wire I9176;
wire g2869;
wire I5397;
wire g3741;
wire g2109;
wire g5266;
wire g5455;
wire I2196;
wire I3626;
wire g1879;
wire g3226;
wire I8144;
wire g1341;
wire g3700;
wire g2378;
wire g4449;
wire g4775;
wire g1246;
wire g3079;
wire g3110;
wire g5770;
wire g4841;
wire g5229;
wire g5635;
wire g4154;
wire I4429;
wire g5300;
wire I8745;
wire g4814;
wire g6149;
wire g6564;
wire g6403;
wire g4942;
wire I8232;
wire g3789;
wire g3316;
wire g3461;
wire g1491;
wire g1646;
wire g1027;
wire g3686;
wire g1715;
wire I8226;
wire g6273;
wire g2857;
wire I3053;
wire g5023;
wire g5414;
wire g2102;
wire g3668;
wire I3590;
wire I3714;
wire g3953;
wire g5144;
wire I9203;
wire g4615;
wire g5919;
wire g3746;
wire g5368;
wire I6280;
wire g2937;
wire I4459;
wire I4176;
wire I2240;
wire g2748;
wire I3355;
wire g4296;
wire g4231;
wire g2699;
wire g6339;
wire g5941;
wire g1812;
wire g5063;
wire I9227;
wire g964;
wire g6887;
wire I5379;
wire g4301;
wire g3551;
wire g6278;
wire g5666;
wire g6103;
wire g4781;
wire I3261;
wire g5316;
wire g2457;
wire g5019;
wire I4337;
wire g6343;
wire g1823;
wire I6786;
wire g4214;
wire g2828;
wire g4167;
wire g3888;
wire g1699;
wire g3976;
wire I3281;
wire I6195;
wire g6607;
wire I1868;
wire g5728;
wire g6285;
wire g1284;
wire I2782;
wire g1109;
wire I3010;
wire g2886;
wire g4937;
wire I4189;
wire g1504;
wire I8005;
wire g2778;
wire g1054;
wire g3832;
wire I2773;
wire g6874;
wire g2194;
wire g4458;
wire g6254;
wire I8555;
wire g1106;
wire g1914;
wire I8356;
wire g4726;
wire I5324;
wire g1064;
wire g4836;
wire g2660;
wire I3422;
wire g3481;
wire I8497;
wire I9047;
wire g6192;
wire g3042;
wire I2873;
wire g3924;
wire g2360;
wire g2080;
wire g4586;
wire g3714;
wire g5348;
wire g6726;
wire I4799;
wire g2722;
wire g2397;
wire I3656;
wire g2801;
wire I3623;
wire I2165;
wire g6540;
wire g6570;
wire g3370;
wire g2604;
wire g6501;
wire g2173;
wire I5750;
wire I4465;
wire g5717;
wire I4285;
wire g766;
wire I8126;
wire I5713;
wire I2506;
wire g3863;
wire g4621;
wire g5493;
wire g5699;
wire g1902;
wire g4344;
wire g3620;
wire g4139;
wire I3022;
wire g5089;
wire g4497;
wire g2353;
wire g941;
wire g980;
wire g4037;
wire I8435;
wire g4807;
wire I8027;
wire g5425;
wire g3485;
wire g2739;
wire g3655;
wire I2269;
wire g4323;
wire I6780;
wire g2512;
wire g5534;
wire g5633;
wire g5957;
wire I2638;
wire g5581;
wire g3546;
wire I5991;
wire I5658;
wire g6161;
wire g2912;
wire g2873;
wire I5511;
wire g6061;
wire g2036;
wire g4773;
wire g2856;
wire g6836;
wire g1053;
wire g4007;
wire g3652;
wire g6769;
wire g5885;
wire g2473;
wire I2147;
wire I6470;
wire g1685;
wire I1996;
wire g5453;
wire g5328;
wire g3122;
wire g4376;
wire g3280;
wire I6425;
wire g853;
wire g2935;
wire I8459;
wire I8438;
wire g5853;
wire I7397;
wire g5430;
wire g6164;
wire g3526;
wire g896;
wire I3665;
wire I2081;
wire g6852;
wire g5113;
wire g4462;
wire I4446;
wire g1075;
wire g2081;
wire g6466;
wire g4767;
wire g3318;
wire g5097;
wire g6552;
wire g3637;
wire g6578;
wire g836;
wire I8761;
wire g905;
wire I4003;
wire g3830;
wire g6918;
wire g4442;
wire I7988;
wire I3198;
wire I2964;
wire g3303;
wire g2491;
wire g5573;
wire g3749;
wire g3134;
wire g2159;
wire g1322;
wire g2449;
wire g1787;
wire g1807;
wire g5625;
wire g5619;
wire g2394;
wire I2225;
wire I5421;
wire g5022;
wire I3144;
wire g3872;
wire I5920;
wire g1325;
wire g4423;
wire g6245;
wire g4562;
wire g2894;
wire I3177;
wire g6935;
wire I5227;
wire g1687;
wire g6702;
wire g3961;
wire g5506;
wire g4911;
wire g6495;
wire g2888;
wire I4752;
wire I7817;
wire I7164;
wire g6934;
wire g1631;
wire g1835;
wire I7404;
wire g5083;
wire g4253;
wire g1947;
wire g2317;
wire g6889;
wire g5093;
wire g1436;
wire g971;
wire g2587;
wire I2857;
wire I8617;
wire g3666;
wire I6635;
wire g5240;
wire g4535;
wire g3456;
wire g6484;
wire I7970;
wire g3702;
wire g4635;
wire I7086;
wire g6631;
wire g5861;
wire g2960;
wire g1305;
wire g4856;
wire I3553;
wire I4270;
wire I7251;
wire I8128;
wire I5106;
wire g4518;
wire g3145;
wire g1898;
wire g2580;
wire I7432;
wire g1811;
wire I5466;
wire I3343;
wire I7051;
wire g4392;
wire g1471;
wire I3875;
wire g5911;
wire g3839;
wire g2283;
wire g1666;
wire I5831;
wire g1777;
wire g2794;
wire g6256;
wire g4473;
wire g4209;
wire g5688;
wire g3331;
wire g2040;
wire g3879;
wire g729;
wire g1587;
wire I1942;
wire I6060;
wire I4527;
wire g1674;
wire g1112;
wire g5647;
wire g4721;
wire I5728;
wire g6891;
wire I5774;
wire g5645;
wire I3979;
wire I3102;
wire g5501;
wire g5043;
wire g3372;
wire g6409;
wire g3241;
wire g3730;
wire g2481;
wire I3819;
wire g2615;
wire g2598;
wire g6718;
wire g4176;
wire I2925;
wire I6737;
wire I9220;
wire I2367;
wire I8051;
wire g3448;
wire g4052;
wire I7695;
wire I4492;
wire g2747;
wire I6795;
wire g6785;
wire g4011;
wire g6537;
wire I3988;
wire g6246;
wire g6211;
wire g5472;
wire g2830;
wire g5123;
wire I9146;
wire g1849;
wire I2933;
wire g4792;
wire g6517;
wire I3868;
wire g2765;
wire g4581;
wire g4448;
wire I6397;
wire g1640;
wire g1176;
wire I5862;
wire g6325;
wire g1286;
wire g6676;
wire I3650;
wire g6418;
wire g4407;
wire I3385;
wire I8721;
wire g1503;
wire I3632;
wire I9066;
wire I3307;
wire g6831;
wire g6096;
wire I7910;
wire g2863;
wire g5419;
wire g4693;
wire g6423;
wire I3736;
wire g5902;
wire g4092;
wire g2464;
wire I6196;
wire I7218;
wire g4368;
wire g6595;
wire g6113;
wire I8387;
wire g6781;
wire g5483;
wire I7805;
wire g5167;
wire g4787;
wire g3477;
wire g4602;
wire g3974;
wire I2327;
wire I7612;
wire g4810;
wire g5361;
wire I5746;
wire g3602;
wire g1119;
wire g5691;
wire g5896;
wire g1372;
wire g3251;
wire g1612;
wire g2169;
wire g5153;
wire g5674;
wire g6649;
wire g5679;
wire g5898;
wire I4192;
wire g1048;
wire g6711;
wire g857;
wire I4441;
wire g1884;
wire g5236;
wire g2232;
wire I2760;
wire g6304;
wire I6027;
wire I3694;
wire I5529;
wire g5905;
wire I2321;
wire g3263;
wire g2998;
wire g4402;
wire g5176;
wire I8208;
wire g6653;
wire g5926;
wire I6366;
wire g4697;
wire I3189;
wire g5539;
wire I6296;
wire g4234;
wire I8252;
wire g4261;
wire I2411;
wire g3449;
wire g5015;
wire I8749;
wire g4815;
wire g4243;
wire g4618;
wire g3339;
wire I3791;
wire g3709;
wire g4198;
wire g5384;
wire g2433;
wire I3972;
wire g6292;
wire g5658;
wire g4843;
wire g6602;
wire I7865;
wire g5891;
wire g4659;
wire I8690;
wire g4358;
wire g4496;
wire g1449;
wire g4903;
wire g3764;
wire g5997;
wire g4799;
wire g3108;
wire I1859;
wire g5371;
wire g5809;
wire I4354;
wire g4862;
wire g5783;
wire g6873;
wire I3797;
wire I4534;
wire g2308;
wire g2837;
wire g4652;
wire g6146;
wire g5753;
wire g2928;
wire g4642;
wire g6772;
wire g2789;
wire g2154;
wire g5549;
wire g3015;
wire I3062;
wire I8346;
wire g4869;
wire I3808;
wire g3694;
wire g4648;
wire g3525;
wire g3295;
wire I8758;
wire g6235;
wire I8135;
wire g3819;
wire g4165;
wire g1764;
wire g5490;
wire g1649;
wire I6946;
wire g3614;
wire I2044;
wire g6882;
wire g5235;
wire g6060;
wire I7276;
wire I6501;
wire g3216;
wire I8342;
wire I6176;
wire g4860;
wire g3305;
wire g2679;
wire g3798;
wire g6612;
wire g5616;
wire g4153;
wire I5854;
wire g6762;
wire I2110;
wire g1338;
wire g4242;
wire g1748;
wire I2154;
wire I2376;
wire I7494;
wire g5636;
wire I2089;
wire g6502;
wire g3388;
wire I2309;
wire g3172;
wire I8357;
wire g4495;
wire g3843;
wire I5577;
wire g5542;
wire g3866;
wire g4359;
wire g5720;
wire g3899;
wire I3836;
wire I2497;
wire g4235;
wire g4822;
wire g4350;
wire g1256;
wire g6194;
wire I2460;
wire g4867;
wire g1156;
wire g917;
wire I1850;
wire I4264;
wire I7557;
wire g5354;
wire g3536;
wire g6833;
wire I8662;
wire I6012;
wire I1847;
wire g2809;
wire g6369;
wire g2976;
wire g2110;
wire g5471;
wire I4235;
wire I2212;
wire g3482;
wire g5596;
wire g5564;
wire I5649;
wire g4529;
wire g6067;
wire I8943;
wire g1771;
wire g3727;
wire I5157;
wire g1806;
wire g6411;
wire g2574;
wire g3634;
wire I9167;
wire g3012;
wire I2402;
wire g6539;
wire g3801;
wire I8506;
wire I6382;
wire I3016;
wire g3910;
wire I4782;
wire g1193;
wire g2841;
wire g4224;
wire I5699;
wire g6721;
wire g5555;
wire g4143;
wire g3856;
wire I2831;
wire I9217;
wire I3611;
wire g3793;
wire g3455;
wire g6905;
wire g2245;
wire g3219;
wire I3672;
wire g3800;
wire I5002;
wire g2948;
wire I3563;
wire g6344;
wire g3599;
wire I6744;
wire g3155;
wire g4223;
wire g1189;
wire g6586;
wire g3998;
wire g5188;
wire g5154;
wire g4674;
wire I6564;
wire g4753;
wire g2700;
wire I4306;
wire g4124;
wire I7520;
wire g6090;
wire I6075;
wire I7349;
wire g6331;
wire g6104;
wire g1738;
wire g3975;
wire g3621;
wire I5352;
wire g4361;
wire g4215;
wire g6328;
wire I6020;
wire g2685;
wire g2885;
wire g6606;
wire I2648;
wire I3431;
wire I3890;
wire g6043;
wire I5182;
wire g5665;
wire g4431;
wire I3705;
wire g1730;
wire g4612;
wire g2381;
wire I2414;
wire I5391;
wire g1740;
wire g6725;
wire g4300;
wire I3025;
wire g3559;
wire g829;
wire I6689;
wire g5181;
wire g5317;
wire g3204;
wire g4770;
wire I3170;
wire I7045;
wire I5657;
wire g6428;
wire g4938;
wire g5420;
wire I7980;
wire g2361;
wire g3345;
wire g6354;
wire g5349;
wire g6479;
wire I3179;
wire g2637;
wire g6509;
wire g2101;
wire I2570;
wire g5727;
wire I2125;
wire g6532;
wire I3447;
wire g2829;
wire g6643;
wire I6430;
wire g5470;
wire g2488;
wire g4943;
wire I8702;
wire g2770;
wire g4049;
wire g1107;
wire g4782;
wire g4171;
wire I6039;
wire g4629;
wire g3043;
wire g4587;
wire g4273;
wire g2951;
wire g4166;
wire g6922;
wire g5494;
wire g5938;
wire I8869;
wire I5337;
wire I5739;
wire g5215;
wire g3278;
wire g1754;
wire I3125;
wire g5088;
wire g2142;
wire g3324;
wire I3895;
wire g4033;
wire I7107;
wire I5033;
wire g6270;
wire g4485;
wire g4438;
wire I6555;
wire I9134;
wire I4976;
wire g5456;
wire g5296;
wire g4833;
wire g3925;
wire I1987;
wire I3605;
wire g6320;
wire I8710;
wire I2033;
wire I7990;
wire g4620;
wire I2115;
wire g1142;
wire I2808;
wire g4980;
wire g2031;
wire I7989;
wire g6404;
wire I8482;
wire I3405;
wire g3361;
wire I3886;
wire g6581;
wire g3227;
wire g5702;
wire I5050;
wire g2266;
wire I4664;
wire g3293;
wire g6719;
wire g3952;
wire g3740;
wire g3381;
wire g1340;
wire g1623;
wire g3739;
wire I7146;
wire g6749;
wire g1263;
wire I8767;
wire I8223;
wire I8162;
wire I5257;
wire g3687;
wire g6079;
wire g1101;
wire g4398;
wire g3810;
wire g6375;
wire g4381;
wire I7814;
wire g1792;
wire I4294;
wire g6929;
wire I7643;
wire g3349;
wire g6845;
wire g1254;
wire g4199;
wire g1355;
wire g842;
wire I3587;
wire g4182;
wire g6119;
wire g6129;
wire g1714;
wire g6610;
wire g3979;
wire I8485;
wire g3281;
wire g4000;
wire I2588;
wire g5194;
wire I8377;
wire g2783;
wire g6563;
wire g6819;
wire I7361;
wire g2197;
wire g4859;
wire g2756;
wire g4680;
wire I5977;
wire g4450;
wire g5024;
wire g5367;
wire g5942;
wire g3774;
wire g2779;
wire I5292;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g678 <= 0;
  else
    g678 <= g4130;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g332 <= 0;
  else
    g332 <= g6823;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g123 <= 0;
  else
    g123 <= g6940;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g207 <= 0;
  else
    g207 <= g6102;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g695 <= 0;
  else
    g695 <= g4147;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g461 <= 0;
  else
    g461 <= g4841;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g18 <= 0;
  else
    g18 <= g6725;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g292 <= 0;
  else
    g292 <= g3232;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g331 <= 0;
  else
    g331 <= g4119;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g689 <= 0;
  else
    g689 <= g4141;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g24 <= 0;
  else
    g24 <= g6726;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g465 <= 0;
  else
    g465 <= g6507;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g84 <= 0;
  else
    g84 <= g6590;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g291 <= 0;
  else
    g291 <= g3231;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g676 <= 0;
  else
    g676 <= g5330;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g622 <= 0;
  else
    g622 <= g5147;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g117 <= 0;
  else
    g117 <= g4839;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g278 <= 0;
  else
    g278 <= g6105;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g128 <= 0;
  else
    g128 <= g5138;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g598 <= 0;
  else
    g598 <= g4122;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g554 <= 0;
  else
    g554 <= g6827;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g496 <= 0;
  else
    g496 <= g6745;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g179 <= 0;
  else
    g179 <= g6405;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g48 <= 0;
  else
    g48 <= g6729;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g590 <= 0;
  else
    g590 <= g6595;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g551 <= 0;
  else
    g551 <= g6826;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g682 <= 0;
  else
    g682 <= g4134;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g11 <= 0;
  else
    g11 <= g6599;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g606 <= 0;
  else
    g606 <= g4857;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g188 <= 0;
  else
    g188 <= g6406;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g646 <= 0;
  else
    g646 <= g5148;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g327 <= 0;
  else
    g327 <= g4117;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g361 <= 0;
  else
    g361 <= g6582;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g289 <= 0;
  else
    g289 <= g3229;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g398 <= 0;
  else
    g398 <= g5700;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g684 <= 0;
  else
    g684 <= g4136;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g619 <= 0;
  else
    g619 <= g4858;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g208 <= 0;
  else
    g208 <= g5876;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g248 <= 0;
  else
    g248 <= g3239;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g390 <= 0;
  else
    g390 <= g5698;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g625 <= 0;
  else
    g625 <= g5328;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g681 <= 0;
  else
    g681 <= g4133;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g437 <= 0;
  else
    g437 <= g4847;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g276 <= 0;
  else
    g276 <= g5877;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3 <= 0;
  else
    g3 <= g6597;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g323 <= 0;
  else
    g323 <= g4120;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g224 <= 0;
  else
    g224 <= g3235;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g685 <= 0;
  else
    g685 <= g4137;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g43 <= 0;
  else
    g43 <= g6407;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g157 <= 0;
  else
    g157 <= g5470;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g282 <= 0;
  else
    g282 <= g6841;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g697 <= 0;
  else
    g697 <= g4149;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g206 <= 0;
  else
    g206 <= g6101;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g449 <= 0;
  else
    g449 <= g4844;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g118 <= 0;
  else
    g118 <= g4113;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g528 <= 0;
  else
    g528 <= g6504;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g284 <= 0;
  else
    g284 <= g3224;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g426 <= 0;
  else
    g426 <= g4855;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g634 <= 0;
  else
    g634 <= g4424;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g669 <= 0;
  else
    g669 <= g5582;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g520 <= 0;
  else
    g520 <= g6502;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g281 <= 0;
  else
    g281 <= g6107;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g175 <= 0;
  else
    g175 <= g5472;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g15 <= 0;
  else
    g15 <= g6602;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g631 <= 0;
  else
    g631 <= g5581;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g69 <= 0;
  else
    g69 <= g6587;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g693 <= 0;
  else
    g693 <= g4145;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g337 <= 0;
  else
    g337 <= g2585;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g457 <= 0;
  else
    g457 <= g4842;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g486 <= 0;
  else
    g486 <= g2586;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g471 <= 0;
  else
    g471 <= g1291;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g328 <= 0;
  else
    g328 <= g4118;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g285 <= 0;
  else
    g285 <= g3225;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g418 <= 0;
  else
    g418 <= g4853;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g402 <= 0;
  else
    g402 <= g4849;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g297 <= 0;
  else
    g297 <= g6512;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g212 <= 0;
  else
    g212 <= g3233;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g410 <= 0;
  else
    g410 <= g4851;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g430 <= 0;
  else
    g430 <= g4856;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g33 <= 0;
  else
    g33 <= g6854;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g662 <= 0;
  else
    g662 <= g1831;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g453 <= 0;
  else
    g453 <= g4843;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g269 <= 0;
  else
    g269 <= g6510;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g574 <= 0;
  else
    g574 <= g6591;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g441 <= 0;
  else
    g441 <= g4846;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g664 <= 0;
  else
    g664 <= g1288;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g349 <= 0;
  else
    g349 <= g5478;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g211 <= 0;
  else
    g211 <= g6840;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g586 <= 0;
  else
    g586 <= g6594;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g571 <= 0;
  else
    g571 <= g5580;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g29 <= 0;
  else
    g29 <= g6853;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g326 <= 0;
  else
    g326 <= g4840;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g698 <= 0;
  else
    g698 <= g4150;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g654 <= 0;
  else
    g654 <= g5490;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g293 <= 0;
  else
    g293 <= g6511;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g690 <= 0;
  else
    g690 <= g4142;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g445 <= 0;
  else
    g445 <= g4845;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g374 <= 0;
  else
    g374 <= g5694;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6 <= 0;
  else
    g6 <= g6722;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g687 <= 0;
  else
    g687 <= g4139;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g357 <= 0;
  else
    g357 <= g5480;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g386 <= 0;
  else
    g386 <= g5697;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g504 <= 0;
  else
    g504 <= g6498;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g665 <= 0;
  else
    g665 <= g4126;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g166 <= 0;
  else
    g166 <= g5471;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g541 <= 0;
  else
    g541 <= g6505;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g74 <= 0;
  else
    g74 <= g6588;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g338 <= 0;
  else
    g338 <= g5475;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g696 <= 0;
  else
    g696 <= g4148;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g516 <= 0;
  else
    g516 <= g6501;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g536 <= 0;
  else
    g536 <= g6506;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g683 <= 0;
  else
    g683 <= g4135;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g353 <= 0;
  else
    g353 <= g5479;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g545 <= 0;
  else
    g545 <= g6824;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g254 <= 0;
  else
    g254 <= g3240;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g341 <= 0;
  else
    g341 <= g5476;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g290 <= 0;
  else
    g290 <= g3230;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2 <= 0;
  else
    g2 <= g6721;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g287 <= 0;
  else
    g287 <= g3227;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g336 <= 0;
  else
    g336 <= g6925;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g345 <= 0;
  else
    g345 <= g5477;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g628 <= 0;
  else
    g628 <= g5489;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g679 <= 0;
  else
    g679 <= g4131;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g28 <= 0;
  else
    g28 <= g6727;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g688 <= 0;
  else
    g688 <= g4140;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g283 <= 0;
  else
    g283 <= g6842;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g613 <= 0;
  else
    g613 <= g4423;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g10 <= 0;
  else
    g10 <= g6723;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g14 <= 0;
  else
    g14 <= g6724;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g680 <= 0;
  else
    g680 <= g4132;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g143 <= 0;
  else
    g143 <= g6401;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g672 <= 0;
  else
    g672 <= g5491;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g667 <= 0;
  else
    g667 <= g4127;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g366 <= 0;
  else
    g366 <= g6278;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g279 <= 0;
  else
    g279 <= g6106;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g492 <= 0;
  else
    g492 <= g6744;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g170 <= 0;
  else
    g170 <= g6404;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g686 <= 0;
  else
    g686 <= g4138;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g288 <= 0;
  else
    g288 <= g3228;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g638 <= 0;
  else
    g638 <= g1289;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g602 <= 0;
  else
    g602 <= g4123;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g642 <= 0;
  else
    g642 <= g4658;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g280 <= 0;
  else
    g280 <= g5878;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g663 <= 0;
  else
    g663 <= g4125;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g610 <= 0;
  else
    g610 <= g4124;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g148 <= 0;
  else
    g148 <= g5874;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g209 <= 0;
  else
    g209 <= g6103;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g675 <= 0;
  else
    g675 <= g1294;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g478 <= 0;
  else
    g478 <= g1292;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g122 <= 0;
  else
    g122 <= g4115;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g54 <= 0;
  else
    g54 <= g6584;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g594 <= 0;
  else
    g594 <= g6596;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g286 <= 0;
  else
    g286 <= g3226;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g489 <= 0;
  else
    g489 <= g2587;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g616 <= 0;
  else
    g616 <= g4657;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g79 <= 0;
  else
    g79 <= g6589;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g218 <= 0;
  else
    g218 <= g3234;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g242 <= 0;
  else
    g242 <= g3238;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g578 <= 0;
  else
    g578 <= g6592;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g184 <= 0;
  else
    g184 <= g5473;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g119 <= 0;
  else
    g119 <= g4114;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g668 <= 0;
  else
    g668 <= g6800;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g139 <= 0;
  else
    g139 <= g5141;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g422 <= 0;
  else
    g422 <= g4854;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g210 <= 0;
  else
    g210 <= g6839;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g394 <= 0;
  else
    g394 <= g5699;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g230 <= 0;
  else
    g230 <= g3236;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g25 <= 0;
  else
    g25 <= g6601;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g204 <= 0;
  else
    g204 <= g5875;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g658 <= 0;
  else
    g658 <= g4425;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g650 <= 0;
  else
    g650 <= g5329;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g378 <= 0;
  else
    g378 <= g5695;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g508 <= 0;
  else
    g508 <= g6499;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g548 <= 0;
  else
    g548 <= g6825;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g370 <= 0;
  else
    g370 <= g5693;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g406 <= 0;
  else
    g406 <= g4850;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g236 <= 0;
  else
    g236 <= g3237;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g500 <= 0;
  else
    g500 <= g6497;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g205 <= 0;
  else
    g205 <= g6100;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g197 <= 0;
  else
    g197 <= g6509;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g666 <= 0;
  else
    g666 <= g4128;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g114 <= 0;
  else
    g114 <= g4116;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g524 <= 0;
  else
    g524 <= g6503;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g260 <= 0;
  else
    g260 <= g3241;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g111 <= 0;
  else
    g111 <= g6277;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g131 <= 0;
  else
    g131 <= g5139;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g7 <= 0;
  else
    g7 <= g6598;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g19 <= 0;
  else
    g19 <= g6600;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g677 <= 0;
  else
    g677 <= g4129;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g582 <= 0;
  else
    g582 <= g6593;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g485 <= 0;
  else
    g485 <= g6801;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g699 <= 0;
  else
    g699 <= g4426;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g193 <= 0;
  else
    g193 <= g5474;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g135 <= 0;
  else
    g135 <= g5140;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g382 <= 0;
  else
    g382 <= g5696;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g414 <= 0;
  else
    g414 <= g4852;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g434 <= 0;
  else
    g434 <= g4848;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g266 <= 0;
  else
    g266 <= g4659;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g49 <= 0;
  else
    g49 <= g6583;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g152 <= 0;
  else
    g152 <= g6402;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g692 <= 0;
  else
    g692 <= g4144;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g277 <= 0;
  else
    g277 <= g6104;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g127 <= 0;
  else
    g127 <= g6941;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g161 <= 0;
  else
    g161 <= g6403;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g512 <= 0;
  else
    g512 <= g6500;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g532 <= 0;
  else
    g532 <= g6508;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g64 <= 0;
  else
    g64 <= g6586;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g694 <= 0;
  else
    g694 <= g4146;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g691 <= 0;
  else
    g691 <= g4143;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1 <= 0;
  else
    g1 <= g6720;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g59 <= 0;
  else
    g59 <= g6585;
assign g2171 = ((~I3304));
assign I2596 = ((~g985));
assign g3491 = ((~g2608));
assign g3610 = (g2397&g3034);
assign g4355 = (g430&g3778);
assign I8764 = ((~g6564));
assign g6579 = ((~g6490));
assign I3711 = ((~g1848));
assign g4610 = ((~I6186))|((~I6187));
assign g3277 = (g2174&g2625);
assign g3892 = ((~g3575));
assign g4396 = (g422&g3801);
assign g4866 = (g4756)|(g4491);
assign g6365 = ((~I8159));
assign g3783 = ((~I4980));
assign g3603 = (g2370&g3019);
assign g4111 = ((~I5415));
assign I5793 = ((~g3803));
assign g2887 = ((~g1858));
assign I5743 = ((~g4022));
assign g6136 = ((~I7856));
assign g1276 = ((~g847));
assign I8494 = ((~g6428));
assign g3885 = ((~I5124));
assign g1946 = ((~I3053));
assign g6034 = ((~g5824));
assign g3034 = ((~I4249));
assign g4847 = ((~I6549));
assign I9085 = ((~g6850));
assign g2776 = ((~g2378));
assign I4667 = ((~g2908));
assign g6542 = ((~I8538));
assign g6426 = (g6288)|(g6119);
assign I7463 = ((~g5622));
assign g5729 = ((~I7494));
assign g6561 = ((~I8567));
assign I4452 = ((~g2117));
assign I7963 = ((~g6276));
assign g2039 = ((~I3148));
assign g5788 = ((~I7587));
assign g6293 = (g6244)|(g6085);
assign g6577 = ((~g6488));
assign g5711 = ((~I7472));
assign I4678 = ((~g2670));
assign I5517 = ((~g3885));
assign I8872 = ((~g6695));
assign I6923 = ((~g5124));
assign g5925 = ((~I7707));
assign g5805 = ((~I7604));
assign g5216 = (g563&g5025);
assign g1110 = ((~I2140));
assign I7333 = ((~g5386));
assign I8491 = ((~g6480));
assign g5025 = ((~g4814));
assign I2753 = ((~g1174));
assign g5119 = ((~I6769));
assign g2098 = ((~g1363));
assign g5099 = ((~I6737));
assign I5526 = ((~g3848));
assign I2479 = ((~g1049));
assign I4961 = ((~g3597));
assign g4342 = (g3978&g3299);
assign g4623 = ((~g4262));
assign g3150 = ((~I4391));
assign g5445 = ((~g5274));
assign g5778 = ((~I7542))|((~I7543));
assign I2442 = ((~g872));
assign g3864 = (g3693)|(g3176);
assign g4432 = ((~g923)&(~g4253));
assign g736 = ((~I1841));
assign g3761 = ((~g3605));
assign I2299 = ((~g830))|((~g341));
assign g4157 = (g3830&g1533);
assign g5680 = (g5562)|(g5429);
assign g4835 = (g4533&g4530);
assign g4136 = ((~I5490));
assign g1628 = (g815&g809);
assign g6544 = ((~I8544));
assign I4173 = ((~g2408));
assign g4276 = ((~I5731));
assign I3556 = ((~g1484));
assign I2150 = ((~g10));
assign g6419 = ((~I8267));
assign g2535 = ((~I3653));
assign I4526 = ((~g2909))|((~g646));
assign I3298 = ((~g1725));
assign g3554 = (g2941&g179);
assign I8335 = ((~g6308));
assign I5195 = ((~g3567))|((~g3571));
assign g6358 = ((~I8126)&(~I8127)&(~I8128)&(~I8129));
assign g2416 = ((~I3556));
assign I2738 = ((~g1236));
assign I8821 = ((~g6691));
assign I2845 = ((~g1193));
assign g6261 = (g5673)|(g5944);
assign g1387 = ((~g862))|((~g314))|((~g301));
assign g3366 = (g248&g2893);
assign I8564 = ((~g6429));
assign g3638 = ((~g3108));
assign g4236 = (g654&g3907);
assign g2859 = (g2112&g1649);
assign g3534 = ((~I4752));
assign I9031 = ((~g6809));
assign I8393 = (g6317)|(g6130)|(g6133)|(g6151);
assign g5498 = (g5449&g3460);
assign g1589 = (g1059)|(g1045);
assign I7039 = ((~g5309));
assign g5874 = ((~I7634));
assign I8209 = (g6015)|(g6212)|(g4950)|(g4877);
assign g4401 = (g426&g3802);
assign I7571 = ((~g5678))|((~I7569));
assign g6890 = ((~I9137));
assign g940 = ((~g64));
assign I6371 = ((~g4569));
assign g2135 = ((~I3261));
assign g3670 = (g2234&g2792);
assign g6114 = (g5904)|(g5604);
assign g3922 = ((~I5157));
assign g4454 = (g4395)|(g4051);
assign g1822 = ((~g1070))|((~g1084));
assign g6847 = (g5861)|(g6837);
assign g6818 = ((~I8991));
assign g5491 = ((~I7193));
assign g1063 = ((~g675));
assign g4830 = (g4529&g4525);
assign g6015 = ((~g5857));
assign I5433 = ((~g3728));
assign I7692 = ((~g5711));
assign g1206 = ((~I2212));
assign I3894 = ((~g286))|((~I3893));
assign g5726 = ((~I7487));
assign g6853 = ((~I9082));
assign I7906 = ((~g5912));
assign g2177 = ((~I3322));
assign g4150 = ((~I5532));
assign g3029 = ((~I4240));
assign I6660 = ((~g4762))|((~I6659));
assign g1925 = ((~I3028));
assign g6827 = ((~I9014));
assign I5603 = ((~g3893));
assign g835 = ((~g345));
assign g4811 = (g4429)|(g4432);
assign g5673 = (g59&g5573);
assign I9116 = ((~g6864));
assign I5023 = ((~g3263));
assign g5329 = ((~I6989));
assign I8196 = ((~g6188))|((~I8194));
assign g5295 = (g5047)|(g4766);
assign I2449 = ((~g971));
assign g6743 = ((~I8907));
assign g6101 = ((~I7799));
assign I7481 = ((~g5629));
assign g3067 = ((~I4294));
assign g3748 = (g3366)|(g2782);
assign g1841 = ((~I2929));
assign I9128 = ((~g6864));
assign g4854 = ((~I6570));
assign I7987 = (g6194)|(g5958)|(g5975)|(g5997);
assign g1829 = ((~I2898))|((~I2899));
assign g6279 = ((~I7969)&(~I7970)&(~I7971)&(~I7972));
assign g6605 = ((~I8681));
assign I9179 = ((~g6875));
assign I3019 = ((~g1755));
assign g5318 = ((~g676))|((~g5060));
assign g6879 = ((~I9104));
assign I6318 = ((~g4447));
assign g6837 = ((~g6822));
assign g6594 = ((~I8650));
assign g6494 = ((~g952)&(~g6348));
assign g3598 = (g2808)|(g2821);
assign I8713 = ((~g6522));
assign g6155 = (g2588&g5997);
assign I6895 = ((~g5010));
assign g1369 = ((~I2405));
assign I5233 = ((~g3571));
assign I8202 = ((~g478))|((~I8201));
assign g5602 = (g594&g5515);
assign I2521 = ((~g1063));
assign I3137 = ((~g1315));
assign I7509 = ((~g5587));
assign g2087 = ((~g1352));
assign g893 = ((~g23));
assign I8370 = (g5214)|(g6358);
assign g6923 = (g6918&g6917);
assign I2716 = ((~g1115));
assign g6333 = (g3896&g6212);
assign g2709 = ((~I3864));
assign g2315 = ((~I3465));
assign g6108 = (g5898)|(g5598);
assign I2420 = ((~g791));
assign g809 = ((~I1874));
assign g5694 = (g5633)|(g5482);
assign g6142 = (g5909)|(g3806);
assign g5135 = ((~I6783));
assign I8110 = ((~g6143));
assign g3755 = (g2604&g3481);
assign I8285 = ((~g6310));
assign g2018 = (g1423&g1254);
assign g5363 = (g4439&g5179);
assign I2073 = ((~g15))|((~I2072));
assign g3848 = ((~I5059));
assign g3128 = ((~I4375));
assign g6364 = ((~I8156));
assign g1567 = ((~I2537));
assign I6386 = ((~g4462));
assign g6587 = ((~I8629));
assign g1784 = (g858&g889);
assign g3931 = ((~g3353)&(~g3361));
assign g3200 = ((~I4437));
assign g5185 = (g524&g4993);
assign g4459 = (g4245&g1899);
assign g6549 = (g6473)|(g4247);
assign g4717 = ((~g4465));
assign I6093 = ((~g4394));
assign g6523 = ((~I8485));
assign g3342 = ((~g3086));
assign I2179 = ((~g293));
assign I3534 = ((~g1295));
assign g4068 = (g3293)|(g2685);
assign g4127 = ((~I5463));
assign g4526 = ((~I6090));
assign g1813 = ((~I2870));
assign g4144 = ((~I5514));
assign g5947 = ((~g5821))|((~g2944));
assign g1366 = ((~I2402));
assign g5946 = ((~g5729));
assign g1982 = ((~I3093));
assign I7433 = ((~g111))|((~I7432));
assign g3619 = (g2449&g3057);
assign g1344 = ((~I2379));
assign g5935 = (g5112&g5784);
assign g2780 = ((~I3971))|((~I3972));
assign g6086 = (g1143&g5742);
assign g4619 = ((~g4248));
assign I3434 = ((~g1627));
assign I9011 = ((~g6819));
assign I6456 = ((~g4633));
assign I3056 = ((~g1519));
assign g2941 = (g2166&g170);
assign I3855 = ((~g2550));
assign I8653 = ((~g6531));
assign g4644 = ((~I6231));
assign g3990 = (g3684)|(g3155);
assign I8626 = ((~g6543));
assign g2727 = ((~g2324));
assign g2340 = (g1398&g1387);
assign I2343 = ((~g1177));
assign I2499 = ((~g1036))|((~I2497));
assign g3851 = (g3681)|(g3146);
assign g2307 = ((~I3446))|((~I3447));
assign g3333 = (g2264&g2728);
assign g3154 = (g2039&g1410);
assign g4756 = (g3816&g4587);
assign g3936 = (g3551&g940);
assign g6556 = (g6339)|(g6467);
assign I4684 = ((~g2687));
assign g4114 = ((~I5424));
assign g3646 = (g2179&g2756);
assign I5944 = ((~g4356));
assign g1192 = ((~g44));
assign g3013 = ((~I4211))|((~I4212));
assign g1665 = ((~g985));
assign g3701 = (g2268&g2838);
assign I2728 = ((~g1232));
assign g4634 = (g4341)|(g3615);
assign I8378 = (g5173)|(g5166)|(g5235)|(g5245);
assign g5478 = ((~I7170));
assign g4839 = ((~I6525));
assign I6311 = ((~g4444));
assign g6822 = ((~g6786));
assign g2767 = ((~g2364));
assign g6401 = ((~I8217));
assign I8056 = ((~g6109));
assign I3358 = ((~g1323));
assign I3620 = ((~g1484));
assign g1922 = ((~I3025));
assign I7593 = ((~g5605));
assign I5783 = ((~g3810))|((~I5782));
assign I4008 = ((~g292))|((~g2568));
assign I4246 = ((~g2194));
assign g5958 = ((~g5818));
assign g4699 = ((~I6289));
assign g5512 = ((~I7254));
assign I5708 = ((~g3942));
assign g4461 = (g4241&g2919);
assign I2284 = ((~g922));
assign g4168 = (g3925&g1355);
assign g6488 = ((~g6367));
assign g4720 = ((~I6340));
assign g6150 = (g3204&g6015);
assign I2608 = ((~g1143));
assign I7143 = ((~g5323));
assign g5489 = ((~I7187));
assign g6269 = (g524&g5908);
assign g3869 = (g3642)|(g3650);
assign I3068 = ((~g1439));
assign g3109 = ((~g2360))|((~g1064));
assign I8800 = ((~g6684));
assign I3028 = ((~g1504));
assign g2688 = ((~I3836));
assign g4178 = (g3959&g2110);
assign I8837 = ((~g6665));
assign I8369 = (g5165)|(g5159)|(g5233)|(g5240);
assign g1853 = ((~I2955));
assign g3768 = (g3448&g1528);
assign I5702 = ((~g3845));
assign I4646 = ((~g2602));
assign I3244 = ((~g1772));
assign g965 = ((~I2033));
assign I4204 = ((~g2255))|((~I4203));
assign g3382 = (g3136&g2934);
assign I5505 = ((~g3860));
assign g5141 = ((~I6801));
assign g2157 = ((~I3278));
assign g1695 = ((~g1106));
assign g2954 = ((~g2381));
assign g5541 = ((~g5388)&(~g1880));
assign I8089 = ((~g6120));
assign g5198 = (g558&g5025);
assign g3912 = ((~g3505));
assign g6691 = (g6275)|(g6603);
assign g3973 = ((~g3368)&(~g3374));
assign I6543 = ((~g4718));
assign I7440 = ((~g5515))|((~I7439));
assign I1980 = ((~g230))|((~I1978));
assign g2356 = (g1603&g269);
assign g5269 = (g557&g5025);
assign g4600 = (g4054&g4289);
assign g6065 = ((~g5784));
assign I4340 = ((~g1935));
assign g5629 = (g5499)|(g3298);
assign g6536 = ((~I8524));
assign g6055 = (g5824&g1696);
assign g4266 = ((~g3757)&(~g3283));
assign g3778 = ((~g3388));
assign g4702 = ((~I6296));
assign g1861 = ((~I2967));
assign g2078 = ((~g1345));
assign I8946 = ((~g6778));
assign I6177 = ((~g571))|((~I6175));
assign I3485 = ((~g1450));
assign g2915 = ((~g1931));
assign g4120 = ((~I5442));
assign g5373 = (g161&g5250);
assign I5427 = ((~g3726));
assign g1847 = ((~I2943));
assign g3958 = ((~g3316)&(~g3326));
assign g3807 = ((~I5006));
assign g6900 = ((~I9167));
assign g5074 = (g4792)|(g4598);
assign g6147 = ((~I7871));
assign g2112 = ((~I3240));
assign g6093 = (g1177&g5742);
assign g4603 = ((~I6170));
assign g6185 = (g6055)|(g5995);
assign I8066 = ((~g6114));
assign g2733 = (g2422&g1943);
assign I6612 = ((~g4660));
assign g2876 = ((~g1943));
assign I2023 = ((~g254))|((~I2021));
assign g5565 = ((~I7312))|((~I7313));
assign I5720 = ((~g4022));
assign g932 = ((~g337));
assign g1675 = ((~g1101));
assign I2278 = ((~g917));
assign I5460 = ((~g3771));
assign I4166 = ((~g2390));
assign g6371 = ((~I8177));
assign I2508 = ((~g1044))|((~I2506));
assign I2324 = ((~g1209));
assign g5047 = (g3954&g4806);
assign g4777 = ((~g4457)&(~g4459));
assign I8500 = ((~g6431));
assign I2825 = ((~g1143));
assign I3340 = ((~g1282));
assign I6819 = ((~g5019));
assign g6654 = ((~I8758));
assign I8997 = ((~g6790));
assign g4249 = ((~I5699));
assign g3991 = (g3685)|(g3156);
assign g3465 = ((~g2986));
assign g2030 = ((~I3137));
assign g4637 = (g4344)|(g3619);
assign g5916 = (g5728)|(g3781);
assign g2025 = ((~g1276));
assign g2265 = ((~I3408));
assign g1887 = ((~I2982));
assign g4285 = (g3490)|(g3887);
assign I2961 = ((~g1731));
assign I7002 = ((~g5308));
assign g5274 = ((~I6933));
assign I5648 = ((~g3974))|((~I5647));
assign g2796 = ((~I3999));
assign g5536 = ((~g5467));
assign I6963 = ((~g4874))|((~I6962));
assign I5400 = ((~g3963));
assign g5159 = (g536&g4967);
assign g5210 = ((~I6874));
assign I5644 = ((~g4059));
assign I3699 = ((~g642))|((~I3697));
assign g3053 = ((~I4276));
assign g4468 = (g4214)|(g3831);
assign g1960 = ((~I3071));
assign I7197 = ((~g5431));
assign I2880 = ((~g1143));
assign g1637 = ((~I2596));
assign g3571 = ((~g3084));
assign g5142 = (g148&g5099);
assign g4803 = ((~I6474))|((~I6475));
assign g6416 = ((~I8258));
assign g3094 = ((~I4337));
assign g3463 = ((~g2682));
assign g6239 = (g2339)|(g6073);
assign g4333 = (g3964&g3284);
assign g4508 = ((~I6036));
assign I5768 = ((~g3957))|((~I5766));
assign I3071 = ((~g1504));
assign g4812 = ((~g4550))|((~g1560))|((~g1559))|((~g2073));
assign I3740 = ((~g2021))|((~I3739));
assign g1219 = ((~I2218));
assign g3377 = (g3118&g2931);
assign I5442 = ((~g3731));
assign I6143 = ((~g4237));
assign I3328 = ((~g1273));
assign I4252 = ((~g2555));
assign g1043 = ((~g486));
assign g6176 = (g6068)|(g6033);
assign g6909 = (g6896&g6894);
assign I7313 = ((~g590))|((~I7311));
assign I2290 = ((~g971));
assign I6475 = ((~g578))|((~I6473));
assign I3954 = ((~g2497))|((~I3952));
assign g3772 = ((~g3466));
assign g4267 = ((~I5720));
assign I5865 = ((~g3743));
assign g2419 = (g1808&g54);
assign g3144 = (g236&g2440);
assign I2134 = ((~g705));
assign g3651 = (g3064&g2766);
assign I2013 = ((~g532))|((~g260));
assign g1899 = ((~I2998));
assign g6884 = ((~I9119));
assign g2712 = ((~g2320));
assign I8476 = ((~g6457));
assign I2143 = ((~g2));
assign g1641 = ((~I2604));
assign g3779 = ((~g3466));
assign g3329 = (g2748&g2907);
assign g1703 = ((~I2707));
assign I2221 = ((~g43));
assign I4623 = ((~g2962));
assign g4628 = ((~g4273));
assign g4566 = ((~g4198));
assign I8730 = ((~g6535));
assign g4698 = (g4586&g2106);
assign g1319 = ((~I2312));
assign I7170 = ((~g5435));
assign g3834 = ((~I5027));
assign g1123 = ((~I2165));
assign I8273 = ((~g6301));
assign g4732 = ((~I6362));
assign I7871 = ((~g6097));
assign I2399 = ((~g729));
assign I2199 = ((~g33));
assign g6327 = (g3884&g6212);
assign g5894 = ((~g5731));
assign g5601 = (g5052&g5518);
assign I5837 = ((~g3850));
assign g2719 = ((~I3875))|((~I3876));
assign I8809 = ((~g6687));
assign I6391 = ((~g4504))|((~I6390));
assign g3697 = (g2796&g2481);
assign g6434 = ((~I8300));
assign g4002 = ((~I5293))|((~I5294));
assign I5214 = ((~g3567));
assign g5527 = ((~I7267));
assign I2109 = ((~g602))|((~I2108));
assign g4661 = (g4637&g4634);
assign I5071 = ((~g3263));
assign I5209 = ((~g3271))|((~I5207));
assign I9098 = ((~g6864));
assign I8512 = ((~g6441));
assign g6252 = (g5905)|(g2381);
assign g4435 = ((~I5944));
assign g5948 = (g5779&g5407);
assign g4824 = ((~g4615));
assign g2864 = ((~g1887));
assign g2781 = (g2544&g1982);
assign g2961 = ((~g1861));
assign I8659 = ((~g6523));
assign g6569 = ((~I8591));
assign g4387 = ((~I5868));
assign g5624 = (g5494)|(g3280);
assign I7097 = ((~g5194))|((~g574));
assign I2334 = ((~g1193));
assign g2771 = (g2497&g1975);
assign I5019 = ((~g3318));
assign I5301 = ((~g471))|((~I5300));
assign g5054 = ((~g4816));
assign g3028 = ((~I4234))|((~I4235));
assign g6301 = (g6254)|(g6092);
assign g5996 = ((~g5824));
assign g5191 = (g461&g4877);
assign g1518 = ((~g980)&(~g965));
assign g5160 = ((~g5099));
assign I1947 = ((~g699));
assign g4900 = ((~I6607));
assign g4219 = (g3911&g1655);
assign g4790 = ((~I6456));
assign I8897 = ((~g6707));
assign g2766 = ((~g2361));
assign g3517 = ((~g3173))|((~g3002))|((~g2976))|((~g2179));
assign g1327 = ((~I2334));
assign g1334 = ((~I2355));
assign I2340 = ((~g1142));
assign g709 = ((~g114));
assign I3112 = ((~g1439));
assign g5454 = (g5256&g4549);
assign I8432 = ((~g6411));
assign g5177 = (g445&g4877);
assign g4170 = (g382&g3900);
assign g2253 = ((~I3388));
assign g3375 = (g260&g2912);
assign g2975 = ((~I4176));
assign g3082 = ((~I4315));
assign I6403 = ((~g4492));
assign I6063 = ((~g4381));
assign g3874 = ((~I5103));
assign I7521 = ((~g361))|((~I7520));
assign g2515 = ((~I3641));
assign I4809 = ((~g2974));
assign I8620 = ((~g6541));
assign g5676 = (g5559)|(g5424);
assign g6899 = ((~I9164));
assign I2349 = ((~g1160));
assign g4382 = ((~I5857));
assign I8650 = ((~g6529));
assign g2850 = (g2018&g1255);
assign I2601 = ((~g1161));
assign g5010 = ((~I6646));
assign I2663 = ((~g1006));
assign g1236 = ((~I2234));
assign g6767 = (g6754&g2986);
assign g6670 = (g6557)|(g6634)|(g4410)|(g2948);
assign I5068 = ((~g3571));
assign g6465 = ((~I8329));
assign g4225 = ((~g4059));
assign g4565 = ((~g4195));
assign g4188 = ((~I5594));
assign g4853 = ((~I6567));
assign g5251 = ((~g5069));
assign I6420 = ((~g4618));
assign g3661 = (g2234&g2778);
assign I3999 = ((~g1837));
assign g2588 = ((~I3717));
assign I6661 = ((~g3541))|((~I6659));
assign I3990 = ((~g2544))|((~I3988));
assign I2611 = ((~g1209));
assign g1583 = ((~g1001));
assign g6420 = ((~I8270));
assign g4678 = ((~g2897))|((~g2101))|((~g1514))|((~g4550));
assign g4222 = ((~I5654));
assign g5630 = (g5501)|(g3309);
assign g3631 = (g2631&g2324);
assign g3726 = (g119&g3251);
assign g2494 = ((~I3623));
assign I7478 = ((~g5628));
assign g3457 = ((~g2653));
assign I7254 = ((~g5458));
assign g4404 = ((~I5907));
assign g5687 = ((~g5567));
assign I6346 = ((~g4563));
assign g5582 = ((~I7342));
assign I7230 = ((~g170))|((~g5372));
assign g3829 = (g3294)|(g3305);
assign g850 = ((~g602));
assign g1046 = ((~g489));
assign I3031 = ((~g1504));
assign g4607 = (g4232)|(g3899);
assign g6260 = (g1703&g6048);
assign I3468 = ((~g1802));
assign g3871 = (g3701)|(g3186);
assign I8834 = ((~g6661));
assign g5554 = ((~g5455));
assign I4009 = ((~g292))|((~I4008));
assign I7570 = ((~g79))|((~I7569));
assign g6679 = (g6637)|(g6558);
assign g6456 = (g6346)|(g5954);
assign I8576 = ((~g6436));
assign g1575 = (g980&g965);
assign g3593 = ((~g2997));
assign g2440 = ((~I3575));
assign g3966 = ((~g3329)&(~g3339));
assign I8255 = ((~g6292));
assign g3177 = ((~I4414));
assign I8074 = ((~g6118));
assign I3540 = ((~g1670));
assign I6659 = ((~g4762))|((~g3541));
assign g2959 = ((~g1861));
assign g4873 = (g4838&g4173);
assign g6444 = (g6338)|(g5936);
assign I6579 = ((~g4798));
assign I8961 = ((~g6778));
assign g6376 = ((~g6267));
assign I4445 = ((~g2092))|((~I4444));
assign g4596 = ((~g4184)&(~g4186));
assign I8441 = ((~g6419));
assign g897 = ((~g41));
assign g4613 = ((~I6195))|((~I6196));
assign g6771 = (g6758&g3483);
assign I6362 = ((~g4569));
assign g3302 = (g212&g2867);
assign g5797 = ((~I7596));
assign I3641 = ((~g1491));
assign I3779 = ((~g2125));
assign g2091 = ((~g1355));
assign I7058 = ((~g5281));
assign g6429 = ((~g6376)&(~g4086)&(~g4074)&(~g4302));
assign g5085 = (g4694)|(g4280);
assign g1293 = ((~I2284));
assign g5515 = (g590&g5364);
assign I8727 = ((~g6536));
assign I7802 = ((~g5920));
assign g1160 = ((~I2179));
assign I2653 = ((~g996));
assign g6553 = ((~I8555));
assign g3986 = (g3667)|(g3133);
assign I3691 = ((~g1732));
assign g2343 = ((~I3493));
assign g4048 = (g414&g3388);
assign g5617 = (g5061&g5524);
assign g1880 = ((~g1603));
assign I3516 = ((~g1295));
assign g5435 = ((~I7113));
assign g3299 = ((~g3049));
assign I8180 = ((~g6176));
assign g6601 = ((~I8671));
assign g4840 = ((~I6528));
assign g4446 = (g4383)|(g4043);
assign g5486 = (g386&g5331);
assign g1116 = ((~I2154));
assign I5532 = ((~g3861));
assign I2943 = ((~g1715));
assign I8423 = ((~g6423));
assign g2647 = ((~I3791));
assign I8524 = ((~g6496));
assign I7972 = (g4915)|(g5025);
assign g3684 = (g2268&g2817);
assign I5382 = ((~g3952));
assign I8479 = ((~g6482));
assign g1684 = ((~I2668));
assign g945 = ((~g536));
assign g6937 = (g4616)|(g6934);
assign g1233 = ((~I2231));
assign g5358 = ((~I7012));
assign g1439 = ((~I2449));
assign g5138 = ((~I6792));
assign I7223 = ((~g161))|((~g5370));
assign g3118 = ((~I4366));
assign I2998 = ((~g1257));
assign g5242 = ((~g5085));
assign g4585 = ((~g4171)&(~g4177));
assign g862 = ((~g319));
assign g4180 = (g3929&g2119);
assign g1484 = ((~I2473));
assign I5760 = ((~g3836))|((~I5759));
assign I6417 = ((~g4617));
assign g3290 = (g2213&g2664);
assign I4123 = ((~g2043));
assign g4502 = ((~I6020));
assign g6308 = ((~I8034));
assign I9170 = ((~g6883));
assign g6044 = ((~g5824));
assign g2541 = ((~I3659));
assign I8913 = ((~g6743));
assign g3658 = (g3118&g2776);
assign g1998 = ((~I3109));
assign g3228 = ((~I4483));
assign g3903 = ((~g3505)&(~g471));
assign g3859 = ((~I5078));
assign g5864 = ((~g5649))|((~g1529))|((~g1088))|((~g2068));
assign g6616 = ((~I8710));
assign I7167 = ((~g5434));
assign g2906 = ((~g1911));
assign g1076 = ((~I2115));
assign g3671 = (g2760&g2405);
assign g2754 = ((~g2347));
assign I5686 = ((~g3942));
assign I1825 = ((~g361));
assign g3782 = ((~g3388));
assign I8860 = ((~g6699));
assign I2630 = ((~g1143));
assign I8079 = (g6194)|(g5958)|(g5975)|(g5997);
assign g3076 = ((~I4309));
assign I2428 = ((~g774));
assign I1874 = ((~g282));
assign I3816 = ((~g2580));
assign I3109 = ((~g1504));
assign g5395 = ((~I7061));
assign g5553 = (g5012&g5440);
assign g3535 = ((~g3216))|((~g2215))|((~g2197))|((~g2968));
assign I3927 = ((~g2245));
assign I8975 = ((~g6791));
assign I8165 = ((~g6189));
assign g5937 = (g5775&g5392);
assign g2720 = (g2422&g1919);
assign g5450 = ((~g5292));
assign g2243 = ((~I3376));
assign I7372 = ((~g5493));
assign g5492 = (g5441&g3452);
assign g3367 = (g2809&g1960);
assign g2608 = ((~I3746));
assign g6812 = ((~I8984));
assign I6549 = ((~g4699));
assign I4334 = ((~g2256));
assign g5310 = ((~g5067));
assign I7686 = ((~g5705));
assign g6102 = ((~I7802));
assign g4103 = ((~I5391));
assign g2179 = ((~I3328));
assign I4159 = ((~g2015))|((~g619));
assign g6402 = ((~I8220));
assign g6828 = (g6803&g5958);
assign g4723 = ((~I6349));
assign I4273 = ((~g2197));
assign I9119 = ((~g6855));
assign g4054 = (g3694&g69);
assign I2627 = ((~g1053));
assign I2721 = ((~g1219));
assign g1821 = ((~I2883));
assign I3575 = ((~g1305));
assign g2158 = ((~I3281));
assign g3600 = ((~I4791));
assign g6848 = (g3741&g328&g6843);
assign I6473 = ((~g4541))|((~g578));
assign g929 = ((~g49));
assign g1581 = ((~g910));
assign I9092 = ((~g6855));
assign g2104 = ((~g1372));
assign I8195 = ((~g471))|((~I8194));
assign g3195 = (g2473&g2541);
assign g6817 = ((~I8988));
assign g3840 = ((~I5043));
assign g4044 = (g410&g3388);
assign I7173 = ((~g5436));
assign g3480 = ((~g2986));
assign g6094 = (g1177&g5753);
assign g4451 = (g4390)|(g4048);
assign g5499 = (g5451&g3462);
assign I6733 = ((~g4773));
assign g3821 = (g2951)|(g3466);
assign g3923 = ((~g3378)&(~g3381));
assign I8656 = ((~g6532));
assign g6535 = ((~I8521));
assign g4213 = ((~I5633));
assign g6924 = (g6920&g6919);
assign I6956 = ((~g5124));
assign g3289 = ((~g3034));
assign g1842 = ((~g1612));
assign I5630 = ((~g3914));
assign g6070 = ((~g5824));
assign g3276 = ((~I4546))|((~I4547));
assign g4730 = (g1423&g4565);
assign g3459 = ((~g2664));
assign g3902 = ((~g3575));
assign g3291 = ((~g3037));
assign g1108 = ((~I2134));
assign g2631 = ((~I3773));
assign I7153 = ((~g5358));
assign g3972 = (g3646)|(g3103);
assign I5328 = ((~g3502));
assign g1820 = ((~I2880));
assign g894 = ((~I1917));
assign g2800 = ((~g2430));
assign g4137 = ((~I5493));
assign g4494 = ((~I6004));
assign g3743 = (g3344)|(g2758);
assign I3313 = ((~g1337));
assign g6541 = ((~I8535));
assign g3611 = (g2370&g3037);
assign g6135 = (g5584&g5958);
assign g6543 = ((~I8541));
assign I7267 = ((~g5458));
assign g1711 = ((~I2712));
assign g5303 = (g5053)|(g4768);
assign I5309 = ((~g3512))|((~I5307));
assign I8203 = ((~g6192))|((~I8201));
assign g1891 = ((~I2986));
assign g4611 = (g3985&g119&g4300);
assign g3490 = (g353&g2959);
assign I5385 = ((~g3962));
assign g5693 = (g5632)|(g5481);
assign g4155 = ((~I5551));
assign g2568 = ((~I3678));
assign g3886 = ((~g3346));
assign g849 = ((~g598));
assign I6933 = ((~g5124));
assign g2891 = ((~g1884));
assign g4156 = (g3926&g2078);
assign I8309 = ((~g6304));
assign I6340 = ((~g4561));
assign g4356 = (g175&g3779);
assign I3528 = ((~g1422));
assign I3833 = ((~g2266));
assign g3379 = (g3104&g1988);
assign g6427 = ((~g6376)&(~g4086)&(~g4074)&(~g4068));
assign I6072 = ((~g4385));
assign I3569 = ((~g1789));
assign g1498 = ((~I2479));
assign I7548 = ((~g64))|((~g5672));
assign g6248 = (g465&g5894);
assign g2607 = ((~I3740))|((~I3741));
assign g4307 = ((~I5774));
assign I5622 = ((~g3914));
assign g6500 = ((~I8420));
assign g4343 = ((~g4011));
assign g5250 = ((~g4929));
assign g6697 = ((~I8809));
assign I2542 = ((~g821))|((~g774));
assign I2408 = ((~g719));
assign g5875 = ((~I7637));
assign g3833 = (g3602)|(g3608);
assign g5777 = ((~I7535))|((~I7536));
assign g4657 = ((~I6244));
assign g2663 = ((~g2308));
assign I6995 = ((~g5220));
assign g749 = ((~I1847));
assign g6896 = ((~I9155));
assign I5177 = ((~g3267));
assign I8573 = ((~g6435));
assign I3629 = ((~g1759));
assign g5682 = (g84&g5578);
assign g6271 = (g2955)|(g5885);
assign I3965 = ((~g2268));
assign g4395 = (g445&g3800);
assign I2620 = ((~g1177));
assign I6615 = ((~g4745));
assign I5109 = ((~g3710));
assign g3685 = (g2256&g2818);
assign g2213 = ((~I3346));
assign g4134 = ((~I5484));
assign g6614 = (g932&g6556);
assign I3614 = ((~g1295));
assign g5087 = ((~g4736));
assign g3343 = ((~g3090));
assign I8150 = ((~g6185));
assign I3419 = ((~g1287));
assign I4347 = ((~g2555));
assign g1052 = ((~g668));
assign g5446 = (g4537&g5241);
assign g5351 = (g5326&g3459);
assign g6309 = (g6265)|(g6098);
assign I9185 = ((~g6877));
assign g5049 = ((~I6685));
assign I5705 = ((~g3942));
assign g2858 = ((~g1815))|((~g2577));
assign g1059 = ((~g702));
assign g1720 = ((~g1111));
assign g760 = ((~I1853));
assign I5264 = ((~g3638));
assign g3984 = ((~g3564));
assign I5654 = ((~g3742));
assign g4057 = (g422&g3388);
assign g1833 = ((~I2913));
assign g4115 = ((~I5427));
assign g1696 = ((~I2700));
assign g3332 = ((~g3079));
assign g5477 = ((~I7167));
assign g3095 = ((~I4340));
assign I2391 = ((~g774));
assign I7576 = ((~g84))|((~g5680));
assign g5062 = (g4661)|(g4666);
assign g3437 = (g837&g2853);
assign g4460 = (g4218&g1539);
assign g6268 = (g5677)|(g5951);
assign I2683 = ((~g613))|((~I2681));
assign g5936 = (g5113&g5788);
assign I8147 = ((~g6182));
assign g1594 = ((~g1143));
assign I4205 = ((~g743))|((~I4203));
assign I4223 = ((~g2176));
assign g5149 = (g4910&g1480);
assign g2059 = ((~g1402));
assign g4160 = (g3923&g1345);
assign I6170 = ((~g4343));
assign g5540 = ((~I7284));
assign g5888 = ((~g5731));
assign I2067 = ((~g686));
assign g3911 = ((~I5148));
assign g4932 = (g157&g4727);
assign g3760 = (g548&g3465);
assign I2014 = ((~g532))|((~I2013));
assign g4321 = ((~I5790));
assign g6770 = (g6754&g3482);
assign I4288 = ((~g2215));
assign I6706 = ((~g4731));
assign g1772 = ((~I2811));
assign I4195 = ((~g2173));
assign g5277 = (g5023)|(g4763);
assign I6444 = ((~g4503));
assign g1762 = ((~I2791));
assign g3767 = (g2706&g3504);
assign I3471 = ((~g1450));
assign I3013 = ((~g1519));
assign I7562 = ((~g74))|((~g5676));
assign g6748 = (g6733&g6732);
assign g6125 = (g5708&g5975);
assign g2701 = ((~I3855));
assign I7587 = ((~g5605));
assign I7336 = ((~g5534));
assign g2839 = ((~g2535));
assign g4179 = (g390&g3902);
assign g5197 = (g465&g4967);
assign g5217 = (g4866&g5092);
assign g3180 = (g260&g2506);
assign I3395 = ((~g1286));
assign g2357 = ((~I3509));
assign g2136 = ((~g1395));
assign g6373 = ((~I8183));
assign g2111 = ((~g1384));
assign g5326 = (g5069)|(g4410)|(g3012);
assign g2015 = (g616&g1419);
assign g6690 = (g6270)|(g6650);
assign g4218 = ((~I5640));
assign g4374 = ((~I5837));
assign I4031 = ((~g1846));
assign g4601 = ((~g4191));
assign g3792 = ((~g3388));
assign g3383 = (g3128&g2004);
assign I5784 = ((~g628))|((~I5782));
assign I7796 = ((~g5917));
assign g4703 = ((~I6299));
assign I3047 = ((~g1426));
assign g6512 = ((~I8456));
assign g5451 = (g5251&g4544);
assign I8888 = ((~g6708));
assign g6738 = (g6713&g809&g5242);
assign g5379 = ((~I7035));
assign g4778 = ((~I6430));
assign I7081 = ((~g5281));
assign g6066 = (g5824&g1721);
assign I3596 = ((~g1305));
assign g5372 = (g5213)|(g4942);
assign g4669 = ((~g4550))|((~g1017))|((~g1680))|((~g2897));
assign g1220 = ((~I2221));
assign I2676 = ((~g131))|((~I2674));
assign g4247 = (g1764&g4007&g1628);
assign g6334 = (g3858&g6212);
assign g4865 = (g4776&g1849);
assign g3901 = ((~g3575));
assign I2358 = ((~g1176));
assign g3963 = ((~I5217));
assign g6588 = ((~I8632));
assign g2079 = ((~g1348));
assign g1848 = ((~I2946));
assign g2585 = ((~I3708));
assign g3327 = (g2772&g2906);
assign I7698 = ((~g5717));
assign g3883 = (g3709)|(g3203);
assign g2053 = (g1094&g1675);
assign g4221 = ((~I5648))|((~I5649));
assign g3683 = (g3150&g2813);
assign g1620 = (g1056&g1084);
assign g1609 = (g760&g754);
assign g6524 = ((~I8488));
assign g1555 = ((~I2521));
assign g6744 = ((~I8910));
assign g2550 = ((~I3665));
assign g6941 = ((~I9236));
assign g6077 = (g5824&g1735);
assign I2898 = ((~g1027))|((~I2897));
assign g4716 = ((~I6330));
assign g4248 = ((~I5696));
assign g6363 = ((~I8153));
assign g3649 = (g3104&g2764);
assign g3127 = (g224&g2394);
assign g5660 = (g4509&g5549);
assign I8638 = ((~g6553));
assign g5387 = ((~I7051));
assign g6685 = (g6256)|(g6644);
assign I3669 = ((~g1739));
assign I8665 = ((~g6527));
assign I6561 = ((~g4707));
assign g2306 = ((~g1743));
assign g710 = ((~g128));
assign I2072 = ((~g15))|((~g11));
assign g4527 = ((~I6093));
assign g6035 = ((~g5824));
assign I2877 = ((~g1123));
assign I7104 = ((~g5273));
assign I2893 = ((~g1236));
assign g4145 = ((~I5517));
assign g3891 = (g3683)|(g3688);
assign g5231 = (g5048)|(g672);
assign I2682 = ((~g918))|((~I2681));
assign I5081 = ((~g3589));
assign g2672 = ((~I3816));
assign g2134 = ((~I3258));
assign g4708 = (g578&g4541);
assign g5186 = (g422&g4950);
assign g4309 = ((~g4074));
assign I8818 = ((~g6690));
assign g2509 = ((~I3635));
assign I8857 = ((~g6698));
assign g5995 = ((~g5824));
assign g5782 = ((~I7570))|((~I7571));
assign g6493 = ((~g6375));
assign g4126 = ((~I5460));
assign g1690 = ((~I2692));
assign I9233 = ((~g6938));
assign g1854 = ((~I2958));
assign g3203 = (g2497&g2565);
assign I3934 = ((~g288))|((~I3933));
assign g1988 = ((~I3099));
assign g4237 = ((~g4049))|((~g4017));
assign I5484 = ((~g3875));
assign g2726 = ((~I3886));
assign I8707 = ((~g6520));
assign g2675 = ((~I3819));
assign g1111 = ((~I2143));
assign I2617 = ((~g1193));
assign g2252 = ((~I3385));
assign g4667 = (g4653&g4651);
assign g5943 = ((~g5818))|((~g2940));
assign g3626 = (g3031&g2727);
assign g6310 = (g6269)|(g6099);
assign I8420 = ((~g6422));
assign I6114 = ((~g4405));
assign I4939 = ((~g3437))|((~g357));
assign g3930 = ((~g3317)&(~g3328));
assign I6534 = ((~g4706));
assign g6530 = ((~I8506));
assign g1797 = ((~g98))|((~g1064))|((~g1070));
assign g1398 = ((~g306))|((~g889));
assign g5069 = (g1595)|(g4688);
assign g6507 = ((~I8441));
assign I2498 = ((~g1042))|((~I2497));
assign g4226 = ((~g4050));
assign I9208 = ((~g6922));
assign g5330 = ((~I6992));
assign I5882 = ((~g3871));
assign g6156 = (g2591&g6015);
assign g6141 = (g3173&g5997);
assign I8379 = (g5212)|(g6357);
assign g2043 = ((~I3158));
assign I4935 = ((~g3369));
assign g6236 = ((~g6070));
assign I9038 = ((~g6833));
assign I5548 = ((~g4059));
assign g1459 = ((~g926)&(~g950)&(~g948));
assign I8159 = ((~g6167));
assign I8411 = ((~g6415));
assign g6322 = ((~I8056));
assign I7556 = ((~g69))|((~I7555));
assign g4597 = (g3694&g4286);
assign g1642 = ((~g809));
assign g1274 = ((~g856));
assign g2882 = ((~g1854));
assign I8044 = ((~g6252));
assign g3704 = (g2276&g2841);
assign g1335 = ((~I2358));
assign I2537 = ((~g971));
assign I2675 = ((~g710))|((~I2674));
assign g4047 = (g453&g3388);
assign g3238 = ((~I4513));
assign I6685 = ((~g4716));
assign g5234 = (g197&g4915);
assign g2370 = ((~I3522));
assign g5863 = ((~g5649))|((~g1076))|((~g1535))|((~g2068));
assign g2554 = ((~I3669));
assign g6417 = ((~I8261));
assign g6698 = ((~I8812));
assign g5924 = ((~I7704));
assign g3326 = (g2734&g1891);
assign I5659 = ((~g3979))|((~I5657));
assign I5252 = ((~g3546));
assign I8541 = ((~g6452));
assign g3376 = (g3104&g1979);
assign I6187 = ((~g3955))|((~I6185));
assign I3083 = ((~g1426));
assign g1122 = ((~I2162));
assign I2053 = ((~g684));
assign g4457 = (g4261&g2902);
assign I5952 = ((~g4367));
assign g6144 = (g3183&g5997);
assign I9101 = ((~g6855));
assign g5574 = ((~g5407));
assign g6669 = (g6613)|(g4679);
assign g2953 = (g2381&g293);
assign g1519 = ((~I2491));
assign I8177 = ((~g6173));
assign I8544 = ((~g6453));
assign g1283 = ((~g853));
assign I3653 = ((~g1305));
assign I3617 = ((~g1305));
assign g5202 = (g4904)|(g4914)|(g4894);
assign g2042 = ((~I3155));
assign g2295 = ((~g1578));
assign g3921 = ((~g3512));
assign g6799 = (g4948&g6782);
assign g1593 = ((~g1054));
assign g6435 = ((~g6376)&(~g4086)&(~g4309)&(~g4302));
assign I8246 = ((~g6290));
assign I7583 = ((~g5605));
assign I5208 = ((~g3267))|((~I5207));
assign I6299 = ((~g4438));
assign I2916 = ((~g1643));
assign g1117 = ((~g32));
assign g6572 = ((~I8600));
assign g1318 = ((~I2309));
assign I3647 = ((~g1747));
assign g1655 = ((~g985));
assign g5485 = (g382&g5331);
assign g1759 = ((~I2782));
assign g6492 = ((~g6348)&(~g1734));
assign I8582 = ((~g6439));
assign g2212 = ((~I3343));
assign g5048 = ((~g4819)&(~g3491)&(~g3559));
assign g6048 = ((~g5824));
assign g5531 = (g5349)|(g3275);
assign I2785 = ((~g1222));
assign g4670 = ((~g4611))|((~g3528));
assign g4513 = ((~I6051));
assign I8290 = ((~g6291));
assign I1995 = ((~g504))|((~I1994));
assign I5692 = ((~g3942));
assign g6883 = ((~I9116));
assign I8916 = ((~g6742));
assign g6302 = (g5740&g6164);
assign g4388 = ((~I5871));
assign g6706 = ((~I8828));
assign g4660 = ((~I6253));
assign g6803 = ((~I8975));
assign I3952 = ((~g289))|((~g2497));
assign g5524 = ((~I7264));
assign I4516 = ((~g2777));
assign g6511 = ((~I8453));
assign I6126 = ((~g4240));
assign I5249 = ((~g3589));
assign g1654 = ((~g878));
assign g2625 = ((~I3767));
assign I3843 = ((~g2145));
assign g5178 = (g516&g4993);
assign I7646 = ((~g5774));
assign I3093 = ((~g1426));
assign g6655 = ((~I8761));
assign I7091 = ((~g5281));
assign g4206 = ((~I5626));
assign g3858 = (g3629)|(g3636);
assign g6710 = ((~I8840));
assign g6754 = (g6676)|(g6625)|(g6737);
assign I3074 = ((~g1426));
assign I6775 = ((~g4790));
assign g4842 = ((~I6534));
assign I5481 = ((~g3866));
assign g6117 = ((~g5880));
assign I5647 = ((~g3974))|((~g3968));
assign I9137 = ((~g6864));
assign g1426 = ((~I2445));
assign g5166 = (g541&g4967);
assign g4161 = (g3931&g2087);
assign g2024 = ((~I3126))|((~I3127));
assign g5228 = (g5096)|(g4800);
assign g6660 = (g6640)|(g6637);
assign I6962 = ((~g4874))|((~g586));
assign g4636 = ((~g4286));
assign g2740 = ((~I3909));
assign I3502 = ((~g1295));
assign g2734 = ((~I3902));
assign g899 = ((~I1924));
assign g6747 = (g6614)|(g6731);
assign g1664 = ((~I2643));
assign g5537 = ((~g5385));
assign I3441 = ((~g1502));
assign g2066 = ((~g1341));
assign g5821 = ((~g5638))|((~g2056))|((~g1076))|((~g1666));
assign g6421 = ((~I8273));
assign g5143 = (g157&g5099);
assign g6930 = (g6740)|(g6928);
assign g5211 = (g4860&g5086);
assign g6314 = ((~I8044));
assign g3052 = ((~I4273));
assign g950 = ((~I2022))|((~I2023));
assign I3158 = ((~g1829));
assign g6368 = ((~I8168));
assign g5120 = ((~I6772));
assign g3192 = ((~I4429));
assign I6102 = ((~g4399));
assign I7535 = ((~g54))|((~I7534));
assign I5403 = ((~g3970));
assign g1769 = ((~I2802));
assign I6099 = ((~g4398));
assign g4948 = (g4834)|(g4836);
assign g4764 = ((~I6400));
assign g4559 = ((~g4187));
assign g830 = ((~g338));
assign I8467 = ((~g6457));
assign g6085 = (g1161&g5731);
assign g6720 = ((~I8854));
assign I2122 = ((~g689));
assign I8881 = ((~g6711));
assign I6084 = ((~g4391));
assign I2207 = ((~g7));
assign g719 = ((~I1835));
assign g4805 = ((~g4473));
assign g5436 = ((~I7116));
assign I3361 = ((~g1331));
assign g6130 = (g5720&g5958);
assign g4503 = ((~I6023));
assign g3223 = ((~I4468));
assign g6554 = (g6337)|(g6466);
assign I7342 = ((~g5579));
assign g1161 = ((~I2182));
assign I8279 = ((~g6307));
assign g3672 = (g3136&g2800);
assign g5245 = (g297&g4915);
assign I4444 = ((~g2092))|((~g606));
assign g3650 = (g2660&g2347);
assign g6450 = (g6341)|(g5940);
assign I6414 = ((~g4497));
assign g6841 = ((~I9044));
assign g1702 = ((~g1107));
assign g5218 = (g564&g5025);
assign g3616 = (g2397&g3049);
assign g6915 = (g6906&g6905);
assign g3301 = (g218&g2866);
assign g4769 = ((~g4606));
assign g4035 = (g437&g3388);
assign I9021 = ((~g6812));
assign g5804 = (g5371)|(g5603);
assign g6617 = ((~I8713));
assign g1292 = ((~I2281));
assign I5520 = ((~g3835));
assign g5787 = ((~g5685));
assign I6105 = ((~g4400));
assign g2936 = ((~g2026));
assign g3054 = ((~I4279));
assign I6231 = ((~g4350));
assign g6167 = (g6056)|(g6039);
assign I5412 = ((~g4034));
assign I7549 = ((~g64))|((~I7548));
assign g3985 = ((~g1138))|((~g3718))|((~g2142));
assign g2933 = ((~I4123));
assign g3176 = (g2422&g2494);
assign g3161 = (g2397&g2470);
assign g898 = ((~g47));
assign g6173 = (g6066)|(g6043);
assign I2883 = ((~g1143));
assign g4189 = ((~I5597));
assign g1683 = ((~g1017));
assign g948 = ((~I2014))|((~I2015));
assign g6736 = (g6712&g754&g5237);
assign g4181 = (g3939&g1381);
assign g834 = ((~g341));
assign g4240 = ((~g1589)&(~g1879)&(~g3793));
assign g3229 = ((~I4486));
assign g5883 = (g5824&g3752);
assign g6701 = ((~I8821));
assign g939 = ((~I1987))|((~I1988));
assign g4662 = ((~g4640));
assign g2907 = ((~g1914));
assign g2875 = ((~g1940));
assign g6255 = (g1335&g5895);
assign g861 = ((~g179));
assign g6792 = (g6770)|(g3321);
assign g6600 = ((~I8668));
assign g4798 = ((~I6464));
assign I7971 = (g5202)|(g4993)|(g4967)|(g4980);
assign I5116 = ((~g3259));
assign g5170 = (g5091&g2111);
assign g4800 = (g4648&g4296);
assign I7073 = ((~g5281));
assign g6768 = (g6750&g3477);
assign g4789 = (g3551&g4632);
assign I6816 = ((~g5111));
assign g5053 = (g4599&g4808);
assign g5854 = ((~g5638))|((~g1683))|((~g1552))|((~g2062));
assign g2174 = ((~I3313));
assign g1411 = ((~g314))|((~g873));
assign g3499 = (g357&g2961);
assign I3346 = ((~g1327));
assign g2819 = ((~g2467));
assign g3729 = (g327&g3441);
assign I7224 = ((~g161))|((~I7223));
assign g4436 = (g4359)|(g4035);
assign g4509 = ((~I6039));
assign g3601 = ((~I4794));
assign g5623 = (g5503)|(g5357);
assign I2835 = ((~g1209));
assign g3845 = ((~I5050));
assign g2656 = ((~I3800));
assign I3776 = ((~g2044));
assign g2137 = (g760&g1638);
assign g6838 = ((~I9035));
assign g5562 = (g5228&g5457);
assign I6525 = ((~g4770));
assign g3992 = (g1555)|(g3559);
assign I6033 = ((~g4179));
assign g3374 = (g2809&g1969);
assign g1001 = ((~I2044));
assign g4403 = ((~I5904));
assign I4229 = ((~g2284));
assign I4267 = ((~g2525));
assign g5209 = (g560&g5025);
assign g4443 = (g4377)|(g4041);
assign g1282 = ((~g849));
assign I3697 = ((~g1570))|((~g642));
assign g3315 = (g2701&g1875);
assign g1729 = ((~I2731));
assign g3629 = (g2809&g2738);
assign I7065 = ((~g5281));
assign g6162 = ((~g5926));
assign g1852 = ((~I2952));
assign g1402 = ((~g310))|((~g866))|((~g873));
assign I6008 = ((~g4163));
assign g4429 = (g923&g4253&g2936);
assign g6604 = ((~I8678));
assign I8030 = ((~g6239));
assign I4940 = ((~g3437))|((~I4939));
assign g3453 = ((~g2628));
assign I7098 = ((~g5194))|((~I7097));
assign I5938 = ((~g4351));
assign I5236 = ((~g3545));
assign g3873 = (g3649)|(g3657);
assign I8894 = ((~g6709));
assign I7683 = ((~g5702));
assign g1546 = ((~g1101));
assign I2989 = ((~g1519));
assign g4804 = ((~g4473));
assign g3089 = (g212&g2336);
assign g2164 = ((~I3291));
assign g5281 = (g5074)|(g5124);
assign I3222 = ((~g1790));
assign I5316 = ((~g3557));
assign g1574 = ((~I2543))|((~I2544));
assign g6622 = ((~I8724));
assign g4545 = ((~g4416));
assign I4240 = ((~g2165));
assign g6109 = (g5900)|(g5599);
assign g1573 = ((~g729))|((~g719))|((~g766));
assign I3493 = ((~g1461));
assign g2125 = ((~I3255));
assign I2791 = ((~g1236));
assign g4472 = ((~g3380))|((~g4253));
assign g6628 = (g2138&g1612&g6540);
assign g6319 = ((~I8051));
assign I3788 = ((~g2554));
assign g4564 = ((~g4192));
assign g5424 = (g390&g5296);
assign I5668 = ((~g3828));
assign I2958 = ((~g1257));
assign g6739 = (g6715&g815&g5242);
assign g5433 = ((~I7107));
assign g1191 = ((~g38));
assign I3893 = ((~g286))|((~g2422));
assign g4328 = ((~g4092));
assign g4606 = ((~g4193));
assign I6054 = ((~g4194));
assign g5406 = (g374&g5270);
assign g3854 = ((~I5071));
assign g3828 = (g3304)|(g1351);
assign g3669 = (g2234&g2790);
assign g5429 = (g398&g5304);
assign I1938 = ((~g332));
assign I6321 = ((~g4559));
assign g3288 = (g2631&g2634);
assign g5583 = (g5569)|(g4020);
assign g3143 = (g242&g2437);
assign g1045 = ((~g699));
assign I8417 = ((~g6420));
assign I3741 = ((~g349))|((~I3739));
assign g1584 = ((~g743));
assign g3458 = ((~g2656));
assign g4053 = (g3387&g1415);
assign I4366 = ((~g2244));
assign g3773 = ((~g3466));
assign g3660 = (g2568&g3110);
assign g2682 = ((~I3826));
assign I2004 = ((~g500))|((~I2003));
assign g3884 = (g3666)|(g3671);
assign g6940 = ((~I9233));
assign I5594 = ((~g3821));
assign g6099 = (g1222&g5753);
assign I6452 = ((~g4629));
assign g6362 = ((~I8150));
assign g5051 = ((~I6689));
assign I5189 = ((~g3593))|((~I5187));
assign g5183 = (g418&g4950);
assign g4712 = ((~I6318));
assign g4715 = ((~I6327));
assign I5609 = ((~g3893));
assign g4758 = ((~I6382));
assign g3757 = (g2619&g3487);
assign g6140 = (g5587&g5975);
assign g1978 = ((~g1387));
assign g6568 = ((~I8588));
assign I5782 = ((~g3810))|((~g628));
assign I4784 = ((~g622))|((~I4782));
assign I2473 = ((~g971));
assign g2586 = ((~I3711));
assign g6529 = ((~I8503));
assign g3529 = ((~g3200))|((~g2215))|((~g2976))|((~g2968));
assign g2705 = ((~I3858));
assign g3718 = (g1743&g3140&g1157);
assign g5992 = ((~g5869));
assign g4363 = (g402&g3786);
assign g6157 = (g3158&g5997);
assign I5084 = ((~g3593));
assign g6335 = ((~I8079)&(~I8080)&(~I8081)&(~I8082));
assign I6630 = ((~g4745));
assign I1969 = ((~g516))|((~g236));
assign I6649 = ((~g4693));
assign g928 = ((~I1962))|((~I1963));
assign I3874 = ((~g285))|((~g2397));
assign g2671 = (g2263&g2296);
assign g6454 = (g6344)|(g5949);
assign g6294 = (g6249)|(g6090);
assign g6250 = (g1692&g6036);
assign g4129 = ((~I5469));
assign g2551 = (g715&g1826);
assign g3084 = ((~I4321));
assign I6531 = ((~g4704));
assign g4116 = ((~I5430));
assign I7543 = ((~g5669))|((~I7541));
assign g2923 = ((~g1969));
assign g5068 = (g4673)|(g4677);
assign g1556 = ((~g878));
assign g6431 = ((~I8295));
assign g6849 = ((~I9074));
assign g5752 = ((~I7509));
assign g3090 = ((~I4331));
assign g6300 = (g6253)|(g6091);
assign g6745 = ((~I8913));
assign g4658 = ((~I6247));
assign I2373 = ((~g1143));
assign g2577 = (g1743&g1797&g1793&g1138);
assign g5994 = ((~g5873));
assign g5151 = ((~I6819));
assign I2405 = ((~g1112));
assign g2524 = ((~I3647));
assign I8138 = (g4980)|(g4915)|(g5025)|(g5054);
assign I9082 = ((~g6849));
assign I2811 = ((~g1209));
assign g3933 = ((~g3327)&(~g3336));
assign g3728 = (g326&g3441);
assign g4786 = ((~I6448));
assign I7550 = ((~g5672))|((~I7548));
assign g4238 = ((~g3755)&(~g3279));
assign I1871 = ((~g281));
assign I1924 = ((~g663));
assign I6567 = ((~g4715));
assign g3357 = (g242&g2889);
assign g1743 = ((~g1064))|((~g94));
assign g2089 = (g1123&g1578);
assign I1856 = ((~g204));
assign g4173 = ((~I5577));
assign I2172 = ((~g691));
assign g5696 = (g5637)|(g5484);
assign g6558 = (g1842&g6474);
assign g1774 = ((~I2817));
assign g5376 = (g170&g5255);
assign g5443 = (g4537&g5251&g2307);
assign I4964 = ((~g3673));
assign I2922 = ((~g1774));
assign I2062 = ((~g3))|((~I2060));
assign I4402 = ((~g2283));
assign I2899 = ((~g634))|((~I2897));
assign g3075 = ((~I4306));
assign I3935 = ((~g2473))|((~I3933));
assign g6731 = (g6717&g4427);
assign I8235 = ((~g6312));
assign g1831 = ((~I2907));
assign g6406 = ((~I8232));
assign g5147 = ((~I6809));
assign g6298 = (g6255)|(g6093);
assign I6976 = ((~g5136));
assign g6864 = (g6852)|(g2089);
assign g5552 = ((~g5354)&(~g5356));
assign g3680 = (g2245&g2805);
assign I7707 = ((~g5701));
assign I4315 = ((~g2245));
assign g1249 = ((~I2240));
assign g3354 = ((~g3096));
assign g6534 = ((~I8518));
assign g2769 = ((~I3953))|((~I3954));
assign g5230 = ((~I6895));
assign g2744 = ((~g2336));
assign I3099 = ((~g1519));
assign g2913 = ((~g1925));
assign I7209 = ((~g143))|((~I7208));
assign g4583 = (g1808&g4267);
assign I6582 = ((~g4765));
assign I6182 = ((~g4249));
assign g6589 = ((~I8635));
assign g4772 = ((~I6420));
assign I5790 = ((~g3803));
assign g5949 = (g5119&g5805);
assign g1529 = ((~g1076));
assign I8535 = ((~g6447));
assign I5436 = ((~g3729));
assign g4631 = (g4340)|(g3611);
assign I6809 = ((~g5051));
assign g1481 = ((~g815)&(~g809));
assign g4722 = ((~I6346));
assign g5668 = (g49&g5571);
assign g4967 = ((~g4674)&(~g952));
assign g3541 = ((~g2643));
assign I2074 = ((~g11))|((~I2072));
assign g3019 = ((~I4226));
assign g1595 = (g729&g719&g766&I2566);
assign g3820 = (g3287)|(g2671);
assign I8755 = ((~g6561));
assign g6593 = ((~I8647));
assign I4802 = ((~g2877));
assign g2230 = ((~I3355));
assign g1721 = ((~I2721));
assign g5476 = ((~I7164));
assign g4246 = ((~I5692));
assign g6230 = ((~g6040));
assign g6259 = (g1699&g6044);
assign g2835 = ((~g2506));
assign g5955 = (g5782&g5420);
assign I4919 = ((~g3522))|((~g650));
assign g6340 = (g6257&g6069);
assign g3690 = (g2276&g2827);
assign g3286 = (g2196&g2656);
assign I7261 = ((~g5458));
assign I8681 = ((~g6566));
assign g5791 = ((~I7590));
assign g2692 = ((~I3840));
assign I3906 = ((~g2234));
assign I8552 = ((~g6455));
assign g5563 = ((~g5381));
assign I2749 = ((~g1209));
assign g6374 = ((~I8186));
assign g4608 = ((~I6176))|((~I6177));
assign I1978 = ((~g512))|((~g230));
assign g5632 = (g4494&g5538);
assign g4560 = ((~g4188));
assign g3209 = ((~I4452));
assign I8093 = ((~g6122));
assign I8360 = (I8356)|(I8357)|(I8358)|(I8359);
assign I6740 = ((~g4781));
assign g6902 = ((~I9173));
assign g1845 = ((~I2934))|((~I2935));
assign g1710 = ((~g1109));
assign g6263 = (g1711&g6052);
assign g4109 = ((~I5409));
assign g4394 = ((~I5885));
assign g996 = ((~I2041));
assign I5308 = ((~g478))|((~I5307));
assign g5681 = (g79&g5577);
assign g3785 = ((~g3466));
assign I9164 = ((~g6885));
assign g1514 = (g1017&g1011);
assign g4933 = ((~I6625));
assign g3275 = (g2172&g2615);
assign g6684 = (g6250)|(g6643);
assign I5451 = ((~g3967));
assign I2979 = ((~g1263));
assign g1826 = (g714&g710);
assign g4292 = ((~g4059));
assign g3928 = (g3512&g478);
assign I7577 = ((~g84))|((~I7576));
assign I2910 = ((~g1645));
assign g6351 = ((~I8107));
assign g2865 = ((~g2296));
assign g3612 = ((~I4809));
assign g4135 = ((~I5487));
assign g5449 = (g4545&g5246);
assign I4324 = ((~g1918));
assign g3320 = ((~g3067));
assign g1359 = ((~g866))|((~g306));
assign I4258 = ((~g2169));
assign g6074 = ((~g5794));
assign I2681 = ((~g918))|((~g613));
assign g1267 = ((~g843));
assign I3206 = ((~g1823));
assign I5948 = ((~g4360));
assign I2244 = ((~g567))|((~g598));
assign g3862 = (g3632)|(g3641);
assign g3364 = ((~g3114));
assign g5386 = (g5227)|(g669);
assign I2417 = ((~g774));
assign I7838 = ((~g5947));
assign I3723 = ((~g2158));
assign g5546 = ((~g5388));
assign g6878 = ((~I9101));
assign g4045 = (g3425&g123);
assign g5309 = ((~g5063));
assign g2160 = (g1624&g929);
assign g3311 = (g218&g2872);
assign I8907 = ((~g6702));
assign g3841 = (g3614)|(g3617);
assign g2787 = ((~g2405));
assign I3942 = ((~g1833));
assign g4162 = ((~I5562));
assign I3007 = ((~g1439));
assign g4871 = ((~I6599));
assign I4537 = ((~g2877));
assign g821 = ((~I1880));
assign g5227 = ((~g5019)&(~g3559));
assign I5320 = ((~g3559));
assign g6505 = ((~I8435));
assign I2724 = ((~g1220));
assign g4378 = (g410&g3792);
assign I8300 = ((~g6299));
assign g4493 = ((~I6001));
assign g4340 = (g3972&g3291);
assign I1841 = ((~g207));
assign I8778 = (g6612)|(g6611)|(g6609)|(g6607);
assign g6281 = ((~I7987)&(~I7988)&(~I7989)&(~I7990));
assign g5776 = ((~I7528))|((~I7529));
assign I4510 = ((~g2753));
assign I9014 = ((~g6820));
assign g6229 = ((~g6036));
assign g5439 = ((~g5261));
assign g3368 = (g2822&g2923);
assign g5418 = ((~g5162)&(~g5169));
assign g5915 = ((~I7679));
assign g2602 = ((~g2061));
assign I4410 = ((~g2088));
assign I5037 = ((~g3705));
assign g6032 = ((~g5770));
assign I4955 = ((~g3673));
assign g2106 = ((~g1378));
assign I3478 = ((~g1450));
assign g3031 = ((~I4246));
assign g2155 = ((~I3274));
assign I6437 = ((~g4501));
assign g2612 = ((~I3752));
assign I7232 = ((~g5372))|((~I7230));
assign g4549 = (g4416)|(g3013);
assign g1060 = ((~g107));
assign g5246 = (g5077)|(g2080);
assign g2687 = ((~I3833));
assign I2992 = ((~g1741));
assign g3186 = (g2449&g2515);
assign I3659 = ((~g1491));
assign g4524 = ((~I6084));
assign I6992 = ((~g5151));
assign g3532 = ((~g3212))|((~g2215))|((~g3007))|((~g2981));
assign g4186 = (g3973&g1395);
assign g5117 = ((~I6763));
assign g4314 = ((~g4080));
assign g2244 = ((~I3379));
assign g2119 = ((~g1391));
assign g2805 = ((~g2443));
assign I5753 = ((~g4022));
assign g3983 = ((~I5270))|((~I5271));
assign I5756 = ((~g3922));
assign g4100 = ((~I5382));
assign g3703 = (g2284&g2840);
assign I9110 = ((~g6864));
assign I2382 = ((~g719));
assign I4040 = (g1279&g2025&g1267);
assign I8863 = ((~g6700));
assign g5327 = (g5077)|(g4416)|(g3028);
assign g4625 = ((~g4267));
assign g1918 = ((~I3019));
assign g1560 = ((~g996)&(~g980));
assign g4837 = ((~g4473));
assign I7514 = ((~g5590));
assign g2653 = ((~I3797));
assign I4151 = ((~g2551))|((~I4150));
assign I2119 = ((~g688));
assign g1773 = ((~I2814));
assign I7042 = ((~g5310));
assign g4832 = (g4517&g4512);
assign I3400 = ((~g135))|((~I3398));
assign g2956 = ((~g1861));
assign I7358 = ((~g5565));
assign g6796 = ((~I8958));
assign g4385 = ((~I5862));
assign I6334 = ((~g4454));
assign g3867 = ((~I5094));
assign I9173 = ((~g6876));
assign I4471 = ((~g3040));
assign g3893 = ((~g3664))|((~g3656))|((~g3647));
assign g2853 = (g836&g2021);
assign I6474 = ((~g4541))|((~I6473));
assign g1706 = (g766&g719&g729);
assign g5452 = (g5315&g4612);
assign g4210 = ((~I5630));
assign g6276 = ((~I7960));
assign I2890 = ((~g1123));
assign g1578 = ((~I2552));
assign I6186 = ((~g4301))|((~I6185));
assign g4372 = (g406&g3790);
assign I7069 = ((~g5281));
assign g3742 = ((~I4920))|((~I4921));
assign g4004 = ((~I5301))|((~I5302));
assign g3538 = ((~g2588))|((~g2215))|((~g2197))|((~g2179));
assign g6118 = (g5911)|(g5619);
assign g3608 = (g2599&g2308);
assign g6829 = (g6806&g5958);
assign g5675 = (g64&g5574);
assign g798 = ((~I1868));
assign g1460 = ((~I2457));
assign g5530 = ((~I7270));
assign g1288 = ((~I2269));
assign I7150 = ((~g5355));
assign g6124 = (g5705&g5958);
assign g5774 = ((~I7517));
assign g3340 = (g2772&g2915);
assign g2752 = ((~g2343));
assign g2609 = ((~I3749));
assign g3777 = ((~g3388));
assign g3969 = ((~I5233));
assign g2175 = ((~I3316));
assign I9095 = ((~g6855));
assign g5140 = ((~I6798));
assign g1734 = ((~g952));
assign g4700 = ((~I6292));
assign g3489 = (g2607&g1861);
assign g6741 = ((~g6705))|((~g6461))|((~g4941));
assign g3190 = (g260&g2535);
assign I3457 = ((~g784))|((~I3455));
assign g6830 = (g6809&g5975);
assign I8488 = ((~g6426));
assign g1679 = ((~g985));
assign I8724 = ((~g6533));
assign g4380 = ((~I5851));
assign g6483 = (I8385)|(I8386)|(I8387);
assign I9158 = ((~g6887));
assign g3633 = (g2497&g3076);
assign I5359 = (g3518&g3521&g3526&g3530);
assign g5045 = ((~I6677));
assign g6931 = (g6741)|(g6929);
assign g6839 = ((~I9038));
assign g3733 = (g3325)|(g2733);
assign g5649 = ((~I7404));
assign g4428 = ((~I5933));
assign g2758 = (g2497&g1963);
assign g2802 = ((~g2437));
assign I4321 = ((~g1917));
assign g3232 = ((~I4495));
assign g1940 = ((~I3047));
assign g5331 = ((~I6995));
assign g4220 = ((~I5644));
assign g3663 = (g2215&g2779);
assign g5857 = ((~g5638))|((~g1552))|((~g1017))|((~g2062));
assign g4488 = (g1633&g4202);
assign g1838 = ((~g1595));
assign g5356 = (g5265&g1902);
assign g4851 = ((~I6561));
assign g5012 = (g4782)|(g4580);
assign g1321 = ((~I2318));
assign g1931 = ((~I3034));
assign I3698 = ((~g1570))|((~I3697));
assign I6078 = ((~g4387));
assign g3876 = ((~I5109));
assign I3413 = ((~g616))|((~I3411));
assign g3498 = ((~g2634));
assign g1011 = ((~I2050));
assign I7536 = ((~g5666))|((~I7534));
assign g5256 = ((~g5077));
assign I8884 = ((~g6704));
assign g2118 = ((~I3247));
assign g5165 = (g508&g4993);
assign g6189 = (g6060)|(g6035);
assign g4456 = (g3829&g4229);
assign I6812 = ((~g5110));
assign g1332 = ((~I2349));
assign I4261 = ((~g1857));
assign g2791 = ((~I3989))|((~I3990));
assign g5505 = ((~I7224))|((~I7225));
assign I6051 = ((~g4185));
assign g2497 = ((~I3626));
assign g5741 = ((~g5602));
assign g938 = ((~g59));
assign g6704 = (g6660)|(g492);
assign g4914 = ((~g4816));
assign I4243 = ((~g1853));
assign I5091 = ((~g3242));
assign g3191 = (g2497&g2538);
assign g4531 = ((~I6105));
assign g5584 = ((~I7346));
assign g1577 = ((~g1001));
assign g4406 = ((~I5913));
assign g6133 = (g5723&g5975);
assign g6913 = (g6900&g6898);
assign I3050 = ((~g1439));
assign g2268 = ((~I3419));
assign I5430 = ((~g3727));
assign g1190 = ((~I2199));
assign g4598 = (g1978&g4253);
assign g3504 = ((~g2675));
assign g6439 = ((~g6385)&(~g3733)&(~g4328)&(~g4314));
assign I4351 = ((~g2233));
assign I5424 = ((~g3725));
assign I2805 = ((~g1205));
assign g4371 = (g461&g3789);
assign g4227 = ((~g4059));
assign g4819 = ((~I6500))|((~I6501));
assign g5407 = ((~I7073));
assign g4701 = (g4596&g1378);
assign g3341 = (g2998&g2709);
assign g4536 = ((~I6118));
assign g2826 = ((~g2481));
assign g3488 = ((~g2728));
assign I5197 = ((~g3571))|((~I5195));
assign I1988 = ((~g224))|((~I1986));
assign g6844 = (I9057)|(I9058)|(I9059);
assign g5391 = ((~I7055));
assign g6893 = ((~I9146));
assign I7099 = ((~g574))|((~I7097));
assign g2934 = ((~g2004));
assign g6618 = ((~I8716));
assign g5061 = ((~I6701));
assign g5923 = ((~I7701));
assign I7245 = ((~g188))|((~I7244));
assign g4195 = ((~I5615));
assign g3421 = (g622&g2846);
assign I8521 = ((~g6495));
assign g2275 = ((~I3422));
assign I2385 = ((~g784));
assign I3268 = ((~g1656));
assign I3678 = ((~g1690));
assign g1328 = ((~I2337));
assign I8081 = (g4894)|(g4904)|(g4993)|(g4967);
assign g6729 = ((~I8881));
assign g6057 = ((~g5824));
assign I5418 = ((~g4036));
assign g5910 = (g5816&g5667);
assign g6571 = ((~I8597));
assign g6504 = ((~I8432));
assign I7528 = ((~g49))|((~I7527));
assign g1682 = ((~g829));
assign g2818 = ((~g2464));
assign g6447 = (g6340)|(g5938);
assign I3399 = ((~g1826))|((~I3398));
assign g6321 = (g3873&g6212);
assign g2813 = ((~g2457));
assign g1928 = ((~I3031));
assign I3755 = ((~g2125));
assign I5243 = ((~g3242))|((~I5242));
assign g5637 = (g4499&g5543);
assign g5233 = (g551&g4980);
assign g1291 = ((~I2278));
assign g2916 = (g1030&g2113);
assign g1969 = ((~I3080));
assign g3751 = (g3375)|(g2807);
assign g6486 = ((~g6363));
assign I6283 = ((~g4613));
assign I3864 = ((~g2044));
assign I4468 = ((~g2583));
assign I6783 = ((~g4822));
assign g1138 = ((~g102))|((~g98));
assign g4349 = (g441&g3775);
assign g4471 = (g4253&g332);
assign I8806 = ((~g6686));
assign g2446 = ((~I3581));
assign I6485 = ((~g4603));
assign g3644 = (g2197&g2755);
assign g3609 = (g2706&g2678);
assign g1935 = ((~I3040));
assign I7029 = ((~g5149));
assign g3522 = (g646&g2909);
assign g3929 = ((~g3373)&(~g3376));
assign g1410 = ((~g1233));
assign I6377 = ((~g4569));
assign I8591 = ((~g6448));
assign g3857 = (g3687)|(g3161);
assign g5171 = (g406&g4950);
assign I5998 = ((~g4157));
assign I7237 = ((~g179))|((~g5374));
assign g3837 = (g3609)|(g3613);
assign g1088 = ((~I2119));
assign I9131 = ((~g6855));
assign g5880 = ((~g5824));
assign g3905 = ((~g3512)&(~g478));
assign g3989 = (g3679)|(g3144);
assign I3505 = ((~g1305));
assign g3434 = (g2850&g857);
assign g2908 = ((~g536)&(~g2010)&(~g541));
assign I5637 = ((~g3914));
assign g3710 = ((~g3029));
assign g2293 = ((~g1567));
assign g3842 = (g3670)|(g3135);
assign g5308 = ((~I6963))|((~I6964));
assign g4353 = (g3989&g3332);
assign g4046 = (I5351&I5352);
assign g6824 = ((~I9005));
assign g1250 = ((~g123));
assign g2544 = ((~I3662));
assign g1290 = ((~I2275));
assign I9028 = ((~g6806));
assign I9035 = ((~g6812));
assign g4845 = ((~I6543));
assign g5468 = ((~I7150));
assign I5394 = ((~g4016));
assign g4511 = ((~I6045));
assign g2892 = ((~g1982));
assign I3059 = ((~g1519));
assign g5112 = ((~I6750));
assign g1395 = ((~I2428));
assign g4017 = ((~g107))|((~g3425));
assign g3971 = (g3644)|(g3099);
assign g2096 = ((~I3212));
assign g6491 = ((~g6373));
assign I3846 = ((~g284))|((~g2370));
assign I2485 = ((~g766));
assign g5813 = ((~I7612));
assign g2743 = ((~g2333));
assign I3970 = ((~g290))|((~g2518));
assign g2166 = (g1633&g161);
assign g4430 = (g4349)|(g4015);
assign g4265 = ((~I5716));
assign I7113 = ((~g5295));
assign g2008 = ((~g866))|((~g873))|((~g1784));
assign g5670 = ((~g5527));
assign I7640 = ((~g5773));
assign g2073 = (g1088&g1499);
assign I2700 = ((~g1173));
assign I3717 = ((~g2154));
assign I9052 = ((~g3598))|((~I9050));
assign g6313 = (g3841&g6194);
assign I4371 = ((~g2555));
assign I4437 = ((~g2108));
assign g4763 = ((~I6397));
assign I7355 = ((~g5535));
assign I6289 = ((~g4433));
assign I6269 = ((~g4655));
assign g3451 = ((~g2615));
assign I7541 = ((~g59))|((~g5669));
assign I4743 = ((~g2594));
assign g2323 = (g471&g1358);
assign g1905 = ((~I3004));
assign g3030 = ((~I4243));
assign g3309 = (g2243&g2695);
assign g4500 = (g4243)|(g2010);
assign I6096 = ((~g4397));
assign I5406 = ((~g3976));
assign I2707 = ((~g1190));
assign I7193 = ((~g5466));
assign g5603 = (g5504&g4911);
assign I2797 = ((~g798))|((~I2795));
assign g4043 = (g457&g3388);
assign g6650 = (g6580&g6235);
assign g4399 = ((~I5896));
assign I6406 = ((~g4473));
assign I6081 = ((~g4388));
assign g930 = ((~I1970))|((~I1971));
assign I4212 = ((~g804))|((~I4210));
assign g5077 = (g1612)|(g4694);
assign g6621 = ((~I8721));
assign I3800 = ((~g2145));
assign I8264 = ((~g6296));
assign I5933 = ((~g4346));
assign I2982 = ((~g1426));
assign I5537 = ((~g654))|((~I5535));
assign g2834 = (g1263&g1257&g1270&I4040);
assign g1586 = ((~g1052));
assign I8644 = ((~g6526));
assign g6243 = (g500&g5890);
assign g1659 = ((~I2638));
assign g6240 = (g4205&g5888);
assign I6315 = ((~g4446));
assign g2995 = ((~I4183))|((~I4184));
assign g6693 = (g6618&g6617);
assign g6468 = (g2032&g6394&g1609);
assign I9122 = ((~g6864));
assign I3148 = ((~g1595));
assign I4501 = ((~g2705));
assign I8594 = ((~g6446));
assign g2067 = ((~I3178))|((~I3179));
assign g2196 = ((~I3337));
assign g4609 = ((~I6182));
assign g3815 = (g3282)|(g2659);
assign g1375 = ((~I2411));
assign I3456 = ((~g1691))|((~I3455));
assign g6673 = (g6559)|(g6640)|(g4416)|(g2950);
assign I4433 = ((~g2103));
assign I5454 = ((~g3874));
assign g848 = ((~g594));
assign I5153 = ((~g3330));
assign g2555 = ((~I3672));
assign I7808 = ((~g5919));
assign g6842 = ((~I9047));
assign I7210 = ((~g5367))|((~I7208));
assign g4205 = (g3843)|(g541);
assign g2845 = ((~g2565));
assign g1534 = ((~I2498))|((~I2499));
assign I6666 = ((~g4740));
assign g3001 = ((~I4198));
assign I8171 = ((~g6170));
assign g4561 = ((~g4189));
assign I5056 = ((~g3567));
assign I5876 = ((~g3870));
assign I5926 = ((~g4153));
assign g6514 = ((~I8462));
assign I5696 = ((~g3942));
assign g3236 = ((~I4507));
assign I2776 = ((~g1192));
assign g5201 = (g4859&g5084);
assign g6151 = (g3209&g5997);
assign g3756 = ((~I4940))|((~I4941));
assign g6361 = ((~I8147));
assign I2854 = ((~g1236));
assign g2721 = (g2397&g1922);
assign g3502 = ((~g1411))|((~g1402))|((~g2795));
assign g2505 = ((~I3629));
assign g1733 = ((~I2741));
assign g1039 = ((~g662));
assign I6570 = ((~g4719));
assign g6644 = (g6575&g6230);
assign I8153 = ((~g6185));
assign g6886 = ((~I9125));
assign g4941 = (g4829)|(g4832);
assign g6084 = (g1123&g5753);
assign I2015 = ((~g260))|((~I2013));
assign g2001 = ((~I3112));
assign g4949 = (g193&g4753);
assign g5059 = ((~I6697));
assign I6918 = ((~g5124));
assign g2413 = ((~I3553));
assign g5381 = ((~I7039));
assign I2674 = ((~g710))|((~g131));
assign I3961 = ((~g1835));
assign g2897 = (g1030&g2062);
assign I6964 = ((~g586))|((~I6962));
assign I5094 = ((~g3705));
assign g3022 = ((~I4229));
assign g2924 = (g2095)|(g1573);
assign I8276 = ((~g6303));
assign g5434 = ((~I7110));
assign I6763 = ((~g4780));
assign I3247 = ((~g1791));
assign g6705 = (g6693)|(g4835);
assign g5193 = (g532&g4967);
assign g1275 = ((~g842));
assign I4495 = ((~g3022));
assign g3117 = (g218&g2367);
assign g2084 = (g1577&g1563);
assign I4920 = ((~g3522))|((~I4919));
assign g4783 = ((~I6441));
assign g6436 = ((~g6385)&(~g3733)&(~g4328)&(~g4080));
assign I3037 = ((~g1769));
assign g2777 = ((~I3965));
assign g5575 = ((~g5411));
assign g6345 = (g6273&g6083);
assign g2460 = ((~I3590));
assign g5695 = (g5635)|(g5483);
assign g3355 = ((~g3100));
assign g4492 = ((~I5998));
assign I5633 = ((~g3768));
assign g6014 = ((~g5824));
assign g3239 = ((~I4516));
assign g6659 = (g6634)|(g6631);
assign g5260 = ((~g4938));
assign I2218 = ((~g11));
assign g5892 = ((~g5742));
assign g2296 = ((~I3441));
assign g2866 = ((~g1905));
assign g2484 = ((~I3611));
assign g6329 = (g3888&g6212);
assign g5628 = (g5498)|(g3292);
assign I9074 = ((~g6844));
assign g4501 = (g4250&g1671);
assign I2287 = ((~g927));
assign I6792 = ((~g5097));
assign I6305 = ((~g4441));
assign g1115 = ((~g40));
assign g4512 = ((~I6048));
assign I7596 = ((~g5605));
assign I8875 = ((~g6697));
assign g1317 = ((~I2306));
assign g6287 = (g6241)|(g6082);
assign g1407 = (g301&g866);
assign g2405 = ((~I3543));
assign g4825 = ((~g4472))|((~g4465));
assign g6715 = ((~g6673));
assign g4622 = ((~g4252));
assign g4422 = ((~g4111));
assign g5052 = ((~I6692));
assign g3136 = ((~I4382));
assign g5908 = ((~g5753));
assign g4010 = ((~g3601));
assign g1222 = ((~I2225));
assign g5444 = (g4545&g5256&g1574);
assign g2768 = ((~g2367));
assign g4706 = ((~I6308));
assign g6521 = ((~I8479));
assign g5148 = ((~I6812));
assign g4874 = (g582&g4708);
assign I1917 = ((~g48));
assign g3040 = ((~I4255));
assign I2970 = ((~g1504));
assign g3618 = (g3016&g2712);
assign g4584 = ((~g4164)&(~g4168));
assign g3259 = ((~g2996));
assign g3540 = ((~I4762));
assign g6299 = (g5530&g6163);
assign g5179 = ((~g5099));
assign g4239 = ((~g3763)&(~g3296));
assign g5350 = (g5325&g3453);
assign I3331 = ((~g1631));
assign g5475 = ((~I7161));
assign I6750 = ((~g4771));
assign g3212 = ((~I4455));
assign g5375 = ((~I7029));
assign g3769 = ((~g3622));
assign I7490 = ((~g5583));
assign I8426 = ((~g6424));
assign g6258 = (g512&g5899);
assign g2138 = (g1639&g809);
assign I4203 = ((~g2255))|((~g743));
assign I2293 = ((~g971));
assign g847 = ((~g590));
assign I8082 = (g4980)|(g4915)|(g5025)|(g5054);
assign g3215 = ((~g2340))|((~g1402));
assign g4630 = (g4339)|(g3610);
assign g3007 = ((~g2197));
assign g3298 = (g2231&g2679);
assign g5545 = ((~g5331));
assign g5374 = (g5215)|(g4947);
assign g5956 = (g5783&g5425);
assign g5199 = ((~I6867));
assign I7856 = ((~g5994));
assign I2973 = ((~g1687));
assign g5812 = (g5376)|(g5618);
assign g1557 = ((~g1017));
assign g6623 = ((~I8727));
assign I8696 = ((~g6569));
assign g5357 = (g398&g5220);
assign g3208 = (g895&g2551);
assign g6262 = (g516&g5901);
assign I3488 = ((~g1295));
assign g3681 = (g2234&g2806);
assign I8368 = (g6148)|(g6321)|(g5176)|(g5184);
assign I3044 = ((~g1257));
assign g6231 = ((~g6044));
assign g5780 = ((~I7556))|((~I7557));
assign g3914 = ((~I5153));
assign g2330 = ((~g1777));
assign g6123 = (g5702&g5958);
assign g6592 = ((~I8644));
assign g5568 = ((~g5423));
assign I8629 = ((~g6544));
assign g6336 = (g6246&g6065);
assign g4228 = ((~I5668));
assign I3086 = ((~g1439));
assign g4491 = (g3554&g4215);
assign g3913 = (g3449)|(g2860);
assign g3678 = (g2256&g2802);
assign g6179 = (g6077)|(g6051);
assign g6798 = (g4946&g6781);
assign g1724 = ((~I2724));
assign g6692 = (g6616&g6615);
assign I3708 = ((~g1946));
assign I6540 = ((~g4714));
assign I6692 = ((~g4720));
assign g5219 = ((~I6885));
assign g1094 = ((~I2122));
assign g6056 = (g5824&g1699);
assign g6489 = ((~g6369));
assign I8674 = ((~g6521));
assign I3560 = ((~g1673));
assign g3114 = ((~I4362));
assign g5164 = (g437&g4877);
assign I3804 = ((~g2575));
assign I6723 = ((~g4761));
assign g6687 = (g6260)|(g6646);
assign g6901 = ((~I9170));
assign g2728 = ((~I3890));
assign g1846 = ((~I2940));
assign g4826 = (g4209&g4463);
assign I7346 = ((~g5531));
assign I1961 = ((~g520))|((~g242));
assign g4757 = (g4456)|(g4158);
assign g5050 = (g4285&g4807);
assign g2086 = ((~I3198));
assign I9077 = ((~g6845));
assign g5184 = (g453&g4877);
assign g3321 = (g2252&g2713);
assign g5794 = ((~I7593));
assign g4863 = (g4777&g2874);
assign I8632 = ((~g6548));
assign g3861 = ((~I5084));
assign g2670 = (g2029&g1503);
assign g4128 = ((~I5466));
assign g3939 = ((~g3340)&(~g3351));
assign g6746 = ((~I8916));
assign I2763 = ((~g1236));
assign g2981 = ((~g2179));
assign g5304 = ((~I6956));
assign g4354 = (g437&g3777);
assign g1979 = ((~I3090));
assign g1330 = ((~I2343));
assign g4117 = ((~I5433));
assign g6107 = ((~I7817));
assign I4681 = ((~g2947));
assign g1957 = ((~I3068));
assign I8693 = ((~g6570));
assign I5597 = ((~g3821));
assign g1894 = ((~I2989));
assign I2457 = ((~g1253));
assign g6158 = (g2594&g6015);
assign I5333 = ((~g3491));
assign I2306 = ((~g896));
assign g5521 = ((~I7261));
assign g4759 = (g536&g4500);
assign I2788 = ((~g1236));
assign g1345 = ((~I2382));
assign g4848 = ((~I6552));
assign I2108 = ((~g602))|((~g610));
assign g4714 = ((~I6324));
assign g6330 = ((~I8070));
assign g6295 = (g5379&g6162);
assign g921 = ((~g111));
assign g2650 = ((~I3794));
assign g4379 = ((~I5848));
assign g4677 = (g4652&g4646);
assign g5488 = (g394&g5331);
assign g3622 = ((~I4821));
assign g5152 = (g430&g4950);
assign g3384 = ((~g2834));
assign g3932 = ((~I5169));
assign I3152 = ((~g1322));
assign g4617 = ((~g4242));
assign g1358 = ((~g1119));
assign g6533 = ((~I8515));
assign I4414 = ((~g2090));
assign g4123 = ((~I5451));
assign g4169 = (g3966&g2099);
assign g6312 = ((~I8040));
assign g4797 = (g4593&g4643);
assign g2618 = ((~I3758));
assign g3356 = (g248&g2888);
assign g2525 = ((~I3650));
assign g2242 = ((~I3373));
assign g5993 = ((~g5872));
assign I8444 = ((~g6421));
assign g4059 = (g3466)|(g3425);
assign g5714 = ((~I7475));
assign g4752 = (g4452)|(g4155);
assign I8229 = ((~g6330));
assign g5060 = (g3491)|(g4819);
assign I3225 = ((~g1813));
assign g5824 = ((~g5631));
assign I1853 = ((~g211));
assign I5910 = ((~g3750));
assign g2695 = ((~I3843));
assign g3334 = (g236&g2883);
assign g4187 = ((~I5591));
assign I2091 = ((~g29))|((~I2089));
assign g6657 = ((~I8767));
assign g4277 = (g3936&g942);
assign g2320 = ((~I3474));
assign I2940 = ((~g1653));
assign g6357 = ((~I8117)&(~I8118)&(~I8119)&(~I8120));
assign g3630 = (g3167&g1756);
assign g3852 = ((~I5065));
assign I4420 = ((~g2096));
assign g6645 = (g6576&g6231);
assign I3352 = ((~g1285));
assign g3628 = (g2449&g3070);
assign g4624 = ((~g4265));
assign I6015 = ((~g4170));
assign I7439 = ((~g5515))|((~g594));
assign g5576 = ((~g5415));
assign g1832 = ((~I2910));
assign g2408 = ((~I3546));
assign I1832 = ((~g143));
assign g3187 = ((~I4424));
assign I3284 = ((~g1702));
assign g5667 = ((~g5524));
assign g6892 = ((~I9143));
assign g2060 = ((~g1369));
assign I5618 = ((~g3821));
assign g3770 = ((~I4961));
assign I2870 = ((~g1161));
assign I7542 = ((~g59))|((~I7541));
assign g5457 = ((~g5304));
assign g5265 = ((~g4863)&(~g4865));
assign I8462 = ((~g6430));
assign I8258 = ((~g6293));
assign g4001 = (g3702)|(g3190);
assign I2593 = ((~g1177));
assign g2686 = ((~I3830));
assign I8940 = ((~g6783));
assign g6400 = ((~I8208)&(~I8209)&(~I8210)&(~I8211));
assign g3806 = (g3384&g2024);
assign I3411 = ((~g1419))|((~g616));
assign I9065 = (g6158)|(g6333)|(g5152)|(g5156);
assign g5018 = (g4791)|(g4597);
assign g2659 = (g1686&g2296);
assign I5767 = ((~g3961))|((~I5766));
assign g2870 = ((~g2296));
assign I5006 = ((~g3604));
assign g4599 = (g3499)|(g4230);
assign g3512 = (g2928&g1764);
assign I7534 = ((~g54))|((~g5666));
assign I2491 = ((~g821));
assign I2967 = ((~g1682));
assign g6316 = (g3855&g6194);
assign g4151 = ((~I5536))|((~I5537));
assign g1477 = ((~g952));
assign g5551 = ((~I7295));
assign g4684 = (g4584&g1341);
assign g6555 = (g1838&g6469);
assign g2753 = ((~I3927));
assign I6185 = ((~g4301))|((~g3955));
assign g3539 = ((~g2591))|((~g2215))|((~g2197))|((~g2981));
assign I6434 = ((~g4622));
assign g4386 = ((~I5865));
assign g5292 = ((~I6942));
assign I1979 = ((~g512))|((~I1978));
assign g2178 = ((~I3325));
assign I9051 = ((~g6832))|((~I9050));
assign I2635 = ((~g1055));
assign g6115 = ((~g5879));
assign g4838 = (g4648&g84);
assign g4146 = ((~I5520));
assign I3105 = ((~g1439));
assign g6926 = (g6798)|(g6923);
assign I6789 = ((~g4871));
assign g6280 = ((~I7978)&(~I7979)&(~I7980)&(~I7981));
assign g4373 = (g4001&g3370);
assign g2333 = ((~I3485));
assign g5698 = (g5648)|(g5486);
assign I6390 = ((~g4504))|((~g4610));
assign g3533 = (g3154)|(g3166);
assign g6877 = ((~I9098));
assign g6480 = (I8360)|(g6359);
assign g3957 = ((~I5196))|((~I5197));
assign g5939 = (g5776&g5395);
assign I3764 = ((~g2044));
assign g927 = ((~I1958));
assign g2955 = (g2381&g297);
assign I9152 = ((~g6889));
assign g4736 = ((~I6366));
assign g6795 = (g4867)|(g6772);
assign g1205 = ((~g45));
assign I3916 = ((~g2449))|((~I3914));
assign g6277 = ((~I7963));
assign I6801 = ((~g5045));
assign g3287 = (g135&g2865);
assign g6148 = (g3196&g6015);
assign g3433 = (g1359&g2831&g905);
assign g5950 = ((~g5730));
assign g2367 = ((~I3519));
assign g2944 = ((~g269))|((~g2381));
assign g4393 = ((~I5882));
assign g3847 = ((~I5056));
assign g4433 = (g4354)|(g4032);
assign g2312 = ((~I3462));
assign I8891 = ((~g6706));
assign g1783 = ((~I2831));
assign g1627 = ((~I2584));
assign g6033 = ((~g5824));
assign g1656 = ((~I2635));
assign g6519 = ((~I8473));
assign I4593 = ((~g2966));
assign g6100 = ((~I7796));
assign I6495 = ((~g4607));
assign g5872 = ((~g5649))|((~g1557))|((~g1564))|((~g2113));
assign g6366 = ((~I8162));
assign g4132 = ((~I5478));
assign I6036 = ((~g4370));
assign g4643 = ((~g4293));
assign I8201 = ((~g478))|((~g6192));
assign I5307 = ((~g478))|((~g3512));
assign I2986 = ((~g1504));
assign g4760 = ((~I6386));
assign g2410 = ((~I3550));
assign I4331 = ((~g2555));
assign g1351 = ((~I2388));
assign I6942 = ((~g5124));
assign g5518 = ((~I7258));
assign g6567 = ((~I8585));
assign g5773 = ((~I7514));
assign I4941 = ((~g357))|((~I4939));
assign g3613 = (g2604&g2312);
assign g2105 = ((~g1375));
assign g4110 = ((~I5412));
assign I2245 = ((~g567))|((~I2244));
assign g5622 = (g5492)|(g3277);
assign g6110 = (g5883)|(g5996);
assign I4398 = ((~g2086));
assign I1844 = ((~g208));
assign I7578 = ((~g5680))|((~I7576));
assign I4424 = ((~g2097));
assign g3365 = (g254&g2892);
assign g6352 = ((~I8110));
assign I4211 = ((~g2294))|((~I4210));
assign g2172 = ((~I3307));
assign I3161 = ((~g1270));
assign g5775 = ((~I7521))|((~I7522));
assign g6076 = ((~g5797));
assign g1875 = ((~I2970));
assign I7966 = ((~g6166));
assign g1814 = ((~I2873));
assign I4358 = ((~g2525));
assign I7116 = ((~g5299));
assign g4341 = (g3977&g3297);
assign g3312 = ((~I4587));
assign I6087 = ((~g4392));
assign g5497 = (g5447&g3458);
assign I3004 = ((~g1426));
assign g2113 = (g1576&g1535);
assign I5169 = ((~g3593));
assign I3425 = ((~g1274));
assign g1030 = ((~I2057));
assign I8614 = ((~g6537));
assign I4455 = ((~g2118));
assign g3023 = ((~g2215));
assign I4226 = ((~g2525));
assign I6677 = ((~g4757));
assign I2735 = ((~g1118));
assign g5226 = (g672&g5054);
assign g3014 = ((~I4217));
assign I5053 = ((~g3710));
assign g6506 = ((~I8438));
assign I6949 = ((~g5050));
assign I8779 = (g6605)|(g6656)|(g6654)|(g6652);
assign g6562 = ((~I8570));
assign g1528 = ((~g878));
assign I1994 = ((~g504))|((~g218));
assign g2156 = (g815&g1642);
assign g3369 = ((~I4646));
assign I2574 = (g804&g798&g791);
assign g5684 = ((~I7440))|((~I7441));
assign g3162 = ((~I4402));
assign g6699 = ((~I8815));
assign I2037 = ((~g679));
assign g5067 = ((~g4801));
assign g4158 = ((~I5556));
assign g3267 = ((~g3030));
assign I3644 = ((~g1685));
assign I3933 = ((~g288))|((~g2473));
assign g4946 = (g4830)|(g4833);
assign I4507 = ((~g2739));
assign I5615 = ((~g3914));
assign g1966 = ((~I3077));
assign g4740 = (g4448)|(g4154);
assign I4587 = ((~g2962));
assign g5247 = ((~g4900));
assign I8647 = ((~g6528));
assign I7799 = ((~g5918));
assign g4080 = (g3302)|(g2700);
assign I7055 = ((~g5318));
assign I5078 = ((~g3719));
assign g3300 = (g2232&g2682);
assign g4308 = ((~I5777));
assign I8588 = ((~g6443));
assign g6499 = ((~I8417));
assign g5953 = (g5781&g5415);
assign I6023 = ((~g4151));
assign g1643 = ((~I2608));
assign g2090 = ((~I3206));
assign I7487 = ((~g5684));
assign g5638 = ((~I7397));
assign g3750 = (g3372)|(g2794);
assign g4434 = (g4355)|(g4033);
assign g2664 = ((~I3808));
assign g6925 = ((~I9208));
assign g1480 = ((~g985));
assign I6874 = ((~g4861));
assign I5388 = ((~g3969));
assign I8189 = ((~g6179));
assign g3926 = ((~g3338)&(~g3350));
assign g6446 = ((~g6385)&(~g4334)&(~g4092)&(~g4314));
assign I5487 = ((~g3881));
assign g3682 = (g2772&g2430);
assign g4445 = (g4235&g1854);
assign I2315 = ((~g1222));
assign I4150 = ((~g2551))|((~g139));
assign g4334 = ((~g3733));
assign g6619 = (g6515&g6115);
assign g5533 = (g5351)|(g3290);
assign g952 = ((~I2029));
assign g5604 = (g5059&g5521);
assign g2409 = ((~g1815));
assign g6160 = ((~g5926));
assign g6075 = ((~g269)&(~g5863));
assign g6914 = (g6895&g6893);
assign g2867 = ((~g1908));
assign g3336 = (g2760&g1911);
assign g5621 = (g5508&g4943);
assign g946 = ((~g361));
assign I7238 = ((~g179))|((~I7237));
assign g2294 = (g1716&g791&g798);
assign I7441 = ((~g594))|((~I7439));
assign I5508 = ((~g3867));
assign g6730 = ((~I8884));
assign g1934 = ((~I3037));
assign g6307 = (g6262)|(g6096);
assign I5242 = ((~g3242))|((~g3247));
assign g5895 = ((~g5742));
assign g2026 = (g1359&g1402&g1398&g901);
assign g4579 = ((~g4206));
assign I5545 = ((~g3814));
assign g6253 = (g508&g5896);
assign g3659 = (g2672&g2361);
assign g3904 = ((~g3575));
assign g900 = ((~I1927));
assign g4108 = ((~I5406));
assign g3836 = ((~I5033));
assign I4276 = ((~g2170));
assign I8220 = ((~g6322));
assign g1678 = ((~I2658));
assign I3140 = ((~g1317));
assign g4915 = ((~g4669));
assign g1782 = ((~I2828));
assign g5467 = (g3868)|(g5318)|(g3992);
assign g1329 = ((~I2340));
assign g3970 = ((~I5236));
assign I3258 = ((~g1760));
assign g2931 = ((~g1988));
assign I3513 = ((~g1450));
assign g2889 = ((~g1975));
assign g1825 = ((~I2893));
assign g6910 = (g6892&g6891);
assign g6437 = (g6302)|(g6121);
assign g3771 = ((~I4964));
assign I6253 = ((~g4608));
assign g2827 = ((~g2485));
assign g1394 = ((~g1206));
assign g6809 = ((~I8981));
assign g2117 = ((~I3244));
assign g1273 = ((~g839));
assign g5011 = ((~I6649));
assign g6821 = ((~g6785));
assign I4300 = ((~g2234));
assign g4058 = (g3424&g1246);
assign g4679 = ((~I6269));
assign I6057 = ((~g4379));
assign g6716 = (g6682&g932);
assign g3881 = ((~I5116));
assign I2995 = ((~g1742));
assign I5119 = ((~g3714));
assign g4550 = ((~I6126));
assign g4537 = ((~g4410));
assign I5493 = ((~g3834));
assign g2803 = ((~g2440));
assign g3784 = (g114&g3251);
assign g1943 = ((~I3050));
assign I8570 = ((~g6433));
assign g5136 = ((~I6786));
assign I3316 = ((~g1344));
assign g1326 = ((~g894));
assign g6742 = ((~g6683))|((~g932))|((~g6716));
assign g6876 = ((~I9095));
assign I5591 = ((~g3821));
assign g5889 = ((~g5742));
assign g4453 = (g4238&g1858);
assign I7811 = ((~g5921));
assign I6400 = ((~g4473));
assign g4364 = ((~I5825));
assign I7689 = ((~g5708));
assign g5364 = (g574&g5194);
assign g4427 = (g4373)|(g3668);
assign I3212 = ((~g1806));
assign g6898 = ((~I9161));
assign g6441 = ((~I8309));
assign g6481 = (I8367)|(I8368)|(I8369)|(I8370);
assign g6457 = (g6352)|(g6347);
assign g5945 = (g5118&g5801);
assign g1576 = (g1101&g1094);
assign I5196 = ((~g3567))|((~I5195));
assign g5662 = (g5553)|(g5402);
assign g6703 = (g6692)|(g4831);
assign g3965 = ((~g3359)&(~g3367));
assign g4515 = ((~I6057));
assign g2790 = ((~g2413));
assign I3675 = ((~g1491));
assign g6126 = (g5711&g5958);
assign g6599 = ((~I8665));
assign g4802 = ((~I6470));
assign I2696 = ((~g1156));
assign g3662 = (g2544&g3114);
assign g6620 = (g6516&g6117);
assign g2254 = ((~I3391));
assign g2461 = ((~I3593));
assign g6451 = ((~g6385)&(~g4334)&(~g4328)&(~g4314));
assign I2949 = ((~g1263));
assign g5431 = ((~I7098))|((~I7099));
assign g937 = ((~I1979))|((~I1980));
assign g3656 = ((~g2769)&(~g2757)&(~g2745));
assign g804 = ((~I1871));
assign g3732 = (g3324)|(g2732);
assign I7501 = ((~g5596));
assign g4405 = ((~I5910));
assign g1638 = ((~g754));
assign g2267 = (g1716&g791);
assign g3093 = ((~I4334));
assign I5351 = (g3511&g3517&g3520&g3525);
assign g3233 = ((~I4498));
assign g6212 = ((~I7910));
assign g5951 = (g5780&g5411);
assign g4489 = (g2166&g4206);
assign g5618 = (g5506&g4933);
assign g4042 = (g406&g3388);
assign g3505 = (g2924&g1749);
assign I6132 = ((~g4219));
assign g4639 = ((~g4289));
assign I3465 = ((~g1724));
assign g3647 = ((~g2731)&(~g2719)&(~g2698));
assign I3455 = ((~g1691))|((~g784));
assign g4779 = ((~g4461)&(~g4464));
assign I2346 = ((~g1193));
assign I5065 = ((~g3714));
assign g2921 = ((~g1950));
assign g4507 = ((~I6033));
assign g2713 = ((~I3868));
assign g2085 = (g1123&g1567);
assign g2214 = ((~I3349));
assign g1917 = ((~I3016));
assign I6701 = ((~g4726));
assign I7246 = ((~g5377))|((~I7244));
assign g6609 = ((~I8693));
assign g2962 = ((~g2008));
assign g6152 = (g3212&g6015);
assign g6885 = ((~I9122));
assign g5066 = (g4668)|(g4672);
assign g4020 = ((~I5324));
assign g6405 = ((~I8229));
assign g2884 = ((~g1957));
assign g3679 = (g2245&g2803);
assign I6349 = ((~g4569));
assign g3135 = (g2370&g2416);
assign I3662 = ((~g1688));
assign g6634 = (g1595&g6545);
assign g6708 = ((~I8834));
assign g5200 = (g559&g5025);
assign I3235 = ((~g1807));
assign g5487 = (g390&g5331);
assign I8984 = ((~g6794));
assign I4921 = ((~g650))|((~I4919));
assign g2619 = ((~I3761));
assign g3237 = ((~I4510));
assign g4731 = ((~I6359));
assign g5157 = (g496&g4904);
assign g5084 = ((~g4727));
assign g6415 = ((~I8255));
assign g2044 = ((~I3161));
assign I7264 = ((~g5458));
assign g6083 = ((~g5809));
assign I3398 = ((~g1826))|((~g135));
assign g6346 = (g6274&g6087);
assign g3328 = (g2701&g1894);
assign g4616 = (g4231&g3761);
assign g6513 = ((~I8459));
assign I4023 = ((~g2315));
assign g6651 = ((~I8749));
assign g3835 = ((~I5030));
assign g5504 = ((~I7217))|((~I7218));
assign I7190 = ((~g5432));
assign g2241 = ((~I3370));
assign g5380 = (g188&g5264);
assign g1333 = ((~I2352));
assign I3364 = ((~g1648));
assign g5627 = (g5497)|(g3286);
assign g4784 = ((~I6444));
assign g4685 = (g4591&g2079);
assign g3896 = (g3689)|(g3697);
assign g6286 = (g6238)|(g6079);
assign g1289 = ((~I2272));
assign g5232 = (g548&g4980);
assign I5302 = ((~g3505))|((~I5300));
assign g5909 = (g5787&g3384);
assign g6938 = ((~I9227));
assign g5192 = (g1046&g4894);
assign g1038 = ((~g127));
assign I5043 = ((~g3247));
assign g6789 = (g3764)|(g6769);
assign g5261 = ((~I6918));
assign g1470 = ((~g937)&(~g930)&(~g928));
assign I8243 = ((~g6286));
assign I4545 = ((~g2853))|((~g353));
assign I2507 = ((~g1047))|((~I2506));
assign I7007 = ((~g5314));
assign g6656 = ((~I8764));
assign g1316 = ((~I2300))|((~I2301));
assign I1865 = ((~g279));
assign I3337 = ((~g1338));
assign I2952 = ((~g1594));
assign I8295 = ((~g6295));
assign g4510 = ((~I6042));
assign g4194 = ((~I5612));
assign g4823 = ((~I6507));
assign I4217 = ((~g2163));
assign g2485 = ((~I3614));
assign g5865 = ((~g5649))|((~g1088))|((~g1076))|((~g2068));
assign I3858 = ((~g2197));
assign g4567 = ((~I6139));
assign g2009 = ((~g901))|((~g1387))|((~g905));
assign I9041 = ((~g6835));
assign g4140 = ((~I5502));
assign g5111 = ((~I6744))|((~I6745));
assign g1221 = ((~g46));
assign g3335 = (g230&g2884);
assign g3452 = ((~g2625));
assign g3002 = ((~g2215));
assign I5188 = ((~g3589))|((~I5187));
assign g6241 = (g1325&g5887);
assign g2145 = ((~I3268));
assign g3466 = ((~I4706));
assign g2437 = ((~I3572));
assign g4284 = ((~I5739));
assign g6766 = (g6750&g2986);
assign g6490 = ((~g6371));
assign I2527 = ((~g766))|((~I2526));
assign g2165 = ((~I3294));
assign I7187 = ((~g5387));
assign I2741 = ((~g1222));
assign I2131 = ((~g24));
assign I8518 = ((~g6494));
assign I3271 = ((~g1748));
assign g5441 = (g4537&g5251&g1558);
assign I4050 = ((~g2059));
assign g2068 = (g1541&g1546);
assign g1857 = ((~I2961));
assign g5098 = (g4021&g4837);
assign g3875 = ((~I5106));
assign g3352 = (g2796&g2920);
assign g5158 = (g504&g4993);
assign I7161 = ((~g5465));
assign g931 = ((~g54));
assign g6082 = (g1123&g5742);
assign I3971 = ((~g290))|((~I3970));
assign g3464 = (g341&g2956);
assign g3982 = (g3663)|(g3127);
assign g2099 = ((~g1366));
assign I6766 = ((~g4783));
assign g5975 = ((~g5821));
assign g6089 = (g1143&g5731);
assign I4986 = ((~g3638));
assign g1535 = ((~g1088));
assign g6777 = (g6762&g3488);
assign g3816 = (g3434&g861);
assign I6798 = ((~g5042));
assign g1044 = ((~I2081))|((~I2082));
assign g3960 = ((~I5204));
assign g4744 = (g3434&g4582);
assign g6797 = ((~I8961));
assign g4852 = ((~I6564));
assign g1950 = ((~I3059));
assign g2391 = ((~I3534));
assign I3720 = ((~g2155));
assign g2430 = ((~I3563));
assign g2950 = (g2156&g1612);
assign g2759 = (g2473&g1966);
assign g5172 = (g441&g4877);
assign I8958 = ((~g6774));
assign g6238 = (g528&g5886);
assign g3759 = (g2644&g3498);
assign I6292 = ((~g4434));
assign I3376 = ((~g1328));
assign g2842 = ((~I4050));
assign g6790 = (g3765)|(g6773);
assign I8854 = ((~g6696));
assign I7352 = ((~g5533));
assign I7339 = ((~g5540));
assign g3359 = (g2822&g2922);
assign g3046 = ((~I4267));
assign g985 = ((~g638));
assign g3104 = ((~I4351));
assign I8267 = ((~g6297));
assign g5912 = ((~g5853));
assign I8120 = (g4915)|(g5025);
assign I3794 = ((~g2044));
assign I3379 = ((~g1647));
assign I3525 = ((~g1461));
assign g4816 = ((~g996))|((~g4550))|((~g1518))|((~g2073));
assign g6713 = ((~g6679));
assign I8774 = (g6655)|(g6653)|(g6651)|(g6649);
assign g5360 = (g4431&g5160);
assign I5568 = ((~g3897));
assign g2095 = ((~g1584))|((~g749))|((~g736));
assign I8981 = ((~g6793));
assign g5570 = ((~g5392));
assign g4021 = (g3558)|(g2949);
assign g1331 = ((~I2346));
assign g5672 = (g5557)|(g5414);
assign g3338 = (g3162&g2914);
assign g6712 = ((~g6676));
assign g3322 = ((~g3070));
assign g3182 = (g2473&g2512);
assign g6686 = (g6259)|(g6645);
assign g5605 = (g3575)|(g5500);
assign g3085 = ((~I4324));
assign I5716 = ((~g3942));
assign I2464 = ((~g850));
assign g6646 = (g6577&g6232);
assign g2860 = (g710&g2296);
assign g4929 = ((~I6621));
assign g4397 = ((~I5890));
assign I3215 = ((~g1820));
assign g6888 = ((~I9131));
assign g4849 = ((~I6555));
assign I2552 = ((~g971));
assign g2920 = ((~g1947));
assign I3096 = ((~g1439));
assign I3169 = ((~g1540))|((~I3168));
assign g3234 = ((~I4501));
assign I8249 = ((~g6289));
assign I3752 = ((~g2044));
assign g1883 = ((~g1797));
assign g3995 = (g3690)|(g3170);
assign I3188 = ((~g1716))|((~g791));
assign g2215 = ((~I3352));
assign I3823 = ((~g2125));
assign g5248 = ((~g4911));
assign g2256 = ((~I3395));
assign I8119 = (g5202)|(g4993)|(g4967)|(g4980);
assign g2997 = ((~I4192));
assign g6695 = ((~I8803));
assign I2364 = ((~g1143));
assign g5110 = ((~I6740));
assign g4633 = ((~g4284));
assign g6825 = ((~I9008));
assign g1036 = ((~I2061))|((~I2062));
assign g4289 = ((~I5746));
assign I8240 = ((~g6287));
assign I7176 = ((~g5437));
assign I5761 = ((~g3503))|((~I5759));
assign g913 = ((~g658));
assign g2434 = ((~g1064))|((~g1070))|((~g1620));
assign g6461 = (g6353)|(g6351);
assign I8515 = ((~g6492));
assign g3133 = (g236&g2410);
assign I8815 = ((~g6689));
assign g2029 = ((~I3134));
assign g6788 = (g3760)|(g6767);
assign g1564 = ((~g1030));
assign I5987 = ((~g4224));
assign I8678 = ((~g6565));
assign I2897 = ((~g1027))|((~g634));
assign I6004 = ((~g4159));
assign I8456 = ((~g6417));
assign g1423 = ((~I2442));
assign g3999 = (g3699)|(g3181);
assign I2821 = ((~g1221));
assign I3080 = ((~g1519));
assign I3382 = ((~g1284));
assign g6522 = ((~I8482));
assign g3371 = (g260&g2904);
assign I3367 = ((~g1283));
assign I6867 = ((~g5082));
assign g5593 = ((~I7355));
assign I3294 = ((~g1720));
assign I7978 = (g6194)|(g5958)|(g5975)|(g5997);
assign g858 = ((~g301));
assign g1348 = ((~I2385));
assign g4904 = ((~g4812));
assign g2061 = ((~I3169))|((~I3170));
assign g6305 = ((~I8027));
assign I2330 = ((~g1122));
assign g4051 = (g449&g3388);
assign g5500 = (g5430&g5074);
assign g5173 = (g512&g4993);
assign g3980 = ((~I5264));
assign g2538 = ((~I3656));
assign g4104 = ((~I5394));
assign g3575 = ((~I4777));
assign I4903 = ((~g3223));
assign I8473 = ((~g6485));
assign I8531 = ((~g6444));
assign I4382 = ((~g2265));
assign I7679 = ((~g5726));
assign I1932 = ((~g667));
assign I2904 = ((~g1256));
assign g5890 = ((~g5753));
assign g6707 = ((~I8831));
assign g1660 = ((~g985));
assign I8156 = ((~g6167));
assign g4793 = (g4277&g4639);
assign g1645 = ((~I2614));
assign I4546 = ((~g2853))|((~I4545));
assign g1175 = ((~g42));
assign g4656 = (g4369)|(g3662);
assign g4202 = ((~I5622));
assign I8107 = ((~g6136));
assign I2703 = ((~g1189));
assign g6516 = ((~g6409));
assign g3643 = (g2518&g3086);
assign I4182 = ((~g2292))|((~g749));
assign g3123 = (g230&g2391);
assign I5640 = ((~g3770));
assign g6469 = (g2121&g2032&g6394);
assign g5708 = ((~I7469));
assign g4683 = (g4585&g2066);
assign g1474 = ((~g760)&(~g754));
assign I8394 = (g6154)|(g6329)|(g5186)|(g5172);
assign g4147 = ((~I5523));
assign I9182 = ((~g6879));
assign I5439 = ((~g3730));
assign g1502 = ((~g709));
assign g4464 = (g4272&g1937);
assign I8453 = ((~g6414));
assign g1047 = ((~I2090))|((~I2091));
assign g4229 = ((~g4059));
assign g5224 = (g5123)|(g3630);
assign I3729 = ((~g2436));
assign g6170 = (g6061)|(g6014);
assign g6116 = (g5910)|(g5617);
assign g6153 = (g3216&g5997);
assign g6424 = ((~I8282));
assign I5360 = (g3532&g3536&g3539&g3544);
assign g5560 = (g5044&g5456);
assign I4757 = ((~g2861));
assign g3049 = ((~I4270));
assign I4019 = ((~g1841));
assign g5264 = ((~g4943));
assign I9230 = ((~g6936));
assign g3196 = ((~I4433));
assign g1731 = ((~I2735));
assign g5723 = ((~I7484));
assign g6242 = (g2356)|(g6075);
assign g5122 = (g193&g4662);
assign g1650 = ((~I2627));
assign g5599 = (g5049&g5512);
assign I2671 = ((~g1017));
assign I3304 = ((~g1740));
assign g1671 = ((~g985));
assign g5509 = ((~I7251));
assign I3334 = ((~g1330));
assign g5503 = (g366&g5384);
assign g6068 = (g5824&g1726);
assign g6324 = (g3880&g6212);
assign g6449 = ((~g6385)&(~g4334)&(~g4328)&(~g4080));
assign g4426 = ((~I5929));
assign g3625 = (g2619&g2320);
assign g873 = ((~g306));
assign I8386 = (g6152)|(g6327)|(g5183)|(g5177);
assign I3848 = ((~g2370))|((~I3846));
assign g3882 = ((~I5119));
assign g1937 = ((~I3044));
assign g6440 = (g6336)|(g5935);
assign g3503 = (g3122)|(g3132);
assign g865 = ((~g188));
assign g3699 = (g2276&g2836);
assign g5873 = ((~g5649))|((~g1017))|((~g1564))|((~g2113));
assign g5678 = (g5560)|(g5428);
assign I6410 = ((~g4473));
assign g2233 = ((~I3364));
assign g6933 = ((~I9220));
assign I2828 = ((~g1193));
assign g3907 = (g650&g3522);
assign I5496 = ((~g3839));
assign g6127 = (g5714&g5975);
assign I6558 = ((~g4705));
assign g3956 = ((~g3337)&(~g3349));
assign I3370 = ((~g1805));
assign g1570 = (g634&g1027);
assign I4255 = ((~g2179));
assign g3283 = (g2609&g2622);
assign g4809 = ((~I6485));
assign I8183 = ((~g6176));
assign I5890 = ((~g3878));
assign g2793 = (g2568&g1991);
assign g854 = ((~g646));
assign g1416 = (g913&g266);
assign g5094 = ((~g4685)&(~g4686));
assign g4788 = ((~I6452));
assign g3242 = ((~g3083));
assign I4220 = ((~g2164));
assign I3126 = ((~g1279))|((~I3125));
assign g5241 = (g5069)|(g2067);
assign g3460 = ((~g2667));
assign g3962 = ((~I5214));
assign g5661 = ((~g5518));
assign g4514 = ((~I6054));
assign I2867 = ((~g1143));
assign g5860 = ((~g5634));
assign g1749 = ((~I2767))|((~I2768));
assign I5027 = ((~g3267));
assign g5432 = ((~I7104));
assign I5293 = ((~g3421))|((~I5292));
assign I2614 = ((~g1123));
assign g5801 = ((~I7600));
assign g6574 = ((~g6484));
assign I7239 = ((~g5374))|((~I7237));
assign g1837 = ((~I2925));
assign g4299 = ((~I5756));
assign g1836 = ((~I2922));
assign g3665 = (g2748&g2378);
assign I8270 = ((~g6300));
assign g5139 = ((~I6795));
assign g1788 = ((~g985));
assign g2968 = ((~g2179));
assign g6040 = ((~g5824));
assign g3813 = ((~g3258));
assign g4592 = (g3147&g4281);
assign g2599 = ((~I3729));
assign g6311 = (g3837&g6194);
assign I8211 = (g4915)|(g5025);
assign g4517 = ((~I6063));
assign g2973 = ((~I4170));
assign g4532 = ((~I6108));
assign I8597 = ((~g6445));
assign g3838 = ((~I5037));
assign I3876 = ((~g2397))|((~I3874));
assign I2029 = ((~g677));
assign I2712 = ((~g1203));
assign g4947 = (g184&g4741);
assign g4250 = ((~I5702));
assign g4666 = (g4630&g4627);
assign I7600 = ((~g5605));
assign g4322 = ((~I5793));
assign g4877 = ((~g952)&(~g4680));
assign g2644 = ((~I3788));
assign g6802 = ((~I8972));
assign I3638 = ((~g1484));
assign g4521 = ((~I6075));
assign I8579 = ((~g6438));
assign g4808 = ((~g4473));
assign I5851 = ((~g3739));
assign g6408 = ((~g6283));
assign g5044 = (g4797)|(g4602);
assign I3989 = ((~g291))|((~I3988));
assign g6288 = (g5615&g6160);
assign g5220 = ((~g4903));
assign I3770 = ((~g2145));
assign g3545 = ((~g3085));
assign I9008 = ((~g6818));
assign g6438 = ((~g6376)&(~g4323)&(~g4074)&(~g4068));
assign g5017 = (g4784&g1679);
assign I9044 = ((~g6836));
assign I3301 = ((~g1730));
assign I5536 = ((~g3907))|((~I5535));
assign I5499 = ((~g3847));
assign g2594 = ((~I3723));
assign g3654 = (g2518&g3100);
assign g3199 = ((~g1861));
assign I8002 = ((~g6110));
assign g846 = ((~g586));
assign I3065 = ((~g1426));
assign g1559 = ((~g965));
assign g6624 = ((~I8730));
assign g4857 = ((~I6579));
assign I8527 = ((~g6440));
assign g5392 = ((~I7058));
assign I8910 = ((~g6730));
assign g6315 = (g3849&g6194);
assign g5886 = ((~g5753));
assign g2565 = ((~I3675));
assign I4210 = ((~g2294))|((~g804));
assign g5014 = (g4785)|(g4583);
assign g3940 = ((~I5177));
assign g2518 = ((~I3644));
assign g4719 = ((~I6337));
assign I7563 = ((~g74))|((~I7562));
assign g6342 = (g6264&g6076);
assign I8878 = ((~g6710));
assign I3412 = ((~g1419))|((~I3411));
assign I2057 = ((~g685));
assign g3484 = (g349&g2958);
assign g5550 = ((~g5331));
assign g5090 = ((~g4741));
assign g5482 = (g370&g5331);
assign I5502 = ((~g3853));
assign g3230 = ((~I4489));
assign g6784 = ((~I8940));
assign I4160 = ((~g2015))|((~I4159));
assign I3155 = ((~g1612));
assign I2768 = ((~g743))|((~I2766));
assign g5569 = (g5348&g3772);
assign g2932 = ((~g1998));
assign g3942 = (g3215)|(g3575);
assign g2909 = (g606&g2092);
assign g4447 = (g4384)|(g4044);
assign g3967 = ((~I5223));
assign I2814 = ((~g1222));
assign g4038 = (g430&g3388);
assign I3608 = ((~g1461));
assign I5226 = ((~g3259))|((~g3263));
assign I9050 = ((~g6832))|((~g3598));
assign g1725 = ((~g1113));
assign g944 = ((~I2004))|((~I2005));
assign g3520 = ((~g3183))|((~g3002))|((~g2197))|((~g2968));
assign g4039 = (g402&g3388);
assign g3224 = ((~I4471));
assign g4766 = ((~I6406));
assign g6443 = ((~g6385)&(~g4334)&(~g4092)&(~g4080));
assign g1543 = ((~g1006));
assign g5428 = (g394&g5300);
assign g1681 = ((~I2663));
assign g1323 = ((~I2324));
assign g949 = ((~g79));
assign g6165 = ((~g5926));
assign g6911 = (g6904&g6902);
assign I5472 = ((~g3846));
assign I8034 = ((~g6242));
assign g4040 = ((~I5343));
assign I4498 = ((~g2686));
assign g3978 = (g3655)|(g3117);
assign g6582 = ((~I8614));
assign g1513 = ((~g878));
assign g6265 = (g520&g5903);
assign g4133 = ((~I5481));
assign g6432 = ((~g6376)&(~g4086)&(~g4309)&(~g4068));
assign g4739 = (g2850&g4579);
assign g6904 = ((~I9179));
assign g5917 = ((~I7683));
assign I3883 = ((~g2574));
assign g3063 = ((~I4288));
assign g4113 = ((~I5421));
assign I2604 = ((~g1222));
assign g2820 = ((~g2470));
assign g1858 = ((~I2964));
assign g2634 = ((~I3776));
assign g5466 = ((~I7146));
assign I3733 = ((~g2031));
assign I5899 = ((~g3748));
assign g1624 = ((~I2581));
assign g4339 = (g3971&g3289);
assign I5626 = ((~g3914));
assign g1608 = ((~I2570));
assign g6359 = ((~I8135)&(~I8136)&(~I8137)&(~I8138));
assign I3915 = ((~g287))|((~I3914));
assign g3898 = ((~g3575));
assign I6930 = ((~g5017));
assign g6560 = ((~I8564));
assign I3923 = ((~g2581));
assign g5116 = ((~g4810));
assign g5952 = (g5120&g5809);
assign g4588 = (g2419&g4273);
assign g1037 = ((~I2067));
assign I6045 = ((~g4375));
assign I1970 = ((~g516))|((~I1969));
assign I2688 = ((~g1030));
assign I2929 = ((~g1659));
assign g2176 = ((~I3319));
assign I6697 = ((~g4722));
assign I3288 = ((~g1710));
assign g1890 = ((~g1359));
assign g4141 = ((~I5505));
assign g3167 = (g1883&g921);
assign g1670 = ((~I2648));
assign g5878 = ((~I7646));
assign I8168 = ((~g6170));
assign g3787 = ((~I4986));
assign g2890 = ((~g1875));
assign I2731 = ((~g1117));
assign I3240 = ((~g1460));
assign I7475 = ((~g5627));
assign g4050 = (I5359&I5360);
assign g3981 = (g3661)|(g3123);
assign g6598 = ((~I8662));
assign g3790 = ((~g3388));
assign g6875 = ((~I9092));
assign I9059 = (g5185)|(g5198)|(g6279);
assign g3855 = (g3626)|(g3631);
assign g3284 = ((~g3019));
assign I3496 = ((~g1326));
assign g1542 = ((~g878));
assign g1056 = ((~g89));
assign g1633 = (g716&g152);
assign g6625 = (g2121&g1595&g6538);
assign g3330 = ((~g1815))|((~g1797))|((~g3109));
assign I5457 = ((~g3766));
assign I8773 = (g6610)|(g6608)|(g6606)|(g6604);
assign g3483 = ((~g2716));
assign g3955 = ((~I5188))|((~I5189));
assign g1253 = ((~I2245))|((~I2246));
assign g1588 = ((~g798));
assign I9107 = ((~g6855));
assign g3745 = (g3356)|(g2770);
assign I4161 = ((~g619))|((~I4159));
assign g6341 = (g6261&g6074);
assign g2108 = ((~I3232));
assign I7529 = ((~g5662))|((~I7527));
assign g5740 = ((~I7501));
assign I1927 = ((~g665));
assign g2010 = ((~g1473))|((~g1470))|((~g1459));
assign I2296 = ((~g893));
assign I5857 = ((~g3740));
assign g6840 = ((~I9041));
assign g6608 = ((~I8690));
assign g5299 = ((~I6949));
assign g872 = ((~g143));
assign g4183 = (g3965&g1391);
assign g6566 = ((~I8582));
assign g1761 = ((~I2788));
assign g2583 = ((~g1830));
assign g2922 = ((~g1960));
assign I6576 = ((~g4700));
assign I7960 = ((~g5925));
assign I8843 = ((~g6658));
assign I7996 = ((~g6137));
assign I6327 = ((~g4451));
assign g1113 = ((~I2147));
assign g5095 = (g4794&g951);
assign g5677 = (g69&g5575);
assign I5030 = ((~g3242));
assign g4346 = (g157&g3773);
assign g6274 = (g5682)|(g5956);
assign I2301 = ((~g341))|((~I2299));
assign I5409 = ((~g3980));
assign g3325 = (g224&g2876);
assign g6247 = (g504&g5893);
assign g2836 = ((~g2509));
assign I7035 = ((~g5150));
assign g2902 = ((~g1899));
assign I6337 = ((~g4455));
assign g6728 = ((~I8878));
assign g926 = ((~I1952))|((~I1953));
assign I8358 = (g5192)|(g5153)|(g5158)|(g5197);
assign g2958 = ((~g1861));
assign I7564 = ((~g5676))|((~I7562));
assign g4834 = (g4534&g4531);
assign g1791 = ((~I2845));
assign I3909 = ((~g2044));
assign g3906 = ((~g3575));
assign g1461 = ((~I2460));
assign g3889 = ((~g3575));
assign g2364 = ((~I3516));
assign I8103 = ((~g6134));
assign g5378 = (g179&g5260);
assign g1975 = ((~I3086));
assign g5182 = (g520&g4993);
assign g5731 = ((~g952)&(~g5688));
assign g6816 = (g6784&g3346);
assign g3558 = (g338&g3199);
assign I8136 = (g6015)|(g6212)|(g4950)|(g4877);
assign I6672 = ((~g4752));
assign g2746 = (g2473&g1954);
assign g2390 = ((~I3531));
assign g3589 = ((~g3094));
assign g6128 = (g5590&g5958);
assign g6283 = ((~I7999));
assign g2581 = ((~I3694));
assign I8118 = (g6015)|(g6212)|(g4950)|(g4877);
assign I7119 = ((~g5303));
assign I6042 = ((~g4374));
assign g3353 = (g3162&g2921);
assign g2678 = ((~g2312));
assign g2603 = ((~I3733));
assign g6640 = (g1612&g6549);
assign g3530 = ((~g3204))|((~g3023))|((~g2197))|((~g2179));
assign g4490 = (g2941&g4210);
assign g3479 = (g345&g2957);
assign g3037 = ((~I4252));
assign g4499 = ((~I6015));
assign I3811 = ((~g2145));
assign g2940 = ((~g197))|((~g2381));
assign g3246 = ((~I4527))|((~I4528));
assign g6794 = (g6777)|(g3333);
assign g2032 = ((~g1749));
assign g4686 = (g4590&g1348);
assign g3865 = (g3637)|(g3648);
assign g4850 = ((~I6558));
assign I4474 = ((~g3052));
assign I7270 = ((~g5352));
assign g6052 = ((~g5824));
assign g3860 = ((~I5081));
assign g5495 = (g5444&g3456);
assign g3849 = (g3618)|(g3625);
assign g5697 = (g5646)|(g5485);
assign g5324 = ((~g5069)&(~g4410)&(~g766));
assign I3635 = ((~g1305));
assign g6832 = ((~I9021));
assign g6498 = ((~I8414));
assign I5059 = ((~g3259));
assign g4272 = ((~g3767)&(~g3319));
assign g5577 = ((~g5420));
assign I2275 = ((~g909));
assign g4525 = ((~I6087));
assign I6607 = ((~g4745));
assign g4152 = ((~I5542));
assign g2883 = ((~g1954));
assign g4107 = ((~I5403));
assign I3408 = ((~g1644));
assign g1419 = (g613&g918);
assign g5065 = (g4667)|(g4671);
assign g2004 = ((~I3115));
assign I2643 = ((~g965));
assign g2706 = ((~I3861));
assign g2575 = ((~I3684));
assign g4638 = (g4345)|(g3620);
assign g4118 = ((~I5436));
assign g3074 = ((~I4303));
assign g6527 = ((~I8497));
assign g5189 = (g528&g4993);
assign I5600 = ((~g3821));
assign g2806 = ((~g2446));
assign g4041 = (g461&g3388);
assign g3802 = ((~g3388));
assign g5818 = ((~g5638))|((~g2056))|((~g1666))|((~g1661));
assign g1563 = ((~g1006));
assign g1422 = ((~g1039)&(~g913));
assign g4671 = (g4645&g4641);
assign I8567 = ((~g6432));
assign g2056 = (g1672&g1675);
assign I5217 = ((~g3673));
assign g3693 = (g2256&g2830);
assign g1315 = ((~I2296));
assign g5922 = ((~I7698));
assign I4234 = ((~g2267))|((~I4233));
assign g6091 = (g1161&g5753);
assign g3158 = ((~I4398));
assign I9161 = ((~g6880));
assign I4303 = ((~g1897));
assign I3687 = ((~g1814));
assign I5187 = ((~g3589))|((~g3593));
assign g4827 = (g4520&g4515);
assign I2185 = ((~g29));
assign g4640 = ((~g4402))|((~g1056));
assign I2955 = ((~g1729));
assign g3362 = (g3031&g2740);
assign g3642 = (g3054&g2754);
assign I5343 = ((~g3599));
assign I2528 = ((~g719))|((~I2526));
assign g5442 = ((~g5270));
assign g6296 = (g6247)|(g6088);
assign I4522 = ((~g2801));
assign I4233 = ((~g2267))|((~g798));
assign I8414 = ((~g6418));
assign I3546 = ((~g1586));
assign g6774 = ((~g6754))|((~g6750));
assign g3878 = (g3703)|(g3191);
assign g1661 = ((~g1076));
assign g2757 = ((~I3934))|((~I3935));
assign I8687 = ((~g6568));
assign I4312 = ((~g2555));
assign g6846 = (g5860)|(g6834);
assign I7208 = ((~g143))|((~g5367));
assign I6247 = ((~g4609));
assign I8503 = ((~g6434));
assign g1006 = ((~I2047));
assign g6778 = ((~g6762))|((~g6758));
assign g3758 = (g545&g3461);
assign g2945 = ((~I4133));
assign g6137 = ((~I7859));
assign I4783 = ((~g2846))|((~I4782));
assign I6448 = ((~g4626));
assign g6347 = ((~I8103));
assign I3274 = ((~g1773));
assign g6289 = (g6240)|(g6081);
assign g6895 = ((~I9152));
assign g2311 = ((~I3456))|((~I3457));
assign I6745 = ((~g582))|((~I6743));
assign g1337 = ((~I2364));
assign g4232 = ((~I5674));
assign g6583 = ((~I8617));
assign g6485 = (I8393)|(I8394)|(I8395);
assign g6412 = ((~I8246));
assign I5562 = ((~g4002));
assign I4777 = ((~g2962));
assign g6385 = ((~g6271));
assign g6591 = ((~I8641));
assign g845 = ((~g582));
assign g3308 = ((~g3060));
assign g6182 = (g6047)|(g6034);
assign g5954 = (g5121&g5813);
assign g3705 = ((~g3014));
assign g6414 = ((~I8252));
assign g6332 = ((~I8074));
assign g5314 = ((~I6972));
assign g3346 = ((~I4623));
assign g1954 = ((~I3065));
assign g4022 = ((~I5328));
assign g3207 = ((~I4445))|((~I4446));
assign g3775 = ((~g3388));
assign g1644 = ((~I2611));
assign g3844 = (g3540&g1665);
assign I4791 = ((~g2814));
assign I8447 = ((~g6410));
assign I3537 = ((~g1305));
assign I7110 = ((~g5291));
assign g3763 = (g3064&g3501);
assign I6937 = ((~g5124));
assign g5155 = ((~g5099));
assign I3310 = ((~g1640));
assign g4713 = ((~I6321));
assign I2802 = ((~g1204));
assign g784 = ((~I1862));
assign I8345 = (g6326)|(g6135)|(g6140)|(g6157);
assign g3183 = ((~I4420));
assign g5145 = (g175&g5099);
assign g4707 = ((~I6311));
assign g4362 = (g3996&g3355);
assign g5659 = (g5551)|(g5398);
assign I2544 = ((~g774))|((~I2542));
assign g4410 = (g3903&g1474);
assign g6232 = ((~g6048));
assign I8994 = ((~g6789));
assign I5551 = ((~g4059));
assign g5559 = (g5024&g5453);
assign g1550 = ((~g996));
assign g6145 = (g3187&g6015);
assign g3258 = ((~I4537));
assign g3935 = (g3464)|(g2868);
assign g4465 = ((~g319))|((~g4253));
assign g791 = ((~I1865));
assign g5664 = ((~g5521));
assign g6122 = ((~I7838));
assign g4164 = (g3958&g2091);
assign g3723 = ((~I4903));
assign g5388 = (g5318)|(g1589)|(g3491);
assign g3358 = (g2842&g1369);
assign I8061 = ((~g6113));
assign I5674 = ((~g4003));
assign g4861 = ((~I6587));
assign g3486 = ((~g2869));
assign g6132 = (g3752&g5880);
assign g5163 = (g402&g4950);
assign g5474 = (g5363)|(g5146);
assign g901 = ((~g314))|((~g310));
assign g3171 = (g248&g2488);
assign g3296 = (g3054&g2650);
assign g5779 = ((~I7549))|((~I7550));
assign g2324 = ((~I3478));
assign I5223 = ((~g3537));
assign g4578 = ((~g4234)&(~g3928));
assign g3799 = ((~g3388));
assign g5852 = ((~g5638))|((~g2053))|((~g1661));
assign I2204 = ((~g694));
assign g3425 = (g2296&g3208);
assign I5736 = ((~g4022));
assign g3927 = ((~g3382)&(~g3383));
assign I4483 = ((~g3082));
assign g6397 = ((~I8202))|((~I8203));
assign g6689 = (g6266)|(g6648);
assign g5440 = ((~g5266));
assign g6733 = ((~I8891));
assign g4034 = ((~I5333));
assign g4377 = (g457&g3791);
assign I5731 = ((~g3942));
assign g6758 = (g6673)|(g6628)|(g6738);
assign g1209 = ((~I2215));
assign g1255 = ((~g161));
assign g6531 = ((~I8509));
assign g2316 = ((~I3468));
assign I8349 = (I8345)|(I8346)|(I8347)|(I8348);
assign I2080 = ((~g25))|((~g19));
assign g3719 = ((~g3053));
assign g3615 = (g2422&g3046);
assign g5212 = (g561&g5025);
assign g4645 = (g4352)|(g3633);
assign g4193 = ((~I5609));
assign I6621 = ((~g4745));
assign I8282 = ((~g6309));
assign I5490 = ((~g3832));
assign I3767 = ((~g2125));
assign I5904 = ((~g3749));
assign g3796 = ((~g3388));
assign I7522 = ((~g5659))|((~I7520));
assign g908 = ((~I1932));
assign I1958 = ((~g702));
assign g4245 = ((~g3759)&(~g3288));
assign g3537 = ((~I4757));
assign g4653 = (g4361)|(g3652);
assign I4547 = ((~g353))|((~I4545));
assign g1378 = ((~I2414));
assign g2339 = (g1603&g197);
assign g6306 = ((~I8030));
assign g2872 = ((~g1922));
assign g4498 = ((~I6012));
assign g878 = ((~g639));
assign g743 = ((~I1844));
assign g6709 = ((~I8837));
assign I6769 = ((~g4786));
assign g3996 = (g3691)|(g3171);
assign g4015 = (g445&g3388);
assign g3519 = ((~g2740));
assign I3349 = ((~g1334));
assign g2506 = ((~I3632));
assign I6302 = ((~g4440));
assign g2350 = ((~I3502));
assign I2864 = ((~g1177));
assign g6580 = ((~g6491));
assign g3360 = (g2783&g1947);
assign g6154 = (g3219&g6015);
assign g4794 = (g4593&g949);
assign I2935 = ((~g345))|((~I2933));
assign g2255 = (g1706&g736);
assign g6081 = (g1177&g5731);
assign g4191 = ((~I5603));
assign I4528 = ((~g646))|((~I4526));
assign I9155 = ((~g6882));
assign I2578 = ((~g1209));
assign I5204 = ((~g3534));
assign g6474 = (g2138&g2036&g6397);
assign I8603 = ((~g6449));
assign g5578 = ((~g5425));
assign I6111 = ((~g4404));
assign g5064 = ((~I6706));
assign I8450 = ((~g6412));
assign I2237 = ((~g465));
assign g5174 = ((~g5099));
assign I2658 = ((~g1001));
assign g1174 = ((~g37));
assign I7216 = ((~g152))|((~g5368));
assign g5866 = ((~g5649))|((~g1529))|((~g2081));
assign g4655 = (g4368)|(g3660);
assign I6194 = ((~g4199))|((~g631));
assign I9057 = (g6320)|(g6828)|(g6830)|(g6153);
assign g1287 = ((~g855));
assign g6826 = ((~I9011));
assign I7451 = ((~g5597));
assign g6370 = ((~I8174));
assign g1802 = (g89&g1064);
assign g3780 = (g3043&g3519);
assign g6348 = (g5869&g6211);
assign I5893 = ((~g3747));
assign I2907 = ((~g1498));
assign g6482 = (I8376)|(I8377)|(I8378)|(I8379);
assign g6318 = (g3865&g6212);
assign g1672 = ((~g1094));
assign g3564 = ((~g2618));
assign g6611 = ((~I8699));
assign g5598 = (g5046&g5509);
assign g4993 = ((~g4674)&(~g1477));
assign g6683 = (g6465)|(g6622)|(g6621);
assign g4463 = ((~g4364));
assign g6337 = ((~I8089));
assign g1473 = ((~g944)&(~g941)&(~g939));
assign I2394 = ((~g719));
assign I4184 = ((~g749))|((~I4182));
assign g4691 = (g4581&g2098);
assign g3691 = (g2268&g2828);
assign g3776 = ((~g3466));
assign I7484 = ((~g5630));
assign I4170 = ((~g2157));
assign g4148 = ((~I5526));
assign g1735 = ((~I2745));
assign g4101 = ((~I5385));
assign I8395 = (g5182)|(g5200)|(g6280);
assign I5848 = ((~g3856));
assign g4541 = (g631&g4199);
assign I3077 = ((~g1439));
assign I7318 = ((~g5452));
assign g1793 = ((~g94))|((~g1084));
assign g5700 = (g5663)|(g5488);
assign g3041 = ((~I4258));
assign I1935 = ((~g666));
assign g6912 = (g6899&g6897);
assign g4262 = ((~I5713));
assign I6175 = ((~g4236))|((~g571));
assign g5121 = ((~I6775));
assign g6515 = ((~g6408));
assign g1636 = ((~I2593));
assign g6442 = ((~g6376)&(~g4323)&(~g4074)&(~g4302));
assign I4309 = ((~g2525));
assign I6343 = ((~g4458));
assign I2842 = ((~g1177));
assign g2007 = ((~g1411));
assign g6880 = ((~I9107));
assign I5923 = ((~g4299));
assign g2807 = (g2568&g2001);
assign g3373 = (g3118&g2927);
assign g3057 = ((~I4282));
assign g6425 = ((~I8285));
assign g5561 = ((~g5391)&(~g1589)&(~g3793)&(~g1880));
assign g4003 = ((~g3441));
assign g6088 = (g1143&g5753);
assign g4504 = ((~I6027))|((~I6028));
assign g951 = ((~g84));
assign g5437 = ((~I7119));
assign I4671 = ((~g2928));
assign I3519 = ((~g1305));
assign g5671 = (g54&g5572);
assign g6854 = ((~I9085));
assign g910 = ((~I1938));
assign I3847 = ((~g284))|((~I3846));
assign g4762 = ((~I6391))|((~I6392));
assign I8210 = (g5202)|(g4993)|(g4967)|(g4980);
assign g1270 = ((~g844));
assign g3797 = ((~g3388));
assign g4928 = (g148&g4723);
assign g5481 = (g366&g5331);
assign I3946 = ((~g2256));
assign g2861 = (g2120&g1654);
assign g2021 = (g835&g1436);
assign g3086 = ((~I4327));
assign I2779 = ((~g1038));
assign I3578 = ((~g1484));
assign I2424 = ((~g719));
assign I3090 = ((~g1504));
assign g6724 = ((~I8866));
assign I8966 = ((~g6796));
assign I3749 = ((~g2484));
assign g4687 = (g4493&g1542);
assign g3450 = ((~I4688));
assign I5868 = ((~g3864));
assign I4980 = ((~g3546));
assign g6073 = ((~g197)&(~g5862));
assign g3988 = (g3678)|(g3143);
assign g3337 = (g2796&g2913);
assign g4785 = (g2160&g4625);
assign I4504 = ((~g2726));
assign g1533 = ((~g878));
assign I2388 = ((~g878));
assign g6750 = (g6670)|(g6625)|(g6736);
assign g6927 = (g6799)|(g6924);
assign g2996 = ((~I4189));
assign I6090 = ((~g4393));
assign I6001 = ((~g4162));
assign g4632 = ((~g4281));
assign g5751 = ((~I7506));
assign I9104 = ((~g6864));
assign g6647 = (g6578&g6233);
assign g6787 = (g3758)|(g6766);
assign g3877 = (g3651)|(g3659);
assign g706 = ((~I1825));
assign g5903 = ((~g5753));
assign I5535 = ((~g3907))|((~g654));
assign I4010 = ((~g2568))|((~I4008));
assign I1953 = ((~g248))|((~I1951));
assign g5566 = ((~I7318));
assign g5169 = (g5093&g1375);
assign I6885 = ((~g4872));
assign g3677 = ((~g3140));
assign I5445 = ((~g4040));
assign g4172 = (g3930&g1366);
assign g6694 = ((~I8800));
assign g6850 = ((~I9077));
assign g1647 = ((~I2620));
assign g2946 = ((~g2296));
assign g4286 = ((~I5743));
assign g6576 = ((~g6487));
assign I8329 = ((~g6305));
assign I5825 = ((~g3914));
assign I8040 = ((~g6142));
assign g5382 = ((~I7042));
assign I3826 = ((~g2145));
assign I3531 = ((~g1593));
assign g2903 = ((~g1902));
assign I4318 = ((~g2171));
assign g3350 = (g3150&g1928);
assign I8129 = (g4915)|(g5025);
assign g3814 = (g913&g3546);
assign I8716 = ((~g6518));
assign g4486 = (g716&g4195);
assign g2814 = ((~I4023));
assign g6407 = ((~I8235));
assign g2467 = ((~I3599));
assign I3445 = ((~g1689))|((~g729));
assign I6552 = ((~g4702));
assign g1742 = ((~I2756));
assign g5887 = ((~g5742));
assign I2021 = ((~g528))|((~g254));
assign g5571 = ((~g5395));
assign g6166 = ((~I7892));
assign I7077 = ((~g5281));
assign g3424 = ((~I4671));
assign g3521 = ((~g3187))|((~g3023))|((~g3007))|((~g2179));
assign g6039 = ((~g5824));
assign I5415 = ((~g3723));
assign I3251 = ((~g1471));
assign g5118 = ((~I6766));
assign g4568 = ((~g4233)&(~g3924));
assign g6906 = ((~I9185));
assign I5244 = ((~g3247))|((~I5242));
assign I3840 = ((~g2125));
assign g4270 = ((~I5723));
assign I4362 = ((~g2555));
assign g1232 = ((~I2228));
assign g4185 = (g398&g3906);
assign g2877 = ((~g2434));
assign g6783 = ((~g6747))|((~g5068))|((~g5066));
assign g4440 = (g4371)|(g4038);
assign I4152 = ((~g139))|((~I4150));
assign g6665 = (I8778)|(I8779);
assign g3140 = ((~g2409))|((~g1060))|((~g1620));
assign I8803 = ((~g6685));
assign g6834 = ((~g6821));
assign g838 = ((~g564));
assign g6188 = ((~g5950));
assign g3657 = (g2734&g2357);
assign g6801 = ((~I8969));
assign g4872 = (g4760&g1549);
assign I5478 = ((~g3859));
assign g5162 = (g5088&g2105);
assign g4858 = ((~I6582));
assign g3752 = ((~I4935));
assign g2914 = ((~g1928));
assign I1838 = ((~g206));
assign g2986 = ((~g2010));
assign I6324 = ((~g4450));
assign g3528 = ((~g1802)&(~g3167));
assign g1558 = ((~I2527))|((~I2528));
assign g5410 = (g378&g5274);
assign g5817 = (g5380)|(g5621);
assign I6743 = ((~g4708))|((~g582));
assign g3868 = ((~g3491));
assign g5532 = (g5350)|(g3278);
assign g1994 = ((~I3105));
assign I3599 = ((~g1484));
assign I8080 = (g6015)|(g6212)|(g4950)|(g4877);
assign g3511 = ((~g3158))|((~g3002))|((~g2976))|((~g2968));
assign g2804 = ((~I4009))|((~I4010));
assign I7981 = (g4915)|(g5025);
assign I5871 = ((~g3744));
assign g4582 = ((~g4210));
assign g2291 = ((~I3434));
assign I2584 = ((~g839));
assign g6105 = ((~I7811));
assign g4771 = ((~I6417));
assign g4577 = ((~g4202));
assign g5398 = (g366&g5261);
assign g4801 = ((~g4487));
assign g6251 = (g5668)|(g5939);
assign g943 = ((~g496));
assign g3941 = (g3479)|(g2873);
assign I7497 = ((~g5687));
assign g5225 = (g669&g5054);
assign g6487 = ((~g6365));
assign I8831 = ((~g6665));
assign g3113 = (g224&g2364);
assign g4086 = (g3310)|(g2720);
assign I4249 = ((~g2525));
assign g2731 = ((~I3894))|((~I3895));
assign g2234 = ((~I3367));
assign I4391 = ((~g2275));
assign g1680 = ((~g1011));
assign g1541 = ((~g1094));
assign g6732 = ((~I8888));
assign g716 = ((~I1832));
assign I8070 = ((~g6116));
assign I5270 = ((~g3705))|((~I5269));
assign g3968 = ((~I5227))|((~I5228));
assign g2121 = (g1632&g754);
assign g6843 = ((~I9051))|((~I9052));
assign g3688 = (g2783&g2457);
assign g6448 = ((~g6376)&(~g4323)&(~g4309)&(~g4302));
assign g2347 = ((~I3499));
assign g1049 = ((~g266));
assign g3282 = (g131&g2863);
assign I5879 = ((~g3745));
assign I7434 = ((~g5554))|((~I7432));
assign g2896 = (g2323)|(g1763);
assign g4765 = ((~I6403));
assign g3597 = ((~I4783))|((~I4784));
assign I6772 = ((~g4788));
assign g2716 = ((~I3871));
assign I8113 = ((~g6147));
assign I3830 = ((~g2179));
assign g4516 = ((~I6060));
assign g5508 = ((~I7245))|((~I7246));
assign g3870 = (g3700)|(g3182);
assign g4425 = ((~I5926));
assign I2817 = ((~g1222));
assign g5620 = (g5507&g4938);
assign g3271 = ((~g3042));
assign I5606 = ((~g3821));
assign I3871 = ((~g2145));
assign g3231 = ((~I4492));
assign g5742 = ((~g5686));
assign g3698 = (g2284&g2835);
assign g5502 = ((~I7209))|((~I7210));
assign g3247 = ((~g2973));
assign I6069 = ((~g4213));
assign I5124 = ((~g3719));
assign I2169 = ((~g269));
assign g4590 = ((~g4169)&(~g4172));
assign I6026 = ((~g4223))|((~g4221));
assign I2795 = ((~g804))|((~g798));
assign I5463 = ((~g3783));
assign g5705 = ((~I7466));
assign I2246 = ((~g598))|((~I2244));
assign g5808 = (g5373)|(g5616);
assign g3850 = (g3680)|(g3145);
assign I7704 = ((~g5723));
assign I7506 = ((~g5584));
assign I8972 = ((~g6795));
assign g5091 = ((~g4698)&(~g4701));
assign g6323 = (g3877&g6194);
assign g1279 = ((~g848));
assign g2745 = ((~I3915))|((~I3916));
assign g6573 = ((~I8603));
assign g3319 = (g2688&g2675);
assign g3664 = ((~g2804)&(~g2791)&(~g2780));
assign g4530 = ((~I6102));
assign g3635 = (g2473&g3079);
assign I2234 = ((~g697));
assign g3500 = ((~g2647));
assign I3861 = ((~g1834));
assign g2967 = ((~I4166));
assign g6134 = ((~I7852));
assign g2849 = ((~g2577));
assign I7061 = ((~g5281));
assign I1877 = ((~g283));
assign I7244 = ((~g188))|((~g5377));
assign g5249 = ((~g4868)&(~g4870));
assign g5800 = (g5369)|(g5600);
assign g2643 = ((~I3785));
assign g2792 = ((~g2416));
assign g4593 = (g4277&g947);
assign g5479 = ((~I7173));
assign g3235 = ((~I4504));
assign g4533 = ((~I6111));
assign g6919 = (g6912)|(g6914);
assign g4351 = (g166&g3776);
assign I7969 = (g6194)|(g5958)|(g5975)|(g5997);
assign g1775 = ((~g952));
assign g6430 = ((~g6385)&(~g3733)&(~g4092)&(~g4080));
assign I4519 = ((~g2788));
assign g1689 = (g766&g719);
assign I2175 = ((~g25));
assign g4520 = ((~I6072));
assign g5402 = (g370&g5266);
assign g2422 = ((~I3560));
assign I3134 = ((~g1336));
assign g3147 = (g2419&g59);
assign g4163 = (g374&g3892);
assign g1789 = ((~I2839));
assign g6557 = (g1595&g6469);
assign I5300 = ((~g471))|((~g3505));
assign g4627 = (g4333)|(g3603);
assign g2584 = ((~I3705));
assign I3572 = ((~g1295));
assign I2300 = ((~g830))|((~I2299));
assign g2772 = ((~I3961));
assign g6275 = (g1735&g6070);
assign g5683 = ((~I7433))|((~I7434));
assign g1815 = ((~g102))|((~g1070));
assign g3744 = (g3345)|(g2759);
assign g2974 = ((~I4173));
assign g6584 = ((~I8620));
assign g4950 = ((~g1472)&(~g4680));
assign g4348 = (g3987&g3322);
assign g3934 = ((~g3377)&(~g3379));
assign g1114 = ((~I2150));
assign I8470 = ((~g6461));
assign g6503 = ((~I8429));
assign g1790 = ((~I2842));
assign g1585 = (g1017&g1011);
assign I6392 = ((~g4610))|((~I6390));
assign g3887 = (g3276&g1861);
assign g923 = ((~g332));
assign I8699 = ((~g6573));
assign g6106 = ((~I7814));
assign g5323 = (g5098)|(g4802);
assign I2379 = ((~g1123));
assign g6326 = (g3833&g6194);
assign g5663 = (g4513&g5550);
assign g1732 = ((~I2738));
assign g6793 = (g6771)|(g3323);
assign I7231 = ((~g170))|((~I7230));
assign g4936 = (g4827)|(g4828);
assign g1919 = ((~I3022));
assign g4251 = ((~I5705));
assign g2582 = ((~I3698))|((~I3699));
assign I9058 = (g6156)|(g6331)|(g5190)|(g5164);
assign I3001 = ((~g1267));
assign g1760 = ((~I2785));
assign g3557 = ((~g2598));
assign g6637 = (g1842&g6549);
assign g6272 = (g5679)|(g5953);
assign I5269 = ((~g3705))|((~g3710));
assign I8538 = ((~g6450));
assign I2767 = ((~g749))|((~I2766));
assign g4831 = (g4528&g4524);
assign g4780 = ((~I6434));
assign g1716 = (g821&g774&g784);
assign g4727 = ((~I6355));
assign g3977 = (g3653)|(g3113);
assign g4487 = ((~I5991));
assign I2272 = ((~g908));
assign g5496 = (g5446&g3457);
assign g5046 = ((~I6680));
assign I6537 = ((~g4711));
assign I6952 = ((~g5124));
assign I3785 = ((~g2346));
assign g3689 = (g3162&g2826);
assign I5040 = ((~g3271));
assign g6282 = ((~I7996));
assign g3531 = ((~g3209))|((~g2215))|((~g2976))|((~g2179));
assign g6727 = ((~I8875));
assign I7517 = ((~g5593));
assign g2957 = ((~g1861));
assign I4282 = ((~g2525));
assign g909 = ((~I1935));
assign g4589 = ((~g4180)&(~g4183));
assign I7608 = ((~g5605));
assign g6920 = (g6915)|(g6916);
assign g6613 = (g932&g6554);
assign g6658 = (g6132)|(g6620);
assign I3726 = ((~g2030));
assign g1824 = ((~I2890));
assign g6051 = ((~g5824));
assign I4477 = ((~g3063));
assign I3773 = ((~g2524));
assign g5213 = (g4862&g5087);
assign g2035 = ((~I3144));
assign g2336 = ((~I3488));
assign g1320 = ((~I2315));
assign I2370 = ((~g1123));
assign g3225 = ((~I4474));
assign I2140 = ((~g28));
assign I6244 = ((~g4519));
assign g6932 = ((~I9217));
assign I2526 = ((~g766))|((~g719));
assign I7637 = ((~g5751));
assign g1418 = ((~g486)&(~g943));
assign g2107 = (g1583&g1543);
assign g5415 = ((~I7081));
assign g3604 = ((~I4799));
assign g4184 = (g3934&g2136);
assign g5567 = ((~g5418));
assign g5325 = ((~g5077)&(~g4416)&(~g821));
assign g866 = ((~g314));
assign g1539 = ((~g878));
assign I2476 = ((~g971));
assign g3170 = (g254&g2485);
assign g6433 = ((~g6385)&(~g3733)&(~g4092)&(~g4314));
assign g6559 = (g1612&g6474);
assign g3897 = ((~g3251));
assign g1756 = ((~I2779));
assign g6565 = ((~I8579));
assign I5523 = ((~g3840));
assign I7295 = ((~g5439));
assign g4383 = (g453&g3796);
assign g3099 = (g218&g2350);
assign g5879 = ((~g5770));
assign I2919 = ((~g1787));
assign g5115 = ((~I6759));
assign I3914 = ((~g287))|((~g2449));
assign g5399 = ((~I7065));
assign g3166 = (g2042&g1233);
assign g4718 = ((~I6334));
assign I3232 = ((~g1782));
assign g839 = ((~g567));
assign g4293 = ((~I5750));
assign g3064 = ((~I4291));
assign g5458 = (g3466)|(g5311);
assign I6927 = ((~g5124));
assign g5465 = ((~I7143));
assign g2097 = ((~I3215));
assign I5929 = ((~g4152));
assign g2698 = ((~I3847))|((~I3848));
assign g2576 = ((~I3687));
assign I2445 = ((~g971));
assign I9002 = ((~g6802));
assign g855 = ((~g650));
assign g4159 = (g370&g3890);
assign g6266 = (g1721&g6057);
assign I8991 = ((~g6788));
assign g3747 = (g3365)|(g2781);
assign I9113 = ((~g6855));
assign g2622 = ((~I3764));
assign g2691 = ((~g2317));
assign g6264 = (g5675)|(g5948);
assign g1499 = (g1101&g1094);
assign g5921 = ((~I7695));
assign g3363 = ((~g3110));
assign g3285 = (g2195&g2653);
assign g5686 = ((~g5546))|((~g1017))|((~g1551))|((~g2916));
assign g3544 = ((~g2594))|((~g2215))|((~g2197))|((~g2179));
assign g2100 = ((~g1588))|((~g804))|((~g791));
assign g3954 = (g3484)|(g3489);
assign I3127 = ((~g1276))|((~I3125));
assign g3880 = (g3658)|(g3665);
assign g4522 = ((~I6078));
assign g5558 = (g5018&g5450);
assign I1880 = ((~g276));
assign I4297 = ((~g2555));
assign g1055 = ((~g269));
assign g4400 = ((~I5899));
assign g4569 = ((~I6143));
assign g5307 = ((~I6959));
assign I5294 = ((~g625))|((~I5292));
assign g1878 = ((~I2973));
assign g6894 = ((~I9149));
assign g5669 = (g5556)|(g5410);
assign g3310 = (g224&g2871);
assign g2276 = ((~I3425));
assign I3474 = ((~g1450));
assign g5940 = (g5115&g5794);
assign I2668 = ((~g1011));
assign I3681 = ((~g1821));
assign g5273 = ((~I6930));
assign I2003 = ((~g500))|((~g212));
assign g6939 = ((~I9230));
assign g2170 = ((~I3301));
assign g4614 = ((~g4308));
assign g5918 = ((~I7686));
assign g4230 = (g3756&g1861);
assign I2162 = ((~g197));
assign g3487 = ((~g2622));
assign g2895 = ((~g1894));
assign g2195 = ((~I3334));
assign g1042 = ((~I2073))|((~I2074));
assign g5377 = (g5217)|(g4949);
assign g4654 = (g4362)|(g3654);
assign g1808 = (g706&g49);
assign I4706 = ((~g2877));
assign g3297 = ((~g3046));
assign g3527 = ((~I4743));
assign g4894 = ((~g4813));
assign I5469 = ((~g3838));
assign I3190 = ((~g791))|((~I3188));
assign g4370 = ((~I5831));
assign g5291 = (g5043)|(g4764);
assign g4138 = ((~I5496));
assign g1997 = ((~g1398));
assign g1336 = ((~I2361));
assign g3791 = ((~g3388));
assign g6233 = ((~g6052));
assign g6688 = (g6263)|(g6647);
assign g6497 = ((~I8411));
assign I3168 = ((~g1540))|((~g1534));
assign g5278 = ((~I6937));
assign g6131 = (g5593&g5975);
assign I3522 = ((~g1664));
assign I7701 = ((~g5720));
assign g1972 = ((~I3083));
assign g4864 = (g4744)|(g4490);
assign I6546 = ((~g4692));
assign g1363 = ((~I2399));
assign I1835 = ((~g205));
assign g6097 = ((~g2954))|((~g5857));
assign g4233 = (g3912)|(g471);
assign g4131 = ((~I5475));
assign I8969 = ((~g6797));
assign I8348 = (g5229)|(g5234)|(g5218)|(g5225);
assign g6121 = ((~I7835));
assign g4192 = ((~I5606));
assign g4244 = (g1749&g4004&g1609);
assign I3202 = ((~g1812));
assign g6823 = ((~I9002));
assign g3124 = ((~I4371));
assign g4106 = ((~I5400));
assign g5383 = ((~I7045));
assign g4352 = (g3988&g3331);
assign I2090 = ((~g33))|((~I2089));
assign I4480 = ((~g3073));
assign g3781 = ((~I4976));
assign g4122 = ((~I5448));
assign I3391 = ((~g1646));
assign g4704 = ((~I6302));
assign g5146 = (g184&g5099);
assign I2128 = ((~g18));
assign g5473 = (g5362)|(g5145);
assign g6193 = ((~g5957));
assign I2543 = ((~g821))|((~I2542));
assign g754 = ((~I1850));
assign I8866 = ((~g6701));
assign I4183 = ((~g2292))|((~I4182));
assign g5900 = (g5804&g5658);
assign g4391 = ((~I5876));
assign I4343 = ((~g2525));
assign g6062 = ((~g5824));
assign g6545 = (g6468)|(g4244);
assign I6359 = ((~g4566));
assign g6903 = ((~I9176));
assign g4347 = (g3986&g3320);
assign I2946 = ((~g1587));
assign I4794 = ((~g2814));
assign g2919 = ((~g1937));
assign g3762 = (g2672&g3500);
assign I9064 = (g6323)|(g6829)|(g6831)|(g6155);
assign g4646 = (g4353)|(g3635);
assign g1776 = ((~I2821));
assign I8668 = ((~g6530));
assign g5876 = ((~I7640));
assign g4119 = ((~I5439));
assign I8752 = ((~g6514));
assign I2060 = ((~g7))|((~g3));
assign g4774 = ((~g4442)&(~g4445));
assign g6740 = ((~g6703))|((~g6457))|((~g4936));
assign I2355 = ((~g1177));
assign I8623 = ((~g6542));
assign g5544 = ((~g5331));
assign g6092 = (g1123&g5731);
assign g2822 = ((~I4031));
assign g3387 = ((~I4664));
assign g3307 = (g2242&g2692);
assign g774 = ((~I1859));
assign I8600 = ((~g6451));
assign g2868 = (g1316&g1861);
assign g3073 = ((~I4300));
assign g6338 = (g6251&g6067);
assign g6590 = ((~I8638));
assign g6714 = ((~g6670));
assign g3632 = (g3043&g2743);
assign g4846 = ((~I6546));
assign I2041 = ((~g680));
assign g3692 = (g2268&g2829);
assign g3803 = ((~I5002));
assign I7555 = ((~g69))|((~g5674));
assign g5634 = ((~g5563))|((~g4767));
assign g714 = ((~g131));
assign g3323 = (g2253&g2716);
assign I9140 = ((~g6888));
assign g5893 = ((~g5753));
assign I5885 = ((~g3746));
assign I8117 = (g6194)|(g5958)|(g5975)|(g5997);
assign I4513 = ((~g2765));
assign I2623 = ((~g1161));
assign g4870 = (g4779&g1884);
assign I2281 = ((~g900));
assign g4455 = (g4396)|(g4052);
assign g2088 = ((~I3202));
assign I3325 = ((~g1340));
assign g1384 = ((~I2420));
assign g6297 = (g6248)|(g6089);
assign I9143 = ((~g6886));
assign g5355 = ((~I7007));
assign g6159 = (g3177&g6015);
assign g5447 = (g4545&g5256&g2311);
assign g3157 = (g2422&g2467);
assign g3083 = ((~I4318));
assign I1952 = ((~g524))|((~I1951));
assign I3388 = ((~g1324));
assign I8585 = ((~g6442));
assign g4672 = (g4635&g4631);
assign I5843 = ((~g3851));
assign g2443 = ((~I3578));
assign I5556 = ((~g4059));
assign g4692 = ((~I6280));
assign I5514 = ((~g3882));
assign g1691 = (g821&g774);
assign g5150 = ((~I6816));
assign g4828 = (g4510&g4508);
assign I7590 = ((~g5605));
assign I7311 = ((~g5364))|((~g590));
assign g5156 = (g434&g4877);
assign I8137 = (g4894)|(g4904)|(g4993)|(g4967);
assign I8828 = ((~g6661));
assign I3115 = ((~g1519));
assign g5370 = (g5211)|(g4937);
assign I8635 = ((~g6552));
assign g6069 = ((~g5791));
assign g6773 = (g6762&g2986);
assign g6908 = (g6907&g3886);
assign g3645 = (g2497&g3090);
assign g2092 = (g642&g1570);
assign g3786 = ((~g3388));
assign g4149 = ((~I5529));
assign I4821 = ((~g2877));
assign g6413 = ((~I8249));
assign I5840 = ((~g3732));
assign g889 = ((~g310));
assign g5631 = ((~g5536));
assign g6528 = ((~I8500));
assign I6756 = ((~g4775));
assign I7829 = ((~g5926));
assign I3428 = ((~g1825));
assign g1830 = ((~I2904));
assign I6959 = ((~g5089));
assign g6455 = (g6345)|(g5952);
assign I2361 = ((~g1075));
assign I2453 = ((~g952));
assign I7466 = ((~g5624));
assign I3481 = ((~g1461));
assign g5315 = ((~g5116));
assign g6525 = ((~I8491));
assign I1963 = ((~g242))|((~I1961));
assign g4910 = ((~I6612));
assign g6723 = ((~I8863));
assign I2193 = ((~g693));
assign I2756 = ((~g1175));
assign I4059 = ((~g1878));
assign I5376 = ((~g4014));
assign g1324 = ((~I2327));
assign g5082 = ((~g4723));
assign g3478 = ((~g2695));
assign g1632 = ((~g760));
assign g6445 = ((~g6376)&(~g4323)&(~g4309)&(~g4068));
assign g2640 = ((~I3782));
assign I5907 = ((~g3883));
assign g1755 = ((~I2776));
assign g4437 = ((~I5948));
assign g3846 = ((~I5053));
assign g6936 = (g5438)|(g6935);
assign g6257 = (g5671)|(g5941);
assign g4688 = (g1474&g4568);
assign g6921 = (g6908)|(g6816);
assign g4563 = ((~g4190));
assign g4252 = ((~I5708));
assign I8641 = ((~g6524));
assign g1472 = ((~g952));
assign g6249 = (g1332&g5892);
assign g6806 = ((~I8978));
assign I8217 = ((~g6319));
assign I2047 = ((~g682));
assign g1834 = ((~I2916));
assign I6488 = ((~g4603));
assign g1294 = ((~I2287));
assign g3501 = ((~g2650));
assign g1084 = ((~g98));
assign g3181 = (g254&g2509);
assign g1688 = ((~I2688));
assign g3648 = (g2722&g2343);
assign I7634 = ((~g5727));
assign I3593 = ((~g1295));
assign I6139 = ((~g4222));
assign g6510 = ((~I8450));
assign I6028 = ((~g4221))|((~I6026));
assign g4813 = ((~g4550))|((~g965))|((~g1560))|((~g2073));
assign g5600 = (g5502&g4900);
assign g1177 = ((~I2193));
assign g1391 = ((~I2424));
assign g5626 = (g5496)|(g3285);
assign g1551 = ((~g1011));
assign g4591 = ((~g4178)&(~g4181));
assign I5228 = ((~g3263))|((~I5226));
assign g4534 = ((~I6114));
assign I8186 = ((~g6179));
assign g3627 = (g2473&g3067);
assign I3509 = ((~g1461));
assign g3462 = ((~g2679));
assign g4519 = ((~I6069));
assign g6496 = ((~g952)&(~g6354));
assign g2795 = ((~g1997))|((~g866));
assign I9024 = ((~g6803));
assign I4688 = ((~g3207));
assign g1908 = ((~I3007));
assign I6989 = ((~g5307));
assign g5016 = (g4789)|(g4592);
assign g4741 = ((~I6371));
assign I6573 = ((~g4721));
assign I3761 = ((~g2505));
assign I4489 = ((~g2975));
assign I3499 = ((~g1450));
assign I5542 = ((~g3984));
assign g3240 = ((~I4519));
assign I7999 = ((~g6137));
assign g5092 = ((~g4753));
assign I1962 = ((~g520))|((~I1961));
assign g3344 = (g242&g2885);
assign g5403 = ((~I7069));
assign g6700 = ((~I8818));
assign g3146 = (g2370&g2446);
assign g6851 = (g6846&g2293);
assign g2966 = ((~I4160))|((~I4161));
assign g5385 = (g3992)|(g5318);
assign I4762 = ((~g2862));
assign g6897 = ((~I9158));
assign g5438 = (g5224&g3769);
assign g2817 = ((~g2461));
assign I3739 = ((~g2021))|((~g349));
assign g5137 = ((~I6789));
assign g5944 = (g5778&g5403);
assign g6237 = (g5912)|(g2381);
assign g6080 = ((~g5805));
assign g5359 = (g4428&g5155);
assign g5352 = ((~I7002));
assign g4345 = (g3982&g3308);
assign g1648 = ((~I2623));
assign I2887 = ((~g1123));
assign g4130 = ((~I5472));
assign I3602 = ((~g1491));
assign g6508 = ((~I8444));
assign g5507 = ((~I7238))|((~I7239));
assign I6986 = ((~g5230));
assign I8127 = (g6015)|(g6212)|(g4950)|(g4877);
assign g6317 = (g3862&g6194);
assign g3653 = (g2215&g2767);
assign g6615 = ((~I8707));
assign g1692 = ((~I2696));
assign g4271 = (g2121&g1749&g4004);
assign I2228 = ((~g15));
assign g4806 = ((~g4473));
assign I3902 = ((~g2576));
assign g6907 = (g6874)|(g3358);
assign I8812 = ((~g6688));
assign g2591 = ((~I3720));
assign g942 = ((~g69));
assign g3518 = ((~g3177))|((~g3023))|((~g3007))|((~g2981));
assign g6163 = ((~g5926));
assign g4036 = ((~I5337));
assign g3667 = (g2245&g2789);
assign g1070 = ((~g94));
assign g3617 = (g2609&g2317);
assign I2692 = ((~g1037));
assign I8385 = (g6316)|(g6128)|(g6131)|(g6149);
assign g2904 = ((~g1991));
assign g2470 = ((~I3602));
assign I2796 = ((~g804))|((~I2795));
assign g1763 = (g478&g1119);
assign I7284 = ((~g5383));
assign g3853 = ((~I5068));
assign I9125 = ((~g6855));
assign I3550 = ((~g1295));
assign I7225 = ((~g5370))|((~I7223));
assign I5766 = ((~g3961))|((~g3957));
assign I5475 = ((~g3852));
assign g5480 = ((~I7176));
assign g2041 = ((~I3152));
assign I7604 = ((~g5605));
assign g4768 = ((~I6410));
assign g5884 = ((~g5864));
assign g6603 = (g6581&g6236);
assign g6800 = ((~I8966));
assign g6087 = ((~g5813));
assign g2905 = ((~g1994));
assign g5423 = ((~g5170)&(~g5175));
assign g2062 = (g1499&g1666);
assign I2337 = ((~g1209));
assign g1295 = ((~I2290));
assign g1726 = ((~I2728));
assign I3543 = ((~g1461));
assign g4319 = ((~I5783))|((~I5784));
assign I2231 = ((~g465));
assign g3096 = ((~I4343));
assign g5161 = (g5095&g4535);
assign g5096 = (g4794&g4647);
assign g1549 = ((~g878));
assign g947 = ((~g74));
assign g4452 = (g3820&g4227);
assign g852 = ((~g634));
assign g6734 = ((~I8894));
assign I7892 = ((~g5916));
assign g3304 = (g2857&g1513);
assign g4694 = (g1481&g4578);
assign I6066 = ((~g4382));
assign g5214 = (g562&g5025);
assign g6737 = (g6714&g760&g5237);
assign g6782 = (g6719)|(g6749);
assign g1911 = ((~I3010));
assign g6036 = ((~g5824));
assign g5114 = ((~I6756));
assign I3178 = ((~g1706))|((~I3177));
assign I2182 = ((~g692));
assign g2231 = ((~I3358));
assign g6820 = ((~I8997));
assign g4375 = ((~I5840));
assign g1963 = ((~I3074));
assign g3788 = ((~g3466));
assign g5311 = (g5013&g4468);
assign I8840 = ((~g6657));
assign g4829 = (g4526&g4522);
assign g5816 = (g5378)|(g5620);
assign I2913 = ((~g1792));
assign g6917 = (g6909)|(g6910);
assign I2766 = ((~g749))|((~g743));
assign I6108 = ((~g4403));
assign g2738 = ((~g2327));
assign I4279 = ((~g2230));
assign g2264 = ((~I3405));
assign g4032 = (g441&g3388);
assign g4855 = ((~I6573));
assign I7472 = ((~g5626));
assign g4424 = ((~I5923));
assign g3317 = (g2722&g2895);
assign g5572 = ((~g5399));
assign g1686 = ((~I2675))|((~I2676));
assign I7312 = ((~g5364))|((~I7311));
assign g5042 = ((~I6672));
assign g895 = ((~g139));
assign g4441 = (g4372)|(g4039);
assign g851 = ((~g606));
assign g1582 = ((~g784))|((~g774))|((~g821));
assign g2874 = ((~g1849));
assign I2352 = ((~g1161));
assign g2120 = ((~I3251));
assign g4761 = (g4567&g1674);
assign g4868 = (g4774&g2891);
assign I3581 = ((~g1491));
assign I3255 = ((~g1650));
assign I3746 = ((~g2035));
assign g1352 = ((~I2391));
assign g2846 = (g619&g2015);
assign g5899 = ((~g5753));
assign g1173 = ((~I2185));
assign g3605 = ((~I4802));
assign g3831 = (g2330&g3425);
assign g815 = ((~I1877));
assign g5579 = ((~I7333));
assign g2346 = ((~I3496));
assign g5535 = (g5353)|(g3300);
assign I2581 = ((~g946));
assign g1417 = ((~g873))|((~g889));
assign I8988 = ((~g6787));
assign g1157 = ((~g89))|((~g107));
assign g5237 = ((~g5083));
assign g6078 = ((~g5801));
assign g3567 = ((~g3074));
assign I2082 = ((~g19))|((~I2080));
assign g5538 = ((~g5331));
assign g1603 = ((~g1039)&(~g658));
assign g5904 = (g5812&g5664);
assign I5448 = ((~g3960));
assign I7527 = ((~g49))|((~g5662));
assign g856 = ((~g654));
assign I6250 = ((~g4514));
assign g3440 = ((~I4678));
assign g3890 = ((~g3575));
assign g5362 = (g4437&g5174);
assign I5259 = ((~g3719))|((~I5257));
assign g1118 = ((~g36));
assign g5897 = ((~g5731));
assign g4190 = ((~I5600));
assign g6648 = (g6579&g6234);
assign g3441 = ((~I4681));
assign I3953 = ((~g289))|((~I3952));
assign I8548 = ((~g6454));
assign I6118 = ((~g4406));
assign g1953 = ((~I3062));
assign g6244 = (g4759&g5891);
assign g4357 = (g3990&g3342);
assign g2284 = ((~I3431));
assign g6143 = ((~I7865));
assign g6303 = (g6258)|(g6094);
assign I9005 = ((~g6817));
assign g1819 = ((~I2877));
assign g1985 = ((~I3096));
assign I6464 = ((~g4562));
assign g3132 = (g2306&g1206);
assign I4375 = ((~g2254));
assign g6696 = ((~I8806));
assign g5869 = ((~g5649))|((~g1076))|((~g2081));
assign g6453 = (g6343)|(g5945);
assign g6575 = ((~g6486));
assign g2292 = (g1706&g736&g743);
assign I5612 = ((~g3910));
assign g5781 = ((~I7563))|((~I7564));
assign I2848 = ((~g1193));
assign g6367 = ((~I8165));
assign g3060 = ((~I4285));
assign I5759 = ((~g3836))|((~g3503));
assign g844 = ((~g578));
assign g6652 = ((~I8752));
assign I4133 = ((~g2040));
assign g6291 = (g5210&g6161);
assign I3373 = ((~g1320));
assign I5103 = ((~g3440));
assign g5587 = ((~I7349));
assign I2318 = ((~g1236));
assign g4444 = (g4378)|(g4042);
assign g6786 = ((~I8946));
assign g2435 = ((~g1138))|((~g1777))|((~g1157));
assign g4776 = ((~g4449)&(~g4453));
assign I6599 = ((~g4823));
assign I3462 = ((~g1450));
assign g3900 = ((~g3575));
assign I8359 = (g5232)|(g5236)|(g5216)|(g5226);
assign g3997 = (g1250&g3425&g2849);
assign g5168 = ((~g5099));
assign g6928 = ((~g4532))|((~g6926));
assign g4844 = ((~I6540));
assign g6596 = ((~I8656));
assign I3452 = ((~g1450));
assign g4580 = (g706&g4262);
assign g5580 = ((~I7336));
assign I2566 = (g749&g743&g736);
assign I8174 = ((~g6173));
assign g4626 = ((~g4270));
assign g2821 = (g1890&g910);
assign g918 = (g610&g602);
assign I1971 = ((~g236))|((~I1969));
assign I2745 = ((~g1249));
assign I5271 = ((~g3710))|((~I5269));
assign g5086 = ((~g4732));
assign g5648 = (g4507&g5545);
assign I3278 = ((~g1695));
assign I5207 = ((~g3267))|((~g3271));
assign g1673 = ((~I2653));
assign g6855 = (g6851)|(g2085);
assign g5190 = (g426&g4950);
assign g3731 = (g331&g3441);
assign I7012 = ((~g5316));
assign I3034 = ((~g1519));
assign g2327 = ((~I3481));
assign g1897 = ((~I2992));
assign g4177 = (g3933&g1372);
assign g2760 = ((~I3942));
assign I9149 = ((~g6884));
assign I4486 = ((~g3093));
assign I4327 = ((~g2525));
assign I2934 = ((~g1436))|((~I2933));
assign g6835 = ((~I9028));
assign g4016 = ((~I5320));
assign g2755 = ((~g2350));
assign g6518 = ((~I8470));
assign g2871 = ((~g1919));
assign g6467 = ((~I8335));
assign I2860 = ((~g1177));
assign I6507 = ((~g4644));
assign g2862 = ((~I4066));
assign g6717 = ((~g6669))|((~g5065))|((~g5062));
assign g6473 = (g2036&g6397&g1628);
assign g5597 = ((~I7361));
assign g1285 = ((~g852));
assign g4389 = (g449&g3798);
assign g5369 = (g143&g5247);
assign g3641 = (g2644&g2333);
assign I2050 = ((~g683));
assign I7569 = ((~g79))|((~g5678));
assign g4302 = ((~g4068));
assign g4014 = ((~I5316));
assign g4102 = ((~I5388));
assign g4735 = (g2018&g4577);
assign g6047 = (g5824&g1692);
assign I6625 = ((~g4745));
assign I6646 = ((~g4687));
assign g4280 = (g2138&g1764&g4007);
assign I5723 = ((~g3942));
assign g5646 = (g4502&g5544);
assign g3987 = (g3669)|(g3134);
assign g3351 = (g2760&g1931);
assign g6682 = (g6478)|(g6624)|(g6623);
assign g837 = ((~g353));
assign g1741 = ((~I2753));
assign g4745 = (g4468)|(g4569);
assign g5411 = ((~I7077));
assign I3322 = ((~g1333));
assign I6680 = ((~g4713));
assign g1639 = ((~g815));
assign g6881 = ((~I9110));
assign I3584 = ((~g1678));
assign g4074 = (g3301)|(g2699);
assign g1450 = ((~I2453));
assign g3378 = (g3136&g2932);
assign g5615 = ((~I7372));
assign I7832 = ((~g5943));
assign g2764 = ((~g2357));
assign g2103 = ((~I3225));
assign I6355 = ((~g4569));
assign I6308 = ((~g4443));
assign I1862 = ((~g278));
assign I5777 = ((~g3807));
assign g4439 = ((~I5952));
assign g4369 = (g3999&g3364);
assign g3636 = (g2701&g2327);
assign g3724 = (g117&g3251);
assign g5124 = ((~I6780));
assign g5590 = ((~I7352));
assign g2732 = (g2449&g1940);
assign g2893 = ((~g1985));
assign g1540 = ((~I2507))|((~I2508));
assign I2022 = ((~g528))|((~I2021));
assign I3446 = ((~g1689))|((~I3445));
assign g1204 = ((~g39));
assign g4791 = (g3936&g4636);
assign I5148 = ((~g3450));
assign g1653 = ((~I2630));
assign g5901 = ((~g5753));
assign I7217 = ((~g152))|((~I7216));
assign g4528 = ((~I6096));
assign I1986 = ((~g508))|((~g224));
assign I3782 = ((~g2145));
assign g6597 = ((~I8659));
assign g3173 = ((~I4410));
assign g5877 = ((~I7643));
assign g3380 = ((~g2831));
assign g3156 = (g242&g2464);
assign I8332 = ((~g6306));
assign g3306 = ((~g3057));
assign g6290 = (g6245)|(g6086);
assign g3765 = (g554&g3485);
assign I7258 = ((~g5458));
assign g3070 = ((~I4297));
assign g4523 = ((~I6081));
assign g6422 = ((~I8276));
assign I6753 = ((~g4772));
assign g6452 = (g6342)|(g5942);
assign g1805 = ((~I2854));
assign g5448 = ((~g5278));
assign g5556 = (g5015&g5445);
assign g6410 = ((~I8240));
assign I8684 = ((~g6567));
assign I5913 = ((~g3751));
assign I8194 = ((~g471))|((~g6188));
assign g5353 = (g5327&g3463);
assign g4384 = (g414&g3797);
assign I3319 = ((~g1636));
assign I9236 = ((~g6939));
assign I8429 = ((~g6425));
assign I6352 = ((~g4564));
assign I7469 = ((~g5625));
assign I7835 = ((~g5926));
assign I6330 = ((~g4560));
assign I7852 = ((~g5993));
assign g4320 = ((~g4011));
assign g2163 = ((~I3288));
assign g2808 = (g2009&g1581);
assign g6095 = ((~g2952))|((~g5854));
assign I6048 = ((~g4376));
assign g5920 = ((~I7692));
assign g6661 = (I8773)|(I8774);
assign g6267 = (g2953)|(g5884);
assign g843 = ((~g574));
assign I6972 = ((~g5135));
assign g4099 = ((~I5379));
assign g6585 = ((~I8623));
assign g3454 = (g2933&g1660);
assign g5175 = (g5094&g1384);
assign g4668 = (g4642&g4638);
assign g3100 = ((~I4347));
assign g4673 = (g4656&g4654);
assign g6520 = ((~I8476));
assign g4142 = ((~I5508));
assign g1770 = ((~I2805));
assign g6098 = (g1209&g5753);
assign g2840 = ((~g2538));
assign g5180 = (g414&g4950);
assign g1017 = ((~I2053));
assign I8671 = ((~g6519));
assign I1951 = ((~g524))|((~g248));
assign g4281 = ((~I5736));
assign g5685 = ((~g5552));
assign g4360 = (g184&g3785);
assign g3964 = (g3634)|(g3089);
assign g6538 = ((~g6469));
assign I3684 = ((~g1733));
assign g3725 = (g118&g3251);
assign g4125 = ((~I5457));
assign I2190 = ((~g297));
assign I6759 = ((~g4778));
assign I8367 = (g6313)|(g6124)|(g6127)|(g6144);
assign I7859 = ((~g6032));
assign I6441 = ((~g4624));
assign g922 = ((~I1947));
assign g6722 = ((~I8860));
assign g5187 = (g457&g4877);
assign g5557 = (g5016&g5448);
assign I5896 = ((~g3879));
assign I8978 = ((~g6792));
assign I8261 = ((~g6298));
assign I4066 = ((~g2582));
assign g1415 = ((~g1246));
assign g5784 = ((~I7583));
assign g3016 = ((~I4223));
assign g4651 = (g4357)|(g3643);
assign g3673 = ((~g3075));
assign g1739 = ((~I2749));
assign g3959 = ((~g3352)&(~g3360));
assign g715 = ((~g135));
assign g1936 = ((~g1756));
assign g5730 = ((~I7497));
assign g4641 = (g4347)|(g3627);
assign I6587 = ((~g4803));
assign I8509 = ((~g6437));
assign g4367 = (g193&g3788);
assign I3758 = ((~g2041));
assign g6353 = ((~I8113));
assign g6735 = ((~I8897));
assign g2949 = (g830&g1861);
assign g6526 = ((~I8494));
assign I2312 = ((~g897));
assign g2838 = ((~g2515));
assign g1781 = ((~I2825));
assign I2005 = ((~g212))|((~I2003));
assign g2782 = (g2518&g1985);
assign I2137 = ((~g1));
assign I4462 = ((~g2135));
assign g6548 = ((~I8548));
assign g3510 = ((~g2709));
assign g2947 = ((~g1411))|((~g2026));
assign g2667 = ((~I3811));
assign g5862 = ((~g5649))|((~g1529))|((~g1535))|((~g2068));
assign g4241 = ((~g3774)&(~g3341));
assign g2788 = ((~I3983));
assign I2839 = ((~g1123));
assign g3279 = (g2599&g2612);
assign g2831 = ((~g2007))|((~g862))|((~g1784));
assign g2927 = ((~g1979));
assign I8347 = (g5188)|(g5157)|(g5154)|(g5193);
assign g6916 = (g6903&g6901);
assign g6120 = ((~I7832));
assign g3294 = (g139&g2870);
assign g6234 = ((~g6057));
assign g5013 = (g4826)|(g4621);
assign I3291 = ((~g1714));
assign g1339 = ((~I2370));
assign g4544 = (g4410)|(g2995);
assign I3983 = ((~g2276));
assign g4647 = ((~g4296));
assign g6791 = (g6768)|(g3307);
assign I4291 = ((~g2241));
assign g4416 = (g3905&g1481);
assign I6499 = ((~g4504))|((~g3541));
assign I6500 = ((~g4504))|((~I6499));
assign I3040 = ((~g1770));
assign g2952 = ((~g2381));
assign g1747 = ((~I2760));
assign I2159 = ((~g465));
assign I8376 = (g6315)|(g6126)|(g6129)|(g6146);
assign g6394 = ((~I8195))|((~I8196));
assign g5692 = ((~I7451));
assign g4705 = ((~I6305));
assign g3766 = ((~I4955));
assign I4198 = ((~g2276));
assign I6528 = ((~g4815));
assign g5701 = (g5683&g3813);
assign g3292 = (g2214&g2667);
assign g5484 = (g378&g5331);
assign g1203 = ((~I2207));
assign g4390 = (g418&g3799);
assign g5543 = ((~g5331));
assign I7979 = (g6015)|(g6212)|(g4950)|(g4877);
assign g6478 = ((~I8342));
assign g1257 = ((~g845));
assign g1552 = ((~g1030));
assign g5255 = ((~g4933));
assign I2061 = ((~g7))|((~I2060));
assign g4711 = ((~I6315));
assign g1991 = ((~I3102));
assign g2436 = ((~I3569));
assign g1381 = ((~I2417));
assign g2628 = ((~I3770));
assign g5270 = ((~I6927));
assign g2263 = ((~I3399))|((~I3400));
assign g1143 = ((~I2172));
assign I2215 = ((~g695));
assign g3103 = (g212&g2353);
assign I5258 = ((~g3714))|((~I5257));
assign I9176 = ((~g6881));
assign g2869 = ((~g2433));
assign I5397 = ((~g3932));
assign g3741 = ((~g901))|((~g3433))|((~g2340));
assign g2109 = ((~I3235));
assign g5266 = ((~I6923));
assign g5455 = ((~g2330))|((~g5311));
assign I3626 = ((~g1684));
assign I2196 = ((~g3));
assign g4105 = ((~I5397));
assign g1879 = ((~g1603)&(~g1416));
assign g3226 = ((~I4477));
assign I8144 = ((~g6182));
assign g3700 = (g2276&g2837);
assign g1341 = ((~I2376));
assign g2378 = ((~I3525));
assign g4449 = (g4266&g2887);
assign g1246 = ((~I2237));
assign g4775 = ((~I6425));
assign g3079 = ((~I4312));
assign g3110 = ((~I4358));
assign g4841 = ((~I6531));
assign g5770 = ((~g5645));
assign g5229 = (g545&g4980);
assign g5635 = (g4498&g5542);
assign g4154 = ((~I5548));
assign I4429 = ((~g2102));
assign g5300 = ((~I6952));
assign I8745 = ((~g6513));
assign g4814 = ((~g4550))|((~g1575))|((~g1550))|((~g2073));
assign g6149 = (g3200&g5997);
assign g6564 = ((~I8576));
assign g6403 = ((~I8223));
assign g4942 = (g175&g4736);
assign I8232 = ((~g6332));
assign g3789 = ((~g3388));
assign g3316 = (g2748&g2894);
assign g3461 = ((~g2986));
assign g1491 = ((~I2476));
assign g1646 = ((~I2617));
assign g1027 = (g598&g567);
assign g1715 = ((~I2716));
assign I8226 = ((~g6328));
assign g3686 = (g2256&g2819);
assign g6273 = (g5681)|(g5955);
assign g2857 = ((~I4059));
assign I3053 = ((~g1407));
assign g5023 = (g3935&g4804);
assign g5414 = (g382&g5278);
assign g2102 = ((~I3222));
assign g3668 = (g2568&g3124);
assign g4098 = ((~I5376));
assign I3590 = ((~g1781));
assign I3714 = ((~g1852));
assign g5144 = (g166&g5099);
assign I9203 = ((~g6921));
assign g3953 = (g3554&g188);
assign g4615 = ((~g4322));
assign g5919 = ((~I7689));
assign g3746 = (g3357)|(g2771);
assign g5368 = (g5201)|(g4932);
assign I6280 = ((~g4430));
assign g2937 = (g2160&g931);
assign I4459 = ((~g2134));
assign I4176 = ((~g2268));
assign I2240 = ((~g19));
assign g2748 = ((~I3923));
assign g4296 = ((~I5753));
assign I3355 = ((~g1608));
assign g4231 = (g3997)|(g4000);
assign g2699 = (g2397&g1905);
assign g6339 = ((~I8093));
assign g5941 = (g5777&g5399);
assign g1812 = ((~I2867));
assign g5063 = ((~g4799));
assign g964 = ((~g357));
assign I9227 = ((~g6937));
assign g6887 = ((~I9128));
assign g3222 = ((~I4465));
assign I5379 = ((~g3940));
assign g4301 = ((~I5767))|((~I5768));
assign g3551 = (g2937&g938);
assign g6278 = ((~I7966));
assign g5666 = (g5555)|(g5406);
assign I3261 = ((~g1783));
assign g4781 = ((~I6437));
assign g6103 = ((~I7805));
assign g5316 = ((~I6976));
assign g2457 = ((~I3587));
assign g5019 = ((~I6660))|((~I6661));
assign g6343 = (g6268&g6078);
assign I4337 = ((~g1934));
assign I6786 = ((~g4824));
assign g1823 = ((~I2887));
assign g4214 = (g1822&g4045);
assign g2828 = ((~g2488));
assign g4167 = (g378&g3898);
assign g3888 = (g3672)|(g3682);
assign g3976 = ((~I5252));
assign g1699 = ((~I2703));
assign I3281 = ((~g1761));
assign I6195 = ((~g4199))|((~I6194));
assign g6607 = ((~I8687));
assign g5728 = (g5623&g3889);
assign I1868 = ((~g280));
assign g6285 = ((~I8005));
assign g1284 = ((~g851));
assign I2782 = ((~g1177));
assign g2886 = ((~g1966));
assign g1109 = ((~I2137));
assign I3010 = ((~g1504));
assign g4937 = (g166&g4732);
assign I4189 = ((~g2159));
assign I8005 = ((~g6110));
assign g1504 = ((~I2485));
assign g1054 = ((~g485));
assign g3832 = ((~I5023));
assign I2773 = ((~g1191));
assign g2778 = ((~g2391));
assign g6874 = (g6873&g2060);
assign g4458 = (g4401)|(g4057);
assign g2194 = ((~I3331));
assign g6254 = (g532&g5897);
assign I8555 = ((~g6456));
assign g1914 = ((~I3013));
assign g1106 = ((~I2128));
assign I8356 = (g6311)|(g6123)|(g6125)|(g6141);
assign I5324 = ((~g3466));
assign g4726 = ((~I6352));
assign g1064 = ((~g102));
assign g4836 = (g4527&g4523);
assign g2660 = ((~I3804));
assign I3422 = ((~g1641));
assign I8497 = ((~g6481));
assign I9047 = ((~g6838));
assign g3481 = ((~g2612));
assign g6192 = ((~g5946));
assign g3042 = ((~I4261));
assign I2873 = ((~g1161));
assign g3924 = (g3505&g471);
assign g2360 = ((~g1793));
assign g2080 = ((~I3189))|((~I3190));
assign g4586 = ((~g4161)&(~g4165));
assign g3714 = ((~g3041));
assign g5348 = (g5317)|(g5122);
assign g6726 = ((~I8872));
assign I4799 = ((~g2967));
assign g2722 = ((~I3883));
assign I3656 = ((~g1484));
assign g2397 = ((~I3540));
assign g2801 = ((~I4003));
assign I3623 = ((~g1491));
assign I2165 = ((~g690));
assign g6570 = ((~I8594));
assign g6540 = ((~g6474));
assign g3370 = ((~g3124));
assign g2604 = ((~I3736));
assign g6501 = ((~I8423));
assign g2173 = ((~I3310));
assign I4465 = ((~g2945));
assign I5750 = ((~g4022));
assign g5717 = ((~I7478));
assign I4285 = ((~g2555));
assign g766 = ((~I1856));
assign I8126 = (g6194)|(g5958)|(g5975)|(g5997);
assign I5713 = ((~g4022));
assign I2506 = ((~g1047))|((~g1044));
assign g3863 = (g3692)|(g3172);
assign g5699 = (g5660)|(g5487);
assign g5493 = ((~I7197));
assign g1902 = ((~I3001));
assign g4621 = (g3953&g4364);
assign g3620 = (g2422&g3060);
assign g4344 = (g3981&g3306);
assign I3022 = ((~g1426));
assign g4139 = ((~I5499));
assign g4497 = (g4166)|(g3784);
assign g5089 = ((~I6723));
assign g2353 = ((~I3505));
assign g941 = ((~I1995))|((~I1996));
assign g980 = ((~I2037));
assign g4037 = (g2896&g3388);
assign I8435 = ((~g6413));
assign g4807 = ((~g4473));
assign I8027 = ((~g6237));
assign g5425 = ((~I7091));
assign g3485 = ((~g2986));
assign g2739 = ((~I3906));
assign g3655 = (g2197&g2768);
assign g4323 = ((~g4086));
assign I2269 = ((~g899));
assign I6780 = ((~g4825));
assign g2512 = ((~I3638));
assign g5534 = ((~I7276));
assign g5633 = (g4496&g5539);
assign g5957 = ((~g5866));
assign I2638 = ((~g1123));
assign g5581 = ((~I7339));
assign g3546 = ((~g3095));
assign I5991 = ((~g4226));
assign I5658 = ((~g3983))|((~I5657));
assign g6161 = ((~g5926));
assign g2912 = ((~g2001));
assign g2873 = (g1845&g1861);
assign I5511 = ((~g3876));
assign g6061 = (g5824&g1711);
assign g2036 = ((~g1764));
assign g2856 = ((~g2010));
assign g4773 = (g4495)|(g4220);
assign g6836 = ((~I9031));
assign g1053 = ((~g197));
assign g4007 = ((~I5308))|((~I5309));
assign g6769 = (g6758&g2986);
assign g3652 = (g2544&g3096);
assign g5885 = ((~g5865));
assign g2473 = ((~I3605));
assign I6470 = ((~g4473));
assign I2147 = ((~g6));
assign g1685 = ((~I2671));
assign I1996 = ((~g218))|((~I1994));
assign g5453 = ((~g5296));
assign g5328 = ((~I6986));
assign g3122 = (g2435&g1394);
assign g4376 = ((~I5843));
assign g3280 = (g2177&g2637);
assign g853 = ((~g642));
assign I6425 = ((~g4619));
assign g2935 = (g2291&g1788);
assign I8459 = ((~g6427));
assign I8438 = ((~g6416));
assign g5853 = ((~g5638))|((~g2053))|((~g1076));
assign I7397 = ((~g5561));
assign g5430 = (g5161)|(g4873);
assign g6164 = ((~g5926));
assign g3526 = ((~g3196))|((~g3023))|((~g2197))|((~g2981));
assign I3665 = ((~g1824));
assign g896 = ((~g22));
assign I2081 = ((~g25))|((~I2080));
assign g6852 = (g6847&g2295);
assign g5113 = ((~I6753));
assign I4446 = ((~g606))|((~I4444));
assign g4462 = ((~I5977));
assign g2081 = (g1094&g1546);
assign g1075 = ((~I2109))|((~I2110));
assign g6466 = ((~I8332));
assign g4767 = ((~g4601));
assign g5097 = ((~I6733));
assign g3318 = ((~I4593));
assign g6552 = ((~I8552));
assign g3637 = (g2822&g2752);
assign g6578 = ((~g6489));
assign g836 = ((~g349));
assign I8761 = ((~g6563));
assign g905 = ((~g301))|((~g319));
assign I4003 = ((~g2284));
assign g3830 = ((~I5019));
assign g6918 = (g6911)|(g6913);
assign g4442 = (g4239&g2882);
assign I7988 = (g6015)|(g6212)|(g4950)|(g4877);
assign I2964 = ((~g1257));
assign I3198 = ((~g1819));
assign g3303 = (g2722&g2890);
assign g2491 = ((~I3620));
assign g5573 = ((~g5403));
assign g3749 = (g3371)|(g2793);
assign g3134 = (g230&g2413);
assign g2159 = ((~I3284));
assign g1322 = ((~I2321));
assign g1787 = ((~I2835));
assign g2449 = ((~I3584));
assign g1807 = ((~I2860));
assign g5625 = (g5495)|(g3281);
assign g5619 = (g5064&g5527);
assign I2225 = ((~g696));
assign g2394 = ((~I3537));
assign g5022 = ((~I6666));
assign I5421 = ((~g3724));
assign I3144 = ((~g1319));
assign g3872 = ((~g3312));
assign I5920 = ((~g4228));
assign g1325 = ((~I2330));
assign g4423 = ((~I5920));
assign g6245 = (g1329&g5889);
assign g4562 = ((~I6132));
assign g2894 = ((~g1891));
assign I3177 = ((~g1706))|((~g736));
assign g6935 = (g6933&g3622);
assign I5227 = ((~g3259))|((~I5226));
assign g1687 = ((~I2682))|((~I2683));
assign g6702 = (g6659)|(g496);
assign g3961 = ((~I5208))|((~I5209));
assign g4911 = ((~I6615));
assign g5506 = ((~I7231))|((~I7232));
assign g6495 = ((~g6354)&(~g1775));
assign I4752 = ((~g2859));
assign g2888 = ((~g1972));
assign I7817 = ((~g5924));
assign I7164 = ((~g5433));
assign g6934 = (g6932&g3605);
assign g1631 = ((~I2588));
assign g1835 = ((~I2919));
assign I7404 = ((~g5541));
assign g4253 = (g1861&g3819);
assign g5083 = (g4688)|(g4271);
assign g1947 = ((~I3056));
assign g2317 = ((~I3471));
assign g6889 = ((~I9134));
assign g5093 = ((~g4683)&(~g4684));
assign g1436 = (g834&g830);
assign g971 = ((~g658));
assign g2587 = ((~I3714));
assign I2857 = ((~g1161));
assign I8617 = ((~g6539));
assign g3666 = (g3128&g2787);
assign I6635 = ((~g4745));
assign g5240 = (g293&g4915);
assign g4535 = ((~g4173));
assign g3456 = ((~g2640));
assign g6484 = ((~g6361));
assign I7970 = (g6015)|(g6212)|(g4950)|(g4877);
assign g3702 = (g2284&g2839);
assign g4635 = (g4342)|(g3616);
assign I7086 = ((~g5281));
assign g6631 = (g1838&g6545);
assign g5861 = ((~g5636));
assign g2960 = ((~I4151))|((~I4152));
assign g1305 = ((~I2293));
assign g4856 = ((~I6576));
assign I3553 = ((~g1305));
assign I4270 = ((~g2555));
assign I7251 = ((~g5458));
assign I8128 = (g5202)|(g4993)|(g4967)|(g4980);
assign g3145 = (g2397&g2443);
assign I5106 = ((~g3247));
assign g4518 = ((~I6066));
assign g2580 = ((~I3691));
assign g1898 = ((~I2995));
assign I7432 = ((~g111))|((~g5554));
assign g1811 = ((~I2864));
assign I5466 = ((~g3787));
assign I3343 = ((~g1623));
assign I7051 = ((~g5219));
assign g4392 = ((~I5879));
assign g1471 = ((~I2464));
assign I3875 = ((~g285))|((~I3874));
assign g5911 = (g5817&g5670);
assign g3839 = ((~I5040));
assign g2283 = ((~I3428));
assign g1666 = ((~g1088));
assign I5831 = ((~g3842));
assign g1777 = ((~g1060))|((~g102))|((~g89));
assign g2794 = (g2544&g1994);
assign g6256 = (g1696&g6040);
assign g4473 = (g3575)|(g4253);
assign g4209 = (g3816&g865);
assign g5688 = ((~g5546))|((~g1585))|((~g2084))|((~g2916));
assign g3331 = ((~g3076));
assign g2040 = ((~g1738));
assign g3879 = (g3704)|(g3195);
assign g729 = ((~I1838));
assign g1587 = ((~g1123));
assign I1942 = ((~g664));
assign I6060 = ((~g4380));
assign I4527 = ((~g2909))|((~I4526));
assign g1674 = ((~g985));
assign g1112 = ((~g336));
assign g5647 = ((~g5509));
assign g4721 = ((~I6343));
assign I5728 = ((~g4022));
assign I5774 = ((~g3807));
assign g6891 = ((~I9140));
assign I3979 = ((~g1836));
assign g5645 = ((~g5537));
assign g5501 = (g5454&g3478);
assign I3102 = ((~g1426));
assign g5043 = (g3941&g4805);
assign g3372 = (g254&g2905);
assign g3241 = ((~I4522));
assign g3730 = (g328&g3441);
assign g6409 = ((~g6285));
assign g2481 = ((~I3608));
assign I3819 = ((~g2044));
assign g2615 = ((~I3755));
assign g2598 = ((~I3726));
assign g6718 = (g4511&g6661);
assign g4176 = (g386&g3901);
assign I2925 = ((~g1762));
assign I6737 = ((~g4662));
assign I9220 = ((~g6930));
assign I8051 = ((~g6108));
assign I2367 = ((~g1161));
assign g3448 = ((~I4684));
assign g4052 = (g418&g3388);
assign I7695 = ((~g5714));
assign I4492 = ((~g3001));
assign g2747 = (g2449&g1957);
assign I6795 = ((~g5022));
assign g6785 = ((~I8943));
assign g6537 = ((~I8527));
assign g4011 = ((~g3486));
assign I3988 = ((~g291))|((~g2544));
assign g6246 = (g5665)|(g5937);
assign g6211 = ((~g5992));
assign g5472 = (g5361)|(g5144);
assign g2830 = ((~g2494));
assign g5123 = (g4670&g1936);
assign I9146 = ((~g6890));
assign g1849 = ((~I2949));
assign I2933 = ((~g1436))|((~g345));
assign g4792 = (g1417&g4471);
assign I3868 = ((~g2125));
assign g6517 = ((~I8467));
assign g2765 = ((~I3946));
assign g4581 = ((~g4156)&(~g4160));
assign g4448 = (g3815&g4225);
assign I6397 = ((~g4473));
assign g1640 = ((~I2601));
assign g1176 = ((~I2190));
assign g6325 = ((~I8061));
assign I5862 = ((~g3863));
assign g1286 = ((~g854));
assign g6676 = (g6631)|(g6555);
assign I3650 = ((~g1650));
assign g6418 = ((~I8264));
assign g4407 = (g4054&g74);
assign I3385 = ((~g1318));
assign I8721 = ((~g6534));
assign I9066 = (g5189)|(g5269)|(g6400);
assign I3632 = ((~g1295));
assign I3307 = ((~g1339));
assign g1503 = ((~g878));
assign g6831 = (g6812&g5975);
assign g6096 = (g1193&g5753);
assign g2863 = ((~g2296));
assign I7910 = ((~g5905));
assign g5419 = (g386&g5292);
assign g4693 = ((~I6283));
assign g6423 = ((~I8279));
assign I3736 = ((~g2460));
assign g5902 = (g5808&g5661);
assign g2464 = ((~I3596));
assign g4092 = (g3311)|(g2721);
assign I6196 = ((~g631))|((~I6194));
assign I7218 = ((~g5368))|((~I7216));
assign g4368 = (g3998&g3363);
assign g6595 = ((~I8653));
assign g6113 = (g5902)|(g5601);
assign I8387 = (g5178)|(g5209)|(g6281);
assign g6781 = (g6718)|(g6748);
assign g5483 = (g374&g5331);
assign I7805 = ((~g5923));
assign g5167 = (g5011&g1556);
assign g4787 = (g2937&g4628);
assign g3477 = ((~g2692));
assign g4602 = (g4407&g4293);
assign g3974 = ((~I5243))|((~I5244));
assign I2327 = ((~g1222));
assign I7612 = ((~g5605));
assign g4810 = ((~I6488));
assign g5361 = (g4435&g5168);
assign I5746 = ((~g4022));
assign g3602 = (g2688&g2663);
assign g1119 = ((~I2159));
assign g5691 = ((~g5568));
assign g5896 = ((~g5753));
assign g1372 = ((~I2408));
assign g3251 = ((~I4534));
assign g1612 = (g784&g774&g821&I2574);
assign g2169 = ((~I3298));
assign g5153 = (g492&g4904);
assign g5674 = (g5558)|(g5419);
assign g6649 = ((~I8745));
assign g5898 = (g5800&g5647);
assign g5679 = (g74&g5576);
assign g1048 = ((~g492));
assign I4192 = ((~g1847));
assign g6711 = ((~I8843));
assign g857 = ((~g170));
assign I4441 = ((~g2109));
assign g1884 = ((~I2979));
assign g5236 = (g269&g4915);
assign g2232 = ((~I3361));
assign I2760 = ((~g1193));
assign g6304 = (g5915&g6165);
assign I6027 = ((~g4223))|((~I6026));
assign I3694 = ((~g1811));
assign I5529 = ((~g3854));
assign g5905 = ((~g5852));
assign I2321 = ((~g898));
assign g3263 = ((~g3015));
assign g2998 = ((~I4195));
assign g4402 = ((~g4017));
assign g5176 = (g410&g4950);
assign I8208 = (g6194)|(g5958)|(g5975)|(g5997);
assign g6653 = ((~I8755));
assign g5926 = ((~g5741))|((~g639));
assign I6366 = ((~g4569));
assign g4697 = (g4589&g1363);
assign I3189 = ((~g1716))|((~I3188));
assign g5539 = ((~g5331));
assign I6296 = ((~g4436));
assign g4234 = (g3921)|(g478);
assign I8252 = ((~g6294));
assign g4261 = ((~g3762)&(~g3295));
assign I2411 = ((~g736));
assign g3449 = (g128&g2946);
assign g5015 = (g4787)|(g4588);
assign I8749 = ((~g6560));
assign g4815 = ((~I6495));
assign g4243 = (g4053)|(g4058);
assign g4618 = ((~g4246));
assign g3339 = (g2734&g1914);
assign I3791 = ((~g2044));
assign g3709 = (g2284&g2845);
assign g4198 = ((~I5618));
assign g5384 = ((~g5220));
assign g2433 = ((~g1418)&(~g1449));
assign I3972 = ((~g2518))|((~I3970));
assign g6292 = (g6243)|(g6084);
assign g5658 = ((~g5512));
assign g6602 = ((~I8674));
assign g4843 = ((~I6537));
assign I7865 = ((~g6095));
assign g5891 = ((~g5731));
assign g4659 = ((~I6250));
assign I8690 = ((~g6571));
assign g4358 = (g3991&g3343);
assign g1449 = ((~g489)&(~g1048));
assign g4496 = ((~I6008));
assign g4903 = ((~g4717))|((~g858));
assign g3764 = (g551&g3480);
assign g5997 = ((~g5854));
assign g4799 = ((~g4485));
assign g3108 = ((~I4354));
assign I1859 = ((~g277));
assign g5371 = (g152&g5248);
assign g5809 = ((~I7608));
assign I4354 = ((~g1953));
assign g4862 = (g4739)|(g4489);
assign g5783 = ((~I7577))|((~I7578));
assign g6873 = ((~g6848))|((~g3621));
assign I4534 = ((~g2858));
assign I3797 = ((~g2125));
assign g2308 = ((~I3452));
assign g2837 = ((~g2512));
assign g4652 = (g4358)|(g3645);
assign g6146 = (g3192&g5997);
assign g2928 = (g2100)|(g1582);
assign g5753 = ((~g1477)&(~g5688));
assign g4642 = (g4348)|(g3628);
assign g6772 = (g6746&g3312);
assign g2789 = ((~g2410));
assign g2154 = ((~I3271));
assign g5549 = ((~g5331));
assign g3015 = ((~I4220));
assign I3062 = ((~g1776));
assign I8346 = (g6159)|(g6334)|(g5163)|(g5191);
assign I3808 = ((~g2125));
assign g4869 = ((~g4662));
assign g3694 = (g3147&g64);
assign g4648 = (g4407&g79);
assign g3525 = ((~g3192))|((~g3002))|((~g2197))|((~g2179));
assign g3295 = (g2660&g2647);
assign I8758 = ((~g6562));
assign g6235 = ((~g6062));
assign I8135 = (g6194)|(g5958)|(g5975)|(g5997);
assign g3819 = (g964&g3437);
assign g4165 = (g3927&g1352);
assign g1764 = ((~I2796))|((~I2797));
assign g5490 = ((~I7190));
assign g1649 = ((~g985));
assign I6946 = ((~g5124));
assign g3614 = (g2998&g2691);
assign I2044 = ((~g681));
assign g6882 = ((~I9113));
assign g5235 = (g554&g4980);
assign g6060 = (g5824&g1703);
assign I7276 = ((~g5375));
assign I6501 = ((~g3541))|((~I6499));
assign g3216 = ((~I4459));
assign I8342 = ((~g6314));
assign I6176 = ((~g4236))|((~I6175));
assign g4860 = (g4735)|(g4488);
assign g3305 = (g2960&g2296);
assign g2679 = ((~I3823));
assign g3798 = ((~g3388));
assign g6612 = ((~I8702));
assign g5616 = (g5505&g4929);
assign g4153 = ((~I5545));
assign g4121 = ((~I5445));
assign g6762 = (g6679)|(g6628)|(g6739);
assign I5854 = ((~g3857));
assign I2110 = ((~g610))|((~I2108));
assign g1338 = ((~I2367));
assign g4242 = ((~I5686));
assign g5469 = ((~I7153));
assign g1748 = ((~I2763));
assign I2154 = ((~g14));
assign I2376 = ((~g729));
assign I7494 = ((~g5691));
assign g5636 = ((~g5564))|((~g4769));
assign I2089 = ((~g33))|((~g29));
assign g6502 = ((~I8426));
assign g3388 = ((~I4667));
assign I2309 = ((~g1236));
assign g3172 = (g2449&g2491);
assign I8357 = (g6145)|(g6318)|(g5171)|(g5187);
assign g4495 = (g3913&g4292);
assign I5577 = ((~g4022));
assign g3843 = (g2856&g945&g3533);
assign g4359 = (g434&g3782);
assign g3866 = ((~I5091));
assign g5542 = ((~g5331));
assign g5720 = ((~I7481));
assign g3899 = (g323&g3441);
assign I3836 = ((~g1832));
assign I2497 = ((~g1042))|((~g1036));
assign g4235 = ((~g3780)&(~g3362));
assign g4822 = ((~g4614));
assign g4350 = ((~g4010));
assign g1256 = ((~g838));
assign g6194 = ((~I7906));
assign g4867 = (g4811&g3872);
assign I2460 = ((~g952));
assign g1156 = ((~I2175));
assign g917 = ((~I1942));
assign I1850 = ((~g210));
assign I4264 = ((~g2212));
assign I7557 = ((~g5674))|((~I7555));
assign g5354 = (g5249&g2903);
assign g3536 = ((~g3219))|((~g2215))|((~g3007))|((~g2179));
assign g6833 = ((~I9024));
assign I8662 = ((~g6525));
assign g6372 = ((~I8180));
assign I6012 = ((~g4167));
assign I1847 = ((~g209));
assign g2809 = ((~I4019));
assign g6369 = ((~I8171));
assign g2976 = ((~g2197));
assign g2110 = ((~g1381));
assign g5471 = (g5360)|(g5143);
assign I4235 = ((~g798))|((~I4233));
assign I2212 = ((~g123));
assign g3482 = ((~g2713));
assign g5596 = ((~I7358));
assign g5564 = ((~g5382));
assign I5649 = ((~g3968))|((~I5647));
assign g4529 = ((~I6099));
assign g6067 = ((~g5788));
assign g3727 = (g122&g3251);
assign g1771 = ((~I2808));
assign I8943 = ((~g6774));
assign I5157 = ((~g3454));
assign g1806 = ((~I2857));
assign g6411 = ((~I8243));
assign g2574 = ((~I3681));
assign g3634 = (g2179&g2744);
assign I9167 = ((~g6878));
assign g3012 = ((~I4204))|((~I4205));
assign I2402 = ((~g774));
assign g6539 = ((~I8531));
assign g3801 = ((~g3388));
assign I8506 = ((~g6483));
assign I6382 = ((~g4460));
assign I3016 = ((~g1754));
assign g3910 = (g3546&g1049);
assign I4782 = ((~g2846))|((~g622));
assign g2841 = ((~g2541));
assign g1193 = ((~I2204));
assign g4224 = ((~g4046));
assign I5699 = ((~g3844));
assign g6721 = ((~I8857));
assign g5555 = (g5014&g5442);
assign g4143 = ((~I5511));
assign I2831 = ((~g1209));
assign g3856 = (g3686)|(g3157);
assign I9217 = ((~g6931));
assign I3611 = ((~g1771));
assign g3793 = ((~g3491));
assign g3455 = ((~g2637));
assign g6905 = ((~I9182));
assign g2245 = ((~I3382));
assign g3219 = ((~I4462));
assign g3800 = ((~g3388));
assign I3672 = ((~g1656));
assign I5002 = ((~g3612));
assign g2948 = (g2137&g1595);
assign I3563 = ((~g1461));
assign g6344 = (g6272&g6080);
assign I6744 = ((~g4708))|((~I6743));
assign g3599 = (g2935)|(g1637);
assign g3155 = (g248&g2461);
assign g4223 = ((~I5658))|((~I5659));
assign g6586 = ((~I8626));
assign g1189 = ((~I2196));
assign g3998 = (g3698)|(g3180);
assign g5188 = (g1043&g4894);
assign g4674 = ((~g4550))|((~g1514))|((~g2107))|((~g2897));
assign g5154 = (g500&g4993);
assign g4753 = ((~I6377));
assign I6564 = ((~g4712));
assign g2700 = (g2370&g1908);
assign I4306 = ((~g1898));
assign g4124 = ((~I5454));
assign I7520 = ((~g361))|((~g5659));
assign g6090 = (g1161&g5742);
assign I7349 = ((~g5532));
assign I6075 = ((~g4386));
assign g6331 = (g3891&g6212);
assign g6104 = ((~I7808));
assign g1738 = ((~g1108));
assign g3975 = ((~I5249));
assign g3621 = ((~g1407)&(~g2842));
assign I5352 = (g3529&g3531&g3535&g3538);
assign g4361 = (g3995&g3354);
assign g4215 = ((~I5637));
assign g6328 = ((~I8066));
assign I6020 = ((~g4176));
assign g2685 = (g2370&g1887);
assign g2885 = ((~g1963));
assign g6606 = ((~I8684));
assign I2648 = ((~g980));
assign I3431 = ((~g1275));
assign I3890 = ((~g2145));
assign g6043 = ((~g5824));
assign I5182 = ((~g3271));
assign g5665 = (g361&g5570);
assign I3705 = ((~g2316));
assign g4431 = ((~I5938));
assign g1730 = ((~g1114));
assign g4612 = ((~g4320));
assign g2381 = ((~I3528));
assign I2414 = ((~g784));
assign I5391 = ((~g3975));
assign g1740 = ((~g1116));
assign g6725 = ((~I8869));
assign I3025 = ((~g1439));
assign g4300 = ((~I5760))|((~I5761));
assign g3559 = ((~g2603));
assign g829 = ((~g323));
assign I6689 = ((~g4758));
assign g5181 = (g449&g4877);
assign g5317 = (g148&g4869);
assign g4770 = ((~I6414));
assign g3204 = ((~I4441));
assign I3170 = ((~g1534))|((~I3168));
assign I7045 = ((~g5167));
assign I5657 = ((~g3983))|((~g3979));
assign g6428 = ((~I8290));
assign g4938 = ((~I6630));
assign g5420 = ((~I7086));
assign I7980 = (g5202)|(g4993)|(g4967)|(g4980);
assign g3345 = (g236&g2886);
assign g2361 = ((~I3513));
assign g6354 = (g5866&g6193);
assign g5349 = (g5324&g3451);
assign g6479 = (I8349)|(g6335);
assign I3179 = ((~g736))|((~I3177));
assign g2637 = ((~I3779));
assign g6509 = ((~I8447));
assign g2101 = (g1001&g1543);
assign I2570 = ((~g1222));
assign I2125 = ((~g698));
assign g6532 = ((~I8512));
assign g5727 = ((~I7490));
assign I3447 = ((~g729))|((~I3445));
assign g6643 = (g6574&g6229);
assign g2829 = ((~g2491));
assign I6430 = ((~g4620));
assign g5470 = (g5359)|(g5142);
assign g2488 = ((~I3617));
assign I8702 = ((~g6572));
assign g4943 = ((~I6635));
assign g4049 = ((~g3677))|((~g3425));
assign g2770 = (g2518&g1972);
assign g1107 = ((~I2131));
assign g4782 = (g1624&g4623);
assign g4171 = (g3956&g2104);
assign I6039 = ((~g4182));
assign g4629 = ((~g4276));
assign g3043 = ((~I4264));
assign g4273 = ((~I5728));
assign g4587 = ((~g4215));
assign g2951 = ((~g2142))|((~g1797));
assign g4166 = ((~I5568));
assign g6922 = ((~I9203));
assign g5494 = (g5443&g3455);
assign g5938 = (g5114&g5791);
assign I5337 = ((~g3564));
assign I5739 = ((~g3942));
assign I8869 = ((~g6694));
assign g5215 = (g4864&g5090);
assign g3278 = (g2175&g2628);
assign g6284 = ((~I8002));
assign g1754 = ((~I2773));
assign I3125 = ((~g1279))|((~g1276));
assign g3324 = (g230&g2875);
assign g5088 = ((~g4691)&(~g4697));
assign g2142 = (g1793&g1777);
assign I3895 = ((~g2422))|((~I3893));
assign g4033 = (g426&g3388);
assign I7107 = ((~g5277));
assign I5033 = ((~g3527));
assign g6270 = (g1726&g6062);
assign g4485 = ((~I5987));
assign g4438 = (g4363)|(g4037);
assign I6555 = ((~g4703));
assign I9134 = ((~g6864));
assign I4976 = ((~g3575));
assign g5296 = ((~I6946));
assign g5456 = ((~g5300));
assign g4833 = (g4521&g4516);
assign g3925 = ((~g3303)&(~g3315));
assign I1987 = ((~g508))|((~I1986));
assign I3605 = ((~g1681));
assign g6320 = (g3869&g6194);
assign I8710 = ((~g6517));
assign I2033 = ((~g678));
assign I7990 = (g4915)|(g5025);
assign g4620 = ((~g4251));
assign I2115 = ((~g687));
assign g1142 = ((~I2169));
assign I2808 = ((~g1161));
assign g2031 = ((~I3140));
assign g4980 = ((~g4678));
assign I7989 = (g5202)|(g4993)|(g4967)|(g4980);
assign I8482 = ((~g6461));
assign g6404 = ((~I8226));
assign I3405 = ((~g1321));
assign g3361 = (g3150&g1950);
assign I3886 = ((~g2215));
assign g3227 = ((~I4480));
assign g6581 = ((~g6493));
assign g5702 = ((~I7463));
assign I5050 = ((~g3246));
assign g2266 = ((~I3412))|((~I3413));
assign g3293 = (g212&g2864);
assign I4664 = ((~g2924));
assign g6719 = (g4518&g6665);
assign g3952 = ((~I5182));
assign g3740 = (g3335)|(g2747);
assign g3381 = (g3128&g1998);
assign g1340 = ((~I2373));
assign g1623 = ((~I2578));
assign I7146 = ((~g5231));
assign g3739 = (g3334)|(g2746);
assign g6749 = (g6735&g6734);
assign g1263 = ((~g846));
assign I8767 = ((~g6619));
assign I8223 = ((~g6325));
assign I8162 = ((~g6189));
assign I5257 = ((~g3714))|((~g3719));
assign g6079 = (g1236&g5753);
assign g3687 = (g2245&g2820);
assign g1101 = ((~I2125));
assign g4398 = ((~I5893));
assign g3810 = (g625&g3421);
assign g6375 = ((~I8189));
assign g4381 = ((~I5854));
assign I7814 = ((~g5922));
assign g1792 = ((~I2848));
assign I4294 = ((~g2525));
assign g6929 = ((~g4536))|((~g6927));
assign I7643 = ((~g5752));
assign g3349 = (g2783&g1925);
assign g6845 = (I9064)|(I9065)|(I9066);
assign g1254 = ((~g152));
assign g4199 = (g628&g3810);
assign g4112 = ((~I5418));
assign g1355 = ((~I2394));
assign g842 = ((~g571));
assign I3587 = ((~g1461));
assign g4182 = (g394&g3904);
assign g6119 = ((~I7829));
assign g6129 = (g5717&g5975);
assign g1714 = ((~g1110));
assign g6610 = ((~I8696));
assign g3979 = ((~I5258))|((~I5259));
assign I8485 = ((~g6479));
assign g3281 = (g2178&g2640);
assign g4000 = ((~g1250)&(~g3425));
assign I2588 = ((~g1193));
assign g5194 = (g586&g4874);
assign I8377 = (g6150)|(g6324)|(g5180)|(g5181);
assign g2783 = ((~I3979));
assign g6819 = ((~I8994));
assign g6563 = ((~I8573));
assign I7361 = ((~g5566));
assign g2197 = ((~I3340));
assign g4859 = (g4730)|(g4486);
assign g2756 = ((~g2353));
assign g4680 = ((~g4550))|((~g1514))|((~g1006))|((~g2897));
assign I5977 = ((~g4319));
assign g6360 = ((~I8144));
assign g4450 = (g4389)|(g4047);
assign g5024 = (g4793)|(g4600);
assign g5367 = (g5199)|(g4928);
assign g5942 = (g5117&g5797);
assign g3774 = (g3016&g3510);
assign g2779 = ((~g2394));
assign I5292 = ((~g3421))|((~g625));
endmodule
