//NOTE: no-implementation module stub

module SW10200C (
    input  wire [4:0] A0,
    input  wire [4:0] A1,
    input  wire [4:0] A2,
    input  wire [4:0] A3,
    input  wire [4:0] A4,
    input  wire [4:0] B0,
    input  wire [4:0] B1,
    input  wire [4:0] B2,
    input  wire [4:0] B3,
    input  wire [4:0] B4,
    input  wire CKA,
    input  wire CKB,
    input  wire CSA,
    input  wire CSB,
    input  wire [11:0] DI0,
    input  wire [11:0] DI1,
    input  wire [11:0] DI2,
    input  wire [11:0] DI3,
    input  wire [11:0] DI4,
    input  wire [11:0] DI5,
    input  wire [11:0] DI6,
    input  wire [11:0] DI7,
    input  wire [11:0] DI8,
    input  wire [11:0] DI9,
    input  wire [11:0] DI10,
    input  wire [11:0] DI11,
    output reg [11:0] DO0,
    output reg [11:0] DO1,
    output reg [11:0] DO2,
    output reg [11:0] DO3,
    output reg [11:0] DO4,
    output reg [11:0] DO5,
    output reg [11:0] DO6,
    output reg [11:0] DO7,
    output reg [11:0] DO8,
    output reg [11:0] DO9,
    output reg [11:0] DO10,
    output reg [11:0] DO11,
    input  wire WEB,
    input  wire OE
);

endmodule
