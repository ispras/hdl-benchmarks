module test ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , 
 n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , 
 n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , 
 n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , 
 n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , 
 n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , 
 n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , 
 n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , 
 n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , 
 n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , 
 n181 , n182 , n183 , n184 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 ;
output n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , 
 n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , 
 n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , 
 n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , 
 n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , 
 n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , 
 n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , 
 n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , 
 n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , 
 n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , 
 n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , 
 n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , 
 n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 ;
wire n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , 
 n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , 
 n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , 
 n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , 
 n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , 
 n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , 
 n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , 
 n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , 
 n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , 
 n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , 
 n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , 
 n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , 
 n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , 
 n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , 
 n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , 
 n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , 
 n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , 
 n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , 
 n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , 
 n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , 
 n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , 
 n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , 
 n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , 
 n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , 
 n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , 
 n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , 
 n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , 
 n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , 
 n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , 
 n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , 
 n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , 
 n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , 
 n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , 
 n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , 
 n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , 
 n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , 
 n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , 
 n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , 
 n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , 
 n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , 
 n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , 
 n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , 
 n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , 
 n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , 
 n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , 
 n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , 
 n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , 
 n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , 
 n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , 
 n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , 
 n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , 
 n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , 
 n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , 
 n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , 
 n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , 
 n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , 
 n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , 
 n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , 
 n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , 
 n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , 
 n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , 
 n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , 
 n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , 
 n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , 
 n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , 
 n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , 
 n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , 
 n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , 
 n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , 
 n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , 
 n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , 
 n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , 
 n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , 
 n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , 
 n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , 
 n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , 
 n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , 
 n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , 
 n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , 
 n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , 
 n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , 
 n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , 
 n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , 
 n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , 
 n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , 
 n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , 
 n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , 
 n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , 
 n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , 
 n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , 
 n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , 
 n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , 
 n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , 
 n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , 
 n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , 
 n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , 
 n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , 
 n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , 
 n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , 
 n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , 
 n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , 
 n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , 
 n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , 
 n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , 
 n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , 
 n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , 
 n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , 
 n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , 
 n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , 
 n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , 
 n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , 
 n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , 
 n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , 
 n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , 
 n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , 
 n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , 
 n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , 
 n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , 
 n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , 
 n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , 
 n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , 
 n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , 
 n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , 
 n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , 
 n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , 
 n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , 
 n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , 
 n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , 
 n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , 
 n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , 
 n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , 
 n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , 
 n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , 
 n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , 
 n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , 
 n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , 
 n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , 
 n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , 
 n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , 
 n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , 
 n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , 
 n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , 
 n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , 
 n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , 
 n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , 
 n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , 
 n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , 
 n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , 
 n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , 
 n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , 
 n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , 
 n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , 
 n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , 
 n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , 
 n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , 
 n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , 
 n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , 
 n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , 
 n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , 
 n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , 
 n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , 
 n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , 
 n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , 
 n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , 
 n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , 
 n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , 
 n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , 
 n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , 
 n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , 
 n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , 
 n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , 
 n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , 
 n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , 
 n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , 
 n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , 
 n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , 
 n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , 
 n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , 
 n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , 
 n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , 
 n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , 
 n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , 
 n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , 
 n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , 
 n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , 
 n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , 
 n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , 
 n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , 
 n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , 
 n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , 
 n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , 
 n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , 
 n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , 
 n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , 
 n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , 
 n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , 
 n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , 
 n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , 
 n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , 
 n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , 
 n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , 
 n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , 
 n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , 
 n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , 
 n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , 
 n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , 
 n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , 
 n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , 
 n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , 
 n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , 
 n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , 
 n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , 
 n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , 
 n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , 
 n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , 
 n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , 
 n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , 
 n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , 
 n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , 
 n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , 
 n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , 
 n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , 
 n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , 
 n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , 
 n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , 
 n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , 
 n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , 
 n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , 
 n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , 
 n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , 
 n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , 
 n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , 
 n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , 
 n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , 
 n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , 
 n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , 
 n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , 
 n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , 
 n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , 
 n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , 
 n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , 
 n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , 
 n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , 
 n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , 
 n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , 
 n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , 
 n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , 
 n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , 
 n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , 
 n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , 
 n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , 
 n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , 
 n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , 
 n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , 
 n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , 
 n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , 
 n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , 
 n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , 
 n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , 
 n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , 
 n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , 
 n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , 
 n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , 
 n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , 
 n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , 
 n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , 
 n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , 
 n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , 
 n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , 
 n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , 
 n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , 
 n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , 
 n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , 
 n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , 
 n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , 
 n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , 
 n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , 
 n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , 
 n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , 
 n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , 
 n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , 
 n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , 
 n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , 
 n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , 
 n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , 
 n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , 
 n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , 
 n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , 
 n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , 
 n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , 
 n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , 
 n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , 
 n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , 
 n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , 
 n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , 
 n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , 
 n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , 
 n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , 
 n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , 
 n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , 
 n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , 
 n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , 
 n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , 
 n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , 
 n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , 
 n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , 
 n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , 
 n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , 
 n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , 
 n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , 
 n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , 
 n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , 
 n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , 
 n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , 
 n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , 
 n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , 
 n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , 
 n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , 
 n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , 
 n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , 
 n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , 
 n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , 
 n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , 
 n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , 
 n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , 
 n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , 
 n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , 
 n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , 
 n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , 
 n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , 
 n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , 
 n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , 
 n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , 
 n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , 
 n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , 
 n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , 
 n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , 
 n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , 
 n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , 
 n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , 
 n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , 
 n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , 
 n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , 
 n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , 
 n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , 
 n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , 
 n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , 
 n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , 
 n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , 
 n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , 
 n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , 
 n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , 
 n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , 
 n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , 
 n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , 
 n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , 
 n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , 
 n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , 
 n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , 
 n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , 
 n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , 
 n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , 
 n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , 
 n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , 
 n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , 
 n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , 
 n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , 
 n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , 
 n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , 
 n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , 
 n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , 
 n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , 
 n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , 
 n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , 
 n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , 
 n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , 
 n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , 
 n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , 
 n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , 
 n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , 
 n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , 
 n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , 
 n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , 
 n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , 
 n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , 
 n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , 
 n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , 
 n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , 
 n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , 
 n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , 
 n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , 
 n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , 
 n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , 
 n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , 
 n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , 
 n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , 
 n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , 
 n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , 
 n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , 
 n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , 
 n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , 
 n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , 
 n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , 
 n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , 
 n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , 
 n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , 
 n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , 
 n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , 
 n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , 
 n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , 
 n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , 
 n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , 
 n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , 
 n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , 
 n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , 
 n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , 
 n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , 
 n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , 
 n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , 
 n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , 
 n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , 
 n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , 
 n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , 
 n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , 
 n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , 
 n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , 
 n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , 
 n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , 
 n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , 
 n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , 
 n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , 
 n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , 
 n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , 
 n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , 
 n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , 
 n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , 
 n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , 
 n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , 
 n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , 
 n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , 
 n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , 
 n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , 
 n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , 
 n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , 
 n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , 
 n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , 
 n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , 
 n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , 
 n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , 
 n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , 
 n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , 
 n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , 
 n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , 
 n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , 
 n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , 
 n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , 
 n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , 
 n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , 
 n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , 
 n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , 
 n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , 
 n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , 
 n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , 
 n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , 
 n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , 
 n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , 
 n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , 
 n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , 
 n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , 
 n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , 
 n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , 
 n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , 
 n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , 
 n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , 
 n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , 
 n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , 
 n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , 
 n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , 
 n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , 
 n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , 
 n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , 
 n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , 
 n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , 
 n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , 
 n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , 
 n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , 
 n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , 
 n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , 
 n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , 
 n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , 
 n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , 
 n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , 
 n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , 
 n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , 
 n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , 
 n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , 
 n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , 
 n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , 
 n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , 
 n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , 
 n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , 
 n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , 
 n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , 
 n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , 
 n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , 
 n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , 
 n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , 
 n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , 
 n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , 
 n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , 
 n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , 
 n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , 
 n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , 
 n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , 
 n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , 
 n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , 
 n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , 
 n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , 
 n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , 
 n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , 
 n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , 
 n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , 
 n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , 
 n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , 
 n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , 
 n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , 
 n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , 
 n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , 
 n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , 
 n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , 
 n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , 
 n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , 
 n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , 
 n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , 
 n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , 
 n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , 
 n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , 
 n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , 
 n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , 
 n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , 
 n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , 
 n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , 
 n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , 
 n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , 
 n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , 
 n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , 
 n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , 
 n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , 
 n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , 
 n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , 
 n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , 
 n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , 
 n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , 
 n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , 
 n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , 
 n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , 
 n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , 
 n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , 
 n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , 
 n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , 
 n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , 
 n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , 
 n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , 
 n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , 
 n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , 
 n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , 
 n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , 
 n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , 
 n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , 
 n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , 
 n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , 
 n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , 
 n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , 
 n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , 
 n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , 
 n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , 
 n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , 
 n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , 
 n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , 
 n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , 
 n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , 
 n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , 
 n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , 
 n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , 
 n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , 
 n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , 
 n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , 
 n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , 
 n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , 
 n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , 
 n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , 
 n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , 
 n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , 
 n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , 
 n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , 
 n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , 
 n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , 
 n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , 
 n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , 
 n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , 
 n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , 
 n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , 
 n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , 
 n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , 
 n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , 
 n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , 
 n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , 
 n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , 
 n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , 
 n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , 
 n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , 
 n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , 
 n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , 
 n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , 
 n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , 
 n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , 
 n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , 
 n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , 
 n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , 
 n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , 
 n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , 
 n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , 
 n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , 
 n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , 
 n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , 
 n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , 
 n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , 
 n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , 
 n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , 
 n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , 
 n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , 
 n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , 
 n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , 
 n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , 
 n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , 
 n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , 
 n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , 
 n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , 
 n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , 
 n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , 
 n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , 
 n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , 
 n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , 
 n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , 
 n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , 
 n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , 
 n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , 
 n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , 
 n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , 
 n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , 
 n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , 
 n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , 
 n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , 
 n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , 
 n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , 
 n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , 
 n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , 
 n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , 
 n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , 
 n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , 
 n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , 
 n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , 
 n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , 
 n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , 
 n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , 
 n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , 
 n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , 
 n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , 
 n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , 
 n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , 
 n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , 
 n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , 
 n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , 
 n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , 
 n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , 
 n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , 
 n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , 
 n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , 
 n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , 
 n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , 
 n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , 
 n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , 
 n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , 
 n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , 
 n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , 
 n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , 
 n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , 
 n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , 
 n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , 
 n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , 
 n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , 
 n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , 
 n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , 
 n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , 
 n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , 
 n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , 
 n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , 
 n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , 
 n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , 
 n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , 
 n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , 
 n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , 
 n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , 
 n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , 
 n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , 
 n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , 
 n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , 
 n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , 
 n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , 
 n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , 
 n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , 
 n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , 
 n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , 
 n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , 
 n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , 
 n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , 
 n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , 
 n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , 
 n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , 
 n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , 
 n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , 
 n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , 
 n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , 
 n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , 
 n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , 
 n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , 
 n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , 
 n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , 
 n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , 
 n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , 
 n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , 
 n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , 
 n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , 
 n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , 
 n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , 
 n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , 
 n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , 
 n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , 
 n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , 
 n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , 
 n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , 
 n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , 
 n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , 
 n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , 
 n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , 
 n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , 
 n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , 
 n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , 
 n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , 
 n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , 
 n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , 
 n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , 
 n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , 
 n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , 
 n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , 
 n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , 
 n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , 
 n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , 
 n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , 
 n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , 
 n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , 
 n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , 
 n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , 
 n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , 
 n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , 
 n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , 
 n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , 
 n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , 
 n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , 
 n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , 
 n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , 
 n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , 
 n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , 
 n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , 
 n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , 
 n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , 
 n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , 
 n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , 
 n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , 
 n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , 
 n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , 
 n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , 
 n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , 
 n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , 
 n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , 
 n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , 
 n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , 
 n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , 
 n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , 
 n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , 
 n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , 
 n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , 
 n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , 
 n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , 
 n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , 
 n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , 
 n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , 
 n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , 
 n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , 
 n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , 
 n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , 
 n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , 
 n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , 
 n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , 
 n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , 
 n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , 
 n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , 
 n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , 
 n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , 
 n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , 
 n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , 
 n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , 
 n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , 
 n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , 
 n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , 
 n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , 
 n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , 
 n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , 
 n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , 
 n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , 
 n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , 
 n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , 
 n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , 
 n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , 
 n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , 
 n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , 
 n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , 
 n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , 
 n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , 
 n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , 
 n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , 
 n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , 
 n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , 
 n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , 
 n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , 
 n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , 
 n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , 
 n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , 
 n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , 
 n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , 
 n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , 
 n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , 
 n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , 
 n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , 
 n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , 
 n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , 
 n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , 
 n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , 
 n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , 
 n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , 
 n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , 
 n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , 
 n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , 
 n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , 
 n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , 
 n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , 
 n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , 
 n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , 
 n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , 
 n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , 
 n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , 
 n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , 
 n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , 
 n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , 
 n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , 
 n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , 
 n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , 
 n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , 
 n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , 
 n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , 
 n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , 
 n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , 
 n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , 
 n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , 
 n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , 
 n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , 
 n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , 
 n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , 
 n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , 
 n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , 
 n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , 
 n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , 
 n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , 
 n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , 
 n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , 
 n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , 
 n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , 
 n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , 
 n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , 
 n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , 
 n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , 
 n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , 
 n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , 
 n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , 
 n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , 
 n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , 
 n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , 
 n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , 
 n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , 
 n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , 
 n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , 
 n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , 
 n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , 
 n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , 
 n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , 
 n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , 
 n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , 
 n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , 
 n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , 
 n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , 
 n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , 
 n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , 
 n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , 
 n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , 
 n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , 
 n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , 
 n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , 
 n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , 
 n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , 
 n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , 
 n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , 
 n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , 
 n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , 
 n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , 
 n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , 
 n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , 
 n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , 
 n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , 
 n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , 
 n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , 
 n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , 
 n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , 
 n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , 
 n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , 
 n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , 
 n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , 
 n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , 
 n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , 
 n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , 
 n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , 
 n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , 
 n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , 
 n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , 
 n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , 
 n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , 
 n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , 
 n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , 
 n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , 
 n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , 
 n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , 
 n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , 
 n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , 
 n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , 
 n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , 
 n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , 
 n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , 
 n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , 
 n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , 
 n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , 
 n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , 
 n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , 
 n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , 
 n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , 
 n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , 
 n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , 
 n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , 
 n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , 
 n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , 
 n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , 
 n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , 
 n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , 
 n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , 
 n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , 
 n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , 
 n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , 
 n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , 
 n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , 
 n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , 
 n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , 
 n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , 
 n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , 
 n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , 
 n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , 
 n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , 
 n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , 
 n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , 
 n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , 
 n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , 
 n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , 
 n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , 
 n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , 
 n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , 
 n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , 
 n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , 
 n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , 
 n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , 
 n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , 
 n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , 
 n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , 
 n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , 
 n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , 
 n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , 
 n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , 
 n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , 
 n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , 
 n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , 
 n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , 
 n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , 
 n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , 
 n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , 
 n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , 
 n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , 
 n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , 
 n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , 
 n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , 
 n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , 
 n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , 
 n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , 
 n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , 
 n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , 
 n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , 
 n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , 
 n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , 
 n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , 
 n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , 
 n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , 
 n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , 
 n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , 
 n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , 
 n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , 
 n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , 
 n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , 
 n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , 
 n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , 
 n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , 
 n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , 
 n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , 
 n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , 
 n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , 
 n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , 
 n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , 
 n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , 
 n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , 
 n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , 
 n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , 
 n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , 
 n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , 
 n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , 
 n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , 
 n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , 
 n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , 
 n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , 
 n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , 
 n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , 
 n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , 
 n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , 
 n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , 
 n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , 
 n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , 
 n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , 
 n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , 
 n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , 
 n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , 
 n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , 
 n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , 
 n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , 
 n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , 
 n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , 
 n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , 
 n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , 
 n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , 
 n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , 
 n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , 
 n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , 
 n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , 
 n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , 
 n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , 
 n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , 
 n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , 
 n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , 
 n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , 
 n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , 
 n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , 
 n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , 
 n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , 
 n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , 
 n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , 
 n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , 
 n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , 
 n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , 
 n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , 
 n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , 
 n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , 
 n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , 
 n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , 
 n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , 
 n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , 
 n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , 
 n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , 
 n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , 
 n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , 
 n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , 
 n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , 
 n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , 
 n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , 
 n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , 
 n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , 
 n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , 
 n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , 
 n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , 
 n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , 
 n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , 
 n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , 
 n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , 
 n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , 
 n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , 
 n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , 
 n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , 
 n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , 
 n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , 
 n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , 
 n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , 
 n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , 
 n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , 
 n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , 
 n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , 
 n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , 
 n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , 
 n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , 
 n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , 
 n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , 
 n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , 
 n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , 
 n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , 
 n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , 
 n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , 
 n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , 
 n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , 
 n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , 
 n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , 
 n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , 
 n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , 
 n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , 
 n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , 
 n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , 
 n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , 
 n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , 
 n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , 
 n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , 
 n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , 
 n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , 
 n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , 
 n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , 
 n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , 
 n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , 
 n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , 
 n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , 
 n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , 
 n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , 
 n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , 
 n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , 
 n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , 
 n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , 
 n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , 
 n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , 
 n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , 
 n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , 
 n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , 
 n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , 
 n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , 
 n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , 
 n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , 
 n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , 
 n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , 
 n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , 
 n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , 
 n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , 
 n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , 
 n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , 
 n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , 
 n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , 
 n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , 
 n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , 
 n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , 
 n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , 
 n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , 
 n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , 
 n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , 
 n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , 
 n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , 
 n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , 
 n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , 
 n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , 
 n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , 
 n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , 
 n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , 
 n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , 
 n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , 
 n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , 
 n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , 
 n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , 
 n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , 
 n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , 
 n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , 
 n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , 
 n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , 
 n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , 
 n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , 
 n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , 
 n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , 
 n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , 
 n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , 
 n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , 
 n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , 
 n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , 
 n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , 
 n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , 
 n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , 
 n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , 
 n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , 
 n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , 
 n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , 
 n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , 
 n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , 
 n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , 
 n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , 
 n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , 
 n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , 
 n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , 
 n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , 
 n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , 
 n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , 
 n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , 
 n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , 
 n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , 
 n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , 
 n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , 
 n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , 
 n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , 
 n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , 
 n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , 
 n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , 
 n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , 
 n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , 
 n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , 
 n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , 
 n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , 
 n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , 
 n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , 
 n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , 
 n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , 
 n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , 
 n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , 
 n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , 
 n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , 
 n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , 
 n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , 
 n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , 
 n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , 
 n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , 
 n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , 
 n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , 
 n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , 
 n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , 
 n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , 
 n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , 
 n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , 
 n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , 
 n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , 
 n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , 
 n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , 
 n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , 
 n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , 
 n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , 
 n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , 
 n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , 
 n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , 
 n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , 
 n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , 
 n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , 
 n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , 
 n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , 
 n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , 
 n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , 
 n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , 
 n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , 
 n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , 
 n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , 
 n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , 
 n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , 
 n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , 
 n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , 
 n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , 
 n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , 
 n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , 
 n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , 
 n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , 
 n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , 
 n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , 
 n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , 
 n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , 
 n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , 
 n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , 
 n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , 
 n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , 
 n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , 
 n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , 
 n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , 
 n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , 
 n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , 
 n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , 
 n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , 
 n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , 
 n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , 
 n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , 
 n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , 
 n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , 
 n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , 
 n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , 
 n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , 
 n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , 
 n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , 
 n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , 
 n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , 
 n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , 
 n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , 
 n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , 
 n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , 
 n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , 
 n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , 
 n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , 
 n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , 
 n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , 
 n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , 
 n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , 
 n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , 
 n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , 
 n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , 
 n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , 
 n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , 
 n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , 
 n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , 
 n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , 
 n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , 
 n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , 
 n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , 
 n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , 
 n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , 
 n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , 
 n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , 
 n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , 
 n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , 
 n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , 
 n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , 
 n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , 
 n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , 
 n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , 
 n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , 
 n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , 
 n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , 
 n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , 
 n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , 
 n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , 
 n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , 
 n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , 
 n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , 
 n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , 
 n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , 
 n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , 
 n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , 
 n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , 
 n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , 
 n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , 
 n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , 
 n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , 
 n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , 
 n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , 
 n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , 
 n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , 
 n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , 
 n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , 
 n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , 
 n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , 
 n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , 
 n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , 
 n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , 
 n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , 
 n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , 
 n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , 
 n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , 
 n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , 
 n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , 
 n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , 
 n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , 
 n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , 
 n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , 
 n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , 
 n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , 
 n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , 
 n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , 
 n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , 
 n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , 
 n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , 
 n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , 
 n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , 
 n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , 
 n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , 
 n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , 
 n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , 
 n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , 
 n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , 
 n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , 
 n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , 
 n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , 
 n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , 
 n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , 
 n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , 
 n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , 
 n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , 
 n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , 
 n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , 
 n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , 
 n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , 
 n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , 
 n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , 
 n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , 
 n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , 
 n14641 , n14642 , n14643 , n14644 , n14645 , C0n , C0 , C1n , C1 ;
buf ( n370 , n0 );
buf ( n371 , n1 );
buf ( n372 , n2 );
buf ( n373 , n3 );
buf ( n374 , n4 );
buf ( n375 , n5 );
buf ( n376 , n6 );
buf ( n377 , n7 );
buf ( n378 , n8 );
buf ( n379 , n9 );
buf ( n380 , n10 );
buf ( n381 , n11 );
buf ( n382 , n12 );
buf ( n383 , n13 );
buf ( n384 , n14 );
buf ( n385 , n15 );
buf ( n386 , n16 );
buf ( n387 , n17 );
buf ( n388 , n18 );
buf ( n389 , n19 );
buf ( n390 , n20 );
buf ( n391 , n21 );
buf ( n392 , n22 );
buf ( n393 , n23 );
buf ( n394 , n24 );
buf ( n395 , n25 );
buf ( n396 , n26 );
buf ( n397 , n27 );
buf ( n398 , n28 );
buf ( n399 , n29 );
buf ( n400 , n30 );
buf ( n401 , n31 );
buf ( n402 , n32 );
buf ( n403 , n33 );
buf ( n404 , n34 );
buf ( n405 , n35 );
buf ( n406 , n36 );
buf ( n407 , n37 );
buf ( n408 , n38 );
buf ( n409 , n39 );
buf ( n410 , n40 );
buf ( n411 , n41 );
buf ( n412 , n42 );
buf ( n413 , n43 );
buf ( n414 , n44 );
buf ( n415 , n45 );
buf ( n416 , n46 );
buf ( n417 , n47 );
buf ( n418 , n48 );
buf ( n419 , n49 );
buf ( n420 , n50 );
buf ( n421 , n51 );
buf ( n422 , n52 );
buf ( n423 , n53 );
buf ( n424 , n54 );
buf ( n425 , n55 );
buf ( n56 , n426 );
buf ( n57 , n427 );
buf ( n58 , n428 );
buf ( n59 , n429 );
buf ( n60 , n430 );
buf ( n61 , n431 );
buf ( n62 , n432 );
buf ( n63 , n433 );
buf ( n64 , n434 );
buf ( n65 , n435 );
buf ( n66 , n436 );
buf ( n67 , n437 );
buf ( n68 , n438 );
buf ( n69 , n439 );
buf ( n70 , n440 );
buf ( n71 , n441 );
buf ( n72 , n442 );
buf ( n73 , n443 );
buf ( n74 , n444 );
buf ( n75 , n445 );
buf ( n76 , n446 );
buf ( n77 , n447 );
buf ( n78 , n448 );
buf ( n79 , n449 );
buf ( n80 , n450 );
buf ( n81 , n451 );
buf ( n82 , n452 );
buf ( n83 , n453 );
buf ( n84 , n454 );
buf ( n85 , n455 );
buf ( n86 , n456 );
buf ( n87 , n457 );
buf ( n88 , n458 );
buf ( n89 , n459 );
buf ( n90 , n460 );
buf ( n91 , n461 );
buf ( n92 , n462 );
buf ( n93 , n463 );
buf ( n94 , n464 );
buf ( n95 , n465 );
buf ( n96 , n466 );
buf ( n97 , n467 );
buf ( n98 , n468 );
buf ( n99 , n469 );
buf ( n100 , n470 );
buf ( n101 , n471 );
buf ( n102 , n472 );
buf ( n103 , n473 );
buf ( n104 , n474 );
buf ( n105 , n475 );
buf ( n106 , n476 );
buf ( n107 , n477 );
buf ( n108 , n478 );
buf ( n109 , n479 );
buf ( n110 , n480 );
buf ( n111 , n481 );
buf ( n112 , n482 );
buf ( n113 , n483 );
buf ( n114 , n484 );
buf ( n115 , n485 );
buf ( n116 , n486 );
buf ( n117 , n487 );
buf ( n118 , n488 );
buf ( n119 , n489 );
buf ( n120 , n490 );
buf ( n121 , n491 );
buf ( n122 , n492 );
buf ( n123 , n493 );
buf ( n124 , n494 );
buf ( n125 , n495 );
buf ( n126 , n496 );
buf ( n127 , n497 );
buf ( n128 , n498 );
buf ( n129 , n499 );
buf ( n130 , n500 );
buf ( n131 , n501 );
buf ( n132 , n502 );
buf ( n133 , n503 );
buf ( n134 , n504 );
buf ( n135 , n505 );
buf ( n136 , n506 );
buf ( n137 , n507 );
buf ( n138 , n508 );
buf ( n139 , n509 );
buf ( n140 , n510 );
buf ( n141 , n511 );
buf ( n142 , n512 );
buf ( n143 , n513 );
buf ( n144 , n514 );
buf ( n145 , n515 );
buf ( n146 , n516 );
buf ( n147 , n517 );
buf ( n148 , n518 );
buf ( n149 , n519 );
buf ( n150 , n520 );
buf ( n151 , n521 );
buf ( n152 , n522 );
buf ( n153 , n523 );
buf ( n154 , n524 );
buf ( n155 , n525 );
buf ( n156 , n526 );
buf ( n157 , n527 );
buf ( n158 , n528 );
buf ( n159 , n529 );
buf ( n160 , n530 );
buf ( n161 , n531 );
buf ( n162 , n532 );
buf ( n163 , n533 );
buf ( n164 , n534 );
buf ( n165 , n535 );
buf ( n166 , n536 );
buf ( n167 , n537 );
buf ( n168 , n538 );
buf ( n169 , n539 );
buf ( n170 , n540 );
buf ( n171 , n541 );
buf ( n172 , n542 );
buf ( n173 , n543 );
buf ( n174 , n544 );
buf ( n175 , n545 );
buf ( n176 , n546 );
buf ( n177 , n547 );
buf ( n178 , n548 );
buf ( n179 , n549 );
buf ( n180 , n550 );
buf ( n181 , n551 );
buf ( n182 , n552 );
buf ( n183 , n553 );
buf ( n184 , n554 );
buf ( n426 , C0 );
buf ( n427 , C0 );
buf ( n428 , C0 );
buf ( n429 , C0 );
buf ( n430 , C0 );
buf ( n431 , C0 );
buf ( n432 , C0 );
buf ( n433 , C0 );
buf ( n434 , C0 );
buf ( n435 , C0 );
buf ( n436 , C0 );
buf ( n437 , C0 );
buf ( n438 , C0 );
buf ( n439 , C0 );
buf ( n440 , C0 );
buf ( n441 , C0 );
buf ( n442 , C0 );
buf ( n443 , C0 );
buf ( n444 , C0 );
buf ( n445 , C0 );
buf ( n446 , C0 );
buf ( n447 , C0 );
buf ( n448 , C0 );
buf ( n449 , C0 );
buf ( n450 , C0 );
buf ( n451 , C0 );
buf ( n452 , C0 );
buf ( n453 , C0 );
buf ( n454 , C0 );
buf ( n455 , C0 );
buf ( n456 , C0 );
buf ( n457 , C0 );
buf ( n458 , C0 );
buf ( n459 , C0 );
buf ( n460 , C0 );
buf ( n461 , C0 );
buf ( n462 , C0 );
buf ( n463 , C0 );
buf ( n464 , C0 );
buf ( n465 , C0 );
buf ( n466 , C0 );
buf ( n467 , C0 );
buf ( n468 , C0 );
buf ( n469 , C0 );
buf ( n470 , C0 );
buf ( n471 , C0 );
buf ( n472 , C0 );
buf ( n473 , C0 );
buf ( n474 , C0 );
buf ( n475 , C0 );
buf ( n476 , C0 );
buf ( n477 , C0 );
buf ( n478 , C0 );
buf ( n479 , C0 );
buf ( n480 , C0 );
buf ( n481 , C0 );
buf ( n482 , C0 );
buf ( n483 , C0 );
buf ( n484 , C0 );
buf ( n485 , C0 );
buf ( n486 , C0 );
buf ( n487 , C0 );
buf ( n488 , C0 );
buf ( n489 , C0 );
buf ( n490 , n14587 );
buf ( n491 , n14555 );
buf ( n492 , n14566 );
buf ( n493 , n14512 );
buf ( n494 , n14640 );
buf ( n495 , n14498 );
buf ( n496 , n14078 );
buf ( n497 , n14614 );
buf ( n498 , n14600 );
buf ( n499 , n14641 );
buf ( n500 , n14641 );
buf ( n501 , n14641 );
buf ( n502 , n14641 );
buf ( n503 , n14641 );
buf ( n504 , n14641 );
buf ( n505 , n14641 );
buf ( n506 , n14562 );
buf ( n507 , n14562 );
buf ( n508 , n14562 );
buf ( n509 , n14562 );
buf ( n510 , n14562 );
buf ( n511 , n14562 );
buf ( n512 , n14562 );
buf ( n513 , n14562 );
buf ( n514 , n14562 );
buf ( n515 , n14562 );
buf ( n516 , n14562 );
buf ( n517 , n14562 );
buf ( n518 , n14563 );
buf ( n519 , n14563 );
buf ( n520 , n14563 );
buf ( n521 , n14563 );
buf ( n522 , n14563 );
buf ( n523 , n14563 );
buf ( n524 , n14563 );
buf ( n525 , n14563 );
buf ( n526 , n14563 );
buf ( n527 , n14563 );
buf ( n528 , n14563 );
buf ( n529 , n14563 );
buf ( n530 , n13586 );
buf ( n531 , n14579 );
buf ( n532 , n14620 );
buf ( n533 , n13635 );
buf ( n534 , n13650 );
buf ( n535 , n14099 );
buf ( n536 , n14136 );
buf ( n537 , n14551 );
buf ( n538 , n14121 );
buf ( n539 , n14199 );
buf ( n540 , n14645 );
buf ( n541 , n14179 );
buf ( n542 , n14606 );
buf ( n543 , n14591 );
buf ( n544 , n14226 );
buf ( n545 , n14250 );
buf ( n546 , n14261 );
buf ( n547 , n14489 );
buf ( n548 , n14435 );
buf ( n549 , n14473 );
buf ( n550 , n14477 );
buf ( n551 , n14537 );
buf ( n552 , n14466 );
buf ( n553 , n14469 );
buf ( n554 , n14630 );
not ( n555 , n370 );
nand ( n556 , n370 , n374 );
not ( n557 , n556 );
nand ( n558 , n371 , n373 );
not ( n559 , n558 );
or ( n560 , n557 , n559 );
and ( n561 , n370 , n375 );
xor ( n562 , n372 , n561 );
and ( n563 , n372 , n373 );
and ( n564 , n562 , n563 );
and ( n565 , n372 , n561 );
or ( n566 , n564 , n565 );
nand ( n567 , n560 , n566 );
nand ( n568 , n370 , n373 );
nand ( n569 , n371 , n372 );
xor ( n570 , n568 , n569 );
not ( n571 , n371 );
xor ( n572 , n570 , n571 );
not ( n573 , n556 );
not ( n574 , n558 );
nand ( n575 , n573 , n574 );
nand ( n576 , n567 , n572 , n575 );
nand ( n577 , n568 , n569 );
nand ( n578 , n568 , n571 );
nand ( n579 , n569 , n571 );
nand ( n580 , n577 , n578 , n579 );
nand ( n581 , n370 , n372 );
nand ( n582 , n580 , n581 );
nand ( n583 , n576 , n582 );
nor ( n584 , n555 , n583 );
not ( n585 , n584 );
nand ( n586 , n371 , n374 );
not ( n587 , n586 );
xor ( n588 , n372 , n561 );
xor ( n589 , n588 , n563 );
not ( n590 , n589 );
not ( n591 , n590 );
or ( n592 , n587 , n591 );
nand ( n593 , n370 , n376 );
not ( n594 , n593 );
not ( n595 , n594 );
nand ( n596 , n371 , n375 );
not ( n597 , n596 );
not ( n598 , n597 );
or ( n599 , n595 , n598 );
not ( n600 , n596 );
not ( n601 , n593 );
or ( n602 , n600 , n601 );
and ( n603 , n372 , n374 );
nand ( n604 , n602 , n603 );
nand ( n605 , n599 , n604 );
nand ( n606 , n592 , n605 );
not ( n607 , n586 );
nand ( n608 , n589 , n607 );
and ( n609 , n606 , n608 );
not ( n610 , n574 );
not ( n611 , n556 );
and ( n612 , n610 , n611 );
and ( n613 , n556 , n574 );
nor ( n614 , n612 , n613 );
xor ( n615 , n566 , n614 );
nand ( n616 , n609 , n615 );
not ( n617 , n616 );
nand ( n618 , n373 , n374 );
not ( n619 , n618 );
not ( n620 , n370 );
not ( n621 , n377 );
or ( n622 , n620 , n621 );
nand ( n623 , n371 , n376 );
nand ( n624 , n622 , n623 );
not ( n625 , n624 );
and ( n626 , n372 , n375 );
not ( n627 , n626 );
or ( n628 , n625 , n627 );
nand ( n629 , n371 , n376 , n370 , n377 );
nand ( n630 , n628 , n629 );
nor ( n631 , n619 , n630 );
nand ( n632 , n372 , n374 );
nand ( n633 , n371 , n375 );
nand ( n634 , n370 , n376 );
and ( n635 , n633 , n634 );
not ( n636 , n633 );
and ( n637 , n636 , n594 );
nor ( n638 , n635 , n637 );
xor ( n639 , n632 , n638 );
or ( n640 , n631 , n639 );
not ( n641 , n618 );
nand ( n642 , n641 , n630 );
nand ( n643 , n640 , n642 );
not ( n644 , n643 );
not ( n645 , n644 );
xor ( n646 , n607 , n605 );
xnor ( n647 , n646 , n589 );
not ( n648 , n647 );
or ( n649 , n645 , n648 );
nand ( n650 , n373 , n375 , n372 , n376 );
not ( n651 , n650 );
nand ( n652 , n618 , n373 );
not ( n653 , n652 );
and ( n654 , n651 , n653 );
nand ( n655 , n372 , n375 );
nand ( n656 , n371 , n376 );
and ( n657 , n655 , n656 );
not ( n658 , n655 );
not ( n659 , n623 );
and ( n660 , n658 , n659 );
nor ( n661 , n657 , n660 );
and ( n662 , n370 , n377 );
xor ( n663 , n661 , n662 );
nand ( n664 , n652 , n650 );
and ( n665 , n663 , n664 );
nor ( n666 , n654 , n665 );
xor ( n667 , n618 , n630 );
xnor ( n668 , n667 , n639 );
nand ( n669 , n666 , n668 );
nand ( n670 , n649 , n669 );
not ( n671 , n670 );
not ( n672 , n671 );
not ( n673 , n663 );
not ( n674 , n650 );
not ( n675 , n374 );
not ( n676 , n373 );
or ( n677 , n675 , n676 );
nand ( n678 , n677 , n373 );
not ( n679 , n678 );
or ( n680 , n674 , n679 );
or ( n681 , n678 , n650 );
nand ( n682 , n680 , n681 );
not ( n683 , n682 );
and ( n684 , n673 , n683 );
and ( n685 , n682 , n663 );
nor ( n686 , n684 , n685 );
nand ( n687 , n374 , n375 );
nand ( n688 , n371 , n377 );
xor ( n689 , n687 , n688 );
nand ( n690 , n373 , n375 );
nand ( n691 , n376 , n372 );
xnor ( n692 , n690 , n691 );
and ( n693 , n689 , n692 );
and ( n694 , n687 , n688 );
or ( n695 , n693 , n694 );
nand ( n696 , n686 , n695 );
not ( n697 , n696 );
xor ( n698 , n687 , n688 );
xor ( n699 , n698 , n692 );
nand ( n700 , n372 , n377 );
not ( n701 , n700 );
nand ( n702 , n373 , n376 );
not ( n703 , n702 );
and ( n704 , n701 , n703 );
nand ( n705 , n700 , n702 );
not ( n706 , n375 );
and ( n707 , n706 , n374 );
and ( n708 , n705 , n707 );
nor ( n709 , n704 , n708 );
nand ( n710 , n699 , n709 );
not ( n711 , n710 );
nand ( n712 , n377 , n374 , n375 );
not ( n713 , n712 );
nand ( n714 , n375 , n377 );
nand ( n715 , n377 , n376 );
nor ( n716 , n714 , n715 );
nand ( n717 , n713 , n716 );
nand ( n718 , n374 , n376 );
not ( n719 , n718 );
nand ( n720 , n373 , n377 );
not ( n721 , n720 );
or ( n722 , n719 , n721 );
nand ( n723 , n374 , n376 );
nand ( n724 , n373 , n377 );
or ( n725 , n723 , n724 );
nand ( n726 , n722 , n725 );
nand ( n727 , n726 , n712 );
and ( n728 , n374 , n377 );
nand ( n729 , n375 , n376 );
nor ( n730 , n728 , n729 );
and ( n731 , n727 , n730 );
nor ( n732 , n712 , n726 );
nor ( n733 , n731 , n732 );
nand ( n734 , n717 , n733 );
not ( n735 , n734 );
or ( n736 , n700 , n702 );
not ( n737 , n373 );
not ( n738 , n376 );
or ( n739 , n737 , n738 );
nand ( n740 , n372 , n377 );
nand ( n741 , n739 , n740 );
nand ( n742 , n736 , n741 );
not ( n743 , n742 );
not ( n744 , n707 );
and ( n745 , n743 , n744 );
and ( n746 , n707 , n742 );
nor ( n747 , n745 , n746 );
not ( n748 , n618 );
and ( n749 , n377 , n376 );
nand ( n750 , n748 , n749 );
nand ( n751 , n747 , n750 );
not ( n752 , n751 );
or ( n753 , n735 , n752 );
not ( n754 , n747 );
not ( n755 , n750 );
nand ( n756 , n754 , n755 );
nand ( n757 , n753 , n756 );
not ( n758 , n757 );
or ( n759 , n711 , n758 );
or ( n760 , n699 , n709 );
nand ( n761 , n759 , n760 );
not ( n762 , n761 );
or ( n763 , n697 , n762 );
not ( n764 , n686 );
not ( n765 , n695 );
nand ( n766 , n764 , n765 );
nand ( n767 , n763 , n766 );
not ( n768 , n767 );
or ( n769 , n672 , n768 );
not ( n770 , n647 );
not ( n771 , n644 );
and ( n772 , n770 , n771 );
nand ( n773 , n647 , n644 );
nor ( n774 , n666 , n668 );
and ( n775 , n773 , n774 );
nor ( n776 , n772 , n775 );
nand ( n777 , n769 , n776 );
not ( n778 , n777 );
or ( n779 , n617 , n778 );
nor ( n780 , n615 , n609 );
not ( n781 , n780 );
nand ( n782 , n779 , n781 );
not ( n783 , n782 );
or ( n784 , n585 , n783 );
not ( n785 , n575 );
not ( n786 , n567 );
or ( n787 , n785 , n786 );
not ( n788 , n572 );
nand ( n789 , n787 , n788 );
not ( n790 , n582 );
or ( n791 , n789 , n790 );
or ( n792 , n580 , n581 );
nand ( n793 , n791 , n792 );
or ( n794 , n793 , n371 );
nand ( n795 , n794 , n370 );
nand ( n796 , n784 , n795 );
buf ( n797 , n796 );
and ( n798 , n715 , n376 );
buf ( n799 , n798 );
and ( n800 , n797 , n799 );
buf ( n801 , n800 );
buf ( n802 , n801 );
buf ( n803 , n767 );
buf ( n804 , n803 );
not ( n805 , n774 );
buf ( n806 , n669 );
nand ( n807 , n805 , n806 );
not ( n808 , n807 );
and ( n809 , n804 , n808 );
not ( n810 , n804 );
and ( n811 , n810 , n807 );
nor ( n812 , n809 , n811 );
buf ( n813 , n812 );
buf ( n814 , n813 );
buf ( n815 , n814 );
buf ( n816 , n815 );
and ( n817 , n802 , n816 );
not ( n818 , n802 );
buf ( n819 , n815 );
not ( n820 , n819 );
buf ( n821 , n820 );
buf ( n822 , n821 );
and ( n823 , n818 , n822 );
nor ( n824 , n817 , n823 );
buf ( n825 , n824 );
not ( n826 , n790 );
nand ( n827 , n826 , n792 );
not ( n828 , n827 );
not ( n829 , n616 );
not ( n830 , n576 );
nor ( n831 , n829 , n830 );
not ( n832 , n831 );
buf ( n833 , n777 );
not ( n834 , n833 );
or ( n835 , n832 , n834 );
and ( n836 , n780 , n576 );
not ( n837 , n789 );
nor ( n838 , n836 , n837 );
nand ( n839 , n835 , n838 );
not ( n840 , n839 );
or ( n841 , n828 , n840 );
or ( n842 , n827 , n839 );
nand ( n843 , n841 , n842 );
buf ( n844 , n843 );
not ( n845 , n844 );
buf ( n846 , n845 );
buf ( n847 , n846 );
not ( n848 , n847 );
buf ( n849 , n848 );
and ( n850 , n714 , n749 );
not ( n851 , n714 );
and ( n852 , n851 , n715 );
or ( n853 , n850 , n852 );
nand ( n854 , n849 , n853 );
buf ( n855 , n854 );
nand ( n856 , n571 , n370 );
not ( n857 , n856 );
not ( n858 , n857 );
nor ( n859 , n829 , n583 );
not ( n860 , n859 );
not ( n861 , n777 );
or ( n862 , n860 , n861 );
not ( n863 , n781 );
not ( n864 , n583 );
and ( n865 , n863 , n864 );
nor ( n866 , n865 , n793 );
nand ( n867 , n862 , n866 );
not ( n868 , n867 );
not ( n869 , n868 );
or ( n870 , n858 , n869 );
nand ( n871 , n867 , n856 );
nand ( n872 , n870 , n871 );
buf ( n873 , n872 );
not ( n874 , n873 );
buf ( n875 , n874 );
buf ( n876 , n875 );
not ( n877 , n876 );
buf ( n878 , n877 );
buf ( n879 , n878 );
buf ( n880 , n798 );
and ( n881 , n879 , n880 );
xor ( n882 , n699 , n709 );
xor ( n883 , n882 , n757 );
nand ( n884 , n812 , n883 );
buf ( n885 , n884 );
not ( n886 , n885 );
buf ( n887 , n886 );
buf ( n888 , n887 );
nor ( n889 , n881 , n888 );
buf ( n890 , n889 );
buf ( n891 , n890 );
or ( n892 , n855 , n891 );
buf ( n893 , n878 );
buf ( n894 , n887 );
buf ( n895 , n798 );
nand ( n896 , n893 , n894 , n895 );
buf ( n897 , n896 );
buf ( n898 , n897 );
nand ( n899 , n892 , n898 );
buf ( n900 , n899 );
buf ( n901 , n900 );
not ( n902 , n901 );
buf ( n903 , n902 );
xor ( n904 , n825 , n903 );
not ( n905 , n830 );
nand ( n906 , n905 , n789 );
xnor ( n907 , n782 , n906 );
buf ( n908 , n907 );
not ( n909 , n730 );
nand ( n910 , n374 , n377 );
xor ( n911 , n910 , n375 );
nand ( n912 , n911 , n729 );
nand ( n913 , n909 , n912 );
and ( n914 , n913 , n716 );
not ( n915 , n913 );
not ( n916 , n716 );
and ( n917 , n915 , n916 );
or ( n918 , n914 , n917 );
nand ( n919 , n908 , n918 );
buf ( n920 , n919 );
not ( n921 , n920 );
not ( n922 , n829 );
nand ( n923 , n922 , n781 );
not ( n924 , n923 );
not ( n925 , n924 );
not ( n926 , n833 );
not ( n927 , n926 );
or ( n928 , n925 , n927 );
nand ( n929 , n833 , n923 );
nand ( n930 , n928 , n929 );
buf ( n931 , n930 );
not ( n932 , n931 );
buf ( n933 , n932 );
buf ( n934 , n933 );
not ( n935 , n934 );
buf ( n936 , n935 );
not ( n937 , n912 );
not ( n938 , n716 );
or ( n939 , n937 , n938 );
nand ( n940 , n939 , n909 );
not ( n941 , n940 );
not ( n942 , n941 );
not ( n943 , n732 );
nand ( n944 , n943 , n727 );
not ( n945 , n944 );
not ( n946 , n945 );
or ( n947 , n942 , n946 );
nand ( n948 , n944 , n940 );
nand ( n949 , n947 , n948 );
nand ( n950 , n936 , n949 );
buf ( n951 , n950 );
not ( n952 , n951 );
or ( n953 , n921 , n952 );
not ( n954 , n806 );
not ( n955 , n803 );
or ( n956 , n954 , n955 );
not ( n957 , n774 );
nand ( n958 , n956 , n957 );
not ( n959 , n958 );
and ( n960 , n647 , n643 );
not ( n961 , n647 );
and ( n962 , n961 , n644 );
nor ( n963 , n960 , n962 );
not ( n964 , n963 );
and ( n965 , n959 , n964 );
and ( n966 , n958 , n963 );
nor ( n967 , n965 , n966 );
not ( n968 , n967 );
nand ( n969 , n756 , n751 );
xnor ( n970 , n734 , n969 );
buf ( n971 , n970 );
buf ( n972 , n971 );
buf ( n973 , n972 );
nand ( n974 , n968 , n973 );
buf ( n975 , n974 );
not ( n976 , n975 );
buf ( n977 , n976 );
buf ( n978 , n977 );
nand ( n979 , n953 , n978 );
buf ( n980 , n979 );
buf ( n981 , n980 );
not ( n982 , n919 );
not ( n983 , n950 );
nand ( n984 , n982 , n983 );
buf ( n985 , n984 );
nand ( n986 , n981 , n985 );
buf ( n987 , n986 );
xnor ( n988 , n904 , n987 );
buf ( n989 , n988 );
not ( n990 , n919 );
and ( n991 , n974 , n990 );
not ( n992 , n974 );
and ( n993 , n992 , n919 );
nor ( n994 , n991 , n993 );
xor ( n995 , n983 , n994 );
buf ( n996 , n995 );
not ( n997 , n996 );
nand ( n998 , n878 , n798 );
xor ( n999 , n884 , n998 );
xnor ( n1000 , n999 , n854 );
not ( n1001 , n1000 );
buf ( n1002 , n1001 );
not ( n1003 , n1002 );
or ( n1004 , n997 , n1003 );
buf ( n1005 , n796 );
buf ( n1006 , n1005 );
buf ( n1007 , n1006 );
buf ( n1008 , n1007 );
buf ( n1009 , n377 );
nand ( n1010 , n1008 , n1009 );
buf ( n1011 , n1010 );
and ( n1012 , n764 , n765 );
not ( n1013 , n764 );
and ( n1014 , n1013 , n695 );
nor ( n1015 , n1012 , n1014 );
not ( n1016 , n1015 );
buf ( n1017 , n761 );
not ( n1018 , n1017 );
not ( n1019 , n1018 );
or ( n1020 , n1016 , n1019 );
not ( n1021 , n1015 );
nand ( n1022 , n1021 , n1017 );
nand ( n1023 , n1020 , n1022 );
buf ( n1024 , n1023 );
buf ( n1025 , n1024 );
buf ( n1026 , n1025 );
and ( n1027 , n1011 , n1026 );
not ( n1028 , n1011 );
buf ( n1029 , n1026 );
not ( n1030 , n1029 );
buf ( n1031 , n1030 );
and ( n1032 , n1028 , n1031 );
nor ( n1033 , n1027 , n1032 );
and ( n1034 , n1023 , n973 );
not ( n1035 , n857 );
not ( n1036 , n868 );
or ( n1037 , n1035 , n1036 );
nand ( n1038 , n1037 , n871 );
buf ( n1039 , n1038 );
nand ( n1040 , n1034 , n377 , n1039 );
nand ( n1041 , n1033 , n1040 );
not ( n1042 , n1041 );
buf ( n1043 , n968 );
not ( n1044 , n1043 );
buf ( n1045 , n918 );
not ( n1046 , n1045 );
buf ( n1047 , n1046 );
buf ( n1048 , n1047 );
nor ( n1049 , n1044 , n1048 );
buf ( n1050 , n1049 );
buf ( n1051 , n1050 );
buf ( n1052 , n936 );
buf ( n1053 , n853 );
and ( n1054 , n1052 , n1053 );
buf ( n1055 , n1054 );
buf ( n1056 , n1055 );
buf ( n1057 , n908 );
buf ( n1058 , n798 );
and ( n1059 , n1057 , n1058 );
buf ( n1060 , n1059 );
buf ( n1061 , n1060 );
and ( n1062 , n1051 , n1056 );
or ( n1063 , C0 , n1062 );
buf ( n1064 , n1063 );
not ( n1065 , n1064 );
or ( n1066 , n1042 , n1065 );
not ( n1067 , n1033 );
not ( n1068 , n1040 );
nand ( n1069 , n1067 , n1068 );
nand ( n1070 , n1066 , n1069 );
buf ( n1071 , n1070 );
nand ( n1072 , n1004 , n1071 );
buf ( n1073 , n1072 );
buf ( n1074 , n1073 );
not ( n1075 , n995 );
nand ( n1076 , n1075 , n1000 );
buf ( n1077 , n1076 );
nand ( n1078 , n1074 , n1077 );
buf ( n1079 , n1078 );
buf ( n1080 , n1079 );
buf ( n1081 , n812 );
not ( n1082 , n1015 );
not ( n1083 , n1018 );
or ( n1084 , n1082 , n1083 );
nand ( n1085 , n1084 , n1022 );
buf ( n1086 , n1085 );
nand ( n1087 , n1081 , n1086 );
buf ( n1088 , n1087 );
and ( n1089 , n968 , n883 );
xor ( n1090 , n1088 , n1089 );
buf ( n1091 , n949 );
buf ( n1092 , n908 );
nand ( n1093 , n1091 , n1092 );
buf ( n1094 , n1093 );
xnor ( n1095 , n1090 , n1094 );
not ( n1096 , n1095 );
buf ( n1097 , n843 );
buf ( n1098 , n918 );
and ( n1099 , n1097 , n1098 );
buf ( n1100 , n1099 );
buf ( n1101 , n933 );
not ( n1102 , n1101 );
buf ( n1103 , n1102 );
buf ( n1104 , n1103 );
buf ( n1105 , n970 );
and ( n1106 , n1104 , n1105 );
buf ( n1107 , n1106 );
xor ( n1108 , n1100 , n1107 );
buf ( n1109 , n1038 );
buf ( n1110 , n853 );
and ( n1111 , n1109 , n1110 );
buf ( n1112 , n1111 );
xor ( n1113 , n1108 , n1112 );
not ( n1114 , n1113 );
or ( n1115 , n1096 , n1114 );
or ( n1116 , n1113 , n1095 );
nand ( n1117 , n1115 , n1116 );
buf ( n1118 , n1085 );
buf ( n1119 , n883 );
nand ( n1120 , n1118 , n1119 );
buf ( n1121 , n1120 );
buf ( n1122 , n1121 );
not ( n1123 , n1122 );
buf ( n1124 , n968 );
buf ( n1125 , n949 );
nand ( n1126 , n1124 , n1125 );
buf ( n1127 , n1126 );
buf ( n1128 , n1127 );
not ( n1129 , n1128 );
or ( n1130 , n1123 , n1129 );
buf ( n1131 , n812 );
buf ( n1132 , n973 );
and ( n1133 , n1131 , n1132 );
buf ( n1134 , n1133 );
buf ( n1135 , n1134 );
nand ( n1136 , n1130 , n1135 );
buf ( n1137 , n1136 );
buf ( n1138 , n1137 );
buf ( n1139 , n1127 );
not ( n1140 , n1139 );
buf ( n1141 , n1121 );
not ( n1142 , n1141 );
buf ( n1143 , n1142 );
buf ( n1144 , n1143 );
nand ( n1145 , n1140 , n1144 );
buf ( n1146 , n1145 );
buf ( n1147 , n1146 );
nand ( n1148 , n1138 , n1147 );
buf ( n1149 , n1148 );
buf ( n1150 , n1149 );
buf ( n1151 , n1007 );
buf ( n1152 , n1026 );
buf ( n1153 , n377 );
and ( n1154 , n1151 , n1152 , n1153 );
buf ( n1155 , n1154 );
buf ( n1156 , n1155 );
xor ( n1157 , n1150 , n1156 );
buf ( n1158 , n908 );
buf ( n1159 , n853 );
nand ( n1160 , n1158 , n1159 );
buf ( n1161 , n1160 );
buf ( n1162 , n1161 );
not ( n1163 , n1162 );
buf ( n1164 , n1163 );
buf ( n1165 , n1164 );
not ( n1166 , n1165 );
buf ( n1167 , n936 );
buf ( n1168 , n918 );
and ( n1169 , n1167 , n1168 );
buf ( n1170 , n1169 );
buf ( n1171 , n1170 );
not ( n1172 , n1171 );
or ( n1173 , n1166 , n1172 );
buf ( n1174 , n798 );
not ( n1175 , n1174 );
buf ( n1176 , n1175 );
buf ( n1177 , C1 );
buf ( n1178 , n1177 );
nand ( n1179 , n1173 , n1178 );
buf ( n1180 , n1179 );
buf ( n1181 , n1180 );
and ( n1182 , n1157 , n1181 );
and ( n1183 , n1150 , n1156 );
or ( n1184 , n1182 , n1183 );
buf ( n1185 , n1184 );
xor ( n1186 , n1117 , n1185 );
buf ( n1187 , n1186 );
xor ( n1188 , n989 , n1080 );
xor ( n1189 , n1188 , n1187 );
buf ( n1190 , n1189 );
xor ( n1191 , n989 , n1080 );
and ( n1192 , n1191 , n1187 );
and ( n1193 , n989 , n1080 );
or ( n1194 , n1192 , n1193 );
buf ( n1195 , n1194 );
and ( n1196 , n815 , n1007 , n798 );
not ( n1197 , n1088 );
nand ( n1198 , n1197 , n1089 );
not ( n1199 , n1198 );
not ( n1200 , n1094 );
or ( n1201 , n1199 , n1200 );
not ( n1202 , n1089 );
nand ( n1203 , n1202 , n1088 );
nand ( n1204 , n1201 , n1203 );
xor ( n1205 , n1196 , n1204 );
xor ( n1206 , n1100 , n1107 );
and ( n1207 , n1206 , n1112 );
and ( n1208 , n1100 , n1107 );
or ( n1209 , n1207 , n1208 );
xnor ( n1210 , n1205 , n1209 );
buf ( n1211 , n1210 );
not ( n1212 , n1113 );
nand ( n1213 , n1212 , n1095 );
buf ( n1214 , n1213 );
not ( n1215 , n1214 );
buf ( n1216 , n1185 );
not ( n1217 , n1216 );
or ( n1218 , n1215 , n1217 );
not ( n1219 , n1095 );
nand ( n1220 , n1219 , n1113 );
buf ( n1221 , n1220 );
nand ( n1222 , n1218 , n1221 );
buf ( n1223 , n1222 );
buf ( n1224 , n1223 );
not ( n1225 , n825 );
nand ( n1226 , n1225 , n903 );
not ( n1227 , n1226 );
not ( n1228 , n987 );
or ( n1229 , n1227 , n1228 );
not ( n1230 , n903 );
nand ( n1231 , n1230 , n825 );
nand ( n1232 , n1229 , n1231 );
buf ( n1233 , n1103 );
buf ( n1234 , n883 );
and ( n1235 , n1233 , n1234 );
buf ( n1236 , n1235 );
buf ( n1237 , n872 );
buf ( n1238 , n918 );
and ( n1239 , n1237 , n1238 );
buf ( n1240 , n1239 );
xor ( n1241 , n1236 , n1240 );
buf ( n1242 , n843 );
buf ( n1243 , n949 );
and ( n1244 , n1242 , n1243 );
buf ( n1245 , n1244 );
xor ( n1246 , n1241 , n1245 );
buf ( n1247 , n1246 );
buf ( n1248 , n968 );
buf ( n1249 , n1085 );
and ( n1250 , n1248 , n1249 );
buf ( n1251 , n1250 );
buf ( n1252 , n1251 );
not ( n1253 , n795 );
nand ( n1254 , n782 , n584 );
not ( n1255 , n1254 );
or ( n1256 , n1253 , n1255 );
nand ( n1257 , n1256 , n853 );
not ( n1258 , n1257 );
buf ( n1259 , n1258 );
xor ( n1260 , n1252 , n1259 );
buf ( n1261 , n908 );
buf ( n1262 , n973 );
and ( n1263 , n1261 , n1262 );
buf ( n1264 , n1263 );
buf ( n1265 , n1264 );
xor ( n1266 , n1260 , n1265 );
buf ( n1267 , n1266 );
buf ( n1268 , n1267 );
not ( n1269 , n1268 );
buf ( n1270 , n1269 );
buf ( n1271 , n1270 );
and ( n1272 , n1247 , n1271 );
not ( n1273 , n1247 );
buf ( n1274 , n1267 );
and ( n1275 , n1273 , n1274 );
nor ( n1276 , n1272 , n1275 );
buf ( n1277 , n1276 );
xnor ( n1278 , n1232 , n1277 );
buf ( n1279 , n1278 );
xor ( n1280 , n1211 , n1224 );
xor ( n1281 , n1280 , n1279 );
buf ( n1282 , n1281 );
xor ( n1283 , n1211 , n1224 );
and ( n1284 , n1283 , n1279 );
and ( n1285 , n1211 , n1224 );
or ( n1286 , n1284 , n1285 );
buf ( n1287 , n1286 );
not ( n1288 , n1070 );
and ( n1289 , n995 , n1001 );
not ( n1290 , n995 );
and ( n1291 , n1290 , n1000 );
nor ( n1292 , n1289 , n1291 );
xor ( n1293 , n1288 , n1292 );
not ( n1294 , n1293 );
xor ( n1295 , n1150 , n1156 );
xor ( n1296 , n1295 , n1181 );
buf ( n1297 , n1296 );
buf ( n1298 , n1297 );
not ( n1299 , n1298 );
buf ( n1300 , n1299 );
not ( n1301 , n1300 );
and ( n1302 , n1294 , n1301 );
buf ( n1303 , n1293 );
buf ( n1304 , n1300 );
nand ( n1305 , n1303 , n1304 );
buf ( n1306 , n1305 );
buf ( n1307 , n1143 );
buf ( n1308 , n1127 );
xor ( n1309 , n1307 , n1308 );
buf ( n1310 , n1134 );
xor ( n1311 , n1309 , n1310 );
buf ( n1312 , n1311 );
buf ( n1313 , n1312 );
not ( n1314 , n1313 );
buf ( n1315 , n1170 );
buf ( n1316 , n1164 );
and ( n1317 , n1315 , n1316 );
not ( n1318 , n1315 );
buf ( n1319 , n1161 );
and ( n1320 , n1318 , n1319 );
nor ( n1321 , n1317 , n1320 );
buf ( n1322 , n1321 );
buf ( n1323 , n849 );
buf ( n1324 , n798 );
and ( n1325 , n1323 , n1324 );
buf ( n1326 , n1325 );
xnor ( n1327 , n1322 , n1326 );
buf ( n1328 , n1327 );
not ( n1329 , n1328 );
buf ( n1330 , n1329 );
buf ( n1331 , n1330 );
nand ( n1332 , n1314 , n1331 );
buf ( n1333 , n1332 );
buf ( n1334 , n1333 );
buf ( n1335 , n1312 );
not ( n1336 , n1335 );
buf ( n1337 , n1327 );
not ( n1338 , n1337 );
or ( n1339 , n1336 , n1338 );
buf ( n1340 , n812 );
buf ( n1341 , n1340 );
buf ( n1342 , n1341 );
buf ( n1343 , n1342 );
buf ( n1344 , n949 );
and ( n1345 , n1343 , n1344 );
buf ( n1346 , n1345 );
buf ( n1347 , n1346 );
buf ( n1348 , n843 );
buf ( n1349 , n1348 );
buf ( n1350 , n1349 );
buf ( n1351 , n1350 );
not ( n1352 , n1351 );
buf ( n1353 , n883 );
buf ( n1354 , n1353 );
buf ( n1355 , n1354 );
buf ( n1356 , n1355 );
buf ( n1357 , n377 );
nand ( n1358 , n1356 , n1357 );
buf ( n1359 , n1358 );
buf ( n1360 , n1359 );
nor ( n1361 , n1352 , n1360 );
buf ( n1362 , n1361 );
buf ( n1363 , n1362 );
xor ( n1364 , n1347 , n1363 );
nand ( n1365 , n377 , n1038 );
xnor ( n1366 , n1365 , n1034 );
buf ( n1367 , n1366 );
and ( n1368 , n1364 , n1367 );
and ( n1369 , n1347 , n1363 );
or ( n1370 , n1368 , n1369 );
buf ( n1371 , n1370 );
buf ( n1372 , n1371 );
nand ( n1373 , n1339 , n1372 );
buf ( n1374 , n1373 );
buf ( n1375 , n1374 );
nand ( n1376 , n1334 , n1375 );
buf ( n1377 , n1376 );
and ( n1378 , n1306 , n1377 );
nor ( n1379 , n1302 , n1378 );
buf ( n1380 , n1379 );
not ( n1381 , n1380 );
buf ( n1382 , n1381 );
xor ( n1383 , n1051 , n1056 );
xor ( n1384 , n1383 , n1061 );
buf ( n1385 , n1384 );
buf ( n1386 , n1385 );
buf ( n1387 , n883 );
buf ( n1388 , n970 );
and ( n1389 , n1387 , n1388 );
buf ( n1390 , n1389 );
buf ( n1391 , n1390 );
buf ( n1392 , n968 );
buf ( n1393 , n853 );
and ( n1394 , n1392 , n1393 );
buf ( n1395 , n1394 );
buf ( n1396 , n1395 );
xor ( n1397 , n1391 , n1396 );
buf ( n1398 , n1103 );
buf ( n1399 , n798 );
and ( n1400 , n1398 , n1399 );
buf ( n1401 , n1400 );
buf ( n1402 , n1401 );
and ( n1403 , n1397 , n1402 );
and ( n1404 , n1391 , n1396 );
or ( n1405 , n1403 , n1404 );
buf ( n1406 , n1405 );
buf ( n1407 , n1406 );
xor ( n1408 , n1386 , n1407 );
buf ( n1409 , n1085 );
buf ( n1410 , n949 );
and ( n1411 , n1409 , n1410 );
buf ( n1412 , n1411 );
buf ( n1413 , n1412 );
buf ( n1414 , n1342 );
not ( n1415 , n1414 );
buf ( n1416 , n1047 );
nor ( n1417 , n1415 , n1416 );
buf ( n1418 , n1417 );
buf ( n1419 , n1418 );
xor ( n1420 , n1413 , n1419 );
buf ( n1421 , n908 );
buf ( n1422 , n1421 );
buf ( n1423 , n377 );
nand ( n1424 , n1422 , n1423 );
buf ( n1425 , n1424 );
buf ( n1426 , n1425 );
buf ( n1427 , n883 );
buf ( n1428 , n949 );
nand ( n1429 , n1427 , n1428 );
buf ( n1430 , n1429 );
buf ( n1431 , n1430 );
nor ( n1432 , n1426 , n1431 );
buf ( n1433 , n1432 );
buf ( n1434 , n1433 );
and ( n1435 , n1420 , n1434 );
and ( n1436 , n1413 , n1419 );
or ( n1437 , n1435 , n1436 );
buf ( n1438 , n1437 );
buf ( n1439 , n1438 );
and ( n1440 , n1408 , n1439 );
and ( n1441 , n1386 , n1407 );
or ( n1442 , n1440 , n1441 );
buf ( n1443 , n1442 );
buf ( n1444 , n1443 );
buf ( n1445 , n1068 );
not ( n1446 , n1445 );
buf ( n1447 , n1033 );
not ( n1448 , n1447 );
or ( n1449 , n1446 , n1448 );
buf ( n1450 , n1068 );
buf ( n1451 , n1033 );
or ( n1452 , n1450 , n1451 );
nand ( n1453 , n1449 , n1452 );
buf ( n1454 , n1453 );
xor ( n1455 , n1064 , n1454 );
buf ( n1456 , n1455 );
buf ( n1457 , n1312 );
buf ( n1458 , n1330 );
xor ( n1459 , n1457 , n1458 );
buf ( n1460 , n1371 );
xnor ( n1461 , n1459 , n1460 );
buf ( n1462 , n1461 );
buf ( n1463 , n1462 );
xor ( n1464 , n1444 , n1456 );
xor ( n1465 , n1464 , n1463 );
buf ( n1466 , n1465 );
xor ( n1467 , n1444 , n1456 );
and ( n1468 , n1467 , n1463 );
and ( n1469 , n1444 , n1456 );
or ( n1470 , n1468 , n1469 );
buf ( n1471 , n1470 );
buf ( n1472 , n1293 );
buf ( n1473 , n1293 );
not ( n1474 , n1473 );
buf ( n1475 , n1474 );
buf ( n1476 , n1475 );
buf ( n1477 , n1377 );
buf ( n1478 , n1297 );
and ( n1479 , n1477 , n1478 );
not ( n1480 , n1477 );
buf ( n1481 , n1300 );
and ( n1482 , n1480 , n1481 );
nor ( n1483 , n1479 , n1482 );
buf ( n1484 , n1483 );
buf ( n1485 , n1484 );
and ( n1486 , n1485 , n1476 );
not ( n1487 , n1485 );
and ( n1488 , n1487 , n1472 );
nor ( n1489 , n1486 , n1488 );
buf ( n1490 , n1489 );
buf ( n1491 , n1421 );
buf ( n1492 , n1007 );
buf ( n1493 , n1026 );
nand ( n1494 , n1492 , n1493 );
buf ( n1495 , n1494 );
buf ( n1496 , n1495 );
xor ( n1497 , n1491 , n1496 );
buf ( n1498 , n936 );
buf ( n1499 , n1498 );
buf ( n1500 , n1499 );
buf ( n1501 , n1500 );
buf ( n1502 , n1421 );
and ( n1503 , n1501 , n1502 );
buf ( n1504 , n1503 );
buf ( n1505 , n1504 );
xnor ( n1506 , n1497 , n1505 );
buf ( n1507 , n1506 );
buf ( n1508 , n1507 );
buf ( n1509 , n1039 );
buf ( n1510 , n815 );
and ( n1511 , n1509 , n1510 );
buf ( n1512 , n1511 );
buf ( n1513 , n1512 );
buf ( n1514 , n849 );
buf ( n1515 , n967 );
not ( n1516 , n1515 );
buf ( n1517 , n1516 );
and ( n1518 , n1514 , n1517 );
buf ( n1519 , n1518 );
buf ( n1520 , n1519 );
xor ( n1521 , n1513 , n1520 );
buf ( n1522 , n1007 );
buf ( n1523 , n1355 );
nand ( n1524 , n1522 , n1523 );
buf ( n1525 , n1524 );
buf ( n1526 , n1525 );
not ( n1527 , n1526 );
buf ( n1528 , n908 );
buf ( n1529 , n1516 );
nand ( n1530 , n1528 , n1529 );
buf ( n1531 , n1530 );
buf ( n1532 , n1531 );
not ( n1533 , n1532 );
or ( n1534 , n1527 , n1533 );
buf ( n1535 , n1039 );
not ( n1536 , n1535 );
buf ( n1537 , n1031 );
nor ( n1538 , n1536 , n1537 );
buf ( n1539 , n1538 );
buf ( n1540 , n1539 );
nand ( n1541 , n1534 , n1540 );
buf ( n1542 , n1541 );
buf ( n1543 , n1542 );
or ( n1544 , n1525 , n1531 );
buf ( n1545 , n1544 );
nand ( n1546 , n1543 , n1545 );
buf ( n1547 , n1546 );
buf ( n1548 , n1547 );
xor ( n1549 , n1521 , n1548 );
buf ( n1550 , n1549 );
buf ( n1551 , n1550 );
buf ( n1552 , n849 );
buf ( n1553 , n1026 );
and ( n1554 , n1552 , n1553 );
buf ( n1555 , n1554 );
not ( n1556 , n1555 );
buf ( n1557 , n878 );
buf ( n1558 , n883 );
nand ( n1559 , n1557 , n1558 );
buf ( n1560 , n1559 );
buf ( n1561 , n1560 );
buf ( n1562 , n936 );
buf ( n1563 , n968 );
and ( n1564 , n1562 , n1563 );
buf ( n1565 , n1564 );
buf ( n1566 , n1565 );
not ( n1567 , n1566 );
buf ( n1568 , n1567 );
buf ( n1569 , n1568 );
nand ( n1570 , n1561 , n1569 );
buf ( n1571 , n1570 );
not ( n1572 , n1571 );
or ( n1573 , n1556 , n1572 );
buf ( n1574 , n1039 );
buf ( n1575 , n1355 );
nand ( n1576 , n1574 , n1575 );
buf ( n1577 , n1576 );
not ( n1578 , n1577 );
nand ( n1579 , n1578 , n1565 );
nand ( n1580 , n1573 , n1579 );
not ( n1581 , n1580 );
buf ( n1582 , n849 );
not ( n1583 , n1582 );
buf ( n1584 , n821 );
nor ( n1585 , n1583 , n1584 );
buf ( n1586 , n1585 );
not ( n1587 , n1586 );
or ( n1588 , n1581 , n1587 );
buf ( n1589 , n1586 );
not ( n1590 , n1589 );
buf ( n1591 , n1590 );
not ( n1592 , n1591 );
buf ( n1593 , n1580 );
not ( n1594 , n1593 );
buf ( n1595 , n1594 );
not ( n1596 , n1595 );
or ( n1597 , n1592 , n1596 );
buf ( n1598 , n1500 );
not ( n1599 , n1598 );
buf ( n1600 , n812 );
not ( n1601 , n1600 );
buf ( n1602 , n1601 );
buf ( n1603 , n1602 );
not ( n1604 , n1603 );
buf ( n1605 , n908 );
nand ( n1606 , n1604 , n1605 );
buf ( n1607 , n1606 );
buf ( n1608 , n1607 );
not ( n1609 , n1608 );
buf ( n1610 , n1609 );
buf ( n1611 , n1610 );
not ( n1612 , n1611 );
or ( n1613 , n1599 , n1612 );
buf ( n1614 , n1607 );
not ( n1615 , n1614 );
buf ( n1616 , n936 );
not ( n1617 , n1616 );
buf ( n1618 , n1617 );
buf ( n1619 , n1618 );
not ( n1620 , n1619 );
or ( n1621 , n1615 , n1620 );
buf ( n1622 , n796 );
buf ( n1623 , n973 );
and ( n1624 , n1622 , n1623 );
buf ( n1625 , n1624 );
buf ( n1626 , n1625 );
nand ( n1627 , n1621 , n1626 );
buf ( n1628 , n1627 );
buf ( n1629 , n1628 );
nand ( n1630 , n1613 , n1629 );
buf ( n1631 , n1630 );
nand ( n1632 , n1597 , n1631 );
nand ( n1633 , n1588 , n1632 );
buf ( n1634 , n1633 );
xor ( n1635 , n1508 , n1551 );
xor ( n1636 , n1635 , n1634 );
buf ( n1637 , n1636 );
xor ( n1638 , n1508 , n1551 );
and ( n1639 , n1638 , n1634 );
and ( n1640 , n1508 , n1551 );
or ( n1641 , n1639 , n1640 );
buf ( n1642 , n1641 );
xor ( n1643 , n1413 , n1419 );
xor ( n1644 , n1643 , n1434 );
buf ( n1645 , n1644 );
buf ( n1646 , n1645 );
buf ( n1647 , n970 );
buf ( n1648 , n949 );
and ( n1649 , n1647 , n1648 );
buf ( n1650 , n1649 );
buf ( n1651 , n1650 );
buf ( n1652 , n1023 );
not ( n1653 , n1652 );
buf ( n1654 , n853 );
not ( n1655 , n1654 );
buf ( n1656 , n1655 );
buf ( n1657 , n1656 );
nor ( n1658 , n1653 , n1657 );
buf ( n1659 , n1658 );
buf ( n1660 , n1659 );
xor ( n1661 , n1651 , n1660 );
buf ( n1662 , n1342 );
not ( n1663 , n1662 );
buf ( n1664 , n1176 );
nor ( n1665 , n1663 , n1664 );
buf ( n1666 , n1665 );
buf ( n1667 , n1666 );
and ( n1668 , n1661 , n1667 );
and ( n1669 , n1651 , n1660 );
or ( n1670 , n1668 , n1669 );
buf ( n1671 , n1670 );
buf ( n1672 , n1671 );
xor ( n1673 , n1430 , n1425 );
buf ( n1674 , n1673 );
xor ( n1675 , n1672 , n1674 );
buf ( n1676 , n973 );
buf ( n1677 , n377 );
not ( n1678 , n1677 );
buf ( n1679 , n1618 );
nor ( n1680 , n1678 , n1679 );
buf ( n1681 , n1680 );
buf ( n1682 , n1681 );
and ( n1683 , n1676 , n1682 );
buf ( n1684 , n1683 );
buf ( n1685 , n1684 );
and ( n1686 , n1675 , n1685 );
and ( n1687 , n1672 , n1674 );
or ( n1688 , n1686 , n1687 );
buf ( n1689 , n1688 );
buf ( n1690 , n1689 );
buf ( n1691 , n1023 );
buf ( n1692 , n918 );
nand ( n1693 , n1691 , n1692 );
buf ( n1694 , n1693 );
buf ( n1695 , n1694 );
not ( n1696 , n1695 );
buf ( n1697 , n968 );
buf ( n1698 , n798 );
nand ( n1699 , n1697 , n1698 );
buf ( n1700 , n1699 );
buf ( n1701 , n1700 );
not ( n1702 , n1701 );
or ( n1703 , n1696 , n1702 );
buf ( n1704 , n1342 );
buf ( n1705 , n853 );
and ( n1706 , n1704 , n1705 );
buf ( n1707 , n1706 );
buf ( n1708 , n1707 );
nand ( n1709 , n1703 , n1708 );
buf ( n1710 , n1709 );
buf ( n1711 , n1710 );
buf ( n1712 , n1694 );
not ( n1713 , n1712 );
buf ( n1714 , n1713 );
buf ( n1715 , C1 );
buf ( n1716 , n1715 );
nand ( n1717 , n1711 , n1716 );
buf ( n1718 , n1717 );
buf ( n1719 , n1718 );
xor ( n1720 , n1391 , n1396 );
xor ( n1721 , n1720 , n1402 );
buf ( n1722 , n1721 );
buf ( n1723 , n1722 );
xor ( n1724 , n1719 , n1723 );
buf ( n1725 , n1350 );
buf ( n1726 , n377 );
nand ( n1727 , n1725 , n1726 );
buf ( n1728 , n1727 );
xnor ( n1729 , n1355 , n1728 );
buf ( n1730 , n1729 );
xor ( n1731 , n1724 , n1730 );
buf ( n1732 , n1731 );
buf ( n1733 , n1732 );
xor ( n1734 , n1646 , n1690 );
xor ( n1735 , n1734 , n1733 );
buf ( n1736 , n1735 );
xor ( n1737 , n1646 , n1690 );
and ( n1738 , n1737 , n1733 );
and ( n1739 , n1646 , n1690 );
or ( n1740 , n1738 , n1739 );
buf ( n1741 , n1740 );
xnor ( n1742 , n1707 , n1714 );
buf ( n1743 , n1742 );
buf ( n1744 , n1700 );
and ( n1745 , n1743 , n1744 );
nor ( n1746 , n1745 , C0 );
buf ( n1747 , n1746 );
buf ( n1748 , n1747 );
buf ( n1749 , n1355 );
buf ( n1750 , n918 );
and ( n1751 , n1749 , n1750 );
buf ( n1752 , n1751 );
buf ( n1753 , n1752 );
nand ( n1754 , n1516 , n377 );
buf ( n1755 , n1754 );
buf ( n1756 , n973 );
buf ( n1757 , n918 );
nand ( n1758 , n1756 , n1757 );
buf ( n1759 , n1758 );
buf ( n1760 , n1759 );
nor ( n1761 , n1755 , n1760 );
buf ( n1762 , n1761 );
buf ( n1763 , n1762 );
xor ( n1764 , n1753 , n1763 );
xor ( n1765 , n1676 , n1682 );
buf ( n1766 , n1765 );
buf ( n1767 , n1766 );
and ( n1768 , n1764 , n1767 );
and ( n1769 , n1753 , n1763 );
or ( n1770 , n1768 , n1769 );
buf ( n1771 , n1770 );
buf ( n1772 , n1771 );
xor ( n1773 , n1672 , n1674 );
xor ( n1774 , n1773 , n1685 );
buf ( n1775 , n1774 );
buf ( n1776 , n1775 );
xor ( n1777 , n1748 , n1772 );
xor ( n1778 , n1777 , n1776 );
buf ( n1779 , n1778 );
xor ( n1780 , n1748 , n1772 );
and ( n1781 , n1780 , n1776 );
and ( n1782 , n1748 , n1772 );
or ( n1783 , n1781 , n1782 );
buf ( n1784 , n1783 );
xor ( n1785 , n1386 , n1407 );
xor ( n1786 , n1785 , n1439 );
buf ( n1787 , n1786 );
buf ( n1788 , n1516 );
buf ( n1789 , n815 );
and ( n1790 , n1788 , n1789 );
buf ( n1791 , n1790 );
buf ( n1792 , n1791 );
xor ( n1793 , n1236 , n1240 );
and ( n1794 , n1793 , n1245 );
and ( n1795 , n1236 , n1240 );
or ( n1796 , n1794 , n1795 );
buf ( n1797 , n1796 );
xor ( n1798 , n1252 , n1259 );
and ( n1799 , n1798 , n1265 );
and ( n1800 , n1252 , n1259 );
or ( n1801 , n1799 , n1800 );
buf ( n1802 , n1801 );
buf ( n1803 , n1802 );
xor ( n1804 , n1792 , n1797 );
xor ( n1805 , n1804 , n1803 );
buf ( n1806 , n1805 );
xor ( n1807 , n1792 , n1797 );
and ( n1808 , n1807 , n1803 );
and ( n1809 , n1792 , n1797 );
or ( n1810 , n1808 , n1809 );
buf ( n1811 , n1810 );
xor ( n1812 , n1651 , n1660 );
xor ( n1813 , n1812 , n1667 );
buf ( n1814 , n1813 );
buf ( n1815 , n1814 );
buf ( n1816 , n1355 );
buf ( n1817 , n853 );
and ( n1818 , n1816 , n1817 );
buf ( n1819 , n1818 );
buf ( n1820 , n1819 );
buf ( n1821 , n1026 );
buf ( n1822 , n798 );
and ( n1823 , n1821 , n1822 );
buf ( n1824 , n1823 );
buf ( n1825 , n1824 );
xor ( n1826 , n1820 , n1825 );
buf ( n1827 , n815 );
buf ( n1828 , n377 );
nand ( n1829 , n1827 , n1828 );
buf ( n1830 , n1829 );
buf ( n1831 , n1830 );
buf ( n1832 , n949 );
not ( n1833 , n1832 );
buf ( n1834 , n1833 );
buf ( n1835 , n1834 );
nor ( n1836 , n1831 , n1835 );
buf ( n1837 , n1836 );
buf ( n1838 , n1837 );
and ( n1839 , n1826 , n1838 );
or ( n1840 , n1839 , C0 );
buf ( n1841 , n1840 );
buf ( n1842 , n1841 );
xor ( n1843 , n1753 , n1763 );
xor ( n1844 , n1843 , n1767 );
buf ( n1845 , n1844 );
buf ( n1846 , n1845 );
xor ( n1847 , n1815 , n1842 );
xor ( n1848 , n1847 , n1846 );
buf ( n1849 , n1848 );
xor ( n1850 , n1815 , n1842 );
and ( n1851 , n1850 , n1846 );
and ( n1852 , n1815 , n1842 );
or ( n1853 , n1851 , n1852 );
buf ( n1854 , n1853 );
buf ( n1855 , n849 );
not ( n1856 , n1855 );
buf ( n1857 , n1856 );
buf ( n1858 , n1857 );
not ( n1859 , n1421 );
buf ( n1860 , n1859 );
nor ( n1861 , n1858 , n1860 );
buf ( n1862 , n1861 );
buf ( n1863 , n1862 );
buf ( n1864 , n1007 );
buf ( n1865 , n815 );
and ( n1866 , n1864 , n1865 );
buf ( n1867 , n1866 );
buf ( n1868 , n1867 );
buf ( n1869 , n849 );
not ( n1870 , n1869 );
buf ( n1871 , n1618 );
nor ( n1872 , n1870 , n1871 );
buf ( n1873 , n1872 );
buf ( n1874 , n1873 );
xor ( n1875 , n1868 , n1874 );
buf ( n1876 , n1039 );
buf ( n1877 , n1516 );
and ( n1878 , n1876 , n1877 );
buf ( n1879 , n1878 );
buf ( n1880 , n1879 );
and ( n1881 , n1875 , n1880 );
and ( n1882 , n1868 , n1874 );
or ( n1883 , n1881 , n1882 );
buf ( n1884 , n1883 );
buf ( n1885 , n1884 );
buf ( n1886 , n1007 );
buf ( n1887 , n1516 );
and ( n1888 , n1886 , n1887 );
buf ( n1889 , n1888 );
buf ( n1890 , n1889 );
buf ( n1891 , n1857 );
not ( n1892 , n1891 );
buf ( n1893 , n1892 );
buf ( n1894 , n1893 );
xor ( n1895 , n1890 , n1894 );
buf ( n1896 , n1039 );
buf ( n1897 , n1500 );
and ( n1898 , n1896 , n1897 );
buf ( n1899 , n1898 );
buf ( n1900 , n1899 );
xor ( n1901 , n1895 , n1900 );
buf ( n1902 , n1901 );
buf ( n1903 , n1902 );
xor ( n1904 , n1863 , n1885 );
xor ( n1905 , n1904 , n1903 );
buf ( n1906 , n1905 );
xor ( n1907 , n1863 , n1885 );
and ( n1908 , n1907 , n1903 );
and ( n1909 , n1863 , n1885 );
or ( n1910 , n1908 , n1909 );
buf ( n1911 , n1910 );
buf ( n1912 , n1421 );
not ( n1913 , n1912 );
buf ( n1914 , n1495 );
not ( n1915 , n1914 );
buf ( n1916 , n1915 );
buf ( n1917 , n1916 );
not ( n1918 , n1917 );
or ( n1919 , n1913 , n1918 );
buf ( n1920 , n1504 );
not ( n1921 , n1920 );
buf ( n1922 , n1921 );
buf ( n1923 , n1922 );
nand ( n1924 , n1919 , n1923 );
buf ( n1925 , n1924 );
buf ( n1926 , n1925 );
xor ( n1927 , n1868 , n1874 );
xor ( n1928 , n1927 , n1880 );
buf ( n1929 , n1928 );
buf ( n1930 , n1929 );
xor ( n1931 , n1513 , n1520 );
and ( n1932 , n1931 , n1548 );
and ( n1933 , n1513 , n1520 );
or ( n1934 , n1932 , n1933 );
buf ( n1935 , n1934 );
buf ( n1936 , n1935 );
xor ( n1937 , n1926 , n1930 );
xor ( n1938 , n1937 , n1936 );
buf ( n1939 , n1938 );
xor ( n1940 , n1926 , n1930 );
and ( n1941 , n1940 , n1936 );
and ( n1942 , n1926 , n1930 );
or ( n1943 , n1941 , n1942 );
buf ( n1944 , n1943 );
buf ( n1945 , n1246 );
not ( n1946 , n1945 );
buf ( n1947 , n1270 );
nand ( n1948 , n1946 , n1947 );
buf ( n1949 , n1948 );
buf ( n1950 , n1949 );
buf ( n1951 , n1232 );
nand ( n1952 , n1267 , n1246 );
buf ( n1953 , n1952 );
not ( n1954 , n1950 );
not ( n1955 , n1951 );
or ( n1956 , n1954 , n1955 );
nand ( n1957 , n1956 , n1953 );
buf ( n1958 , n1957 );
xor ( n1959 , n1719 , n1723 );
and ( n1960 , n1959 , n1730 );
and ( n1961 , n1719 , n1723 );
or ( n1962 , n1960 , n1961 );
buf ( n1963 , n1962 );
buf ( n1964 , n1355 );
buf ( n1965 , n798 );
nand ( n1966 , n1964 , n1965 );
buf ( n1967 , n1966 );
buf ( n1968 , n1967 );
buf ( n1969 , n973 );
buf ( n1970 , n853 );
nand ( n1971 , n1969 , n1970 );
buf ( n1972 , n1971 );
buf ( n1973 , n1972 );
nand ( n1974 , n1968 , n1973 );
buf ( n1975 , n1974 );
not ( n1976 , n1975 );
buf ( n1977 , n949 );
buf ( n1978 , n918 );
and ( n1979 , n1977 , n1978 );
buf ( n1980 , n1979 );
not ( n1981 , n1980 );
or ( n1982 , n1976 , n1981 );
nand ( n1983 , n1982 , C1 );
buf ( n1984 , n1983 );
xor ( n1985 , n1759 , n1754 );
buf ( n1986 , n1985 );
xor ( n1987 , n1820 , n1825 );
xor ( n1988 , n1987 , n1838 );
buf ( n1989 , n1988 );
buf ( n1990 , n1989 );
xor ( n1991 , n1984 , n1986 );
xor ( n1992 , n1991 , n1990 );
buf ( n1993 , n1992 );
xor ( n1994 , n1984 , n1986 );
and ( n1995 , n1994 , n1990 );
and ( n1996 , n1984 , n1986 );
or ( n1997 , n1995 , n1996 );
buf ( n1998 , n1997 );
xor ( n1999 , n1531 , n1525 );
xor ( n2000 , n1999 , n1539 );
buf ( n2001 , n2000 );
and ( n2002 , n1631 , n1586 );
not ( n2003 , n1631 );
or ( n2004 , n1857 , n821 );
and ( n2005 , n2003 , n2004 );
nor ( n2006 , n2002 , n2005 );
buf ( n2007 , n2006 );
not ( n2008 , n2007 );
buf ( n2009 , n1595 );
not ( n2010 , n2009 );
and ( n2011 , n2008 , n2010 );
buf ( n2012 , n1595 );
buf ( n2013 , n2006 );
and ( n2014 , n2012 , n2013 );
nor ( n2015 , n2011 , n2014 );
buf ( n2016 , n2015 );
buf ( n2017 , n2016 );
nand ( n2018 , n2001 , n2017 );
buf ( n2019 , n2018 );
buf ( n2020 , n1967 );
not ( n2021 , n2020 );
buf ( n2022 , n1980 );
not ( n2023 , n2022 );
buf ( n2024 , n1972 );
not ( n2025 , n2024 );
or ( n2026 , n2023 , n2025 );
buf ( n2027 , n1972 );
buf ( n2028 , n1980 );
or ( n2029 , n2027 , n2028 );
nand ( n2030 , n2026 , n2029 );
buf ( n2031 , n2030 );
buf ( n2032 , n2031 );
not ( n2033 , n2032 );
or ( n2034 , n2021 , n2033 );
buf ( n2035 , n2031 );
buf ( n2036 , n1967 );
or ( n2037 , n2035 , n2036 );
nand ( n2038 , n2034 , n2037 );
buf ( n2039 , n2038 );
buf ( n2040 , n2039 );
buf ( n2041 , n949 );
buf ( n2042 , n853 );
and ( n2043 , n2041 , n2042 );
buf ( n2044 , n2043 );
buf ( n2045 , n2044 );
buf ( n2046 , n1026 );
buf ( n2047 , n377 );
and ( n2048 , n2046 , n2047 );
buf ( n2049 , n2048 );
buf ( n2050 , n2049 );
and ( n2051 , n2045 , n2050 );
buf ( n2052 , n2051 );
buf ( n2053 , n2052 );
buf ( n2054 , n1830 );
buf ( n2055 , n1834 );
and ( n2056 , n2054 , n2055 );
not ( n2057 , n2054 );
buf ( n2058 , n949 );
and ( n2059 , n2057 , n2058 );
nor ( n2060 , n2056 , n2059 );
buf ( n2061 , n2060 );
buf ( n2062 , n2061 );
xor ( n2063 , n2040 , n2053 );
xor ( n2064 , n2063 , n2062 );
buf ( n2065 , n2064 );
xor ( n2066 , n2040 , n2053 );
and ( n2067 , n2066 , n2062 );
and ( n2068 , n2040 , n2053 );
or ( n2069 , n2067 , n2068 );
buf ( n2070 , n2069 );
buf ( n2071 , n402 );
buf ( n2072 , n970 );
buf ( n2073 , n377 );
and ( n2074 , n2072 , n2073 );
buf ( n2075 , n2074 );
buf ( n2076 , n2075 );
and ( n2077 , n2071 , n2076 );
buf ( n2078 , n2077 );
buf ( n2079 , n2078 );
buf ( n2080 , n949 );
buf ( n2081 , n798 );
and ( n2082 , n2080 , n2081 );
buf ( n2083 , n2082 );
buf ( n2084 , n2083 );
buf ( n2085 , n918 );
buf ( n2086 , n918 );
buf ( n2087 , n853 );
nand ( n2088 , n2086 , n2087 );
buf ( n2089 , n2088 );
buf ( n2090 , n2089 );
xor ( n2091 , n2085 , n2090 );
buf ( n2092 , n1359 );
xor ( n2093 , n2091 , n2092 );
buf ( n2094 , n2093 );
buf ( n2095 , n2094 );
xor ( n2096 , n2079 , n2084 );
xor ( n2097 , n2096 , n2095 );
buf ( n2098 , n2097 );
xor ( n2099 , n2079 , n2084 );
and ( n2100 , n2099 , n2095 );
or ( n2101 , n2100 , C0 );
buf ( n2102 , n2101 );
buf ( n2103 , n973 );
buf ( n2104 , n798 );
and ( n2105 , n2103 , n2104 );
buf ( n2106 , n2105 );
buf ( n2107 , n2106 );
buf ( n2108 , n1359 );
not ( n2109 , n2108 );
buf ( n2110 , n918 );
nand ( n2111 , n2109 , n2110 );
buf ( n2112 , n2111 );
buf ( n2113 , n2112 );
buf ( n2114 , n2089 );
nand ( n2115 , n2113 , n2114 );
buf ( n2116 , n2115 );
buf ( n2117 , n2116 );
xor ( n2118 , n2045 , n2050 );
buf ( n2119 , n2118 );
buf ( n2120 , n2119 );
xor ( n2121 , n2107 , n2117 );
xor ( n2122 , n2121 , n2120 );
buf ( n2123 , n2122 );
xor ( n2124 , n2107 , n2117 );
and ( n2125 , n2124 , n2120 );
or ( n2126 , n2125 , C0 );
buf ( n2127 , n2126 );
buf ( n2128 , n1039 );
buf ( n2129 , n1421 );
and ( n2130 , n2128 , n2129 );
buf ( n2131 , n2130 );
buf ( n2132 , n2131 );
buf ( n2133 , n1500 );
buf ( n2134 , n1007 );
and ( n2135 , n2133 , n2134 );
buf ( n2136 , n2135 );
buf ( n2137 , n2136 );
xor ( n2138 , n1890 , n1894 );
and ( n2139 , n2138 , n1900 );
and ( n2140 , n1890 , n1894 );
or ( n2141 , n2139 , n2140 );
buf ( n2142 , n2141 );
buf ( n2143 , n2142 );
xor ( n2144 , n2132 , n2137 );
xor ( n2145 , n2144 , n2143 );
buf ( n2146 , n2145 );
xor ( n2147 , n2132 , n2137 );
and ( n2148 , n2147 , n2143 );
and ( n2149 , n2132 , n2137 );
or ( n2150 , n2148 , n2149 );
buf ( n2151 , n2150 );
xor ( n2152 , n1347 , n1363 );
xor ( n2153 , n2152 , n1367 );
buf ( n2154 , n2153 );
buf ( n2155 , n796 );
buf ( n2156 , n949 );
and ( n2157 , n2155 , n2156 );
buf ( n2158 , n2157 );
buf ( n2159 , n2158 );
buf ( n2160 , n936 );
buf ( n2161 , n1342 );
and ( n2162 , n2160 , n2161 );
buf ( n2163 , n2162 );
buf ( n2164 , n2163 );
xor ( n2165 , n2159 , n2164 );
buf ( n2166 , n908 );
buf ( n2167 , n1023 );
and ( n2168 , n2166 , n2167 );
buf ( n2169 , n2168 );
buf ( n2170 , n2169 );
xor ( n2171 , n2165 , n2170 );
buf ( n2172 , n2171 );
buf ( n2173 , n2172 );
not ( n2174 , n2173 );
buf ( n2175 , n2174 );
buf ( n2176 , n2175 );
buf ( n2177 , n1516 );
buf ( n2178 , n796 );
buf ( n2179 , n918 );
and ( n2180 , n2178 , n2179 );
buf ( n2181 , n2180 );
buf ( n2182 , n2181 );
xor ( n2183 , n2177 , n2182 );
buf ( n2184 , n908 );
buf ( n2185 , n883 );
and ( n2186 , n2184 , n2185 );
buf ( n2187 , n2186 );
buf ( n2188 , n2187 );
and ( n2189 , n2183 , n2188 );
and ( n2190 , n2177 , n2182 );
or ( n2191 , n2189 , n2190 );
buf ( n2192 , n2191 );
buf ( n2193 , n2192 );
buf ( n2194 , n2175 );
buf ( n2195 , n2192 );
not ( n2196 , n2176 );
not ( n2197 , n2193 );
and ( n2198 , n2196 , n2197 );
and ( n2199 , n2194 , n2195 );
nor ( n2200 , n2198 , n2199 );
buf ( n2201 , n2200 );
buf ( n2202 , n2000 );
not ( n2203 , n2202 );
buf ( n2204 , n2203 );
and ( n2205 , n1103 , n1085 );
buf ( n2206 , n2205 );
buf ( n2207 , n872 );
buf ( n2208 , n949 );
and ( n2209 , n2207 , n2208 );
buf ( n2210 , n2209 );
buf ( n2211 , n2210 );
buf ( n2212 , n849 );
buf ( n2213 , n973 );
and ( n2214 , n2212 , n2213 );
buf ( n2215 , n2214 );
buf ( n2216 , n2215 );
xor ( n2217 , n2206 , n2211 );
xor ( n2218 , n2217 , n2216 );
buf ( n2219 , n2218 );
xor ( n2220 , n2206 , n2211 );
and ( n2221 , n2220 , n2216 );
and ( n2222 , n2206 , n2211 );
or ( n2223 , n2221 , n2222 );
buf ( n2224 , n2223 );
buf ( n2225 , n2175 );
buf ( n2226 , n2192 );
not ( n2227 , n2226 );
buf ( n2228 , n2227 );
buf ( n2229 , n2228 );
nand ( n2230 , n2225 , n2229 );
buf ( n2231 , n2230 );
xor ( n2232 , n2159 , n2164 );
and ( n2233 , n2232 , n2170 );
and ( n2234 , n2159 , n2164 );
or ( n2235 , n2233 , n2234 );
buf ( n2236 , n2235 );
buf ( n2237 , n1039 );
buf ( n2238 , n1859 );
not ( n2239 , n2238 );
buf ( n2240 , n1007 );
nand ( n2241 , n2239 , n2240 );
buf ( n2242 , n2241 );
buf ( n2243 , n2242 );
not ( n2244 , n2243 );
buf ( n2245 , n2244 );
buf ( n2246 , n2245 );
buf ( n2247 , n1893 );
buf ( n2248 , n1039 );
nand ( n2249 , n2247 , n2248 );
buf ( n2250 , n2249 );
buf ( n2251 , n2250 );
not ( n2252 , n2237 );
not ( n2253 , n2246 );
or ( n2254 , n2252 , n2253 );
nand ( n2255 , n2254 , n2251 );
buf ( n2256 , n2255 );
xor ( n2257 , n2071 , n2076 );
buf ( n2258 , n2257 );
buf ( n2259 , n404 );
buf ( n2260 , n918 );
buf ( n2261 , n377 );
and ( n2262 , n2260 , n2261 );
buf ( n2263 , n2262 );
buf ( n2264 , n2263 );
xor ( n2265 , n2259 , n2264 );
buf ( n2266 , n2265 );
and ( n2267 , n2259 , n2264 );
buf ( n2268 , n2267 );
buf ( n2269 , n405 );
buf ( n2270 , n798 );
xor ( n2271 , n2269 , n2270 );
buf ( n2272 , n2271 );
and ( n2273 , n2269 , n2270 );
buf ( n2274 , n2273 );
buf ( n2275 , n403 );
buf ( n2276 , n853 );
xor ( n2277 , n2275 , n2276 );
buf ( n2278 , n2277 );
and ( n2279 , n2275 , n2276 );
buf ( n2280 , n2279 );
buf ( n2281 , n1565 );
buf ( n2282 , n1560 );
buf ( n2283 , n1577 );
buf ( n2284 , n1565 );
not ( n2285 , n2281 );
not ( n2286 , n2282 );
or ( n2287 , n2285 , n2286 );
or ( n2288 , n2283 , n2284 );
nand ( n2289 , n2287 , n2288 );
buf ( n2290 , n2289 );
buf ( n2291 , n1893 );
buf ( n2292 , n1007 );
and ( n2293 , n2291 , n2292 );
buf ( n2294 , n2293 );
buf ( n2295 , n949 );
buf ( n2296 , n377 );
and ( n2297 , n2295 , n2296 );
buf ( n2298 , n2297 );
buf ( n2299 , n1039 );
buf ( n2300 , n973 );
and ( n2301 , n2299 , n2300 );
buf ( n2302 , n2301 );
buf ( n2303 , n1893 );
buf ( n2304 , n1355 );
and ( n2305 , n2303 , n2304 );
buf ( n2306 , n2305 );
buf ( n2307 , n2175 );
buf ( n2308 , n2228 );
or ( n2309 , n2307 , n2308 );
buf ( n2310 , n2309 );
buf ( n2311 , n1500 );
buf ( n2312 , n1625 );
buf ( n2313 , n1610 );
xor ( n2314 , n2311 , n2312 );
xor ( n2315 , n2314 , n2313 );
buf ( n2316 , n2315 );
buf ( n2317 , n377 );
buf ( n2318 , n1656 );
not ( n2319 , n2317 );
nor ( n2320 , n2319 , n2318 );
buf ( n2321 , n2320 );
not ( n2322 , n2302 );
xor ( n2323 , n2322 , n2306 );
xnor ( n2324 , n2323 , n2224 );
not ( n2325 , n1196 );
nand ( n2326 , n2325 , n1204 );
not ( n2327 , n2326 );
not ( n2328 , n1209 );
or ( n2329 , n2327 , n2328 );
not ( n2330 , n1204 );
nand ( n2331 , n2330 , n1196 );
nand ( n2332 , n2329 , n2331 );
not ( n2333 , n2332 );
xor ( n2334 , n2177 , n2182 );
xor ( n2335 , n2334 , n2188 );
buf ( n2336 , n2335 );
not ( n2337 , n2336 );
not ( n2338 , n2219 );
nand ( n2339 , n2337 , n2338 );
not ( n2340 , n2339 );
or ( n2341 , n2333 , n2340 );
not ( n2342 , n2338 );
nand ( n2343 , n2342 , n2336 );
nand ( n2344 , n2341 , n2343 );
xor ( n2345 , n2324 , n2344 );
not ( n2346 , n2201 );
not ( n2347 , n2346 );
not ( n2348 , n1811 );
not ( n2349 , n2348 );
or ( n2350 , n2347 , n2349 );
nand ( n2351 , n1811 , n2201 );
nand ( n2352 , n2350 , n2351 );
xor ( n2353 , n2345 , n2352 );
buf ( n2354 , n2353 );
not ( n2355 , n1958 );
not ( n2356 , n1806 );
nand ( n2357 , n2355 , n2356 );
not ( n2358 , n2357 );
xor ( n2359 , n2337 , n2342 );
xnor ( n2360 , n2359 , n2332 );
not ( n2361 , n2360 );
or ( n2362 , n2358 , n2361 );
nand ( n2363 , n1958 , n1806 );
nand ( n2364 , n2362 , n2363 );
buf ( n2365 , n2364 );
nor ( n2366 , n2354 , n2365 );
buf ( n2367 , n2366 );
buf ( n2368 , n2367 );
not ( n2369 , n2368 );
not ( n2370 , n2204 );
not ( n2371 , n2016 );
not ( n2372 , n2371 );
or ( n2373 , n2370 , n2372 );
nand ( n2374 , n2373 , n2019 );
xor ( n2375 , n2236 , n2316 );
xor ( n2376 , n2290 , n1555 );
and ( n2377 , n2375 , n2376 );
and ( n2378 , n2236 , n2316 );
or ( n2379 , n2377 , n2378 );
xor ( n2380 , n2374 , n2379 );
not ( n2381 , n2302 );
not ( n2382 , n2306 );
or ( n2383 , n2381 , n2382 );
not ( n2384 , n2322 );
not ( n2385 , n2306 );
not ( n2386 , n2385 );
or ( n2387 , n2384 , n2386 );
nand ( n2388 , n2387 , n2224 );
nand ( n2389 , n2383 , n2388 );
xor ( n2390 , n2236 , n2316 );
xor ( n2391 , n2390 , n2376 );
xor ( n2392 , n2389 , n2391 );
not ( n2393 , n2231 );
not ( n2394 , n1811 );
or ( n2395 , n2393 , n2394 );
nand ( n2396 , n2395 , n2310 );
and ( n2397 , n2392 , n2396 );
and ( n2398 , n2389 , n2391 );
or ( n2399 , n2397 , n2398 );
nor ( n2400 , n2380 , n2399 );
buf ( n2401 , n2400 );
not ( n2402 , n2401 );
not ( n2403 , n1287 );
not ( n2404 , n1806 );
not ( n2405 , n2355 );
or ( n2406 , n2404 , n2405 );
nand ( n2407 , n1958 , n2356 );
nand ( n2408 , n2406 , n2407 );
and ( n2409 , n2408 , n2360 );
not ( n2410 , n2408 );
not ( n2411 , n2360 );
and ( n2412 , n2410 , n2411 );
nor ( n2413 , n2409 , n2412 );
not ( n2414 , n2413 );
nand ( n2415 , n2403 , n2414 );
buf ( n2416 , n2415 );
xor ( n2417 , n2389 , n2391 );
xor ( n2418 , n2417 , n2396 );
buf ( n2419 , n2418 );
not ( n2420 , n2419 );
buf ( n2421 , n2324 );
or ( n2422 , n2352 , n2421 );
buf ( n2423 , n2344 );
and ( n2424 , n2422 , n2423 );
and ( n2425 , n2352 , n2421 );
nor ( n2426 , n2424 , n2425 );
buf ( n2427 , n2426 );
nand ( n2428 , n2420 , n2427 );
buf ( n2429 , n2428 );
buf ( n2430 , n2429 );
nand ( n2431 , n2369 , n2402 , n2416 , n2430 );
buf ( n2432 , n2431 );
buf ( n2433 , n2432 );
buf ( n2434 , n1642 );
not ( n2435 , n2434 );
buf ( n2436 , n2435 );
buf ( n2437 , n2436 );
buf ( n2438 , n1939 );
not ( n2439 , n2438 );
buf ( n2440 , n2439 );
buf ( n2441 , n2440 );
or ( n2442 , n2437 , n2441 );
buf ( n2443 , n2442 );
not ( n2444 , n2443 );
not ( n2445 , n2371 );
not ( n2446 , n2000 );
or ( n2447 , n2445 , n2446 );
not ( n2448 , n2204 );
not ( n2449 , n2016 );
or ( n2450 , n2448 , n2449 );
nand ( n2451 , n2450 , n2379 );
nand ( n2452 , n2447 , n2451 );
buf ( n2453 , n2452 );
buf ( n2454 , n1637 );
nand ( n2455 , n2453 , n2454 );
buf ( n2456 , n2455 );
buf ( n2457 , n2456 );
not ( n2458 , n2457 );
buf ( n2459 , n2436 );
buf ( n2460 , n2440 );
nand ( n2461 , n2459 , n2460 );
buf ( n2462 , n2461 );
buf ( n2463 , n2462 );
nand ( n2464 , n2458 , n2463 );
buf ( n2465 , n2464 );
not ( n2466 , n2465 );
or ( n2467 , n2444 , n2466 );
or ( n2468 , n2146 , n1911 );
not ( n2469 , n1906 );
not ( n2470 , n1944 );
nand ( n2471 , n2469 , n2470 );
nand ( n2472 , n2468 , n2471 );
not ( n2473 , n2472 );
nand ( n2474 , n2467 , n2473 );
buf ( n2475 , n2474 );
nand ( n2476 , n1944 , n1906 );
not ( n2477 , n2468 );
or ( n2478 , n2476 , n2477 );
nand ( n2479 , n2146 , n1911 );
nand ( n2480 , n2478 , n2479 );
buf ( n2481 , n2480 );
xor ( n2482 , n2250 , n1039 );
xor ( n2483 , n2482 , n2242 );
nand ( n2484 , n2151 , n2483 );
buf ( n2485 , n2484 );
buf ( n2486 , n2256 );
buf ( n2487 , n2294 );
nor ( n2488 , n2486 , n2487 );
buf ( n2489 , n2488 );
buf ( n2490 , n2489 );
or ( n2491 , n2485 , n2490 );
buf ( n2492 , n2256 );
buf ( n2493 , n2294 );
nand ( n2494 , n2492 , n2493 );
buf ( n2495 , n2494 );
buf ( n2496 , n2495 );
nand ( n2497 , n2491 , n2496 );
buf ( n2498 , n2497 );
buf ( n2499 , n2498 );
nor ( n2500 , n2481 , n2499 );
buf ( n2501 , n2500 );
buf ( n2502 , n2501 );
nand ( n2503 , n2433 , n2475 , n2502 );
buf ( n2504 , n2503 );
buf ( n2505 , n2504 );
buf ( n2506 , n1195 );
not ( n2507 , n2506 );
buf ( n2508 , n1282 );
not ( n2509 , n2508 );
and ( n2510 , n2507 , n2509 );
buf ( n2511 , n1190 );
not ( n2512 , n2511 );
buf ( n2513 , n2512 );
buf ( n2514 , n2513 );
buf ( n2515 , n1382 );
not ( n2516 , n2515 );
buf ( n2517 , n2516 );
buf ( n2518 , n2517 );
and ( n2519 , n2514 , n2518 );
nor ( n2520 , n2510 , n2519 );
buf ( n2521 , n2520 );
buf ( n2522 , n1490 );
buf ( n2523 , n1471 );
nor ( n2524 , n2522 , n2523 );
buf ( n2525 , n2524 );
buf ( n2526 , n2525 );
buf ( n2527 , n1466 );
xor ( n2528 , n2154 , n1963 );
and ( n2529 , n2528 , n1787 );
and ( n2530 , n2154 , n1963 );
or ( n2531 , n2529 , n2530 );
buf ( n2532 , n2531 );
nor ( n2533 , n2527 , n2532 );
buf ( n2534 , n2533 );
buf ( n2535 , n2534 );
nor ( n2536 , n2526 , n2535 );
buf ( n2537 , n2536 );
nand ( n2538 , n2521 , n2537 );
nand ( n2539 , n2538 , n2474 , n2501 );
buf ( n2540 , n2539 );
buf ( n2541 , n2498 );
not ( n2542 , n2541 );
buf ( n2543 , n2489 );
not ( n2544 , n2543 );
buf ( n2545 , n2151 );
buf ( n2546 , n2483 );
or ( n2547 , n2545 , n2546 );
buf ( n2548 , n2547 );
buf ( n2549 , n2548 );
nand ( n2550 , n2544 , n2549 );
buf ( n2551 , n2550 );
buf ( n2552 , n2551 );
nand ( n2553 , n2542 , n2552 );
buf ( n2554 , n2553 );
buf ( n2555 , n2554 );
and ( n2556 , n2505 , n2540 , n2555 );
buf ( n2557 , n2556 );
buf ( n2558 , n2557 );
not ( n2559 , n1741 );
xor ( n2560 , n2154 , n1963 );
xor ( n2561 , n2560 , n1787 );
not ( n2562 , n2561 );
and ( n2563 , n2559 , n2562 );
nor ( n2564 , n1736 , n1784 );
nor ( n2565 , n2563 , n2564 );
not ( n2566 , n2565 );
buf ( n2567 , n1779 );
buf ( n2568 , n1854 );
nor ( n2569 , n2567 , n2568 );
buf ( n2570 , n2569 );
buf ( n2571 , n1849 );
buf ( n2572 , n1998 );
nand ( n2573 , n2571 , n2572 );
buf ( n2574 , n2573 );
or ( n2575 , n2570 , n2574 );
buf ( n2576 , n1779 );
buf ( n2577 , n1854 );
nand ( n2578 , n2576 , n2577 );
buf ( n2579 , n2578 );
nand ( n2580 , n2575 , n2579 );
not ( n2581 , n2580 );
or ( n2582 , n2566 , n2581 );
not ( n2583 , n2561 );
not ( n2584 , n1741 );
nand ( n2585 , n2583 , n2584 );
and ( n2586 , n1736 , n1784 );
and ( n2587 , n2585 , n2586 );
buf ( n2588 , n2561 );
buf ( n2589 , n1741 );
and ( n2590 , n2588 , n2589 );
buf ( n2591 , n2590 );
nor ( n2592 , n2587 , n2591 );
nand ( n2593 , n2582 , n2592 );
buf ( n2594 , n2593 );
buf ( n2595 , n2501 );
not ( n2596 , n2595 );
buf ( n2597 , n2596 );
buf ( n2598 , n2597 );
nor ( n2599 , n2594 , n2598 );
buf ( n2600 , n2599 );
buf ( n2601 , n2600 );
not ( n2602 , n2570 );
not ( n2603 , n2602 );
buf ( n2604 , n1849 );
buf ( n2605 , n1998 );
nor ( n2606 , n2604 , n2605 );
buf ( n2607 , n2606 );
buf ( n2608 , n2607 );
nor ( n2609 , n2603 , n2608 );
buf ( n2610 , n2123 );
buf ( n2611 , n2102 );
nor ( n2612 , n2610 , n2611 );
buf ( n2613 , n2612 );
buf ( n2614 , n2613 );
buf ( n2615 , n2098 );
and ( n2616 , n2280 , n2258 );
buf ( n2617 , n2616 );
nand ( n2618 , n2615 , n2617 );
buf ( n2619 , n2618 );
buf ( n2620 , n2619 );
or ( n2621 , n2614 , n2620 );
buf ( n2622 , n2123 );
buf ( n2623 , n2102 );
nand ( n2624 , n2622 , n2623 );
buf ( n2625 , n2624 );
buf ( n2626 , n2625 );
nand ( n2627 , n2621 , n2626 );
buf ( n2628 , n2627 );
not ( n2629 , n2628 );
buf ( n2630 , n1993 );
buf ( n2631 , n2070 );
nor ( n2632 , n2630 , n2631 );
buf ( n2633 , n2632 );
buf ( n2634 , n2633 );
buf ( n2635 , n2065 );
buf ( n2636 , n2127 );
nor ( n2637 , n2635 , n2636 );
buf ( n2638 , n2637 );
buf ( n2639 , n2638 );
nor ( n2640 , n2634 , n2639 );
buf ( n2641 , n2640 );
not ( n2642 , n2641 );
or ( n2643 , n2629 , n2642 );
buf ( n2644 , n2633 );
not ( n2645 , n2644 );
buf ( n2646 , n2645 );
buf ( n2647 , n2646 );
buf ( n2648 , n2127 );
buf ( n2649 , n2065 );
and ( n2650 , n2648 , n2649 );
buf ( n2651 , n2650 );
buf ( n2652 , n2651 );
and ( n2653 , n2647 , n2652 );
buf ( n2654 , n1993 );
buf ( n2655 , n2070 );
and ( n2656 , n2654 , n2655 );
nor ( n2657 , n2653 , n2656 );
buf ( n2658 , n2657 );
nand ( n2659 , n2643 , n2658 );
nand ( n2660 , n2565 , n2609 , n2659 );
buf ( n2661 , n2660 );
buf ( n2662 , n2474 );
nor ( n2663 , n2570 , n2608 );
not ( n2664 , n2638 );
or ( n2665 , n2098 , n2616 );
or ( n2666 , n2123 , n2102 );
xor ( n2667 , n2278 , n2298 );
buf ( n2668 , n2667 );
not ( n2669 , n2668 );
buf ( n2670 , n2268 );
not ( n2671 , n2670 );
and ( n2672 , n2669 , n2671 );
xor ( n2673 , n2280 , n2258 );
buf ( n2674 , n2673 );
and ( n2675 , n2278 , n2298 );
buf ( n2676 , n2675 );
nor ( n2677 , n2674 , n2676 );
buf ( n2678 , n2677 );
buf ( n2679 , n2678 );
nor ( n2680 , n2672 , n2679 );
buf ( n2681 , n2680 );
buf ( n2682 , n2681 );
buf ( n2683 , n2266 );
buf ( n2684 , n2274 );
nor ( n2685 , n2683 , n2684 );
buf ( n2686 , n2685 );
buf ( n2687 , n2686 );
buf ( n2688 , n406 );
not ( n2689 , n2688 );
and ( n2690 , C1 , n2689 );
buf ( n2691 , n407 );
buf ( n2692 , n408 );
buf ( n2693 , n377 );
buf ( n2694 , n409 );
nand ( n2695 , n2691 , n2692 , n2693 , n2694 );
buf ( n2696 , n2695 );
buf ( n2697 , n2696 );
nor ( n2698 , n2690 , n2697 );
buf ( n2699 , n2698 );
buf ( n2700 , n2699 );
nor ( n2701 , C0 , n2700 );
buf ( n2702 , n2701 );
buf ( n2703 , n2702 );
buf ( n2704 , n2321 );
buf ( n2705 , n2272 );
nor ( n2706 , n2704 , n2705 );
buf ( n2707 , n2706 );
buf ( n2708 , n2707 );
nor ( n2709 , n2687 , n2703 , n2708 );
buf ( n2710 , n2709 );
buf ( n2711 , n2710 );
nand ( n2712 , n2682 , n2711 );
buf ( n2713 , n2712 );
buf ( n2714 , n2713 );
buf ( n2715 , n2686 );
not ( n2716 , n2715 );
buf ( n2717 , n2716 );
buf ( n2718 , n2717 );
buf ( n2719 , n2321 );
buf ( n2720 , n2272 );
and ( n2721 , n2718 , n2719 , n2720 );
buf ( n2722 , n2266 );
buf ( n2723 , n2274 );
and ( n2724 , n2722 , n2723 );
nor ( n2725 , n2721 , n2724 );
buf ( n2726 , n2725 );
buf ( n2727 , n2726 );
not ( n2728 , n2727 );
buf ( n2729 , n2681 );
nand ( n2730 , n2728 , n2729 );
buf ( n2731 , n2730 );
buf ( n2732 , n2731 );
buf ( n2733 , n2678 );
not ( n2734 , n2733 );
buf ( n2735 , n2734 );
buf ( n2736 , n2735 );
buf ( n2737 , n2667 );
buf ( n2738 , n2268 );
and ( n2739 , n2736 , n2737 , n2738 );
buf ( n2740 , n2673 );
buf ( n2741 , n2675 );
and ( n2742 , n2740 , n2741 );
nor ( n2743 , n2739 , n2742 );
buf ( n2744 , n2743 );
buf ( n2745 , n2744 );
nand ( n2746 , n2714 , n2732 , n2745 );
buf ( n2747 , n2746 );
nand ( n2748 , n2665 , n2666 , n2747 );
nor ( n2749 , n2748 , n2633 );
nand ( n2750 , n2664 , n2749 );
nor ( n2751 , n2564 , n2750 );
nand ( n2752 , n2663 , n2751 , n2585 );
buf ( n2753 , n2752 );
nand ( n2754 , n2601 , n2661 , n2662 , n2753 );
buf ( n2755 , n2754 );
buf ( n2756 , n2755 );
buf ( n2757 , n2474 );
buf ( n2758 , n2452 );
buf ( n2759 , n1637 );
or ( n2760 , n2758 , n2759 );
buf ( n2761 , n2760 );
buf ( n2762 , n2761 );
buf ( n2763 , n2462 );
nand ( n2764 , n2762 , n2763 );
buf ( n2765 , n2764 );
buf ( n2766 , n2765 );
buf ( n2767 , n2472 );
nor ( n2768 , n2766 , n2767 );
buf ( n2769 , n2768 );
buf ( n2770 , n2769 );
buf ( n2771 , n2597 );
nor ( n2772 , n2770 , n2771 );
buf ( n2773 , n2772 );
buf ( n2774 , n2773 );
nand ( n2775 , n2757 , n2774 );
buf ( n2776 , n2775 );
buf ( n2777 , n2776 );
and ( n2778 , n2756 , n2777 );
buf ( n2779 , n2778 );
buf ( n2780 , n2779 );
nand ( n2781 , n2558 , n2780 );
buf ( n2782 , n2781 );
not ( n2783 , n2593 );
and ( n2784 , n2609 , n2751 , n2585 );
not ( n2785 , n2480 );
nand ( n2786 , n2785 , n2484 );
nor ( n2787 , n2784 , n2786 );
nand ( n2788 , n2474 , n2783 , n2660 , n2787 );
buf ( n2789 , n2788 );
buf ( n2790 , n2465 );
not ( n2791 , n2790 );
buf ( n2792 , n2791 );
buf ( n2793 , n2792 );
not ( n2794 , n2793 );
buf ( n2795 , n2479 );
buf ( n2796 , n2484 );
and ( n2797 , n2795 , n2796 );
buf ( n2798 , n2797 );
buf ( n2799 , n2798 );
buf ( n2800 , n2443 );
buf ( n2801 , n2476 );
nand ( n2802 , n2799 , n2800 , n2801 );
buf ( n2803 , n2802 );
buf ( n2804 , n2803 );
not ( n2805 , n2804 );
and ( n2806 , n2794 , n2805 );
buf ( n2807 , n2472 );
buf ( n2808 , n2798 );
and ( n2809 , n2807 , n2808 );
nor ( n2810 , n2806 , n2809 );
buf ( n2811 , n2810 );
buf ( n2812 , n2811 );
not ( n2813 , n2812 );
buf ( n2814 , n2769 );
not ( n2815 , n2814 );
and ( n2816 , n2813 , n2815 );
buf ( n2817 , n2367 );
not ( n2818 , n2817 );
buf ( n2819 , n2400 );
not ( n2820 , n2819 );
buf ( n2821 , n2415 );
buf ( n2822 , n2429 );
nand ( n2823 , n2818 , n2820 , n2821 , n2822 );
buf ( n2824 , n2823 );
buf ( n2825 , n2824 );
buf ( n2826 , n2811 );
not ( n2827 , n2826 );
buf ( n2828 , n2827 );
buf ( n2829 , n2828 );
and ( n2830 , n2825 , n2829 );
nor ( n2831 , n2816 , n2830 );
buf ( n2832 , n2831 );
buf ( n2833 , n2832 );
and ( n2834 , n2828 , n2538 );
buf ( n2835 , n2548 );
not ( n2836 , n2835 );
buf ( n2837 , n2836 );
nor ( n2838 , n2834 , n2837 );
buf ( n2839 , n2838 );
nand ( n2840 , n2789 , n2833 , n2839 );
buf ( n2841 , n2840 );
buf ( n2842 , n2761 );
buf ( n2843 , n2432 );
not ( n2844 , n2843 );
buf ( n2845 , n2844 );
not ( n2846 , n2845 );
buf ( n2847 , n1490 );
buf ( n2848 , n1471 );
nand ( n2849 , n2847 , n2848 );
buf ( n2850 , n2849 );
nand ( n2851 , n1466 , n2531 );
and ( n2852 , n2850 , n2851 );
nor ( n2853 , n2852 , n2525 );
buf ( n2854 , n2853 );
not ( n2855 , n2854 );
buf ( n2856 , n2521 );
not ( n2857 , n2856 );
or ( n2858 , n2855 , n2857 );
buf ( n2859 , n1195 );
not ( n2860 , n2859 );
buf ( n2861 , n1282 );
not ( n2862 , n2861 );
buf ( n2863 , n2862 );
buf ( n2864 , n2863 );
nand ( n2865 , n2860 , n2864 );
buf ( n2866 , n2865 );
buf ( n2867 , n2866 );
buf ( n2868 , n1190 );
buf ( n2869 , n1382 );
and ( n2870 , n2868 , n2869 );
buf ( n2871 , n2870 );
buf ( n2872 , n2871 );
and ( n2873 , n2867 , n2872 );
buf ( n2874 , n2863 );
not ( n2875 , n2874 );
buf ( n2876 , n2875 );
buf ( n2877 , n2876 );
buf ( n2878 , n1195 );
and ( n2879 , n2877 , n2878 );
nor ( n2880 , n2873 , n2879 );
buf ( n2881 , n2880 );
buf ( n2882 , n2881 );
nand ( n2883 , n2858 , n2882 );
buf ( n2884 , n2883 );
not ( n2885 , n2884 );
or ( n2886 , n2846 , n2885 );
buf ( n2887 , n2400 );
not ( n2888 , n2887 );
buf ( n2889 , n2888 );
nand ( n2890 , n2889 , n2429 );
not ( n2891 , n2890 );
not ( n2892 , n2367 );
buf ( n2893 , n1287 );
not ( n2894 , n2893 );
buf ( n2895 , n2413 );
not ( n2896 , n2895 );
or ( n2897 , n2894 , n2896 );
buf ( n2898 , n2353 );
buf ( n2899 , n2364 );
nand ( n2900 , n2898 , n2899 );
buf ( n2901 , n2900 );
buf ( n2902 , n2901 );
nand ( n2903 , n2897 , n2902 );
buf ( n2904 , n2903 );
nand ( n2905 , n2892 , n2904 );
not ( n2906 , n2905 );
and ( n2907 , n2891 , n2906 );
not ( n2908 , n2400 );
not ( n2909 , n2908 );
and ( n2910 , n2422 , n2423 );
nor ( n2911 , n2910 , n2425 );
not ( n2912 , n2418 );
nor ( n2913 , n2911 , n2912 );
not ( n2914 , n2913 );
or ( n2915 , n2909 , n2914 );
nand ( n2916 , n2380 , n2399 );
nand ( n2917 , n2915 , n2916 );
nor ( n2918 , n2907 , n2917 );
nand ( n2919 , n2886 , n2918 );
buf ( n2920 , n2919 );
nand ( n2921 , n2842 , n2920 );
buf ( n2922 , n2921 );
buf ( n2923 , n2922 );
nand ( n2924 , n2783 , n2752 , n2660 );
buf ( n2925 , n2924 );
buf ( n2926 , n2925 );
buf ( n2927 , n2521 );
not ( n2928 , n2927 );
buf ( n2929 , n2525 );
buf ( n2930 , n2534 );
or ( n2931 , n2929 , n2930 );
buf ( n2932 , n2931 );
buf ( n2933 , n2932 );
nor ( n2934 , n2928 , n2933 );
buf ( n2935 , n2934 );
and ( n2936 , n2845 , n2935 );
buf ( n2937 , n2936 );
buf ( n2938 , n2761 );
nand ( n2939 , n2926 , n2937 , n2938 );
buf ( n2940 , n2939 );
buf ( n2941 , n2940 );
buf ( n2942 , n2456 );
nand ( n2943 , n2923 , n2941 , n2942 );
buf ( n2944 , n2943 );
buf ( n2945 , n2925 );
not ( n2946 , n2415 );
buf ( n2947 , n2367 );
nor ( n2948 , n2946 , n2947 );
not ( n2949 , n2948 );
nor ( n2950 , n2949 , n2538 );
buf ( n2951 , n2950 );
nand ( n2952 , n2945 , n2951 );
buf ( n2953 , n2952 );
buf ( n2954 , C1 );
buf ( n2955 , n2769 );
not ( n2956 , n2955 );
buf ( n2957 , n2956 );
buf ( n2958 , n2957 );
buf ( n2959 , n2551 );
not ( n2960 , n2959 );
buf ( n2961 , n1007 );
nand ( n2962 , n2960 , n2961 );
buf ( n2963 , n2962 );
buf ( n2964 , n2963 );
nor ( n2965 , n2958 , n2964 );
buf ( n2966 , n2965 );
buf ( n2967 , C1 );
buf ( n2968 , n2919 );
not ( n2969 , n2765 );
buf ( n2970 , n2969 );
nand ( n2971 , n2968 , n2970 );
buf ( n2972 , n2971 );
buf ( n2973 , n2919 );
buf ( n2974 , n2769 );
nand ( n2975 , n2973 , n2974 );
buf ( n2976 , n2975 );
not ( n2977 , n2845 );
not ( n2978 , n2884 );
or ( n2979 , n2977 , n2978 );
nand ( n2980 , n2979 , n2918 );
buf ( n2981 , n2980 );
buf ( n2982 , n2966 );
nand ( n2983 , n2981 , n2982 );
buf ( n2984 , n2983 );
buf ( n2985 , n2919 );
not ( n2986 , n2985 );
buf ( n2987 , n2986 );
not ( n2988 , n2947 );
not ( n2989 , n2415 );
not ( n2990 , n2429 );
nor ( n2991 , n2989 , n2990 );
nand ( n2992 , n2988 , n2991 );
not ( n2993 , n2992 );
buf ( n2994 , n2993 );
buf ( n2995 , n2884 );
or ( n2996 , n2990 , n2905 );
not ( n2997 , n2913 );
nand ( n2998 , n2996 , n2997 );
buf ( n2999 , n2998 );
and ( n3000 , n2994 , n2995 );
nor ( n3001 , n3000 , n2999 );
buf ( n3002 , n3001 );
buf ( n3003 , n2480 );
not ( n3004 , n3003 );
buf ( n3005 , n2474 );
nand ( n3006 , n3004 , n3005 );
buf ( n3007 , n3006 );
buf ( n3008 , n3007 );
buf ( n3009 , n2963 );
not ( n3010 , n3009 );
buf ( n3011 , n3010 );
buf ( n3012 , n3011 );
buf ( n3013 , n1007 );
not ( n3014 , n3013 );
buf ( n3015 , n2498 );
not ( n3016 , n3015 );
or ( n3017 , n3014 , n3016 );
nand ( n3018 , n1039 , n1007 );
buf ( n3019 , n3018 );
nand ( n3020 , n3017 , n3019 );
buf ( n3021 , n3020 );
buf ( n3022 , n3021 );
and ( n3023 , n3008 , n3012 );
nor ( n3024 , n3023 , n3022 );
buf ( n3025 , n3024 );
buf ( n3026 , n2957 );
buf ( n3027 , n2551 );
nor ( n3028 , n3026 , n3027 );
buf ( n3029 , n3028 );
buf ( n3030 , n2957 );
buf ( n3031 , n2837 );
nor ( n3032 , n3030 , n3031 );
buf ( n3033 , n3032 );
not ( n3034 , n2990 );
nand ( n3035 , n3034 , n2997 );
buf ( n3036 , n3035 );
not ( n3037 , n3036 );
buf ( n3038 , n3037 );
buf ( n3039 , n2462 );
buf ( n3040 , n2443 );
nand ( n3041 , n3039 , n3040 );
buf ( n3042 , n3041 );
buf ( n3043 , n2944 );
buf ( n3044 , n3042 );
xnor ( n3045 , n3043 , n3044 );
buf ( n3046 , n3045 );
buf ( n3047 , n409 );
buf ( n3048 , n415 );
and ( n3049 , n3047 , n3048 );
buf ( n3050 , n3049 );
buf ( n3051 , n3050 );
buf ( n3052 , n407 );
buf ( n3053 , n417 );
and ( n3054 , n3052 , n3053 );
buf ( n3055 , n3054 );
buf ( n3056 , n3055 );
buf ( n3057 , n408 );
buf ( n3058 , n416 );
and ( n3059 , n3057 , n3058 );
buf ( n3060 , n3059 );
buf ( n3061 , n3060 );
xor ( n3062 , n3051 , n3056 );
xor ( n3063 , n3062 , n3061 );
buf ( n3064 , n3063 );
xor ( n3065 , n3051 , n3056 );
and ( n3066 , n3065 , n3061 );
and ( n3067 , n3051 , n3056 );
or ( n3068 , n3066 , n3067 );
buf ( n3069 , n3068 );
buf ( n3070 , n391 );
buf ( n3071 , n393 );
and ( n3072 , n3070 , n3071 );
buf ( n3073 , n3072 );
buf ( n3074 , n3073 );
buf ( n3075 , n392 );
buf ( n3076 , n393 );
nand ( n3077 , n3075 , n3076 );
buf ( n3078 , n3077 );
buf ( n3079 , n3078 );
buf ( n3080 , n409 );
buf ( n3081 , n416 );
nand ( n3082 , n3080 , n3081 );
buf ( n3083 , n3082 );
buf ( n3084 , n3083 );
nor ( n3085 , n3079 , n3084 );
buf ( n3086 , n3085 );
buf ( n3087 , n3086 );
buf ( n3088 , C0 );
xor ( n3089 , n3074 , n3087 );
xor ( n3090 , n3089 , n3088 );
buf ( n3091 , n3090 );
and ( n3092 , n3074 , n3087 );
or ( n3093 , C0 , n3092 );
buf ( n3094 , n3093 );
buf ( n3095 , n408 );
buf ( n3096 , n415 );
and ( n3097 , n3095 , n3096 );
buf ( n3098 , n3097 );
buf ( n3099 , n3098 );
buf ( n3100 , n407 );
buf ( n3101 , n416 );
and ( n3102 , n3100 , n3101 );
buf ( n3103 , n3102 );
buf ( n3104 , n3103 );
buf ( n3105 , n406 );
buf ( n3106 , n417 );
and ( n3107 , n3105 , n3106 );
buf ( n3108 , n3107 );
buf ( n3109 , n3108 );
xor ( n3110 , n3099 , n3104 );
xor ( n3111 , n3110 , n3109 );
buf ( n3112 , n3111 );
xor ( n3113 , n3099 , n3104 );
and ( n3114 , n3113 , n3109 );
and ( n3115 , n3099 , n3104 );
or ( n3116 , n3114 , n3115 );
buf ( n3117 , n3116 );
not ( n3118 , n392 );
nand ( n3119 , n3118 , n391 , n393 );
not ( n3120 , n391 );
nand ( n3121 , n3120 , n392 , n393 );
nand ( n3122 , n3119 , n3121 );
buf ( n3123 , n3122 );
buf ( n3124 , n409 );
buf ( n3125 , n414 );
nand ( n3126 , n3124 , n3125 );
buf ( n3127 , n3126 );
buf ( n3128 , n390 );
buf ( n3129 , n393 );
nand ( n3130 , n3128 , n3129 );
buf ( n3131 , n3130 );
xor ( n3132 , n3127 , n3131 );
buf ( n3133 , n3132 );
not ( n3134 , n392 );
nor ( n3135 , n3134 , n393 );
buf ( n3136 , n3135 );
xor ( n3137 , n3123 , n3133 );
xor ( n3138 , n3137 , n3136 );
buf ( n3139 , n3138 );
xor ( n3140 , n3123 , n3133 );
and ( n3141 , n3140 , n3136 );
and ( n3142 , n3123 , n3133 );
or ( n3143 , n3141 , n3142 );
buf ( n3144 , n3143 );
buf ( n3145 , n3069 );
buf ( n3146 , n3112 );
buf ( n3147 , n3094 );
xor ( n3148 , n3145 , n3146 );
xor ( n3149 , n3148 , n3147 );
buf ( n3150 , n3149 );
xor ( n3151 , n3145 , n3146 );
and ( n3152 , n3151 , n3147 );
and ( n3153 , n3145 , n3146 );
or ( n3154 , n3152 , n3153 );
buf ( n3155 , n3154 );
buf ( n3156 , n407 );
buf ( n3157 , n415 );
and ( n3158 , n3156 , n3157 );
buf ( n3159 , n3158 );
buf ( n3160 , n3159 );
buf ( n3161 , n409 );
buf ( n3162 , n413 );
and ( n3163 , n3161 , n3162 );
buf ( n3164 , n3163 );
buf ( n3165 , n3164 );
buf ( n3166 , n406 );
buf ( n3167 , n416 );
and ( n3168 , n3166 , n3167 );
buf ( n3169 , n3168 );
buf ( n3170 , n3169 );
xor ( n3171 , n3160 , n3165 );
xor ( n3172 , n3171 , n3170 );
buf ( n3173 , n3172 );
xor ( n3174 , n3160 , n3165 );
and ( n3175 , n3174 , n3170 );
and ( n3176 , n3160 , n3165 );
or ( n3177 , n3175 , n3176 );
buf ( n3178 , n3177 );
buf ( n3179 , n405 );
buf ( n3180 , n417 );
and ( n3181 , n3179 , n3180 );
buf ( n3182 , n3181 );
buf ( n3183 , n3182 );
buf ( n3184 , n408 );
buf ( n3185 , n414 );
and ( n3186 , n3184 , n3185 );
buf ( n3187 , n3186 );
buf ( n3188 , n3187 );
buf ( n3189 , n389 );
buf ( n3190 , n393 );
and ( n3191 , n3189 , n3190 );
buf ( n3192 , n3191 );
buf ( n3193 , n3192 );
xor ( n3194 , n3188 , n3193 );
buf ( n3195 , n3194 );
buf ( n3196 , n3195 );
buf ( n3197 , n3135 );
buf ( n3198 , n391 );
and ( n3199 , n3197 , n3198 );
buf ( n3200 , n3199 );
buf ( n3201 , n3200 );
xor ( n3202 , n3183 , n3196 );
xor ( n3203 , n3202 , n3201 );
buf ( n3204 , n3203 );
xor ( n3205 , n3183 , n3196 );
and ( n3206 , n3205 , n3201 );
and ( n3207 , n3183 , n3196 );
or ( n3208 , n3206 , n3207 );
buf ( n3209 , n3208 );
buf ( n3210 , n3131 );
buf ( n3211 , n3127 );
nor ( n3212 , n3210 , n3211 );
buf ( n3213 , n3212 );
buf ( n3214 , n3213 );
buf ( n3215 , n3122 );
buf ( n3216 , n392 );
and ( n3217 , n3215 , n3216 );
buf ( n3218 , n3217 );
buf ( n3219 , n3218 );
buf ( n3220 , n3117 );
xor ( n3221 , n3214 , n3219 );
xor ( n3222 , n3221 , n3220 );
buf ( n3223 , n3222 );
xor ( n3224 , n3214 , n3219 );
and ( n3225 , n3224 , n3220 );
and ( n3226 , n3214 , n3219 );
or ( n3227 , n3225 , n3226 );
buf ( n3228 , n3227 );
buf ( n3229 , n3173 );
buf ( n3230 , n3144 );
buf ( n3231 , n3204 );
xor ( n3232 , n3229 , n3230 );
xor ( n3233 , n3232 , n3231 );
buf ( n3234 , n3233 );
xor ( n3235 , n3229 , n3230 );
and ( n3236 , n3235 , n3231 );
and ( n3237 , n3229 , n3230 );
or ( n3238 , n3236 , n3237 );
buf ( n3239 , n3238 );
nand ( n3240 , n392 , n391 );
not ( n3241 , n3240 );
nand ( n3242 , n390 , n393 );
and ( n3243 , n3242 , n3120 );
not ( n3244 , n3242 );
and ( n3245 , n3244 , n391 );
or ( n3246 , n3243 , n3245 );
not ( n3247 , n3246 );
or ( n3248 , n3241 , n3247 );
and ( n3249 , n391 , n392 );
nand ( n3250 , n3249 , n3242 );
nand ( n3251 , n3248 , n3250 );
nand ( n3252 , n392 , n393 , n391 );
and ( n3253 , n3251 , n3252 );
not ( n3254 , n3251 );
not ( n3255 , n3252 );
and ( n3256 , n3254 , n3255 );
nor ( n3257 , n3253 , n3256 );
buf ( n3258 , n3257 );
buf ( n3259 , n3258 );
buf ( n3260 , n393 );
and ( n3261 , n3259 , n3260 );
buf ( n3262 , n3261 );
buf ( n3263 , n3262 );
buf ( n3264 , n3223 );
buf ( n3265 , n3155 );
xor ( n3266 , n3263 , n3264 );
xor ( n3267 , n3266 , n3265 );
buf ( n3268 , n3267 );
xor ( n3269 , n3263 , n3264 );
and ( n3270 , n3269 , n3265 );
and ( n3271 , n3263 , n3264 );
or ( n3272 , n3270 , n3271 );
buf ( n3273 , n3272 );
buf ( n3274 , n407 );
buf ( n3275 , n414 );
and ( n3276 , n3274 , n3275 );
buf ( n3277 , n3276 );
buf ( n3278 , n3277 );
buf ( n3279 , n408 );
buf ( n3280 , n413 );
and ( n3281 , n3279 , n3280 );
buf ( n3282 , n3281 );
buf ( n3283 , n3282 );
buf ( n3284 , n409 );
buf ( n3285 , n412 );
and ( n3286 , n3284 , n3285 );
buf ( n3287 , n3286 );
buf ( n3288 , n3287 );
xor ( n3289 , n3278 , n3283 );
xor ( n3290 , n3289 , n3288 );
buf ( n3291 , n3290 );
xor ( n3292 , n3278 , n3283 );
and ( n3293 , n3292 , n3288 );
and ( n3294 , n3278 , n3283 );
or ( n3295 , n3293 , n3294 );
buf ( n3296 , n3295 );
buf ( n3297 , n388 );
buf ( n3298 , n393 );
and ( n3299 , n3297 , n3298 );
buf ( n3300 , n3299 );
buf ( n3301 , n3300 );
buf ( n3302 , n404 );
buf ( n3303 , n417 );
and ( n3304 , n3302 , n3303 );
buf ( n3305 , n3304 );
buf ( n3306 , n3305 );
buf ( n3307 , n3135 );
buf ( n3308 , n390 );
and ( n3309 , n3307 , n3308 );
buf ( n3310 , n3309 );
buf ( n3311 , n3310 );
xor ( n3312 , n3301 , n3306 );
xor ( n3313 , n3312 , n3311 );
buf ( n3314 , n3313 );
xor ( n3315 , n3301 , n3306 );
and ( n3316 , n3315 , n3311 );
and ( n3317 , n3301 , n3306 );
or ( n3318 , n3316 , n3317 );
buf ( n3319 , n3318 );
buf ( n3320 , n405 );
buf ( n3321 , n416 );
and ( n3322 , n3320 , n3321 );
buf ( n3323 , n3322 );
buf ( n3324 , n3323 );
buf ( n3325 , n406 );
buf ( n3326 , n415 );
and ( n3327 , n3325 , n3326 );
buf ( n3328 , n3327 );
buf ( n3329 , n3328 );
xor ( n3330 , n3324 , n3329 );
buf ( n3331 , n3330 );
buf ( n3332 , n3331 );
buf ( n3333 , n3122 );
buf ( n3334 , n391 );
and ( n3335 , n3333 , n3334 );
buf ( n3336 , n3335 );
buf ( n3337 , n3336 );
and ( n3338 , n3188 , n3193 );
buf ( n3339 , n3338 );
buf ( n3340 , n3339 );
xor ( n3341 , n3332 , n3337 );
xor ( n3342 , n3341 , n3340 );
buf ( n3343 , n3342 );
xor ( n3344 , n3332 , n3337 );
and ( n3345 , n3344 , n3340 );
and ( n3346 , n3332 , n3337 );
or ( n3347 , n3345 , n3346 );
buf ( n3348 , n3347 );
buf ( n3349 , n3178 );
buf ( n3350 , n3291 );
buf ( n3351 , n3314 );
xor ( n3352 , n3349 , n3350 );
xor ( n3353 , n3352 , n3351 );
buf ( n3354 , n3353 );
xor ( n3355 , n3349 , n3350 );
and ( n3356 , n3355 , n3351 );
and ( n3357 , n3349 , n3350 );
or ( n3358 , n3356 , n3357 );
buf ( n3359 , n3358 );
buf ( n3360 , n3209 );
buf ( n3361 , n3228 );
buf ( n3362 , n3343 );
xor ( n3363 , n3360 , n3361 );
xor ( n3364 , n3363 , n3362 );
buf ( n3365 , n3364 );
xor ( n3366 , n3360 , n3361 );
and ( n3367 , n3366 , n3362 );
and ( n3368 , n3360 , n3361 );
or ( n3369 , n3367 , n3368 );
buf ( n3370 , n3369 );
buf ( n3371 , n3258 );
buf ( n3372 , n392 );
and ( n3373 , n3371 , n3372 );
buf ( n3374 , n3373 );
buf ( n3375 , n3374 );
nand ( n3376 , n392 , n390 );
nand ( n3377 , n393 , n389 );
or ( n3378 , n3376 , n3377 );
not ( n3379 , n393 );
not ( n3380 , n389 );
or ( n3381 , n3379 , n3380 );
nand ( n3382 , n392 , n390 );
nand ( n3383 , n3381 , n3382 );
nand ( n3384 , n3378 , n3383 );
buf ( n3385 , n3384 );
nand ( n3386 , n393 , n390 , n391 );
or ( n3387 , n3385 , n3386 );
nand ( n3388 , n3384 , n3386 );
buf ( n3389 , n3388 );
nand ( n3390 , n3387 , n3389 );
nand ( n3391 , n393 , n392 , n391 );
nand ( n3392 , n3391 , n3250 );
not ( n3393 , n3392 );
and ( n3394 , n3390 , n3393 );
not ( n3395 , n3390 );
and ( n3396 , n3395 , n3392 );
nor ( n3397 , n3394 , n3396 );
buf ( n3398 , n3397 );
buf ( n3399 , n393 );
and ( n3400 , n3398 , n3399 );
buf ( n3401 , n3400 );
buf ( n3402 , n3401 );
buf ( n3403 , n3354 );
xor ( n3404 , n3375 , n3402 );
xor ( n3405 , n3404 , n3403 );
buf ( n3406 , n3405 );
xor ( n3407 , n3375 , n3402 );
and ( n3408 , n3407 , n3403 );
and ( n3409 , n3375 , n3402 );
or ( n3410 , n3408 , n3409 );
buf ( n3411 , n3410 );
buf ( n3412 , n3239 );
buf ( n3413 , n3365 );
buf ( n3414 , n3406 );
xor ( n3415 , n3412 , n3413 );
xor ( n3416 , n3415 , n3414 );
buf ( n3417 , n3416 );
xor ( n3418 , n3412 , n3413 );
and ( n3419 , n3418 , n3414 );
and ( n3420 , n3412 , n3413 );
or ( n3421 , n3419 , n3420 );
buf ( n3422 , n3421 );
buf ( n3423 , n409 );
buf ( n3424 , n411 );
and ( n3425 , n3423 , n3424 );
buf ( n3426 , n3425 );
buf ( n3427 , n3426 );
buf ( n3428 , n387 );
buf ( n3429 , n393 );
and ( n3430 , n3428 , n3429 );
buf ( n3431 , n3430 );
buf ( n3432 , n3431 );
buf ( n3433 , n405 );
buf ( n3434 , n415 );
and ( n3435 , n3433 , n3434 );
buf ( n3436 , n3435 );
buf ( n3437 , n3436 );
xor ( n3438 , n3427 , n3432 );
xor ( n3439 , n3438 , n3437 );
buf ( n3440 , n3439 );
xor ( n3441 , n3427 , n3432 );
and ( n3442 , n3441 , n3437 );
and ( n3443 , n3427 , n3432 );
or ( n3444 , n3442 , n3443 );
buf ( n3445 , n3444 );
buf ( n3446 , n407 );
buf ( n3447 , n413 );
and ( n3448 , n3446 , n3447 );
buf ( n3449 , n3448 );
buf ( n3450 , n3449 );
buf ( n3451 , n408 );
buf ( n3452 , n412 );
and ( n3453 , n3451 , n3452 );
buf ( n3454 , n3453 );
buf ( n3455 , n3454 );
buf ( n3456 , n406 );
buf ( n3457 , n414 );
and ( n3458 , n3456 , n3457 );
buf ( n3459 , n3458 );
buf ( n3460 , n3459 );
xor ( n3461 , n3450 , n3455 );
xor ( n3462 , n3461 , n3460 );
buf ( n3463 , n3462 );
xor ( n3464 , n3450 , n3455 );
and ( n3465 , n3464 , n3460 );
and ( n3466 , n3450 , n3455 );
or ( n3467 , n3465 , n3466 );
buf ( n3468 , n3467 );
buf ( n3469 , n3122 );
buf ( n3470 , n390 );
and ( n3471 , n3469 , n3470 );
buf ( n3472 , n3471 );
buf ( n3473 , n3472 );
buf ( n3474 , n403 );
buf ( n3475 , n417 );
and ( n3476 , n3474 , n3475 );
buf ( n3477 , n3476 );
buf ( n3478 , n3477 );
buf ( n3479 , n404 );
buf ( n3480 , n416 );
and ( n3481 , n3479 , n3480 );
buf ( n3482 , n3481 );
buf ( n3483 , n3482 );
xor ( n3484 , n3478 , n3483 );
buf ( n3485 , n3484 );
buf ( n3486 , n3485 );
buf ( n3487 , n3135 );
buf ( n3488 , n389 );
and ( n3489 , n3487 , n3488 );
buf ( n3490 , n3489 );
buf ( n3491 , n3490 );
xor ( n3492 , n3473 , n3486 );
xor ( n3493 , n3492 , n3491 );
buf ( n3494 , n3493 );
xor ( n3495 , n3473 , n3486 );
and ( n3496 , n3495 , n3491 );
and ( n3497 , n3473 , n3486 );
or ( n3498 , n3496 , n3497 );
buf ( n3499 , n3498 );
and ( n3500 , n3324 , n3329 );
buf ( n3501 , n3500 );
buf ( n3502 , n3501 );
buf ( n3503 , n3296 );
buf ( n3504 , n3440 );
xor ( n3505 , n3502 , n3503 );
xor ( n3506 , n3505 , n3504 );
buf ( n3507 , n3506 );
xor ( n3508 , n3502 , n3503 );
and ( n3509 , n3508 , n3504 );
and ( n3510 , n3502 , n3503 );
or ( n3511 , n3509 , n3510 );
buf ( n3512 , n3511 );
buf ( n3513 , n3463 );
buf ( n3514 , n3319 );
buf ( n3515 , n3348 );
xor ( n3516 , n3513 , n3514 );
xor ( n3517 , n3516 , n3515 );
buf ( n3518 , n3517 );
xor ( n3519 , n3513 , n3514 );
and ( n3520 , n3519 , n3515 );
and ( n3521 , n3513 , n3514 );
or ( n3522 , n3520 , n3521 );
buf ( n3523 , n3522 );
buf ( n3524 , n3257 );
buf ( n3525 , n391 );
and ( n3526 , n3524 , n3525 );
buf ( n3527 , n3526 );
buf ( n3528 , n3527 );
buf ( n3529 , n3494 );
not ( n3530 , n3397 );
buf ( n3531 , n392 );
not ( n3532 , n3531 );
buf ( n3533 , n3532 );
nor ( n3534 , n3530 , n3533 );
buf ( n3535 , n3534 );
xor ( n3536 , n3528 , n3529 );
xor ( n3537 , n3536 , n3535 );
buf ( n3538 , n3537 );
xor ( n3539 , n3528 , n3529 );
and ( n3540 , n3539 , n3535 );
and ( n3541 , n3528 , n3529 );
or ( n3542 , n3540 , n3541 );
buf ( n3543 , n3542 );
buf ( n3544 , n3507 );
nand ( n3545 , n389 , n392 , n390 , n393 );
nand ( n3546 , n388 , n393 );
not ( n3547 , n3546 );
and ( n3548 , n389 , n392 );
xor ( n3549 , n3547 , n3548 );
not ( n3550 , n390 );
nor ( n3551 , n3550 , n391 );
xor ( n3552 , n3549 , n3551 );
xor ( n3553 , n3545 , n3552 );
not ( n3554 , n3250 );
not ( n3555 , n3554 );
not ( n3556 , n3388 );
or ( n3557 , n3555 , n3556 );
not ( n3558 , n3384 );
not ( n3559 , n3386 );
and ( n3560 , n3558 , n3559 );
not ( n3561 , n3391 );
and ( n3562 , n3388 , n3561 );
nor ( n3563 , n3560 , n3562 );
nand ( n3564 , n3557 , n3563 );
xnor ( n3565 , n3553 , n3564 );
buf ( n3566 , n3565 );
buf ( n3567 , n393 );
and ( n3568 , n3566 , n3567 );
buf ( n3569 , n3568 );
buf ( n3570 , n3569 );
buf ( n3571 , n3359 );
xor ( n3572 , n3544 , n3570 );
xor ( n3573 , n3572 , n3571 );
buf ( n3574 , n3573 );
xor ( n3575 , n3544 , n3570 );
and ( n3576 , n3575 , n3571 );
and ( n3577 , n3544 , n3570 );
or ( n3578 , n3576 , n3577 );
buf ( n3579 , n3578 );
buf ( n3580 , n3370 );
buf ( n3581 , n3518 );
buf ( n3582 , n3538 );
xor ( n3583 , n3580 , n3581 );
xor ( n3584 , n3583 , n3582 );
buf ( n3585 , n3584 );
xor ( n3586 , n3580 , n3581 );
and ( n3587 , n3586 , n3582 );
and ( n3588 , n3580 , n3581 );
or ( n3589 , n3587 , n3588 );
buf ( n3590 , n3589 );
buf ( n3591 , n3411 );
buf ( n3592 , n3574 );
buf ( n3593 , n3585 );
xor ( n3594 , n3591 , n3592 );
xor ( n3595 , n3594 , n3593 );
buf ( n3596 , n3595 );
xor ( n3597 , n3591 , n3592 );
and ( n3598 , n3597 , n3593 );
and ( n3599 , n3591 , n3592 );
or ( n3600 , n3598 , n3599 );
buf ( n3601 , n3600 );
buf ( n3602 , n406 );
buf ( n3603 , n413 );
and ( n3604 , n3602 , n3603 );
buf ( n3605 , n3604 );
buf ( n3606 , n3605 );
buf ( n3607 , n403 );
buf ( n3608 , n416 );
and ( n3609 , n3607 , n3608 );
buf ( n3610 , n3609 );
buf ( n3611 , n3610 );
buf ( n3612 , n404 );
buf ( n3613 , n415 );
and ( n3614 , n3612 , n3613 );
buf ( n3615 , n3614 );
buf ( n3616 , n3615 );
xor ( n3617 , n3606 , n3611 );
xor ( n3618 , n3617 , n3616 );
buf ( n3619 , n3618 );
xor ( n3620 , n3606 , n3611 );
and ( n3621 , n3620 , n3616 );
and ( n3622 , n3606 , n3611 );
or ( n3623 , n3621 , n3622 );
buf ( n3624 , n3623 );
buf ( n3625 , n409 );
buf ( n3626 , n410 );
and ( n3627 , n3625 , n3626 );
buf ( n3628 , n3627 );
buf ( n3629 , n3628 );
and ( n3630 , n405 , n414 );
buf ( n3631 , n3630 );
buf ( n3632 , n407 );
buf ( n3633 , n412 );
and ( n3634 , n3632 , n3633 );
buf ( n3635 , n3634 );
buf ( n3636 , n3635 );
xor ( n3637 , n3629 , n3631 );
xor ( n3638 , n3637 , n3636 );
buf ( n3639 , n3638 );
xor ( n3640 , n3629 , n3631 );
and ( n3641 , n3640 , n3636 );
and ( n3642 , n3629 , n3631 );
or ( n3643 , n3641 , n3642 );
buf ( n3644 , n3643 );
buf ( n3645 , n3590 );
buf ( n3646 , n3543 );
not ( n3647 , n3545 );
not ( n3648 , n3647 );
not ( n3649 , n3552 );
not ( n3650 , n3649 );
not ( n3651 , n3650 );
or ( n3652 , n3648 , n3651 );
not ( n3653 , n3545 );
not ( n3654 , n3649 );
or ( n3655 , n3653 , n3654 );
nand ( n3656 , n3655 , n3564 );
nand ( n3657 , n3652 , n3656 );
not ( n3658 , n3657 );
nand ( n3659 , n389 , n391 );
not ( n3660 , n3659 );
and ( n3661 , n388 , n392 );
xor ( n3662 , n3660 , n3661 );
xor ( n3663 , n3431 , n3662 );
and ( n3664 , n390 , n391 );
xor ( n3665 , n3663 , n3664 );
not ( n3666 , n3665 );
xor ( n3667 , n3547 , n3548 );
and ( n3668 , n3667 , n3551 );
and ( n3669 , n3547 , n3548 );
or ( n3670 , n3668 , n3669 );
and ( n3671 , n3666 , n3670 );
nand ( n3672 , n3658 , n3671 );
not ( n3673 , n3647 );
not ( n3674 , n3552 );
or ( n3675 , n3673 , n3674 );
or ( n3676 , n3552 , n3647 );
nand ( n3677 , n3676 , n3564 );
nand ( n3678 , n3675 , n3677 );
not ( n3679 , n3678 );
not ( n3680 , n3670 );
and ( n3681 , n3665 , n3680 );
nand ( n3682 , n3679 , n3681 );
nand ( n3683 , n3665 , n3670 );
not ( n3684 , n3683 );
nand ( n3685 , n3666 , n3680 );
not ( n3686 , n3685 );
or ( n3687 , n3684 , n3686 );
nand ( n3688 , n3687 , n3657 );
nand ( n3689 , n3672 , n3682 , n3688 );
buf ( n3690 , n3689 );
buf ( n3691 , n393 );
and ( n3692 , n3690 , n3691 );
buf ( n3693 , n3692 );
buf ( n3694 , n3693 );
xor ( n3695 , n3646 , n3694 );
buf ( n3696 , n3499 );
buf ( n3697 , n3258 );
buf ( n3698 , n390 );
and ( n3699 , n3697 , n3698 );
buf ( n3700 , n3699 );
buf ( n3701 , n3700 );
xor ( n3702 , n3696 , n3701 );
buf ( n3703 , n3135 );
buf ( n3704 , n388 );
and ( n3705 , n3703 , n3704 );
buf ( n3706 , n3705 );
buf ( n3707 , n3706 );
not ( n3708 , n3122 );
not ( n3709 , n389 );
nor ( n3710 , n3708 , n3709 );
buf ( n3711 , n3710 );
xor ( n3712 , n3707 , n3711 );
buf ( n3713 , n3445 );
xor ( n3714 , n3712 , n3713 );
buf ( n3715 , n3714 );
buf ( n3716 , n3715 );
xor ( n3717 , n3702 , n3716 );
buf ( n3718 , n3717 );
buf ( n3719 , n3718 );
xor ( n3720 , n3695 , n3719 );
buf ( n3721 , n3720 );
buf ( n3722 , n3721 );
buf ( n3723 , n3579 );
buf ( n3724 , n408 );
buf ( n3725 , n411 );
and ( n3726 , n3724 , n3725 );
buf ( n3727 , n3726 );
buf ( n3728 , n3727 );
buf ( n3729 , n402 );
buf ( n3730 , n417 );
nand ( n3731 , n3729 , n3730 );
buf ( n3732 , n3731 );
buf ( n3733 , n386 );
buf ( n3734 , n393 );
nand ( n3735 , n3733 , n3734 );
buf ( n3736 , n3735 );
xor ( n3737 , n3732 , n3736 );
buf ( n3738 , n3737 );
xor ( n3739 , n3728 , n3738 );
and ( n3740 , n3478 , n3483 );
buf ( n3741 , n3740 );
buf ( n3742 , n3741 );
xor ( n3743 , n3739 , n3742 );
buf ( n3744 , n3743 );
buf ( n3745 , n3744 );
buf ( n3746 , n3397 );
buf ( n3747 , n391 );
and ( n3748 , n3746 , n3747 );
buf ( n3749 , n3748 );
buf ( n3750 , n3749 );
xor ( n3751 , n3745 , n3750 );
buf ( n3752 , n3512 );
xor ( n3753 , n3751 , n3752 );
buf ( n3754 , n3753 );
buf ( n3755 , n3754 );
xor ( n3756 , n3723 , n3755 );
buf ( n3757 , n3523 );
buf ( n3758 , n3565 );
buf ( n3759 , n392 );
and ( n3760 , n3758 , n3759 );
buf ( n3761 , n3760 );
buf ( n3762 , n3761 );
xor ( n3763 , n3757 , n3762 );
buf ( n3764 , n3468 );
buf ( n3765 , n3639 );
xor ( n3766 , n3764 , n3765 );
buf ( n3767 , n3619 );
xor ( n3768 , n3766 , n3767 );
buf ( n3769 , n3768 );
buf ( n3770 , n3769 );
xor ( n3771 , n3763 , n3770 );
buf ( n3772 , n3771 );
buf ( n3773 , n3772 );
xor ( n3774 , n3756 , n3773 );
buf ( n3775 , n3774 );
buf ( n3776 , n3775 );
xor ( n3777 , n3645 , n3722 );
xor ( n3778 , n3777 , n3776 );
buf ( n3779 , n3778 );
xor ( n3780 , n3645 , n3722 );
and ( n3781 , n3780 , n3776 );
and ( n3782 , n3645 , n3722 );
or ( n3783 , n3781 , n3782 );
buf ( n3784 , n3783 );
xor ( n3785 , n3728 , n3738 );
and ( n3786 , n3785 , n3742 );
and ( n3787 , n3728 , n3738 );
or ( n3788 , n3786 , n3787 );
buf ( n3789 , n3788 );
xor ( n3790 , n3707 , n3711 );
and ( n3791 , n3790 , n3713 );
or ( n3792 , n3791 , C0 );
buf ( n3793 , n3792 );
xor ( n3794 , n3764 , n3765 );
and ( n3795 , n3794 , n3767 );
and ( n3796 , n3764 , n3765 );
or ( n3797 , n3795 , n3796 );
buf ( n3798 , n3797 );
xor ( n3799 , n3696 , n3701 );
and ( n3800 , n3799 , n3716 );
and ( n3801 , n3696 , n3701 );
or ( n3802 , n3800 , n3801 );
buf ( n3803 , n3802 );
xor ( n3804 , n3745 , n3750 );
and ( n3805 , n3804 , n3752 );
and ( n3806 , n3745 , n3750 );
or ( n3807 , n3805 , n3806 );
buf ( n3808 , n3807 );
xor ( n3809 , n3757 , n3762 );
and ( n3810 , n3809 , n3770 );
and ( n3811 , n3757 , n3762 );
or ( n3812 , n3810 , n3811 );
buf ( n3813 , n3812 );
xor ( n3814 , n3646 , n3694 );
and ( n3815 , n3814 , n3719 );
and ( n3816 , n3646 , n3694 );
or ( n3817 , n3815 , n3816 );
buf ( n3818 , n3817 );
xor ( n3819 , n3723 , n3755 );
and ( n3820 , n3819 , n3773 );
and ( n3821 , n3723 , n3755 );
or ( n3822 , n3820 , n3821 );
buf ( n3823 , n3822 );
buf ( n3824 , n408 );
buf ( n3825 , n410 );
and ( n3826 , n3824 , n3825 );
buf ( n3827 , n3826 );
buf ( n3828 , n3827 );
buf ( n3829 , n403 );
buf ( n3830 , n415 );
and ( n3831 , n3829 , n3830 );
buf ( n3832 , n3831 );
buf ( n3833 , n3832 );
buf ( n3834 , n404 );
buf ( n3835 , n414 );
and ( n3836 , n3834 , n3835 );
buf ( n3837 , n3836 );
buf ( n3838 , n3837 );
xor ( n3839 , n3828 , n3833 );
xor ( n3840 , n3839 , n3838 );
buf ( n3841 , n3840 );
xor ( n3842 , n3828 , n3833 );
and ( n3843 , n3842 , n3838 );
and ( n3844 , n3828 , n3833 );
or ( n3845 , n3843 , n3844 );
buf ( n3846 , n3845 );
buf ( n3847 , n402 );
buf ( n3848 , n416 );
and ( n3849 , n3847 , n3848 );
buf ( n3850 , n3849 );
buf ( n3851 , n3850 );
buf ( n3852 , n407 );
buf ( n3853 , n411 );
and ( n3854 , n3852 , n3853 );
buf ( n3855 , n3854 );
buf ( n3856 , n3855 );
buf ( n3857 , n405 );
buf ( n3858 , n413 );
and ( n3859 , n3857 , n3858 );
buf ( n3860 , n3859 );
buf ( n3861 , n3860 );
xor ( n3862 , n3851 , n3856 );
xor ( n3863 , n3862 , n3861 );
buf ( n3864 , n3863 );
xor ( n3865 , n3851 , n3856 );
and ( n3866 , n3865 , n3861 );
and ( n3867 , n3851 , n3856 );
or ( n3868 , n3866 , n3867 );
buf ( n3869 , n3868 );
buf ( n3870 , n3864 );
buf ( n3871 , n3841 );
xor ( n3872 , n3870 , n3871 );
buf ( n3873 , n3789 );
xor ( n3874 , n3872 , n3873 );
buf ( n3875 , n3874 );
buf ( n3876 , n3875 );
buf ( n3877 , n3565 );
buf ( n3878 , n391 );
and ( n3879 , n3877 , n3878 );
buf ( n3880 , n3879 );
buf ( n3881 , n3880 );
xor ( n3882 , n3876 , n3881 );
buf ( n3883 , n3803 );
xor ( n3884 , n3882 , n3883 );
buf ( n3885 , n3884 );
buf ( n3886 , n3885 );
buf ( n3887 , n3818 );
buf ( n3888 , n3689 );
buf ( n3889 , n392 );
and ( n3890 , n3888 , n3889 );
buf ( n3891 , n3890 );
buf ( n3892 , n3891 );
buf ( n3893 , n3808 );
xor ( n3894 , n3892 , n3893 );
buf ( n3895 , n406 );
buf ( n3896 , n412 );
and ( n3897 , n3895 , n3896 );
buf ( n3898 , n3897 );
buf ( n3899 , n3898 );
buf ( n3900 , n3736 );
buf ( n3901 , n3732 );
nor ( n3902 , n3900 , n3901 );
buf ( n3903 , n3902 );
buf ( n3904 , n3903 );
xor ( n3905 , n3899 , n3904 );
buf ( n3906 , n3122 );
not ( n3907 , n3906 );
buf ( n3908 , n388 );
not ( n3909 , n3908 );
buf ( n3910 , n3909 );
buf ( n3911 , n3910 );
nor ( n3912 , n3907 , n3911 );
buf ( n3913 , n3912 );
buf ( n3914 , n3913 );
xor ( n3915 , n3905 , n3914 );
buf ( n3916 , n3915 );
buf ( n3917 , n3916 );
buf ( n3918 , n3793 );
xor ( n3919 , n3917 , n3918 );
not ( n3920 , n3258 );
buf ( n3921 , n3920 );
buf ( n3922 , n3709 );
nor ( n3923 , n3921 , n3922 );
buf ( n3924 , n3923 );
buf ( n3925 , n3924 );
xor ( n3926 , n3919 , n3925 );
buf ( n3927 , n3926 );
buf ( n3928 , n3927 );
xor ( n3929 , n3894 , n3928 );
buf ( n3930 , n3929 );
buf ( n3931 , n3930 );
xor ( n3932 , n3886 , n3887 );
xor ( n3933 , n3932 , n3931 );
buf ( n3934 , n3933 );
xor ( n3935 , n3886 , n3887 );
and ( n3936 , n3935 , n3931 );
and ( n3937 , n3886 , n3887 );
or ( n3938 , n3936 , n3937 );
buf ( n3939 , n3938 );
xor ( n3940 , n3431 , n3662 );
and ( n3941 , n3940 , n3664 );
and ( n3942 , n3431 , n3662 );
or ( n3943 , n3941 , n3942 );
and ( n3944 , n389 , n390 );
xor ( n3945 , n389 , n3944 );
and ( n3946 , n3660 , n3661 );
xor ( n3947 , n3945 , n3946 );
nand ( n3948 , n387 , n392 );
not ( n3949 , n3948 );
and ( n3950 , n386 , n393 );
xor ( n3951 , n3949 , n3950 );
and ( n3952 , n388 , n391 );
xor ( n3953 , n3951 , n3952 );
xor ( n3954 , n3947 , n3953 );
not ( n3955 , n3954 );
xor ( n3956 , n3943 , n3955 );
not ( n3957 , n3685 );
not ( n3958 , n3678 );
or ( n3959 , n3957 , n3958 );
buf ( n3960 , n3683 );
nand ( n3961 , n3959 , n3960 );
xnor ( n3962 , n3956 , n3961 );
buf ( n3963 , n3962 );
buf ( n3964 , n3963 );
buf ( n3965 , n393 );
and ( n3966 , n3964 , n3965 );
buf ( n3967 , n3966 );
buf ( n3968 , n3967 );
buf ( n3969 , n3798 );
buf ( n3970 , n3397 );
buf ( n3971 , n390 );
and ( n3972 , n3970 , n3971 );
buf ( n3973 , n3972 );
buf ( n3974 , n3973 );
xor ( n3975 , n3969 , n3974 );
buf ( n3976 , n3135 );
buf ( n3977 , n387 );
and ( n3978 , n3976 , n3977 );
buf ( n3979 , n3978 );
buf ( n3980 , n3979 );
buf ( n3981 , n3624 );
xor ( n3982 , n3980 , n3981 );
buf ( n3983 , n3644 );
xor ( n3984 , n3982 , n3983 );
buf ( n3985 , n3984 );
buf ( n3986 , n3985 );
xor ( n3987 , n3975 , n3986 );
buf ( n3988 , n3987 );
buf ( n3989 , n3988 );
xor ( n3990 , n3968 , n3989 );
buf ( n3991 , n3813 );
xor ( n3992 , n3990 , n3991 );
buf ( n3993 , n3992 );
buf ( n3994 , n3993 );
buf ( n3995 , n3823 );
buf ( n3996 , n3934 );
xor ( n3997 , n3994 , n3995 );
xor ( n3998 , n3997 , n3996 );
buf ( n3999 , n3998 );
xor ( n4000 , n3994 , n3995 );
and ( n4001 , n4000 , n3996 );
and ( n4002 , n3994 , n3995 );
or ( n4003 , n4001 , n4002 );
buf ( n4004 , n4003 );
xor ( n4005 , n3899 , n3904 );
and ( n4006 , n4005 , n3914 );
and ( n4007 , n3899 , n3904 );
or ( n4008 , n4006 , n4007 );
buf ( n4009 , n4008 );
xor ( n4010 , n3980 , n3981 );
and ( n4011 , n4010 , n3983 );
and ( n4012 , n3980 , n3981 );
or ( n4013 , n4011 , n4012 );
buf ( n4014 , n4013 );
xor ( n4015 , n3870 , n3871 );
and ( n4016 , n4015 , n3873 );
and ( n4017 , n3870 , n3871 );
or ( n4018 , n4016 , n4017 );
buf ( n4019 , n4018 );
xor ( n4020 , n3917 , n3918 );
and ( n4021 , n4020 , n3925 );
and ( n4022 , n3917 , n3918 );
or ( n4023 , n4021 , n4022 );
buf ( n4024 , n4023 );
xor ( n4025 , n3969 , n3974 );
and ( n4026 , n4025 , n3986 );
and ( n4027 , n3969 , n3974 );
or ( n4028 , n4026 , n4027 );
buf ( n4029 , n4028 );
xor ( n4030 , n3876 , n3881 );
and ( n4031 , n4030 , n3883 );
and ( n4032 , n3876 , n3881 );
or ( n4033 , n4031 , n4032 );
buf ( n4034 , n4033 );
xor ( n4035 , n3892 , n3893 );
and ( n4036 , n4035 , n3928 );
and ( n4037 , n3892 , n3893 );
or ( n4038 , n4036 , n4037 );
buf ( n4039 , n4038 );
xor ( n4040 , n3968 , n3989 );
and ( n4041 , n4040 , n3991 );
and ( n4042 , n3968 , n3989 );
or ( n4043 , n4041 , n4042 );
buf ( n4044 , n4043 );
buf ( n4045 , n402 );
buf ( n4046 , n415 );
and ( n4047 , n4045 , n4046 );
buf ( n4048 , n4047 );
buf ( n4049 , n4048 );
buf ( n4050 , n403 );
buf ( n4051 , n414 );
and ( n4052 , n4050 , n4051 );
buf ( n4053 , n4052 );
buf ( n4054 , n4053 );
buf ( n4055 , n406 );
buf ( n4056 , n411 );
and ( n4057 , n4055 , n4056 );
buf ( n4058 , n4057 );
buf ( n4059 , n4058 );
xor ( n4060 , n4049 , n4054 );
xor ( n4061 , n4060 , n4059 );
buf ( n4062 , n4061 );
xor ( n4063 , n4049 , n4054 );
and ( n4064 , n4063 , n4059 );
and ( n4065 , n4049 , n4054 );
or ( n4066 , n4064 , n4065 );
buf ( n4067 , n4066 );
buf ( n4068 , n404 );
buf ( n4069 , n413 );
and ( n4070 , n4068 , n4069 );
buf ( n4071 , n4070 );
buf ( n4072 , n4071 );
buf ( n4073 , n405 );
buf ( n4074 , n412 );
and ( n4075 , n4073 , n4074 );
buf ( n4076 , n4075 );
buf ( n4077 , n4076 );
buf ( n4078 , n407 );
buf ( n4079 , n410 );
and ( n4080 , n4078 , n4079 );
buf ( n4081 , n4080 );
buf ( n4082 , n4081 );
xor ( n4083 , n4072 , n4077 );
xor ( n4084 , n4083 , n4082 );
buf ( n4085 , n4084 );
xor ( n4086 , n4072 , n4077 );
and ( n4087 , n4086 , n4082 );
and ( n4088 , n4072 , n4077 );
or ( n4089 , n4087 , n4088 );
buf ( n4090 , n4089 );
buf ( n4091 , n4044 );
buf ( n4092 , n4029 );
buf ( n4093 , n3689 );
buf ( n4094 , n391 );
and ( n4095 , n4093 , n4094 );
buf ( n4096 , n4095 );
buf ( n4097 , n4096 );
xor ( n4098 , n4092 , n4097 );
buf ( n4099 , n4009 );
buf ( n4100 , n3135 );
buf ( n4101 , n386 );
and ( n4102 , n4100 , n4101 );
buf ( n4103 , n4102 );
buf ( n4104 , n4103 );
buf ( n4105 , n3122 );
buf ( n4106 , n387 );
and ( n4107 , n4105 , n4106 );
buf ( n4108 , n4107 );
buf ( n4109 , n4108 );
xor ( n4110 , n4104 , n4109 );
buf ( n4111 , n3869 );
xor ( n4112 , n4110 , n4111 );
buf ( n4113 , n4112 );
buf ( n4114 , n4113 );
xor ( n4115 , n4099 , n4114 );
buf ( n4116 , n3920 );
buf ( n4117 , n3910 );
nor ( n4118 , n4116 , n4117 );
buf ( n4119 , n4118 );
buf ( n4120 , n4119 );
xor ( n4121 , n4115 , n4120 );
buf ( n4122 , n4121 );
buf ( n4123 , n4122 );
xor ( n4124 , n4098 , n4123 );
buf ( n4125 , n4124 );
buf ( n4126 , n4125 );
buf ( n4127 , n3963 );
buf ( n4128 , n392 );
and ( n4129 , n4127 , n4128 );
buf ( n4130 , n4129 );
buf ( n4131 , n4130 );
buf ( n4132 , n4014 );
buf ( n4133 , n3397 );
buf ( n4134 , n389 );
and ( n4135 , n4133 , n4134 );
buf ( n4136 , n4135 );
buf ( n4137 , n4136 );
xor ( n4138 , n4132 , n4137 );
buf ( n4139 , n4019 );
xor ( n4140 , n4138 , n4139 );
buf ( n4141 , n4140 );
buf ( n4142 , n4141 );
xor ( n4143 , n4131 , n4142 );
not ( n4144 , n3954 );
not ( n4145 , n3943 );
nand ( n4146 , n4144 , n4145 );
not ( n4147 , n4146 );
not ( n4148 , n3961 );
or ( n4149 , n4147 , n4148 );
nand ( n4150 , n3954 , n3943 );
nand ( n4151 , n4149 , n4150 );
buf ( n4152 , n4151 );
and ( n4153 , n389 , n3944 );
xor ( n4154 , n3949 , n3950 );
and ( n4155 , n4154 , n3952 );
and ( n4156 , n3949 , n3950 );
or ( n4157 , n4155 , n4156 );
xor ( n4158 , n4153 , n4157 );
and ( n4159 , n388 , n390 );
and ( n4160 , n387 , n391 );
xor ( n4161 , n4159 , n4160 );
and ( n4162 , n386 , n392 );
xor ( n4163 , n4161 , n4162 );
xor ( n4164 , n4158 , n4163 );
not ( n4165 , n4164 );
xor ( n4166 , n3945 , n3946 );
and ( n4167 , n4166 , n3953 );
and ( n4168 , n3945 , n3946 );
or ( n4169 , n4167 , n4168 );
not ( n4170 , n4169 );
nand ( n4171 , n4165 , n4170 );
nand ( n4172 , n4164 , n4169 );
nand ( n4173 , n4171 , n4172 );
not ( n4174 , n4173 );
and ( n4175 , n4152 , n4174 );
not ( n4176 , n4152 );
and ( n4177 , n4176 , n4173 );
nor ( n4178 , n4175 , n4177 );
buf ( n4179 , n4178 );
buf ( n4180 , n4179 );
buf ( n4181 , n4180 );
buf ( n4182 , n4181 );
buf ( n4183 , n393 );
and ( n4184 , n4182 , n4183 );
buf ( n4185 , n4184 );
buf ( n4186 , n4185 );
xor ( n4187 , n4143 , n4186 );
buf ( n4188 , n4187 );
buf ( n4189 , n4188 );
xor ( n4190 , n4091 , n4126 );
xor ( n4191 , n4190 , n4189 );
buf ( n4192 , n4191 );
xor ( n4193 , n4091 , n4126 );
and ( n4194 , n4193 , n4189 );
and ( n4195 , n4091 , n4126 );
or ( n4196 , n4194 , n4195 );
buf ( n4197 , n4196 );
buf ( n4198 , n4034 );
buf ( n4199 , n3846 );
buf ( n4200 , n4085 );
xor ( n4201 , n4199 , n4200 );
buf ( n4202 , n4062 );
xor ( n4203 , n4201 , n4202 );
buf ( n4204 , n4203 );
buf ( n4205 , n4204 );
buf ( n4206 , n3565 );
buf ( n4207 , n390 );
and ( n4208 , n4206 , n4207 );
buf ( n4209 , n4208 );
buf ( n4210 , n4209 );
xor ( n4211 , n4205 , n4210 );
buf ( n4212 , n4024 );
xor ( n4213 , n4211 , n4212 );
buf ( n4214 , n4213 );
buf ( n4215 , n4214 );
xor ( n4216 , n4198 , n4215 );
buf ( n4217 , n4039 );
xor ( n4218 , n4216 , n4217 );
buf ( n4219 , n4218 );
buf ( n4220 , n4219 );
buf ( n4221 , n3939 );
buf ( n4222 , n4192 );
xor ( n4223 , n4220 , n4221 );
xor ( n4224 , n4223 , n4222 );
buf ( n4225 , n4224 );
xor ( n4226 , n4220 , n4221 );
and ( n4227 , n4226 , n4222 );
and ( n4228 , n4220 , n4221 );
or ( n4229 , n4227 , n4228 );
buf ( n4230 , n4229 );
xor ( n4231 , n4104 , n4109 );
and ( n4232 , n4231 , n4111 );
or ( n4233 , n4232 , C0 );
buf ( n4234 , n4233 );
xor ( n4235 , n4199 , n4200 );
and ( n4236 , n4235 , n4202 );
and ( n4237 , n4199 , n4200 );
or ( n4238 , n4236 , n4237 );
buf ( n4239 , n4238 );
xor ( n4240 , n4099 , n4114 );
and ( n4241 , n4240 , n4120 );
and ( n4242 , n4099 , n4114 );
or ( n4243 , n4241 , n4242 );
buf ( n4244 , n4243 );
xor ( n4245 , n4132 , n4137 );
and ( n4246 , n4245 , n4139 );
and ( n4247 , n4132 , n4137 );
or ( n4248 , n4246 , n4247 );
buf ( n4249 , n4248 );
xor ( n4250 , n4205 , n4210 );
and ( n4251 , n4250 , n4212 );
and ( n4252 , n4205 , n4210 );
or ( n4253 , n4251 , n4252 );
buf ( n4254 , n4253 );
xor ( n4255 , n4092 , n4097 );
and ( n4256 , n4255 , n4123 );
and ( n4257 , n4092 , n4097 );
or ( n4258 , n4256 , n4257 );
buf ( n4259 , n4258 );
xor ( n4260 , n4131 , n4142 );
and ( n4261 , n4260 , n4186 );
and ( n4262 , n4131 , n4142 );
or ( n4263 , n4261 , n4262 );
buf ( n4264 , n4263 );
xor ( n4265 , n4198 , n4215 );
and ( n4266 , n4265 , n4217 );
and ( n4267 , n4198 , n4215 );
or ( n4268 , n4266 , n4267 );
buf ( n4269 , n4268 );
buf ( n4270 , n406 );
buf ( n4271 , n410 );
and ( n4272 , n4270 , n4271 );
buf ( n4273 , n4272 );
buf ( n4274 , n4273 );
buf ( n4275 , n404 );
buf ( n4276 , n412 );
and ( n4277 , n4275 , n4276 );
buf ( n4278 , n4277 );
buf ( n4279 , n4278 );
buf ( n4280 , n405 );
buf ( n4281 , n411 );
and ( n4282 , n4280 , n4281 );
buf ( n4283 , n4282 );
buf ( n4284 , n4283 );
xor ( n4285 , n4274 , n4279 );
xor ( n4286 , n4285 , n4284 );
buf ( n4287 , n4286 );
xor ( n4288 , n4274 , n4279 );
and ( n4289 , n4288 , n4284 );
and ( n4290 , n4274 , n4279 );
or ( n4291 , n4289 , n4290 );
buf ( n4292 , n4291 );
buf ( n4293 , n3122 );
buf ( n4294 , n386 );
and ( n4295 , n4293 , n4294 );
buf ( n4296 , n4295 );
buf ( n4297 , n4296 );
buf ( n4298 , n402 );
buf ( n4299 , n414 );
and ( n4300 , n4298 , n4299 );
buf ( n4301 , n4300 );
buf ( n4302 , n4301 );
buf ( n4303 , n403 );
buf ( n4304 , n413 );
and ( n4305 , n4303 , n4304 );
buf ( n4306 , n4305 );
buf ( n4307 , n4306 );
xor ( n4308 , n4302 , n4307 );
buf ( n4309 , n4308 );
buf ( n4310 , n4309 );
buf ( n4311 , n4090 );
xor ( n4312 , n4297 , n4310 );
xor ( n4313 , n4312 , n4311 );
buf ( n4314 , n4313 );
xor ( n4315 , n4297 , n4310 );
and ( n4316 , n4315 , n4311 );
and ( n4317 , n4297 , n4310 );
or ( n4318 , n4316 , n4317 );
buf ( n4319 , n4318 );
buf ( n4320 , n4259 );
buf ( n4321 , n4244 );
buf ( n4322 , n3257 );
not ( n4323 , n4322 );
buf ( n4324 , n387 );
not ( n4325 , n4324 );
buf ( n4326 , n4325 );
buf ( n4327 , n4326 );
nor ( n4328 , n4323 , n4327 );
buf ( n4329 , n4328 );
buf ( n4330 , n4329 );
buf ( n4331 , n4314 );
xor ( n4332 , n4330 , n4331 );
buf ( n4333 , n4239 );
xor ( n4334 , n4332 , n4333 );
buf ( n4335 , n4334 );
buf ( n4336 , n4335 );
xor ( n4337 , n4321 , n4336 );
not ( n4338 , n390 );
buf ( n4339 , n3689 );
not ( n4340 , n4339 );
buf ( n4341 , n4340 );
nor ( n4342 , n4338 , n4341 );
buf ( n4343 , n4342 );
xor ( n4344 , n4337 , n4343 );
buf ( n4345 , n4344 );
buf ( n4346 , n4345 );
xor ( n4347 , n4320 , n4346 );
buf ( n4348 , n4264 );
xor ( n4349 , n4347 , n4348 );
buf ( n4350 , n4349 );
buf ( n4351 , n4350 );
buf ( n4352 , n4197 );
buf ( n4353 , n3962 );
buf ( n4354 , n391 );
and ( n4355 , n4353 , n4354 );
buf ( n4356 , n4355 );
buf ( n4357 , n4356 );
buf ( n4358 , n4249 );
xor ( n4359 , n4357 , n4358 );
buf ( n4360 , n4254 );
xor ( n4361 , n4359 , n4360 );
buf ( n4362 , n4361 );
buf ( n4363 , n4362 );
buf ( n4364 , n4181 );
buf ( n4365 , n392 );
and ( n4366 , n4364 , n4365 );
buf ( n4367 , n4366 );
buf ( n4368 , n4367 );
buf ( n4369 , n3397 );
buf ( n4370 , n388 );
and ( n4371 , n4369 , n4370 );
buf ( n4372 , n4371 );
buf ( n4373 , n4372 );
buf ( n4374 , n3565 );
buf ( n4375 , n389 );
and ( n4376 , n4374 , n4375 );
buf ( n4377 , n4376 );
buf ( n4378 , n4377 );
xor ( n4379 , n4373 , n4378 );
buf ( n4380 , n4067 );
buf ( n4381 , n4287 );
xor ( n4382 , n4380 , n4381 );
buf ( n4383 , n4234 );
xor ( n4384 , n4382 , n4383 );
buf ( n4385 , n4384 );
buf ( n4386 , n4385 );
xor ( n4387 , n4379 , n4386 );
buf ( n4388 , n4387 );
buf ( n4389 , n4388 );
xor ( n4390 , n4368 , n4389 );
not ( n4391 , n4171 );
not ( n4392 , n4152 );
or ( n4393 , n4391 , n4392 );
nand ( n4394 , n4393 , n4172 );
xor ( n4395 , n4153 , n4157 );
and ( n4396 , n4395 , n4163 );
and ( n4397 , n4153 , n4157 );
or ( n4398 , n4396 , n4397 );
and ( n4399 , n387 , n390 );
xor ( n4400 , n4159 , n4160 );
and ( n4401 , n4400 , n4162 );
and ( n4402 , n4159 , n4160 );
or ( n4403 , n4401 , n4402 );
xor ( n4404 , n4399 , n4403 );
and ( n4405 , n388 , n389 );
xor ( n4406 , n388 , n4405 );
and ( n4407 , n386 , n391 );
xor ( n4408 , n4406 , n4407 );
xor ( n4409 , n4404 , n4408 );
buf ( n4410 , n4409 );
xor ( n4411 , n4398 , n4410 );
buf ( n4412 , n4411 );
and ( n4413 , n4394 , n4412 );
not ( n4414 , n4394 );
not ( n4415 , n4411 );
and ( n4416 , n4414 , n4415 );
nor ( n4417 , n4413 , n4416 );
buf ( n4418 , n4417 );
buf ( n4419 , n393 );
and ( n4420 , n4418 , n4419 );
buf ( n4421 , n4420 );
buf ( n4422 , n4421 );
xor ( n4423 , n4390 , n4422 );
buf ( n4424 , n4423 );
buf ( n4425 , n4424 );
xor ( n4426 , n4363 , n4425 );
buf ( n4427 , n4269 );
xor ( n4428 , n4426 , n4427 );
buf ( n4429 , n4428 );
buf ( n4430 , n4429 );
xor ( n4431 , n4351 , n4352 );
xor ( n4432 , n4431 , n4430 );
buf ( n4433 , n4432 );
xor ( n4434 , n4351 , n4352 );
and ( n4435 , n4434 , n4430 );
and ( n4436 , n4351 , n4352 );
or ( n4437 , n4435 , n4436 );
buf ( n4438 , n4437 );
xor ( n4439 , n4380 , n4381 );
and ( n4440 , n4439 , n4383 );
and ( n4441 , n4380 , n4381 );
or ( n4442 , n4440 , n4441 );
buf ( n4443 , n4442 );
xor ( n4444 , n4330 , n4331 );
and ( n4445 , n4444 , n4333 );
and ( n4446 , n4330 , n4331 );
or ( n4447 , n4445 , n4446 );
buf ( n4448 , n4447 );
xor ( n4449 , n4373 , n4378 );
and ( n4450 , n4449 , n4386 );
and ( n4451 , n4373 , n4378 );
or ( n4452 , n4450 , n4451 );
buf ( n4453 , n4452 );
xor ( n4454 , n4321 , n4336 );
and ( n4455 , n4454 , n4343 );
and ( n4456 , n4321 , n4336 );
or ( n4457 , n4455 , n4456 );
buf ( n4458 , n4457 );
xor ( n4459 , n4357 , n4358 );
and ( n4460 , n4459 , n4360 );
and ( n4461 , n4357 , n4358 );
or ( n4462 , n4460 , n4461 );
buf ( n4463 , n4462 );
xor ( n4464 , n4368 , n4389 );
and ( n4465 , n4464 , n4422 );
and ( n4466 , n4368 , n4389 );
or ( n4467 , n4465 , n4466 );
buf ( n4468 , n4467 );
xor ( n4469 , n4320 , n4346 );
and ( n4470 , n4469 , n4348 );
and ( n4471 , n4320 , n4346 );
or ( n4472 , n4470 , n4471 );
buf ( n4473 , n4472 );
xor ( n4474 , n4363 , n4425 );
and ( n4475 , n4474 , n4427 );
and ( n4476 , n4363 , n4425 );
or ( n4477 , n4475 , n4476 );
buf ( n4478 , n4477 );
buf ( n4479 , n402 );
buf ( n4480 , n413 );
and ( n4481 , n4479 , n4480 );
buf ( n4482 , n4481 );
buf ( n4483 , n4482 );
buf ( n4484 , n403 );
buf ( n4485 , n412 );
and ( n4486 , n4484 , n4485 );
buf ( n4487 , n4486 );
buf ( n4488 , n4487 );
buf ( n4489 , n404 );
buf ( n4490 , n411 );
and ( n4491 , n4489 , n4490 );
buf ( n4492 , n4491 );
buf ( n4493 , n4492 );
xor ( n4494 , n4483 , n4488 );
xor ( n4495 , n4494 , n4493 );
buf ( n4496 , n4495 );
xor ( n4497 , n4483 , n4488 );
and ( n4498 , n4497 , n4493 );
and ( n4499 , n4483 , n4488 );
or ( n4500 , n4498 , n4499 );
buf ( n4501 , n4500 );
buf ( n4502 , n405 );
buf ( n4503 , n410 );
and ( n4504 , n4502 , n4503 );
buf ( n4505 , n4504 );
buf ( n4506 , n4505 );
and ( n4507 , n4302 , n4307 );
buf ( n4508 , n4507 );
buf ( n4509 , n4508 );
buf ( n4510 , n4292 );
xor ( n4511 , n4506 , n4509 );
xor ( n4512 , n4511 , n4510 );
buf ( n4513 , n4512 );
xor ( n4514 , n4506 , n4509 );
and ( n4515 , n4514 , n4510 );
and ( n4516 , n4506 , n4509 );
or ( n4517 , n4515 , n4516 );
buf ( n4518 , n4517 );
buf ( n4519 , n4463 );
buf ( n4520 , n4448 );
buf ( n4521 , n3257 );
buf ( n4522 , n386 );
and ( n4523 , n4521 , n4522 );
buf ( n4524 , n4523 );
buf ( n4525 , n4524 );
buf ( n4526 , n3397 );
buf ( n4527 , n387 );
and ( n4528 , n4526 , n4527 );
buf ( n4529 , n4528 );
buf ( n4530 , n4529 );
xor ( n4531 , n4525 , n4530 );
buf ( n4532 , n3565 );
buf ( n4533 , n388 );
and ( n4534 , n4532 , n4533 );
buf ( n4535 , n4534 );
buf ( n4536 , n4535 );
xor ( n4537 , n4531 , n4536 );
buf ( n4538 , n4537 );
buf ( n4539 , n4538 );
xor ( n4540 , n4520 , n4539 );
and ( n4541 , n390 , n3962 );
buf ( n4542 , n4541 );
xor ( n4543 , n4540 , n4542 );
buf ( n4544 , n4543 );
buf ( n4545 , n4544 );
xor ( n4546 , n4519 , n4545 );
buf ( n4547 , n4468 );
xor ( n4548 , n4546 , n4547 );
buf ( n4549 , n4548 );
buf ( n4550 , n4549 );
buf ( n4551 , n4478 );
buf ( n4552 , n4453 );
buf ( n4553 , n4181 );
buf ( n4554 , n391 );
and ( n4555 , n4553 , n4554 );
buf ( n4556 , n4555 );
buf ( n4557 , n4556 );
xor ( n4558 , n4552 , n4557 );
buf ( n4559 , n4417 );
buf ( n4560 , n392 );
and ( n4561 , n4559 , n4560 );
buf ( n4562 , n4561 );
buf ( n4563 , n4562 );
xor ( n4564 , n4558 , n4563 );
buf ( n4565 , n4564 );
buf ( n4566 , n4565 );
buf ( n4567 , n4458 );
not ( n4568 , n4164 );
not ( n4569 , n4169 );
and ( n4570 , n4568 , n4569 );
nor ( n4571 , n4409 , n4398 );
nor ( n4572 , n4570 , n4571 );
not ( n4573 , n4572 );
not ( n4574 , n4151 );
or ( n4575 , n4573 , n4574 );
not ( n4576 , n4409 );
not ( n4577 , n4398 );
nand ( n4578 , n4576 , n4577 );
not ( n4579 , n4164 );
nor ( n4580 , n4579 , n4170 );
and ( n4581 , n4578 , n4580 );
nor ( n4582 , n4576 , n4577 );
nor ( n4583 , n4581 , n4582 );
nand ( n4584 , n4575 , n4583 );
buf ( n4585 , n4584 );
and ( n4586 , n387 , n389 );
and ( n4587 , n386 , n390 );
xor ( n4588 , n4586 , n4587 );
xor ( n4589 , n388 , n4405 );
and ( n4590 , n4589 , n4407 );
and ( n4591 , n388 , n4405 );
or ( n4592 , n4590 , n4591 );
xor ( n4593 , n4588 , n4592 );
xor ( n4594 , n4399 , n4403 );
and ( n4595 , n4594 , n4408 );
and ( n4596 , n4399 , n4403 );
or ( n4597 , n4595 , n4596 );
not ( n4598 , n4597 );
and ( n4599 , n4593 , n4598 );
not ( n4600 , n4593 );
and ( n4601 , n4600 , n4597 );
nor ( n4602 , n4599 , n4601 );
not ( n4603 , n4602 );
and ( n4604 , n4585 , n4603 );
not ( n4605 , n4585 );
and ( n4606 , n4605 , n4602 );
nor ( n4607 , n4604 , n4606 );
buf ( n4608 , n4607 );
buf ( n4609 , n393 );
and ( n4610 , n4608 , n4609 );
buf ( n4611 , n4610 );
buf ( n4612 , n4611 );
xor ( n4613 , n4567 , n4612 );
buf ( n4614 , n4443 );
buf ( n4615 , n4496 );
buf ( n4616 , n4319 );
xor ( n4617 , n4615 , n4616 );
buf ( n4618 , n4513 );
xor ( n4619 , n4617 , n4618 );
buf ( n4620 , n4619 );
buf ( n4621 , n4620 );
xor ( n4622 , n4614 , n4621 );
buf ( n4623 , n4341 );
buf ( n4624 , n3709 );
nor ( n4625 , n4623 , n4624 );
buf ( n4626 , n4625 );
buf ( n4627 , n4626 );
xor ( n4628 , n4622 , n4627 );
buf ( n4629 , n4628 );
buf ( n4630 , n4629 );
xor ( n4631 , n4613 , n4630 );
buf ( n4632 , n4631 );
buf ( n4633 , n4632 );
xor ( n4634 , n4566 , n4633 );
buf ( n4635 , n4473 );
xor ( n4636 , n4634 , n4635 );
buf ( n4637 , n4636 );
buf ( n4638 , n4637 );
xor ( n4639 , n4550 , n4551 );
xor ( n4640 , n4639 , n4638 );
buf ( n4641 , n4640 );
xor ( n4642 , n4550 , n4551 );
and ( n4643 , n4642 , n4638 );
and ( n4644 , n4550 , n4551 );
or ( n4645 , n4643 , n4644 );
buf ( n4646 , n4645 );
xor ( n4647 , n4615 , n4616 );
and ( n4648 , n4647 , n4618 );
and ( n4649 , n4615 , n4616 );
or ( n4650 , n4648 , n4649 );
buf ( n4651 , n4650 );
xor ( n4652 , n4525 , n4530 );
and ( n4653 , n4652 , n4536 );
and ( n4654 , n4525 , n4530 );
or ( n4655 , n4653 , n4654 );
buf ( n4656 , n4655 );
xor ( n4657 , n4614 , n4621 );
and ( n4658 , n4657 , n4627 );
and ( n4659 , n4614 , n4621 );
or ( n4660 , n4658 , n4659 );
buf ( n4661 , n4660 );
xor ( n4662 , n4520 , n4539 );
and ( n4663 , n4662 , n4542 );
and ( n4664 , n4520 , n4539 );
or ( n4665 , n4663 , n4664 );
buf ( n4666 , n4665 );
xor ( n4667 , n4552 , n4557 );
and ( n4668 , n4667 , n4563 );
and ( n4669 , n4552 , n4557 );
or ( n4670 , n4668 , n4669 );
buf ( n4671 , n4670 );
xor ( n4672 , n4567 , n4612 );
and ( n4673 , n4672 , n4630 );
and ( n4674 , n4567 , n4612 );
or ( n4675 , n4673 , n4674 );
buf ( n4676 , n4675 );
xor ( n4677 , n4519 , n4545 );
and ( n4678 , n4677 , n4547 );
and ( n4679 , n4519 , n4545 );
or ( n4680 , n4678 , n4679 );
buf ( n4681 , n4680 );
xor ( n4682 , n4566 , n4633 );
and ( n4683 , n4682 , n4635 );
and ( n4684 , n4566 , n4633 );
or ( n4685 , n4683 , n4684 );
buf ( n4686 , n4685 );
buf ( n4687 , n402 );
buf ( n4688 , n412 );
and ( n4689 , n4687 , n4688 );
buf ( n4690 , n4689 );
buf ( n4691 , n4690 );
buf ( n4692 , n403 );
buf ( n4693 , n411 );
and ( n4694 , n4692 , n4693 );
buf ( n4695 , n4694 );
buf ( n4696 , n4695 );
buf ( n4697 , n404 );
buf ( n4698 , n410 );
and ( n4699 , n4697 , n4698 );
buf ( n4700 , n4699 );
buf ( n4701 , n4700 );
xor ( n4702 , n4691 , n4696 );
xor ( n4703 , n4702 , n4701 );
buf ( n4704 , n4703 );
xor ( n4705 , n4691 , n4696 );
and ( n4706 , n4705 , n4701 );
and ( n4707 , n4691 , n4696 );
or ( n4708 , n4706 , n4707 );
buf ( n4709 , n4708 );
buf ( n4710 , n4501 );
buf ( n4711 , n4704 );
buf ( n4712 , n4518 );
xor ( n4713 , n4710 , n4711 );
xor ( n4714 , n4713 , n4712 );
buf ( n4715 , n4714 );
xor ( n4716 , n4710 , n4711 );
and ( n4717 , n4716 , n4712 );
and ( n4718 , n4710 , n4711 );
or ( n4719 , n4717 , n4718 );
buf ( n4720 , n4719 );
buf ( n4721 , n3397 );
buf ( n4722 , n386 );
and ( n4723 , n4721 , n4722 );
buf ( n4724 , n4723 );
buf ( n4725 , n4724 );
buf ( n4726 , n3565 );
buf ( n4727 , n387 );
and ( n4728 , n4726 , n4727 );
buf ( n4729 , n4728 );
buf ( n4730 , n4729 );
buf ( n4731 , n4651 );
xor ( n4732 , n4725 , n4730 );
xor ( n4733 , n4732 , n4731 );
buf ( n4734 , n4733 );
xor ( n4735 , n4725 , n4730 );
and ( n4736 , n4735 , n4731 );
and ( n4737 , n4725 , n4730 );
or ( n4738 , n4736 , n4737 );
buf ( n4739 , n4738 );
buf ( n4740 , n4715 );
buf ( n4741 , n3689 );
buf ( n4742 , n388 );
and ( n4743 , n4741 , n4742 );
buf ( n4744 , n4743 );
buf ( n4745 , n4744 );
buf ( n4746 , n4656 );
xor ( n4747 , n4740 , n4745 );
xor ( n4748 , n4747 , n4746 );
buf ( n4749 , n4748 );
xor ( n4750 , n4740 , n4745 );
and ( n4751 , n4750 , n4746 );
and ( n4752 , n4740 , n4745 );
or ( n4753 , n4751 , n4752 );
buf ( n4754 , n4753 );
and ( n4755 , n3963 , n389 );
buf ( n4756 , n4755 );
buf ( n4757 , n4734 );
buf ( n4758 , n4181 );
buf ( n4759 , n390 );
and ( n4760 , n4758 , n4759 );
buf ( n4761 , n4760 );
buf ( n4762 , n4761 );
xor ( n4763 , n4756 , n4757 );
xor ( n4764 , n4763 , n4762 );
buf ( n4765 , n4764 );
xor ( n4766 , n4756 , n4757 );
and ( n4767 , n4766 , n4762 );
and ( n4768 , n4756 , n4757 );
or ( n4769 , n4767 , n4768 );
buf ( n4770 , n4769 );
buf ( n4771 , n4661 );
and ( n4772 , n4417 , n391 );
buf ( n4773 , n4772 );
buf ( n4774 , n4749 );
xor ( n4775 , n4771 , n4773 );
xor ( n4776 , n4775 , n4774 );
buf ( n4777 , n4776 );
xor ( n4778 , n4771 , n4773 );
and ( n4779 , n4778 , n4774 );
and ( n4780 , n4771 , n4773 );
or ( n4781 , n4779 , n4780 );
buf ( n4782 , n4781 );
buf ( n4783 , n4666 );
not ( n4784 , n4593 );
nand ( n4785 , n4784 , n4598 );
not ( n4786 , n4785 );
not ( n4787 , n4584 );
or ( n4788 , n4786 , n4787 );
nand ( n4789 , n4593 , n4597 );
buf ( n4790 , n4789 );
nand ( n4791 , n4788 , n4790 );
and ( n4792 , n387 , n388 );
xor ( n4793 , n387 , n4792 );
and ( n4794 , n386 , n389 );
xor ( n4795 , n4793 , n4794 );
not ( n4796 , n4795 );
xor ( n4797 , n4586 , n4587 );
and ( n4798 , n4797 , n4592 );
and ( n4799 , n4586 , n4587 );
or ( n4800 , n4798 , n4799 );
not ( n4801 , n4800 );
or ( n4802 , n4796 , n4801 );
or ( n4803 , n4795 , n4800 );
nand ( n4804 , n4802 , n4803 );
not ( n4805 , n4804 );
and ( n4806 , n4791 , n4805 );
not ( n4807 , n4791 );
buf ( n4808 , n4804 );
and ( n4809 , n4807 , n4808 );
nor ( n4810 , n4806 , n4809 );
buf ( n4811 , n4810 );
buf ( n4812 , n4811 );
buf ( n4813 , n4812 );
buf ( n4814 , n4813 );
buf ( n4815 , n393 );
nand ( n4816 , n4814 , n4815 );
buf ( n4817 , n4816 );
buf ( n4818 , n4817 );
not ( n4819 , n4818 );
buf ( n4820 , n4819 );
buf ( n4821 , n4820 );
buf ( n4822 , n4607 );
not ( n4823 , n4822 );
buf ( n4824 , n3533 );
nor ( n4825 , n4823 , n4824 );
buf ( n4826 , n4825 );
buf ( n4827 , n4826 );
xor ( n4828 , n4783 , n4821 );
xor ( n4829 , n4828 , n4827 );
buf ( n4830 , n4829 );
xor ( n4831 , n4783 , n4821 );
and ( n4832 , n4831 , n4827 );
and ( n4833 , n4783 , n4821 );
or ( n4834 , n4832 , n4833 );
buf ( n4835 , n4834 );
buf ( n4836 , n4765 );
buf ( n4837 , n4671 );
buf ( n4838 , n4676 );
xor ( n4839 , n4836 , n4837 );
xor ( n4840 , n4839 , n4838 );
buf ( n4841 , n4840 );
xor ( n4842 , n4836 , n4837 );
and ( n4843 , n4842 , n4838 );
and ( n4844 , n4836 , n4837 );
or ( n4845 , n4843 , n4844 );
buf ( n4846 , n4845 );
buf ( n4847 , n4777 );
buf ( n4848 , n4830 );
buf ( n4849 , n4681 );
xor ( n4850 , n4847 , n4848 );
xor ( n4851 , n4850 , n4849 );
buf ( n4852 , n4851 );
xor ( n4853 , n4847 , n4848 );
and ( n4854 , n4853 , n4849 );
and ( n4855 , n4847 , n4848 );
or ( n4856 , n4854 , n4855 );
buf ( n4857 , n4856 );
buf ( n4858 , n4841 );
buf ( n4859 , n4686 );
buf ( n4860 , n4852 );
xor ( n4861 , n4858 , n4859 );
xor ( n4862 , n4861 , n4860 );
buf ( n4863 , n4862 );
xor ( n4864 , n4858 , n4859 );
and ( n4865 , n4864 , n4860 );
and ( n4866 , n4858 , n4859 );
or ( n4867 , n4865 , n4866 );
buf ( n4868 , n4867 );
buf ( n4869 , n402 );
buf ( n4870 , n411 );
and ( n4871 , n4869 , n4870 );
buf ( n4872 , n4871 );
buf ( n4873 , n4872 );
buf ( n4874 , n403 );
buf ( n4875 , n410 );
and ( n4876 , n4874 , n4875 );
buf ( n4877 , n4876 );
buf ( n4878 , n4877 );
buf ( n4879 , n4709 );
xor ( n4880 , n4873 , n4878 );
xor ( n4881 , n4880 , n4879 );
buf ( n4882 , n4881 );
xor ( n4883 , n4873 , n4878 );
and ( n4884 , n4883 , n4879 );
and ( n4885 , n4873 , n4878 );
or ( n4886 , n4884 , n4885 );
buf ( n4887 , n4886 );
buf ( n4888 , n4882 );
buf ( n4889 , n3565 );
buf ( n4890 , n386 );
and ( n4891 , n4889 , n4890 );
buf ( n4892 , n4891 );
buf ( n4893 , n4892 );
buf ( n4894 , n4720 );
xor ( n4895 , n4888 , n4893 );
xor ( n4896 , n4895 , n4894 );
buf ( n4897 , n4896 );
xor ( n4898 , n4888 , n4893 );
and ( n4899 , n4898 , n4894 );
and ( n4900 , n4888 , n4893 );
or ( n4901 , n4899 , n4900 );
buf ( n4902 , n4901 );
buf ( n4903 , n3689 );
buf ( n4904 , n387 );
and ( n4905 , n4903 , n4904 );
buf ( n4906 , n4905 );
buf ( n4907 , n4906 );
and ( n4908 , n3963 , n388 );
buf ( n4909 , n4908 );
buf ( n4910 , n4739 );
xor ( n4911 , n4907 , n4909 );
xor ( n4912 , n4911 , n4910 );
buf ( n4913 , n4912 );
xor ( n4914 , n4907 , n4909 );
and ( n4915 , n4914 , n4910 );
and ( n4916 , n4907 , n4909 );
or ( n4917 , n4915 , n4916 );
buf ( n4918 , n4917 );
buf ( n4919 , n4178 );
buf ( n4920 , n389 );
and ( n4921 , n4919 , n4920 );
buf ( n4922 , n4921 );
buf ( n4923 , n4922 );
buf ( n4924 , n4897 );
and ( n4925 , n4394 , n4412 );
not ( n4926 , n4394 );
and ( n4927 , n4926 , n4415 );
nor ( n4928 , n4925 , n4927 );
buf ( n4929 , n4928 );
buf ( n4930 , n390 );
and ( n4931 , n4929 , n4930 );
buf ( n4932 , n4931 );
buf ( n4933 , n4932 );
xor ( n4934 , n4923 , n4924 );
xor ( n4935 , n4934 , n4933 );
buf ( n4936 , n4935 );
xor ( n4937 , n4923 , n4924 );
and ( n4938 , n4937 , n4933 );
and ( n4939 , n4923 , n4924 );
or ( n4940 , n4938 , n4939 );
buf ( n4941 , n4940 );
buf ( n4942 , n4810 );
buf ( n4943 , n392 );
and ( n4944 , n4942 , n4943 );
buf ( n4945 , n4944 );
buf ( n4946 , n4945 );
buf ( n4947 , n4607 );
buf ( n4948 , n391 );
and ( n4949 , n4947 , n4948 );
buf ( n4950 , n4949 );
buf ( n4951 , n4950 );
buf ( n4952 , n4754 );
xor ( n4953 , n4946 , n4951 );
xor ( n4954 , n4953 , n4952 );
buf ( n4955 , n4954 );
xor ( n4956 , n4946 , n4951 );
and ( n4957 , n4956 , n4952 );
and ( n4958 , n4946 , n4951 );
or ( n4959 , n4957 , n4958 );
buf ( n4960 , n4959 );
buf ( n4961 , n4913 );
buf ( n4962 , n4770 );
not ( n4963 , n4803 );
not ( n4964 , n4785 );
not ( n4965 , n4584 );
or ( n4966 , n4964 , n4965 );
nand ( n4967 , n4966 , n4789 );
not ( n4968 , n4967 );
or ( n4969 , n4963 , n4968 );
nand ( n4970 , n4800 , n4795 );
nand ( n4971 , n4969 , n4970 );
xor ( n4972 , n387 , n4792 );
and ( n4973 , n4972 , n4794 );
and ( n4974 , n387 , n4792 );
or ( n4975 , n4973 , n4974 );
and ( n4976 , n386 , n388 );
nor ( n4977 , n4975 , n4976 );
not ( n4978 , n4977 );
nand ( n4979 , n4975 , n4976 );
nand ( n4980 , n4978 , n4979 );
not ( n4981 , n4980 );
and ( n4982 , n4971 , n4981 );
not ( n4983 , n4971 );
and ( n4984 , n4983 , n4980 );
nor ( n4985 , n4982 , n4984 );
buf ( n4986 , n4985 );
buf ( n4987 , n393 );
and ( n4988 , n4986 , n4987 );
buf ( n4989 , n4988 );
buf ( n4990 , n4989 );
xor ( n4991 , n4961 , n4962 );
xor ( n4992 , n4991 , n4990 );
buf ( n4993 , n4992 );
xor ( n4994 , n4961 , n4962 );
and ( n4995 , n4994 , n4990 );
and ( n4996 , n4961 , n4962 );
or ( n4997 , n4995 , n4996 );
buf ( n4998 , n4997 );
buf ( n4999 , n4936 );
buf ( n5000 , n4835 );
buf ( n5001 , n4782 );
xor ( n5002 , n4999 , n5000 );
xor ( n5003 , n5002 , n5001 );
buf ( n5004 , n5003 );
xor ( n5005 , n4999 , n5000 );
and ( n5006 , n5005 , n5001 );
and ( n5007 , n4999 , n5000 );
or ( n5008 , n5006 , n5007 );
buf ( n5009 , n5008 );
buf ( n5010 , n4955 );
buf ( n5011 , n4993 );
buf ( n5012 , n4846 );
xor ( n5013 , n5010 , n5011 );
xor ( n5014 , n5013 , n5012 );
buf ( n5015 , n5014 );
xor ( n5016 , n5010 , n5011 );
and ( n5017 , n5016 , n5012 );
and ( n5018 , n5010 , n5011 );
or ( n5019 , n5017 , n5018 );
buf ( n5020 , n5019 );
buf ( n5021 , n5004 );
buf ( n5022 , n4857 );
buf ( n5023 , n5015 );
xor ( n5024 , n5021 , n5022 );
xor ( n5025 , n5024 , n5023 );
buf ( n5026 , n5025 );
xor ( n5027 , n5021 , n5022 );
and ( n5028 , n5027 , n5023 );
and ( n5029 , n5021 , n5022 );
or ( n5030 , n5028 , n5029 );
buf ( n5031 , n5030 );
buf ( n5032 , n402 );
buf ( n5033 , n410 );
and ( n5034 , n5032 , n5033 );
buf ( n5035 , n5034 );
buf ( n5036 , n5035 );
buf ( n5037 , n4887 );
buf ( n5038 , n386 );
not ( n5039 , n5038 );
buf ( n5040 , n4341 );
nor ( n5041 , n5039 , n5040 );
buf ( n5042 , n5041 );
buf ( n5043 , n5042 );
xor ( n5044 , n5036 , n5037 );
xor ( n5045 , n5044 , n5043 );
buf ( n5046 , n5045 );
xor ( n5047 , n5036 , n5037 );
and ( n5048 , n5047 , n5043 );
and ( n5049 , n5036 , n5037 );
or ( n5050 , n5048 , n5049 );
buf ( n5051 , n5050 );
buf ( n5052 , n3962 );
not ( n5053 , n5052 );
buf ( n5054 , n4326 );
nor ( n5055 , n5053 , n5054 );
buf ( n5056 , n5055 );
buf ( n5057 , n5056 );
buf ( n5058 , n4178 );
buf ( n5059 , n388 );
and ( n5060 , n5058 , n5059 );
buf ( n5061 , n5060 );
buf ( n5062 , n5061 );
buf ( n5063 , n4902 );
xor ( n5064 , n5057 , n5062 );
xor ( n5065 , n5064 , n5063 );
buf ( n5066 , n5065 );
xor ( n5067 , n5057 , n5062 );
and ( n5068 , n5067 , n5063 );
and ( n5069 , n5057 , n5062 );
or ( n5070 , n5068 , n5069 );
buf ( n5071 , n5070 );
buf ( n5072 , n5046 );
buf ( n5073 , n4417 );
buf ( n5074 , n389 );
and ( n5075 , n5073 , n5074 );
buf ( n5076 , n5075 );
buf ( n5077 , n5076 );
and ( n5078 , n4585 , n4603 );
not ( n5079 , n4585 );
and ( n5080 , n5079 , n4602 );
nor ( n5081 , n5078 , n5080 );
buf ( n5082 , n5081 );
buf ( n5083 , n390 );
and ( n5084 , n5082 , n5083 );
buf ( n5085 , n5084 );
buf ( n5086 , n5085 );
xor ( n5087 , n5072 , n5077 );
xor ( n5088 , n5087 , n5086 );
buf ( n5089 , n5088 );
xor ( n5090 , n5072 , n5077 );
and ( n5091 , n5090 , n5086 );
and ( n5092 , n5072 , n5077 );
or ( n5093 , n5091 , n5092 );
buf ( n5094 , n5093 );
buf ( n5095 , n4810 );
buf ( n5096 , n391 );
and ( n5097 , n5095 , n5096 );
buf ( n5098 , n5097 );
buf ( n5099 , n5098 );
not ( n5100 , n393 );
and ( n5101 , n4326 , n386 );
nor ( n5102 , n5100 , n5101 );
not ( n5103 , n5102 );
not ( n5104 , n4795 );
not ( n5105 , n4800 );
and ( n5106 , n5104 , n5105 );
nor ( n5107 , n5106 , n4977 );
not ( n5108 , n5107 );
not ( n5109 , n4967 );
or ( n5110 , n5108 , n5109 );
not ( n5111 , n4970 );
not ( n5112 , n4977 );
and ( n5113 , n5111 , n5112 );
not ( n5114 , n4979 );
nor ( n5115 , n5113 , n5114 );
nand ( n5116 , n5110 , n5115 );
not ( n5117 , n5116 );
or ( n5118 , n5103 , n5117 );
nand ( n5119 , n4967 , n5107 );
and ( n5120 , n5101 , n393 );
nand ( n5121 , n5119 , n5115 , n5120 );
nand ( n5122 , n5118 , n5121 );
buf ( n5123 , n5122 );
buf ( n5124 , n4918 );
xor ( n5125 , n5099 , n5123 );
xor ( n5126 , n5125 , n5124 );
buf ( n5127 , n5126 );
xor ( n5128 , n5099 , n5123 );
and ( n5129 , n5128 , n5124 );
and ( n5130 , n5099 , n5123 );
or ( n5131 , n5129 , n5130 );
buf ( n5132 , n5131 );
buf ( n5133 , n4941 );
and ( n5134 , n4985 , n392 );
buf ( n5135 , n5134 );
buf ( n5136 , n5066 );
xor ( n5137 , n5133 , n5135 );
xor ( n5138 , n5137 , n5136 );
buf ( n5139 , n5138 );
xor ( n5140 , n5133 , n5135 );
and ( n5141 , n5140 , n5136 );
and ( n5142 , n5133 , n5135 );
or ( n5143 , n5141 , n5142 );
buf ( n5144 , n5143 );
buf ( n5145 , n4960 );
buf ( n5146 , n5089 );
buf ( n5147 , n4998 );
xor ( n5148 , n5145 , n5146 );
xor ( n5149 , n5148 , n5147 );
buf ( n5150 , n5149 );
xor ( n5151 , n5145 , n5146 );
and ( n5152 , n5151 , n5147 );
and ( n5153 , n5145 , n5146 );
or ( n5154 , n5152 , n5153 );
buf ( n5155 , n5154 );
buf ( n5156 , n5127 );
buf ( n5157 , n5139 );
buf ( n5158 , n5009 );
xor ( n5159 , n5156 , n5157 );
xor ( n5160 , n5159 , n5158 );
buf ( n5161 , n5160 );
xor ( n5162 , n5156 , n5157 );
and ( n5163 , n5162 , n5158 );
and ( n5164 , n5156 , n5157 );
or ( n5165 , n5163 , n5164 );
buf ( n5166 , n5165 );
buf ( n5167 , n5150 );
buf ( n5168 , n5020 );
buf ( n5169 , n5161 );
xor ( n5170 , n5167 , n5168 );
xor ( n5171 , n5170 , n5169 );
buf ( n5172 , n5171 );
xor ( n5173 , n5167 , n5168 );
and ( n5174 , n5173 , n5169 );
and ( n5175 , n5167 , n5168 );
or ( n5176 , n5174 , n5175 );
buf ( n5177 , n5176 );
and ( n5178 , n386 , n3963 );
buf ( n5179 , n5178 );
buf ( n5180 , n4181 );
buf ( n5181 , n387 );
and ( n5182 , n5180 , n5181 );
buf ( n5183 , n5182 );
buf ( n5184 , n5183 );
buf ( n5185 , n4928 );
buf ( n5186 , n388 );
and ( n5187 , n5185 , n5186 );
buf ( n5188 , n5187 );
buf ( n5189 , n5188 );
xor ( n5190 , n5179 , n5184 );
xor ( n5191 , n5190 , n5189 );
buf ( n5192 , n5191 );
xor ( n5193 , n5179 , n5184 );
and ( n5194 , n5193 , n5189 );
and ( n5195 , n5179 , n5184 );
or ( n5196 , n5194 , n5195 );
buf ( n5197 , n5196 );
buf ( n5198 , n5051 );
buf ( n5199 , n4813 );
buf ( n5200 , n390 );
nand ( n5201 , n5199 , n5200 );
buf ( n5202 , n5201 );
buf ( n5203 , n5202 );
not ( n5204 , n5203 );
buf ( n5205 , n5204 );
buf ( n5206 , n5205 );
buf ( n5207 , n4607 );
buf ( n5208 , n389 );
and ( n5209 , n5207 , n5208 );
buf ( n5210 , n5209 );
buf ( n5211 , n5210 );
xor ( n5212 , n5198 , n5206 );
xor ( n5213 , n5212 , n5211 );
buf ( n5214 , n5213 );
xor ( n5215 , n5198 , n5206 );
and ( n5216 , n5215 , n5211 );
and ( n5217 , n5198 , n5206 );
or ( n5218 , n5216 , n5217 );
buf ( n5219 , n5218 );
and ( n5220 , n5107 , n386 );
not ( n5221 , n5220 );
not ( n5222 , n4791 );
or ( n5223 , n5221 , n5222 );
not ( n5224 , n4326 );
not ( n5225 , n5115 );
or ( n5226 , n5224 , n5225 );
nand ( n5227 , n5226 , n386 );
nand ( n5228 , n5223 , n5227 );
buf ( n5229 , n5228 );
buf ( n5230 , n393 );
and ( n5231 , n5229 , n5230 );
buf ( n5232 , n5231 );
buf ( n5233 , n5232 );
buf ( n5234 , n5071 );
xnor ( n5235 , n5116 , n5101 );
nor ( n5236 , n5235 , n3533 );
buf ( n5237 , n5236 );
xor ( n5238 , n5233 , n5234 );
xor ( n5239 , n5238 , n5237 );
buf ( n5240 , n5239 );
xor ( n5241 , n5233 , n5234 );
and ( n5242 , n5241 , n5237 );
and ( n5243 , n5233 , n5234 );
or ( n5244 , n5242 , n5243 );
buf ( n5245 , n5244 );
buf ( n5246 , n5192 );
buf ( n5247 , n4985 );
buf ( n5248 , n391 );
and ( n5249 , n5247 , n5248 );
buf ( n5250 , n5249 );
buf ( n5251 , n5250 );
buf ( n5252 , n5094 );
xor ( n5253 , n5246 , n5251 );
xor ( n5254 , n5253 , n5252 );
buf ( n5255 , n5254 );
xor ( n5256 , n5246 , n5251 );
and ( n5257 , n5256 , n5252 );
and ( n5258 , n5246 , n5251 );
or ( n5259 , n5257 , n5258 );
buf ( n5260 , n5259 );
buf ( n5261 , n5132 );
buf ( n5262 , n5214 );
buf ( n5263 , n5240 );
xor ( n5264 , n5261 , n5262 );
xor ( n5265 , n5264 , n5263 );
buf ( n5266 , n5265 );
xor ( n5267 , n5261 , n5262 );
and ( n5268 , n5267 , n5263 );
and ( n5269 , n5261 , n5262 );
or ( n5270 , n5268 , n5269 );
buf ( n5271 , n5270 );
buf ( n5272 , n5144 );
buf ( n5273 , n5255 );
buf ( n5274 , n5155 );
xor ( n5275 , n5272 , n5273 );
xor ( n5276 , n5275 , n5274 );
buf ( n5277 , n5276 );
xor ( n5278 , n5272 , n5273 );
and ( n5279 , n5278 , n5274 );
and ( n5280 , n5272 , n5273 );
or ( n5281 , n5279 , n5280 );
buf ( n5282 , n5281 );
buf ( n5283 , n5266 );
buf ( n5284 , n5166 );
buf ( n5285 , n5277 );
xor ( n5286 , n5283 , n5284 );
xor ( n5287 , n5286 , n5285 );
buf ( n5288 , n5287 );
xor ( n5289 , n5283 , n5284 );
and ( n5290 , n5289 , n5285 );
and ( n5291 , n5283 , n5284 );
or ( n5292 , n5290 , n5291 );
buf ( n5293 , n5292 );
buf ( n5294 , n4181 );
buf ( n5295 , n386 );
and ( n5296 , n5294 , n5295 );
buf ( n5297 , n5296 );
buf ( n5298 , n5297 );
buf ( n5299 , n4928 );
buf ( n5300 , n387 );
and ( n5301 , n5299 , n5300 );
buf ( n5302 , n5301 );
buf ( n5303 , n5302 );
buf ( n5304 , n5228 );
buf ( n5305 , n392 );
and ( n5306 , n5304 , n5305 );
buf ( n5307 , n5306 );
buf ( n5308 , n5307 );
xor ( n5309 , n5298 , n5303 );
xor ( n5310 , n5309 , n5308 );
buf ( n5311 , n5310 );
xor ( n5312 , n5298 , n5303 );
and ( n5313 , n5312 , n5308 );
and ( n5314 , n5298 , n5303 );
or ( n5315 , n5313 , n5314 );
buf ( n5316 , n5315 );
buf ( n5317 , n4813 );
buf ( n5318 , n389 );
and ( n5319 , n5317 , n5318 );
buf ( n5320 , n5319 );
buf ( n5321 , n5320 );
buf ( n5322 , n5081 );
buf ( n5323 , n388 );
and ( n5324 , n5322 , n5323 );
buf ( n5325 , n5324 );
buf ( n5326 , n5325 );
not ( n5327 , n5101 );
not ( n5328 , n5116 );
not ( n5329 , n5328 );
or ( n5330 , n5327 , n5329 );
or ( n5331 , n5328 , n5101 );
nand ( n5332 , n5330 , n5331 );
buf ( n5333 , n5332 );
buf ( n5334 , n391 );
and ( n5335 , n5333 , n5334 );
buf ( n5336 , n5335 );
buf ( n5337 , n5336 );
xor ( n5338 , n5321 , n5326 );
xor ( n5339 , n5338 , n5337 );
buf ( n5340 , n5339 );
xor ( n5341 , n5321 , n5326 );
and ( n5342 , n5341 , n5337 );
and ( n5343 , n5321 , n5326 );
or ( n5344 , n5342 , n5343 );
buf ( n5345 , n5344 );
and ( n5346 , n4985 , n390 );
buf ( n5347 , n5346 );
buf ( n5348 , n5197 );
buf ( n5349 , n5219 );
xor ( n5350 , n5347 , n5348 );
xor ( n5351 , n5350 , n5349 );
buf ( n5352 , n5351 );
xor ( n5353 , n5347 , n5348 );
and ( n5354 , n5353 , n5349 );
and ( n5355 , n5347 , n5348 );
or ( n5356 , n5354 , n5355 );
buf ( n5357 , n5356 );
buf ( n5358 , n5311 );
buf ( n5359 , n5245 );
buf ( n5360 , n5340 );
xor ( n5361 , n5358 , n5359 );
xor ( n5362 , n5361 , n5360 );
buf ( n5363 , n5362 );
xor ( n5364 , n5358 , n5359 );
and ( n5365 , n5364 , n5360 );
and ( n5366 , n5358 , n5359 );
or ( n5367 , n5365 , n5366 );
buf ( n5368 , n5367 );
buf ( n5369 , n5352 );
buf ( n5370 , n5260 );
buf ( n5371 , n5271 );
xor ( n5372 , n5369 , n5370 );
xor ( n5373 , n5372 , n5371 );
buf ( n5374 , n5373 );
xor ( n5375 , n5369 , n5370 );
and ( n5376 , n5375 , n5371 );
and ( n5377 , n5369 , n5370 );
or ( n5378 , n5376 , n5377 );
buf ( n5379 , n5378 );
buf ( n5380 , n5363 );
buf ( n5381 , n5374 );
buf ( n5382 , n5282 );
xor ( n5383 , n5380 , n5381 );
xor ( n5384 , n5383 , n5382 );
buf ( n5385 , n5384 );
xor ( n5386 , n5380 , n5381 );
and ( n5387 , n5386 , n5382 );
and ( n5388 , n5380 , n5381 );
or ( n5389 , n5387 , n5388 );
buf ( n5390 , n5389 );
buf ( n5391 , n4417 );
buf ( n5392 , n386 );
and ( n5393 , n5391 , n5392 );
buf ( n5394 , n5393 );
buf ( n5395 , n5394 );
buf ( n5396 , n4813 );
buf ( n5397 , n5396 );
buf ( n5398 , n5397 );
buf ( n5399 , n5398 );
buf ( n5400 , n388 );
nand ( n5401 , n5399 , n5400 );
buf ( n5402 , n5401 );
buf ( n5403 , n5402 );
not ( n5404 , n5403 );
buf ( n5405 , n5404 );
buf ( n5406 , n5405 );
buf ( n5407 , n5081 );
not ( n5408 , n5407 );
buf ( n5409 , n4326 );
nor ( n5410 , n5408 , n5409 );
buf ( n5411 , n5410 );
buf ( n5412 , n5411 );
xor ( n5413 , n5395 , n5406 );
xor ( n5414 , n5413 , n5412 );
buf ( n5415 , n5414 );
xor ( n5416 , n5395 , n5406 );
and ( n5417 , n5416 , n5412 );
and ( n5418 , n5395 , n5406 );
or ( n5419 , n5417 , n5418 );
buf ( n5420 , n5419 );
buf ( n5421 , n5228 );
buf ( n5422 , n5421 );
buf ( n5423 , n5422 );
buf ( n5424 , n5423 );
buf ( n5425 , n391 );
and ( n5426 , n5424 , n5425 );
buf ( n5427 , n5426 );
buf ( n5428 , n5427 );
and ( n5429 , n5332 , n390 );
buf ( n5430 , n5429 );
buf ( n5431 , n4985 );
buf ( n5432 , n389 );
and ( n5433 , n5431 , n5432 );
buf ( n5434 , n5433 );
buf ( n5435 , n5434 );
xor ( n5436 , n5428 , n5430 );
xor ( n5437 , n5436 , n5435 );
buf ( n5438 , n5437 );
xor ( n5439 , n5428 , n5430 );
and ( n5440 , n5439 , n5435 );
and ( n5441 , n5428 , n5430 );
or ( n5442 , n5440 , n5441 );
buf ( n5443 , n5442 );
buf ( n5444 , n5316 );
buf ( n5445 , n5345 );
buf ( n5446 , n5415 );
xor ( n5447 , n5444 , n5445 );
xor ( n5448 , n5447 , n5446 );
buf ( n5449 , n5448 );
xor ( n5450 , n5444 , n5445 );
and ( n5451 , n5450 , n5446 );
and ( n5452 , n5444 , n5445 );
or ( n5453 , n5451 , n5452 );
buf ( n5454 , n5453 );
buf ( n5455 , n5438 );
buf ( n5456 , n5357 );
buf ( n5457 , n5368 );
xor ( n5458 , n5455 , n5456 );
xor ( n5459 , n5458 , n5457 );
buf ( n5460 , n5459 );
xor ( n5461 , n5455 , n5456 );
and ( n5462 , n5461 , n5457 );
and ( n5463 , n5455 , n5456 );
or ( n5464 , n5462 , n5463 );
buf ( n5465 , n5464 );
buf ( n5466 , n5449 );
buf ( n5467 , n5460 );
buf ( n5468 , n5379 );
xor ( n5469 , n5466 , n5467 );
xor ( n5470 , n5469 , n5468 );
buf ( n5471 , n5470 );
xor ( n5472 , n5466 , n5467 );
and ( n5473 , n5472 , n5468 );
and ( n5474 , n5466 , n5467 );
or ( n5475 , n5473 , n5474 );
buf ( n5476 , n5475 );
buf ( n5477 , n5423 );
buf ( n5478 , n390 );
and ( n5479 , n5477 , n5478 );
buf ( n5480 , n5479 );
buf ( n5481 , n5480 );
buf ( n5482 , n5081 );
buf ( n5483 , n386 );
and ( n5484 , n5482 , n5483 );
buf ( n5485 , n5484 );
buf ( n5486 , n5485 );
buf ( n5487 , n5398 );
buf ( n5488 , n387 );
and ( n5489 , n5487 , n5488 );
buf ( n5490 , n5489 );
buf ( n5491 , n5490 );
xor ( n5492 , n5481 , n5486 );
xor ( n5493 , n5492 , n5491 );
buf ( n5494 , n5493 );
xor ( n5495 , n5481 , n5486 );
and ( n5496 , n5495 , n5491 );
and ( n5497 , n5481 , n5486 );
or ( n5498 , n5496 , n5497 );
buf ( n5499 , n5498 );
buf ( n5500 , n5332 );
buf ( n5501 , n389 );
and ( n5502 , n5500 , n5501 );
buf ( n5503 , n5502 );
buf ( n5504 , n5503 );
and ( n5505 , n4985 , n388 );
buf ( n5506 , n5505 );
buf ( n5507 , n5420 );
xor ( n5508 , n5504 , n5506 );
xor ( n5509 , n5508 , n5507 );
buf ( n5510 , n5509 );
xor ( n5511 , n5504 , n5506 );
and ( n5512 , n5511 , n5507 );
and ( n5513 , n5504 , n5506 );
or ( n5514 , n5512 , n5513 );
buf ( n5515 , n5514 );
buf ( n5516 , n5494 );
buf ( n5517 , n5443 );
buf ( n5518 , n5510 );
xor ( n5519 , n5516 , n5517 );
xor ( n5520 , n5519 , n5518 );
buf ( n5521 , n5520 );
xor ( n5522 , n5516 , n5517 );
and ( n5523 , n5522 , n5518 );
and ( n5524 , n5516 , n5517 );
or ( n5525 , n5523 , n5524 );
buf ( n5526 , n5525 );
buf ( n5527 , n5454 );
buf ( n5528 , n5521 );
buf ( n5529 , n5465 );
xor ( n5530 , n5527 , n5528 );
xor ( n5531 , n5530 , n5529 );
buf ( n5532 , n5531 );
xor ( n5533 , n5527 , n5528 );
and ( n5534 , n5533 , n5529 );
and ( n5535 , n5527 , n5528 );
or ( n5536 , n5534 , n5535 );
buf ( n5537 , n5536 );
buf ( n5538 , n5423 );
buf ( n5539 , n389 );
and ( n5540 , n5538 , n5539 );
buf ( n5541 , n5540 );
buf ( n5542 , n5541 );
buf ( n5543 , n5398 );
buf ( n5544 , n386 );
and ( n5545 , n5543 , n5544 );
buf ( n5546 , n5545 );
buf ( n5547 , n5546 );
buf ( n5548 , n5332 );
buf ( n5549 , n388 );
and ( n5550 , n5548 , n5549 );
buf ( n5551 , n5550 );
buf ( n5552 , n5551 );
xor ( n5553 , n5542 , n5547 );
xor ( n5554 , n5553 , n5552 );
buf ( n5555 , n5554 );
xor ( n5556 , n5542 , n5547 );
and ( n5557 , n5556 , n5552 );
and ( n5558 , n5542 , n5547 );
or ( n5559 , n5557 , n5558 );
buf ( n5560 , n5559 );
buf ( n5561 , n4985 );
buf ( n5562 , n387 );
and ( n5563 , n5561 , n5562 );
buf ( n5564 , n5563 );
buf ( n5565 , n5564 );
buf ( n5566 , n5499 );
buf ( n5567 , n5555 );
xor ( n5568 , n5565 , n5566 );
xor ( n5569 , n5568 , n5567 );
buf ( n5570 , n5569 );
xor ( n5571 , n5565 , n5566 );
and ( n5572 , n5571 , n5567 );
and ( n5573 , n5565 , n5566 );
or ( n5574 , n5572 , n5573 );
buf ( n5575 , n5574 );
buf ( n5576 , n5515 );
buf ( n5577 , n5570 );
buf ( n5578 , n5526 );
xor ( n5579 , n5576 , n5577 );
xor ( n5580 , n5579 , n5578 );
buf ( n5581 , n5580 );
xor ( n5582 , n5576 , n5577 );
and ( n5583 , n5582 , n5578 );
and ( n5584 , n5576 , n5577 );
or ( n5585 , n5583 , n5584 );
buf ( n5586 , n5585 );
buf ( n5587 , n5423 );
buf ( n5588 , n388 );
and ( n5589 , n5587 , n5588 );
buf ( n5590 , n5589 );
buf ( n5591 , n5590 );
buf ( n5592 , n5332 );
buf ( n5593 , n387 );
and ( n5594 , n5592 , n5593 );
buf ( n5595 , n5594 );
buf ( n5596 , n5595 );
buf ( n5597 , n4985 );
buf ( n5598 , n386 );
and ( n5599 , n5597 , n5598 );
buf ( n5600 , n5599 );
buf ( n5601 , n5600 );
xor ( n5602 , n5591 , n5596 );
xor ( n5603 , n5602 , n5601 );
buf ( n5604 , n5603 );
and ( n5605 , n5591 , n5596 );
or ( n5606 , C0 , n5605 );
buf ( n5607 , n5606 );
buf ( n5608 , n5560 );
buf ( n5609 , n5604 );
buf ( n5610 , n5575 );
xor ( n5611 , n5608 , n5609 );
xor ( n5612 , n5611 , n5610 );
buf ( n5613 , n5612 );
xor ( n5614 , n5608 , n5609 );
and ( n5615 , n5614 , n5610 );
and ( n5616 , n5608 , n5609 );
or ( n5617 , n5615 , n5616 );
buf ( n5618 , n5617 );
buf ( n5619 , n5423 );
buf ( n5620 , n387 );
and ( n5621 , n5619 , n5620 );
buf ( n5622 , n5621 );
buf ( n5623 , n5622 );
buf ( n5624 , n5332 );
buf ( n5625 , n386 );
and ( n5626 , n5624 , n5625 );
buf ( n5627 , n5626 );
buf ( n5628 , n5627 );
buf ( n5629 , n5607 );
xor ( n5630 , n5623 , n5628 );
xor ( n5631 , n5630 , n5629 );
buf ( n5632 , n5631 );
and ( n5633 , n5623 , n5628 );
or ( n5634 , C0 , n5633 );
buf ( n5635 , n5634 );
not ( n5636 , n5390 );
not ( n5637 , n5636 );
not ( n5638 , n5471 );
not ( n5639 , n5638 );
or ( n5640 , n5637 , n5639 );
not ( n5641 , n5471 );
not ( n5642 , n5390 );
or ( n5643 , n5641 , n5642 );
nand ( n5644 , n5385 , n5293 );
nand ( n5645 , n5643 , n5644 );
nand ( n5646 , n5640 , n5645 );
not ( n5647 , n5646 );
not ( n5648 , n5476 );
not ( n5649 , n5532 );
nand ( n5650 , n5648 , n5649 );
not ( n5651 , n5537 );
not ( n5652 , n5581 );
nand ( n5653 , n5651 , n5652 );
and ( n5654 , n5650 , n5653 );
and ( n5655 , n5647 , n5654 );
not ( n5656 , n5537 );
nand ( n5657 , n5656 , n5652 );
not ( n5658 , n5657 );
nand ( n5659 , n5532 , n5476 );
not ( n5660 , n5659 );
not ( n5661 , n5660 );
or ( n5662 , n5658 , n5661 );
not ( n5663 , n5652 );
nand ( n5664 , n5663 , n5537 );
nand ( n5665 , n5662 , n5664 );
nor ( n5666 , n5655 , n5665 );
buf ( n5667 , n5666 );
not ( n5668 , n5667 );
buf ( n5669 , n5668 );
not ( n5670 , n5636 );
not ( n5671 , n5638 );
or ( n5672 , n5670 , n5671 );
buf ( n5673 , n5385 );
not ( n5674 , n5673 );
buf ( n5675 , n5674 );
buf ( n5676 , n5293 );
not ( n5677 , n5676 );
buf ( n5678 , n5677 );
nand ( n5679 , n5675 , n5678 );
nand ( n5680 , n5672 , n5679 );
not ( n5681 , n5680 );
buf ( n5682 , n5681 );
buf ( n5683 , n5654 );
or ( n5684 , n5613 , n5586 );
buf ( n5685 , n5618 );
buf ( n5686 , n5632 );
or ( n5687 , n5685 , n5686 );
buf ( n5688 , n5687 );
nand ( n5689 , n5684 , n5688 );
not ( n5690 , n5635 );
buf ( n5691 , n5423 );
buf ( n5692 , n386 );
nand ( n5693 , n5691 , n5692 );
buf ( n5694 , n5693 );
nand ( n5695 , n5690 , n5694 );
not ( n5696 , n5695 );
nor ( n5697 , n5689 , n5696 );
buf ( n5698 , n5697 );
and ( n5699 , n5682 , n5683 , n5698 );
buf ( n5700 , n5699 );
buf ( n5701 , n5675 );
not ( n5702 , n5701 );
buf ( n5703 , n5293 );
nand ( n5704 , n5702 , n5703 );
buf ( n5705 , n5704 );
buf ( n5706 , n5705 );
buf ( n5707 , n5679 );
and ( n5708 , n5706 , n5707 );
buf ( n5709 , n5708 );
buf ( n5710 , n5705 );
not ( n5711 , n5710 );
buf ( n5712 , n5711 );
nand ( n5713 , n5177 , n5288 );
buf ( n5714 , n5713 );
not ( n5715 , n5714 );
buf ( n5716 , n5715 );
buf ( n5717 , n5026 );
buf ( n5718 , n4868 );
nand ( n5719 , n5717 , n5718 );
buf ( n5720 , n5719 );
buf ( n5721 , n4863 );
not ( n5722 , n5721 );
buf ( n5723 , n5722 );
or ( n5724 , n4641 , n4438 );
buf ( n5725 , n5724 );
nand ( n5726 , n4641 , n4438 );
buf ( n5727 , n5726 );
buf ( n5728 , n5727 );
nand ( n5729 , n5725 , n5728 );
buf ( n5730 , n5729 );
not ( n5731 , n3422 );
not ( n5732 , n3596 );
or ( n5733 , n5731 , n5732 );
not ( n5734 , n3268 );
not ( n5735 , n3150 );
buf ( n5736 , n3078 );
buf ( n5737 , n3083 );
xnor ( n5738 , n5736 , n5737 );
buf ( n5739 , n5738 );
buf ( n5740 , n5739 );
buf ( n5741 , n393 );
buf ( n5742 , n409 );
nand ( n5743 , n5741 , n5742 );
buf ( n5744 , n5743 );
buf ( n5745 , n5744 );
not ( n5746 , n5745 );
buf ( n5747 , n408 );
nand ( n5748 , n5746 , n5747 );
buf ( n5749 , n5748 );
buf ( n5750 , n5749 );
nand ( n5751 , n5740 , n5750 );
buf ( n5752 , n5751 );
buf ( n5753 , n5752 );
buf ( n5754 , n408 );
not ( n5755 , n5754 );
buf ( n5756 , n5744 );
nand ( n5757 , n5755 , n5756 );
buf ( n5758 , n5757 );
buf ( n5759 , n5758 );
buf ( n5760 , n417 );
and ( n5761 , n5753 , n5759 , n5760 );
buf ( n5762 , n5761 );
buf ( n5763 , n5762 );
not ( n5764 , n5763 );
buf ( n5765 , n3091 );
not ( n5766 , n5765 );
or ( n5767 , n5764 , n5766 );
buf ( n5768 , n3064 );
not ( n5769 , n5768 );
buf ( n5770 , n5769 );
buf ( n5771 , n5770 );
nand ( n5772 , n5767 , n5771 );
buf ( n5773 , n5772 );
buf ( n5774 , n3091 );
buf ( n5775 , n5762 );
or ( n5776 , n5774 , n5775 );
buf ( n5777 , n5776 );
and ( n5778 , n3139 , n5773 , n5777 );
not ( n5779 , n5778 );
and ( n5780 , n5735 , n5779 );
buf ( n5781 , n5773 );
buf ( n5782 , n5777 );
and ( n5783 , n5781 , n5782 );
buf ( n5784 , n3139 );
nor ( n5785 , n5783 , n5784 );
buf ( n5786 , n5785 );
nor ( n5787 , n5780 , n5786 );
nand ( n5788 , n5787 , n3234 );
nand ( n5789 , n5734 , n5788 );
or ( n5790 , n5787 , n3234 );
and ( n5791 , n5789 , n5790 , n3273 );
or ( n5792 , n5791 , n3417 );
not ( n5793 , n3273 );
nand ( n5794 , n5789 , n5790 );
nand ( n5795 , n5793 , n5794 );
nand ( n5796 , n5792 , n5795 );
nand ( n5797 , n5733 , n5796 );
buf ( n5798 , n5797 );
buf ( n5799 , n3596 );
buf ( n5800 , n3422 );
or ( n5801 , n5799 , n5800 );
buf ( n5802 , n5801 );
buf ( n5803 , n5802 );
buf ( n5804 , n3601 );
and ( n5805 , n5798 , n5803 );
nor ( n5806 , n5805 , n5804 );
buf ( n5807 , n5806 );
buf ( n5808 , n5618 );
buf ( n5809 , n5632 );
nand ( n5810 , n5808 , n5809 );
buf ( n5811 , n5810 );
buf ( n5812 , n5811 );
not ( n5813 , n5812 );
buf ( n5814 , n5813 );
buf ( n5815 , n5635 );
not ( n5816 , n5815 );
buf ( n5817 , n5816 );
buf ( n5818 , n5817 );
buf ( n5819 , n5694 );
nor ( n5820 , n5818 , n5819 );
buf ( n5821 , n5820 );
nand ( n5822 , n5684 , n5650 , n5653 );
buf ( n5823 , n5822 );
buf ( n5824 , n5681 );
not ( n5825 , n5823 );
nand ( n5826 , n5825 , n5824 );
buf ( n5827 , n5826 );
buf ( n5828 , n5636 );
buf ( n5829 , n5638 );
or ( n5830 , n5828 , n5829 );
buf ( n5831 , n5830 );
xnor ( n5832 , n413 , n412 );
buf ( n5833 , n411 );
buf ( n5834 , n412 );
xor ( n5835 , n5833 , n5834 );
buf ( n5836 , n5835 );
and ( n5837 , n5832 , n5836 );
buf ( n5838 , n5837 );
not ( n5839 , n5838 );
buf ( n5840 , n5839 );
nand ( n5841 , n5840 , n5832 );
not ( n5842 , n411 );
and ( n5843 , n421 , n425 );
buf ( n5844 , n422 );
buf ( n5845 , n423 );
or ( n5846 , n5844 , n5845 );
buf ( n5847 , n373 );
not ( n5848 , n5847 );
buf ( n5849 , n5848 );
buf ( n5850 , n5849 );
nand ( n5851 , n5846 , n5850 );
buf ( n5852 , n5851 );
nand ( n5853 , n422 , n423 );
nand ( n5854 , n5852 , n5853 );
xor ( n5855 , n5843 , n5854 );
buf ( n5856 , n372 );
not ( n5857 , n5856 );
buf ( n5858 , n421 );
not ( n5859 , n5858 );
and ( n5860 , n5857 , n5859 );
buf ( n5861 , n372 );
buf ( n5862 , n421 );
and ( n5863 , n5861 , n5862 );
nor ( n5864 , n5860 , n5863 );
buf ( n5865 , n5864 );
nand ( n5866 , n424 , n422 );
and ( n5867 , n5865 , n5866 );
not ( n5868 , n5865 );
not ( n5869 , n5866 );
and ( n5870 , n5868 , n5869 );
nor ( n5871 , n5867 , n5870 );
xor ( n5872 , n5855 , n5871 );
buf ( n5873 , n422 );
buf ( n5874 , n425 );
nand ( n5875 , n5873 , n5874 );
buf ( n5876 , n5875 );
buf ( n5877 , n5876 );
not ( n5878 , n5877 );
buf ( n5879 , n424 );
buf ( n5880 , n423 );
nand ( n5881 , n5879 , n5880 );
buf ( n5882 , n5881 );
buf ( n5883 , n5882 );
not ( n5884 , n5883 );
or ( n5885 , n5878 , n5884 );
buf ( n5886 , n424 );
buf ( n5887 , n423 );
nor ( n5888 , n5886 , n5887 );
buf ( n5889 , n5888 );
buf ( n5890 , n5889 );
buf ( n5891 , n374 );
or ( n5892 , n5890 , n5891 );
buf ( n5893 , n5882 );
nand ( n5894 , n5892 , n5893 );
buf ( n5895 , n5894 );
buf ( n5896 , n5895 );
nand ( n5897 , n5885 , n5896 );
buf ( n5898 , n5897 );
buf ( n5899 , n5898 );
not ( n5900 , n5899 );
buf ( n5901 , n5900 );
nor ( n5902 , n5872 , n5901 );
buf ( n5903 , n5902 );
buf ( n5904 , n424 );
buf ( n5905 , n423 );
and ( n5906 , n5904 , n5905 );
buf ( n5907 , n5906 );
buf ( n5908 , n5907 );
buf ( n5909 , n5876 );
and ( n5910 , n5908 , n5909 );
not ( n5911 , n5908 );
buf ( n5912 , n5876 );
not ( n5913 , n5912 );
buf ( n5914 , n5913 );
buf ( n5915 , n5914 );
and ( n5916 , n5911 , n5915 );
nor ( n5917 , n5910 , n5916 );
buf ( n5918 , n5917 );
xnor ( n5919 , n5918 , n5895 );
buf ( n5920 , n5919 );
xor ( n5921 , n423 , n373 );
xnor ( n5922 , n5921 , n422 );
buf ( n5923 , n5922 );
nor ( n5924 , n5920 , n5923 );
buf ( n5925 , n5924 );
buf ( n5926 , n5925 );
nor ( n5927 , n5903 , n5926 );
buf ( n5928 , n5927 );
buf ( n5929 , n5928 );
xor ( n5930 , n5843 , n5854 );
and ( n5931 , n5930 , n5871 );
and ( n5932 , n5843 , n5854 );
or ( n5933 , n5931 , n5932 );
not ( n5934 , n5933 );
not ( n5935 , n421 );
nand ( n5936 , n5935 , n372 );
not ( n5937 , n5936 );
and ( n5938 , n422 , n424 );
not ( n5939 , n5938 );
or ( n5940 , n5937 , n5939 );
not ( n5941 , n372 );
nand ( n5942 , n5941 , n421 );
nand ( n5943 , n5940 , n5942 );
not ( n5944 , n5943 );
xor ( n5945 , n371 , n420 );
and ( n5946 , n5945 , n422 );
not ( n5947 , n5945 );
not ( n5948 , n422 );
and ( n5949 , n5947 , n5948 );
nor ( n5950 , n5946 , n5949 );
not ( n5951 , n5950 );
not ( n5952 , n5951 );
or ( n5953 , n5944 , n5952 );
or ( n5954 , n5943 , n5951 );
nand ( n5955 , n5953 , n5954 );
not ( n5956 , n5955 );
and ( n5957 , n422 , n423 );
buf ( n5958 , n420 );
buf ( n5959 , n425 );
and ( n5960 , n5958 , n5959 );
buf ( n5961 , n5960 );
nand ( n5962 , n424 , n421 );
and ( n5963 , n5961 , n5962 );
not ( n5964 , n5961 );
not ( n5965 , n5962 );
and ( n5966 , n5964 , n5965 );
or ( n5967 , n5963 , n5966 );
xor ( n5968 , n5957 , n5967 );
not ( n5969 , n5968 );
or ( n5970 , n5956 , n5969 );
or ( n5971 , n5955 , n5968 );
nand ( n5972 , n5970 , n5971 );
not ( n5973 , n5972 );
nand ( n5974 , n5934 , n5973 );
buf ( n5975 , n5974 );
not ( n5976 , n425 );
nand ( n5977 , n5976 , n419 );
and ( n5978 , n5977 , n370 );
not ( n5979 , n5977 );
not ( n5980 , n370 );
and ( n5981 , n5979 , n5980 );
nor ( n5982 , n5978 , n5981 );
buf ( n5983 , n5982 );
not ( n5984 , n5957 );
not ( n5985 , n5965 );
or ( n5986 , n5984 , n5985 );
not ( n5987 , n5853 );
not ( n5988 , n5962 );
or ( n5989 , n5987 , n5988 );
nand ( n5990 , n5989 , n5961 );
nand ( n5991 , n5986 , n5990 );
buf ( n5992 , n5991 );
xor ( n5993 , n5983 , n5992 );
buf ( n5994 , n424 );
buf ( n5995 , n420 );
nand ( n5996 , n5994 , n5995 );
buf ( n5997 , n5996 );
buf ( n5998 , n5997 );
not ( n5999 , n5998 );
buf ( n6000 , n5999 );
buf ( n6001 , n6000 );
buf ( n6002 , n421 );
buf ( n6003 , n423 );
and ( n6004 , n6002 , n6003 );
buf ( n6005 , n6004 );
buf ( n6006 , n6005 );
xor ( n6007 , n6001 , n6006 );
buf ( n6008 , n420 );
buf ( n6009 , n422 );
nor ( n6010 , n6008 , n6009 );
buf ( n6011 , n6010 );
buf ( n6012 , n6011 );
buf ( n6013 , n371 );
or ( n6014 , n6012 , n6013 );
buf ( n6015 , n420 );
buf ( n6016 , n422 );
nand ( n6017 , n6015 , n6016 );
buf ( n6018 , n6017 );
buf ( n6019 , n6018 );
nand ( n6020 , n6014 , n6019 );
buf ( n6021 , n6020 );
buf ( n6022 , n6021 );
xor ( n6023 , n6007 , n6022 );
buf ( n6024 , n6023 );
buf ( n6025 , n6024 );
xor ( n6026 , n5993 , n6025 );
buf ( n6027 , n6026 );
buf ( n6028 , n6027 );
not ( n6029 , n6028 );
buf ( n6030 , n5943 );
not ( n6031 , n6030 );
buf ( n6032 , n5950 );
buf ( n6033 , n6032 );
nand ( n6034 , n6031 , n6033 );
buf ( n6035 , n6034 );
and ( n6036 , n5968 , n6035 );
not ( n6037 , n5943 );
nor ( n6038 , n6037 , n6032 );
nor ( n6039 , n6036 , n6038 );
buf ( n6040 , n6039 );
nand ( n6041 , n6029 , n6040 );
buf ( n6042 , n6041 );
buf ( n6043 , n6042 );
xor ( n6044 , n424 , n374 );
not ( n6045 , n423 );
xor ( n6046 , n6044 , n6045 );
buf ( n6047 , n6046 );
buf ( n6048 , n423 );
buf ( n6049 , n425 );
and ( n6050 , n6048 , n6049 );
buf ( n6051 , n6050 );
buf ( n6052 , n6051 );
or ( n6053 , n6047 , n6052 );
not ( n6054 , n376 );
not ( n6055 , n377 );
and ( n6056 , n6054 , n6055 );
nor ( n6057 , n6056 , n425 );
buf ( n6058 , n6057 );
and ( n6059 , n424 , n425 );
nor ( n6060 , n6059 , n706 );
buf ( n6061 , n6060 );
nor ( n6062 , n6058 , n6061 );
buf ( n6063 , n6062 );
buf ( n6064 , n6063 );
nand ( n6065 , n6053 , n6064 );
buf ( n6066 , n6065 );
buf ( n6067 , n6046 );
buf ( n6068 , n6051 );
nand ( n6069 , n6067 , n6068 );
buf ( n6070 , n6069 );
nand ( n6071 , n6066 , n6070 );
buf ( n6072 , n6071 );
nand ( n6073 , n5929 , n5975 , n6043 , n6072 );
buf ( n6074 , n6073 );
buf ( n6075 , n5972 );
buf ( n6076 , n5933 );
nor ( n6077 , n6075 , n6076 );
buf ( n6078 , n6077 );
buf ( n6079 , n6078 );
buf ( n6080 , n5902 );
nor ( n6081 , n6079 , n6080 );
buf ( n6082 , n6081 );
buf ( n6083 , n6082 );
buf ( n6084 , n6042 );
nand ( n6085 , n5872 , n5901 );
buf ( n6086 , n6085 );
nand ( n6087 , n5919 , n5922 );
buf ( n6088 , n6087 );
nand ( n6089 , n6086 , n6088 );
buf ( n6090 , n6089 );
buf ( n6091 , n6090 );
nand ( n6092 , n6083 , n6084 , n6091 );
buf ( n6093 , n6092 );
buf ( n6094 , n6027 );
not ( n6095 , n6094 );
buf ( n6096 , n6039 );
nand ( n6097 , n6095 , n6096 );
buf ( n6098 , n6097 );
buf ( n6099 , n6098 );
buf ( n6100 , n5972 );
buf ( n6101 , n5933 );
and ( n6102 , n6100 , n6101 );
buf ( n6103 , n6102 );
buf ( n6104 , n6103 );
nand ( n6105 , n6099 , n6104 );
buf ( n6106 , n6105 );
buf ( n6107 , n6039 );
not ( n6108 , n6107 );
buf ( n6109 , n6027 );
buf ( n6110 , n6109 );
buf ( n6111 , n6110 );
buf ( n6112 , n6111 );
nand ( n6113 , n6108 , n6112 );
buf ( n6114 , n6113 );
nand ( n6115 , n6074 , n6093 , n6106 , n6114 );
buf ( n6116 , n6115 );
buf ( n6117 , n419 );
not ( n6118 , n6117 );
buf ( n6119 , n418 );
buf ( n6120 , n420 );
nand ( n6121 , n6119 , n6120 );
buf ( n6122 , n6121 );
buf ( n6123 , n6122 );
nand ( n6124 , n6118 , n6123 );
buf ( n6125 , n6124 );
buf ( n6126 , n419 );
not ( n6127 , n6126 );
buf ( n6128 , n418 );
nand ( n6129 , n6127 , n6128 );
buf ( n6130 , n6129 );
or ( n6131 , n6125 , n6130 );
not ( n6132 , n6131 );
buf ( n6133 , n418 );
buf ( n6134 , n422 );
nand ( n6135 , n6133 , n6134 );
buf ( n6136 , n6135 );
buf ( n6137 , n419 );
buf ( n6138 , n421 );
nand ( n6139 , n6137 , n6138 );
buf ( n6140 , n6139 );
nand ( n6141 , n6136 , n6140 );
buf ( n6142 , n6141 );
not ( n6143 , n6142 );
buf ( n6144 , n419 );
not ( n6145 , n6144 );
buf ( n6146 , n420 );
nor ( n6147 , n6145 , n6146 );
buf ( n6148 , n6147 );
buf ( n6149 , n6148 );
not ( n6150 , n6149 );
buf ( n6151 , n6150 );
buf ( n6152 , n6151 );
not ( n6153 , n6152 );
or ( n6154 , n6143 , n6153 );
buf ( n6155 , n418 );
buf ( n6156 , n421 );
nand ( n6157 , n6155 , n6156 );
buf ( n6158 , n6157 );
buf ( n6159 , n6158 );
nand ( n6160 , n6154 , n6159 );
buf ( n6161 , n6160 );
buf ( n6162 , n6161 );
buf ( n6163 , n419 );
not ( n6164 , n6163 );
buf ( n6165 , n6122 );
nor ( n6166 , n6164 , n6165 );
buf ( n6167 , n6166 );
buf ( n6168 , n6167 );
not ( n6169 , n6168 );
buf ( n6170 , n6125 );
nand ( n6171 , n6169 , n6170 );
buf ( n6172 , n6171 );
buf ( n6173 , n6172 );
nor ( n6174 , n6162 , n6173 );
buf ( n6175 , n6174 );
not ( n6176 , n6175 );
not ( n6177 , n420 );
buf ( n6178 , n418 );
buf ( n6179 , n423 );
nand ( n6180 , n6178 , n6179 );
buf ( n6181 , n6180 );
nand ( n6182 , n6177 , n6181 );
not ( n6183 , n6140 );
not ( n6184 , n6136 );
or ( n6185 , n6183 , n6184 );
buf ( n6186 , n419 );
buf ( n6187 , n422 );
nand ( n6188 , n6186 , n6187 );
buf ( n6189 , n6188 );
not ( n6190 , n6189 );
not ( n6191 , n6158 );
nand ( n6192 , n6190 , n6191 );
nand ( n6193 , n6185 , n6192 );
xor ( n6194 , n6182 , n6193 );
buf ( n6195 , n420 );
buf ( n6196 , n421 );
nand ( n6197 , n6195 , n6196 );
buf ( n6198 , n6197 );
buf ( n6199 , n6198 );
buf ( n6200 , n6189 );
nand ( n6201 , n6199 , n6200 );
buf ( n6202 , n6201 );
buf ( n6203 , n6018 );
buf ( n6204 , n419 );
buf ( n6205 , n423 );
nand ( n6206 , n6204 , n6205 );
buf ( n6207 , n6206 );
buf ( n6208 , n6207 );
nand ( n6209 , n6203 , n6208 );
buf ( n6210 , n6209 );
and ( n6211 , n6202 , n6210 );
and ( n6212 , n6194 , n6211 );
and ( n6213 , n6182 , n6193 );
or ( n6214 , n6212 , n6213 );
xor ( n6215 , n6191 , n6148 );
xnor ( n6216 , n6215 , n6141 );
or ( n6217 , n6214 , n6216 );
nand ( n6218 , n6176 , n6217 );
nor ( n6219 , n6132 , n6218 );
xor ( n6220 , n6001 , n6006 );
and ( n6221 , n6220 , n6022 );
and ( n6222 , n6001 , n6006 );
or ( n6223 , n6221 , n6222 );
buf ( n6224 , n6223 );
buf ( n6225 , n6224 );
nand ( n6226 , n421 , n422 );
nand ( n6227 , n420 , n423 );
xor ( n6228 , n6226 , n6227 );
nand ( n6229 , n424 , n419 );
xnor ( n6230 , n6228 , n6229 );
buf ( n6231 , n6230 );
xor ( n6232 , n6225 , n6231 );
buf ( n6233 , n425 );
buf ( n6234 , n418 );
nand ( n6235 , n6233 , n6234 );
buf ( n6236 , n6235 );
buf ( n6237 , n6236 );
not ( n6238 , n6237 );
buf ( n6239 , n6238 );
buf ( n6240 , n6239 );
buf ( n6241 , n418 );
buf ( n6242 , n421 );
xnor ( n6243 , n6241 , n6242 );
buf ( n6244 , n6243 );
buf ( n6245 , n6244 );
xor ( n6246 , n6240 , n6245 );
not ( n6247 , n419 );
not ( n6248 , n5980 );
or ( n6249 , n6247 , n6248 );
nand ( n6250 , n419 , n425 );
nand ( n6251 , n6249 , n6250 );
buf ( n6252 , n6251 );
xor ( n6253 , n6246 , n6252 );
buf ( n6254 , n6253 );
buf ( n6255 , n6254 );
and ( n6256 , n6232 , n6255 );
and ( n6257 , n6225 , n6231 );
or ( n6258 , n6256 , n6257 );
buf ( n6259 , n6258 );
buf ( n6260 , n6259 );
not ( n6261 , n6260 );
or ( n6262 , n6207 , n6018 );
nand ( n6263 , n6262 , n6210 );
xor ( n6264 , n6240 , n6245 );
and ( n6265 , n6264 , n6252 );
and ( n6266 , n6240 , n6245 );
or ( n6267 , n6265 , n6266 );
buf ( n6268 , n6267 );
xor ( n6269 , n6263 , n6268 );
and ( n6270 , n424 , n419 );
not ( n6271 , n6270 );
not ( n6272 , n420 );
not ( n6273 , n423 );
or ( n6274 , n6272 , n6273 );
nand ( n6275 , n421 , n422 );
nand ( n6276 , n6274 , n6275 );
not ( n6277 , n6276 );
or ( n6278 , n6271 , n6277 );
nand ( n6279 , n421 , n422 , n420 , n423 );
nand ( n6280 , n6278 , n6279 );
buf ( n6281 , n418 );
not ( n6282 , n6281 );
buf ( n6283 , n421 );
not ( n6284 , n6283 );
and ( n6285 , n6282 , n6284 );
buf ( n6286 , n424 );
buf ( n6287 , n418 );
and ( n6288 , n6286 , n6287 );
nor ( n6289 , n6285 , n6288 );
buf ( n6290 , n6289 );
and ( n6291 , n6280 , n6290 );
not ( n6292 , n6280 );
not ( n6293 , n6290 );
and ( n6294 , n6292 , n6293 );
nor ( n6295 , n6291 , n6294 );
xor ( n6296 , n6269 , n6295 );
buf ( n6297 , n6296 );
not ( n6298 , n6297 );
and ( n6299 , n6261 , n6298 );
xor ( n6300 , n5983 , n5992 );
and ( n6301 , n6300 , n6025 );
and ( n6302 , n5983 , n5992 );
or ( n6303 , n6301 , n6302 );
buf ( n6304 , n6303 );
xor ( n6305 , n6225 , n6231 );
xor ( n6306 , n6305 , n6255 );
buf ( n6307 , n6306 );
nor ( n6308 , n6304 , n6307 );
buf ( n6309 , n6308 );
nor ( n6310 , n6299 , n6309 );
buf ( n6311 , n6310 );
buf ( n6312 , n6311 );
buf ( n6313 , n423 );
not ( n6314 , n6313 );
buf ( n6315 , n6122 );
not ( n6316 , n6315 );
buf ( n6317 , n6316 );
buf ( n6318 , n6317 );
not ( n6319 , n6318 );
or ( n6320 , n6314 , n6319 );
buf ( n6321 , n6182 );
nand ( n6322 , n6320 , n6321 );
buf ( n6323 , n6322 );
buf ( n6324 , n6323 );
not ( n6325 , n6198 );
not ( n6326 , n6190 );
or ( n6327 , n6325 , n6326 );
nand ( n6328 , n419 , n422 );
nand ( n6329 , n6328 , n420 , n421 );
nand ( n6330 , n6327 , n6329 );
xor ( n6331 , n6330 , n6210 );
buf ( n6332 , n6331 );
xor ( n6333 , n6324 , n6332 );
buf ( n6334 , n421 );
not ( n6335 , n6334 );
buf ( n6336 , n6280 );
not ( n6337 , n6336 );
or ( n6338 , n6335 , n6337 );
buf ( n6339 , n424 );
buf ( n6340 , n418 );
nand ( n6341 , n6339 , n6340 );
buf ( n6342 , n6341 );
buf ( n6343 , n6342 );
nand ( n6344 , n6338 , n6343 );
buf ( n6345 , n6344 );
buf ( n6346 , n6345 );
xor ( n6347 , n6333 , n6346 );
buf ( n6348 , n6347 );
buf ( n6349 , n6295 );
not ( n6350 , n6349 );
buf ( n6351 , n6350 );
not ( n6352 , n6351 );
buf ( n6353 , n6263 );
not ( n6354 , n6353 );
buf ( n6355 , n6354 );
not ( n6356 , n6355 );
and ( n6357 , n6352 , n6356 );
buf ( n6358 , n6351 );
buf ( n6359 , n6355 );
nand ( n6360 , n6358 , n6359 );
buf ( n6361 , n6360 );
buf ( n6362 , n6268 );
buf ( n6363 , n6362 );
buf ( n6364 , n6363 );
and ( n6365 , n6361 , n6364 );
nor ( n6366 , n6357 , n6365 );
buf ( n6367 , n6366 );
not ( n6368 , n6367 );
buf ( n6369 , n6368 );
nor ( n6370 , n6348 , n6369 );
xor ( n6371 , n6324 , n6332 );
and ( n6372 , n6371 , n6346 );
and ( n6373 , n6324 , n6332 );
or ( n6374 , n6372 , n6373 );
buf ( n6375 , n6374 );
xor ( n6376 , n6182 , n6193 );
xor ( n6377 , n6376 , n6211 );
nor ( n6378 , n6375 , n6377 );
nor ( n6379 , n6370 , n6378 );
buf ( n6380 , n6379 );
nand ( n6381 , n6116 , n6219 , n6312 , n6380 );
buf ( n6382 , n6381 );
not ( n6383 , n6379 );
or ( n6384 , n6259 , n6296 );
nand ( n6385 , n6307 , n6304 );
not ( n6386 , n6385 );
nand ( n6387 , n6384 , n6386 );
nand ( n6388 , n6259 , n6296 );
nand ( n6389 , n6387 , n6388 );
not ( n6390 , n6389 );
or ( n6391 , n6383 , n6390 );
nand ( n6392 , n6375 , n6377 );
not ( n6393 , n6392 );
nand ( n6394 , n6348 , n6369 );
nor ( n6395 , n6378 , n6394 );
nor ( n6396 , n6393 , n6395 );
nand ( n6397 , n6391 , n6396 );
nand ( n6398 , n6397 , n6219 );
buf ( n6399 , n6398 );
buf ( n6400 , n6214 );
buf ( n6401 , n6216 );
nand ( n6402 , n6400 , n6401 );
buf ( n6403 , n6402 );
buf ( n6404 , n6403 );
buf ( n6405 , n6175 );
or ( n6406 , n6404 , n6405 );
buf ( n6407 , n6161 );
buf ( n6408 , n6172 );
nand ( n6409 , n6407 , n6408 );
buf ( n6410 , n6409 );
buf ( n6411 , n6410 );
nand ( n6412 , n6406 , n6411 );
buf ( n6413 , n6412 );
and ( n6414 , n6413 , n6131 );
buf ( n6415 , n6414 );
buf ( n6416 , n418 );
not ( n6417 , n6416 );
buf ( n6418 , n6125 );
buf ( n6419 , n6130 );
nand ( n6420 , n6418 , n6419 );
buf ( n6421 , n6420 );
buf ( n6422 , n6421 );
nand ( n6423 , n6417 , n6422 );
buf ( n6424 , n6423 );
buf ( n6425 , n6424 );
nor ( n6426 , n6415 , n6425 );
buf ( n6427 , n6426 );
buf ( n6428 , n6427 );
nand ( n6429 , n6382 , n6399 , n6428 );
buf ( n6430 , n6429 );
buf ( n6431 , n6430 );
not ( n6432 , n6431 );
buf ( n6433 , n6432 );
buf ( n6434 , n6433 );
not ( n6435 , n6434 );
buf ( n6436 , n6435 );
not ( n6437 , n6436 );
or ( n6438 , n5842 , n6437 );
buf ( n6439 , n411 );
not ( n6440 , n6439 );
buf ( n6441 , n6433 );
nand ( n6442 , n6440 , n6441 );
buf ( n6443 , n6442 );
nand ( n6444 , n6438 , n6443 );
nand ( n6445 , n5841 , n6444 );
not ( n6446 , n6445 );
buf ( n6447 , n6433 );
not ( n6448 , n6447 );
buf ( n6449 , n416 );
not ( n6450 , n6449 );
buf ( n6451 , n6450 );
buf ( n6452 , n6451 );
buf ( n6453 , n415 );
and ( n6454 , n6452 , n6453 );
buf ( n6455 , n6454 );
buf ( n6456 , n6455 );
nand ( n6457 , n6448 , n6456 );
buf ( n6458 , n6457 );
buf ( n6459 , n415 );
not ( n6460 , n6459 );
buf ( n6461 , n6430 );
not ( n6462 , n6461 );
or ( n6463 , n6460 , n6462 );
buf ( n6464 , n6433 );
buf ( n6465 , n415 );
not ( n6466 , n6465 );
buf ( n6467 , n6466 );
buf ( n6468 , n6467 );
nand ( n6469 , n6464 , n6468 );
buf ( n6470 , n6469 );
buf ( n6471 , n6470 );
nand ( n6472 , n6463 , n6471 );
buf ( n6473 , n6472 );
buf ( n6474 , n6473 );
buf ( n6475 , n416 );
nand ( n6476 , n6474 , n6475 );
buf ( n6477 , n6476 );
nand ( n6478 , n6458 , n6477 );
not ( n6479 , n6478 );
or ( n6480 , n6446 , n6479 );
buf ( n6481 , n6477 );
buf ( n6482 , n6458 );
nand ( n6483 , n6481 , n6482 );
buf ( n6484 , n6483 );
buf ( n6485 , n6484 );
not ( n6486 , n6485 );
and ( n6487 , n6444 , n5841 );
buf ( n6488 , n6487 );
nand ( n6489 , n6486 , n6488 );
buf ( n6490 , n6489 );
nand ( n6491 , n6480 , n6490 );
not ( n6492 , n413 );
not ( n6493 , n6436 );
or ( n6494 , n6492 , n6493 );
buf ( n6495 , n6433 );
not ( n6496 , n413 );
buf ( n6497 , n6496 );
nand ( n6498 , n6495 , n6497 );
buf ( n6499 , n6498 );
nand ( n6500 , n6494 , n6499 );
buf ( n6501 , n6496 );
buf ( n6502 , n414 );
not ( n6503 , n6502 );
buf ( n6504 , n6503 );
buf ( n6505 , n6504 );
and ( n6506 , n6501 , n6505 );
buf ( n6507 , n413 );
buf ( n6508 , n414 );
and ( n6509 , n6507 , n6508 );
nor ( n6510 , n6506 , n6509 );
buf ( n6511 , n6510 );
not ( n6512 , n415 );
not ( n6513 , n414 );
or ( n6514 , n6512 , n6513 );
buf ( n6515 , n6467 );
buf ( n6516 , n6504 );
nand ( n6517 , n6515 , n6516 );
buf ( n6518 , n6517 );
nand ( n6519 , n6514 , n6518 );
and ( n6520 , n6511 , n6519 );
buf ( n6521 , n6520 );
not ( n6522 , n6521 );
buf ( n6523 , n6522 );
nand ( n6524 , n6523 , n6519 );
nand ( n6525 , n6500 , n6524 );
buf ( n6526 , n6525 );
buf ( n6527 , n6433 );
xor ( n6528 , n410 , n411 );
buf ( n6529 , n6528 );
nand ( n6530 , n6527 , n6529 );
buf ( n6531 , n6530 );
not ( n6532 , n6531 );
buf ( n6533 , n6528 );
not ( n6534 , n6533 );
buf ( n6535 , n6534 );
buf ( n6536 , n6535 );
buf ( n6537 , n410 );
and ( n6538 , n6536 , n6537 );
buf ( n6539 , n6538 );
and ( n6540 , n6539 , n6433 );
nor ( n6541 , n6532 , n6540 );
buf ( n6542 , n6541 );
nand ( n6543 , n6526 , n6542 );
and ( n6544 , n6491 , n6543 );
not ( n6545 , n6491 );
not ( n6546 , n6543 );
and ( n6547 , n6545 , n6546 );
nor ( n6548 , n6544 , n6547 );
not ( n6549 , n6548 );
not ( n6550 , n6525 );
not ( n6551 , n6541 );
nor ( n6552 , n6550 , n6551 );
not ( n6553 , n6552 );
not ( n6554 , n6519 );
not ( n6555 , n6523 );
or ( n6556 , n6554 , n6555 );
nand ( n6557 , n6556 , n6500 );
buf ( n6558 , n6557 );
not ( n6559 , n6558 );
buf ( n6560 , n6559 );
buf ( n6561 , n6560 );
buf ( n6562 , n6551 );
nand ( n6563 , n6561 , n6562 );
buf ( n6564 , n6563 );
nand ( n6565 , n6553 , n6564 );
not ( n6566 , n6565 );
nand ( n6567 , n6549 , n6566 );
not ( n6568 , n6567 );
buf ( n6569 , n6445 );
buf ( n6570 , n6552 );
nand ( n6571 , n6569 , n6570 );
buf ( n6572 , n6571 );
not ( n6573 , n6572 );
buf ( n6574 , n6478 );
not ( n6575 , n6574 );
or ( n6576 , n6573 , n6575 );
not ( n6577 , n6552 );
buf ( n6578 , n6577 );
buf ( n6579 , n6487 );
buf ( n6580 , n6579 );
buf ( n6581 , n6580 );
buf ( n6582 , n6581 );
nand ( n6583 , n6578 , n6582 );
buf ( n6584 , n6583 );
nand ( n6585 , n6576 , n6584 );
not ( n6586 , n6585 );
or ( n6587 , n6568 , n6586 );
nand ( n6588 , n6548 , n6565 );
nand ( n6589 , n6587 , n6588 );
buf ( n6590 , n6589 );
not ( n6591 , n6590 );
buf ( n6592 , n6591 );
buf ( n6593 , n6585 );
not ( n6594 , n6593 );
not ( n6595 , n6549 );
not ( n6596 , n6565 );
or ( n6597 , n6595 , n6596 );
nand ( n6598 , n6548 , n6566 );
nand ( n6599 , n6597 , n6598 );
not ( n6600 , n6599 );
buf ( n6601 , n6600 );
not ( n6602 , n6601 );
or ( n6603 , n6594 , n6602 );
buf ( n6604 , n6599 );
buf ( n6605 , n6585 );
not ( n6606 , n6605 );
buf ( n6607 , n6606 );
buf ( n6608 , n6607 );
nand ( n6609 , n6604 , n6608 );
buf ( n6610 , n6609 );
buf ( n6611 , n6610 );
nand ( n6612 , n6603 , n6611 );
buf ( n6613 , n6612 );
buf ( n6614 , n376 );
buf ( n6615 , n382 );
nand ( n6616 , n6614 , n6615 );
buf ( n6617 , n6616 );
nand ( n6618 , n374 , n380 );
or ( n6619 , n6617 , n6618 );
nand ( n6620 , n377 , n379 );
not ( n6621 , n6620 );
nand ( n6622 , n375 , n381 );
not ( n6623 , n6622 );
or ( n6624 , n6621 , n6623 );
or ( n6625 , n6620 , n6622 );
nand ( n6626 , n372 , n384 );
nand ( n6627 , n6625 , n6626 );
nand ( n6628 , n6624 , n6627 );
xor ( n6629 , n6619 , n6628 );
buf ( n6630 , n374 );
buf ( n6631 , n381 );
nand ( n6632 , n6630 , n6631 );
buf ( n6633 , n6632 );
buf ( n6634 , n373 );
buf ( n6635 , n382 );
nand ( n6636 , n6634 , n6635 );
buf ( n6637 , n6636 );
buf ( n6638 , n370 );
buf ( n6639 , n385 );
nand ( n6640 , n6638 , n6639 );
buf ( n6641 , n6640 );
nand ( n6642 , n6633 , n6637 , n6641 );
not ( n6643 , n6633 );
not ( n6644 , n6641 );
nand ( n6645 , n6643 , n6637 , n6644 );
not ( n6646 , n6637 );
nand ( n6647 , n6646 , n6641 , n6643 );
nand ( n6648 , n6644 , n6646 , n6633 );
nand ( n6649 , n6642 , n6645 , n6647 , n6648 );
xor ( n6650 , n6629 , n6649 );
buf ( n6651 , n6619 );
buf ( n6652 , n376 );
buf ( n6653 , n380 );
nand ( n6654 , n6652 , n6653 );
buf ( n6655 , n6654 );
buf ( n6656 , n6655 );
buf ( n6657 , n374 );
buf ( n6658 , n382 );
nand ( n6659 , n6657 , n6658 );
buf ( n6660 , n6659 );
buf ( n6661 , n6660 );
nand ( n6662 , n6656 , n6661 );
buf ( n6663 , n6662 );
buf ( n6664 , n6663 );
nand ( n6665 , n6651 , n6664 );
buf ( n6666 , n6665 );
not ( n6667 , n6666 );
nand ( n6668 , n375 , n381 );
xor ( n6669 , n6668 , n6620 );
xor ( n6670 , n6669 , n6626 );
buf ( n6671 , n372 );
buf ( n6672 , n385 );
nand ( n6673 , n6671 , n6672 );
buf ( n6674 , n6673 );
not ( n6675 , n6674 );
buf ( n6676 , n376 );
buf ( n6677 , n381 );
nand ( n6678 , n6676 , n6677 );
buf ( n6679 , n6678 );
not ( n6680 , n6679 );
or ( n6681 , n6675 , n6680 );
not ( n6682 , n6674 );
not ( n6683 , n6682 );
not ( n6684 , n6679 );
not ( n6685 , n6684 );
or ( n6686 , n6683 , n6685 );
nand ( n6687 , n374 , n383 );
nand ( n6688 , n6686 , n6687 );
nand ( n6689 , n6681 , n6688 );
or ( n6690 , n6670 , n6689 );
not ( n6691 , n6690 );
or ( n6692 , n6667 , n6691 );
nand ( n6693 , n6670 , n6689 );
nand ( n6694 , n6692 , n6693 );
xor ( n6695 , n6650 , n6694 );
buf ( n6696 , n372 );
buf ( n6697 , n383 );
nand ( n6698 , n6696 , n6697 );
buf ( n6699 , n6698 );
not ( n6700 , n6699 );
buf ( n6701 , n371 );
buf ( n6702 , n384 );
nand ( n6703 , n6701 , n6702 );
buf ( n6704 , n6703 );
not ( n6705 , n6704 );
or ( n6706 , n6700 , n6705 );
nand ( n6707 , n371 , n383 );
not ( n6708 , n6707 );
nand ( n6709 , n6708 , n372 , n384 );
nand ( n6710 , n6706 , n6709 );
nand ( n6711 , n376 , n379 );
nand ( n6712 , n377 , n378 );
xor ( n6713 , n6711 , n6712 );
buf ( n6714 , n375 );
buf ( n6715 , n380 );
nand ( n6716 , n6714 , n6715 );
buf ( n6717 , n6716 );
not ( n6718 , n6717 );
and ( n6719 , n6713 , n6718 );
not ( n6720 , n6713 );
and ( n6721 , n6720 , n6717 );
or ( n6722 , n6719 , n6721 );
xor ( n6723 , n6710 , n6722 );
nand ( n6724 , n377 , n380 );
buf ( n6725 , n6724 );
buf ( n6726 , n373 );
buf ( n6727 , n383 );
nand ( n6728 , n6726 , n6727 );
buf ( n6729 , n6728 );
buf ( n6730 , n6729 );
or ( n6731 , n6725 , n6730 );
buf ( n6732 , n371 );
buf ( n6733 , n385 );
nand ( n6734 , n6732 , n6733 );
buf ( n6735 , n6734 );
buf ( n6736 , n6735 );
nand ( n6737 , n6731 , n6736 );
buf ( n6738 , n6737 );
buf ( n6739 , n6724 );
buf ( n6740 , n6729 );
nand ( n6741 , n6739 , n6740 );
buf ( n6742 , n6741 );
nand ( n6743 , n6738 , n6742 );
xor ( n6744 , n6723 , n6743 );
and ( n6745 , n6695 , n6744 );
and ( n6746 , n6650 , n6694 );
or ( n6747 , n6745 , n6746 );
buf ( n6748 , n6747 );
xor ( n6749 , n6710 , n6722 );
and ( n6750 , n6749 , n6743 );
and ( n6751 , n6710 , n6722 );
or ( n6752 , n6750 , n6751 );
nand ( n6753 , n6633 , n6637 );
not ( n6754 , n6643 );
not ( n6755 , n6646 );
or ( n6756 , n6754 , n6755 );
nand ( n6757 , n6756 , n6641 );
nand ( n6758 , n6753 , n6757 );
nand ( n6759 , n371 , n383 );
xor ( n6760 , n6759 , n6618 );
nand ( n6761 , n376 , n378 );
xor ( n6762 , n6760 , n6761 );
not ( n6763 , n6762 );
not ( n6764 , n6709 );
nand ( n6765 , n6763 , n6764 );
nand ( n6766 , n6762 , n6709 );
nand ( n6767 , n6765 , n6766 );
and ( n6768 , n6758 , n6767 );
not ( n6769 , n6758 );
and ( n6770 , n6762 , n6709 );
not ( n6771 , n6762 );
and ( n6772 , n6771 , n6764 );
nor ( n6773 , n6770 , n6772 );
and ( n6774 , n6769 , n6773 );
or ( n6775 , n6768 , n6774 );
xor ( n6776 , n6752 , n6775 );
buf ( n6777 , n372 );
buf ( n6778 , n382 );
nand ( n6779 , n6777 , n6778 );
buf ( n6780 , n6779 );
buf ( n6781 , n6780 );
not ( n6782 , n6781 );
buf ( n6783 , n6782 );
buf ( n6784 , n370 );
buf ( n6785 , n384 );
nand ( n6786 , n6784 , n6785 );
buf ( n6787 , n6786 );
xor ( n6788 , n6783 , n6787 );
nand ( n6789 , n376 , n379 );
not ( n6790 , n6789 );
not ( n6791 , n6790 );
not ( n6792 , n6718 );
or ( n6793 , n6791 , n6792 );
nand ( n6794 , n6793 , n6712 );
nand ( n6795 , n6717 , n6789 );
nand ( n6796 , n6794 , n6795 );
xnor ( n6797 , n6788 , n6796 );
buf ( n6798 , n373 );
buf ( n6799 , n381 );
nand ( n6800 , n6798 , n6799 );
buf ( n6801 , n6800 );
buf ( n6802 , n6801 );
not ( n6803 , n6802 );
buf ( n6804 , n375 );
buf ( n6805 , n379 );
nand ( n6806 , n6804 , n6805 );
buf ( n6807 , n6806 );
buf ( n6808 , n6807 );
not ( n6809 , n6808 );
or ( n6810 , n6803 , n6809 );
nand ( n6811 , n373 , n379 );
not ( n6812 , n6811 );
nand ( n6813 , n6812 , n375 , n381 );
buf ( n6814 , n6813 );
nand ( n6815 , n6810 , n6814 );
buf ( n6816 , n6815 );
buf ( n6817 , n6816 );
not ( n6818 , n6817 );
buf ( n6819 , n6818 );
xor ( n6820 , n6797 , n6819 );
xor ( n6821 , n6619 , n6628 );
and ( n6822 , n6821 , n6649 );
and ( n6823 , n6619 , n6628 );
or ( n6824 , n6822 , n6823 );
not ( n6825 , n6824 );
xor ( n6826 , n6820 , n6825 );
xor ( n6827 , n6776 , n6826 );
buf ( n6828 , n6827 );
xor ( n6829 , n6748 , n6828 );
not ( n6830 , n6528 );
nand ( n6831 , n5973 , n5934 );
not ( n6832 , n6087 );
not ( n6833 , n5872 );
nand ( n6834 , n6833 , n5898 );
nand ( n6835 , n6832 , n6834 );
nand ( n6836 , n6835 , n6085 );
nand ( n6837 , n6831 , n6836 );
buf ( n6838 , n6831 );
buf ( n6839 , n5928 );
buf ( n6840 , n6071 );
nand ( n6841 , n6838 , n6839 , n6840 );
buf ( n6842 , n6841 );
buf ( n6843 , n6103 );
not ( n6844 , n6843 );
buf ( n6845 , n6844 );
nand ( n6846 , n6837 , n6842 , n6845 );
nand ( n6847 , n6098 , n6114 );
and ( n6848 , n6846 , n6847 );
not ( n6849 , n6846 );
not ( n6850 , n6847 );
and ( n6851 , n6849 , n6850 );
nor ( n6852 , n6848 , n6851 );
buf ( n6853 , n6852 );
not ( n6854 , n6853 );
buf ( n6855 , n6854 );
not ( n6856 , n6855 );
or ( n6857 , n6830 , n6856 );
buf ( n6858 , n6831 );
buf ( n6859 , n6845 );
and ( n6860 , n6858 , n6859 );
buf ( n6861 , n6860 );
not ( n6862 , n6836 );
buf ( n6863 , n5928 );
buf ( n6864 , n6071 );
nand ( n6865 , n6863 , n6864 );
buf ( n6866 , n6865 );
nand ( n6867 , n6862 , n6866 );
xor ( n6868 , n6861 , n6867 );
buf ( n6869 , n6868 );
buf ( n6870 , n6539 );
nand ( n6871 , n6869 , n6870 );
buf ( n6872 , n6871 );
nand ( n6873 , n6857 , n6872 );
buf ( n6874 , n6873 );
xor ( n6875 , n6829 , n6874 );
buf ( n6876 , n6875 );
buf ( n6877 , n6876 );
xor ( n6878 , n6650 , n6694 );
xor ( n6879 , n6878 , n6744 );
buf ( n6880 , n6879 );
not ( n6881 , n6880 );
xor ( n6882 , n6729 , n6735 );
not ( n6883 , n6724 );
xor ( n6884 , n6882 , n6883 );
not ( n6885 , n6884 );
buf ( n6886 , n375 );
buf ( n6887 , n382 );
nand ( n6888 , n6886 , n6887 );
buf ( n6889 , n6888 );
buf ( n6890 , n6889 );
not ( n6891 , n6890 );
buf ( n6892 , n6724 );
nand ( n6893 , n6891 , n6892 );
buf ( n6894 , n6893 );
buf ( n6895 , n6894 );
buf ( n6896 , n373 );
buf ( n6897 , n384 );
nand ( n6898 , n6896 , n6897 );
buf ( n6899 , n6898 );
buf ( n6900 , n6899 );
and ( n6901 , n6895 , n6900 );
buf ( n6902 , n6889 );
not ( n6903 , n6902 );
buf ( n6904 , n6724 );
nor ( n6905 , n6903 , n6904 );
buf ( n6906 , n6905 );
buf ( n6907 , n6906 );
nor ( n6908 , n6901 , n6907 );
buf ( n6909 , n6908 );
not ( n6910 , n6909 );
and ( n6911 , n6885 , n6910 );
xor ( n6912 , n6687 , n6682 );
xnor ( n6913 , n6912 , n6679 );
not ( n6914 , n6913 );
buf ( n6915 , n6637 );
not ( n6916 , n6915 );
buf ( n6917 , n376 );
buf ( n6918 , n385 );
nand ( n6919 , n6917 , n6918 );
buf ( n6920 , n6919 );
buf ( n6921 , n6920 );
not ( n6922 , n6921 );
buf ( n6923 , n6922 );
buf ( n6924 , n6923 );
nand ( n6925 , n6916 , n6924 );
buf ( n6926 , n6925 );
not ( n6927 , n6926 );
nand ( n6928 , n374 , n384 );
not ( n6929 , n6928 );
nand ( n6930 , n377 , n381 );
not ( n6931 , n6930 );
or ( n6932 , n6929 , n6931 );
buf ( n6933 , n375 );
buf ( n6934 , n383 );
nand ( n6935 , n6933 , n6934 );
buf ( n6936 , n6935 );
not ( n6937 , n6936 );
nor ( n6938 , n6928 , n6930 );
or ( n6939 , n6937 , n6938 );
nand ( n6940 , n6932 , n6939 );
not ( n6941 , n6940 );
nand ( n6942 , n6927 , n6941 );
not ( n6943 , n6942 );
or ( n6944 , n6914 , n6943 );
nand ( n6945 , n6926 , n6940 );
nand ( n6946 , n6944 , n6945 );
nand ( n6947 , n6909 , n6884 );
and ( n6948 , n6946 , n6947 );
nor ( n6949 , n6911 , n6948 );
buf ( n6950 , n6949 );
nand ( n6951 , n6881 , n6950 );
buf ( n6952 , n6951 );
buf ( n6953 , n6952 );
not ( n6954 , n6953 );
xor ( n6955 , n6670 , n6689 );
xor ( n6956 , n6955 , n6666 );
buf ( n6957 , n6956 );
not ( n6958 , n6957 );
not ( n6959 , n6071 );
buf ( n6960 , n5925 );
not ( n6961 , n6960 );
buf ( n6962 , n6961 );
not ( n6963 , n6962 );
or ( n6964 , n6959 , n6963 );
nand ( n6965 , n6964 , n6087 );
not ( n6966 , n6965 );
nor ( n6967 , n5872 , n5901 );
not ( n6968 , n6967 );
nand ( n6969 , n6968 , n6085 );
not ( n6970 , n6969 );
or ( n6971 , n6966 , n6970 );
or ( n6972 , n6965 , n6969 );
nand ( n6973 , n6971 , n6972 );
buf ( n6974 , n6973 );
buf ( n6975 , n6528 );
nand ( n6976 , n6974 , n6975 );
buf ( n6977 , n6976 );
buf ( n6978 , n6977 );
not ( n6979 , n6978 );
buf ( n6980 , n6979 );
buf ( n6981 , n6980 );
not ( n6982 , n6981 );
or ( n6983 , n6958 , n6982 );
buf ( n6984 , n6956 );
not ( n6985 , n6984 );
buf ( n6986 , n6985 );
buf ( n6987 , n6986 );
not ( n6988 , n6987 );
buf ( n6989 , n6977 );
not ( n6990 , n6989 );
or ( n6991 , n6988 , n6990 );
xor ( n6992 , n6909 , n6884 );
xor ( n6993 , n6992 , n6946 );
buf ( n6994 , n6993 );
nand ( n6995 , n6991 , n6994 );
buf ( n6996 , n6995 );
buf ( n6997 , n6996 );
nand ( n6998 , n6983 , n6997 );
buf ( n6999 , n6998 );
buf ( n7000 , n6999 );
not ( n7001 , n7000 );
or ( n7002 , n6954 , n7001 );
buf ( n7003 , n6879 );
not ( n7004 , n6949 );
buf ( n7005 , n7004 );
nand ( n7006 , n7003 , n7005 );
buf ( n7007 , n7006 );
buf ( n7008 , n7007 );
nand ( n7009 , n7002 , n7008 );
buf ( n7010 , n7009 );
buf ( n7011 , n7010 );
xor ( n7012 , n6877 , n7011 );
not ( n7013 , n5832 );
buf ( n7014 , n7013 );
not ( n7015 , n7014 );
or ( n7016 , n6307 , n6304 );
not ( n7017 , n7016 );
not ( n7018 , n6115 );
or ( n7019 , n7017 , n7018 );
nand ( n7020 , n6307 , n6304 );
nand ( n7021 , n7019 , n7020 );
buf ( n7022 , n6259 );
buf ( n7023 , n6296 );
or ( n7024 , n7022 , n7023 );
buf ( n7025 , n7024 );
nand ( n7026 , n7025 , n6388 );
not ( n7027 , n7026 );
and ( n7028 , n7021 , n7027 );
not ( n7029 , n7021 );
and ( n7030 , n7029 , n7026 );
nor ( n7031 , n7028 , n7030 );
buf ( n7032 , n7031 );
not ( n7033 , n7032 );
buf ( n7034 , n7033 );
and ( n7035 , n411 , n7034 );
not ( n7036 , n411 );
and ( n7037 , n7036 , n7031 );
or ( n7038 , n7035 , n7037 );
buf ( n7039 , n7038 );
not ( n7040 , n7039 );
or ( n7041 , n7015 , n7040 );
buf ( n7042 , n411 );
and ( n7043 , n7016 , n7020 );
xor ( n7044 , n7043 , n6116 );
buf ( n7045 , n7044 );
and ( n7046 , n7042 , n7045 );
not ( n7047 , n7042 );
buf ( n7048 , n7044 );
not ( n7049 , n7048 );
buf ( n7050 , n7049 );
buf ( n7051 , n7050 );
and ( n7052 , n7047 , n7051 );
nor ( n7053 , n7046 , n7052 );
buf ( n7054 , n7053 );
buf ( n7055 , n7054 );
buf ( n7056 , n5837 );
nand ( n7057 , n7055 , n7056 );
buf ( n7058 , n7057 );
buf ( n7059 , n7058 );
nand ( n7060 , n7041 , n7059 );
buf ( n7061 , n7060 );
buf ( n7062 , n7061 );
xor ( n7063 , n7012 , n7062 );
buf ( n7064 , n7063 );
buf ( n7065 , n7064 );
xor ( n7066 , n6899 , n6889 );
and ( n7067 , n7066 , n6883 );
not ( n7068 , n7066 );
and ( n7069 , n7068 , n6724 );
nor ( n7070 , n7067 , n7069 );
buf ( n7071 , n7070 );
not ( n7072 , n6941 );
not ( n7073 , n6926 );
or ( n7074 , n7072 , n7073 );
nand ( n7075 , n6927 , n6940 );
nand ( n7076 , n7074 , n7075 );
and ( n7077 , n7076 , n6913 );
not ( n7078 , n7076 );
not ( n7079 , n6913 );
and ( n7080 , n7078 , n7079 );
nor ( n7081 , n7077 , n7080 );
buf ( n7082 , n7081 );
xor ( n7083 , n7071 , n7082 );
buf ( n7084 , n374 );
buf ( n7085 , n385 );
nand ( n7086 , n7084 , n7085 );
buf ( n7087 , n7086 );
buf ( n7088 , n7087 );
not ( n7089 , n7088 );
buf ( n7090 , n7089 );
buf ( n7091 , n7090 );
not ( n7092 , n7091 );
xor ( n7093 , n6930 , n6936 );
buf ( n7094 , n7093 );
buf ( n7095 , n6928 );
xnor ( n7096 , n7094 , n7095 );
buf ( n7097 , n7096 );
buf ( n7098 , n7097 );
not ( n7099 , n7098 );
or ( n7100 , n7092 , n7099 );
buf ( n7101 , n377 );
buf ( n7102 , n382 );
nand ( n7103 , n7101 , n7102 );
buf ( n7104 , n7103 );
buf ( n7105 , n375 );
buf ( n7106 , n384 );
nand ( n7107 , n7105 , n7106 );
buf ( n7108 , n7107 );
xor ( n7109 , n7104 , n7108 );
nand ( n7110 , n376 , n383 );
and ( n7111 , n7109 , n7110 );
and ( n7112 , n7104 , n7108 );
nor ( n7113 , n7111 , n7112 );
not ( n7114 , n7113 );
buf ( n7115 , n7114 );
nand ( n7116 , n7100 , n7115 );
buf ( n7117 , n7116 );
buf ( n7118 , n7117 );
buf ( n7119 , n7097 );
not ( n7120 , n7119 );
buf ( n7121 , n7120 );
buf ( n7122 , n7121 );
buf ( n7123 , n7087 );
nand ( n7124 , n7122 , n7123 );
buf ( n7125 , n7124 );
buf ( n7126 , n7125 );
nand ( n7127 , n7118 , n7126 );
buf ( n7128 , n7127 );
buf ( n7129 , n7128 );
and ( n7130 , n7083 , n7129 );
and ( n7131 , n7071 , n7082 );
or ( n7132 , n7130 , n7131 );
buf ( n7133 , n7132 );
buf ( n7134 , n7133 );
buf ( n7135 , n7108 );
buf ( n7136 , n6920 );
nor ( n7137 , n7135 , n7136 );
buf ( n7138 , n7137 );
buf ( n7139 , n7138 );
buf ( n7140 , n7087 );
nand ( n7141 , n7139 , n7140 );
buf ( n7142 , n7141 );
not ( n7143 , n7142 );
xor ( n7144 , n7104 , n7108 );
xor ( n7145 , n7144 , n7110 );
not ( n7146 , n7145 );
or ( n7147 , n7143 , n7146 );
buf ( n7148 , n7138 );
not ( n7149 , n7148 );
buf ( n7150 , n7149 );
buf ( n7151 , n7150 );
buf ( n7152 , n7090 );
nand ( n7153 , n7151 , n7152 );
buf ( n7154 , n7153 );
nand ( n7155 , n7147 , n7154 );
buf ( n7156 , n373 );
buf ( n7157 , n385 );
nand ( n7158 , n7156 , n7157 );
buf ( n7159 , n7158 );
buf ( n7160 , n7159 );
not ( n7161 , n7160 );
buf ( n7162 , n6617 );
not ( n7163 , n7162 );
or ( n7164 , n7161 , n7163 );
buf ( n7165 , n6926 );
nand ( n7166 , n7164 , n7165 );
buf ( n7167 , n7166 );
and ( n7168 , n7155 , n7167 );
not ( n7169 , n7090 );
not ( n7170 , n7113 );
or ( n7171 , n7169 , n7170 );
nand ( n7172 , n7114 , n7087 );
nand ( n7173 , n7171 , n7172 );
xnor ( n7174 , n7173 , n7121 );
or ( n7175 , n7168 , n7174 );
or ( n7176 , n7155 , n7167 );
nand ( n7177 , n7175 , n7176 );
buf ( n7178 , n7177 );
not ( n7179 , n7178 );
buf ( n7180 , n412 );
not ( n7181 , n7180 );
buf ( n7182 , n6496 );
nand ( n7183 , n7181 , n7182 );
buf ( n7184 , n7183 );
buf ( n7185 , n7184 );
not ( n7186 , n7185 );
buf ( n7187 , n6973 );
not ( n7188 , n7187 );
or ( n7189 , n7186 , n7188 );
buf ( n7190 , n412 );
buf ( n7191 , n413 );
and ( n7192 , n7190 , n7191 );
buf ( n7193 , n411 );
not ( n7194 , n7193 );
buf ( n7195 , n7194 );
buf ( n7196 , n7195 );
nor ( n7197 , n7192 , n7196 );
buf ( n7198 , n7197 );
buf ( n7199 , n7198 );
nand ( n7200 , n7189 , n7199 );
buf ( n7201 , n7200 );
buf ( n7202 , n7201 );
not ( n7203 , n7202 );
or ( n7204 , n7179 , n7203 );
xor ( n7205 , n7071 , n7082 );
xor ( n7206 , n7205 , n7129 );
buf ( n7207 , n7206 );
buf ( n7208 , n7207 );
nand ( n7209 , n7204 , n7208 );
buf ( n7210 , n7209 );
buf ( n7211 , n7210 );
buf ( n7212 , n7201 );
buf ( n7213 , n7177 );
or ( n7214 , n7212 , n7213 );
buf ( n7215 , n7214 );
buf ( n7216 , n7215 );
nand ( n7217 , n7211 , n7216 );
buf ( n7218 , n7217 );
buf ( n7219 , n7218 );
xor ( n7220 , n7134 , n7219 );
buf ( n7221 , n6956 );
buf ( n7222 , n6993 );
xor ( n7223 , n7221 , n7222 );
buf ( n7224 , n6977 );
xnor ( n7225 , n7223 , n7224 );
buf ( n7226 , n7225 );
buf ( n7227 , n7226 );
and ( n7228 , n7220 , n7227 );
and ( n7229 , n7134 , n7219 );
or ( n7230 , n7228 , n7229 );
buf ( n7231 , n7230 );
buf ( n7232 , n7231 );
buf ( n7233 , n6520 );
not ( n7234 , n7233 );
xnor ( n7235 , n6496 , n7031 );
buf ( n7236 , n7235 );
not ( n7237 , n7236 );
or ( n7238 , n7234 , n7237 );
buf ( n7239 , n6496 );
not ( n7240 , n7239 );
not ( n7241 , n6115 );
not ( n7242 , n6311 );
or ( n7243 , n7241 , n7242 );
buf ( n7244 , n6389 );
not ( n7245 , n7244 );
buf ( n7246 , n7245 );
nand ( n7247 , n7243 , n7246 );
not ( n7248 , n6394 );
nor ( n7249 , n6370 , n7248 );
xor ( n7250 , n7247 , n7249 );
buf ( n7251 , n7250 );
not ( n7252 , n7251 );
or ( n7253 , n7240 , n7252 );
buf ( n7254 , n7250 );
buf ( n7255 , n6496 );
or ( n7256 , n7254 , n7255 );
nand ( n7257 , n7253 , n7256 );
buf ( n7258 , n7257 );
buf ( n7259 , n7258 );
not ( n7260 , n6519 );
buf ( n7261 , n7260 );
nand ( n7262 , n7259 , n7261 );
buf ( n7263 , n7262 );
buf ( n7264 , n7263 );
nand ( n7265 , n7238 , n7264 );
buf ( n7266 , n7265 );
buf ( n7267 , n7266 );
xor ( n7268 , n7232 , n7267 );
buf ( n7269 , n415 );
not ( n7270 , n7269 );
not ( n7271 , n6378 );
nand ( n7272 , n7271 , n6392 );
not ( n7273 , n7272 );
not ( n7274 , n6311 );
not ( n7275 , n6366 );
nor ( n7276 , n7275 , n6348 );
nor ( n7277 , n7274 , n7276 );
not ( n7278 , n7277 );
not ( n7279 , n6116 );
or ( n7280 , n7278 , n7279 );
nand ( n7281 , n6387 , n6388 );
buf ( n7282 , n7281 );
buf ( n7283 , n6370 );
not ( n7284 , n7283 );
buf ( n7285 , n7284 );
buf ( n7286 , n7285 );
and ( n7287 , n7282 , n7286 );
buf ( n7288 , n7248 );
nor ( n7289 , n7287 , n7288 );
buf ( n7290 , n7289 );
nand ( n7291 , n7280 , n7290 );
not ( n7292 , n7291 );
or ( n7293 , n7273 , n7292 );
or ( n7294 , n7272 , n7291 );
nand ( n7295 , n7293 , n7294 );
buf ( n7296 , n7295 );
not ( n7297 , n7296 );
buf ( n7298 , n7297 );
buf ( n7299 , n7298 );
not ( n7300 , n7299 );
or ( n7301 , n7270 , n7300 );
and ( n7302 , n7291 , n7272 );
not ( n7303 , n7291 );
not ( n7304 , n7272 );
and ( n7305 , n7303 , n7304 );
nor ( n7306 , n7302 , n7305 );
buf ( n7307 , n7306 );
not ( n7308 , n7307 );
buf ( n7309 , n6467 );
nand ( n7310 , n7308 , n7309 );
buf ( n7311 , n7310 );
buf ( n7312 , n7311 );
nand ( n7313 , n7301 , n7312 );
buf ( n7314 , n7313 );
not ( n7315 , n7314 );
not ( n7316 , n6455 );
or ( n7317 , n7315 , n7316 );
buf ( n7318 , n415 );
and ( n7319 , n6311 , n6379 );
not ( n7320 , n7319 );
not ( n7321 , n6116 );
or ( n7322 , n7320 , n7321 );
buf ( n7323 , n6397 );
not ( n7324 , n7323 );
buf ( n7325 , n7324 );
nand ( n7326 , n7322 , n7325 );
nand ( n7327 , n6217 , n6403 );
not ( n7328 , n7327 );
and ( n7329 , n7326 , n7328 );
not ( n7330 , n7326 );
and ( n7331 , n7330 , n7327 );
nor ( n7332 , n7329 , n7331 );
buf ( n7333 , n7332 );
not ( n7334 , n7333 );
buf ( n7335 , n7334 );
buf ( n7336 , n7335 );
and ( n7337 , n7318 , n7336 );
not ( n7338 , n7318 );
buf ( n7339 , n7332 );
not ( n7340 , n7339 );
buf ( n7341 , n7340 );
buf ( n7342 , n7341 );
not ( n7343 , n7342 );
buf ( n7344 , n7343 );
buf ( n7345 , n7344 );
and ( n7346 , n7338 , n7345 );
nor ( n7347 , n7337 , n7346 );
buf ( n7348 , n7347 );
or ( n7349 , n7348 , n6451 );
nand ( n7350 , n7317 , n7349 );
buf ( n7351 , n7350 );
and ( n7352 , n7268 , n7351 );
and ( n7353 , n7232 , n7267 );
or ( n7354 , n7352 , n7353 );
buf ( n7355 , n7354 );
buf ( n7356 , n7355 );
and ( n7357 , n7065 , n7356 );
not ( n7358 , n7065 );
buf ( n7359 , n7355 );
not ( n7360 , n7359 );
buf ( n7361 , n7360 );
buf ( n7362 , n7361 );
and ( n7363 , n7358 , n7362 );
nor ( n7364 , n7357 , n7363 );
buf ( n7365 , n7364 );
not ( n7366 , n7260 );
and ( n7367 , n413 , n7306 );
not ( n7368 , n413 );
and ( n7369 , n7368 , n7295 );
or ( n7370 , n7367 , n7369 );
not ( n7371 , n7370 );
or ( n7372 , n7366 , n7371 );
buf ( n7373 , n7258 );
buf ( n7374 , n6520 );
nand ( n7375 , n7373 , n7374 );
buf ( n7376 , n7375 );
nand ( n7377 , n7372 , n7376 );
buf ( n7378 , n7377 );
buf ( n7379 , n7013 );
not ( n7380 , n7379 );
buf ( n7381 , n7054 );
not ( n7382 , n7381 );
or ( n7383 , n7380 , n7382 );
and ( n7384 , n411 , n6852 );
not ( n7385 , n411 );
and ( n7386 , n7385 , n6855 );
or ( n7387 , n7384 , n7386 );
buf ( n7388 , n7387 );
buf ( n7389 , n5837 );
nand ( n7390 , n7388 , n7389 );
buf ( n7391 , n7390 );
buf ( n7392 , n7391 );
nand ( n7393 , n7383 , n7392 );
buf ( n7394 , n7393 );
buf ( n7395 , n6528 );
not ( n7396 , n7395 );
buf ( n7397 , n6868 );
not ( n7398 , n7397 );
or ( n7399 , n7396 , n7398 );
buf ( n7400 , n6973 );
buf ( n7401 , n7400 );
buf ( n7402 , n7401 );
buf ( n7403 , n7402 );
buf ( n7404 , n6539 );
nand ( n7405 , n7403 , n7404 );
buf ( n7406 , n7405 );
buf ( n7407 , n7406 );
nand ( n7408 , n7399 , n7407 );
buf ( n7409 , n7408 );
or ( n7410 , n7394 , n7409 );
and ( n7411 , n6879 , n6949 );
not ( n7412 , n6879 );
and ( n7413 , n7412 , n7004 );
nor ( n7414 , n7411 , n7413 );
buf ( n7415 , n7414 );
not ( n7416 , n6999 );
and ( n7417 , n7415 , n7416 );
not ( n7418 , n7415 );
and ( n7419 , n7418 , n6999 );
nor ( n7420 , n7417 , n7419 );
nand ( n7421 , n7410 , n7420 );
nand ( n7422 , n7394 , n7409 );
nand ( n7423 , n7421 , n7422 );
buf ( n7424 , n7423 );
xor ( n7425 , n7378 , n7424 );
not ( n7426 , n416 );
not ( n7427 , n6410 );
nor ( n7428 , n7427 , n6175 );
not ( n7429 , n7428 );
buf ( n7430 , n6397 );
buf ( n7431 , n6217 );
nand ( n7432 , n7430 , n7431 );
buf ( n7433 , n7432 );
buf ( n7434 , n7319 );
buf ( n7435 , n6116 );
buf ( n7436 , n6217 );
nand ( n7437 , n7434 , n7435 , n7436 );
buf ( n7438 , n7437 );
nand ( n7439 , n7433 , n7438 , n6403 );
not ( n7440 , n7439 );
not ( n7441 , n7440 );
or ( n7442 , n7429 , n7441 );
not ( n7443 , n7428 );
nand ( n7444 , n7439 , n7443 );
nand ( n7445 , n7442 , n7444 );
xor ( n7446 , n415 , n7445 );
not ( n7447 , n7446 );
or ( n7448 , n7426 , n7447 );
not ( n7449 , n7348 );
nand ( n7450 , n7449 , n6455 );
nand ( n7451 , n7448 , n7450 );
buf ( n7452 , n7451 );
xnor ( n7453 , n7425 , n7452 );
buf ( n7454 , n7453 );
xor ( n7455 , n7365 , n7454 );
buf ( n7456 , n7455 );
xor ( n7457 , n7232 , n7267 );
xor ( n7458 , n7457 , n7351 );
buf ( n7459 , n7458 );
buf ( n7460 , n7459 );
not ( n7461 , n7460 );
buf ( n7462 , n7461 );
not ( n7463 , n7462 );
buf ( n7464 , n7414 );
buf ( n7465 , n7409 );
xor ( n7466 , n7464 , n7465 );
buf ( n7467 , n6999 );
xor ( n7468 , n7466 , n7467 );
buf ( n7469 , n7468 );
buf ( n7470 , n7469 );
buf ( n7471 , n7394 );
not ( n7472 , n7471 );
buf ( n7473 , n7472 );
buf ( n7474 , n7473 );
and ( n7475 , n7470 , n7474 );
not ( n7476 , n7470 );
buf ( n7477 , n7394 );
and ( n7478 , n7476 , n7477 );
nor ( n7479 , n7475 , n7478 );
buf ( n7480 , n7479 );
buf ( n7481 , n7480 );
not ( n7482 , n7481 );
buf ( n7483 , n7482 );
not ( n7484 , n7483 );
and ( n7485 , n7463 , n7484 );
buf ( n7486 , n7462 );
buf ( n7487 , n7483 );
nand ( n7488 , n7486 , n7487 );
buf ( n7489 , n7488 );
buf ( n7490 , n7013 );
not ( n7491 , n7490 );
buf ( n7492 , n7387 );
not ( n7493 , n7492 );
or ( n7494 , n7491 , n7493 );
buf ( n7495 , n6868 );
not ( n7496 , n7495 );
buf ( n7497 , n7496 );
and ( n7498 , n411 , n7497 );
not ( n7499 , n411 );
and ( n7500 , n7499 , n6868 );
or ( n7501 , n7498 , n7500 );
buf ( n7502 , n7501 );
buf ( n7503 , n5837 );
nand ( n7504 , n7502 , n7503 );
buf ( n7505 , n7504 );
buf ( n7506 , n7505 );
nand ( n7507 , n7494 , n7506 );
buf ( n7508 , n7507 );
buf ( n7509 , n7508 );
xor ( n7510 , n7134 , n7219 );
xor ( n7511 , n7510 , n7227 );
buf ( n7512 , n7511 );
buf ( n7513 , n7512 );
xor ( n7514 , n7509 , n7513 );
buf ( n7515 , n7260 );
not ( n7516 , n7515 );
buf ( n7517 , n7235 );
not ( n7518 , n7517 );
or ( n7519 , n7516 , n7518 );
buf ( n7520 , n413 );
not ( n7521 , n7520 );
buf ( n7522 , n7050 );
not ( n7523 , n7522 );
or ( n7524 , n7521 , n7523 );
buf ( n7525 , n7044 );
buf ( n7526 , n6496 );
nand ( n7527 , n7525 , n7526 );
buf ( n7528 , n7527 );
buf ( n7529 , n7528 );
nand ( n7530 , n7524 , n7529 );
buf ( n7531 , n7530 );
buf ( n7532 , n7531 );
buf ( n7533 , n6520 );
nand ( n7534 , n7532 , n7533 );
buf ( n7535 , n7534 );
buf ( n7536 , n7535 );
nand ( n7537 , n7519 , n7536 );
buf ( n7538 , n7537 );
buf ( n7539 , n7538 );
and ( n7540 , n7514 , n7539 );
and ( n7541 , n7509 , n7513 );
or ( n7542 , n7540 , n7541 );
buf ( n7543 , n7542 );
and ( n7544 , n7489 , n7543 );
nor ( n7545 , n7485 , n7544 );
buf ( n7546 , n7545 );
nand ( n7547 , n7456 , n7546 );
buf ( n7548 , n7547 );
buf ( n7549 , n7548 );
buf ( n7550 , n7549 );
buf ( n7551 , n7550 );
buf ( n7552 , n7551 );
not ( n7553 , n7552 );
xor ( n7554 , n7201 , n7177 );
xor ( n7555 , n7554 , n7207 );
buf ( n7556 , n7555 );
buf ( n7557 , n7013 );
not ( n7558 , n7557 );
buf ( n7559 , n7501 );
not ( n7560 , n7559 );
or ( n7561 , n7558 , n7560 );
buf ( n7562 , n7402 );
not ( n7563 , n7562 );
buf ( n7564 , n7563 );
and ( n7565 , n411 , n7564 );
not ( n7566 , n411 );
and ( n7567 , n7566 , n7402 );
or ( n7568 , n7565 , n7567 );
buf ( n7569 , n7568 );
buf ( n7570 , n5837 );
nand ( n7571 , n7569 , n7570 );
buf ( n7572 , n7571 );
buf ( n7573 , n7572 );
nand ( n7574 , n7561 , n7573 );
buf ( n7575 , n7574 );
buf ( n7576 , n7575 );
xor ( n7577 , n7556 , n7576 );
buf ( n7578 , n7260 );
not ( n7579 , n7578 );
buf ( n7580 , n7531 );
not ( n7581 , n7580 );
or ( n7582 , n7579 , n7581 );
buf ( n7583 , n413 );
not ( n7584 , n7583 );
buf ( n7585 , n6852 );
not ( n7586 , n7585 );
or ( n7587 , n7584 , n7586 );
nand ( n7588 , n6855 , n6496 );
buf ( n7589 , n7588 );
nand ( n7590 , n7587 , n7589 );
buf ( n7591 , n7590 );
buf ( n7592 , n7591 );
buf ( n7593 , n6520 );
nand ( n7594 , n7592 , n7593 );
buf ( n7595 , n7594 );
buf ( n7596 , n7595 );
nand ( n7597 , n7582 , n7596 );
buf ( n7598 , n7597 );
buf ( n7599 , n7598 );
and ( n7600 , n7577 , n7599 );
and ( n7601 , n7556 , n7576 );
or ( n7602 , n7600 , n7601 );
buf ( n7603 , n7602 );
buf ( n7604 , n7603 );
not ( n7605 , n7604 );
buf ( n7606 , n416 );
not ( n7607 , n7606 );
buf ( n7608 , n7314 );
not ( n7609 , n7608 );
or ( n7610 , n7607 , n7609 );
buf ( n7611 , n415 );
buf ( n7612 , n7250 );
and ( n7613 , n7611 , n7612 );
not ( n7614 , n7611 );
buf ( n7615 , n7250 );
not ( n7616 , n7615 );
buf ( n7617 , n7616 );
buf ( n7618 , n7617 );
and ( n7619 , n7614 , n7618 );
nor ( n7620 , n7613 , n7619 );
buf ( n7621 , n7620 );
buf ( n7622 , n7621 );
buf ( n7623 , n6455 );
nand ( n7624 , n7622 , n7623 );
buf ( n7625 , n7624 );
buf ( n7626 , n7625 );
nand ( n7627 , n7610 , n7626 );
buf ( n7628 , n7627 );
buf ( n7629 , n7628 );
not ( n7630 , n7629 );
buf ( n7631 , n7630 );
buf ( n7632 , n7631 );
nand ( n7633 , n7605 , n7632 );
buf ( n7634 , n7633 );
buf ( n7635 , n7634 );
not ( n7636 , n7635 );
xor ( n7637 , n7509 , n7513 );
xor ( n7638 , n7637 , n7539 );
buf ( n7639 , n7638 );
buf ( n7640 , n7639 );
not ( n7641 , n7640 );
or ( n7642 , n7636 , n7641 );
buf ( n7643 , n7631 );
not ( n7644 , n7643 );
buf ( n7645 , n7603 );
nand ( n7646 , n7644 , n7645 );
buf ( n7647 , n7646 );
buf ( n7648 , n7647 );
nand ( n7649 , n7642 , n7648 );
buf ( n7650 , n7649 );
buf ( n7651 , n7650 );
not ( n7652 , n7651 );
buf ( n7653 , n7480 );
buf ( n7654 , n7543 );
xor ( n7655 , n7653 , n7654 );
buf ( n7656 , n7459 );
xnor ( n7657 , n7655 , n7656 );
buf ( n7658 , n7657 );
buf ( n7659 , n7658 );
nand ( n7660 , n7652 , n7659 );
buf ( n7661 , n7660 );
buf ( n7662 , n7661 );
buf ( n7663 , n416 );
not ( n7664 , n7663 );
buf ( n7665 , n415 );
not ( n7666 , n7665 );
buf ( n7667 , n7034 );
not ( n7668 , n7667 );
or ( n7669 , n7666 , n7668 );
buf ( n7670 , n6467 );
buf ( n7671 , n7031 );
nand ( n7672 , n7670 , n7671 );
buf ( n7673 , n7672 );
buf ( n7674 , n7673 );
nand ( n7675 , n7669 , n7674 );
buf ( n7676 , n7675 );
buf ( n7677 , n7676 );
not ( n7678 , n7677 );
or ( n7679 , n7664 , n7678 );
buf ( n7680 , n415 );
buf ( n7681 , n7044 );
and ( n7682 , n7680 , n7681 );
not ( n7683 , n7680 );
buf ( n7684 , n7050 );
and ( n7685 , n7683 , n7684 );
nor ( n7686 , n7682 , n7685 );
buf ( n7687 , n7686 );
buf ( n7688 , n7687 );
buf ( n7689 , n6455 );
nand ( n7690 , n7688 , n7689 );
buf ( n7691 , n7690 );
buf ( n7692 , n7691 );
nand ( n7693 , n7679 , n7692 );
buf ( n7694 , n7693 );
buf ( n7695 , n7694 );
xor ( n7696 , n6868 , n6496 );
not ( n7697 , n7696 );
not ( n7698 , n6523 );
and ( n7699 , n7697 , n7698 );
and ( n7700 , n7591 , n7260 );
nor ( n7701 , n7699 , n7700 );
buf ( n7702 , n7701 );
not ( n7703 , n7702 );
buf ( n7704 , n7703 );
buf ( n7705 , n7704 );
nor ( n7706 , n7695 , n7705 );
buf ( n7707 , n7706 );
buf ( n7708 , n7707 );
buf ( n7709 , n7174 );
not ( n7710 , n7709 );
buf ( n7711 , n7155 );
buf ( n7712 , n7167 );
not ( n7713 , n7712 );
xor ( n7714 , n7711 , n7713 );
buf ( n7715 , n7714 );
buf ( n7716 , n7715 );
not ( n7717 , n7716 );
or ( n7718 , n7710 , n7717 );
buf ( n7719 , n7715 );
buf ( n7720 , n7174 );
or ( n7721 , n7719 , n7720 );
nand ( n7722 , n7718 , n7721 );
buf ( n7723 , n7722 );
not ( n7724 , n7723 );
buf ( n7725 , n7402 );
buf ( n7726 , n7013 );
nand ( n7727 , n7725 , n7726 );
buf ( n7728 , n7727 );
not ( n7729 , n7728 );
and ( n7730 , n7724 , n7729 );
and ( n7731 , n7723 , n7728 );
nor ( n7732 , n7730 , n7731 );
buf ( n7733 , n7145 );
buf ( n7734 , n7150 );
buf ( n7735 , n7090 );
and ( n7736 , n7734 , n7735 );
not ( n7737 , n7734 );
buf ( n7738 , n7087 );
and ( n7739 , n7737 , n7738 );
nor ( n7740 , n7736 , n7739 );
buf ( n7741 , n7740 );
buf ( n7742 , n7741 );
xnor ( n7743 , n7733 , n7742 );
buf ( n7744 , n7743 );
not ( n7745 , n7744 );
buf ( n7746 , n375 );
buf ( n7747 , n385 );
and ( n7748 , n7746 , n7747 );
buf ( n7749 , n376 );
buf ( n7750 , n384 );
and ( n7751 , n7749 , n7750 );
nor ( n7752 , n7748 , n7751 );
buf ( n7753 , n7752 );
buf ( n7754 , n7753 );
not ( n7755 , n7754 );
buf ( n7756 , n7150 );
nand ( n7757 , n7755 , n7756 );
buf ( n7758 , n7757 );
buf ( n7759 , n7758 );
buf ( n7760 , n377 );
buf ( n7761 , n383 );
nand ( n7762 , n7760 , n7761 );
buf ( n7763 , n7762 );
buf ( n7764 , n7763 );
buf ( n7765 , n6920 );
or ( n7766 , n7764 , n7765 );
buf ( n7767 , n7766 );
buf ( n7768 , n7767 );
and ( n7769 , n7759 , n7768 );
buf ( n7770 , n7763 );
buf ( n7771 , n6920 );
and ( n7772 , n7770 , n7771 );
nor ( n7773 , n7769 , n7772 );
buf ( n7774 , n7773 );
not ( n7775 , n7774 );
nand ( n7776 , n7745 , n7775 );
not ( n7777 , n7776 );
buf ( n7778 , n6518 );
not ( n7779 , n7778 );
buf ( n7780 , n6973 );
not ( n7781 , n7780 );
or ( n7782 , n7779 , n7781 );
buf ( n7783 , n414 );
buf ( n7784 , n415 );
and ( n7785 , n7783 , n7784 );
buf ( n7786 , n6496 );
nor ( n7787 , n7785 , n7786 );
buf ( n7788 , n7787 );
buf ( n7789 , n7788 );
nand ( n7790 , n7782 , n7789 );
buf ( n7791 , n7790 );
not ( n7792 , n7791 );
or ( n7793 , n7777 , n7792 );
nand ( n7794 , n7744 , n7774 );
nand ( n7795 , n7793 , n7794 );
and ( n7796 , n7732 , n7795 );
not ( n7797 , n7732 );
not ( n7798 , n7795 );
and ( n7799 , n7797 , n7798 );
nor ( n7800 , n7796 , n7799 );
not ( n7801 , n7800 );
buf ( n7802 , n7801 );
or ( n7803 , n7708 , n7802 );
buf ( n7804 , n7694 );
buf ( n7805 , n7704 );
nand ( n7806 , n7804 , n7805 );
buf ( n7807 , n7806 );
buf ( n7808 , n7807 );
nand ( n7809 , n7803 , n7808 );
buf ( n7810 , n7809 );
not ( n7811 , n7810 );
buf ( n7812 , n7723 );
not ( n7813 , n7812 );
buf ( n7814 , n7728 );
nand ( n7815 , n7813 , n7814 );
buf ( n7816 , n7815 );
buf ( n7817 , n7816 );
not ( n7818 , n7817 );
buf ( n7819 , n7798 );
not ( n7820 , n7819 );
or ( n7821 , n7818 , n7820 );
buf ( n7822 , n7728 );
not ( n7823 , n7822 );
buf ( n7824 , n7723 );
nand ( n7825 , n7823 , n7824 );
buf ( n7826 , n7825 );
buf ( n7827 , n7826 );
nand ( n7828 , n7821 , n7827 );
buf ( n7829 , n7828 );
buf ( n7830 , n7829 );
buf ( n7831 , n6455 );
not ( n7832 , n7831 );
buf ( n7833 , n7676 );
not ( n7834 , n7833 );
or ( n7835 , n7832 , n7834 );
buf ( n7836 , n7621 );
buf ( n7837 , n416 );
nand ( n7838 , n7836 , n7837 );
buf ( n7839 , n7838 );
buf ( n7840 , n7839 );
nand ( n7841 , n7835 , n7840 );
buf ( n7842 , n7841 );
buf ( n7843 , n7842 );
xor ( n7844 , n7830 , n7843 );
xor ( n7845 , n7556 , n7576 );
xor ( n7846 , n7845 , n7599 );
buf ( n7847 , n7846 );
buf ( n7848 , n7847 );
xnor ( n7849 , n7844 , n7848 );
buf ( n7850 , n7849 );
nand ( n7851 , n7811 , n7850 );
not ( n7852 , n7851 );
buf ( n7853 , n413 );
not ( n7854 , n7853 );
buf ( n7855 , n7564 );
not ( n7856 , n7855 );
or ( n7857 , n7854 , n7856 );
buf ( n7858 , n7402 );
buf ( n7859 , n6496 );
nand ( n7860 , n7858 , n7859 );
buf ( n7861 , n7860 );
buf ( n7862 , n7861 );
nand ( n7863 , n7857 , n7862 );
buf ( n7864 , n7863 );
not ( n7865 , n7864 );
not ( n7866 , n6520 );
or ( n7867 , n7865 , n7866 );
or ( n7868 , n7696 , n6519 );
nand ( n7869 , n7867 , n7868 );
buf ( n7870 , n7869 );
not ( n7871 , n7870 );
buf ( n7872 , n7871 );
buf ( n7873 , n7872 );
not ( n7874 , n7873 );
buf ( n7875 , n416 );
not ( n7876 , n7875 );
buf ( n7877 , n7687 );
not ( n7878 , n7877 );
or ( n7879 , n7876 , n7878 );
buf ( n7880 , n415 );
buf ( n7881 , n6855 );
and ( n7882 , n7880 , n7881 );
not ( n7883 , n7880 );
buf ( n7884 , n6852 );
and ( n7885 , n7883 , n7884 );
nor ( n7886 , n7882 , n7885 );
buf ( n7887 , n7886 );
buf ( n7888 , n7887 );
buf ( n7889 , n6455 );
nand ( n7890 , n7888 , n7889 );
buf ( n7891 , n7890 );
buf ( n7892 , n7891 );
nand ( n7893 , n7879 , n7892 );
buf ( n7894 , n7893 );
buf ( n7895 , n7894 );
not ( n7896 , n7895 );
buf ( n7897 , n7896 );
buf ( n7898 , n7897 );
not ( n7899 , n7898 );
or ( n7900 , n7874 , n7899 );
not ( n7901 , n7791 );
not ( n7902 , n7775 );
not ( n7903 , n7744 );
or ( n7904 , n7902 , n7903 );
nand ( n7905 , n7745 , n7774 );
nand ( n7906 , n7904 , n7905 );
and ( n7907 , n7901 , n7906 );
not ( n7908 , n7901 );
not ( n7909 , n7906 );
and ( n7910 , n7908 , n7909 );
nor ( n7911 , n7907 , n7910 );
buf ( n7912 , n7911 );
nand ( n7913 , n7900 , n7912 );
buf ( n7914 , n7913 );
buf ( n7915 , n7914 );
buf ( n7916 , n7897 );
not ( n7917 , n7916 );
buf ( n7918 , n7869 );
nand ( n7919 , n7917 , n7918 );
buf ( n7920 , n7919 );
buf ( n7921 , n7920 );
nand ( n7922 , n7915 , n7921 );
buf ( n7923 , n7922 );
buf ( n7924 , n7923 );
not ( n7925 , n7924 );
buf ( n7926 , n7694 );
not ( n7927 , n7926 );
not ( n7928 , n7701 );
not ( n7929 , n7801 );
or ( n7930 , n7928 , n7929 );
or ( n7931 , n7801 , n7701 );
nand ( n7932 , n7930 , n7931 );
buf ( n7933 , n7932 );
not ( n7934 , n7933 );
and ( n7935 , n7927 , n7934 );
buf ( n7936 , n7694 );
buf ( n7937 , n7932 );
and ( n7938 , n7936 , n7937 );
nor ( n7939 , n7935 , n7938 );
buf ( n7940 , n7939 );
buf ( n7941 , n7940 );
nand ( n7942 , n7925 , n7941 );
buf ( n7943 , n7942 );
not ( n7944 , n7943 );
xor ( n7945 , n7911 , n7869 );
xnor ( n7946 , n7945 , n7897 );
buf ( n7947 , n7946 );
buf ( n7948 , n377 );
buf ( n7949 , n384 );
nand ( n7950 , n7948 , n7949 );
buf ( n7951 , n7950 );
buf ( n7952 , n7951 );
not ( n7953 , n7952 );
buf ( n7954 , n6920 );
nand ( n7955 , n7953 , n7954 );
buf ( n7956 , n7955 );
buf ( n7957 , n7956 );
not ( n7958 , n7957 );
buf ( n7959 , n7402 );
buf ( n7960 , n416 );
nand ( n7961 , n7959 , n7960 );
buf ( n7962 , n7961 );
buf ( n7963 , n7962 );
buf ( n7964 , n415 );
nand ( n7965 , n7963 , n7964 );
buf ( n7966 , n7965 );
buf ( n7967 , n7966 );
not ( n7968 , n7967 );
buf ( n7969 , n7968 );
buf ( n7970 , n7969 );
not ( n7971 , n7970 );
or ( n7972 , n7958 , n7971 );
buf ( n7973 , n6923 );
buf ( n7974 , n7951 );
nand ( n7975 , n7973 , n7974 );
buf ( n7976 , n7975 );
buf ( n7977 , n7976 );
nand ( n7978 , n7972 , n7977 );
buf ( n7979 , n7978 );
not ( n7980 , n7979 );
buf ( n7981 , n7402 );
buf ( n7982 , n7260 );
nand ( n7983 , n7981 , n7982 );
buf ( n7984 , n7983 );
or ( n7985 , n7980 , n7984 );
buf ( n7986 , n7984 );
not ( n7987 , n7986 );
buf ( n7988 , n7980 );
not ( n7989 , n7988 );
or ( n7990 , n7987 , n7989 );
buf ( n7991 , n7763 );
buf ( n7992 , n6920 );
and ( n7993 , n7991 , n7992 );
not ( n7994 , n7991 );
buf ( n7995 , n6923 );
and ( n7996 , n7994 , n7995 );
nor ( n7997 , n7993 , n7996 );
buf ( n7998 , n7997 );
buf ( n7999 , n7998 );
not ( n8000 , n7999 );
buf ( n8001 , n7758 );
not ( n8002 , n8001 );
buf ( n8003 , n8002 );
buf ( n8004 , n8003 );
not ( n8005 , n8004 );
or ( n8006 , n8000 , n8005 );
buf ( n8007 , n8003 );
buf ( n8008 , n7998 );
or ( n8009 , n8007 , n8008 );
nand ( n8010 , n8006 , n8009 );
buf ( n8011 , n8010 );
buf ( n8012 , n8011 );
nand ( n8013 , n7990 , n8012 );
buf ( n8014 , n8013 );
nand ( n8015 , n7985 , n8014 );
buf ( n8016 , n8015 );
nor ( n8017 , n7947 , n8016 );
buf ( n8018 , n8017 );
buf ( n8019 , n8018 );
xor ( n8020 , n8011 , n7984 );
and ( n8021 , n8020 , n7979 );
not ( n8022 , n8020 );
and ( n8023 , n8022 , n7980 );
nor ( n8024 , n8021 , n8023 );
buf ( n8025 , n7887 );
buf ( n8026 , n416 );
nand ( n8027 , n8025 , n8026 );
buf ( n8028 , n8027 );
buf ( n8029 , n415 );
not ( n8030 , n8029 );
buf ( n8031 , n7497 );
not ( n8032 , n8031 );
or ( n8033 , n8030 , n8032 );
buf ( n8034 , n6868 );
buf ( n8035 , n6467 );
nand ( n8036 , n8034 , n8035 );
buf ( n8037 , n8036 );
buf ( n8038 , n8037 );
nand ( n8039 , n8033 , n8038 );
buf ( n8040 , n8039 );
buf ( n8041 , n8040 );
buf ( n8042 , n6455 );
nand ( n8043 , n8041 , n8042 );
buf ( n8044 , n8043 );
nand ( n8045 , n8024 , n8028 , n8044 );
buf ( n8046 , n416 );
not ( n8047 , n8046 );
buf ( n8048 , n8040 );
not ( n8049 , n8048 );
or ( n8050 , n8047 , n8049 );
buf ( n8051 , n7564 );
buf ( n8052 , n6455 );
nand ( n8053 , n8051 , n8052 );
buf ( n8054 , n8053 );
buf ( n8055 , n8054 );
nand ( n8056 , n8050 , n8055 );
buf ( n8057 , n8056 );
buf ( n8058 , n8057 );
buf ( n8059 , n7951 );
not ( n8060 , n8059 );
buf ( n8061 , n6920 );
not ( n8062 , n8061 );
and ( n8063 , n8060 , n8062 );
buf ( n8064 , n7951 );
buf ( n8065 , n6920 );
and ( n8066 , n8064 , n8065 );
nor ( n8067 , n8063 , n8066 );
buf ( n8068 , n8067 );
buf ( n8069 , n8068 );
not ( n8070 , n8069 );
buf ( n8071 , n7969 );
not ( n8072 , n8071 );
or ( n8073 , n8070 , n8072 );
buf ( n8074 , n7969 );
buf ( n8075 , n8068 );
or ( n8076 , n8074 , n8075 );
nand ( n8077 , n8073 , n8076 );
buf ( n8078 , n8077 );
buf ( n8079 , n8078 );
nor ( n8080 , n8058 , n8079 );
buf ( n8081 , n8080 );
buf ( n8082 , n8081 );
buf ( n8083 , n7962 );
buf ( n8084 , n377 );
buf ( n8085 , n385 );
and ( n8086 , n8084 , n8085 );
buf ( n8087 , n8086 );
buf ( n8088 , n8087 );
nand ( n8089 , n8083 , n8088 );
buf ( n8090 , n8089 );
buf ( n8091 , n8090 );
not ( n8092 , n8091 );
buf ( n8093 , n8092 );
buf ( n8094 , n8093 );
or ( n8095 , n8082 , n8094 );
buf ( n8096 , n8057 );
buf ( n8097 , n8078 );
nand ( n8098 , n8096 , n8097 );
buf ( n8099 , n8098 );
buf ( n8100 , n8099 );
nand ( n8101 , n8095 , n8100 );
buf ( n8102 , n8101 );
and ( n8103 , n8045 , n8102 );
buf ( n8104 , n8024 );
not ( n8105 , n8104 );
buf ( n8106 , n8105 );
and ( n8107 , n7887 , n416 );
and ( n8108 , n8040 , n6455 );
nor ( n8109 , n8107 , n8108 );
buf ( n8110 , n8109 );
not ( n8111 , n8110 );
buf ( n8112 , n8111 );
and ( n8113 , n8106 , n8112 );
nor ( n8114 , n8103 , n8113 );
buf ( n8115 , n8114 );
or ( n8116 , n8019 , n8115 );
buf ( n8117 , n7946 );
buf ( n8118 , n8015 );
nand ( n8119 , n8117 , n8118 );
buf ( n8120 , n8119 );
buf ( n8121 , n8120 );
nand ( n8122 , n8116 , n8121 );
buf ( n8123 , n8122 );
not ( n8124 , n8123 );
or ( n8125 , n7944 , n8124 );
not ( n8126 , n7940 );
nand ( n8127 , n8126 , n7923 );
nand ( n8128 , n8125 , n8127 );
not ( n8129 , n8128 );
or ( n8130 , n7852 , n8129 );
not ( n8131 , n7850 );
buf ( n8132 , n7707 );
buf ( n8133 , n7801 );
or ( n8134 , n8132 , n8133 );
buf ( n8135 , n7807 );
nand ( n8136 , n8134 , n8135 );
buf ( n8137 , n8136 );
nand ( n8138 , n8131 , n8137 );
nand ( n8139 , n8130 , n8138 );
buf ( n8140 , n8139 );
not ( n8141 , n7829 );
buf ( n8142 , n6455 );
not ( n8143 , n8142 );
buf ( n8144 , n7676 );
not ( n8145 , n8144 );
or ( n8146 , n8143 , n8145 );
buf ( n8147 , n7839 );
nand ( n8148 , n8146 , n8147 );
buf ( n8149 , n8148 );
not ( n8150 , n8149 );
nand ( n8151 , n8141 , n8150 );
not ( n8152 , n8151 );
not ( n8153 , n7847 );
or ( n8154 , n8152 , n8153 );
not ( n8155 , n8150 );
nand ( n8156 , n8155 , n7829 );
nand ( n8157 , n8154 , n8156 );
buf ( n8158 , n8157 );
not ( n8159 , n8158 );
not ( n8160 , n7631 );
and ( n8161 , n7603 , n8160 );
not ( n8162 , n7603 );
and ( n8163 , n8162 , n7631 );
nor ( n8164 , n8161 , n8163 );
not ( n8165 , n7639 );
and ( n8166 , n8164 , n8165 );
not ( n8167 , n8164 );
and ( n8168 , n8167 , n7639 );
nor ( n8169 , n8166 , n8168 );
buf ( n8170 , n8169 );
nand ( n8171 , n8159 , n8170 );
buf ( n8172 , n8171 );
buf ( n8173 , n8172 );
nand ( n8174 , n8140 , n8173 );
buf ( n8175 , n8174 );
buf ( n8176 , n8175 );
not ( n8177 , n8169 );
nand ( n8178 , n8177 , n8157 );
buf ( n8179 , n8178 );
nand ( n8180 , n8176 , n8179 );
buf ( n8181 , n8180 );
buf ( n8182 , n8181 );
and ( n8183 , n7662 , n8182 );
buf ( n8184 , n8183 );
buf ( n8185 , n8184 );
not ( n8186 , n8185 );
or ( n8187 , n7553 , n8186 );
not ( n8188 , n7548 );
buf ( n8189 , n7650 );
not ( n8190 , n8189 );
buf ( n8191 , n7658 );
nor ( n8192 , n8190 , n8191 );
buf ( n8193 , n8192 );
not ( n8194 , n8193 );
or ( n8195 , n8188 , n8194 );
buf ( n8196 , n7455 );
not ( n8197 , n8196 );
buf ( n8198 , n8197 );
buf ( n8199 , n8198 );
buf ( n8200 , n7545 );
not ( n8201 , n8200 );
buf ( n8202 , n8201 );
buf ( n8203 , n8202 );
nand ( n8204 , n8199 , n8203 );
buf ( n8205 , n8204 );
nand ( n8206 , n8195 , n8205 );
buf ( n8207 , n8206 );
not ( n8208 , n8207 );
buf ( n8209 , n8208 );
buf ( n8210 , n8209 );
nand ( n8211 , n8187 , n8210 );
buf ( n8212 , n8211 );
not ( n8213 , n8212 );
not ( n8214 , n6520 );
not ( n8215 , n413 );
not ( n8216 , n7341 );
or ( n8217 , n8215 , n8216 );
buf ( n8218 , n6496 );
buf ( n8219 , n7332 );
nand ( n8220 , n8218 , n8219 );
buf ( n8221 , n8220 );
nand ( n8222 , n8217 , n8221 );
not ( n8223 , n8222 );
or ( n8224 , n8214 , n8223 );
xnor ( n8225 , n7428 , n413 );
and ( n8226 , n8225 , n7439 );
not ( n8227 , n8225 );
and ( n8228 , n8227 , n7440 );
or ( n8229 , n8226 , n8228 );
nand ( n8230 , n8229 , n7260 );
nand ( n8231 , n8224 , n8230 );
not ( n8232 , n8231 );
xor ( n8233 , n6752 , n6775 );
and ( n8234 , n8233 , n6826 );
and ( n8235 , n6752 , n6775 );
or ( n8236 , n8234 , n8235 );
not ( n8237 , n8236 );
nand ( n8238 , n381 , n372 );
not ( n8239 , n8238 );
nand ( n8240 , n373 , n380 );
nand ( n8241 , n383 , n370 );
nor ( n8242 , n8239 , n8240 , n8241 );
not ( n8243 , n8242 );
nand ( n8244 , n381 , n372 );
nand ( n8245 , n8240 , n8244 , n8241 );
not ( n8246 , n8241 );
nand ( n8247 , n8246 , n8239 , n8240 );
not ( n8248 , n8240 );
not ( n8249 , n8244 );
nand ( n8250 , n8248 , n8249 , n8241 );
nand ( n8251 , n8243 , n8245 , n8247 , n8250 );
not ( n8252 , n8251 );
not ( n8253 , n6813 );
not ( n8254 , n6759 );
nand ( n8255 , n374 , n380 );
not ( n8256 , n8255 );
or ( n8257 , n8254 , n8256 );
or ( n8258 , n8255 , n6707 );
nand ( n8259 , n8258 , n6761 );
nand ( n8260 , n8257 , n8259 );
and ( n8261 , n8253 , n8260 );
and ( n8262 , n8252 , n8261 );
not ( n8263 , n8252 );
nor ( n8264 , n6813 , n8260 );
and ( n8265 , n8263 , n8264 );
nor ( n8266 , n8262 , n8265 );
nand ( n8267 , n8251 , n8260 );
or ( n8268 , n8267 , n8253 );
not ( n8269 , n8260 );
nand ( n8270 , n8269 , n8252 , n6813 );
and ( n8271 , n8266 , n8268 , n8270 );
not ( n8272 , n6819 );
not ( n8273 , n6797 );
not ( n8274 , n8273 );
or ( n8275 , n8272 , n8274 );
nand ( n8276 , n8275 , n6824 );
not ( n8277 , n6819 );
nand ( n8278 , n8277 , n6797 );
nand ( n8279 , n8276 , n8278 );
xor ( n8280 , n8271 , n8279 );
buf ( n8281 , n6787 );
not ( n8282 , n8281 );
buf ( n8283 , n6783 );
nand ( n8284 , n8282 , n8283 );
buf ( n8285 , n8284 );
buf ( n8286 , n8285 );
not ( n8287 , n8286 );
buf ( n8288 , n6796 );
not ( n8289 , n8288 );
or ( n8290 , n8287 , n8289 );
buf ( n8291 , n6780 );
buf ( n8292 , n6787 );
nand ( n8293 , n8291 , n8292 );
buf ( n8294 , n8293 );
buf ( n8295 , n8294 );
nand ( n8296 , n8290 , n8295 );
buf ( n8297 , n8296 );
not ( n8298 , n8297 );
buf ( n8299 , n374 );
buf ( n8300 , n379 );
nand ( n8301 , n8299 , n8300 );
buf ( n8302 , n8301 );
buf ( n8303 , n375 );
buf ( n8304 , n378 );
nand ( n8305 , n8303 , n8304 );
buf ( n8306 , n8305 );
xor ( n8307 , n8302 , n8306 );
buf ( n8308 , n371 );
buf ( n8309 , n382 );
nand ( n8310 , n8308 , n8309 );
buf ( n8311 , n8310 );
xnor ( n8312 , n8307 , n8311 );
xor ( n8313 , n8298 , n8312 );
not ( n8314 , n6758 );
not ( n8315 , n6765 );
or ( n8316 , n8314 , n8315 );
nand ( n8317 , n8316 , n6766 );
xor ( n8318 , n8313 , n8317 );
xnor ( n8319 , n8280 , n8318 );
not ( n8320 , n8319 );
nand ( n8321 , n8237 , n8320 );
not ( n8322 , n8321 );
buf ( n8323 , n6528 );
not ( n8324 , n8323 );
buf ( n8325 , n7044 );
not ( n8326 , n8325 );
or ( n8327 , n8324 , n8326 );
buf ( n8328 , n6855 );
buf ( n8329 , n6539 );
nand ( n8330 , n8328 , n8329 );
buf ( n8331 , n8330 );
buf ( n8332 , n8331 );
nand ( n8333 , n8327 , n8332 );
buf ( n8334 , n8333 );
not ( n8335 , n8334 );
or ( n8336 , n8322 , n8335 );
nand ( n8337 , n8319 , n8236 );
nand ( n8338 , n8336 , n8337 );
not ( n8339 , n8338 );
not ( n8340 , n6528 );
not ( n8341 , n7031 );
or ( n8342 , n8340 , n8341 );
buf ( n8343 , n7044 );
buf ( n8344 , n6539 );
nand ( n8345 , n8343 , n8344 );
buf ( n8346 , n8345 );
nand ( n8347 , n8342 , n8346 );
not ( n8348 , n8347 );
not ( n8349 , n8348 );
and ( n8350 , n8339 , n8349 );
and ( n8351 , n8338 , n8348 );
nor ( n8352 , n8350 , n8351 );
not ( n8353 , n8352 );
or ( n8354 , n8232 , n8353 );
or ( n8355 , n8231 , n8352 );
nand ( n8356 , n8354 , n8355 );
not ( n8357 , n8356 );
xor ( n8358 , n8236 , n8320 );
xnor ( n8359 , n8358 , n8334 );
buf ( n8360 , n8359 );
buf ( n8361 , n6455 );
not ( n8362 , n8361 );
buf ( n8363 , n7446 );
not ( n8364 , n8363 );
or ( n8365 , n8362 , n8364 );
nand ( n8366 , n6131 , n6421 );
xor ( n8367 , n8366 , n415 );
not ( n8368 , n6218 );
nand ( n8369 , n6116 , n7319 , n8368 );
nand ( n8370 , n8368 , n6397 );
not ( n8371 , n6413 );
nand ( n8372 , n8369 , n8370 , n8371 );
xnor ( n8373 , n8367 , n8372 );
buf ( n8374 , n8373 );
buf ( n8375 , n416 );
nand ( n8376 , n8374 , n8375 );
buf ( n8377 , n8376 );
buf ( n8378 , n8377 );
nand ( n8379 , n8365 , n8378 );
buf ( n8380 , n8379 );
buf ( n8381 , n8380 );
or ( n8382 , n8360 , n8381 );
xor ( n8383 , n6877 , n7011 );
and ( n8384 , n8383 , n7062 );
and ( n8385 , n6877 , n7011 );
or ( n8386 , n8384 , n8385 );
buf ( n8387 , n8386 );
buf ( n8388 , n8387 );
nand ( n8389 , n8382 , n8388 );
buf ( n8390 , n8389 );
buf ( n8391 , n8390 );
buf ( n8392 , n8380 );
buf ( n8393 , n8359 );
nand ( n8394 , n8392 , n8393 );
buf ( n8395 , n8394 );
buf ( n8396 , n8395 );
nand ( n8397 , n8391 , n8396 );
buf ( n8398 , n8397 );
buf ( n8399 , n8398 );
not ( n8400 , n8399 );
buf ( n8401 , n8400 );
not ( n8402 , n8401 );
or ( n8403 , n8357 , n8402 );
not ( n8404 , n8356 );
nand ( n8405 , n8398 , n8404 );
nand ( n8406 , n8403 , n8405 );
buf ( n8407 , n416 );
not ( n8408 , n8407 );
buf ( n8409 , n415 );
not ( n8410 , n8409 );
buf ( n8411 , n418 );
not ( n8412 , n8411 );
buf ( n8413 , n6398 );
buf ( n8414 , n6381 );
buf ( n8415 , n6421 );
not ( n8416 , n8415 );
buf ( n8417 , n6414 );
nor ( n8418 , n8416 , n8417 );
buf ( n8419 , n8418 );
buf ( n8420 , n8419 );
nand ( n8421 , n8413 , n8414 , n8420 );
buf ( n8422 , n8421 );
buf ( n8423 , n8422 );
not ( n8424 , n8423 );
or ( n8425 , n8412 , n8424 );
buf ( n8426 , n6398 );
buf ( n8427 , n6427 );
buf ( n8428 , n6381 );
nand ( n8429 , n8426 , n8427 , n8428 );
buf ( n8430 , n8429 );
buf ( n8431 , n8430 );
nand ( n8432 , n8425 , n8431 );
buf ( n8433 , n8432 );
buf ( n8434 , n8433 );
not ( n8435 , n8434 );
buf ( n8436 , n8435 );
buf ( n8437 , n8436 );
not ( n8438 , n8437 );
or ( n8439 , n8410 , n8438 );
buf ( n8440 , n8433 );
buf ( n8441 , n6467 );
nand ( n8442 , n8440 , n8441 );
buf ( n8443 , n8442 );
buf ( n8444 , n8443 );
nand ( n8445 , n8439 , n8444 );
buf ( n8446 , n8445 );
buf ( n8447 , n8446 );
not ( n8448 , n8447 );
or ( n8449 , n8408 , n8448 );
buf ( n8450 , n8373 );
buf ( n8451 , n6455 );
nand ( n8452 , n8450 , n8451 );
buf ( n8453 , n8452 );
buf ( n8454 , n8453 );
nand ( n8455 , n8449 , n8454 );
buf ( n8456 , n8455 );
not ( n8457 , n8271 );
not ( n8458 , n8279 );
not ( n8459 , n8458 );
or ( n8460 , n8457 , n8459 );
nand ( n8461 , n8460 , n8318 );
or ( n8462 , n8458 , n8271 );
nand ( n8463 , n8461 , n8462 );
not ( n8464 , n8298 );
not ( n8465 , n8312 );
or ( n8466 , n8464 , n8465 );
nand ( n8467 , n8466 , n8317 );
not ( n8468 , n8312 );
nand ( n8469 , n8468 , n8297 );
nand ( n8470 , n8467 , n8469 );
buf ( n8471 , n8311 );
buf ( n8472 , n8302 );
or ( n8473 , n8471 , n8472 );
buf ( n8474 , n8306 );
nand ( n8475 , n8473 , n8474 );
buf ( n8476 , n8475 );
buf ( n8477 , n8476 );
buf ( n8478 , n8302 );
buf ( n8479 , n8311 );
nand ( n8480 , n8478 , n8479 );
buf ( n8481 , n8480 );
buf ( n8482 , n8481 );
nand ( n8483 , n8477 , n8482 );
buf ( n8484 , n8483 );
buf ( n8485 , n8484 );
nand ( n8486 , n370 , n382 );
buf ( n8487 , n8486 );
not ( n8488 , n8487 );
and ( n8489 , n373 , n379 );
buf ( n8490 , n8489 );
not ( n8491 , n8490 );
or ( n8492 , n8488 , n8491 );
buf ( n8493 , n8486 );
buf ( n8494 , n8489 );
or ( n8495 , n8493 , n8494 );
nand ( n8496 , n8492 , n8495 );
buf ( n8497 , n8496 );
buf ( n8498 , n8497 );
nand ( n8499 , n371 , n381 );
buf ( n8500 , n8499 );
xor ( n8501 , n8498 , n8500 );
buf ( n8502 , n8501 );
buf ( n8503 , n8502 );
xor ( n8504 , n8485 , n8503 );
buf ( n8505 , n372 );
buf ( n8506 , n380 );
nand ( n8507 , n8505 , n8506 );
buf ( n8508 , n8507 );
buf ( n8509 , n374 );
buf ( n8510 , n378 );
nand ( n8511 , n8509 , n8510 );
buf ( n8512 , n8511 );
xor ( n8513 , n8508 , n8512 );
or ( n8514 , n8238 , n8241 );
nand ( n8515 , n8514 , n8240 );
nand ( n8516 , n8244 , n8241 );
nand ( n8517 , n8515 , n8516 );
xor ( n8518 , n8513 , n8517 );
buf ( n8519 , n8518 );
xor ( n8520 , n8504 , n8519 );
buf ( n8521 , n8520 );
not ( n8522 , n8521 );
or ( n8523 , n8251 , n8260 );
nand ( n8524 , n8523 , n6813 );
nand ( n8525 , n8524 , n8267 );
or ( n8526 , n8470 , n8522 , n8525 );
nand ( n8527 , n8522 , n8525 );
or ( n8528 , n8527 , n8470 );
nand ( n8529 , n8526 , n8528 );
not ( n8530 , n8529 );
not ( n8531 , n8525 );
nand ( n8532 , n8531 , n8522 );
not ( n8533 , n8532 );
and ( n8534 , n8533 , n8470 );
and ( n8535 , n8521 , n8525 );
and ( n8536 , n8535 , n8470 );
nor ( n8537 , n8534 , n8536 );
nand ( n8538 , n8530 , n8537 );
xor ( n8539 , n8463 , n8538 );
not ( n8540 , n8539 );
not ( n8541 , n8540 );
buf ( n8542 , n411 );
buf ( n8543 , n7250 );
xor ( n8544 , n8542 , n8543 );
buf ( n8545 , n8544 );
not ( n8546 , n8545 );
not ( n8547 , n8546 );
not ( n8548 , n5840 );
and ( n8549 , n8547 , n8548 );
not ( n8550 , n411 );
not ( n8551 , n7306 );
or ( n8552 , n8550 , n8551 );
nand ( n8553 , n7295 , n7195 );
nand ( n8554 , n8552 , n8553 );
and ( n8555 , n8554 , n7013 );
nor ( n8556 , n8549 , n8555 );
not ( n8557 , n8556 );
not ( n8558 , n8557 );
or ( n8559 , n8541 , n8558 );
nand ( n8560 , n8556 , n8539 );
nand ( n8561 , n8559 , n8560 );
xor ( n8562 , n8456 , n8561 );
buf ( n8563 , n5837 );
not ( n8564 , n8563 );
buf ( n8565 , n7038 );
not ( n8566 , n8565 );
or ( n8567 , n8564 , n8566 );
buf ( n8568 , n8545 );
buf ( n8569 , n7013 );
nand ( n8570 , n8568 , n8569 );
buf ( n8571 , n8570 );
buf ( n8572 , n8571 );
nand ( n8573 , n8567 , n8572 );
buf ( n8574 , n8573 );
not ( n8575 , n8574 );
xor ( n8576 , n6748 , n6828 );
and ( n8577 , n8576 , n6874 );
and ( n8578 , n6748 , n6828 );
or ( n8579 , n8577 , n8578 );
buf ( n8580 , n8579 );
not ( n8581 , n8580 );
nand ( n8582 , n8575 , n8581 );
not ( n8583 , n8582 );
not ( n8584 , n7260 );
not ( n8585 , n8222 );
or ( n8586 , n8584 , n8585 );
nand ( n8587 , n7370 , n6520 );
nand ( n8588 , n8586 , n8587 );
not ( n8589 , n8588 );
or ( n8590 , n8583 , n8589 );
nand ( n8591 , n8580 , n8574 );
nand ( n8592 , n8590 , n8591 );
xor ( n8593 , n8562 , n8592 );
not ( n8594 , n8593 );
and ( n8595 , n8406 , n8594 );
not ( n8596 , n8406 );
and ( n8597 , n8596 , n8593 );
nor ( n8598 , n8595 , n8597 );
not ( n8599 , n7377 );
not ( n8600 , n7451 );
or ( n8601 , n8599 , n8600 );
not ( n8602 , n7422 );
not ( n8603 , n7421 );
or ( n8604 , n8602 , n8603 );
or ( n8605 , n7451 , n7377 );
nand ( n8606 , n8604 , n8605 );
nand ( n8607 , n8601 , n8606 );
not ( n8608 , n8607 );
xor ( n8609 , n8581 , n8574 );
xnor ( n8610 , n8609 , n8588 );
buf ( n8611 , n8610 );
not ( n8612 , n8611 );
or ( n8613 , n8608 , n8612 );
or ( n8614 , n8611 , n8607 );
xor ( n8615 , n8359 , n8380 );
xor ( n8616 , n8615 , n8387 );
nand ( n8617 , n8614 , n8616 );
nand ( n8618 , n8613 , n8617 );
not ( n8619 , n8618 );
nand ( n8620 , n8598 , n8619 );
buf ( n8621 , n8620 );
not ( n8622 , n8621 );
xor ( n8623 , n8610 , n8607 );
xnor ( n8624 , n8623 , n8616 );
not ( n8625 , n8624 );
buf ( n8626 , n7361 );
not ( n8627 , n8626 );
buf ( n8628 , n7064 );
nor ( n8629 , n8627 , n8628 );
buf ( n8630 , n8629 );
buf ( n8631 , n8630 );
buf ( n8632 , n7454 );
or ( n8633 , n8631 , n8632 );
buf ( n8634 , n7361 );
not ( n8635 , n8634 );
buf ( n8636 , n7064 );
nand ( n8637 , n8635 , n8636 );
buf ( n8638 , n8637 );
buf ( n8639 , n8638 );
nand ( n8640 , n8633 , n8639 );
buf ( n8641 , n8640 );
nor ( n8642 , n8625 , n8641 );
buf ( n8643 , n8642 );
nor ( n8644 , n8622 , n8643 );
buf ( n8645 , n8644 );
buf ( n8646 , n8645 );
not ( n8647 , n5837 );
not ( n8648 , n8554 );
or ( n8649 , n8647 , n8648 );
xor ( n8650 , n7327 , n411 );
xnor ( n8651 , n8650 , n7326 );
nand ( n8652 , n7013 , n8651 );
nand ( n8653 , n8649 , n8652 );
buf ( n8654 , n8653 );
buf ( n8655 , n6455 );
not ( n8656 , n8655 );
buf ( n8657 , n8446 );
not ( n8658 , n8657 );
or ( n8659 , n8656 , n8658 );
buf ( n8660 , n6477 );
buf ( n8661 , n8660 );
nand ( n8662 , n8659 , n8661 );
buf ( n8663 , n8662 );
buf ( n8664 , n8663 );
xor ( n8665 , n8654 , n8664 );
buf ( n8666 , n7260 );
not ( n8667 , n8666 );
not ( n8668 , n8366 );
not ( n8669 , n6496 );
and ( n8670 , n8668 , n8669 );
not ( n8671 , n8668 );
not ( n8672 , n413 );
and ( n8673 , n8671 , n8672 );
or ( n8674 , n8670 , n8673 );
and ( n8675 , n8372 , n8674 );
not ( n8676 , n8372 );
not ( n8677 , n6496 );
and ( n8678 , n8366 , n8677 );
not ( n8679 , n8366 );
not ( n8680 , n413 );
and ( n8681 , n8679 , n8680 );
or ( n8682 , n8678 , n8681 );
and ( n8683 , n8676 , n8682 );
or ( n8684 , n8675 , n8683 );
buf ( n8685 , n8684 );
not ( n8686 , n8685 );
or ( n8687 , n8667 , n8686 );
nand ( n8688 , n8229 , n6520 );
buf ( n8689 , n8688 );
nand ( n8690 , n8687 , n8689 );
buf ( n8691 , n8690 );
buf ( n8692 , n8691 );
not ( n8693 , n8692 );
buf ( n8694 , n8693 );
buf ( n8695 , n8694 );
xnor ( n8696 , n8665 , n8695 );
buf ( n8697 , n8696 );
buf ( n8698 , n8697 );
xor ( n8699 , n8456 , n8561 );
and ( n8700 , n8699 , n8592 );
and ( n8701 , n8456 , n8561 );
or ( n8702 , n8700 , n8701 );
buf ( n8703 , n8702 );
xor ( n8704 , n8698 , n8703 );
buf ( n8705 , n6539 );
not ( n8706 , n8705 );
buf ( n8707 , n7031 );
not ( n8708 , n8707 );
or ( n8709 , n8706 , n8708 );
buf ( n8710 , n7617 );
not ( n8711 , n8710 );
buf ( n8712 , n8711 );
buf ( n8713 , n8712 );
buf ( n8714 , n6528 );
nand ( n8715 , n8713 , n8714 );
buf ( n8716 , n8715 );
buf ( n8717 , n8716 );
nand ( n8718 , n8709 , n8717 );
buf ( n8719 , n8718 );
xor ( n8720 , n8508 , n8512 );
and ( n8721 , n8720 , n8517 );
and ( n8722 , n8508 , n8512 );
or ( n8723 , n8721 , n8722 );
nand ( n8724 , n371 , n380 );
nand ( n8725 , n370 , n382 );
not ( n8726 , n8725 );
not ( n8727 , n8499 );
or ( n8728 , n8726 , n8727 );
or ( n8729 , n8499 , n8725 );
nand ( n8730 , n8729 , n6811 );
nand ( n8731 , n8728 , n8730 );
xor ( n8732 , n8724 , n8731 );
nand ( n8733 , n372 , n379 );
nand ( n8734 , n373 , n378 );
xor ( n8735 , n8733 , n8734 );
nand ( n8736 , n370 , n381 );
xor ( n8737 , n8735 , n8736 );
xor ( n8738 , n8732 , n8737 );
buf ( n8739 , n8738 );
not ( n8740 , n8739 );
buf ( n8741 , n8740 );
and ( n8742 , n8723 , n8741 );
not ( n8743 , n8723 );
and ( n8744 , n8743 , n8738 );
or ( n8745 , n8742 , n8744 );
buf ( n8746 , n8745 );
xor ( n8747 , n8485 , n8503 );
and ( n8748 , n8747 , n8519 );
and ( n8749 , n8485 , n8503 );
or ( n8750 , n8748 , n8749 );
buf ( n8751 , n8750 );
buf ( n8752 , n8751 );
xnor ( n8753 , n8746 , n8752 );
buf ( n8754 , n8753 );
not ( n8755 , n8470 );
not ( n8756 , n8532 );
or ( n8757 , n8755 , n8756 );
not ( n8758 , n8535 );
nand ( n8759 , n8757 , n8758 );
xnor ( n8760 , n8754 , n8759 );
xnor ( n8761 , n8719 , n8760 );
buf ( n8762 , n8761 );
or ( n8763 , n8463 , n8538 );
not ( n8764 , n8763 );
not ( n8765 , n8557 );
or ( n8766 , n8764 , n8765 );
nand ( n8767 , n8463 , n8538 );
nand ( n8768 , n8766 , n8767 );
buf ( n8769 , n8768 );
xor ( n8770 , n8762 , n8769 );
or ( n8771 , n8347 , n8231 );
nand ( n8772 , n8771 , n8338 );
buf ( n8773 , n8772 );
nand ( n8774 , n8347 , n8231 );
buf ( n8775 , n8774 );
nand ( n8776 , n8773 , n8775 );
buf ( n8777 , n8776 );
buf ( n8778 , n8777 );
xnor ( n8779 , n8770 , n8778 );
buf ( n8780 , n8779 );
buf ( n8781 , n8780 );
xnor ( n8782 , n8704 , n8781 );
buf ( n8783 , n8782 );
buf ( n8784 , n8783 );
not ( n8785 , n8404 );
not ( n8786 , n8594 );
or ( n8787 , n8785 , n8786 );
buf ( n8788 , n8398 );
buf ( n8789 , n8788 );
buf ( n8790 , n8789 );
nand ( n8791 , n8787 , n8790 );
buf ( n8792 , n8791 );
nand ( n8793 , n8593 , n8356 );
buf ( n8794 , n8793 );
nand ( n8795 , n8792 , n8794 );
buf ( n8796 , n8795 );
not ( n8797 , n8796 );
buf ( n8798 , n8797 );
nand ( n8799 , n8784 , n8798 );
buf ( n8800 , n8799 );
buf ( n8801 , n8800 );
and ( n8802 , n8646 , n8801 );
buf ( n8803 , n8802 );
not ( n8804 , n8803 );
or ( n8805 , n8213 , n8804 );
buf ( n8806 , n8598 );
not ( n8807 , n8806 );
buf ( n8808 , n8618 );
nand ( n8809 , n8807 , n8808 );
buf ( n8810 , n8809 );
buf ( n8811 , n8810 );
not ( n8812 , n8811 );
not ( n8813 , n8641 );
nor ( n8814 , n8624 , n8813 );
buf ( n8815 , n8814 );
buf ( n8816 , n8620 );
nand ( n8817 , n8815 , n8816 );
buf ( n8818 , n8817 );
buf ( n8819 , n8818 );
not ( n8820 , n8819 );
or ( n8821 , n8812 , n8820 );
buf ( n8822 , n8796 );
not ( n8823 , n8822 );
buf ( n8824 , n8783 );
nand ( n8825 , n8823 , n8824 );
buf ( n8826 , n8825 );
buf ( n8827 , n8826 );
nand ( n8828 , n8821 , n8827 );
buf ( n8829 , n8828 );
buf ( n8830 , n8829 );
not ( n8831 , n8783 );
buf ( n8832 , n8796 );
nand ( n8833 , n8831 , n8832 );
buf ( n8834 , n8833 );
nand ( n8835 , n8830 , n8834 );
buf ( n8836 , n8835 );
buf ( n8837 , n8836 );
not ( n8838 , n8837 );
buf ( n8839 , n8838 );
nand ( n8840 , n8805 , n8839 );
buf ( n8841 , n371 );
buf ( n8842 , n379 );
nand ( n8843 , n8841 , n8842 );
buf ( n8844 , n8843 );
buf ( n8845 , n370 );
buf ( n8846 , n380 );
nand ( n8847 , n8845 , n8846 );
buf ( n8848 , n8847 );
xor ( n8849 , n8844 , n8848 );
buf ( n8850 , n372 );
buf ( n8851 , n378 );
nand ( n8852 , n8850 , n8851 );
buf ( n8853 , n8852 );
xor ( n8854 , n8849 , n8853 );
xor ( n8855 , n8733 , n8734 );
and ( n8856 , n8855 , n8736 );
and ( n8857 , n8733 , n8734 );
or ( n8858 , n8856 , n8857 );
xor ( n8859 , n8724 , n8731 );
and ( n8860 , n8859 , n8737 );
and ( n8861 , n8724 , n8731 );
or ( n8862 , n8860 , n8861 );
xor ( n8863 , n8858 , n8862 );
xor ( n8864 , n8854 , n8863 );
not ( n8865 , n8864 );
not ( n8866 , n7298 );
nand ( n8867 , n8866 , n6528 );
not ( n8868 , n7617 );
nand ( n8869 , n8868 , n6539 );
nand ( n8870 , n8867 , n8869 );
not ( n8871 , n8870 );
or ( n8872 , n8865 , n8871 );
not ( n8873 , n8864 );
and ( n8874 , n8869 , n8873 );
not ( n8875 , n8874 );
not ( n8876 , n8867 );
or ( n8877 , n8875 , n8876 );
not ( n8878 , n8723 );
not ( n8879 , n8738 );
or ( n8880 , n8878 , n8879 );
buf ( n8881 , n8751 );
buf ( n8882 , n8723 );
not ( n8883 , n8882 );
buf ( n8884 , n8741 );
nand ( n8885 , n8883 , n8884 );
buf ( n8886 , n8885 );
buf ( n8887 , n8886 );
nand ( n8888 , n8881 , n8887 );
buf ( n8889 , n8888 );
nand ( n8890 , n8880 , n8889 );
nand ( n8891 , n8877 , n8890 );
nand ( n8892 , n8872 , n8891 );
buf ( n8893 , n8892 );
buf ( n8894 , n7013 );
not ( n8895 , n8894 );
xor ( n8896 , n8668 , n8372 );
xor ( n8897 , n8896 , n411 );
buf ( n8898 , n8897 );
not ( n8899 , n8898 );
or ( n8900 , n8895 , n8899 );
not ( n8901 , n411 );
buf ( n8902 , n7445 );
not ( n8903 , n8902 );
buf ( n8904 , n8903 );
not ( n8905 , n8904 );
or ( n8906 , n8901 , n8905 );
buf ( n8907 , n411 );
not ( n8908 , n8907 );
buf ( n8909 , n7445 );
nand ( n8910 , n8908 , n8909 );
buf ( n8911 , n8910 );
nand ( n8912 , n8906 , n8911 );
buf ( n8913 , n8912 );
buf ( n8914 , n5837 );
nand ( n8915 , n8913 , n8914 );
buf ( n8916 , n8915 );
buf ( n8917 , n8916 );
nand ( n8918 , n8900 , n8917 );
buf ( n8919 , n8918 );
buf ( n8920 , n8919 );
xor ( n8921 , n8893 , n8920 );
not ( n8922 , n7013 );
not ( n8923 , n8912 );
or ( n8924 , n8922 , n8923 );
nand ( n8925 , n8651 , n5837 );
nand ( n8926 , n8924 , n8925 );
not ( n8927 , n8926 );
not ( n8928 , n6478 );
and ( n8929 , n8433 , n6496 );
not ( n8930 , n8433 );
and ( n8931 , n8930 , n413 );
or ( n8932 , n8929 , n8931 );
nand ( n8933 , n8932 , n7260 );
buf ( n8934 , n8684 );
buf ( n8935 , n6520 );
nand ( n8936 , n8934 , n8935 );
buf ( n8937 , n8936 );
nand ( n8938 , n8928 , n8933 , n8937 );
not ( n8939 , n8938 );
or ( n8940 , n8927 , n8939 );
buf ( n8941 , n6574 );
nand ( n8942 , n8933 , n8937 );
buf ( n8943 , n8942 );
nand ( n8944 , n8941 , n8943 );
buf ( n8945 , n8944 );
nand ( n8946 , n8940 , n8945 );
buf ( n8947 , n8946 );
xor ( n8948 , n8921 , n8947 );
buf ( n8949 , n8948 );
not ( n8950 , n8890 );
not ( n8951 , n8864 );
and ( n8952 , n8950 , n8951 );
and ( n8953 , n8890 , n8864 );
nor ( n8954 , n8952 , n8953 );
not ( n8955 , n8954 );
not ( n8956 , n8870 );
or ( n8957 , n8955 , n8956 );
or ( n8958 , n8870 , n8954 );
nand ( n8959 , n8957 , n8958 );
buf ( n8960 , n8959 );
buf ( n8961 , n8754 );
not ( n8962 , n8961 );
buf ( n8963 , n8962 );
buf ( n8964 , n8963 );
not ( n8965 , n8964 );
buf ( n8966 , n8719 );
not ( n8967 , n8966 );
or ( n8968 , n8965 , n8967 );
buf ( n8969 , n8719 );
buf ( n8970 , n8963 );
or ( n8971 , n8969 , n8970 );
buf ( n8972 , n8759 );
nand ( n8973 , n8971 , n8972 );
buf ( n8974 , n8973 );
buf ( n8975 , n8974 );
nand ( n8976 , n8968 , n8975 );
buf ( n8977 , n8976 );
buf ( n8978 , n8977 );
not ( n8979 , n8978 );
buf ( n8980 , n8979 );
buf ( n8981 , n8980 );
xor ( n8982 , n8960 , n8981 );
not ( n8983 , n8694 );
buf ( n8984 , n8663 );
not ( n8985 , n8984 );
buf ( n8986 , n8985 );
not ( n8987 , n8986 );
and ( n8988 , n8983 , n8987 );
buf ( n8989 , n8694 );
buf ( n8990 , n8986 );
nand ( n8991 , n8989 , n8990 );
buf ( n8992 , n8991 );
and ( n8993 , n8992 , n8653 );
nor ( n8994 , n8988 , n8993 );
buf ( n8995 , n8994 );
and ( n8996 , n8982 , n8995 );
and ( n8997 , n8960 , n8981 );
or ( n8998 , n8996 , n8997 );
buf ( n8999 , n8998 );
xor ( n9000 , n8949 , n8999 );
buf ( n9001 , n7298 );
not ( n9002 , n9001 );
buf ( n9003 , n6539 );
not ( n9004 , n9003 );
buf ( n9005 , n9004 );
buf ( n9006 , n9005 );
not ( n9007 , n9006 );
and ( n9008 , n9002 , n9007 );
buf ( n9009 , n7335 );
not ( n9010 , n9009 );
buf ( n9011 , n9010 );
buf ( n9012 , n9011 );
buf ( n9013 , n6528 );
and ( n9014 , n9012 , n9013 );
nor ( n9015 , n9008 , n9014 );
buf ( n9016 , n9015 );
buf ( n9017 , n9016 );
buf ( n9018 , n6520 );
not ( n9019 , n9018 );
buf ( n9020 , n8932 );
not ( n9021 , n9020 );
or ( n9022 , n9019 , n9021 );
nand ( n9023 , n6500 , n7260 );
buf ( n9024 , n9023 );
nand ( n9025 , n9022 , n9024 );
buf ( n9026 , n9025 );
buf ( n9027 , n9026 );
not ( n9028 , n9027 );
buf ( n9029 , n9028 );
buf ( n9030 , n9029 );
xor ( n9031 , n9017 , n9030 );
buf ( n9032 , n371 );
buf ( n9033 , n378 );
nand ( n9034 , n9032 , n9033 );
buf ( n9035 , n9034 );
buf ( n9036 , n370 );
buf ( n9037 , n379 );
nand ( n9038 , n9036 , n9037 );
buf ( n9039 , n9038 );
xor ( n9040 , n9035 , n9039 );
xor ( n9041 , n8844 , n8848 );
and ( n9042 , n9041 , n8853 );
and ( n9043 , n8844 , n8848 );
or ( n9044 , n9042 , n9043 );
xor ( n9045 , n9040 , n9044 );
xor ( n9046 , n8844 , n8848 );
xor ( n9047 , n9046 , n8853 );
and ( n9048 , n8858 , n9047 );
xor ( n9049 , n8844 , n8848 );
xor ( n9050 , n9049 , n8853 );
and ( n9051 , n8862 , n9050 );
and ( n9052 , n8858 , n8862 );
or ( n9053 , n9048 , n9051 , n9052 );
xor ( n9054 , n9053 , n6484 );
xor ( n9055 , n9045 , n9054 );
buf ( n9056 , n9055 );
xnor ( n9057 , n9031 , n9056 );
buf ( n9058 , n9057 );
buf ( n9059 , n9058 );
not ( n9060 , n9059 );
buf ( n9061 , n9060 );
and ( n9062 , n9000 , n9061 );
not ( n9063 , n9000 );
and ( n9064 , n9063 , n9058 );
nor ( n9065 , n9062 , n9064 );
buf ( n9066 , n9065 );
xor ( n9067 , n8960 , n8981 );
xor ( n9068 , n9067 , n8995 );
buf ( n9069 , n9068 );
not ( n9070 , n9069 );
xor ( n9071 , n8926 , n8942 );
not ( n9072 , n6574 );
and ( n9073 , n9071 , n9072 );
not ( n9074 , n9071 );
and ( n9075 , n9074 , n6574 );
nor ( n9076 , n9073 , n9075 );
not ( n9077 , n9076 );
and ( n9078 , n9070 , n9077 );
nand ( n9079 , n9069 , n9076 );
not ( n9080 , n8768 );
nand ( n9081 , n9080 , n8761 );
not ( n9082 , n9081 );
not ( n9083 , n8777 );
or ( n9084 , n9082 , n9083 );
buf ( n9085 , n8761 );
not ( n9086 , n9085 );
buf ( n9087 , n8768 );
nand ( n9088 , n9086 , n9087 );
buf ( n9089 , n9088 );
nand ( n9090 , n9084 , n9089 );
and ( n9091 , n9079 , n9090 );
nor ( n9092 , n9078 , n9091 );
buf ( n9093 , n9092 );
nand ( n9094 , n9066 , n9093 );
buf ( n9095 , n9094 );
buf ( n9096 , n9095 );
not ( n9097 , n9076 );
not ( n9098 , n9097 );
not ( n9099 , n9090 );
not ( n9100 , n9099 );
or ( n9101 , n9098 , n9100 );
nand ( n9102 , n9076 , n9090 );
nand ( n9103 , n9101 , n9102 );
not ( n9104 , n9069 );
and ( n9105 , n9103 , n9104 );
not ( n9106 , n9103 );
and ( n9107 , n9106 , n9069 );
nor ( n9108 , n9105 , n9107 );
buf ( n9109 , n9108 );
not ( n9110 , n9109 );
buf ( n9111 , n9110 );
buf ( n9112 , n9111 );
buf ( n9113 , n8697 );
not ( n9114 , n9113 );
buf ( n9115 , n9114 );
buf ( n9116 , n9115 );
not ( n9117 , n9116 );
buf ( n9118 , n8780 );
not ( n9119 , n9118 );
buf ( n9120 , n9119 );
buf ( n9121 , n9120 );
not ( n9122 , n9121 );
or ( n9123 , n9117 , n9122 );
buf ( n9124 , n8702 );
nand ( n9125 , n9123 , n9124 );
buf ( n9126 , n9125 );
buf ( n9127 , n9126 );
buf ( n9128 , n9120 );
buf ( n9129 , n9115 );
or ( n9130 , n9128 , n9129 );
buf ( n9131 , n9130 );
buf ( n9132 , n9131 );
nand ( n9133 , n9127 , n9132 );
buf ( n9134 , n9133 );
buf ( n9135 , n9134 );
not ( n9136 , n9135 );
buf ( n9137 , n9136 );
buf ( n9138 , n9137 );
nand ( n9139 , n9112 , n9138 );
buf ( n9140 , n9139 );
buf ( n9141 , n9140 );
and ( n9142 , n9096 , n9141 );
buf ( n9143 , n9142 );
xor ( n9144 , n8893 , n8920 );
and ( n9145 , n9144 , n8947 );
and ( n9146 , n8893 , n8920 );
or ( n9147 , n9145 , n9146 );
buf ( n9148 , n9147 );
buf ( n9149 , n9029 );
buf ( n9150 , n9016 );
nand ( n9151 , n9149 , n9150 );
buf ( n9152 , n9151 );
buf ( n9153 , n9152 );
not ( n9154 , n9153 );
buf ( n9155 , n9055 );
not ( n9156 , n9155 );
or ( n9157 , n9154 , n9156 );
buf ( n9158 , n9016 );
not ( n9159 , n9158 );
buf ( n9160 , n9026 );
nand ( n9161 , n9159 , n9160 );
buf ( n9162 , n9161 );
buf ( n9163 , n9162 );
nand ( n9164 , n9157 , n9163 );
buf ( n9165 , n9164 );
buf ( n9166 , n9165 );
not ( n9167 , n9166 );
buf ( n9168 , n9167 );
xor ( n9169 , n9148 , n9168 );
xor ( n9170 , n9035 , n9039 );
xor ( n9171 , n9170 , n9044 );
and ( n9172 , n9053 , n9171 );
xor ( n9173 , n9035 , n9039 );
xor ( n9174 , n9173 , n9044 );
and ( n9175 , n6484 , n9174 );
and ( n9176 , n9053 , n6484 );
or ( n9177 , n9172 , n9175 , n9176 );
xor ( n9178 , n6560 , n9177 );
buf ( n9179 , n370 );
buf ( n9180 , n378 );
nand ( n9181 , n9179 , n9180 );
buf ( n9182 , n9181 );
buf ( n9183 , n9182 );
xor ( n9184 , n9035 , n9039 );
and ( n9185 , n9184 , n9044 );
and ( n9186 , n9035 , n9039 );
or ( n9187 , n9185 , n9186 );
buf ( n9188 , n9187 );
xor ( n9189 , n9183 , n9188 );
buf ( n9190 , n6484 );
xor ( n9191 , n9189 , n9190 );
buf ( n9192 , n9191 );
xor ( n9193 , n9178 , n9192 );
buf ( n9194 , n6528 );
not ( n9195 , n9194 );
buf ( n9196 , n8904 );
not ( n9197 , n9196 );
buf ( n9198 , n9197 );
buf ( n9199 , n9198 );
not ( n9200 , n9199 );
or ( n9201 , n9195 , n9200 );
buf ( n9202 , n9011 );
buf ( n9203 , n6539 );
nand ( n9204 , n9202 , n9203 );
buf ( n9205 , n9204 );
buf ( n9206 , n9205 );
nand ( n9207 , n9201 , n9206 );
buf ( n9208 , n9207 );
buf ( n9209 , n9208 );
not ( n9210 , n9209 );
buf ( n9211 , n7013 );
not ( n9212 , n9211 );
and ( n9213 , n411 , n8436 );
not ( n9214 , n411 );
buf ( n9215 , n8436 );
not ( n9216 , n9215 );
buf ( n9217 , n9216 );
and ( n9218 , n9214 , n9217 );
or ( n9219 , n9213 , n9218 );
buf ( n9220 , n9219 );
not ( n9221 , n9220 );
or ( n9222 , n9212 , n9221 );
buf ( n9223 , n8897 );
buf ( n9224 , n5837 );
nand ( n9225 , n9223 , n9224 );
buf ( n9226 , n9225 );
buf ( n9227 , n9226 );
nand ( n9228 , n9222 , n9227 );
buf ( n9229 , n9228 );
buf ( n9230 , n9229 );
not ( n9231 , n9230 );
buf ( n9232 , n9231 );
buf ( n9233 , n9232 );
not ( n9234 , n9233 );
or ( n9235 , n9210 , n9234 );
buf ( n9236 , n9232 );
buf ( n9237 , n9208 );
or ( n9238 , n9236 , n9237 );
nand ( n9239 , n9235 , n9238 );
buf ( n9240 , n9239 );
xor ( n9241 , n9193 , n9240 );
xnor ( n9242 , n9169 , n9241 );
not ( n9243 , n9242 );
buf ( n9244 , n8949 );
not ( n9245 , n9244 );
buf ( n9246 , n9245 );
buf ( n9247 , n9246 );
not ( n9248 , n9247 );
buf ( n9249 , n9058 );
not ( n9250 , n9249 );
or ( n9251 , n9248 , n9250 );
buf ( n9252 , n8999 );
not ( n9253 , n9252 );
buf ( n9254 , n9253 );
buf ( n9255 , n9254 );
nand ( n9256 , n9251 , n9255 );
buf ( n9257 , n9256 );
buf ( n9258 , n9257 );
buf ( n9259 , n9246 );
not ( n9260 , n9259 );
buf ( n9261 , n9061 );
nand ( n9262 , n9260 , n9261 );
buf ( n9263 , n9262 );
buf ( n9264 , n9263 );
nand ( n9265 , n9258 , n9264 );
buf ( n9266 , n9265 );
buf ( n9267 , n9266 );
not ( n9268 , n9267 );
buf ( n9269 , n9268 );
nand ( n9270 , n9243 , n9269 );
xor ( n9271 , n6560 , n9177 );
and ( n9272 , n9271 , n9192 );
and ( n9273 , n6560 , n9177 );
or ( n9274 , n9272 , n9273 );
buf ( n9275 , n9208 );
not ( n9276 , n9275 );
buf ( n9277 , n9232 );
nand ( n9278 , n9276 , n9277 );
buf ( n9279 , n9278 );
not ( n9280 , n9279 );
not ( n9281 , n9193 );
or ( n9282 , n9280 , n9281 );
buf ( n9283 , n9229 );
buf ( n9284 , n9208 );
nand ( n9285 , n9283 , n9284 );
buf ( n9286 , n9285 );
nand ( n9287 , n9282 , n9286 );
xor ( n9288 , n9274 , n9287 );
buf ( n9289 , n6484 );
not ( n9290 , n9289 );
buf ( n9291 , n9290 );
xor ( n9292 , n6557 , n9291 );
buf ( n9293 , n9292 );
xor ( n9294 , n9183 , n9188 );
and ( n9295 , n9294 , n9190 );
and ( n9296 , n9183 , n9188 );
or ( n9297 , n9295 , n9296 );
buf ( n9298 , n9297 );
buf ( n9299 , n9298 );
xor ( n9300 , n9293 , n9299 );
buf ( n9301 , n9300 );
buf ( n9302 , n9301 );
not ( n9303 , n9302 );
buf ( n9304 , n9303 );
not ( n9305 , n9304 );
buf ( n9306 , n5837 );
not ( n9307 , n9306 );
buf ( n9308 , n9219 );
not ( n9309 , n9308 );
or ( n9310 , n9307 , n9309 );
nand ( n9311 , n6444 , n7013 );
buf ( n9312 , n9311 );
nand ( n9313 , n9310 , n9312 );
buf ( n9314 , n9313 );
buf ( n9315 , n9314 );
not ( n9316 , n9315 );
buf ( n9317 , n6539 );
not ( n9318 , n9317 );
buf ( n9319 , n9198 );
not ( n9320 , n9319 );
or ( n9321 , n9318 , n9320 );
buf ( n9322 , n8896 );
buf ( n9323 , n6528 );
nand ( n9324 , n9322 , n9323 );
buf ( n9325 , n9324 );
buf ( n9326 , n9325 );
nand ( n9327 , n9321 , n9326 );
buf ( n9328 , n9327 );
buf ( n9329 , n9328 );
not ( n9330 , n9329 );
buf ( n9331 , n9330 );
buf ( n9332 , n9331 );
not ( n9333 , n9332 );
and ( n9334 , n9316 , n9333 );
buf ( n9335 , n9314 );
buf ( n9336 , n9331 );
and ( n9337 , n9335 , n9336 );
nor ( n9338 , n9334 , n9337 );
buf ( n9339 , n9338 );
buf ( n9340 , n9339 );
not ( n9341 , n9340 );
buf ( n9342 , n9341 );
not ( n9343 , n9342 );
or ( n9344 , n9305 , n9343 );
buf ( n9345 , n9301 );
buf ( n9346 , n9339 );
nand ( n9347 , n9345 , n9346 );
buf ( n9348 , n9347 );
nand ( n9349 , n9344 , n9348 );
xor ( n9350 , n9288 , n9349 );
not ( n9351 , n9350 );
buf ( n9352 , n9148 );
not ( n9353 , n9352 );
buf ( n9354 , n9168 );
nand ( n9355 , n9353 , n9354 );
buf ( n9356 , n9355 );
not ( n9357 , n9356 );
not ( n9358 , n9241 );
or ( n9359 , n9357 , n9358 );
buf ( n9360 , n9148 );
buf ( n9361 , n9165 );
nand ( n9362 , n9360 , n9361 );
buf ( n9363 , n9362 );
nand ( n9364 , n9359 , n9363 );
not ( n9365 , n9364 );
nand ( n9366 , n9351 , n9365 );
and ( n9367 , n8840 , n9143 , n9270 , n9366 );
buf ( n9368 , n9314 );
not ( n9369 , n9368 );
buf ( n9370 , n9331 );
nand ( n9371 , n9369 , n9370 );
buf ( n9372 , n9371 );
not ( n9373 , n9372 );
not ( n9374 , n9301 );
or ( n9375 , n9373 , n9374 );
buf ( n9376 , n9331 );
not ( n9377 , n9376 );
buf ( n9378 , n9314 );
nand ( n9379 , n9377 , n9378 );
buf ( n9380 , n9379 );
nand ( n9381 , n9375 , n9380 );
not ( n9382 , n9381 );
not ( n9383 , n9382 );
not ( n9384 , n9383 );
not ( n9385 , n6445 );
and ( n9386 , n6557 , n9291 );
buf ( n9387 , n9386 );
not ( n9388 , n9387 );
buf ( n9389 , n6574 );
buf ( n9390 , n6560 );
nand ( n9391 , n9389 , n9390 );
buf ( n9392 , n9391 );
buf ( n9393 , n9392 );
nand ( n9394 , n9388 , n9393 );
buf ( n9395 , n9394 );
xor ( n9396 , n9385 , n9395 );
not ( n9397 , n9386 );
buf ( n9398 , n9397 );
not ( n9399 , n9398 );
buf ( n9400 , n9298 );
not ( n9401 , n9400 );
or ( n9402 , n9399 , n9401 );
buf ( n9403 , n9392 );
nand ( n9404 , n9402 , n9403 );
buf ( n9405 , n9404 );
xnor ( n9406 , n9396 , n9405 );
not ( n9407 , n9406 );
not ( n9408 , n9407 );
or ( n9409 , n9384 , n9408 );
not ( n9410 , n9382 );
not ( n9411 , n9406 );
or ( n9412 , n9410 , n9411 );
not ( n9413 , n6528 );
not ( n9414 , n9217 );
or ( n9415 , n9413 , n9414 );
buf ( n9416 , n8896 );
buf ( n9417 , n6539 );
nand ( n9418 , n9416 , n9417 );
buf ( n9419 , n9418 );
nand ( n9420 , n9415 , n9419 );
nand ( n9421 , n9412 , n9420 );
nand ( n9422 , n9409 , n9421 );
or ( n9423 , n9405 , n6581 );
nand ( n9424 , n9423 , n9395 );
buf ( n9425 , n9405 );
buf ( n9426 , n6581 );
nand ( n9427 , n9425 , n9426 );
buf ( n9428 , n9427 );
nand ( n9429 , n9424 , n9428 );
not ( n9430 , n9429 );
buf ( n9431 , n6539 );
not ( n9432 , n9431 );
buf ( n9433 , n9217 );
not ( n9434 , n9433 );
or ( n9435 , n9432 , n9434 );
buf ( n9436 , n6531 );
nand ( n9437 , n9435 , n9436 );
buf ( n9438 , n9437 );
not ( n9439 , n9438 );
not ( n9440 , n9439 );
buf ( n9441 , n9072 );
buf ( n9442 , n9397 );
nand ( n9443 , n9441 , n9442 );
buf ( n9444 , n9443 );
not ( n9445 , n6557 );
not ( n9446 , n6487 );
or ( n9447 , n9445 , n9446 );
buf ( n9448 , n6550 );
buf ( n9449 , n6445 );
nand ( n9450 , n9448 , n9449 );
buf ( n9451 , n9450 );
nand ( n9452 , n9447 , n9451 );
buf ( n9453 , n9452 );
not ( n9454 , n9453 );
buf ( n9455 , n9454 );
xor ( n9456 , n9444 , n9455 );
not ( n9457 , n9456 );
or ( n9458 , n9440 , n9457 );
or ( n9459 , n9456 , n9439 );
nand ( n9460 , n9458 , n9459 );
not ( n9461 , n9460 );
or ( n9462 , n9430 , n9461 );
or ( n9463 , n9429 , n9460 );
nand ( n9464 , n9462 , n9463 );
nor ( n9465 , n9422 , n9464 );
not ( n9466 , n9465 );
not ( n9467 , n9429 );
buf ( n9468 , n9438 );
not ( n9469 , n9468 );
buf ( n9470 , n9456 );
nand ( n9471 , n9469 , n9470 );
buf ( n9472 , n9471 );
not ( n9473 , n9472 );
or ( n9474 , n9467 , n9473 );
buf ( n9475 , n9456 );
not ( n9476 , n9475 );
buf ( n9477 , n9438 );
nand ( n9478 , n9476 , n9477 );
buf ( n9479 , n9478 );
nand ( n9480 , n9474 , n9479 );
buf ( n9481 , n9480 );
not ( n9482 , n9481 );
not ( n9483 , n9072 );
buf ( n9484 , n6550 );
not ( n9485 , n9484 );
buf ( n9486 , n6445 );
nand ( n9487 , n9485 , n9486 );
buf ( n9488 , n9487 );
not ( n9489 , n9488 );
or ( n9490 , n9483 , n9489 );
buf ( n9491 , n9488 );
not ( n9492 , n9491 );
buf ( n9493 , n9492 );
nand ( n9494 , n6574 , n9493 );
nand ( n9495 , n9490 , n9494 );
not ( n9496 , n9452 );
and ( n9497 , n9495 , n9496 );
not ( n9498 , n9495 );
and ( n9499 , n9498 , n9452 );
nor ( n9500 , n9497 , n9499 );
buf ( n9501 , n9500 );
not ( n9502 , n9501 );
buf ( n9503 , n6542 );
not ( n9504 , n9503 );
and ( n9505 , n9502 , n9504 );
buf ( n9506 , n9500 );
buf ( n9507 , n6542 );
and ( n9508 , n9506 , n9507 );
nor ( n9509 , n9505 , n9508 );
buf ( n9510 , n9509 );
buf ( n9511 , n9510 );
buf ( n9512 , n9072 );
buf ( n9513 , n9452 );
nand ( n9514 , n9512 , n9513 );
buf ( n9515 , n9514 );
buf ( n9516 , n9515 );
buf ( n9517 , n9397 );
nand ( n9518 , n9516 , n9517 );
buf ( n9519 , n9518 );
buf ( n9520 , n9519 );
and ( n9521 , n9511 , n9520 );
not ( n9522 , n9511 );
buf ( n9523 , n9519 );
not ( n9524 , n9523 );
buf ( n9525 , n9524 );
buf ( n9526 , n9525 );
and ( n9527 , n9522 , n9526 );
nor ( n9528 , n9521 , n9527 );
buf ( n9529 , n9528 );
buf ( n9530 , n9529 );
not ( n9531 , n9530 );
buf ( n9532 , n9531 );
buf ( n9533 , n9532 );
nand ( n9534 , n9482 , n9533 );
buf ( n9535 , n9534 );
nand ( n9536 , n9466 , n9535 );
buf ( n9537 , n9536 );
not ( n9538 , n9349 );
not ( n9539 , n9274 );
or ( n9540 , n9538 , n9539 );
nor ( n9541 , n9349 , n9274 );
not ( n9542 , n9287 );
or ( n9543 , n9541 , n9542 );
nand ( n9544 , n9540 , n9543 );
xor ( n9545 , n9420 , n9381 );
xnor ( n9546 , n9545 , n9406 );
nor ( n9547 , n9544 , n9546 );
buf ( n9548 , n9547 );
buf ( n9549 , n6542 );
not ( n9550 , n9549 );
buf ( n9551 , n9519 );
not ( n9552 , n9551 );
or ( n9553 , n9550 , n9552 );
buf ( n9554 , n9500 );
nand ( n9555 , n9553 , n9554 );
buf ( n9556 , n9555 );
buf ( n9557 , n9556 );
buf ( n9558 , n9525 );
not ( n9559 , n6542 );
buf ( n9560 , n9559 );
nand ( n9561 , n9558 , n9560 );
buf ( n9562 , n9561 );
buf ( n9563 , n9562 );
nand ( n9564 , n9557 , n9563 );
buf ( n9565 , n9564 );
buf ( n9566 , n6566 );
and ( n9567 , n6491 , n9493 );
not ( n9568 , n6491 );
and ( n9569 , n9568 , n9488 );
or ( n9570 , n9567 , n9569 );
buf ( n9571 , n9570 );
xor ( n9572 , n9566 , n9571 );
not ( n9573 , n9515 );
not ( n9574 , n9488 );
or ( n9575 , n9573 , n9574 );
buf ( n9576 , n9455 );
buf ( n9577 , n6574 );
nand ( n9578 , n9576 , n9577 );
buf ( n9579 , n9578 );
nand ( n9580 , n9575 , n9579 );
buf ( n9581 , n9580 );
xor ( n9582 , n9572 , n9581 );
buf ( n9583 , n9582 );
buf ( n9584 , C1 );
buf ( n9585 , C0 );
buf ( n9586 , n9585 );
nand ( n9587 , n9570 , n6565 );
buf ( n9588 , n9587 );
buf ( n9589 , n6566 );
not ( n9590 , n9589 );
buf ( n9591 , n9570 );
not ( n9592 , n9591 );
buf ( n9593 , n9592 );
buf ( n9594 , n9593 );
not ( n9595 , n9594 );
or ( n9596 , n9590 , n9595 );
buf ( n9597 , n9580 );
nand ( n9598 , n9596 , n9597 );
buf ( n9599 , n9598 );
buf ( n9600 , n9599 );
nand ( n9601 , n9588 , n9600 );
buf ( n9602 , n9601 );
buf ( n9603 , n6574 );
buf ( n9604 , n6581 );
nor ( n9605 , n9603 , n9604 );
buf ( n9606 , n9605 );
or ( n9607 , n9606 , n9493 );
not ( n9608 , n9607 );
not ( n9609 , n6599 );
or ( n9610 , n9608 , n9609 );
buf ( n9611 , n6599 );
or ( n9612 , n9611 , n9607 );
nand ( n9613 , n9610 , n9612 );
buf ( n9614 , n6567 );
nor ( n9615 , n9606 , n9493 );
buf ( n9616 , n9615 );
nand ( n9617 , n9614 , n9616 );
buf ( n9618 , n9617 );
nand ( n9619 , n9618 , n6588 );
buf ( n9620 , C0 );
buf ( n9621 , n9620 );
nor ( n9622 , n9537 , n9548 , n9586 , n9621 );
buf ( n9623 , n9622 );
nand ( n9624 , n9367 , n9623 );
nand ( n9625 , n9546 , n9544 );
nand ( n9626 , n9422 , n9464 );
buf ( n9627 , n9480 );
buf ( n9628 , n9529 );
nand ( n9629 , n9627 , n9628 );
buf ( n9630 , n9629 );
nand ( n9631 , n9625 , n9626 , n9630 );
buf ( n9632 , n6613 );
buf ( n9633 , n9619 );
nand ( n9634 , n9632 , n9633 );
buf ( n9635 , n9634 );
buf ( n9636 , C1 );
and ( n9637 , n9631 , n9636 , n9584 );
buf ( n9638 , n9637 );
buf ( n9639 , n9536 );
buf ( n9640 , n9630 );
nand ( n9641 , n9639 , n9640 );
buf ( n9642 , n9641 );
buf ( n9643 , n9642 );
and ( n9644 , n9638 , n9643 );
buf ( n9645 , n9602 );
not ( n9646 , n9645 );
buf ( n9647 , n9613 );
not ( n9648 , n9647 );
or ( n9649 , n9646 , n9648 );
buf ( n9650 , n9583 );
not ( n9651 , n9650 );
buf ( n9652 , n9565 );
nand ( n9653 , n9651 , n9652 );
buf ( n9654 , n9653 );
buf ( n9655 , n9654 );
nand ( n9656 , n9649 , n9655 );
buf ( n9657 , n9656 );
not ( n9658 , n9657 );
nand ( n9659 , n9658 , n9635 );
not ( n9660 , n9659 );
or ( n9661 , n9660 , C0 );
buf ( n9662 , n6613 );
buf ( n9663 , n6589 );
nand ( n9664 , n9662 , n9663 );
buf ( n9665 , n9664 );
nand ( n9666 , n9661 , n9665 );
buf ( n9667 , n9666 );
nor ( n9668 , n9644 , n9667 );
buf ( n9669 , n9668 );
buf ( n9670 , n9108 );
buf ( n9671 , n9134 );
nand ( n9672 , n9670 , n9671 );
buf ( n9673 , n9672 );
buf ( n9674 , n9673 );
not ( n9675 , n9674 );
buf ( n9676 , n9095 );
nand ( n9677 , n9675 , n9676 );
buf ( n9678 , n9677 );
buf ( n9679 , n9678 );
buf ( n9680 , n9065 );
not ( n9681 , n9680 );
buf ( n9682 , n9681 );
buf ( n9683 , n9682 );
buf ( n9684 , n9092 );
not ( n9685 , n9684 );
buf ( n9686 , n9685 );
buf ( n9687 , n9686 );
nand ( n9688 , n9683 , n9687 );
buf ( n9689 , n9688 );
buf ( n9690 , n9689 );
nand ( n9691 , n9679 , n9690 );
buf ( n9692 , n9691 );
not ( n9693 , n9692 );
not ( n9694 , n9270 );
or ( n9695 , n9693 , n9694 );
buf ( n9696 , n9350 );
buf ( n9697 , n9364 );
nand ( n9698 , n9696 , n9697 );
buf ( n9699 , n9698 );
buf ( n9700 , n9269 );
not ( n9701 , n9700 );
buf ( n9702 , n9242 );
nand ( n9703 , n9701 , n9702 );
buf ( n9704 , n9703 );
nand ( n9705 , n9699 , n9704 );
not ( n9706 , n9705 );
nand ( n9707 , n9695 , n9706 );
not ( n9708 , n9480 );
not ( n9709 , n9529 );
and ( n9710 , n9708 , n9709 );
nor ( n9711 , n9710 , n9585 );
and ( n9712 , n9711 , n9366 );
not ( n9713 , n9547 );
and ( n9714 , n9636 , n9713 , n9466 );
nand ( n9715 , n9707 , n9712 , n9714 );
nand ( n9716 , n9624 , n9669 , n9715 );
not ( n9717 , n9716 );
not ( n9718 , n9717 );
or ( n9719 , C0 , n9718 );
buf ( n9720 , n9665 );
not ( n9721 , n9720 );
or ( n9722 , C0 , n9721 );
not ( n9723 , n9669 );
buf ( n9724 , n9723 );
nand ( n9725 , n9722 , n9724 );
buf ( n9726 , n9725 );
nand ( n9727 , n9719 , n9726 );
buf ( n9728 , n9727 );
buf ( n9729 , n381 );
not ( n9730 , n9729 );
buf ( n9731 , n9730 );
not ( n9732 , n380 );
and ( n9733 , n9731 , n9732 );
and ( n9734 , n380 , n381 );
nor ( n9735 , n9733 , n9734 );
buf ( n9736 , n382 );
not ( n9737 , n9736 );
buf ( n9738 , n9737 );
and ( n9739 , n381 , n9738 );
not ( n9740 , n381 );
and ( n9741 , n9740 , n382 );
nor ( n9742 , n9739 , n9741 );
and ( n9743 , n9735 , n9742 );
buf ( n9744 , n9743 );
not ( n9745 , n9742 );
buf ( n9746 , n9745 );
nor ( n9747 , n9744 , n9746 );
buf ( n9748 , n9747 );
buf ( n9749 , n9748 );
buf ( n9750 , n9732 );
or ( n9751 , n9749 , n9750 );
buf ( n9752 , n9751 );
buf ( n9753 , n9752 );
not ( n9754 , n9753 );
buf ( n9755 , n9754 );
buf ( n9756 , n9755 );
and ( n9757 , n9728 , n9756 );
buf ( n9758 , n9757 );
buf ( n9759 , n9758 );
buf ( n9760 , n9759 );
buf ( n9761 , n9760 );
buf ( n9762 , n9761 );
not ( n9763 , n9762 );
buf ( n9764 , n9763 );
buf ( n9765 , n9764 );
not ( n9766 , n9717 );
or ( n9767 , C0 , n9766 );
nand ( n9768 , n9767 , n9726 );
buf ( n9769 , n9768 );
and ( n9770 , n379 , n9732 );
not ( n9771 , n379 );
and ( n9772 , n9771 , n380 );
or ( n9773 , n9770 , n9772 );
not ( n9774 , n9773 );
buf ( n9775 , n9774 );
not ( n9776 , n378 );
buf ( n9777 , n9776 );
buf ( n9778 , n379 );
not ( n9779 , n9778 );
buf ( n9780 , n9779 );
buf ( n9781 , n9780 );
and ( n9782 , n9777 , n9781 );
buf ( n9783 , n378 );
buf ( n9784 , n379 );
and ( n9785 , n9783 , n9784 );
nor ( n9786 , n9782 , n9785 );
buf ( n9787 , n9786 );
buf ( n9788 , n9787 );
and ( n9789 , n9775 , n9788 );
buf ( n9790 , n9789 );
buf ( n9791 , n9790 );
not ( n9792 , n9791 );
buf ( n9793 , n9792 );
buf ( n9794 , n9793 );
buf ( n9795 , n9774 );
nand ( n9796 , n9794 , n9795 );
buf ( n9797 , n9796 );
buf ( n9798 , n9797 );
buf ( n9799 , n378 );
and ( n9800 , n9798 , n9799 );
buf ( n9801 , n9800 );
buf ( n9802 , n9801 );
nand ( n9803 , n9769 , n9802 );
buf ( n9804 , n9803 );
buf ( n9805 , n9804 );
buf ( n9806 , n9755 );
buf ( n9807 , n9801 );
nand ( n9808 , n9806 , n9807 );
buf ( n9809 , n9808 );
buf ( n9810 , n9809 );
and ( n9811 , n9765 , n9805 , n9810 );
buf ( n9812 , n9811 );
buf ( n9813 , n9812 );
not ( n9814 , n9813 );
buf ( n9815 , n9717 );
not ( n9816 , n9815 );
or ( n9817 , C0 , n9816 );
buf ( n9818 , n9726 );
nand ( n9819 , n9817 , n9818 );
buf ( n9820 , n9819 );
or ( n9821 , n9820 , n9755 );
nand ( n9822 , n9727 , n9755 );
nand ( n9823 , n9821 , n9822 );
buf ( n9824 , n9823 );
buf ( n9825 , n384 );
buf ( n9826 , n9801 );
not ( n9827 , n9826 );
buf ( n9828 , n9827 );
buf ( n9829 , n9828 );
and ( n9830 , n9825 , n9829 );
not ( n9831 , n9825 );
buf ( n9832 , n9801 );
and ( n9833 , n9831 , n9832 );
nor ( n9834 , n9830 , n9833 );
buf ( n9835 , n9834 );
xor ( n9836 , n383 , n384 );
buf ( n9837 , n9836 );
not ( n9838 , n9837 );
buf ( n9839 , n9838 );
buf ( n9840 , n9839 );
not ( n9841 , n9840 );
buf ( n9842 , n9738 );
buf ( n9843 , n383 );
not ( n9844 , n9843 );
buf ( n9845 , n9844 );
buf ( n9846 , n9845 );
and ( n9847 , n9842 , n9846 );
buf ( n9848 , n382 );
buf ( n9849 , n383 );
and ( n9850 , n9848 , n9849 );
nor ( n9851 , n9847 , n9850 );
buf ( n9852 , n9851 );
and ( n9853 , n9839 , n9852 );
not ( n9854 , n9853 );
buf ( n9855 , n9854 );
not ( n9856 , n9855 );
or ( n9857 , n9841 , n9856 );
buf ( n9858 , n382 );
nand ( n9859 , n9857 , n9858 );
buf ( n9860 , n9859 );
buf ( n9861 , n9860 );
not ( n9862 , n9861 );
buf ( n9863 , n9862 );
and ( n9864 , n9835 , n9863 );
not ( n9865 , n9835 );
and ( n9866 , n9865 , n9860 );
or ( n9867 , n9864 , n9866 );
not ( n9868 , n9867 );
buf ( n9869 , n9868 );
nand ( n9870 , n9824 , n9869 );
buf ( n9871 , n9870 );
buf ( n9872 , n9871 );
nand ( n9873 , n9814 , n9872 );
buf ( n9874 , n9873 );
buf ( n9875 , n9874 );
buf ( n9876 , n9868 );
not ( n9877 , n9876 );
buf ( n9878 , n9823 );
not ( n9879 , n9878 );
buf ( n9880 , n9879 );
buf ( n9881 , n9880 );
nand ( n9882 , n9877 , n9881 );
buf ( n9883 , n9882 );
buf ( n9884 , n9883 );
nand ( n9885 , n9875 , n9884 );
buf ( n9886 , n9885 );
buf ( n9887 , n9880 );
not ( n9888 , n9887 );
buf ( n9889 , n9888 );
not ( n9890 , n9889 );
buf ( n9891 , n9758 );
not ( n9892 , n9891 );
buf ( n9893 , n9863 );
buf ( n9894 , n384 );
and ( n9895 , n9893 , n9894 );
buf ( n9896 , n9895 );
buf ( n9897 , n9896 );
not ( n9898 , n9897 );
buf ( n9899 , n9898 );
buf ( n9900 , n384 );
not ( n9901 , n9900 );
buf ( n9902 , n9860 );
nand ( n9903 , n9901 , n9902 );
buf ( n9904 , n9903 );
nand ( n9905 , n9904 , n9801 );
and ( n9906 , n9899 , n9905 );
buf ( n9907 , n9906 );
not ( n9908 , n9907 );
and ( n9909 , n9892 , n9908 );
buf ( n9910 , n9758 );
buf ( n9911 , n9906 );
and ( n9912 , n9910 , n9911 );
nor ( n9913 , n9909 , n9912 );
buf ( n9914 , n9913 );
buf ( n9915 , n9914 );
not ( n9916 , n9915 );
buf ( n9917 , n9916 );
not ( n9918 , n9917 );
or ( n9919 , n9890 , n9918 );
buf ( n9920 , n9914 );
buf ( n9921 , n9880 );
nand ( n9922 , n9920 , n9921 );
buf ( n9923 , n9922 );
nand ( n9924 , n9919 , n9923 );
not ( n9925 , n9867 );
or ( n9926 , n9924 , n9925 );
nand ( n9927 , n9924 , n9868 );
nand ( n9928 , n9926 , n9927 );
buf ( n9929 , n9928 );
not ( n9930 , n9929 );
buf ( n9931 , n9930 );
and ( n9932 , n9886 , n9931 );
not ( n9933 , n9886 );
and ( n9934 , n9933 , n9928 );
or ( n9935 , n9932 , n9934 );
buf ( n9936 , n9904 );
not ( n9937 , n9936 );
buf ( n9938 , n9761 );
not ( n9939 , n9938 );
or ( n9940 , n9937 , n9939 );
buf ( n9941 , n9899 );
nand ( n9942 , n9940 , n9941 );
buf ( n9943 , n9942 );
not ( n9944 , n9812 );
not ( n9945 , n9944 );
and ( n9946 , n9867 , n9889 );
not ( n9947 , n9867 );
and ( n9948 , n9947 , n9880 );
or ( n9949 , n9946 , n9948 );
not ( n9950 , n9949 );
not ( n9951 , n9950 );
or ( n9952 , n9945 , n9951 );
nand ( n9953 , n9949 , n9812 );
nand ( n9954 , n9952 , n9953 );
xor ( n9955 , n9943 , n9954 );
buf ( n9956 , n384 );
buf ( n9957 , n9860 );
and ( n9958 , n9956 , n9957 );
not ( n9959 , n9956 );
buf ( n9960 , n9863 );
and ( n9961 , n9959 , n9960 );
nor ( n9962 , n9958 , n9961 );
buf ( n9963 , n9962 );
not ( n9964 , n9963 );
not ( n9965 , n9764 );
or ( n9966 , n9964 , n9965 );
buf ( n9967 , n9963 );
not ( n9968 , n9967 );
buf ( n9969 , n9968 );
nand ( n9970 , n9969 , n9761 );
nand ( n9971 , n9966 , n9970 );
buf ( n9972 , n9971 );
not ( n9973 , n9972 );
not ( n9974 , n9801 );
not ( n9975 , n9823 );
or ( n9976 , n9974 , n9975 );
buf ( n9977 , n9880 );
buf ( n9978 , n9828 );
nand ( n9979 , n9977 , n9978 );
buf ( n9980 , n9979 );
nand ( n9981 , n9976 , n9980 );
buf ( n9982 , n9981 );
not ( n9983 , n9982 );
buf ( n9984 , n9983 );
buf ( n9985 , n9984 );
not ( n9986 , n9985 );
or ( n9987 , n9973 , n9986 );
not ( n9988 , n9906 );
buf ( n9989 , n9988 );
nand ( n9990 , n9987 , n9989 );
buf ( n9991 , n9990 );
buf ( n9992 , n9991 );
buf ( n9993 , n9971 );
not ( n9994 , n9993 );
buf ( n9995 , n9981 );
nand ( n9996 , n9994 , n9995 );
buf ( n9997 , n9996 );
buf ( n9998 , n9997 );
nand ( n9999 , n9992 , n9998 );
buf ( n10000 , n9999 );
and ( n10001 , n9955 , n10000 );
and ( n10002 , n9943 , n9954 );
or ( n10003 , n10001 , n10002 );
buf ( n10004 , C0 );
nor ( n10005 , n9935 , n10003 );
buf ( n10006 , n10005 );
nor ( n10007 , n10004 , n10006 );
buf ( n10008 , n10007 );
buf ( n10009 , n10008 );
not ( n10010 , n10009 );
buf ( n10011 , n10010 );
buf ( n10012 , n10011 );
buf ( n10013 , n10008 );
xor ( n10014 , n9943 , n9954 );
xor ( n10015 , n10014 , n10000 );
not ( n10016 , n9871 );
not ( n10017 , n9896 );
or ( n10018 , n10016 , n10017 );
nand ( n10019 , n10018 , n9883 );
buf ( n10020 , n10019 );
not ( n10021 , n10020 );
buf ( n10022 , n10021 );
buf ( n10023 , n10022 );
not ( n10024 , n10023 );
xor ( n10025 , n9906 , n9981 );
xnor ( n10026 , n10025 , n9971 );
buf ( n10027 , n10026 );
not ( n10028 , n10027 );
or ( n10029 , n10024 , n10028 );
buf ( n10030 , n9969 );
buf ( n10031 , n9896 );
nor ( n10032 , n10030 , n10031 );
buf ( n10033 , n10032 );
buf ( n10034 , n10033 );
buf ( n10035 , n9752 );
or ( n10036 , n10034 , n10035 );
buf ( n10037 , n10036 );
buf ( n10038 , n10037 );
buf ( n10039 , n9969 );
not ( n10040 , n10039 );
buf ( n10041 , n9896 );
buf ( n10042 , n9752 );
and ( n10043 , n10041 , n10042 );
buf ( n10044 , n9899 );
buf ( n10045 , n9755 );
and ( n10046 , n10044 , n10045 );
nor ( n10047 , n10043 , n10046 );
buf ( n10048 , n10047 );
buf ( n10049 , n10048 );
not ( n10050 , n10049 );
or ( n10051 , n10040 , n10050 );
buf ( n10052 , n10048 );
buf ( n10053 , n9969 );
or ( n10054 , n10052 , n10053 );
nand ( n10055 , n10051 , n10054 );
buf ( n10056 , n10055 );
buf ( n10057 , n10056 );
not ( n10058 , n10057 );
buf ( n10059 , n10037 );
nand ( n10060 , n10058 , n10059 );
buf ( n10061 , n10060 );
nand ( n10062 , n10061 , n9768 );
buf ( n10063 , n10062 );
xor ( n10064 , n10038 , n10063 );
buf ( n10065 , n9896 );
buf ( n10066 , n9867 );
xor ( n10067 , n10065 , n10066 );
buf ( n10068 , n9880 );
xnor ( n10069 , n10067 , n10068 );
buf ( n10070 , n10069 );
buf ( n10071 , n10070 );
and ( n10072 , n10064 , n10071 );
and ( n10073 , n10038 , n10063 );
or ( n10074 , n10072 , n10073 );
buf ( n10075 , n10074 );
buf ( n10076 , n10075 );
not ( n10077 , n10076 );
buf ( n10078 , n10077 );
buf ( n10079 , n10078 );
nand ( n10080 , n10029 , n10079 );
buf ( n10081 , n10080 );
buf ( n10082 , n10081 );
buf ( n10083 , n10026 );
not ( n10084 , n10083 );
buf ( n10085 , n10019 );
nand ( n10086 , n10084 , n10085 );
buf ( n10087 , n10086 );
buf ( n10088 , n10087 );
nand ( n10089 , n10082 , n10088 );
buf ( n10090 , n10089 );
or ( n10091 , n10015 , n10090 );
not ( n10092 , n5695 );
not ( n10093 , n5689 );
not ( n10094 , n10093 );
not ( n10095 , n5669 );
or ( n10096 , n10094 , n10095 );
buf ( n10097 , n5613 );
and ( n10098 , n5688 , n10097 , n5586 );
nor ( n10099 , n10098 , n5814 );
buf ( n10100 , n10099 );
nand ( n10101 , n10096 , n10100 );
not ( n10102 , n10101 );
or ( n10103 , n10092 , n10102 );
not ( n10104 , n5031 );
not ( n10105 , n5172 );
or ( n10106 , n10104 , n10105 );
nand ( n10107 , n10106 , n5720 );
not ( n10108 , n10107 );
buf ( n10109 , n10108 );
not ( n10110 , n5723 );
not ( n10111 , n4646 );
not ( n10112 , n10111 );
or ( n10113 , n10110 , n10112 );
or ( n10114 , n5026 , n4868 );
nand ( n10115 , n10113 , n10114 );
not ( n10116 , n10115 );
not ( n10117 , n4646 );
not ( n10118 , n4863 );
or ( n10119 , n10117 , n10118 );
nand ( n10120 , n10119 , n5726 );
not ( n10121 , n10120 );
buf ( n10122 , n4438 );
not ( n10123 , n10122 );
buf ( n10124 , n10123 );
not ( n10125 , n10124 );
not ( n10126 , n4641 );
not ( n10127 , n10126 );
or ( n10128 , n10125 , n10127 );
nor ( n10129 , n4433 , n4230 );
and ( n10130 , n3999 , n3784 );
nor ( n10131 , n10130 , n4004 );
or ( n10132 , n3999 , n3784 );
not ( n10133 , n3596 );
not ( n10134 , n3422 );
and ( n10135 , n10133 , n10134 );
not ( n10136 , n3601 );
nor ( n10137 , n10135 , n10136 );
and ( n10138 , n5797 , n10137 );
nor ( n10139 , n10138 , n3779 );
nor ( n10140 , n10139 , n5807 );
nand ( n10141 , n10132 , n10140 );
nand ( n10142 , n10131 , n10141 );
and ( n10143 , n10142 , n4225 );
nand ( n10144 , n3999 , n3784 );
and ( n10145 , n10141 , n10144 );
not ( n10146 , n4004 );
nor ( n10147 , n10145 , n10146 );
nor ( n10148 , n10143 , n10147 );
or ( n10149 , n10129 , n10148 );
buf ( n10150 , n4433 );
buf ( n10151 , n4230 );
nand ( n10152 , n10150 , n10151 );
buf ( n10153 , n10152 );
nand ( n10154 , n10149 , n10153 );
nand ( n10155 , n10128 , n10154 );
nand ( n10156 , n10121 , n10155 );
nand ( n10157 , n10116 , n10156 );
buf ( n10158 , n10157 );
and ( n10159 , n10109 , n10158 );
not ( n10160 , n5288 );
not ( n10161 , n5177 );
and ( n10162 , n10160 , n10161 );
nor ( n10163 , n5031 , n5172 );
nor ( n10164 , n10162 , n10163 );
not ( n10165 , n10164 );
nor ( n10166 , n10159 , n10165 );
nor ( n10167 , n10166 , n5716 );
not ( n10168 , n10167 );
and ( n10169 , n5700 , n10168 );
nor ( n10170 , n10169 , n5821 );
nand ( n10171 , n10103 , n10170 );
not ( n10172 , n10171 );
not ( n10173 , n10172 );
buf ( n10174 , n10173 );
buf ( n10175 , n378 );
nand ( n10176 , n10174 , n10175 );
buf ( n10177 , n10176 );
buf ( n10178 , n10177 );
not ( n10179 , n10178 );
xor ( n10180 , n10038 , n10063 );
xor ( n10181 , n10180 , n10071 );
buf ( n10182 , n10181 );
buf ( n10183 , n10182 );
not ( n10184 , n10183 );
or ( n10185 , n10179 , n10184 );
buf ( n10186 , n9790 );
not ( n10187 , n10186 );
buf ( n10188 , n378 );
not ( n10189 , n10188 );
nand ( n10190 , n5694 , n5817 );
not ( n10191 , n10190 );
not ( n10192 , n10101 );
or ( n10193 , n10191 , n10192 );
nand ( n10194 , n10193 , n10170 );
not ( n10195 , n10194 );
buf ( n10196 , n10195 );
not ( n10197 , n10196 );
or ( n10198 , n10189 , n10197 );
buf ( n10199 , n10173 );
buf ( n10200 , n9776 );
nand ( n10201 , n10199 , n10200 );
buf ( n10202 , n10201 );
buf ( n10203 , n10202 );
nand ( n10204 , n10198 , n10203 );
buf ( n10205 , n10204 );
buf ( n10206 , n10205 );
not ( n10207 , n10206 );
or ( n10208 , n10187 , n10207 );
buf ( n10209 , n9773 );
buf ( n10210 , n378 );
nand ( n10211 , n10209 , n10210 );
buf ( n10212 , n10211 );
buf ( n10213 , n10212 );
nand ( n10214 , n10208 , n10213 );
buf ( n10215 , n10214 );
buf ( n10216 , n10215 );
not ( n10217 , n10093 );
nor ( n10218 , n5532 , n5476 );
not ( n10219 , n10218 );
not ( n10220 , n5471 );
nand ( n10221 , n10220 , n5636 );
nand ( n10222 , n10219 , n10221 , n5653 );
buf ( n10223 , n5679 );
not ( n10224 , n10223 );
buf ( n10225 , n10224 );
nor ( n10226 , n10222 , n10225 );
not ( n10227 , n10226 );
not ( n10228 , n10108 );
not ( n10229 , n10115 );
nand ( n10230 , n10229 , n10156 );
not ( n10231 , n10230 );
or ( n10232 , n10228 , n10231 );
nand ( n10233 , n10232 , n10164 );
buf ( n10234 , n5713 );
nand ( n10235 , n10233 , n10234 );
not ( n10236 , n10235 );
or ( n10237 , n10227 , n10236 );
nand ( n10238 , n10237 , n5666 );
not ( n10239 , n10238 );
or ( n10240 , n10217 , n10239 );
nand ( n10241 , n10240 , n10100 );
not ( n10242 , n5821 );
nand ( n10243 , n10242 , n5695 );
not ( n10244 , n10243 );
and ( n10245 , n10241 , n10244 );
not ( n10246 , n10241 );
and ( n10247 , n10246 , n10243 );
nor ( n10248 , n10245 , n10247 );
not ( n10249 , n10248 );
buf ( n10250 , n10249 );
not ( n10251 , n10250 );
buf ( n10252 , n378 );
nand ( n10253 , n10251 , n10252 );
buf ( n10254 , n10253 );
buf ( n10255 , n10254 );
not ( n10256 , n10255 );
buf ( n10257 , n10256 );
buf ( n10258 , n10257 );
or ( n10259 , n10216 , n10258 );
buf ( n10260 , n10061 );
buf ( n10261 , n9768 );
and ( n10262 , n10260 , n10261 );
not ( n10263 , n10260 );
not ( n10264 , n9717 );
or ( n10265 , C0 , n10264 );
nand ( n10266 , n10265 , n9726 );
not ( n10267 , n10266 );
buf ( n10268 , n10267 );
and ( n10269 , n10263 , n10268 );
nor ( n10270 , n10262 , n10269 );
buf ( n10271 , n10270 );
buf ( n10272 , n10271 );
nand ( n10273 , n10259 , n10272 );
buf ( n10274 , n10273 );
buf ( n10275 , n10274 );
buf ( n10276 , n10215 );
buf ( n10277 , n10257 );
nand ( n10278 , n10276 , n10277 );
buf ( n10279 , n10278 );
buf ( n10280 , n10279 );
nand ( n10281 , n10275 , n10280 );
buf ( n10282 , n10281 );
buf ( n10283 , n10282 );
nand ( n10284 , n10185 , n10283 );
buf ( n10285 , n10284 );
buf ( n10286 , n10177 );
not ( n10287 , n10286 );
buf ( n10288 , n10182 );
not ( n10289 , n10288 );
buf ( n10290 , n10289 );
buf ( n10291 , n10290 );
nand ( n10292 , n10287 , n10291 );
buf ( n10293 , n10292 );
nand ( n10294 , n10285 , n10293 );
not ( n10295 , n10294 );
not ( n10296 , n10022 );
not ( n10297 , n10078 );
or ( n10298 , n10296 , n10297 );
nand ( n10299 , n10075 , n10019 );
nand ( n10300 , n10298 , n10299 );
not ( n10301 , n10300 );
and ( n10302 , n10301 , n10026 );
nor ( n10303 , C0 , n10302 );
not ( n10304 , n10303 );
nand ( n10305 , n10295 , n10304 );
buf ( n10306 , n10305 );
and ( n10307 , n10091 , n10306 );
not ( n10308 , n10307 );
buf ( n10309 , n9969 );
buf ( n10310 , n378 );
buf ( n10311 , n5476 );
not ( n10312 , n10311 );
buf ( n10313 , n5532 );
buf ( n10314 , n10313 );
buf ( n10315 , n10314 );
not ( n10316 , n10315 );
and ( n10317 , n10312 , n10316 );
not ( n10318 , n10233 );
nand ( n10319 , n10318 , n5681 );
not ( n10320 , n5471 );
not ( n10321 , n5390 );
and ( n10322 , n10320 , n10321 );
buf ( n10323 , n5288 );
buf ( n10324 , n5177 );
nand ( n10325 , n10323 , n10324 );
buf ( n10326 , n10325 );
nor ( n10327 , n10322 , n10326 );
not ( n10328 , n10327 );
not ( n10329 , n5679 );
or ( n10330 , n10328 , n10329 );
nand ( n10331 , n10330 , n5646 );
nor ( n10332 , n10331 , n5660 );
and ( n10333 , n10319 , n10332 );
nor ( n10334 , n10317 , n10333 );
nand ( n10335 , n5664 , n5657 );
and ( n10336 , n10334 , n10335 );
not ( n10337 , n10334 );
not ( n10338 , n10335 );
and ( n10339 , n10337 , n10338 );
nor ( n10340 , n10336 , n10339 );
not ( n10341 , n10340 );
buf ( n10342 , n10341 );
and ( n10343 , n10310 , n10342 );
buf ( n10344 , n10343 );
buf ( n10345 , n10344 );
xor ( n10346 , n10309 , n10345 );
not ( n10347 , n9713 );
buf ( n10348 , n9367 );
not ( n10349 , n10348 );
buf ( n10350 , n10349 );
buf ( n10351 , n10350 );
not ( n10352 , n10351 );
buf ( n10353 , n10352 );
buf ( n10354 , n9692 );
buf ( n10355 , n9366 );
buf ( n10356 , n9270 );
and ( n10357 , n10354 , n10355 , n10356 );
buf ( n10358 , n10357 );
buf ( n10359 , n10358 );
not ( n10360 , n10359 );
buf ( n10361 , n9705 );
buf ( n10362 , n9366 );
nand ( n10363 , n10361 , n10362 );
buf ( n10364 , n10363 );
buf ( n10365 , n10364 );
nand ( n10366 , n10360 , n10365 );
buf ( n10367 , n10366 );
or ( n10368 , n10353 , n10367 );
not ( n10369 , n10368 );
or ( n10370 , n10347 , n10369 );
nand ( n10371 , n10370 , n9625 );
buf ( n10372 , n10371 );
buf ( n10373 , n9466 );
buf ( n10374 , n9626 );
nand ( n10375 , n10373 , n10374 );
buf ( n10376 , n10375 );
buf ( n10377 , n10376 );
not ( n10378 , n10377 );
buf ( n10379 , n10378 );
buf ( n10380 , n10379 );
and ( n10381 , n10372 , n10380 );
not ( n10382 , n10372 );
buf ( n10383 , n10376 );
and ( n10384 , n10382 , n10383 );
nor ( n10385 , n10381 , n10384 );
buf ( n10386 , n10385 );
buf ( n10387 , n10386 );
and ( n10388 , n10346 , n10387 );
and ( n10389 , n10309 , n10345 );
or ( n10390 , n10388 , n10389 );
buf ( n10391 , n10390 );
not ( n10392 , n9743 );
not ( n10393 , n380 );
not ( n10394 , n10195 );
or ( n10395 , n10393 , n10394 );
or ( n10396 , n10195 , n380 );
nand ( n10397 , n10395 , n10396 );
not ( n10398 , n10397 );
or ( n10399 , n10392 , n10398 );
nand ( n10400 , n9745 , n380 );
nand ( n10401 , n10399 , n10400 );
not ( n10402 , n10401 );
xor ( n10403 , n10391 , n10402 );
not ( n10404 , n9625 );
nor ( n10405 , n9547 , n10404 );
not ( n10406 , n10405 );
not ( n10407 , n10406 );
not ( n10408 , n10368 );
or ( n10409 , n10407 , n10408 );
not ( n10410 , n10353 );
not ( n10411 , n10367 );
nand ( n10412 , n10410 , n10411 , n10405 );
nand ( n10413 , n10409 , n10412 );
and ( n10414 , n384 , n10413 );
not ( n10415 , n10414 );
buf ( n10416 , n9743 );
not ( n10417 , n10416 );
not ( n10418 , n10241 );
not ( n10419 , n9732 );
nor ( n10420 , n10419 , n10243 );
nand ( n10421 , n10418 , n10420 );
and ( n10422 , n10243 , n380 );
nand ( n10423 , n10418 , n10422 );
and ( n10424 , n10243 , n9732 );
nand ( n10425 , n10424 , n10241 );
not ( n10426 , n380 );
nor ( n10427 , n10426 , n10243 );
nand ( n10428 , n10427 , n10241 );
nand ( n10429 , n10421 , n10423 , n10425 , n10428 );
buf ( n10430 , n10429 );
not ( n10431 , n10430 );
or ( n10432 , n10417 , n10431 );
nand ( n10433 , n10397 , n9745 );
buf ( n10434 , n10433 );
nand ( n10435 , n10432 , n10434 );
buf ( n10436 , n10435 );
not ( n10437 , n10436 );
or ( n10438 , n10415 , n10437 );
buf ( n10439 , n10436 );
buf ( n10440 , n10414 );
or ( n10441 , n10439 , n10440 );
buf ( n10442 , n9773 );
not ( n10443 , n10442 );
buf ( n10444 , n378 );
and ( n10445 , n5811 , n5688 );
not ( n10446 , n10445 );
or ( n10447 , n5827 , n10167 );
not ( n10448 , n5822 );
not ( n10449 , n5647 );
not ( n10450 , n10449 );
and ( n10451 , n10448 , n10450 );
not ( n10452 , n5586 );
not ( n10453 , n5613 );
or ( n10454 , n10452 , n10453 );
nand ( n10455 , n5665 , n5684 );
nand ( n10456 , n10454 , n10455 );
nor ( n10457 , n10451 , n10456 );
nand ( n10458 , n10447 , n10457 );
not ( n10459 , n10458 );
or ( n10460 , n10446 , n10459 );
or ( n10461 , n5827 , n10167 );
not ( n10462 , n10445 );
nand ( n10463 , n10461 , n10457 , n10462 );
nand ( n10464 , n10460 , n10463 );
not ( n10465 , n10464 );
buf ( n10466 , n10465 );
not ( n10467 , n10466 );
buf ( n10468 , n10467 );
buf ( n10469 , n10468 );
and ( n10470 , n10444 , n10469 );
not ( n10471 , n10444 );
buf ( n10472 , n10465 );
and ( n10473 , n10471 , n10472 );
nor ( n10474 , n10470 , n10473 );
buf ( n10475 , n10474 );
buf ( n10476 , n10475 );
not ( n10477 , n10476 );
buf ( n10478 , n10477 );
buf ( n10479 , n10478 );
not ( n10480 , n10479 );
or ( n10481 , n10443 , n10480 );
buf ( n10482 , n378 );
nand ( n10483 , n10097 , n5586 );
and ( n10484 , n10483 , n5684 );
xor ( n10485 , n10238 , n10484 );
buf ( n10486 , n10485 );
xor ( n10487 , n10482 , n10486 );
buf ( n10488 , n10487 );
buf ( n10489 , n10488 );
buf ( n10490 , n9790 );
nand ( n10491 , n10489 , n10490 );
buf ( n10492 , n10491 );
buf ( n10493 , n10492 );
nand ( n10494 , n10481 , n10493 );
buf ( n10495 , n10494 );
buf ( n10496 , n10495 );
nand ( n10497 , n10441 , n10496 );
buf ( n10498 , n10497 );
nand ( n10499 , n10438 , n10498 );
xnor ( n10500 , n10403 , n10499 );
buf ( n10501 , n10500 );
not ( n10502 , n5660 );
not ( n10503 , n10502 );
buf ( n10504 , n10311 );
buf ( n10505 , n10315 );
nor ( n10506 , n10504 , n10505 );
buf ( n10507 , n10506 );
nor ( n10508 , n10503 , n10507 );
not ( n10509 , n10508 );
buf ( n10510 , n5031 );
buf ( n10511 , n5172 );
nor ( n10512 , n10510 , n10511 );
buf ( n10513 , n10512 );
not ( n10514 , n10513 );
not ( n10515 , n10514 );
not ( n10516 , n10107 );
or ( n10517 , n10515 , n10516 );
not ( n10518 , n10163 );
nand ( n10519 , n10518 , n10156 , n10229 );
nand ( n10520 , n10517 , n10519 );
not ( n10521 , n10520 );
not ( n10522 , n5288 );
not ( n10523 , n5177 );
nand ( n10524 , n10522 , n10523 );
not ( n10525 , n10524 );
nor ( n10526 , n5680 , n10525 );
not ( n10527 , n10526 );
or ( n10528 , n10521 , n10527 );
not ( n10529 , n10331 );
nand ( n10530 , n10528 , n10529 );
not ( n10531 , n10530 );
not ( n10532 , n10531 );
or ( n10533 , n10509 , n10532 );
not ( n10534 , n10507 );
nand ( n10535 , n10534 , n10502 );
nand ( n10536 , n10535 , n10530 );
nand ( n10537 , n10533 , n10536 );
buf ( n10538 , n10537 );
buf ( n10539 , n378 );
nand ( n10540 , n10538 , n10539 );
buf ( n10541 , n10540 );
nand ( n10542 , n9366 , n9699 );
not ( n10543 , n10542 );
not ( n10544 , n9143 );
not ( n10545 , n8840 );
or ( n10546 , n10544 , n10545 );
buf ( n10547 , n9692 );
not ( n10548 , n10547 );
buf ( n10549 , n10548 );
nand ( n10550 , n10546 , n10549 );
not ( n10551 , n10550 );
not ( n10552 , n9270 );
or ( n10553 , n10551 , n10552 );
buf ( n10554 , n9704 );
nand ( n10555 , n10553 , n10554 );
not ( n10556 , n10555 );
or ( n10557 , n10543 , n10556 );
or ( n10558 , n10542 , n10555 );
nand ( n10559 , n10557 , n10558 );
nand ( n10560 , n10559 , n384 );
nand ( n10561 , n10541 , n10560 );
buf ( n10562 , n10561 );
not ( n10563 , n10562 );
not ( n10564 , n9773 );
not ( n10565 , n10488 );
or ( n10566 , n10564 , n10565 );
xor ( n10567 , n10310 , n10342 );
buf ( n10568 , n10567 );
nand ( n10569 , n10568 , n9790 );
nand ( n10570 , n10566 , n10569 );
buf ( n10571 , n10570 );
not ( n10572 , n10571 );
or ( n10573 , n10563 , n10572 );
not ( n10574 , n10560 );
buf ( n10575 , n10541 );
not ( n10576 , n10575 );
buf ( n10577 , n10576 );
nand ( n10578 , n10574 , n10577 );
buf ( n10579 , n10578 );
nand ( n10580 , n10573 , n10579 );
buf ( n10581 , n10580 );
buf ( n10582 , n10581 );
xor ( n10583 , n10309 , n10345 );
xor ( n10584 , n10583 , n10387 );
buf ( n10585 , n10584 );
buf ( n10586 , n10585 );
xor ( n10587 , n10582 , n10586 );
xor ( n10588 , n384 , n10413 );
buf ( n10589 , n10588 );
buf ( n10590 , n9853 );
not ( n10591 , n10590 );
not ( n10592 , n382 );
not ( n10593 , n10171 );
not ( n10594 , n10593 );
or ( n10595 , n10592 , n10594 );
or ( n10596 , n10172 , n382 );
nand ( n10597 , n10595 , n10596 );
buf ( n10598 , n10597 );
not ( n10599 , n10598 );
or ( n10600 , n10591 , n10599 );
buf ( n10601 , n9836 );
buf ( n10602 , n382 );
nand ( n10603 , n10601 , n10602 );
buf ( n10604 , n10603 );
buf ( n10605 , n10604 );
nand ( n10606 , n10600 , n10605 );
buf ( n10607 , n10606 );
buf ( n10608 , n10607 );
xor ( n10609 , n10589 , n10608 );
buf ( n10610 , n9745 );
not ( n10611 , n10610 );
buf ( n10612 , n10429 );
not ( n10613 , n10612 );
or ( n10614 , n10611 , n10613 );
buf ( n10615 , n380 );
not ( n10616 , n10615 );
buf ( n10617 , n10468 );
not ( n10618 , n10617 );
or ( n10619 , n10616 , n10618 );
not ( n10620 , n10464 );
nand ( n10621 , n10620 , n9732 );
buf ( n10622 , n10621 );
nand ( n10623 , n10619 , n10622 );
buf ( n10624 , n10623 );
buf ( n10625 , n10624 );
buf ( n10626 , n9743 );
nand ( n10627 , n10625 , n10626 );
buf ( n10628 , n10627 );
buf ( n10629 , n10628 );
nand ( n10630 , n10614 , n10629 );
buf ( n10631 , n10630 );
buf ( n10632 , n10631 );
and ( n10633 , n10609 , n10632 );
and ( n10634 , n10589 , n10608 );
or ( n10635 , n10633 , n10634 );
buf ( n10636 , n10635 );
buf ( n10637 , n10636 );
and ( n10638 , n10587 , n10637 );
and ( n10639 , n10582 , n10586 );
or ( n10640 , n10638 , n10639 );
buf ( n10641 , n10640 );
buf ( n10642 , n10641 );
or ( n10643 , n10501 , n10642 );
and ( n10644 , n10482 , n10486 );
buf ( n10645 , n10644 );
buf ( n10646 , n10645 );
buf ( n10647 , n9630 );
buf ( n10648 , n9535 );
nand ( n10649 , n10647 , n10648 );
buf ( n10650 , n10649 );
buf ( n10651 , n10650 );
buf ( n10652 , n10353 );
buf ( n10653 , n10358 );
or ( n10654 , n10652 , n10653 );
buf ( n10655 , n9713 );
buf ( n10656 , n9466 );
nand ( n10657 , n10655 , n10656 );
buf ( n10658 , n10657 );
buf ( n10659 , n10658 );
not ( n10660 , n10659 );
buf ( n10661 , n10660 );
buf ( n10662 , n10661 );
nand ( n10663 , n10654 , n10662 );
buf ( n10664 , n10663 );
buf ( n10665 , n10664 );
not ( n10666 , n10364 );
not ( n10667 , n10658 );
and ( n10668 , n10666 , n10667 );
nand ( n10669 , n9466 , n10404 );
buf ( n10670 , n10669 );
buf ( n10671 , n9626 );
nand ( n10672 , n10670 , n10671 );
buf ( n10673 , n10672 );
nor ( n10674 , n10668 , n10673 );
buf ( n10675 , n10674 );
nand ( n10676 , n10665 , n10675 );
buf ( n10677 , n10676 );
buf ( n10678 , n10677 );
or ( n10679 , n10651 , n10678 );
buf ( n10680 , n10677 );
buf ( n10681 , n10650 );
nand ( n10682 , n10680 , n10681 );
buf ( n10683 , n10682 );
buf ( n10684 , n10683 );
nand ( n10685 , n10679 , n10684 );
buf ( n10686 , n10685 );
buf ( n10687 , n10686 );
buf ( n10688 , n10033 );
xnor ( n10689 , n10687 , n10688 );
buf ( n10690 , n10689 );
buf ( n10691 , n10690 );
xor ( n10692 , n10646 , n10691 );
not ( n10693 , n9773 );
buf ( n10694 , n378 );
not ( n10695 , n10694 );
buf ( n10696 , n10249 );
not ( n10697 , n10696 );
or ( n10698 , n10695 , n10697 );
not ( n10699 , n10244 );
not ( n10700 , n10418 );
or ( n10701 , n10699 , n10700 );
nand ( n10702 , n10243 , n10241 );
nand ( n10703 , n10701 , n10702 );
nand ( n10704 , n10703 , n9776 );
buf ( n10705 , n10704 );
nand ( n10706 , n10698 , n10705 );
buf ( n10707 , n10706 );
not ( n10708 , n10707 );
or ( n10709 , n10693 , n10708 );
or ( n10710 , n10475 , n9793 );
nand ( n10711 , n10709 , n10710 );
buf ( n10712 , n10711 );
xor ( n10713 , n10692 , n10712 );
buf ( n10714 , n10713 );
buf ( n10715 , n10714 );
nand ( n10716 , n10643 , n10715 );
buf ( n10717 , n10716 );
buf ( n10718 , n10717 );
buf ( n10719 , n10641 );
buf ( n10720 , n10500 );
nand ( n10721 , n10719 , n10720 );
buf ( n10722 , n10721 );
buf ( n10723 , n10722 );
nand ( n10724 , n10718 , n10723 );
buf ( n10725 , n10724 );
buf ( n10726 , n10725 );
not ( n10727 , n10726 );
and ( n10728 , n10465 , n378 );
not ( n10729 , n10728 );
xor ( n10730 , n10056 , n10729 );
buf ( n10731 , n9654 );
buf ( n10732 , n9584 );
nand ( n10733 , n10731 , n10732 );
buf ( n10734 , n10733 );
buf ( n10735 , n10734 );
not ( n10736 , n10735 );
not ( n10737 , n9535 );
not ( n10738 , n10677 );
or ( n10739 , n10737 , n10738 );
nand ( n10740 , n10739 , n9630 );
buf ( n10741 , n10740 );
not ( n10742 , n10741 );
or ( n10743 , n10736 , n10742 );
buf ( n10744 , n10740 );
buf ( n10745 , n10734 );
or ( n10746 , n10744 , n10745 );
nand ( n10747 , n10743 , n10746 );
buf ( n10748 , n10747 );
xnor ( n10749 , n10730 , n10748 );
not ( n10750 , n10401 );
not ( n10751 , n10391 );
or ( n10752 , n10750 , n10751 );
not ( n10753 , n10402 );
not ( n10754 , n10391 );
not ( n10755 , n10754 );
or ( n10756 , n10753 , n10755 );
nand ( n10757 , n10756 , n10499 );
nand ( n10758 , n10752 , n10757 );
xor ( n10759 , n10749 , n10758 );
buf ( n10760 , n9790 );
not ( n10761 , n10760 );
buf ( n10762 , n10707 );
not ( n10763 , n10762 );
or ( n10764 , n10761 , n10763 );
buf ( n10765 , n10205 );
buf ( n10766 , n9773 );
nand ( n10767 , n10765 , n10766 );
buf ( n10768 , n10767 );
buf ( n10769 , n10768 );
nand ( n10770 , n10764 , n10769 );
buf ( n10771 , n10770 );
buf ( n10772 , n10771 );
not ( n10773 , n10772 );
buf ( n10774 , n10033 );
not ( n10775 , n10774 );
buf ( n10776 , n10686 );
nand ( n10777 , n10775 , n10776 );
buf ( n10778 , n10777 );
buf ( n10779 , n10778 );
not ( n10780 , n10779 );
and ( n10781 , n10773 , n10780 );
buf ( n10782 , n10771 );
buf ( n10783 , n10778 );
and ( n10784 , n10782 , n10783 );
nor ( n10785 , n10781 , n10784 );
buf ( n10786 , n10785 );
xor ( n10787 , n10646 , n10691 );
and ( n10788 , n10787 , n10712 );
and ( n10789 , n10646 , n10691 );
or ( n10790 , n10788 , n10789 );
buf ( n10791 , n10790 );
xor ( n10792 , n10786 , n10791 );
xnor ( n10793 , n10759 , n10792 );
buf ( n10794 , n10793 );
not ( n10795 , n10794 );
buf ( n10796 , n10795 );
buf ( n10797 , n10796 );
nand ( n10798 , n10727 , n10797 );
buf ( n10799 , n10798 );
buf ( n10800 , n10177 );
buf ( n10801 , n10290 );
xor ( n10802 , n10800 , n10801 );
buf ( n10803 , n10282 );
xor ( n10804 , n10802 , n10803 );
buf ( n10805 , n10804 );
or ( n10806 , n10056 , n10748 );
nand ( n10807 , n10806 , n10728 );
nand ( n10808 , n10748 , n10056 );
nand ( n10809 , n10807 , n10808 );
buf ( n10810 , n10809 );
not ( n10811 , n10810 );
buf ( n10812 , n10811 );
not ( n10813 , n10812 );
buf ( n10814 , n10771 );
not ( n10815 , n10814 );
buf ( n10816 , n10778 );
nand ( n10817 , n10815 , n10816 );
buf ( n10818 , n10817 );
buf ( n10819 , n10818 );
not ( n10820 , n10819 );
buf ( n10821 , n10791 );
not ( n10822 , n10821 );
or ( n10823 , n10820 , n10822 );
buf ( n10824 , n10778 );
not ( n10825 , n10824 );
buf ( n10826 , n10771 );
nand ( n10827 , n10825 , n10826 );
buf ( n10828 , n10827 );
buf ( n10829 , n10828 );
nand ( n10830 , n10823 , n10829 );
buf ( n10831 , n10830 );
buf ( n10832 , n10831 );
not ( n10833 , n10832 );
buf ( n10834 , n10833 );
not ( n10835 , n10834 );
or ( n10836 , n10813 , n10835 );
xor ( n10837 , n10271 , n10254 );
xor ( n10838 , n10837 , n10215 );
not ( n10839 , n10838 );
nand ( n10840 , n10836 , n10839 );
nand ( n10841 , n10831 , n10809 );
nand ( n10842 , n10805 , n10840 , n10841 );
nand ( n10843 , n10799 , n10842 );
not ( n10844 , n10838 );
not ( n10845 , n10809 );
or ( n10846 , n10844 , n10845 );
or ( n10847 , n10838 , n10809 );
nand ( n10848 , n10846 , n10847 );
xor ( n10849 , n10831 , n10848 );
buf ( n10850 , n10849 );
not ( n10851 , n10850 );
buf ( n10852 , n10851 );
not ( n10853 , n10792 );
not ( n10854 , n10853 );
not ( n10855 , n10749 );
not ( n10856 , n10758 );
nand ( n10857 , n10855 , n10856 );
not ( n10858 , n10857 );
or ( n10859 , n10854 , n10858 );
not ( n10860 , n10856 );
nand ( n10861 , n10860 , n10749 );
nand ( n10862 , n10859 , n10861 );
not ( n10863 , n10862 );
nand ( n10864 , n10852 , n10863 );
buf ( n10865 , n10864 );
buf ( n10866 , n10414 );
buf ( n10867 , n10495 );
xor ( n10868 , n10866 , n10867 );
buf ( n10869 , n10436 );
xnor ( n10870 , n10868 , n10869 );
buf ( n10871 , n10870 );
buf ( n10872 , n10871 );
not ( n10873 , n10872 );
buf ( n10874 , n10235 );
buf ( n10875 , n5709 );
xor ( n10876 , n10874 , n10875 );
buf ( n10877 , n10876 );
buf ( n10878 , n10877 );
not ( n10879 , n10878 );
buf ( n10880 , n10879 );
buf ( n10881 , n10880 );
not ( n10882 , n10881 );
buf ( n10883 , n10882 );
buf ( n10884 , n9704 );
buf ( n10885 , n9270 );
nand ( n10886 , n10884 , n10885 );
buf ( n10887 , n10886 );
xnor ( n10888 , n10550 , n10887 );
nand ( n10889 , n378 , n10883 , n10888 );
buf ( n10890 , n10889 );
not ( n10891 , n10890 );
buf ( n10892 , n10891 );
buf ( n10893 , n10892 );
not ( n10894 , n10893 );
and ( n10895 , n9853 , n382 );
and ( n10896 , n10249 , n10895 );
and ( n10897 , n10597 , n9836 );
nor ( n10898 , n10896 , n10897 );
nand ( n10899 , n10703 , n9738 , n9853 );
nand ( n10900 , n10898 , n10899 );
buf ( n10901 , n10900 );
not ( n10902 , n10901 );
or ( n10903 , n10894 , n10902 );
buf ( n10904 , n10900 );
buf ( n10905 , n10892 );
or ( n10906 , n10904 , n10905 );
buf ( n10907 , n9745 );
not ( n10908 , n10907 );
buf ( n10909 , n10624 );
not ( n10910 , n10909 );
or ( n10911 , n10908 , n10910 );
buf ( n10912 , n10485 );
not ( n10913 , n10912 );
buf ( n10914 , n10913 );
nand ( n10915 , n380 , n10914 );
not ( n10916 , n10915 );
not ( n10917 , n380 );
nand ( n10918 , n10917 , n10485 );
not ( n10919 , n10918 );
or ( n10920 , n10916 , n10919 );
nand ( n10921 , n10920 , n9743 );
buf ( n10922 , n10921 );
nand ( n10923 , n10911 , n10922 );
buf ( n10924 , n10923 );
buf ( n10925 , n10924 );
nand ( n10926 , n10906 , n10925 );
buf ( n10927 , n10926 );
buf ( n10928 , n10927 );
nand ( n10929 , n10903 , n10928 );
buf ( n10930 , n10929 );
buf ( n10931 , n10930 );
not ( n10932 , n10931 );
not ( n10933 , n10570 );
not ( n10934 , n10933 );
and ( n10935 , n10560 , n10577 );
not ( n10936 , n10560 );
and ( n10937 , n10936 , n10541 );
nor ( n10938 , n10935 , n10937 );
not ( n10939 , n10938 );
not ( n10940 , n10939 );
or ( n10941 , n10934 , n10940 );
nand ( n10942 , n10938 , n10570 );
nand ( n10943 , n10941 , n10942 );
buf ( n10944 , n10943 );
buf ( n10945 , n10944 );
buf ( n10946 , n10945 );
buf ( n10947 , n10946 );
not ( n10948 , n10947 );
buf ( n10949 , n10948 );
buf ( n10950 , n10949 );
and ( n10951 , n10524 , n5679 );
not ( n10952 , n10951 );
not ( n10953 , n10520 );
or ( n10954 , n10952 , n10953 );
not ( n10955 , n10225 );
not ( n10956 , n5713 );
and ( n10957 , n10955 , n10956 );
nor ( n10958 , n10957 , n5712 );
nand ( n10959 , n10954 , n10958 );
buf ( n10960 , n10959 );
buf ( n10961 , n10221 );
buf ( n10962 , n5831 );
nand ( n10963 , n10961 , n10962 );
buf ( n10964 , n10963 );
buf ( n10965 , n10964 );
not ( n10966 , n10965 );
buf ( n10967 , n10966 );
buf ( n10968 , n10967 );
and ( n10969 , n10960 , n10968 );
not ( n10970 , n10960 );
buf ( n10971 , n10964 );
and ( n10972 , n10970 , n10971 );
nor ( n10973 , n10969 , n10972 );
buf ( n10974 , n10973 );
buf ( n10975 , n10974 );
not ( n10976 , n10975 );
buf ( n10977 , n10976 );
buf ( n10978 , n10977 );
not ( n10979 , n10978 );
buf ( n10980 , n10979 );
buf ( n10981 , n10980 );
buf ( n10982 , n378 );
nand ( n10983 , n10981 , n10982 );
buf ( n10984 , n10983 );
xor ( n10985 , n384 , n10542 );
xor ( n10986 , n10985 , n10555 );
nand ( n10987 , n10984 , n10986 );
not ( n10988 , n10987 );
buf ( n10989 , n9773 );
not ( n10990 , n10989 );
buf ( n10991 , n10568 );
not ( n10992 , n10991 );
or ( n10993 , n10990 , n10992 );
and ( n10994 , n10535 , n9776 );
not ( n10995 , n10535 );
and ( n10996 , n10995 , n378 );
nor ( n10997 , n10994 , n10996 );
buf ( n10998 , n10531 );
not ( n10999 , n10998 );
and ( n11000 , n10997 , n10999 );
not ( n11001 , n10997 );
and ( n11002 , n11001 , n10998 );
nor ( n11003 , n11000 , n11002 );
nand ( n11004 , n11003 , n9790 );
buf ( n11005 , n11004 );
nand ( n11006 , n10993 , n11005 );
buf ( n11007 , n11006 );
not ( n11008 , n11007 );
or ( n11009 , n10988 , n11008 );
or ( n11010 , n10986 , n10984 );
nand ( n11011 , n11009 , n11010 );
not ( n11012 , n11011 );
buf ( n11013 , n11012 );
nand ( n11014 , n10950 , n11013 );
buf ( n11015 , n11014 );
buf ( n11016 , n11015 );
not ( n11017 , n11016 );
or ( n11018 , n10932 , n11017 );
not ( n11019 , n10987 );
not ( n11020 , n11007 );
or ( n11021 , n11019 , n11020 );
nand ( n11022 , n11021 , n11010 );
nand ( n11023 , n10946 , n11022 );
buf ( n11024 , n11023 );
nand ( n11025 , n11018 , n11024 );
buf ( n11026 , n11025 );
buf ( n11027 , n11026 );
not ( n11028 , n11027 );
buf ( n11029 , n11028 );
buf ( n11030 , n11029 );
not ( n11031 , n11030 );
or ( n11032 , n10873 , n11031 );
xor ( n11033 , n10582 , n10586 );
xor ( n11034 , n11033 , n10637 );
buf ( n11035 , n11034 );
buf ( n11036 , n11035 );
buf ( n11037 , n11036 );
buf ( n11038 , n11037 );
buf ( n11039 , n11038 );
nand ( n11040 , n11032 , n11039 );
buf ( n11041 , n11040 );
buf ( n11042 , n11041 );
buf ( n11043 , n10871 );
not ( n11044 , n11043 );
buf ( n11045 , n11026 );
nand ( n11046 , n11044 , n11045 );
buf ( n11047 , n11046 );
buf ( n11048 , n11047 );
and ( n11049 , n11042 , n11048 );
buf ( n11050 , n11049 );
buf ( n11051 , n10714 );
buf ( n11052 , n10641 );
xor ( n11053 , n11051 , n11052 );
buf ( n11054 , n10500 );
xnor ( n11055 , n11053 , n11054 );
buf ( n11056 , n11055 );
nand ( n11057 , n11050 , n11056 );
buf ( n11058 , n11057 );
nand ( n11059 , n10865 , n11058 );
buf ( n11060 , n11059 );
nor ( n11061 , n10843 , n11060 );
not ( n11062 , n11061 );
xor ( n11063 , n10889 , n10924 );
xnor ( n11064 , n11063 , n10900 );
nand ( n11065 , n10524 , n5713 );
not ( n11066 , n11065 );
not ( n11067 , n11066 );
not ( n11068 , n10520 );
not ( n11069 , n11068 );
or ( n11070 , n11067 , n11069 );
nand ( n11071 , n10520 , n11065 );
nand ( n11072 , n11070 , n11071 );
buf ( n11073 , n11072 );
buf ( n11074 , n378 );
and ( n11075 , n11073 , n11074 );
buf ( n11076 , n11075 );
buf ( n11077 , n11076 );
and ( n11078 , n9689 , n9095 );
buf ( n11079 , n9140 );
not ( n11080 , n11079 );
buf ( n11081 , n8840 );
buf ( n11082 , n11081 );
buf ( n11083 , n11082 );
buf ( n11084 , n11083 );
not ( n11085 , n11084 );
or ( n11086 , n11080 , n11085 );
buf ( n11087 , n9673 );
buf ( n11088 , n11087 );
buf ( n11089 , n11088 );
buf ( n11090 , n11089 );
nand ( n11091 , n11086 , n11090 );
buf ( n11092 , n11091 );
xor ( n11093 , n11078 , n11092 );
buf ( n11094 , n11093 );
xor ( n11095 , n11077 , n11094 );
and ( n11096 , n11089 , n9140 );
xor ( n11097 , n11096 , n11083 );
nand ( n11098 , n2967 , n2984 , n3025 );
and ( n11099 , n11097 , n11098 );
buf ( n11100 , n11099 );
xor ( n11101 , n11095 , n11100 );
buf ( n11102 , n11101 );
buf ( n11103 , n11102 );
buf ( n11104 , n9836 );
not ( n11105 , n11104 );
not ( n11106 , n382 );
not ( n11107 , n10468 );
or ( n11108 , n11106 , n11107 );
nand ( n11109 , n10465 , n9738 );
nand ( n11110 , n11108 , n11109 );
buf ( n11111 , n11110 );
not ( n11112 , n11111 );
or ( n11113 , n11105 , n11112 );
buf ( n11114 , n382 );
buf ( n11115 , n10914 );
and ( n11116 , n11114 , n11115 );
not ( n11117 , n11114 );
buf ( n11118 , n10485 );
and ( n11119 , n11117 , n11118 );
nor ( n11120 , n11116 , n11119 );
buf ( n11121 , n11120 );
not ( n11122 , n11121 );
nand ( n11123 , n11122 , n9853 );
buf ( n11124 , n11123 );
nand ( n11125 , n11113 , n11124 );
buf ( n11126 , n11125 );
buf ( n11127 , n11126 );
xor ( n11128 , n11103 , n11127 );
buf ( n11129 , n9790 );
not ( n11130 , n11129 );
buf ( n11131 , n378 );
buf ( n11132 , n11072 );
and ( n11133 , n11131 , n11132 );
not ( n11134 , n11131 );
buf ( n11135 , n11072 );
not ( n11136 , n11135 );
buf ( n11137 , n11136 );
buf ( n11138 , n11137 );
and ( n11139 , n11134 , n11138 );
nor ( n11140 , n11133 , n11139 );
buf ( n11141 , n11140 );
buf ( n11142 , n11141 );
not ( n11143 , n11142 );
or ( n11144 , n11130 , n11143 );
buf ( n11145 , n378 );
not ( n11146 , n11145 );
buf ( n11147 , n10880 );
not ( n11148 , n11147 );
or ( n11149 , n11146 , n11148 );
buf ( n11150 , n9776 );
buf ( n11151 , n10877 );
nand ( n11152 , n11150 , n11151 );
buf ( n11153 , n11152 );
buf ( n11154 , n11153 );
nand ( n11155 , n11149 , n11154 );
buf ( n11156 , n11155 );
buf ( n11157 , n11156 );
buf ( n11158 , n9773 );
nand ( n11159 , n11157 , n11158 );
buf ( n11160 , n11159 );
buf ( n11161 , n11160 );
nand ( n11162 , n11144 , n11161 );
buf ( n11163 , n11162 );
not ( n11164 , n11163 );
buf ( n11165 , n380 );
not ( n11166 , n11165 );
buf ( n11167 , n10537 );
not ( n11168 , n11167 );
buf ( n11169 , n11168 );
buf ( n11170 , n11169 );
not ( n11171 , n11170 );
or ( n11172 , n11166 , n11171 );
buf ( n11173 , n10537 );
buf ( n11174 , n9732 );
nand ( n11175 , n11173 , n11174 );
buf ( n11176 , n11175 );
buf ( n11177 , n11176 );
nand ( n11178 , n11172 , n11177 );
buf ( n11179 , n11178 );
nand ( n11180 , n11179 , n9745 );
not ( n11181 , n9732 );
and ( n11182 , n10959 , n10964 );
not ( n11183 , n10959 );
and ( n11184 , n11183 , n10967 );
nor ( n11185 , n11182 , n11184 );
not ( n11186 , n11185 );
not ( n11187 , n11186 );
or ( n11188 , n11181 , n11187 );
or ( n11189 , n9732 , n11186 );
nand ( n11190 , n11188 , n11189 );
nand ( n11191 , n11190 , n9743 );
nand ( n11192 , n11164 , n11180 , n11191 );
not ( n11193 , n11192 );
buf ( n11194 , n382 );
not ( n11195 , n11194 );
buf ( n11196 , n10340 );
not ( n11197 , n11196 );
or ( n11198 , n11195 , n11197 );
buf ( n11199 , n10341 );
buf ( n11200 , n9738 );
nand ( n11201 , n11199 , n11200 );
buf ( n11202 , n11201 );
buf ( n11203 , n11202 );
nand ( n11204 , n11198 , n11203 );
buf ( n11205 , n11204 );
not ( n11206 , n11205 );
not ( n11207 , n9853 );
or ( n11208 , n11206 , n11207 );
or ( n11209 , n11121 , n9839 );
nand ( n11210 , n11208 , n11209 );
not ( n11211 , n11210 );
or ( n11212 , n11193 , n11211 );
not ( n11213 , n11191 );
not ( n11214 , n11180 );
or ( n11215 , n11213 , n11214 );
nand ( n11216 , n11215 , n11163 );
nand ( n11217 , n11212 , n11216 );
buf ( n11218 , n11217 );
and ( n11219 , n11128 , n11218 );
and ( n11220 , n11103 , n11127 );
or ( n11221 , n11219 , n11220 );
buf ( n11222 , n11221 );
not ( n11223 , n11222 );
nand ( n11224 , n10883 , n378 );
not ( n11225 , n10888 );
and ( n11226 , n11224 , n11225 );
not ( n11227 , n11224 );
and ( n11228 , n11227 , n10888 );
nor ( n11229 , n11226 , n11228 );
not ( n11230 , n9790 );
not ( n11231 , n378 );
not ( n11232 , n11185 );
or ( n11233 , n11231 , n11232 );
buf ( n11234 , n10974 );
buf ( n11235 , n9776 );
nand ( n11236 , n11234 , n11235 );
buf ( n11237 , n11236 );
nand ( n11238 , n11233 , n11237 );
not ( n11239 , n11238 );
or ( n11240 , n11230 , n11239 );
nand ( n11241 , n11003 , n9773 );
nand ( n11242 , n11240 , n11241 );
xor ( n11243 , n11229 , n11242 );
xor ( n11244 , n10335 , n380 );
not ( n11245 , n10311 );
not ( n11246 , n10315 );
and ( n11247 , n11245 , n11246 );
and ( n11248 , n10319 , n10332 );
nor ( n11249 , n11247 , n11248 );
xnor ( n11250 , n11244 , n11249 );
not ( n11251 , n11250 );
not ( n11252 , n9743 );
or ( n11253 , n11251 , n11252 );
not ( n11254 , n10915 );
not ( n11255 , n10918 );
or ( n11256 , n11254 , n11255 );
nand ( n11257 , n11256 , n9745 );
nand ( n11258 , n11253 , n11257 );
xor ( n11259 , n11243 , n11258 );
not ( n11260 , n11259 );
not ( n11261 , n11179 );
not ( n11262 , n9743 );
or ( n11263 , n11261 , n11262 );
nand ( n11264 , n11250 , n9745 );
nand ( n11265 , n11263 , n11264 );
not ( n11266 , n11265 );
nand ( n11267 , n10157 , n5720 );
not ( n11268 , n11267 );
not ( n11269 , n10513 );
nand ( n11270 , n5172 , n5031 );
nand ( n11271 , n11269 , n11270 );
not ( n11272 , n11271 );
or ( n11273 , n11268 , n11272 );
not ( n11274 , n11267 );
not ( n11275 , n11270 );
nor ( n11276 , n11275 , n10513 );
nand ( n11277 , n11274 , n11276 );
nand ( n11278 , n11273 , n11277 );
and ( n11279 , n378 , n11278 );
not ( n11280 , n11279 );
not ( n11281 , n11280 );
buf ( n11282 , n8620 );
buf ( n11283 , n11282 );
buf ( n11284 , n11283 );
buf ( n11285 , n11284 );
not ( n11286 , n11285 );
buf ( n11287 , n8642 );
not ( n11288 , n11287 );
buf ( n11289 , n11288 );
buf ( n11290 , n11289 );
not ( n11291 , n11290 );
buf ( n11292 , n8212 );
not ( n11293 , n11292 );
or ( n11294 , n11291 , n11293 );
buf ( n11295 , n8814 );
not ( n11296 , n11295 );
buf ( n11297 , n11296 );
buf ( n11298 , n11297 );
nand ( n11299 , n11294 , n11298 );
buf ( n11300 , n11299 );
buf ( n11301 , n11300 );
not ( n11302 , n11301 );
or ( n11303 , n11286 , n11302 );
buf ( n11304 , n8810 );
not ( n11305 , n11304 );
buf ( n11306 , n11305 );
buf ( n11307 , n11306 );
not ( n11308 , n11307 );
buf ( n11309 , n11308 );
buf ( n11310 , n11309 );
nand ( n11311 , n11303 , n11310 );
buf ( n11312 , n11311 );
buf ( n11313 , n8833 );
buf ( n11314 , n8800 );
nand ( n11315 , n11313 , n11314 );
buf ( n11316 , n11315 );
not ( n11317 , n11316 );
and ( n11318 , n11312 , n11317 );
not ( n11319 , n11312 );
and ( n11320 , n11319 , n11316 );
nor ( n11321 , n11318 , n11320 );
nand ( n11322 , n5723 , n10111 );
not ( n11323 , n11322 );
not ( n11324 , n10120 );
or ( n11325 , n11323 , n11324 );
nand ( n11326 , n5724 , n10154 , n11322 );
nand ( n11327 , n11325 , n11326 );
not ( n11328 , n4868 );
not ( n11329 , n11328 );
not ( n11330 , n5026 );
not ( n11331 , n11330 );
or ( n11332 , n11329 , n11331 );
nand ( n11333 , n11332 , n5720 );
not ( n11334 , n11333 );
and ( n11335 , n11327 , n11334 );
not ( n11336 , n11327 );
not ( n11337 , n11328 );
not ( n11338 , n11330 );
or ( n11339 , n11337 , n11338 );
nand ( n11340 , n11339 , n5720 );
and ( n11341 , n11336 , n11340 );
nor ( n11342 , n11335 , n11341 );
nand ( n11343 , n11342 , n378 );
not ( n11344 , n11343 );
nand ( n11345 , n11321 , n11344 );
not ( n11346 , n11345 );
or ( n11347 , n11281 , n11346 );
xor ( n11348 , n11097 , n11098 );
nand ( n11349 , n11347 , n11348 );
not ( n11350 , n11345 );
nand ( n11351 , n11350 , n11279 );
nand ( n11352 , n11349 , n11351 );
not ( n11353 , n11352 );
not ( n11354 , n9773 );
not ( n11355 , n11238 );
or ( n11356 , n11354 , n11355 );
nand ( n11357 , n11156 , n9790 );
nand ( n11358 , n11356 , n11357 );
not ( n11359 , n11358 );
nand ( n11360 , n11353 , n11359 );
not ( n11361 , n11360 );
or ( n11362 , n11266 , n11361 );
nand ( n11363 , n11358 , n11352 );
nand ( n11364 , n11362 , n11363 );
buf ( n11365 , n11364 );
not ( n11366 , n11365 );
buf ( n11367 , n11366 );
nand ( n11368 , n11260 , n11367 );
not ( n11369 , n11368 );
or ( n11370 , n11223 , n11369 );
buf ( n11371 , n11260 );
not ( n11372 , n11371 );
buf ( n11373 , n11372 );
buf ( n11374 , n11373 );
buf ( n11375 , n11364 );
nand ( n11376 , n11374 , n11375 );
buf ( n11377 , n11376 );
nand ( n11378 , n11370 , n11377 );
xor ( n11379 , n11064 , n11378 );
xor ( n11380 , n11229 , n11242 );
and ( n11381 , n11380 , n11258 );
and ( n11382 , n11229 , n11242 );
or ( n11383 , n11381 , n11382 );
buf ( n11384 , n11383 );
not ( n11385 , n11384 );
buf ( n11386 , n10984 );
buf ( n11387 , n10986 );
xor ( n11388 , n11386 , n11387 );
buf ( n11389 , n11007 );
xnor ( n11390 , n11388 , n11389 );
buf ( n11391 , n11390 );
buf ( n11392 , n11391 );
not ( n11393 , n11392 );
or ( n11394 , n11385 , n11393 );
buf ( n11395 , n11391 );
buf ( n11396 , n11383 );
or ( n11397 , n11395 , n11396 );
nand ( n11398 , n11394 , n11397 );
buf ( n11399 , n11398 );
not ( n11400 , n9853 );
not ( n11401 , n11110 );
or ( n11402 , n11400 , n11401 );
xor ( n11403 , n10243 , n382 );
xnor ( n11404 , n11403 , n10241 );
nand ( n11405 , n11404 , n9836 );
nand ( n11406 , n11402 , n11405 );
not ( n11407 , n11406 );
not ( n11408 , n385 );
and ( n11409 , n11408 , n384 );
buf ( n11410 , n11409 );
not ( n11411 , n11410 );
buf ( n11412 , n10195 );
not ( n11413 , n11412 );
or ( n11414 , n11411 , n11413 );
buf ( n11415 , n384 );
buf ( n11416 , n385 );
nand ( n11417 , n11415 , n11416 );
buf ( n11418 , n11417 );
buf ( n11419 , n11418 );
nand ( n11420 , n11414 , n11419 );
buf ( n11421 , n11420 );
not ( n11422 , n11421 );
or ( n11423 , n11407 , n11422 );
buf ( n11424 , n11421 );
not ( n11425 , n11424 );
buf ( n11426 , n11425 );
nand ( n11427 , n9853 , n11110 );
and ( n11428 , n11426 , n11427 , n11405 );
xor ( n11429 , n11077 , n11094 );
and ( n11430 , n11429 , n11100 );
and ( n11431 , n11077 , n11094 );
or ( n11432 , n11430 , n11431 );
buf ( n11433 , n11432 );
buf ( n11434 , n11433 );
not ( n11435 , n11434 );
buf ( n11436 , n11435 );
or ( n11437 , n11428 , n11436 );
nand ( n11438 , n11423 , n11437 );
and ( n11439 , n11399 , n11438 );
not ( n11440 , n11399 );
not ( n11441 , n11438 );
and ( n11442 , n11440 , n11441 );
nor ( n11443 , n11439 , n11442 );
xor ( n11444 , n11379 , n11443 );
buf ( n11445 , n11444 );
not ( n11446 , n11445 );
buf ( n11447 , n11446 );
and ( n11448 , n11436 , n11426 );
not ( n11449 , n11436 );
and ( n11450 , n11449 , n11421 );
nor ( n11451 , n11448 , n11450 );
not ( n11452 , n11451 );
not ( n11453 , n11406 );
and ( n11454 , n11452 , n11453 );
and ( n11455 , n11451 , n11406 );
nor ( n11456 , n11454 , n11455 );
buf ( n11457 , n11409 );
not ( n11458 , n11457 );
and ( n11459 , n384 , n10249 );
not ( n11460 , n384 );
and ( n11461 , n11460 , n10248 );
or ( n11462 , n11459 , n11461 );
buf ( n11463 , n11462 );
not ( n11464 , n11463 );
or ( n11465 , n11458 , n11464 );
buf ( n11466 , n384 );
buf ( n11467 , n10173 );
and ( n11468 , n11466 , n11467 );
not ( n11469 , n11466 );
buf ( n11470 , n10195 );
and ( n11471 , n11469 , n11470 );
nor ( n11472 , n11468 , n11471 );
buf ( n11473 , n11472 );
buf ( n11474 , n11473 );
buf ( n11475 , n385 );
nand ( n11476 , n11474 , n11475 );
buf ( n11477 , n11476 );
buf ( n11478 , n11477 );
nand ( n11479 , n11465 , n11478 );
buf ( n11480 , n11479 );
not ( n11481 , n11480 );
and ( n11482 , n11358 , n11352 );
not ( n11483 , n11358 );
and ( n11484 , n11483 , n11353 );
nor ( n11485 , n11482 , n11484 );
not ( n11486 , n11265 );
and ( n11487 , n11485 , n11486 );
not ( n11488 , n11485 );
and ( n11489 , n11488 , n11265 );
nor ( n11490 , n11487 , n11489 );
buf ( n11491 , n11490 );
not ( n11492 , n11491 );
buf ( n11493 , n11492 );
not ( n11494 , n11493 );
or ( n11495 , n11481 , n11494 );
buf ( n11496 , n11493 );
buf ( n11497 , n11480 );
or ( n11498 , n11496 , n11497 );
xor ( n11499 , n11280 , n11350 );
xnor ( n11500 , n11499 , n11348 );
not ( n11501 , n11500 );
buf ( n11502 , n11306 );
not ( n11503 , n11502 );
buf ( n11504 , n11284 );
nand ( n11505 , n11503 , n11504 );
buf ( n11506 , n11505 );
xnor ( n11507 , n11300 , n11506 );
buf ( n11508 , n11507 );
nand ( n11509 , n10155 , n5727 );
not ( n11510 , n4646 );
not ( n11511 , n4863 );
or ( n11512 , n11510 , n11511 );
nand ( n11513 , n11512 , n11322 );
not ( n11514 , n11513 );
and ( n11515 , n11509 , n11514 );
not ( n11516 , n11509 );
and ( n11517 , n11516 , n11513 );
nor ( n11518 , n11515 , n11517 );
and ( n11519 , n11518 , n378 );
buf ( n11520 , n11519 );
and ( n11521 , n11508 , n11520 );
buf ( n11522 , n11521 );
buf ( n11523 , n11522 );
not ( n11524 , n11523 );
nand ( n11525 , n3018 , n1007 );
not ( n11526 , n11525 );
nand ( n11527 , n2980 , n3029 );
nand ( n11528 , n11527 , n2782 );
not ( n11529 , n11528 );
or ( n11530 , n11526 , n11529 );
not ( n11531 , n11525 );
nand ( n11532 , n11531 , n2782 , n11527 );
nand ( n11533 , n11530 , n11532 );
buf ( n11534 , n11533 );
not ( n11535 , n11534 );
or ( n11536 , n11524 , n11535 );
not ( n11537 , n11522 );
not ( n11538 , n11537 );
not ( n11539 , n11533 );
not ( n11540 , n11539 );
or ( n11541 , n11538 , n11540 );
buf ( n11542 , n11321 );
buf ( n11543 , n11343 );
and ( n11544 , n11542 , n11543 );
not ( n11545 , n11542 );
buf ( n11546 , n11344 );
and ( n11547 , n11545 , n11546 );
nor ( n11548 , n11544 , n11547 );
buf ( n11549 , n11548 );
buf ( n11550 , n11549 );
not ( n11551 , n11550 );
buf ( n11552 , n11551 );
nand ( n11553 , n11541 , n11552 );
buf ( n11554 , n11553 );
nand ( n11555 , n11536 , n11554 );
buf ( n11556 , n11555 );
buf ( n11557 , n11556 );
not ( n11558 , n11557 );
buf ( n11559 , n11558 );
nand ( n11560 , n11501 , n11559 );
not ( n11561 , n11560 );
not ( n11562 , n9773 );
not ( n11563 , n11141 );
or ( n11564 , n11562 , n11563 );
xor ( n11565 , n378 , n11278 );
buf ( n11566 , n11565 );
buf ( n11567 , n9790 );
nand ( n11568 , n11566 , n11567 );
buf ( n11569 , n11568 );
nand ( n11570 , n11564 , n11569 );
not ( n11571 , n11570 );
not ( n11572 , n11571 );
buf ( n11573 , n9773 );
not ( n11574 , n11573 );
buf ( n11575 , n11565 );
not ( n11576 , n11575 );
or ( n11577 , n11574 , n11576 );
xor ( n11578 , n378 , n11340 );
xnor ( n11579 , n11578 , n11327 );
buf ( n11580 , n11579 );
buf ( n11581 , n9790 );
nand ( n11582 , n11580 , n11581 );
buf ( n11583 , n11582 );
buf ( n11584 , n11583 );
nand ( n11585 , n11577 , n11584 );
buf ( n11586 , n11585 );
not ( n11587 , n11586 );
buf ( n11588 , n11519 );
buf ( n11589 , n11507 );
not ( n11590 , n11589 );
buf ( n11591 , n11590 );
buf ( n11592 , n11591 );
and ( n11593 , n11588 , n11592 );
not ( n11594 , n11588 );
buf ( n11595 , n11507 );
and ( n11596 , n11594 , n11595 );
nor ( n11597 , n11593 , n11596 );
buf ( n11598 , n11597 );
buf ( n11599 , n11598 );
xor ( n11600 , n4230 , n4433 );
not ( n11601 , n10147 );
nand ( n11602 , n10142 , n4225 );
nand ( n11603 , n11601 , n11602 );
xor ( n11604 , n11600 , n11603 );
buf ( n11605 , n11604 );
buf ( n11606 , n11605 );
buf ( n11607 , n11606 );
nand ( n11608 , n11607 , n378 );
not ( n11609 , n11608 );
not ( n11610 , n8205 );
nor ( n11611 , n11610 , n8184 );
not ( n11612 , n11611 );
buf ( n11613 , n8193 );
not ( n11614 , n11613 );
buf ( n11615 , n11614 );
and ( n11616 , n11615 , n7551 );
not ( n11617 , n11616 );
or ( n11618 , n11612 , n11617 );
not ( n11619 , n8184 );
not ( n11620 , n11619 );
not ( n11621 , n11615 );
or ( n11622 , n11620 , n11621 );
nand ( n11623 , n7551 , n8205 );
nand ( n11624 , n11622 , n11623 );
nand ( n11625 , n11618 , n11624 );
nand ( n11626 , n11609 , n11625 );
buf ( n11627 , n11626 );
not ( n11628 , n11627 );
buf ( n11629 , n11297 );
buf ( n11630 , n11289 );
nand ( n11631 , n11629 , n11630 );
buf ( n11632 , n11631 );
buf ( n11633 , n11632 );
not ( n11634 , n11633 );
buf ( n11635 , n7551 );
not ( n11636 , n11635 );
buf ( n11637 , n8184 );
not ( n11638 , n11637 );
or ( n11639 , n11636 , n11638 );
buf ( n11640 , n8209 );
nand ( n11641 , n11639 , n11640 );
buf ( n11642 , n11641 );
buf ( n11643 , n11642 );
not ( n11644 , n11643 );
or ( n11645 , n11634 , n11644 );
buf ( n11646 , n11642 );
buf ( n11647 , n11632 );
or ( n11648 , n11646 , n11647 );
buf ( n11649 , n11648 );
buf ( n11650 , n11649 );
nand ( n11651 , n11645 , n11650 );
buf ( n11652 , n11651 );
buf ( n11653 , n11652 );
nand ( n11654 , n11628 , n11653 );
buf ( n11655 , n11654 );
buf ( n11656 , n11655 );
nand ( n11657 , n11599 , n11656 );
buf ( n11658 , n11657 );
not ( n11659 , n11658 );
or ( n11660 , n11587 , n11659 );
buf ( n11661 , n11655 );
not ( n11662 , n11661 );
buf ( n11663 , n11598 );
not ( n11664 , n11663 );
buf ( n11665 , n11664 );
buf ( n11666 , n11665 );
nand ( n11667 , n11662 , n11666 );
buf ( n11668 , n11667 );
nand ( n11669 , n11660 , n11668 );
buf ( n11670 , n11669 );
or ( n11671 , n11572 , n11670 );
not ( n11672 , n9745 );
not ( n11673 , n11190 );
or ( n11674 , n11672 , n11673 );
and ( n11675 , n10877 , n9732 );
not ( n11676 , n10877 );
and ( n11677 , n11676 , n380 );
or ( n11678 , n11675 , n11677 );
nand ( n11679 , n11678 , n9743 );
nand ( n11680 , n11674 , n11679 );
nand ( n11681 , n11671 , n11680 );
nand ( n11682 , n11670 , n11572 );
nand ( n11683 , n11681 , n11682 );
not ( n11684 , n11683 );
or ( n11685 , n11561 , n11684 );
nand ( n11686 , n11556 , n11500 );
nand ( n11687 , n11685 , n11686 );
buf ( n11688 , n11687 );
nand ( n11689 , n11498 , n11688 );
buf ( n11690 , n11689 );
nand ( n11691 , n11495 , n11690 );
xor ( n11692 , n11456 , n11691 );
and ( n11693 , n11259 , n11364 );
not ( n11694 , n11259 );
and ( n11695 , n11694 , n11367 );
nor ( n11696 , n11693 , n11695 );
and ( n11697 , n11222 , n11696 );
not ( n11698 , n11222 );
not ( n11699 , n11696 );
and ( n11700 , n11698 , n11699 );
nor ( n11701 , n11697 , n11700 );
and ( n11702 , n11692 , n11701 );
and ( n11703 , n11456 , n11691 );
or ( n11704 , n11702 , n11703 );
not ( n11705 , n11704 );
nand ( n11706 , n11447 , n11705 );
xor ( n11707 , n11456 , n11691 );
xor ( n11708 , n11707 , n11701 );
not ( n11709 , n11708 );
not ( n11710 , n11490 );
not ( n11711 , n11710 );
buf ( n11712 , n11480 );
not ( n11713 , n11712 );
buf ( n11714 , n11713 );
not ( n11715 , n11714 );
or ( n11716 , n11711 , n11715 );
buf ( n11717 , n11480 );
buf ( n11718 , n11490 );
nand ( n11719 , n11717 , n11718 );
buf ( n11720 , n11719 );
nand ( n11721 , n11716 , n11720 );
buf ( n11722 , n11687 );
not ( n11723 , n11722 );
buf ( n11724 , n11723 );
and ( n11725 , n11721 , n11724 );
not ( n11726 , n11721 );
and ( n11727 , n11726 , n11687 );
nor ( n11728 , n11725 , n11727 );
buf ( n11729 , n11728 );
xor ( n11730 , n11103 , n11127 );
xor ( n11731 , n11730 , n11218 );
buf ( n11732 , n11731 );
buf ( n11733 , n11732 );
not ( n11734 , n11733 );
buf ( n11735 , n11734 );
buf ( n11736 , n11735 );
nand ( n11737 , n11729 , n11736 );
buf ( n11738 , n11737 );
not ( n11739 , n11738 );
buf ( n11740 , n385 );
not ( n11741 , n11740 );
buf ( n11742 , n11462 );
not ( n11743 , n11742 );
or ( n11744 , n11741 , n11743 );
not ( n11745 , n384 );
not ( n11746 , n10468 );
or ( n11747 , n11745 , n11746 );
not ( n11748 , n384 );
nand ( n11749 , n11748 , n10465 );
nand ( n11750 , n11747 , n11749 );
buf ( n11751 , n11750 );
buf ( n11752 , n11409 );
nand ( n11753 , n11751 , n11752 );
buf ( n11754 , n11753 );
buf ( n11755 , n11754 );
nand ( n11756 , n11744 , n11755 );
buf ( n11757 , n11756 );
buf ( n11758 , n9836 );
not ( n11759 , n11758 );
buf ( n11760 , n11205 );
not ( n11761 , n11760 );
or ( n11762 , n11759 , n11761 );
not ( n11763 , n9738 );
not ( n11764 , n10508 );
not ( n11765 , n10531 );
or ( n11766 , n11764 , n11765 );
nand ( n11767 , n11766 , n10536 );
not ( n11768 , n11767 );
or ( n11769 , n11763 , n11768 );
or ( n11770 , n9738 , n10537 );
nand ( n11771 , n11769 , n11770 );
buf ( n11772 , n11771 );
buf ( n11773 , n9853 );
nand ( n11774 , n11772 , n11773 );
buf ( n11775 , n11774 );
buf ( n11776 , n11775 );
nand ( n11777 , n11762 , n11776 );
buf ( n11778 , n11777 );
not ( n11779 , n11778 );
buf ( n11780 , n11522 );
buf ( n11781 , n11533 );
xor ( n11782 , n11780 , n11781 );
buf ( n11783 , n11549 );
xor ( n11784 , n11782 , n11783 );
buf ( n11785 , n11784 );
not ( n11786 , n11785 );
not ( n11787 , n11786 );
or ( n11788 , n11779 , n11787 );
not ( n11789 , n11785 );
not ( n11790 , n11775 );
and ( n11791 , n9836 , n11205 );
nor ( n11792 , n11790 , n11791 );
not ( n11793 , n11792 );
or ( n11794 , n11789 , n11793 );
not ( n11795 , n2980 );
not ( n11796 , n3033 );
or ( n11797 , n11795 , n11796 );
nand ( n11798 , n11797 , n2841 );
buf ( n11799 , n2489 );
not ( n11800 , n11799 );
buf ( n11801 , n2495 );
nand ( n11802 , n11800 , n11801 );
buf ( n11803 , n11802 );
buf ( n11804 , n11803 );
not ( n11805 , n11804 );
buf ( n11806 , n11805 );
and ( n11807 , n11798 , n11806 );
not ( n11808 , n11798 );
and ( n11809 , n11808 , n11803 );
nor ( n11810 , n11807 , n11809 );
not ( n11811 , n11810 );
buf ( n11812 , n9743 );
not ( n11813 , n11812 );
not ( n11814 , n9732 );
not ( n11815 , n11072 );
or ( n11816 , n11814 , n11815 );
nand ( n11817 , n380 , n11137 );
nand ( n11818 , n11816 , n11817 );
buf ( n11819 , n11818 );
not ( n11820 , n11819 );
or ( n11821 , n11813 , n11820 );
buf ( n11822 , n11678 );
buf ( n11823 , n9745 );
nand ( n11824 , n11822 , n11823 );
buf ( n11825 , n11824 );
buf ( n11826 , n11825 );
nand ( n11827 , n11821 , n11826 );
buf ( n11828 , n11827 );
not ( n11829 , n11828 );
or ( n11830 , n11811 , n11829 );
buf ( n11831 , n11828 );
buf ( n11832 , n11798 );
buf ( n11833 , n11806 );
and ( n11834 , n11832 , n11833 );
not ( n11835 , n11832 );
buf ( n11836 , n11803 );
and ( n11837 , n11835 , n11836 );
nor ( n11838 , n11834 , n11837 );
buf ( n11839 , n11838 );
buf ( n11840 , n11839 );
or ( n11841 , n11831 , n11840 );
buf ( n11842 , n378 );
not ( n11843 , n10154 );
and ( n11844 , n11843 , n5730 );
not ( n11845 , n11843 );
not ( n11846 , n5730 );
and ( n11847 , n11845 , n11846 );
nor ( n11848 , n11844 , n11847 );
buf ( n11849 , n11848 );
and ( n11850 , n11842 , n11849 );
buf ( n11851 , n11850 );
buf ( n11852 , n11851 );
buf ( n11853 , n11626 );
not ( n11854 , n11853 );
buf ( n11855 , n11652 );
not ( n11856 , n11855 );
or ( n11857 , n11854 , n11856 );
buf ( n11858 , n11652 );
buf ( n11859 , n11626 );
or ( n11860 , n11858 , n11859 );
nand ( n11861 , n11857 , n11860 );
buf ( n11862 , n11861 );
buf ( n11863 , n11862 );
xor ( n11864 , n11852 , n11863 );
buf ( n11865 , n9773 );
not ( n11866 , n11865 );
buf ( n11867 , n11579 );
not ( n11868 , n11867 );
or ( n11869 , n11866 , n11868 );
buf ( n11870 , n378 );
not ( n11871 , n11870 );
buf ( n11872 , n11518 );
not ( n11873 , n11872 );
buf ( n11874 , n11873 );
buf ( n11875 , n11874 );
not ( n11876 , n11875 );
or ( n11877 , n11871 , n11876 );
buf ( n11878 , n11518 );
buf ( n11879 , n9776 );
nand ( n11880 , n11878 , n11879 );
buf ( n11881 , n11880 );
buf ( n11882 , n11881 );
nand ( n11883 , n11877 , n11882 );
buf ( n11884 , n11883 );
buf ( n11885 , n11884 );
buf ( n11886 , n9790 );
nand ( n11887 , n11885 , n11886 );
buf ( n11888 , n11887 );
buf ( n11889 , n11888 );
nand ( n11890 , n11869 , n11889 );
buf ( n11891 , n11890 );
buf ( n11892 , n11891 );
and ( n11893 , n11864 , n11892 );
and ( n11894 , n11852 , n11863 );
or ( n11895 , n11893 , n11894 );
buf ( n11896 , n11895 );
buf ( n11897 , n11896 );
nand ( n11898 , n11841 , n11897 );
buf ( n11899 , n11898 );
nand ( n11900 , n11830 , n11899 );
nand ( n11901 , n11794 , n11900 );
nand ( n11902 , n11788 , n11901 );
xor ( n11903 , n11757 , n11902 );
nand ( n11904 , n11191 , n11180 );
xor ( n11905 , n11164 , n11904 );
xnor ( n11906 , n11905 , n11210 );
and ( n11907 , n11903 , n11906 );
and ( n11908 , n11757 , n11902 );
or ( n11909 , n11907 , n11908 );
not ( n11910 , n11909 );
or ( n11911 , n11739 , n11910 );
not ( n11912 , n11735 );
buf ( n11913 , n11728 );
not ( n11914 , n11913 );
buf ( n11915 , n11914 );
nand ( n11916 , n11912 , n11915 );
nand ( n11917 , n11911 , n11916 );
buf ( n11918 , n11917 );
not ( n11919 , n11918 );
buf ( n11920 , n11919 );
nand ( n11921 , n11709 , n11920 );
and ( n11922 , n11706 , n11921 );
buf ( n11923 , n10871 );
buf ( n11924 , n11035 );
xor ( n11925 , n11923 , n11924 );
buf ( n11926 , n11026 );
xor ( n11927 , n11925 , n11926 );
buf ( n11928 , n11927 );
buf ( n11929 , n11928 );
xor ( n11930 , n10589 , n10608 );
xor ( n11931 , n11930 , n10632 );
buf ( n11932 , n11931 );
buf ( n11933 , n11932 );
not ( n11934 , n11933 );
buf ( n11935 , n10930 );
not ( n11936 , n11935 );
buf ( n11937 , n11936 );
buf ( n11938 , n11937 );
not ( n11939 , n11938 );
not ( n11940 , n11022 );
and ( n11941 , n11940 , n10943 );
not ( n11942 , n11940 );
not ( n11943 , n10943 );
and ( n11944 , n11942 , n11943 );
nor ( n11945 , n11941 , n11944 );
not ( n11946 , n11945 );
buf ( n11947 , n11946 );
not ( n11948 , n11947 );
or ( n11949 , n11939 , n11948 );
buf ( n11950 , n10930 );
buf ( n11951 , n11945 );
nand ( n11952 , n11950 , n11951 );
buf ( n11953 , n11952 );
buf ( n11954 , n11953 );
nand ( n11955 , n11949 , n11954 );
buf ( n11956 , n11955 );
buf ( n11957 , n11956 );
not ( n11958 , n11957 );
or ( n11959 , n11934 , n11958 );
buf ( n11960 , n11932 );
buf ( n11961 , n11937 );
not ( n11962 , n11961 );
buf ( n11963 , n11946 );
not ( n11964 , n11963 );
or ( n11965 , n11962 , n11964 );
buf ( n11966 , n11953 );
nand ( n11967 , n11965 , n11966 );
buf ( n11968 , n11967 );
buf ( n11969 , n11968 );
or ( n11970 , n11960 , n11969 );
buf ( n11971 , n11383 );
not ( n11972 , n11971 );
buf ( n11973 , n11391 );
nand ( n11974 , n11972 , n11973 );
buf ( n11975 , n11974 );
buf ( n11976 , n11975 );
not ( n11977 , n11976 );
buf ( n11978 , n11438 );
not ( n11979 , n11978 );
or ( n11980 , n11977 , n11979 );
buf ( n11981 , n11391 );
not ( n11982 , n11981 );
buf ( n11983 , n11383 );
nand ( n11984 , n11982 , n11983 );
buf ( n11985 , n11984 );
buf ( n11986 , n11985 );
nand ( n11987 , n11980 , n11986 );
buf ( n11988 , n11987 );
buf ( n11989 , n11988 );
nand ( n11990 , n11970 , n11989 );
buf ( n11991 , n11990 );
buf ( n11992 , n11991 );
nand ( n11993 , n11959 , n11992 );
buf ( n11994 , n11993 );
buf ( n11995 , n11994 );
not ( n11996 , n11995 );
buf ( n11997 , n11996 );
buf ( n11998 , n11997 );
nand ( n11999 , n11929 , n11998 );
buf ( n12000 , n11999 );
buf ( n12001 , n12000 );
xor ( n12002 , n11932 , n11956 );
xnor ( n12003 , n12002 , n11988 );
xor ( n12004 , n11064 , n11378 );
and ( n12005 , n12004 , n11443 );
and ( n12006 , n11064 , n11378 );
or ( n12007 , n12005 , n12006 );
buf ( n12008 , n12007 );
not ( n12009 , n12008 );
buf ( n12010 , n12009 );
nand ( n12011 , n12003 , n12010 );
buf ( n12012 , n12011 );
and ( n12013 , n12001 , n12012 );
buf ( n12014 , n12013 );
nand ( n12015 , n11922 , n12014 );
buf ( n12016 , n12015 );
not ( n12017 , n12016 );
buf ( n12018 , n12017 );
not ( n12019 , n11665 );
not ( n12020 , n11655 );
not ( n12021 , n12020 );
and ( n12022 , n12019 , n12021 );
and ( n12023 , n11665 , n12020 );
nor ( n12024 , n12022 , n12023 );
and ( n12025 , n12024 , n11586 );
not ( n12026 , n12024 );
not ( n12027 , n11586 );
and ( n12028 , n12026 , n12027 );
nor ( n12029 , n12025 , n12028 );
buf ( n12030 , n12029 );
buf ( n12031 , n9853 );
not ( n12032 , n12031 );
buf ( n12033 , n382 );
not ( n12034 , n12033 );
buf ( n12035 , n10977 );
not ( n12036 , n12035 );
or ( n12037 , n12034 , n12036 );
buf ( n12038 , n10980 );
buf ( n12039 , n9738 );
nand ( n12040 , n12038 , n12039 );
buf ( n12041 , n12040 );
buf ( n12042 , n12041 );
nand ( n12043 , n12037 , n12042 );
buf ( n12044 , n12043 );
buf ( n12045 , n12044 );
not ( n12046 , n12045 );
or ( n12047 , n12032 , n12046 );
buf ( n12048 , n11771 );
buf ( n12049 , n9836 );
nand ( n12050 , n12048 , n12049 );
buf ( n12051 , n12050 );
buf ( n12052 , n12051 );
nand ( n12053 , n12047 , n12052 );
buf ( n12054 , n12053 );
buf ( n12055 , n12054 );
xor ( n12056 , n12030 , n12055 );
buf ( n12057 , n385 );
not ( n12058 , n12057 );
and ( n12059 , n384 , n10914 );
not ( n12060 , n384 );
and ( n12061 , n12060 , n10485 );
or ( n12062 , n12059 , n12061 );
buf ( n12063 , n12062 );
not ( n12064 , n12063 );
or ( n12065 , n12058 , n12064 );
xor ( n12066 , n384 , n10341 );
buf ( n12067 , n12066 );
buf ( n12068 , n11409 );
nand ( n12069 , n12067 , n12068 );
buf ( n12070 , n12069 );
buf ( n12071 , n12070 );
nand ( n12072 , n12065 , n12071 );
buf ( n12073 , n12072 );
buf ( n12074 , n12073 );
xnor ( n12075 , n12056 , n12074 );
buf ( n12076 , n12075 );
buf ( n12077 , n12076 );
not ( n12078 , n12077 );
buf ( n12079 , n385 );
not ( n12080 , n12079 );
buf ( n12081 , n12066 );
not ( n12082 , n12081 );
or ( n12083 , n12080 , n12082 );
and ( n12084 , n11767 , n384 );
not ( n12085 , n11767 );
not ( n12086 , n384 );
and ( n12087 , n12085 , n12086 );
nor ( n12088 , n12084 , n12087 );
nand ( n12089 , n11409 , n12088 );
buf ( n12090 , n12089 );
nand ( n12091 , n12083 , n12090 );
buf ( n12092 , n12091 );
buf ( n12093 , n12092 );
not ( n12094 , n2837 );
nand ( n12095 , n12094 , n2484 );
not ( n12096 , n12095 );
not ( n12097 , n3007 );
nand ( n12098 , n2954 , n2976 , n12097 );
not ( n12099 , n12098 );
or ( n12100 , n12096 , n12099 );
nor ( n12101 , n3007 , n12095 );
nand ( n12102 , n2954 , n2976 , n12101 );
nand ( n12103 , n12100 , n12102 );
buf ( n12104 , n8181 );
buf ( n12105 , n12104 );
buf ( n12106 , n12105 );
not ( n12107 , n12106 );
buf ( n12108 , n11615 );
buf ( n12109 , n7661 );
nand ( n12110 , n12108 , n12109 );
buf ( n12111 , n12110 );
not ( n12112 , n12111 );
not ( n12113 , n12112 );
or ( n12114 , n12107 , n12113 );
not ( n12115 , n12111 );
or ( n12116 , n12106 , n12115 );
nand ( n12117 , n12114 , n12116 );
not ( n12118 , n394 );
nor ( n12119 , n12117 , n12118 );
buf ( n12120 , n12119 );
not ( n12121 , n11608 );
not ( n12122 , n11625 );
or ( n12123 , n12121 , n12122 );
or ( n12124 , n11608 , n11625 );
nand ( n12125 , n12123 , n12124 );
buf ( n12126 , n12125 );
xor ( n12127 , n12120 , n12126 );
buf ( n12128 , n9773 );
not ( n12129 , n12128 );
buf ( n12130 , n11884 );
not ( n12131 , n12130 );
or ( n12132 , n12129 , n12131 );
xor ( n12133 , n11842 , n11849 );
buf ( n12134 , n12133 );
buf ( n12135 , n12134 );
buf ( n12136 , n9790 );
nand ( n12137 , n12135 , n12136 );
buf ( n12138 , n12137 );
buf ( n12139 , n12138 );
nand ( n12140 , n12132 , n12139 );
buf ( n12141 , n12140 );
buf ( n12142 , n12141 );
and ( n12143 , n12127 , n12142 );
and ( n12144 , n12120 , n12126 );
or ( n12145 , n12143 , n12144 );
buf ( n12146 , n12145 );
not ( n12147 , n12146 );
xor ( n12148 , n12103 , n12147 );
not ( n12149 , n9745 );
not ( n12150 , n11818 );
or ( n12151 , n12149 , n12150 );
not ( n12152 , n11267 );
not ( n12153 , n11271 );
or ( n12154 , n12152 , n12153 );
nand ( n12155 , n12154 , n11277 );
and ( n12156 , n12155 , n380 );
not ( n12157 , n12155 );
not ( n12158 , n380 );
and ( n12159 , n12157 , n12158 );
nor ( n12160 , n12156 , n12159 );
nand ( n12161 , n9743 , n12160 );
nand ( n12162 , n12151 , n12161 );
xnor ( n12163 , n12148 , n12162 );
buf ( n12164 , n12163 );
xor ( n12165 , n12093 , n12164 );
xor ( n12166 , n12120 , n12126 );
xor ( n12167 , n12166 , n12142 );
buf ( n12168 , n12167 );
buf ( n12169 , n12168 );
buf ( n12170 , n9773 );
not ( n12171 , n12170 );
buf ( n12172 , n12134 );
not ( n12173 , n12172 );
or ( n12174 , n12171 , n12173 );
buf ( n12175 , n378 );
not ( n12176 , n12175 );
buf ( n12177 , n11607 );
not ( n12178 , n12177 );
buf ( n12179 , n12178 );
buf ( n12180 , n12179 );
not ( n12181 , n12180 );
or ( n12182 , n12176 , n12181 );
buf ( n12183 , n11604 );
buf ( n12184 , n12183 );
buf ( n12185 , n12184 );
buf ( n12186 , n12185 );
buf ( n12187 , n9776 );
nand ( n12188 , n12186 , n12187 );
buf ( n12189 , n12188 );
buf ( n12190 , n12189 );
nand ( n12191 , n12182 , n12190 );
buf ( n12192 , n12191 );
buf ( n12193 , n12192 );
buf ( n12194 , n9790 );
nand ( n12195 , n12193 , n12194 );
buf ( n12196 , n12195 );
buf ( n12197 , n12196 );
nand ( n12198 , n12174 , n12197 );
buf ( n12199 , n12198 );
buf ( n12200 , n12199 );
buf ( n12201 , n7850 );
not ( n12202 , n12201 );
buf ( n12203 , n7810 );
nand ( n12204 , n12202 , n12203 );
buf ( n12205 , n12204 );
and ( n12206 , n12205 , n7851 );
buf ( n12207 , n8128 );
xor ( n12208 , n12206 , n12207 );
and ( n12209 , n396 , n12208 );
buf ( n12210 , n395 );
and ( n12211 , n8178 , n8172 );
buf ( n12212 , n8139 );
xor ( n12213 , n12211 , n12212 );
buf ( n12214 , n12213 );
xor ( n12215 , n12210 , n12214 );
buf ( n12216 , n11604 );
not ( n12217 , n12216 );
buf ( n12218 , n9774 );
nor ( n12219 , n12217 , n12218 );
buf ( n12220 , n12219 );
buf ( n12221 , n12220 );
xor ( n12222 , n12215 , n12221 );
buf ( n12223 , n12222 );
xor ( n12224 , n12209 , n12223 );
xor ( n12225 , n396 , n12208 );
not ( n12226 , n12225 );
buf ( n12227 , n398 );
not ( n12228 , n8112 );
not ( n12229 , n8106 );
or ( n12230 , n12228 , n12229 );
nand ( n12231 , n12230 , n8045 );
nand ( n12232 , n8102 , n399 );
and ( n12233 , n12231 , n12232 );
not ( n12234 , n12231 );
not ( n12235 , n8102 );
nand ( n12236 , n12235 , n399 );
and ( n12237 , n12234 , n12236 );
nor ( n12238 , n12233 , n12237 );
buf ( n12239 , n12238 );
xor ( n12240 , n12227 , n12239 );
buf ( n12241 , n8018 );
not ( n12242 , n12241 );
buf ( n12243 , n8120 );
nand ( n12244 , n12242 , n12243 );
buf ( n12245 , n12244 );
xor ( n12246 , n8114 , n12245 );
buf ( n12247 , n12246 );
and ( n12248 , n12240 , n12247 );
and ( n12249 , n12227 , n12239 );
or ( n12250 , n12248 , n12249 );
buf ( n12251 , n12250 );
and ( n12252 , n397 , n12251 );
not ( n12253 , n12252 );
nand ( n12254 , n12226 , n12253 );
not ( n12255 , n12254 );
buf ( n12256 , n9738 );
buf ( n12257 , n9731 );
nand ( n12258 , n12256 , n12257 );
buf ( n12259 , n12258 );
not ( n12260 , n12259 );
not ( n12261 , n11607 );
or ( n12262 , n12260 , n12261 );
buf ( n12263 , n381 );
buf ( n12264 , n382 );
and ( n12265 , n12263 , n12264 );
buf ( n12266 , n9732 );
nor ( n12267 , n12265 , n12266 );
buf ( n12268 , n12267 );
nand ( n12269 , n12262 , n12268 );
not ( n12270 , n12269 );
not ( n12271 , n12270 );
or ( n12272 , n12255 , n12271 );
nand ( n12273 , n12225 , n12252 );
nand ( n12274 , n12272 , n12273 );
and ( n12275 , n12224 , n12274 );
and ( n12276 , n12209 , n12223 );
or ( n12277 , n12275 , n12276 );
buf ( n12278 , n12277 );
xor ( n12279 , n12200 , n12278 );
buf ( n12280 , n9732 );
buf ( n12281 , n9780 );
nand ( n12282 , n12280 , n12281 );
buf ( n12283 , n12282 );
buf ( n12284 , n12283 );
not ( n12285 , n12284 );
buf ( n12286 , n11607 );
not ( n12287 , n12286 );
or ( n12288 , n12285 , n12287 );
buf ( n12289 , n379 );
buf ( n12290 , n380 );
and ( n12291 , n12289 , n12290 );
buf ( n12292 , n9776 );
nor ( n12293 , n12291 , n12292 );
buf ( n12294 , n12293 );
buf ( n12295 , n12294 );
nand ( n12296 , n12288 , n12295 );
buf ( n12297 , n12296 );
not ( n12298 , n12118 );
not ( n12299 , n12106 );
not ( n12300 , n12112 );
or ( n12301 , n12299 , n12300 );
or ( n12302 , n12106 , n12115 );
nand ( n12303 , n12301 , n12302 );
not ( n12304 , n12303 );
or ( n12305 , n12298 , n12304 );
or ( n12306 , n12117 , n12118 );
nand ( n12307 , n12305 , n12306 );
not ( n12308 , n12307 );
xor ( n12309 , n12297 , n12308 );
xor ( n12310 , n12210 , n12214 );
and ( n12311 , n12310 , n12221 );
and ( n12312 , n12210 , n12214 );
or ( n12313 , n12311 , n12312 );
buf ( n12314 , n12313 );
xnor ( n12315 , n12309 , n12314 );
buf ( n12316 , n12315 );
and ( n12317 , n12279 , n12316 );
and ( n12318 , n12200 , n12278 );
or ( n12319 , n12317 , n12318 );
buf ( n12320 , n12319 );
buf ( n12321 , n12320 );
xor ( n12322 , n12169 , n12321 );
not ( n12323 , n9836 );
buf ( n12324 , n382 );
not ( n12325 , n12324 );
buf ( n12326 , n10880 );
not ( n12327 , n12326 );
or ( n12328 , n12325 , n12327 );
buf ( n12329 , n10883 );
buf ( n12330 , n9738 );
nand ( n12331 , n12329 , n12330 );
buf ( n12332 , n12331 );
buf ( n12333 , n12332 );
nand ( n12334 , n12328 , n12333 );
buf ( n12335 , n12334 );
not ( n12336 , n12335 );
or ( n12337 , n12323 , n12336 );
not ( n12338 , n382 );
not ( n12339 , n11137 );
or ( n12340 , n12338 , n12339 );
buf ( n12341 , n11072 );
buf ( n12342 , n9738 );
nand ( n12343 , n12341 , n12342 );
buf ( n12344 , n12343 );
nand ( n12345 , n12340 , n12344 );
nand ( n12346 , n12345 , n9853 );
nand ( n12347 , n12337 , n12346 );
buf ( n12348 , n12347 );
and ( n12349 , n12322 , n12348 );
and ( n12350 , n12169 , n12321 );
or ( n12351 , n12349 , n12350 );
buf ( n12352 , n12351 );
buf ( n12353 , n12352 );
and ( n12354 , n12165 , n12353 );
and ( n12355 , n12093 , n12164 );
or ( n12356 , n12354 , n12355 );
buf ( n12357 , n12356 );
buf ( n12358 , n12357 );
not ( n12359 , n12358 );
or ( n12360 , n12078 , n12359 );
buf ( n12361 , n12357 );
buf ( n12362 , n12076 );
or ( n12363 , n12361 , n12362 );
nand ( n12364 , n12360 , n12363 );
buf ( n12365 , n12364 );
buf ( n12366 , n12365 );
not ( n12367 , n12103 );
not ( n12368 , n12367 );
not ( n12369 , n12147 );
or ( n12370 , n12368 , n12369 );
nand ( n12371 , n12370 , n12162 );
nand ( n12372 , n12146 , n12103 );
nand ( n12373 , n12371 , n12372 );
buf ( n12374 , n12373 );
xor ( n12375 , n11810 , n11896 );
xnor ( n12376 , n12375 , n11828 );
buf ( n12377 , n12376 );
xor ( n12378 , n12374 , n12377 );
xor ( n12379 , n11852 , n11863 );
xor ( n12380 , n12379 , n11892 );
buf ( n12381 , n12380 );
buf ( n12382 , n12381 );
buf ( n12383 , n9836 );
not ( n12384 , n12383 );
buf ( n12385 , n12044 );
not ( n12386 , n12385 );
or ( n12387 , n12384 , n12386 );
buf ( n12388 , n12335 );
buf ( n12389 , n9853 );
nand ( n12390 , n12388 , n12389 );
buf ( n12391 , n12390 );
buf ( n12392 , n12391 );
nand ( n12393 , n12387 , n12392 );
buf ( n12394 , n12393 );
buf ( n12395 , n12394 );
xor ( n12396 , n12382 , n12395 );
not ( n12397 , n9745 );
not ( n12398 , n12160 );
or ( n12399 , n12397 , n12398 );
buf ( n12400 , n380 );
not ( n12401 , n12400 );
not ( n12402 , n11342 );
buf ( n12403 , n12402 );
not ( n12404 , n12403 );
or ( n12405 , n12401 , n12404 );
buf ( n12406 , n11342 );
buf ( n12407 , n9732 );
nand ( n12408 , n12406 , n12407 );
buf ( n12409 , n12408 );
buf ( n12410 , n12409 );
nand ( n12411 , n12405 , n12410 );
buf ( n12412 , n12411 );
buf ( n12413 , n12412 );
buf ( n12414 , n9743 );
nand ( n12415 , n12413 , n12414 );
buf ( n12416 , n12415 );
nand ( n12417 , n12399 , n12416 );
not ( n12418 , n12417 );
not ( n12419 , n2479 );
nor ( n12420 , n12419 , n2477 );
not ( n12421 , n12420 );
not ( n12422 , n2905 );
nor ( n12423 , n12422 , n2917 );
not ( n12424 , n12423 );
nand ( n12425 , n2884 , n2948 );
not ( n12426 , n12425 );
or ( n12427 , n12424 , n12426 );
not ( n12428 , n2890 );
nor ( n12429 , n2917 , n12428 );
nand ( n12430 , n2969 , n2471 );
nor ( n12431 , n12429 , n12430 );
nand ( n12432 , n12427 , n12431 );
not ( n12433 , n2471 );
nand ( n12434 , n2465 , n2443 );
not ( n12435 , n12434 );
or ( n12436 , n12433 , n12435 );
nand ( n12437 , n12436 , n2476 );
nor ( n12438 , C0 , n12437 );
nand ( n12439 , n12432 , n12438 );
not ( n12440 , n12439 );
or ( n12441 , n12421 , n12440 );
not ( n12442 , n12420 );
nand ( n12443 , n12438 , n12432 , n12442 );
nand ( n12444 , n12441 , n12443 );
nand ( n12445 , n12418 , n12444 );
not ( n12446 , n12445 );
not ( n12447 , n12308 );
not ( n12448 , n12297 );
not ( n12449 , n12448 );
or ( n12450 , n12447 , n12449 );
not ( n12451 , n12297 );
not ( n12452 , n12307 );
or ( n12453 , n12451 , n12452 );
nand ( n12454 , n12453 , n12314 );
nand ( n12455 , n12450 , n12454 );
not ( n12456 , n12455 );
or ( n12457 , n12446 , n12456 );
not ( n12458 , n12444 );
nand ( n12459 , n12458 , n12417 );
nand ( n12460 , n12457 , n12459 );
buf ( n12461 , n12460 );
and ( n12462 , n12396 , n12461 );
and ( n12463 , n12382 , n12395 );
or ( n12464 , n12462 , n12463 );
buf ( n12465 , n12464 );
buf ( n12466 , n12465 );
xor ( n12467 , n12378 , n12466 );
buf ( n12468 , n12467 );
buf ( n12469 , n12468 );
and ( n12470 , n12366 , n12469 );
not ( n12471 , n12366 );
buf ( n12472 , n12468 );
not ( n12473 , n12472 );
buf ( n12474 , n12473 );
buf ( n12475 , n12474 );
and ( n12476 , n12471 , n12475 );
nor ( n12477 , n12470 , n12476 );
buf ( n12478 , n12477 );
buf ( n12479 , n12478 );
xor ( n12480 , n12382 , n12395 );
xor ( n12481 , n12480 , n12461 );
buf ( n12482 , n12481 );
buf ( n12483 , n12482 );
not ( n12484 , n12483 );
buf ( n12485 , n12484 );
buf ( n12486 , n12485 );
not ( n12487 , n12486 );
not ( n12488 , n385 );
not ( n12489 , n12088 );
or ( n12490 , n12488 , n12489 );
not ( n12491 , n384 );
not ( n12492 , n10977 );
or ( n12493 , n12491 , n12492 );
buf ( n12494 , n384 );
not ( n12495 , n12494 );
buf ( n12496 , n12495 );
nand ( n12497 , n11186 , n12496 );
nand ( n12498 , n12493 , n12497 );
nand ( n12499 , n12498 , n11409 );
nand ( n12500 , n12490 , n12499 );
not ( n12501 , n12500 );
buf ( n12502 , n9745 );
not ( n12503 , n12502 );
buf ( n12504 , n12412 );
not ( n12505 , n12504 );
or ( n12506 , n12503 , n12505 );
buf ( n12507 , n380 );
buf ( n12508 , n11518 );
and ( n12509 , n12507 , n12508 );
not ( n12510 , n12507 );
buf ( n12511 , n11874 );
and ( n12512 , n12510 , n12511 );
nor ( n12513 , n12509 , n12512 );
buf ( n12514 , n12513 );
buf ( n12515 , n12514 );
buf ( n12516 , n9743 );
nand ( n12517 , n12515 , n12516 );
buf ( n12518 , n12517 );
buf ( n12519 , n12518 );
nand ( n12520 , n12506 , n12519 );
buf ( n12521 , n12520 );
buf ( n12522 , n12521 );
nand ( n12523 , n2925 , n2969 , n2936 );
not ( n12524 , n12434 );
nand ( n12525 , n2972 , n12523 , n12524 );
nand ( n12526 , n2471 , n2476 );
xnor ( n12527 , n12525 , n12526 );
buf ( n12528 , n12527 );
xor ( n12529 , n12522 , n12528 );
buf ( n12530 , n9836 );
not ( n12531 , n12530 );
buf ( n12532 , n12345 );
not ( n12533 , n12532 );
or ( n12534 , n12531 , n12533 );
not ( n12535 , n382 );
not ( n12536 , n12155 );
not ( n12537 , n12536 );
or ( n12538 , n12535 , n12537 );
buf ( n12539 , n9738 );
buf ( n12540 , n12155 );
nand ( n12541 , n12539 , n12540 );
buf ( n12542 , n12541 );
nand ( n12543 , n12538 , n12542 );
buf ( n12544 , n12543 );
buf ( n12545 , n9853 );
nand ( n12546 , n12544 , n12545 );
buf ( n12547 , n12546 );
buf ( n12548 , n12547 );
nand ( n12549 , n12534 , n12548 );
buf ( n12550 , n12549 );
buf ( n12551 , n12550 );
and ( n12552 , n12529 , n12551 );
and ( n12553 , n12522 , n12528 );
or ( n12554 , n12552 , n12553 );
buf ( n12555 , n12554 );
not ( n12556 , n12555 );
or ( n12557 , n12501 , n12556 );
buf ( n12558 , n12555 );
buf ( n12559 , n12500 );
or ( n12560 , n12558 , n12559 );
xor ( n12561 , n12455 , n12444 );
xnor ( n12562 , n12561 , n12417 );
buf ( n12563 , n12562 );
nand ( n12564 , n12560 , n12563 );
buf ( n12565 , n12564 );
nand ( n12566 , n12557 , n12565 );
not ( n12567 , n12566 );
buf ( n12568 , n12567 );
not ( n12569 , n12568 );
or ( n12570 , n12487 , n12569 );
xor ( n12571 , n12093 , n12164 );
xor ( n12572 , n12571 , n12353 );
buf ( n12573 , n12572 );
buf ( n12574 , n12573 );
nand ( n12575 , n12570 , n12574 );
buf ( n12576 , n12575 );
buf ( n12577 , n12576 );
buf ( n12578 , n12485 );
buf ( n12579 , n12567 );
or ( n12580 , n12578 , n12579 );
buf ( n12581 , n12580 );
buf ( n12582 , n12581 );
and ( n12583 , n12577 , n12582 );
buf ( n12584 , n12583 );
buf ( n12585 , n12584 );
nand ( n12586 , n12479 , n12585 );
buf ( n12587 , n12586 );
not ( n12588 , n12587 );
buf ( n12589 , n11607 );
buf ( n12590 , n9745 );
and ( n12591 , n12589 , n12590 );
buf ( n12592 , n12591 );
buf ( n12593 , n8127 );
buf ( n12594 , n7923 );
not ( n12595 , n12594 );
buf ( n12596 , n7940 );
nand ( n12597 , n12595 , n12596 );
buf ( n12598 , n12597 );
buf ( n12599 , n12598 );
nand ( n12600 , n12593 , n12599 );
buf ( n12601 , n12600 );
buf ( n12602 , n12601 );
buf ( n12603 , n8123 );
xnor ( n12604 , n12602 , n12603 );
buf ( n12605 , n12604 );
xor ( n12606 , n397 , n12251 );
and ( n12607 , n12605 , n12606 );
not ( n12608 , n12605 );
not ( n12609 , n12606 );
and ( n12610 , n12608 , n12609 );
nor ( n12611 , n12607 , n12610 );
xor ( n12612 , n12592 , n12611 );
not ( n12613 , n9836 );
not ( n12614 , n382 );
not ( n12615 , n11874 );
or ( n12616 , n12614 , n12615 );
buf ( n12617 , n11518 );
buf ( n12618 , n9738 );
nand ( n12619 , n12617 , n12618 );
buf ( n12620 , n12619 );
nand ( n12621 , n12616 , n12620 );
not ( n12622 , n12621 );
or ( n12623 , n12613 , n12622 );
buf ( n12624 , n382 );
not ( n12625 , n12624 );
buf ( n12626 , n11848 );
not ( n12627 , n12626 );
buf ( n12628 , n12627 );
buf ( n12629 , n12628 );
not ( n12630 , n12629 );
or ( n12631 , n12625 , n12630 );
buf ( n12632 , n9738 );
buf ( n12633 , n11848 );
nand ( n12634 , n12632 , n12633 );
buf ( n12635 , n12634 );
buf ( n12636 , n12635 );
nand ( n12637 , n12631 , n12636 );
buf ( n12638 , n12637 );
buf ( n12639 , n12638 );
buf ( n12640 , n9853 );
nand ( n12641 , n12639 , n12640 );
buf ( n12642 , n12641 );
nand ( n12643 , n12623 , n12642 );
xor ( n12644 , n12612 , n12643 );
nand ( n12645 , C1 , n3002 );
nand ( n12646 , n2889 , n2916 );
not ( n12647 , n12646 );
and ( n12648 , n12645 , n12647 );
not ( n12649 , n12645 );
and ( n12650 , n12649 , n12646 );
nor ( n12651 , n12648 , n12650 );
and ( n12652 , n12644 , n12651 );
and ( n12653 , n12612 , n12643 );
or ( n12654 , n12652 , n12653 );
not ( n12655 , n12654 );
nand ( n12656 , n2761 , n2456 );
nand ( n12657 , C1 , n2987 );
or ( n12658 , n12656 , n12657 );
nand ( n12659 , n12657 , n12656 );
nand ( n12660 , n12658 , n12659 );
not ( n12661 , n12660 );
buf ( n12662 , n382 );
not ( n12663 , n12662 );
buf ( n12664 , n12402 );
not ( n12665 , n12664 );
or ( n12666 , n12663 , n12665 );
buf ( n12667 , n9738 );
buf ( n12668 , n11342 );
nand ( n12669 , n12667 , n12668 );
buf ( n12670 , n12669 );
buf ( n12671 , n12670 );
nand ( n12672 , n12666 , n12671 );
buf ( n12673 , n12672 );
and ( n12674 , n12673 , n9836 );
and ( n12675 , n12621 , n9853 );
nor ( n12676 , n12674 , n12675 );
nand ( n12677 , n12661 , n12676 );
not ( n12678 , n12677 );
or ( n12679 , n12655 , n12678 );
not ( n12680 , n12676 );
nand ( n12681 , n12680 , n12660 );
nand ( n12682 , n12679 , n12681 );
not ( n12683 , n12682 );
buf ( n12684 , n12683 );
not ( n12685 , n12684 );
not ( n12686 , n9836 );
not ( n12687 , n12543 );
or ( n12688 , n12686 , n12687 );
nand ( n12689 , n12673 , n9853 );
nand ( n12690 , n12688 , n12689 );
buf ( n12691 , n12690 );
not ( n12692 , n12605 );
nand ( n12693 , n12692 , n12609 );
not ( n12694 , n12693 );
not ( n12695 , n12592 );
or ( n12696 , n12694 , n12695 );
nand ( n12697 , n12606 , n12605 );
nand ( n12698 , n12696 , n12697 );
buf ( n12699 , n12698 );
not ( n12700 , n12699 );
buf ( n12701 , n9745 );
not ( n12702 , n12701 );
buf ( n12703 , n380 );
not ( n12704 , n12703 );
buf ( n12705 , n12628 );
not ( n12706 , n12705 );
or ( n12707 , n12704 , n12706 );
buf ( n12708 , n9732 );
buf ( n12709 , n11848 );
nand ( n12710 , n12708 , n12709 );
buf ( n12711 , n12710 );
buf ( n12712 , n12711 );
nand ( n12713 , n12707 , n12712 );
buf ( n12714 , n12713 );
buf ( n12715 , n12714 );
not ( n12716 , n12715 );
or ( n12717 , n12702 , n12716 );
buf ( n12718 , n12185 );
buf ( n12719 , n9732 );
nand ( n12720 , n12718 , n12719 );
buf ( n12721 , n12720 );
buf ( n12722 , n12721 );
not ( n12723 , n12722 );
not ( n12724 , n12185 );
buf ( n12725 , n12724 );
buf ( n12726 , n380 );
nand ( n12727 , n12725 , n12726 );
buf ( n12728 , n12727 );
buf ( n12729 , n12728 );
not ( n12730 , n12729 );
or ( n12731 , n12723 , n12730 );
buf ( n12732 , n9743 );
nand ( n12733 , n12731 , n12732 );
buf ( n12734 , n12733 );
buf ( n12735 , n12734 );
nand ( n12736 , n12717 , n12735 );
buf ( n12737 , n12736 );
buf ( n12738 , n12737 );
not ( n12739 , n12738 );
or ( n12740 , n12700 , n12739 );
or ( n12741 , n12737 , n12698 );
xor ( n12742 , n12225 , n12253 );
xnor ( n12743 , n12742 , n12269 );
not ( n12744 , n12743 );
nand ( n12745 , n12741 , n12744 );
buf ( n12746 , n12745 );
nand ( n12747 , n12740 , n12746 );
buf ( n12748 , n12747 );
buf ( n12749 , n12748 );
xnor ( n12750 , n12691 , n12749 );
buf ( n12751 , n12750 );
buf ( n12752 , n12751 );
not ( n12753 , n12752 );
not ( n12754 , n385 );
and ( n12755 , n384 , n10880 );
not ( n12756 , n384 );
and ( n12757 , n12756 , n10883 );
or ( n12758 , n12755 , n12757 );
not ( n12759 , n12758 );
or ( n12760 , n12754 , n12759 );
not ( n12761 , n384 );
not ( n12762 , n11137 );
or ( n12763 , n12761 , n12762 );
not ( n12764 , n384 );
nand ( n12765 , n12764 , n11072 );
nand ( n12766 , n12763 , n12765 );
nand ( n12767 , n12766 , n11409 );
nand ( n12768 , n12760 , n12767 );
buf ( n12769 , n12768 );
not ( n12770 , n12769 );
and ( n12771 , n12753 , n12770 );
buf ( n12772 , n12768 );
buf ( n12773 , n12751 );
and ( n12774 , n12772 , n12773 );
nor ( n12775 , n12771 , n12774 );
buf ( n12776 , n12775 );
buf ( n12777 , n12776 );
not ( n12778 , n12777 );
or ( n12779 , n12685 , n12778 );
buf ( n12780 , n9745 );
not ( n12781 , n12780 );
buf ( n12782 , n12514 );
not ( n12783 , n12782 );
or ( n12784 , n12781 , n12783 );
buf ( n12785 , n12714 );
buf ( n12786 , n9743 );
nand ( n12787 , n12785 , n12786 );
buf ( n12788 , n12787 );
buf ( n12789 , n12788 );
nand ( n12790 , n12784 , n12789 );
buf ( n12791 , n12790 );
xor ( n12792 , n12209 , n12223 );
xor ( n12793 , n12792 , n12274 );
xor ( n12794 , n12791 , n12793 );
xnor ( n12795 , n12794 , n3046 );
not ( n12796 , n12795 );
buf ( n12797 , n12796 );
nand ( n12798 , n12779 , n12797 );
buf ( n12799 , n12798 );
buf ( n12800 , n12799 );
buf ( n12801 , n12776 );
not ( n12802 , n12801 );
buf ( n12803 , n12682 );
nand ( n12804 , n12802 , n12803 );
buf ( n12805 , n12804 );
buf ( n12806 , n12805 );
nand ( n12807 , n12800 , n12806 );
buf ( n12808 , n12807 );
buf ( n12809 , n12808 );
xor ( n12810 , n12522 , n12528 );
xor ( n12811 , n12810 , n12551 );
buf ( n12812 , n12811 );
buf ( n12813 , n12812 );
buf ( n12814 , n12690 );
buf ( n12815 , n12814 );
buf ( n12816 , n12815 );
buf ( n12817 , n12816 );
not ( n12818 , n12817 );
buf ( n12819 , n12768 );
not ( n12820 , n12819 );
or ( n12821 , n12818 , n12820 );
buf ( n12822 , n12768 );
buf ( n12823 , n12816 );
or ( n12824 , n12822 , n12823 );
buf ( n12825 , n12748 );
nand ( n12826 , n12824 , n12825 );
buf ( n12827 , n12826 );
buf ( n12828 , n12827 );
nand ( n12829 , n12821 , n12828 );
buf ( n12830 , n12829 );
buf ( n12831 , n12830 );
xor ( n12832 , n12813 , n12831 );
xor ( n12833 , n12200 , n12278 );
xor ( n12834 , n12833 , n12316 );
buf ( n12835 , n12834 );
buf ( n12836 , n12835 );
not ( n12837 , n12791 );
not ( n12838 , n12793 );
or ( n12839 , n12837 , n12838 );
or ( n12840 , n12791 , n12793 );
nand ( n12841 , n12840 , n3046 );
nand ( n12842 , n12839 , n12841 );
buf ( n12843 , n12842 );
xor ( n12844 , n12836 , n12843 );
buf ( n12845 , n385 );
not ( n12846 , n12845 );
buf ( n12847 , n12498 );
not ( n12848 , n12847 );
or ( n12849 , n12846 , n12848 );
buf ( n12850 , n12758 );
buf ( n12851 , n11409 );
nand ( n12852 , n12850 , n12851 );
buf ( n12853 , n12852 );
buf ( n12854 , n12853 );
nand ( n12855 , n12849 , n12854 );
buf ( n12856 , n12855 );
buf ( n12857 , n12856 );
xor ( n12858 , n12844 , n12857 );
buf ( n12859 , n12858 );
buf ( n12860 , n12859 );
xor ( n12861 , n12832 , n12860 );
buf ( n12862 , n12861 );
buf ( n12863 , n12862 );
xor ( n12864 , n12809 , n12863 );
not ( n12865 , n12744 );
buf ( n12866 , n12698 );
not ( n12867 , n12866 );
buf ( n12868 , n12867 );
not ( n12869 , n12868 );
or ( n12870 , n12865 , n12869 );
nand ( n12871 , n12743 , n12698 );
nand ( n12872 , n12870 , n12871 );
not ( n12873 , n12737 );
and ( n12874 , n12872 , n12873 );
not ( n12875 , n12872 );
and ( n12876 , n12875 , n12737 );
nor ( n12877 , n12874 , n12876 );
not ( n12878 , n12877 );
buf ( n12879 , n12878 );
not ( n12880 , n12879 );
not ( n12881 , n385 );
not ( n12882 , n12766 );
or ( n12883 , n12881 , n12882 );
and ( n12884 , n384 , n12536 );
not ( n12885 , n384 );
and ( n12886 , n12885 , n12155 );
or ( n12887 , n12884 , n12886 );
nand ( n12888 , n12887 , n11409 );
nand ( n12889 , n12883 , n12888 );
buf ( n12890 , n12889 );
not ( n12891 , n12890 );
or ( n12892 , n12880 , n12891 );
buf ( n12893 , n12889 );
not ( n12894 , n12893 );
buf ( n12895 , n12877 );
nand ( n12896 , n12894 , n12895 );
buf ( n12897 , n12896 );
not ( n12898 , n385 );
not ( n12899 , n12887 );
or ( n12900 , n12898 , n12899 );
buf ( n12901 , n384 );
buf ( n12902 , n11342 );
and ( n12903 , n12901 , n12902 );
not ( n12904 , n12901 );
buf ( n12905 , n12402 );
and ( n12906 , n12904 , n12905 );
nor ( n12907 , n12903 , n12906 );
buf ( n12908 , n12907 );
buf ( n12909 , n12908 );
buf ( n12910 , n11409 );
nand ( n12911 , n12909 , n12910 );
buf ( n12912 , n12911 );
nand ( n12913 , n12900 , n12912 );
not ( n12914 , n12913 );
xor ( n12915 , n12227 , n12239 );
xor ( n12916 , n12915 , n12247 );
buf ( n12917 , n12916 );
buf ( n12918 , n12917 );
buf ( n12919 , n384 );
not ( n12920 , n12919 );
buf ( n12921 , n9845 );
nand ( n12922 , n12920 , n12921 );
buf ( n12923 , n12922 );
buf ( n12924 , n12923 );
not ( n12925 , n12924 );
buf ( n12926 , n12185 );
not ( n12927 , n12926 );
or ( n12928 , n12925 , n12927 );
buf ( n12929 , n383 );
buf ( n12930 , n384 );
and ( n12931 , n12929 , n12930 );
buf ( n12932 , n9738 );
nor ( n12933 , n12931 , n12932 );
buf ( n12934 , n12933 );
buf ( n12935 , n12934 );
nand ( n12936 , n12928 , n12935 );
buf ( n12937 , n12936 );
buf ( n12938 , n12937 );
not ( n12939 , n12938 );
buf ( n12940 , n12939 );
buf ( n12941 , n12940 );
xor ( n12942 , n12918 , n12941 );
buf ( n12943 , n9836 );
not ( n12944 , n12943 );
buf ( n12945 , n12638 );
not ( n12946 , n12945 );
or ( n12947 , n12944 , n12946 );
not ( n12948 , n12185 );
nand ( n12949 , n12948 , n382 );
not ( n12950 , n12949 );
buf ( n12951 , n12185 );
buf ( n12952 , n9738 );
nand ( n12953 , n12951 , n12952 );
buf ( n12954 , n12953 );
not ( n12955 , n12954 );
or ( n12956 , n12950 , n12955 );
nand ( n12957 , n12956 , n9853 );
buf ( n12958 , n12957 );
nand ( n12959 , n12947 , n12958 );
buf ( n12960 , n12959 );
buf ( n12961 , n12960 );
and ( n12962 , n12942 , n12961 );
and ( n12963 , n12918 , n12941 );
or ( n12964 , n12962 , n12963 );
buf ( n12965 , n12964 );
not ( n12966 , n12965 );
or ( n12967 , n12914 , n12966 );
buf ( n12968 , n12965 );
buf ( n12969 , n12913 );
or ( n12970 , n12968 , n12969 );
xor ( n12971 , n12612 , n12643 );
xor ( n12972 , n12971 , n12651 );
buf ( n12973 , n12972 );
nand ( n12974 , n12970 , n12973 );
buf ( n12975 , n12974 );
nand ( n12976 , n12967 , n12975 );
nand ( n12977 , n12897 , n12976 );
buf ( n12978 , n12977 );
nand ( n12979 , n12892 , n12978 );
buf ( n12980 , n12979 );
buf ( n12981 , n12980 );
not ( n12982 , n12981 );
xnor ( n12983 , n12795 , n12682 );
buf ( n12984 , n12983 );
not ( n12985 , n12984 );
buf ( n12986 , n12776 );
not ( n12987 , n12986 );
and ( n12988 , n12985 , n12987 );
buf ( n12989 , n12983 );
buf ( n12990 , n12776 );
and ( n12991 , n12989 , n12990 );
nor ( n12992 , n12988 , n12991 );
buf ( n12993 , n12992 );
buf ( n12994 , n12993 );
nand ( n12995 , n12982 , n12994 );
buf ( n12996 , n12995 );
buf ( n12997 , n12996 );
not ( n12998 , n12997 );
not ( n12999 , n12889 );
not ( n13000 , n12878 );
or ( n13001 , n12999 , n13000 );
not ( n13002 , n12889 );
nand ( n13003 , n13002 , n12877 );
nand ( n13004 , n13001 , n13003 );
not ( n13005 , n13004 );
not ( n13006 , n12976 );
or ( n13007 , n13005 , n13006 );
not ( n13008 , n12660 );
not ( n13009 , n12676 );
not ( n13010 , n13009 );
or ( n13011 , n13008 , n13010 );
or ( n13012 , n12660 , n13009 );
nand ( n13013 , n13011 , n13012 );
buf ( n13014 , n13013 );
buf ( n13015 , n12654 );
xor ( n13016 , n13014 , n13015 );
buf ( n13017 , n13016 );
nand ( n13018 , n13007 , n13017 );
not ( n13019 , n13018 );
not ( n13020 , n12976 );
not ( n13021 , n13004 );
nand ( n13022 , n13020 , n13021 );
nand ( n13023 , n13019 , n13022 );
not ( n13024 , n13023 );
buf ( n13025 , n11409 );
not ( n13026 , n13025 );
buf ( n13027 , n384 );
not ( n13028 , n13027 );
buf ( n13029 , n12628 );
not ( n13030 , n13029 );
or ( n13031 , n13028 , n13030 );
buf ( n13032 , n384 );
not ( n13033 , n13032 );
buf ( n13034 , n11848 );
nand ( n13035 , n13033 , n13034 );
buf ( n13036 , n13035 );
buf ( n13037 , n13036 );
nand ( n13038 , n13031 , n13037 );
buf ( n13039 , n13038 );
buf ( n13040 , n13039 );
not ( n13041 , n13040 );
or ( n13042 , n13026 , n13041 );
buf ( n13043 , n384 );
buf ( n13044 , n11874 );
and ( n13045 , n13043 , n13044 );
not ( n13046 , n13043 );
buf ( n13047 , n11518 );
and ( n13048 , n13046 , n13047 );
nor ( n13049 , n13045 , n13048 );
buf ( n13050 , n13049 );
buf ( n13051 , n13050 );
buf ( n13052 , n11408 );
or ( n13053 , n13051 , n13052 );
nand ( n13054 , n13042 , n13053 );
buf ( n13055 , n13054 );
buf ( n13056 , n13055 );
not ( n13057 , n8102 );
not ( n13058 , n12231 );
or ( n13059 , n13057 , n13058 );
or ( n13060 , n12231 , n8102 );
nand ( n13061 , n13059 , n13060 );
buf ( n13062 , n13061 );
buf ( n13063 , n399 );
xor ( n13064 , n13062 , n13063 );
buf ( n13065 , n13064 );
buf ( n13066 , n13065 );
buf ( n13067 , n12185 );
buf ( n13068 , n9836 );
and ( n13069 , n13067 , n13068 );
buf ( n13070 , n13069 );
buf ( n13071 , n13070 );
xor ( n13072 , n13066 , n13071 );
buf ( n13073 , n400 );
buf ( n13074 , n8081 );
not ( n13075 , n13074 );
buf ( n13076 , n8099 );
nand ( n13077 , n13075 , n13076 );
buf ( n13078 , n13077 );
buf ( n13079 , n13078 );
buf ( n13080 , n8093 );
xor ( n13081 , n13079 , n13080 );
buf ( n13082 , n13081 );
buf ( n13083 , n13082 );
xor ( n13084 , n13073 , n13083 );
buf ( n13085 , n11604 );
buf ( n13086 , n385 );
nand ( n13087 , n13085 , n13086 );
buf ( n13088 , n13087 );
buf ( n13089 , n13088 );
buf ( n13090 , n384 );
and ( n13091 , n13089 , n13090 );
buf ( n13092 , n13091 );
buf ( n13093 , n13092 );
and ( n13094 , n13084 , n13093 );
and ( n13095 , n13073 , n13083 );
or ( n13096 , n13094 , n13095 );
buf ( n13097 , n13096 );
buf ( n13098 , n13097 );
xor ( n13099 , n13072 , n13098 );
buf ( n13100 , n13099 );
buf ( n13101 , n13100 );
xor ( n13102 , n13056 , n13101 );
buf ( n13103 , n401 );
not ( n13104 , n13103 );
or ( n13105 , n7962 , n8087 );
nand ( n13106 , n13105 , n8090 );
buf ( n13107 , n13106 );
not ( n13108 , n13107 );
or ( n13109 , n13104 , n13108 );
buf ( n13110 , n13088 );
buf ( n13111 , n13106 );
buf ( n13112 , n401 );
nor ( n13113 , n13111 , n13112 );
buf ( n13114 , n13113 );
buf ( n13115 , n13114 );
or ( n13116 , n13110 , n13115 );
nand ( n13117 , n13109 , n13116 );
buf ( n13118 , n13117 );
buf ( n13119 , n13118 );
xor ( n13120 , n13073 , n13083 );
xor ( n13121 , n13120 , n13093 );
buf ( n13122 , n13121 );
buf ( n13123 , n13122 );
xor ( n13124 , n13119 , n13123 );
not ( n13125 , n385 );
not ( n13126 , n13039 );
or ( n13127 , n13125 , n13126 );
nand ( n13128 , n12724 , n11409 );
nand ( n13129 , n13127 , n13128 );
buf ( n13130 , n13129 );
and ( n13131 , n13124 , n13130 );
and ( n13132 , n13119 , n13123 );
or ( n13133 , n13131 , n13132 );
buf ( n13134 , n13133 );
buf ( n13135 , n13134 );
and ( n13136 , n13102 , n13135 );
and ( n13137 , n13056 , n13101 );
or ( n13138 , n13136 , n13137 );
buf ( n13139 , n13138 );
xor ( n13140 , n12918 , n12941 );
xor ( n13141 , n13140 , n12961 );
buf ( n13142 , n13141 );
nor ( n13143 , n13139 , n13142 );
not ( n13144 , n12422 );
and ( n13145 , n12425 , n13144 );
nand ( n13146 , n13145 , n2953 );
and ( n13147 , n13146 , n3038 );
not ( n13148 , n13146 );
and ( n13149 , n13148 , n3035 );
nor ( n13150 , n13147 , n13149 );
xor ( n13151 , n13066 , n13071 );
and ( n13152 , n13151 , n13098 );
and ( n13153 , n13066 , n13071 );
or ( n13154 , n13152 , n13153 );
buf ( n13155 , n13154 );
xor ( n13156 , n13150 , n13155 );
buf ( n13157 , n385 );
not ( n13158 , n13157 );
buf ( n13159 , n12908 );
not ( n13160 , n13159 );
or ( n13161 , n13158 , n13160 );
buf ( n13162 , n13050 );
not ( n13163 , n13162 );
buf ( n13164 , n11409 );
nand ( n13165 , n13163 , n13164 );
buf ( n13166 , n13165 );
buf ( n13167 , n13166 );
nand ( n13168 , n13161 , n13167 );
buf ( n13169 , n13168 );
xor ( n13170 , n13156 , n13169 );
not ( n13171 , n13170 );
or ( n13172 , n13143 , n13171 );
nand ( n13173 , n13139 , n13142 );
nand ( n13174 , n13172 , n13173 );
not ( n13175 , n13174 );
xor ( n13176 , n13150 , n13155 );
and ( n13177 , n13176 , n13169 );
and ( n13178 , n13150 , n13155 );
or ( n13179 , n13177 , n13178 );
not ( n13180 , n13179 );
buf ( n13181 , n12965 );
buf ( n13182 , n12913 );
xor ( n13183 , n13181 , n13182 );
buf ( n13184 , n12972 );
xnor ( n13185 , n13183 , n13184 );
buf ( n13186 , n13185 );
nand ( n13187 , n13180 , n13186 );
not ( n13188 , n13187 );
or ( n13189 , n13175 , n13188 );
not ( n13190 , n13186 );
nand ( n13191 , n13190 , n13179 );
nand ( n13192 , n13189 , n13191 );
not ( n13193 , n13192 );
or ( n13194 , n13024 , n13193 );
buf ( n13195 , n13017 );
not ( n13196 , n13195 );
buf ( n13197 , n13196 );
not ( n13198 , n13020 );
nand ( n13199 , n13198 , n13021 );
not ( n13200 , n12976 );
nand ( n13201 , n13200 , n13004 );
nand ( n13202 , n13197 , n13199 , n13201 );
nand ( n13203 , n13194 , n13202 );
buf ( n13204 , n13203 );
not ( n13205 , n13204 );
or ( n13206 , n12998 , n13205 );
buf ( n13207 , n12993 );
not ( n13208 , n13207 );
buf ( n13209 , n12980 );
nand ( n13210 , n13208 , n13209 );
buf ( n13211 , n13210 );
buf ( n13212 , n13211 );
nand ( n13213 , n13206 , n13212 );
buf ( n13214 , n13213 );
buf ( n13215 , n13214 );
and ( n13216 , n12864 , n13215 );
and ( n13217 , n12809 , n12863 );
or ( n13218 , n13216 , n13217 );
buf ( n13219 , n13218 );
buf ( n13220 , n13219 );
not ( n13221 , n13220 );
buf ( n13222 , n12482 );
buf ( n13223 , n12566 );
and ( n13224 , n13222 , n13223 );
not ( n13225 , n13222 );
buf ( n13226 , n12567 );
and ( n13227 , n13225 , n13226 );
nor ( n13228 , n13224 , n13227 );
buf ( n13229 , n13228 );
buf ( n13230 , n12573 );
not ( n13231 , n13230 );
buf ( n13232 , n13231 );
and ( n13233 , n13229 , n13232 );
not ( n13234 , n13229 );
and ( n13235 , n13234 , n12573 );
nor ( n13236 , n13233 , n13235 );
xor ( n13237 , n12169 , n12321 );
xor ( n13238 , n13237 , n12348 );
buf ( n13239 , n13238 );
xor ( n13240 , n12836 , n12843 );
and ( n13241 , n13240 , n12857 );
and ( n13242 , n12836 , n12843 );
or ( n13243 , n13241 , n13242 );
buf ( n13244 , n13243 );
xor ( n13245 , n13239 , n13244 );
buf ( n13246 , n12562 );
not ( n13247 , n13246 );
buf ( n13248 , n12500 );
not ( n13249 , n13248 );
buf ( n13250 , n13249 );
buf ( n13251 , n13250 );
not ( n13252 , n13251 );
or ( n13253 , n13247 , n13252 );
not ( n13254 , n12562 );
buf ( n13255 , n13254 );
buf ( n13256 , n12500 );
nand ( n13257 , n13255 , n13256 );
buf ( n13258 , n13257 );
buf ( n13259 , n13258 );
nand ( n13260 , n13253 , n13259 );
buf ( n13261 , n13260 );
buf ( n13262 , n13261 );
buf ( n13263 , n12555 );
and ( n13264 , n13262 , n13263 );
not ( n13265 , n13262 );
buf ( n13266 , n12555 );
not ( n13267 , n13266 );
buf ( n13268 , n13267 );
buf ( n13269 , n13268 );
and ( n13270 , n13265 , n13269 );
nor ( n13271 , n13264 , n13270 );
buf ( n13272 , n13271 );
and ( n13273 , n13245 , n13272 );
and ( n13274 , n13239 , n13244 );
or ( n13275 , n13273 , n13274 );
not ( n13276 , n13275 );
nand ( n13277 , n13236 , n13276 );
buf ( n13278 , n13277 );
xor ( n13279 , n12813 , n12831 );
and ( n13280 , n13279 , n12860 );
and ( n13281 , n12813 , n12831 );
or ( n13282 , n13280 , n13281 );
buf ( n13283 , n13282 );
not ( n13284 , n13283 );
xor ( n13285 , n13239 , n13244 );
xor ( n13286 , n13285 , n13272 );
not ( n13287 , n13286 );
nand ( n13288 , n13284 , n13287 );
buf ( n13289 , n13288 );
and ( n13290 , n13278 , n13289 );
buf ( n13291 , n13290 );
buf ( n13292 , n13291 );
not ( n13293 , n13292 );
or ( n13294 , n13221 , n13293 );
buf ( n13295 , n13286 );
buf ( n13296 , n13283 );
nand ( n13297 , n13295 , n13296 );
buf ( n13298 , n13297 );
buf ( n13299 , n13298 );
not ( n13300 , n13299 );
buf ( n13301 , n13277 );
nand ( n13302 , n13300 , n13301 );
buf ( n13303 , n13302 );
not ( n13304 , n13236 );
buf ( n13305 , n13275 );
nand ( n13306 , n13304 , n13305 );
nand ( n13307 , n13303 , n13306 );
buf ( n13308 , n13307 );
not ( n13309 , n13308 );
buf ( n13310 , n13309 );
buf ( n13311 , n13310 );
nand ( n13312 , n13294 , n13311 );
buf ( n13313 , n13312 );
not ( n13314 , n13313 );
or ( n13315 , n12588 , n13314 );
buf ( n13316 , n12478 );
buf ( n13317 , n12584 );
or ( n13318 , n13316 , n13317 );
buf ( n13319 , n13318 );
nand ( n13320 , n13315 , n13319 );
not ( n13321 , n13320 );
buf ( n13322 , n11732 );
buf ( n13323 , n11909 );
xor ( n13324 , n13322 , n13323 );
buf ( n13325 , n11915 );
xnor ( n13326 , n13324 , n13325 );
buf ( n13327 , n13326 );
xor ( n13328 , n11757 , n11902 );
xor ( n13329 , n13328 , n11906 );
buf ( n13330 , n13329 );
not ( n13331 , n13330 );
buf ( n13332 , n13331 );
not ( n13333 , n13332 );
buf ( n13334 , n11683 );
and ( n13335 , n11500 , n11556 );
not ( n13336 , n11500 );
and ( n13337 , n13336 , n11559 );
nor ( n13338 , n13335 , n13337 );
buf ( n13339 , n13338 );
xnor ( n13340 , n13334 , n13339 );
buf ( n13341 , n13340 );
not ( n13342 , n13341 );
and ( n13343 , n13333 , n13342 );
buf ( n13344 , n13332 );
buf ( n13345 , n13341 );
nand ( n13346 , n13344 , n13345 );
buf ( n13347 , n13346 );
and ( n13348 , n11571 , n11669 );
not ( n13349 , n11571 );
not ( n13350 , n11669 );
and ( n13351 , n13349 , n13350 );
nor ( n13352 , n13348 , n13351 );
and ( n13353 , n13352 , n11680 );
not ( n13354 , n13352 );
not ( n13355 , n11680 );
and ( n13356 , n13354 , n13355 );
nor ( n13357 , n13353 , n13356 );
buf ( n13358 , n13357 );
not ( n13359 , n13358 );
not ( n13360 , n11409 );
not ( n13361 , n12062 );
or ( n13362 , n13360 , n13361 );
nand ( n13363 , n11750 , n385 );
nand ( n13364 , n13362 , n13363 );
not ( n13365 , n13364 );
buf ( n13366 , n13365 );
not ( n13367 , n13366 );
or ( n13368 , n13359 , n13367 );
not ( n13369 , n12054 );
not ( n13370 , n12073 );
or ( n13371 , n13369 , n13370 );
buf ( n13372 , n12073 );
buf ( n13373 , n12054 );
or ( n13374 , n13372 , n13373 );
buf ( n13375 , n12029 );
nand ( n13376 , n13374 , n13375 );
buf ( n13377 , n13376 );
nand ( n13378 , n13371 , n13377 );
buf ( n13379 , n13378 );
nand ( n13380 , n13368 , n13379 );
buf ( n13381 , n13380 );
buf ( n13382 , n13381 );
buf ( n13383 , n13357 );
not ( n13384 , n13383 );
buf ( n13385 , n13364 );
nand ( n13386 , n13384 , n13385 );
buf ( n13387 , n13386 );
buf ( n13388 , n13387 );
nand ( n13389 , n13382 , n13388 );
buf ( n13390 , n13389 );
and ( n13391 , n13347 , n13390 );
nor ( n13392 , n13343 , n13391 );
nand ( n13393 , n13327 , n13392 );
buf ( n13394 , n13393 );
not ( n13395 , n11900 );
not ( n13396 , n11786 );
not ( n13397 , n11778 );
not ( n13398 , n13397 );
or ( n13399 , n13396 , n13398 );
nand ( n13400 , n11785 , n11778 );
nand ( n13401 , n13399 , n13400 );
xnor ( n13402 , n13395 , n13401 );
not ( n13403 , n13402 );
buf ( n13404 , n12373 );
not ( n13405 , n13404 );
buf ( n13406 , n13405 );
not ( n13407 , n13406 );
not ( n13408 , n12376 );
or ( n13409 , n13407 , n13408 );
nand ( n13410 , n13409 , n12465 );
not ( n13411 , n12376 );
nand ( n13412 , n13411 , n12373 );
nand ( n13413 , n13410 , n13412 );
not ( n13414 , n13413 );
or ( n13415 , n13403 , n13414 );
not ( n13416 , n13365 );
not ( n13417 , n13357 );
not ( n13418 , n13417 );
or ( n13419 , n13416 , n13418 );
nand ( n13420 , n13357 , n13364 );
nand ( n13421 , n13419 , n13420 );
and ( n13422 , n13421 , n13378 );
not ( n13423 , n13421 );
not ( n13424 , n13378 );
and ( n13425 , n13423 , n13424 );
nor ( n13426 , n13422 , n13425 );
not ( n13427 , n13426 );
not ( n13428 , n13395 );
not ( n13429 , n13401 );
not ( n13430 , n13429 );
or ( n13431 , n13428 , n13430 );
nand ( n13432 , n13401 , n11900 );
nand ( n13433 , n13431 , n13432 );
not ( n13434 , n13433 );
nor ( n13435 , n13434 , n13413 );
or ( n13436 , n13427 , n13435 );
nand ( n13437 , n13415 , n13436 );
not ( n13438 , n13437 );
not ( n13439 , n13341 );
not ( n13440 , n13390 );
not ( n13441 , n13440 );
or ( n13442 , n13439 , n13441 );
not ( n13443 , n13341 );
nand ( n13444 , n13443 , n13390 );
nand ( n13445 , n13442 , n13444 );
and ( n13446 , n13445 , n13329 );
not ( n13447 , n13445 );
not ( n13448 , n13329 );
and ( n13449 , n13447 , n13448 );
nor ( n13450 , n13446 , n13449 );
nand ( n13451 , n13438 , n13450 );
buf ( n13452 , n13451 );
not ( n13453 , n13452 );
buf ( n13454 , n13453 );
buf ( n13455 , n13454 );
and ( n13456 , n13413 , n13402 );
not ( n13457 , n13413 );
and ( n13458 , n13457 , n13433 );
nor ( n13459 , n13456 , n13458 );
and ( n13460 , n13459 , n13427 );
not ( n13461 , n13459 );
and ( n13462 , n13461 , n13426 );
nor ( n13463 , n13460 , n13462 );
not ( n13464 , n13463 );
not ( n13465 , n12076 );
not ( n13466 , n13465 );
not ( n13467 , n12474 );
or ( n13468 , n13466 , n13467 );
not ( n13469 , n12076 );
not ( n13470 , n12468 );
or ( n13471 , n13469 , n13470 );
nand ( n13472 , n13471 , n12357 );
nand ( n13473 , n13468 , n13472 );
nor ( n13474 , n13464 , n13473 );
buf ( n13475 , n13474 );
nor ( n13476 , n13455 , n13475 );
buf ( n13477 , n13476 );
buf ( n13478 , n13477 );
and ( n13479 , n13394 , n13478 );
buf ( n13480 , n13479 );
not ( n13481 , n13480 );
or ( n13482 , n13321 , n13481 );
not ( n13483 , n13393 );
not ( n13484 , n13465 );
not ( n13485 , n12474 );
or ( n13486 , n13484 , n13485 );
nand ( n13487 , n13486 , n13472 );
not ( n13488 , n13487 );
nor ( n13489 , n13488 , n13463 );
not ( n13490 , n13489 );
not ( n13491 , n13451 );
or ( n13492 , n13490 , n13491 );
buf ( n13493 , n13450 );
not ( n13494 , n13493 );
buf ( n13495 , n13437 );
buf ( n13496 , n13495 );
nand ( n13497 , n13494 , n13496 );
buf ( n13498 , n13497 );
nand ( n13499 , n13492 , n13498 );
not ( n13500 , n13499 );
or ( n13501 , n13483 , n13500 );
buf ( n13502 , n13327 );
not ( n13503 , n13502 );
buf ( n13504 , n13503 );
buf ( n13505 , n13392 );
not ( n13506 , n13505 );
buf ( n13507 , n13506 );
nand ( n13508 , n13504 , n13507 );
nand ( n13509 , n13501 , n13508 );
not ( n13510 , n13509 );
nand ( n13511 , n13482 , n13510 );
and ( n13512 , n12018 , n13511 );
not ( n13513 , n13512 );
or ( n13514 , n11062 , n13513 );
not ( n13515 , n10834 );
not ( n13516 , n10812 );
and ( n13517 , n13515 , n13516 );
and ( n13518 , n10834 , n10812 );
nor ( n13519 , n13518 , n10838 );
nor ( n13520 , n13517 , n13519 );
nor ( n13521 , n10805 , n13520 );
not ( n13522 , n13521 );
buf ( n13523 , n10793 );
buf ( n13524 , n10725 );
nand ( n13525 , n13523 , n13524 );
buf ( n13526 , n13525 );
buf ( n13527 , n13526 );
nand ( n13528 , n10849 , n10862 );
buf ( n13529 , n13528 );
and ( n13530 , n13527 , n13529 );
buf ( n13531 , n13530 );
not ( n13532 , n13531 );
buf ( n13533 , n10725 );
not ( n13534 , n13533 );
buf ( n13535 , n10796 );
nand ( n13536 , n13534 , n13535 );
buf ( n13537 , n13536 );
buf ( n13538 , n11056 );
buf ( n13539 , n11050 );
nor ( n13540 , n13538 , n13539 );
buf ( n13541 , n13540 );
nand ( n13542 , n13537 , n13541 );
not ( n13543 , n13542 );
or ( n13544 , n13532 , n13543 );
and ( n13545 , n10842 , n10864 );
nand ( n13546 , n13544 , n13545 );
nand ( n13547 , n13522 , n13546 );
nor ( n13548 , n12010 , n12003 );
not ( n13549 , n13548 );
not ( n13550 , n12000 );
or ( n13551 , n13549 , n13550 );
buf ( n13552 , n11928 );
not ( n13553 , n13552 );
buf ( n13554 , n13553 );
buf ( n13555 , n13554 );
buf ( n13556 , n11994 );
nand ( n13557 , n13555 , n13556 );
buf ( n13558 , n13557 );
nand ( n13559 , n13551 , n13558 );
not ( n13560 , n13559 );
nand ( n13561 , n11708 , n11917 );
nand ( n13562 , n11444 , n11704 );
nand ( n13563 , n13561 , n13562 );
nand ( n13564 , n13563 , n11706 , n12011 , n12000 );
nand ( n13565 , n13560 , n13564 );
nor ( n13566 , n10843 , n11060 );
nand ( n13567 , n13565 , n13566 );
not ( n13568 , n13567 );
nor ( n13569 , n13547 , n13568 );
nand ( n13570 , n13514 , n13569 );
not ( n13571 , n13570 );
or ( n13572 , n10308 , n13571 );
nor ( n13573 , n10090 , n10015 );
nand ( n13574 , n10294 , n10303 );
or ( n13575 , n13573 , n13574 );
nand ( n13576 , n13575 , C1 );
buf ( n13577 , n13576 );
not ( n13578 , n13577 );
buf ( n13579 , n13578 );
nand ( n13580 , n13572 , n13579 );
buf ( n13581 , n13580 );
and ( n13582 , n13581 , n10013 );
not ( n13583 , n13581 );
and ( n13584 , n13583 , n10012 );
nor ( n13585 , n13582 , n13584 );
buf ( n13586 , n13585 );
buf ( n13587 , n13521 );
not ( n13588 , n13587 );
buf ( n13589 , n10842 );
nand ( n13590 , n13588 , n13589 );
buf ( n13591 , n13590 );
buf ( n13592 , n13591 );
buf ( n13593 , n13591 );
not ( n13594 , n13593 );
buf ( n13595 , n13594 );
buf ( n13596 , n13595 );
buf ( n13597 , n10864 );
not ( n13598 , n13597 );
buf ( n13599 , n11057 );
not ( n13600 , n13599 );
buf ( n13601 , n10796 );
not ( n13602 , n13601 );
buf ( n13603 , n10725 );
nor ( n13604 , n13602 , n13603 );
buf ( n13605 , n13604 );
buf ( n13606 , n13605 );
nor ( n13607 , n13600 , n13606 );
buf ( n13608 , n13607 );
buf ( n13609 , n13608 );
not ( n13610 , n13609 );
not ( n13611 , n13511 );
not ( n13612 , n12018 );
or ( n13613 , n13611 , n13612 );
not ( n13614 , n13565 );
nand ( n13615 , n13613 , n13614 );
buf ( n13616 , n13615 );
not ( n13617 , n13616 );
or ( n13618 , n13610 , n13617 );
buf ( n13619 , n13526 );
buf ( n13620 , n13619 );
buf ( n13621 , n13620 );
and ( n13622 , n13542 , n13621 );
buf ( n13623 , n13622 );
nand ( n13624 , n13618 , n13623 );
buf ( n13625 , n13624 );
not ( n13626 , n13625 );
or ( n13627 , n13598 , n13626 );
buf ( n13628 , n13528 );
nand ( n13629 , n13627 , n13628 );
buf ( n13630 , n13629 );
and ( n13631 , n13630 , n13596 );
not ( n13632 , n13630 );
and ( n13633 , n13632 , n13592 );
nor ( n13634 , n13631 , n13633 );
buf ( n13635 , n13634 );
buf ( n13636 , n10864 );
buf ( n13637 , n13628 );
nand ( n13638 , n13636 , n13637 );
buf ( n13639 , n13638 );
buf ( n13640 , n13639 );
buf ( n13641 , n13639 );
not ( n13642 , n13641 );
buf ( n13643 , n13642 );
buf ( n13644 , n13643 );
buf ( n13645 , n13625 );
and ( n13646 , n13645 , n13644 );
not ( n13647 , n13645 );
and ( n13648 , n13647 , n13640 );
nor ( n13649 , n13646 , n13648 );
buf ( n13650 , n13649 );
buf ( n13651 , n9755 );
buf ( n13652 , n9863 );
and ( n13653 , n13651 , n13652 );
buf ( n13654 , n9752 );
buf ( n13655 , n9860 );
and ( n13656 , n13654 , n13655 );
nor ( n13657 , n13653 , n13656 );
buf ( n13658 , n13657 );
buf ( n13659 , n13658 );
buf ( n13660 , n9828 );
and ( n13661 , n13659 , n13660 );
not ( n13662 , n13659 );
buf ( n13663 , n9801 );
and ( n13664 , n13662 , n13663 );
or ( n13665 , n13661 , n13664 );
buf ( n13666 , n13665 );
buf ( n13667 , n13666 );
buf ( n13668 , n9755 );
and ( n13669 , n13667 , n13668 );
not ( n13670 , n13667 );
buf ( n13671 , n9752 );
and ( n13672 , n13670 , n13671 );
nor ( n13673 , n13669 , n13672 );
buf ( n13674 , n13673 );
buf ( n13675 , n13674 );
not ( n13676 , n13675 );
buf ( n13677 , n9755 );
buf ( n13678 , n9860 );
or ( n13679 , n13677 , n13678 );
buf ( n13680 , n9752 );
buf ( n13681 , n9863 );
or ( n13682 , n13680 , n13681 );
buf ( n13683 , n9801 );
nand ( n13684 , n13682 , n13683 );
buf ( n13685 , n13684 );
buf ( n13686 , n13685 );
nand ( n13687 , n13679 , n13686 );
buf ( n13688 , n13687 );
buf ( n13689 , n13688 );
not ( n13690 , n13689 );
and ( n13691 , n13676 , n13690 );
buf ( n13692 , n13674 );
buf ( n13693 , n13688 );
and ( n13694 , n13692 , n13693 );
nor ( n13695 , n13691 , n13694 );
buf ( n13696 , n13695 );
buf ( n13697 , n10267 );
buf ( n13698 , n9860 );
nand ( n13699 , n13697 , n13698 );
buf ( n13700 , n13699 );
buf ( n13701 , n13700 );
not ( n13702 , n13701 );
buf ( n13703 , n13702 );
not ( n13704 , n13703 );
not ( n13705 , n13666 );
and ( n13706 , n13704 , n13705 );
buf ( n13707 , n13666 );
buf ( n13708 , n13703 );
nand ( n13709 , n13707 , n13708 );
buf ( n13710 , n13709 );
buf ( n13711 , n12086 );
not ( n13712 , n13711 );
buf ( n13713 , n9752 );
buf ( n13714 , n9828 );
nand ( n13715 , n13713 , n13714 );
buf ( n13716 , n13715 );
buf ( n13717 , n13716 );
not ( n13718 , n13717 );
or ( n13719 , n13712 , n13718 );
buf ( n13720 , n9809 );
nand ( n13721 , n13719 , n13720 );
buf ( n13722 , n13721 );
and ( n13723 , n13710 , n13722 );
nor ( n13724 , n13706 , n13723 );
buf ( n13725 , n9758 );
not ( n13726 , n13725 );
buf ( n13727 , n9906 );
nand ( n13728 , n13726 , n13727 );
buf ( n13729 , n13728 );
not ( n13730 , n13729 );
not ( n13731 , n10266 );
not ( n13732 , n9863 );
or ( n13733 , n13731 , n13732 );
nand ( n13734 , n13733 , n13700 );
not ( n13735 , n13734 );
or ( n13736 , n13730 , n13735 );
buf ( n13737 , n9761 );
buf ( n13738 , n9988 );
nand ( n13739 , n13737 , n13738 );
buf ( n13740 , n13739 );
nand ( n13741 , n13736 , n13740 );
buf ( n13742 , n13741 );
buf ( n13743 , n13722 );
buf ( n13744 , n13666 );
xor ( n13745 , n13743 , n13744 );
buf ( n13746 , n13700 );
xnor ( n13747 , n13745 , n13746 );
buf ( n13748 , n13747 );
buf ( n13749 , n13748 );
or ( n13750 , n13742 , n13749 );
buf ( n13751 , n13750 );
buf ( n13752 , n13751 );
not ( n13753 , n13752 );
buf ( n13754 , n9835 );
buf ( n13755 , n9755 );
and ( n13756 , n13754 , n13755 );
not ( n13757 , n13754 );
buf ( n13758 , n9752 );
and ( n13759 , n13757 , n13758 );
nor ( n13760 , n13756 , n13759 );
buf ( n13761 , n13760 );
buf ( n13762 , n13761 );
buf ( n13763 , n13729 );
buf ( n13764 , n9880 );
nand ( n13765 , n13763 , n13764 );
buf ( n13766 , n13765 );
buf ( n13767 , n13766 );
buf ( n13768 , n13740 );
nand ( n13769 , n13767 , n13768 );
buf ( n13770 , n13769 );
buf ( n13771 , n13770 );
xor ( n13772 , n13762 , n13771 );
buf ( n13773 , n13734 );
not ( n13774 , n13773 );
buf ( n13775 , n13774 );
buf ( n13776 , n13775 );
not ( n13777 , n13776 );
buf ( n13778 , n9917 );
not ( n13779 , n13778 );
or ( n13780 , n13777 , n13779 );
buf ( n13781 , n9917 );
buf ( n13782 , n13775 );
or ( n13783 , n13781 , n13782 );
nand ( n13784 , n13780 , n13783 );
buf ( n13785 , n13784 );
buf ( n13786 , n13785 );
and ( n13787 , n13772 , n13786 );
and ( n13788 , n13762 , n13771 );
or ( n13789 , n13787 , n13788 );
buf ( n13790 , n13789 );
buf ( n13791 , n13790 );
not ( n13792 , n13791 );
or ( n13793 , n13753 , n13792 );
buf ( n13794 , n13741 );
buf ( n13795 , n13748 );
nand ( n13796 , n13794 , n13795 );
buf ( n13797 , n13796 );
buf ( n13798 , n13797 );
nand ( n13799 , n13793 , n13798 );
buf ( n13800 , n13799 );
buf ( n13801 , n13800 );
not ( n13802 , n13801 );
or ( n13803 , C0 , n13802 );
buf ( n13804 , n13724 );
buf ( n13805 , n13696 );
nor ( n13806 , n13804 , n13805 );
buf ( n13807 , n13806 );
buf ( n13808 , n13807 );
not ( n13809 , n13808 );
buf ( n13810 , n13809 );
buf ( n13811 , n13810 );
nand ( n13812 , n13803 , n13811 );
buf ( n13813 , n13812 );
buf ( n13814 , n6572 );
not ( n13815 , n13814 );
buf ( n13816 , n13815 );
buf ( n13817 , n13816 );
buf ( n13818 , n415 );
buf ( n13819 , n416 );
and ( n13820 , n13818 , n13819 );
buf ( n13821 , n6458 );
not ( n13822 , n13821 );
buf ( n13823 , n13822 );
buf ( n13824 , n13823 );
nor ( n13825 , n13820 , n13824 );
buf ( n13826 , n13825 );
buf ( n13827 , n13826 );
or ( n13828 , n13817 , n13827 );
buf ( n13829 , n6584 );
nand ( n13830 , n13828 , n13829 );
buf ( n13831 , n13830 );
buf ( n13832 , n13831 );
buf ( n13833 , n6577 );
xor ( n13834 , n13832 , n13833 );
buf ( n13835 , n9559 );
buf ( n13836 , n415 );
and ( n13837 , n13835 , n13836 );
not ( n13838 , n13835 );
buf ( n13839 , n6467 );
and ( n13840 , n13838 , n13839 );
nor ( n13841 , n13837 , n13840 );
buf ( n13842 , n13841 );
buf ( n13843 , n13842 );
not ( n13844 , n13843 );
buf ( n13845 , n9452 );
not ( n13846 , n13845 );
or ( n13847 , n13844 , n13846 );
buf ( n13848 , n9452 );
buf ( n13849 , n13842 );
or ( n13850 , n13848 , n13849 );
nand ( n13851 , n13847 , n13850 );
buf ( n13852 , n13851 );
buf ( n13853 , n13852 );
and ( n13854 , n13834 , n13853 );
and ( n13855 , n13832 , n13833 );
or ( n13856 , n13854 , n13855 );
buf ( n13857 , n13856 );
buf ( n13858 , n13857 );
buf ( n13859 , n9493 );
buf ( n13860 , n13842 );
or ( n13861 , n13859 , n13860 );
buf ( n13862 , n6445 );
buf ( n13863 , n6557 );
or ( n13864 , n13862 , n13863 );
nand ( n13865 , n13861 , n13864 );
buf ( n13866 , n13865 );
buf ( n13867 , n13866 );
buf ( n13868 , n6542 );
xor ( n13869 , n13867 , n13868 );
buf ( n13870 , n6581 );
not ( n13871 , n6500 );
buf ( n13872 , n13871 );
buf ( n13873 , n6523 );
or ( n13874 , n13872 , n13873 );
buf ( n13875 , n6519 );
buf ( n13876 , n6496 );
or ( n13877 , n13875 , n13876 );
nand ( n13878 , n13874 , n13877 );
buf ( n13879 , n13878 );
buf ( n13880 , n13879 );
xor ( n13881 , n13870 , n13880 );
buf ( n13882 , n6542 );
buf ( n13883 , n415 );
nor ( n13884 , n13882 , n13883 );
buf ( n13885 , n13884 );
buf ( n13886 , n13885 );
xor ( n13887 , n13881 , n13886 );
buf ( n13888 , n13887 );
buf ( n13889 , n13888 );
xor ( n13890 , n13869 , n13889 );
buf ( n13891 , n13890 );
buf ( n13892 , n13891 );
xor ( n13893 , n13858 , n13892 );
xor ( n13894 , n13832 , n13833 );
xor ( n13895 , n13894 , n13853 );
buf ( n13896 , n13895 );
buf ( n13897 , n13896 );
not ( n13898 , n13897 );
buf ( n13899 , n13826 );
buf ( n13900 , n6581 );
and ( n13901 , n13899 , n13900 );
not ( n13902 , n13899 );
buf ( n13903 , n6445 );
and ( n13904 , n13902 , n13903 );
nor ( n13905 , n13901 , n13904 );
buf ( n13906 , n13905 );
xor ( n13907 , n13906 , n6577 );
buf ( n13908 , n13907 );
buf ( n13909 , n6566 );
xor ( n13910 , n13908 , n13909 );
buf ( n13911 , n6607 );
and ( n13912 , n13910 , n13911 );
and ( n13913 , n13908 , n13909 );
or ( n13914 , n13912 , n13913 );
buf ( n13915 , n13914 );
buf ( n13916 , n13915 );
nand ( n13917 , n13898 , n13916 );
buf ( n13918 , n13917 );
buf ( n13919 , n13918 );
not ( n13920 , n13919 );
xor ( n13921 , n13908 , n13909 );
xor ( n13922 , n13921 , n13911 );
buf ( n13923 , n13922 );
buf ( n13924 , n13923 );
buf ( n13925 , n6592 );
nand ( n13926 , n13924 , n13925 );
buf ( n13927 , n13926 );
not ( n13928 , n13927 );
buf ( n13929 , n9716 );
buf ( n13930 , n13929 );
buf ( n13931 , n13930 );
not ( n13932 , n13931 );
or ( n13933 , n13928 , n13932 );
buf ( n13934 , n13923 );
not ( n13935 , n13934 );
buf ( n13936 , n6589 );
nand ( n13937 , n13935 , n13936 );
buf ( n13938 , n13937 );
nand ( n13939 , n13933 , n13938 );
buf ( n13940 , n13939 );
not ( n13941 , n13940 );
or ( n13942 , n13920 , n13941 );
buf ( n13943 , n13915 );
not ( n13944 , n13943 );
buf ( n13945 , n13896 );
nand ( n13946 , n13944 , n13945 );
buf ( n13947 , n13946 );
buf ( n13948 , n13947 );
nand ( n13949 , n13942 , n13948 );
buf ( n13950 , n13949 );
buf ( n13951 , n13950 );
xor ( n13952 , n13893 , n13951 );
buf ( n13953 , n13952 );
not ( n13954 , n13953 );
buf ( n13955 , C1 );
buf ( n13956 , n13955 );
buf ( n13957 , n13813 );
buf ( n13958 , n13954 );
nand ( n13959 , n13957 , n13958 );
buf ( n13960 , n13959 );
buf ( n13961 , n13960 );
nand ( n13962 , n13956 , n13961 );
buf ( n13963 , n13962 );
buf ( n13964 , n13963 );
buf ( n13965 , n13963 );
not ( n13966 , n13965 );
buf ( n13967 , n13966 );
buf ( n13968 , n13967 );
buf ( n13969 , n13947 );
buf ( n13970 , n13918 );
nand ( n13971 , n13969 , n13970 );
buf ( n13972 , n13971 );
xnor ( n13973 , n13972 , n13939 );
buf ( n13974 , n13973 );
not ( n13975 , n13974 );
xor ( n13976 , n13696 , n13724 );
xnor ( n13977 , n13976 , n13800 );
buf ( n13978 , n13977 );
nand ( n13979 , n13975 , n13978 );
buf ( n13980 , n13979 );
buf ( n13981 , n13980 );
and ( n13982 , n13938 , n13927 );
xor ( n13983 , n13982 , n13931 );
buf ( n13984 , n13983 );
not ( n13985 , n13984 );
buf ( n13986 , n13790 );
buf ( n13987 , n13986 );
buf ( n13988 , n13987 );
buf ( n13989 , n13988 );
buf ( n13990 , n13741 );
buf ( n13991 , n13748 );
xor ( n13992 , n13990 , n13991 );
buf ( n13993 , n13992 );
buf ( n13994 , n13993 );
xnor ( n13995 , n13989 , n13994 );
buf ( n13996 , n13995 );
buf ( n13997 , n13996 );
nand ( n13998 , n13985 , n13997 );
buf ( n13999 , n13998 );
buf ( n14000 , n13999 );
not ( n14001 , n9889 );
not ( n14002 , n9917 );
or ( n14003 , n14001 , n14002 );
nand ( n14004 , n14003 , n9923 );
not ( n14005 , n14004 );
nand ( n14006 , n14005 , n9868 );
not ( n14007 , n14006 );
buf ( n14008 , n13770 );
buf ( n14009 , n14008 );
buf ( n14010 , n14009 );
not ( n14011 , n14010 );
or ( n14012 , n14007 , n14011 );
buf ( n14013 , n14004 );
buf ( n14014 , n9867 );
nand ( n14015 , n14013 , n14014 );
buf ( n14016 , n14015 );
nand ( n14017 , n14012 , n14016 );
xor ( n14018 , n13762 , n13771 );
xor ( n14019 , n14018 , n13786 );
buf ( n14020 , n14019 );
or ( n14021 , n14017 , n14020 );
buf ( n14022 , n14021 );
and ( n14023 , n13981 , n14000 , n14022 );
buf ( n14024 , n14023 );
not ( n14025 , n14024 );
not ( n14026 , n14006 );
not ( n14027 , n9886 );
or ( n14028 , n14026 , n14027 );
nand ( n14029 , n14028 , n14016 );
not ( n14030 , n14029 );
not ( n14031 , n14010 );
not ( n14032 , n9931 );
or ( n14033 , n14031 , n14032 );
buf ( n14034 , n14010 );
not ( n14035 , n14034 );
buf ( n14036 , n9928 );
nand ( n14037 , n14035 , n14036 );
buf ( n14038 , n14037 );
nand ( n14039 , n14033 , n14038 );
not ( n14040 , n14039 );
and ( n14041 , n14030 , n14040 );
not ( n14042 , n9935 );
not ( n14043 , n10003 );
and ( n14044 , n14042 , n14043 );
nor ( n14045 , n14041 , n14044 );
and ( n14046 , n10091 , n14045 , n10305 );
not ( n14047 , n14046 );
nor ( n14048 , n14047 , n10843 );
nor ( n14049 , n12015 , n11060 );
nand ( n14050 , n13511 , n14048 , n14049 );
not ( n14051 , n14045 );
not ( n14052 , n13576 );
or ( n14053 , n14051 , n14052 );
nand ( n14054 , n14053 , C1 );
buf ( n14055 , n14054 );
buf ( n14056 , n13521 );
nor ( n14057 , n14055 , n14056 );
buf ( n14058 , n14057 );
nand ( n14059 , n13546 , n14058 );
or ( n14060 , n13568 , n14059 );
not ( n14061 , n14054 );
not ( n14062 , n14046 );
and ( n14063 , n14061 , n14062 );
nor ( n14064 , n14017 , n14039 );
nor ( n14065 , n14063 , n14064 );
nand ( n14066 , n14060 , n14065 );
nand ( n14067 , n14050 , n14066 );
not ( n14068 , n14067 );
or ( n14069 , n14025 , n14068 );
buf ( n14070 , C0 );
buf ( n14071 , C1 );
nand ( n14072 , n14069 , C1 );
buf ( n14073 , n14072 );
and ( n14074 , n14073 , n13968 );
not ( n14075 , n14073 );
and ( n14076 , n14075 , n13964 );
nor ( n14077 , n14074 , n14076 );
buf ( n14078 , n14077 );
buf ( n14079 , n13605 );
not ( n14080 , n14079 );
buf ( n14081 , n13621 );
nand ( n14082 , n14080 , n14081 );
buf ( n14083 , n14082 );
buf ( n14084 , n14083 );
buf ( n14085 , n14083 );
not ( n14086 , n14085 );
buf ( n14087 , n14086 );
buf ( n14088 , n14087 );
not ( n14089 , n11057 );
not ( n14090 , n13615 );
or ( n14091 , n14089 , n14090 );
not ( n14092 , n13541 );
nand ( n14093 , n14091 , n14092 );
buf ( n14094 , n14093 );
and ( n14095 , n14094 , n14088 );
not ( n14096 , n14094 );
and ( n14097 , n14096 , n14084 );
nor ( n14098 , n14095 , n14097 );
buf ( n14099 , n14098 );
buf ( n14100 , n13548 );
not ( n14101 , n14100 );
buf ( n14102 , n12011 );
nand ( n14103 , n14101 , n14102 );
buf ( n14104 , n14103 );
buf ( n14105 , n14103 );
not ( n14106 , n14105 );
buf ( n14107 , n14106 );
buf ( n14108 , n14107 );
not ( n14109 , n13511 );
not ( n14110 , n11922 );
or ( n14111 , n14109 , n14110 );
buf ( n14112 , n11706 );
buf ( n14113 , n13563 );
nand ( n14114 , n14112 , n14113 );
nand ( n14115 , n14111 , n14114 );
buf ( n14116 , n14115 );
and ( n14117 , n14116 , n14108 );
not ( n14118 , n14116 );
and ( n14119 , n14118 , n14104 );
nor ( n14120 , n14117 , n14119 );
buf ( n14121 , n14120 );
buf ( n14122 , n14092 );
buf ( n14123 , n11057 );
nand ( n14124 , n14122 , n14123 );
buf ( n14125 , n14124 );
buf ( n14126 , n14125 );
buf ( n14127 , n14125 );
not ( n14128 , n14127 );
buf ( n14129 , n14128 );
buf ( n14130 , n14129 );
buf ( n14131 , n13615 );
and ( n14132 , n14131 , n14130 );
not ( n14133 , n14131 );
and ( n14134 , n14133 , n14126 );
nor ( n14135 , n14132 , n14134 );
buf ( n14136 , n14135 );
buf ( n14137 , n13393 );
buf ( n14138 , n13508 );
nand ( n14139 , n14137 , n14138 );
buf ( n14140 , n14139 );
buf ( n14141 , n14140 );
buf ( n14142 , n14140 );
not ( n14143 , n14142 );
buf ( n14144 , n14143 );
buf ( n14145 , n14144 );
buf ( n14146 , n13454 );
not ( n14147 , n14146 );
buf ( n14148 , n14147 );
buf ( n14149 , n14148 );
not ( n14150 , n14149 );
buf ( n14151 , n13474 );
not ( n14152 , n14151 );
buf ( n14153 , n14152 );
not ( n14154 , n14153 );
not ( n14155 , n12587 );
not ( n14156 , n13313 );
or ( n14157 , n14155 , n14156 );
nand ( n14158 , n14157 , n13319 );
not ( n14159 , n14158 );
or ( n14160 , n14154 , n14159 );
buf ( n14161 , n13489 );
not ( n14162 , n14161 );
buf ( n14163 , n14162 );
nand ( n14164 , n14160 , n14163 );
buf ( n14165 , n14164 );
not ( n14166 , n14165 );
or ( n14167 , n14150 , n14166 );
buf ( n14168 , n13498 );
buf ( n14169 , n14168 );
buf ( n14170 , n14169 );
buf ( n14171 , n14170 );
nand ( n14172 , n14167 , n14171 );
buf ( n14173 , n14172 );
buf ( n14174 , n14173 );
and ( n14175 , n14174 , n14145 );
not ( n14176 , n14174 );
and ( n14177 , n14176 , n14141 );
nor ( n14178 , n14175 , n14177 );
buf ( n14179 , n14178 );
nand ( n14180 , n14112 , n13562 );
buf ( n14181 , n14180 );
buf ( n14182 , n14180 );
not ( n14183 , n14182 );
buf ( n14184 , n14183 );
buf ( n14185 , n14184 );
buf ( n14186 , n11921 );
buf ( n14187 , n14186 );
not ( n14188 , n14187 );
buf ( n14189 , n13511 );
not ( n14190 , n14189 );
or ( n14191 , n14188 , n14190 );
buf ( n14192 , n13561 );
nand ( n14193 , n14191 , n14192 );
buf ( n14194 , n14193 );
and ( n14195 , n14194 , n14185 );
not ( n14196 , n14194 );
and ( n14197 , n14196 , n14181 );
nor ( n14198 , n14195 , n14197 );
buf ( n14199 , n14198 );
buf ( n14200 , n13319 );
buf ( n14201 , n12587 );
buf ( n14202 , n14201 );
nand ( n14203 , n14200 , n14202 );
buf ( n14204 , n14203 );
buf ( n14205 , n14204 );
not ( n14206 , n14205 );
buf ( n14207 , n14206 );
buf ( n14208 , n14207 );
buf ( n14209 , n14204 );
buf ( n14210 , n13219 );
not ( n14211 , n14210 );
buf ( n14212 , n13291 );
not ( n14213 , n14212 );
or ( n14214 , n14211 , n14213 );
buf ( n14215 , n13310 );
nand ( n14216 , n14214 , n14215 );
buf ( n14217 , n14216 );
buf ( n14218 , n14217 );
not ( n14219 , n14218 );
buf ( n14220 , n14219 );
buf ( n14221 , n14220 );
and ( n14222 , n14221 , n14209 );
not ( n14223 , n14221 );
and ( n14224 , n14223 , n14208 );
nor ( n14225 , n14222 , n14224 );
buf ( n14226 , n14225 );
nand ( n14227 , n13306 , n13277 );
buf ( n14228 , n14227 );
buf ( n14229 , n13288 );
buf ( n14230 , n14229 );
not ( n14231 , n14230 );
buf ( n14232 , n13219 );
buf ( n14233 , n14232 );
buf ( n14234 , n14233 );
buf ( n14235 , n14234 );
not ( n14236 , n14235 );
or ( n14237 , n14231 , n14236 );
buf ( n14238 , n13298 );
buf ( n14239 , n14238 );
nand ( n14240 , n14237 , n14239 );
buf ( n14241 , n14240 );
buf ( n14242 , n14241 );
buf ( n14243 , n14227 );
buf ( n14244 , n14241 );
not ( n14245 , n14228 );
not ( n14246 , n14242 );
or ( n14247 , n14245 , n14246 );
or ( n14248 , n14243 , n14244 );
nand ( n14249 , n14247 , n14248 );
buf ( n14250 , n14249 );
nand ( n14251 , n14229 , n14238 );
buf ( n14252 , n14251 );
buf ( n14253 , n14234 );
buf ( n14254 , n14234 );
buf ( n14255 , n14251 );
not ( n14256 , n14252 );
not ( n14257 , n14253 );
or ( n14258 , n14256 , n14257 );
or ( n14259 , n14254 , n14255 );
nand ( n14260 , n14258 , n14259 );
buf ( n14261 , n14260 );
or ( n14262 , n5832 , n7195 );
not ( n14263 , n6444 );
or ( n14264 , n14263 , n5840 );
nand ( n14265 , n14262 , n14264 );
xor ( n14266 , n14265 , n6542 );
nand ( n14267 , n6524 , n413 );
xor ( n14268 , n9559 , n14267 );
and ( n14269 , n14268 , n6581 );
and ( n14270 , n9559 , n14267 );
or ( n14271 , n14269 , n14270 );
and ( n14272 , n14266 , n14271 );
and ( n14273 , n14265 , n6542 );
or ( n14274 , n14272 , n14273 );
nand ( n14275 , n5841 , n411 );
xnor ( n14276 , n14274 , n14275 );
not ( n14277 , n14276 );
xor ( n14278 , n9559 , n14267 );
xor ( n14279 , n14278 , n6581 );
xor ( n14280 , n14279 , n9559 );
xor ( n14281 , n13870 , n13880 );
and ( n14282 , n14281 , n13886 );
and ( n14283 , n13870 , n13880 );
or ( n14284 , n14282 , n14283 );
buf ( n14285 , n14284 );
and ( n14286 , n14280 , n14285 );
and ( n14287 , n14279 , n9559 );
or ( n14288 , n14286 , n14287 );
xor ( n14289 , n14265 , n6542 );
xor ( n14290 , n14289 , n14271 );
nor ( n14291 , n14288 , n14290 );
not ( n14292 , n14291 );
xor ( n14293 , n13858 , n13892 );
and ( n14294 , n14293 , n13951 );
and ( n14295 , n13858 , n13892 );
or ( n14296 , n14294 , n14295 );
buf ( n14297 , n14296 );
buf ( n14298 , n14297 );
xor ( n14299 , n13867 , n13868 );
and ( n14300 , n14299 , n13889 );
and ( n14301 , n13867 , n13868 );
or ( n14302 , n14300 , n14301 );
buf ( n14303 , n14302 );
not ( n14304 , n14303 );
xor ( n14305 , n14279 , n9559 );
xor ( n14306 , n14305 , n14285 );
not ( n14307 , n14306 );
nand ( n14308 , n14304 , n14307 );
nand ( n14309 , n14292 , n14298 , n14308 );
not ( n14310 , n14291 );
nand ( n14311 , n14310 , n14303 , n14306 );
nand ( n14312 , n14288 , n14290 );
nand ( n14313 , n14309 , n14311 , n14312 );
not ( n14314 , n14313 );
or ( n14315 , n14277 , n14314 );
or ( n14316 , n14313 , n14276 );
nand ( n14317 , n14315 , n14316 );
not ( n14318 , n14317 );
not ( n14319 , n13800 );
or ( n14320 , C0 , n14319 );
nor ( n14321 , C0 , n13807 );
nand ( n14322 , n14320 , n14321 );
nand ( n14323 , n14318 , n14322 );
buf ( n14324 , n14323 );
not ( n14325 , n14308 );
not ( n14326 , n14298 );
or ( n14327 , n14325 , n14326 );
nand ( n14328 , n14303 , n14306 );
nand ( n14329 , n14327 , n14328 );
not ( n14330 , n14290 );
nand ( n14331 , n14330 , n14288 );
nor ( n14332 , n14329 , n14331 );
not ( n14333 , n14288 );
nand ( n14334 , n14333 , n14290 );
nor ( n14335 , n14329 , n14334 );
nor ( n14336 , n14332 , n14335 );
not ( n14337 , n14312 );
or ( n14338 , n14337 , n14291 );
nand ( n14339 , n14338 , n14329 );
nand ( n14340 , n14336 , n14339 );
not ( n14341 , n14340 );
nand ( n14342 , n14341 , n14322 );
buf ( n14343 , n14342 );
nand ( n14344 , n14324 , n14343 );
buf ( n14345 , n14344 );
nand ( n14346 , n14298 , n14303 , n14306 );
not ( n14347 , n14308 );
nand ( n14348 , n14347 , n14298 );
not ( n14349 , n14298 );
nand ( n14350 , n14349 , n14303 , n14307 );
nand ( n14351 , n14349 , n14304 , n14306 );
nand ( n14352 , n14346 , n14348 , n14350 , n14351 );
buf ( n14353 , n14352 );
not ( n14354 , n14353 );
buf ( n14355 , n14322 );
nand ( n14356 , n14354 , n14355 );
buf ( n14357 , n14356 );
buf ( n14358 , n14357 );
buf ( n14359 , n13960 );
nand ( n14360 , n14358 , n14359 );
buf ( n14361 , n14360 );
buf ( n14362 , n14361 );
not ( n14363 , n14362 );
buf ( n14364 , n14363 );
not ( n14365 , n14322 );
buf ( n14366 , C1 );
buf ( n14367 , C1 );
or ( n14368 , n14274 , n14275 );
not ( n14369 , n14368 );
not ( n14370 , n14313 );
or ( n14371 , n14369 , n14370 );
nand ( n14372 , n14274 , n14275 );
nand ( n14373 , n14371 , n14372 );
not ( n14374 , n6540 );
and ( n14375 , n9559 , n14374 );
nor ( n14376 , n14373 , n14375 );
buf ( n14377 , n14376 );
not ( n14378 , n14377 );
buf ( n14379 , n14373 );
buf ( n14380 , n14375 );
nand ( n14381 , n14379 , n14380 );
buf ( n14382 , n14381 );
buf ( n14383 , n14382 );
nand ( n14384 , n14378 , n14383 );
buf ( n14385 , n14384 );
xnor ( n14386 , n14374 , n14376 );
or ( n14387 , n14386 , n14365 );
buf ( n14388 , n14387 );
buf ( n14389 , n14365 );
buf ( n14390 , n14385 );
or ( n14391 , n14389 , n14390 );
buf ( n14392 , n14391 );
buf ( n14393 , n14392 );
nand ( n14394 , n14388 , n14393 );
buf ( n14395 , n14394 );
buf ( n14396 , C1 );
buf ( n14397 , n14153 );
buf ( n14398 , n14163 );
nand ( n14399 , n14397 , n14398 );
buf ( n14400 , n14399 );
buf ( n14401 , n14400 );
not ( n14402 , n14401 );
buf ( n14403 , n14402 );
nor ( n14404 , n14345 , n14361 );
buf ( n14405 , n14404 );
buf ( n14406 , n14024 );
nand ( n14407 , n14405 , n14406 );
buf ( n14408 , n14407 );
buf ( n14409 , n14408 );
buf ( n14410 , n14395 );
nor ( n14411 , n14409 , n14410 );
buf ( n14412 , n14411 );
buf ( n14413 , n14408 );
not ( n14414 , n14413 );
buf ( n14415 , n14414 );
buf ( n14416 , C0 );
nor ( n14417 , C0 , n14416 );
buf ( n14418 , n14417 );
buf ( n14419 , n13211 );
buf ( n14420 , n12996 );
nand ( n14421 , n14419 , n14420 );
buf ( n14422 , n14421 );
buf ( n14423 , n14422 );
buf ( n14424 , n13203 );
buf ( n14425 , n14424 );
buf ( n14426 , n14425 );
buf ( n14427 , n14426 );
buf ( n14428 , n14426 );
buf ( n14429 , n14422 );
not ( n14430 , n14423 );
not ( n14431 , n14427 );
or ( n14432 , n14430 , n14431 );
or ( n14433 , n14428 , n14429 );
nand ( n14434 , n14432 , n14433 );
buf ( n14435 , n14434 );
buf ( n14436 , n14366 );
buf ( n14437 , n14357 );
nand ( n14438 , n14436 , n14437 );
buf ( n14439 , n14438 );
buf ( n14440 , n14439 );
not ( n14441 , n14440 );
buf ( n14442 , n14441 );
buf ( n14443 , n14323 );
buf ( n14444 , C1 );
nand ( n14445 , n14443 , n14444 );
buf ( n14446 , n14445 );
buf ( n14447 , n14446 );
not ( n14448 , n14447 );
buf ( n14449 , n14448 );
buf ( n14450 , C1 );
buf ( n14451 , n13202 );
buf ( n14452 , n13023 );
and ( n14453 , n14451 , n14452 );
buf ( n14454 , n14453 );
buf ( n14455 , n13191 );
buf ( n14456 , n13187 );
nand ( n14457 , n14455 , n14456 );
buf ( n14458 , n14457 );
buf ( n14459 , C1 );
buf ( n14460 , n14021 );
buf ( n14461 , C1 );
nand ( n14462 , n14460 , n14461 );
buf ( n14463 , n14462 );
xor ( n14464 , n13056 , n13101 );
xor ( n14465 , n14464 , n13135 );
buf ( n14466 , n14465 );
xor ( n14467 , n13119 , n13123 );
xor ( n14468 , n14467 , n13130 );
buf ( n14469 , n14468 );
buf ( n14470 , n14454 );
buf ( n14471 , n13192 );
xor ( n14472 , n14470 , n14471 );
buf ( n14473 , n14472 );
buf ( n14474 , n14458 );
buf ( n14475 , n13174 );
xnor ( n14476 , n14474 , n14475 );
buf ( n14477 , n14476 );
buf ( n14478 , n12000 );
buf ( n14479 , n13558 );
nand ( n14480 , n14478 , n14479 );
buf ( n14481 , n14480 );
buf ( n14482 , n14064 );
buf ( n14483 , C1 );
not ( n14484 , n14482 );
nand ( n14485 , n14484 , n14483 );
buf ( n14486 , n14485 );
xor ( n14487 , n12809 , n12863 );
xor ( n14488 , n14487 , n13215 );
buf ( n14489 , n14488 );
not ( n14490 , n14439 );
nand ( n14491 , n14490 , n13955 );
or ( n14492 , n14072 , n14491 );
not ( n14493 , n13960 );
nor ( n14494 , n14493 , n14442 );
nand ( n14495 , n14072 , n14494 );
nor ( n14496 , n14439 , C0 , n13960 );
nor ( n14497 , C0 , n14496 );
nand ( n14498 , n14492 , n14495 , n14497 );
buf ( n14499 , n14024 );
buf ( n14500 , n14364 );
and ( n14501 , n14499 , n14500 );
buf ( n14502 , n14501 );
and ( n14503 , n14502 , n14342 );
not ( n14504 , n14503 );
not ( n14505 , n14067 );
or ( n14506 , n14504 , n14505 );
nor ( n14507 , C0 , C0 );
nand ( n14508 , n14506 , n14507 );
and ( n14509 , n14508 , n14449 );
not ( n14510 , n14508 );
and ( n14511 , n14510 , n14446 );
nor ( n14512 , n14509 , n14511 );
and ( n14513 , n14387 , C1 );
not ( n14514 , n14415 );
not ( n14515 , n12587 );
not ( n14516 , n13313 );
or ( n14517 , n14515 , n14516 );
nand ( n14518 , n14517 , n13319 );
not ( n14519 , n14518 );
not ( n14520 , n13480 );
or ( n14521 , n14519 , n14520 );
nand ( n14522 , n14521 , n13510 );
and ( n14523 , n14049 , n14522 , n14048 );
nor ( n14524 , n14523 , C0 );
nand ( n14525 , n14066 , n14524 );
not ( n14526 , n14525 );
or ( n14527 , n14514 , n14526 );
nand ( n14528 , n14527 , n14367 );
not ( n14529 , n13142 );
nand ( n14530 , n13170 , n14529 );
or ( n14531 , n14530 , n13139 );
or ( n14532 , n13171 , n13173 );
and ( n14533 , n13171 , n13139 , n14529 );
not ( n14534 , n13139 );
and ( n14535 , n13171 , n14534 , n13142 );
nor ( n14536 , n14533 , n14535 );
nand ( n14537 , n14531 , n14532 , n14536 );
nand ( n14538 , n14071 , n13980 );
not ( n14539 , n14538 );
not ( n14540 , n14486 );
not ( n14541 , n14115 );
nor ( n14542 , n14100 , n14481 );
nand ( n14543 , n14541 , n14542 );
and ( n14544 , n14100 , n14481 );
not ( n14545 , n14100 );
nor ( n14546 , n14481 , n14102 );
and ( n14547 , n14545 , n14546 );
nor ( n14548 , n14544 , n14547 );
and ( n14549 , n14102 , n14481 );
nand ( n14550 , n14549 , n14115 );
nand ( n14551 , n14543 , n14548 , n14550 );
not ( n14552 , n14528 );
and ( n14553 , n14513 , n14450 );
nand ( n14554 , n14552 , n14553 );
nand ( n14555 , n14554 , C1 , C1 );
not ( n14556 , n13999 );
nor ( n14557 , n14556 , n14539 );
nor ( n14558 , n14538 , n14070 , n13999 );
not ( n14559 , n14525 );
and ( n14560 , n14559 , n14540 );
nor ( n14561 , n14560 , C0 );
not ( n14562 , n14561 );
not ( n14563 , n14561 );
or ( n14564 , n14365 , n14385 );
nand ( n14565 , n14564 , n14450 );
xnor ( n14566 , n14565 , n14528 );
and ( n14567 , n10091 , C1 );
not ( n14568 , n10306 );
not ( n14569 , n13570 );
or ( n14570 , n14568 , n14569 );
nand ( n14571 , n10294 , n10303 );
nand ( n14572 , n14570 , n14571 );
and ( n14573 , n14567 , n14572 );
not ( n14574 , n14567 );
and ( n14575 , n13570 , n10306 );
not ( n14576 , n14571 );
nor ( n14577 , n14575 , n14576 );
and ( n14578 , n14574 , n14577 );
nor ( n14579 , n14573 , n14578 );
not ( n14580 , n14412 );
not ( n14581 , n14525 );
or ( n14582 , n14580 , n14581 );
nand ( n14583 , n14582 , n14396 );
and ( n14584 , n14583 , n14365 );
not ( n14585 , n14583 );
and ( n14586 , n14585 , n14322 );
nor ( n14587 , n14584 , n14586 );
and ( n14588 , n14158 , n14403 );
not ( n14589 , n14158 );
and ( n14590 , n14589 , n14400 );
nor ( n14591 , n14588 , n14590 );
nand ( n14592 , n14525 , n14021 );
nand ( n14593 , n14192 , n14187 );
nand ( n14594 , n14592 , n14459 );
nand ( n14595 , C1 , n13999 );
not ( n14596 , n14595 );
and ( n14597 , n14594 , n14596 );
not ( n14598 , n14594 );
and ( n14599 , n14598 , n14595 );
nor ( n14600 , n14597 , n14599 );
nand ( n14601 , n14170 , n14148 );
not ( n14602 , n14601 );
and ( n14603 , n14164 , n14602 );
not ( n14604 , n14164 );
and ( n14605 , n14604 , n14601 );
nor ( n14606 , n14603 , n14605 );
not ( n14607 , n14557 );
or ( n14608 , n14592 , n14607 );
nor ( n14609 , C0 , n14538 );
nand ( n14610 , n14592 , n14609 );
not ( n14611 , n14539 );
and ( n14612 , n14611 , C0 );
nor ( n14613 , n14612 , n14558 );
nand ( n14614 , n14608 , n14610 , n14613 );
nand ( n14615 , n10306 , n14571 );
not ( n14616 , n14615 );
and ( n14617 , n13570 , n14616 );
not ( n14618 , n13570 );
and ( n14619 , n14618 , n14615 );
nor ( n14620 , n14617 , n14619 );
not ( n14621 , n13106 );
not ( n14622 , n401 );
and ( n14623 , n14621 , n14622 );
and ( n14624 , n13106 , n401 );
nor ( n14625 , n14623 , n14624 );
not ( n14626 , n14625 );
not ( n14627 , n13088 );
or ( n14628 , n14626 , n14627 );
or ( n14629 , n13088 , n14625 );
nand ( n14630 , n14628 , n14629 );
not ( n14631 , n14502 );
not ( n14632 , n14067 );
or ( n14633 , n14631 , n14632 );
nand ( n14634 , n14633 , n14418 );
nand ( n14635 , C1 , n14342 );
not ( n14636 , n14635 );
and ( n14637 , n14634 , n14636 );
not ( n14638 , n14634 );
and ( n14639 , n14638 , n14635 );
nor ( n14640 , n14637 , n14639 );
xor ( n14641 , n14559 , n14463 );
buf ( n14642 , n14189 );
buf ( n14643 , n14593 );
xnor ( n14644 , n14642 , n14643 );
buf ( n14645 , n14644 );
not ( C0n , n0 );
and ( C0 , C0n , n0 );
not ( C1n , n0 );
or ( C1 , C1n , n0 );
endmodule
