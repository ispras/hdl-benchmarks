// IWLS benchmark module "decod" printed on Wed May 29 16:32:29 2002
module decod(a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u);
input
  a,
  b,
  c,
  d,
  e;
output
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r,
  s,
  t,
  u;
wire
  \[13] ,
  \[14] ,
  \[15] ,
  n0,
  \[16] ,
  o0,
  \[17] ,
  \[18] ,
  \[19] ,
  \[0] ,
  \[1] ,
  \[2] ,
  \[3] ,
  \[4] ,
  \[5] ,
  \[20] ,
  \[6] ,
  \[21] ,
  \[7] ,
  \[22] ,
  \[8] ,
  \[10] ,
  \[23] ,
  \[9] ,
  \[11] ,
  \[12] ;
assign
  \[13]  = \[18]  & \[17] ,
  \[14]  = \[23]  & \[20] ,
  \[15]  = \[20]  & \[17] ,
  n0 = e & ~a,
  \[16]  = c & b,
  o0 = e & a,
  \[17]  = n0 & ~d,
  \[18]  = c & ~b,
  f = \[0] ,
  g = \[1] ,
  h = \[2] ,
  i = \[3] ,
  j = \[4] ,
  k = \[5] ,
  l = \[6] ,
  m = \[7] ,
  n = \[8] ,
  o = \[9] ,
  \[19]  = ~c & b,
  p = \[10] ,
  q = \[11] ,
  r = \[12] ,
  s = \[13] ,
  t = \[14] ,
  u = \[15] ,
  \[0]  = \[21]  & \[16] ,
  \[1]  = \[22]  & \[16] ,
  \[2]  = \[21]  & \[19] ,
  \[3]  = \[22]  & \[19] ,
  \[4]  = \[21]  & \[18] ,
  \[5]  = \[22]  & \[18] ,
  \[20]  = ~c & ~b,
  \[6]  = \[21]  & \[20] ,
  \[21]  = o0 & d,
  \[7]  = \[22]  & \[20] ,
  \[22]  = o0 & ~d,
  \[8]  = \[23]  & \[16] ,
  \[10]  = \[23]  & \[19] ,
  \[23]  = n0 & d,
  \[9]  = \[17]  & \[16] ,
  \[11]  = \[19]  & \[17] ,
  \[12]  = \[23]  & \[18] ;
endmodule

