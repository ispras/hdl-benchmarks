//NOTE: no-implementation module stub

module DMDbuf (
    input wire [15:0] DMDin,
    output reg [15:0] DMDin1
);

endmodule
