// IWLS benchmark module "MultiplierB_16" printed on Wed May 29 22:12:32 2002
module MultiplierB_16(\1 , \3 , \4 , \5 , \6 , \7 , \8 , \9 , \10 , \11 , \12 , \13 , \14 , \15 , \16 , \17 , \18 , \50 );
input
  \1 ,
  \3 ,
  \4 ,
  \5 ,
  \6 ,
  \7 ,
  \8 ,
  \9 ,
  \10 ,
  \11 ,
  \12 ,
  \13 ,
  \14 ,
  \15 ,
  \16 ,
  \17 ,
  \18 ;
output
  \50 ;
reg
  \2 ,
  \20 ,
  \21 ,
  \22 ,
  \23 ,
  \24 ,
  \25 ,
  \26 ,
  \27 ,
  \28 ,
  \29 ,
  \30 ,
  \31 ,
  \32 ,
  \33 ,
  \34 ,
  \35 ,
  \36 ,
  \37 ,
  \38 ,
  \39 ,
  \40 ,
  \41 ,
  \42 ,
  \43 ,
  \44 ,
  \45 ,
  \46 ,
  \47 ,
  \48 ;
wire
  \[59] ,
  \[60] ,
  \114 ,
  \115 ,
  \116 ,
  \117 ,
  \118 ,
  \119 ,
  \120 ,
  \121 ,
  \122 ,
  \123 ,
  \124 ,
  \125 ,
  \126 ,
  \127 ,
  \128 ,
  \129 ,
  \130 ,
  \131 ,
  \132 ,
  \133 ,
  \134 ,
  \135 ,
  \136 ,
  \137 ,
  \138 ,
  \139 ,
  \140 ,
  \141 ,
  \142 ,
  \143 ,
  \144 ,
  \145 ,
  \146 ,
  \147 ,
  \148 ,
  \149 ,
  \150 ,
  \151 ,
  \152 ,
  \153 ,
  \154 ,
  \155 ,
  \156 ,
  \157 ,
  \158 ,
  \159 ,
  \160 ,
  \161 ,
  \162 ,
  \163 ,
  \164 ,
  \165 ,
  \166 ,
  \167 ,
  \168 ,
  \169 ,
  \170 ,
  \171 ,
  \172 ,
  \173 ,
  \174 ,
  \175 ,
  \176 ,
  \177 ,
  \178 ,
  \179 ,
  \180 ,
  \181 ,
  \182 ,
  \183 ,
  \184 ,
  \185 ,
  \186 ,
  \187 ,
  \188 ,
  \191 ,
  \192 ,
  \194 ,
  \195 ,
  \197 ,
  \198 ,
  \[31] ,
  \[32] ,
  \[33] ,
  \[34] ,
  \[35] ,
  \200 ,
  \201 ,
  \203 ,
  \204 ,
  \206 ,
  \207 ,
  \209 ,
  \[36] ,
  \210 ,
  \212 ,
  \213 ,
  \215 ,
  \216 ,
  \218 ,
  \219 ,
  \[37] ,
  \221 ,
  \222 ,
  \224 ,
  \225 ,
  \227 ,
  \228 ,
  \[38] ,
  \230 ,
  \231 ,
  \233 ,
  \234 ,
  \235 ,
  \237 ,
  \239 ,
  \[39] ,
  \241 ,
  \243 ,
  \245 ,
  \247 ,
  \249 ,
  \251 ,
  \253 ,
  \255 ,
  \257 ,
  \259 ,
  \261 ,
  \263 ,
  \265 ,
  \[40] ,
  \[41] ,
  \[42] ,
  \[43] ,
  \[44] ,
  \[45] ,
  \[46] ,
  \[47] ,
  \[48] ,
  \[49] ,
  \[50] ,
  \[51] ,
  \[52] ,
  \[53] ,
  \[54] ,
  \[55] ,
  \[56] ,
  \[57] ,
  \[58] ;
assign
  \[59]  = \183 ,
  \[60]  = \188 ,
  \114  = (~\265  & \191 ) | (\265  & ~\191 ),
  \115  = \265  & \20 ,
  \116  = \265  & \34 ,
  \117  = \20  & \34 ,
  \118  = \192  | \117 ,
  \119  = (~\263  & \194 ) | (\263  & ~\194 ),
  \120  = \263  & \21 ,
  \121  = \263  & \35 ,
  \122  = \21  & \35 ,
  \123  = \195  | \122 ,
  \124  = (~\261  & \197 ) | (\261  & ~\197 ),
  \125  = \261  & \22 ,
  \126  = \261  & \36 ,
  \127  = \22  & \36 ,
  \128  = \198  | \127 ,
  \129  = (~\259  & \200 ) | (\259  & ~\200 ),
  \130  = \259  & \23 ,
  \131  = \259  & \37 ,
  \132  = \23  & \37 ,
  \133  = \201  | \132 ,
  \134  = (~\257  & \203 ) | (\257  & ~\203 ),
  \135  = \257  & \24 ,
  \136  = \257  & \38 ,
  \137  = \24  & \38 ,
  \138  = \204  | \137 ,
  \139  = (~\255  & \206 ) | (\255  & ~\206 ),
  \140  = \255  & \25 ,
  \141  = \255  & \39 ,
  \142  = \25  & \39 ,
  \143  = \207  | \142 ,
  \144  = (~\253  & \209 ) | (\253  & ~\209 ),
  \145  = \253  & \26 ,
  \146  = \253  & \40 ,
  \147  = \26  & \40 ,
  \148  = \210  | \147 ,
  \149  = (~\251  & \212 ) | (\251  & ~\212 ),
  \150  = \251  & \27 ,
  \151  = \251  & \41 ,
  \152  = \27  & \41 ,
  \153  = \213  | \152 ,
  \154  = (~\249  & \215 ) | (\249  & ~\215 ),
  \155  = \249  & \28 ,
  \156  = \249  & \42 ,
  \157  = \28  & \42 ,
  \158  = \216  | \157 ,
  \159  = (~\247  & \218 ) | (\247  & ~\218 ),
  \160  = \247  & \29 ,
  \161  = \247  & \43 ,
  \162  = \29  & \43 ,
  \163  = \219  | \162 ,
  \164  = (~\245  & \221 ) | (\245  & ~\221 ),
  \165  = \245  & \30 ,
  \166  = \245  & \44 ,
  \167  = \30  & \44 ,
  \168  = \222  | \167 ,
  \169  = (~\243  & \224 ) | (\243  & ~\224 ),
  \170  = \243  & \31 ,
  \171  = \243  & \45 ,
  \172  = \31  & \45 ,
  \173  = \225  | \172 ,
  \174  = (~\241  & \227 ) | (\241  & ~\227 ),
  \175  = \241  & \32 ,
  \176  = \241  & \46 ,
  \177  = \32  & \46 ,
  \178  = \228  | \177 ,
  \179  = (~\239  & \230 ) | (\239  & ~\230 ),
  \180  = \239  & \33 ,
  \181  = \239  & \47 ,
  \182  = \33  & \47 ,
  \183  = \231  | \182 ,
  \184  = (~\237  & \233 ) | (\237  & ~\233 ),
  \185  = \237  & \2 ,
  \186  = \237  & \48 ,
  \187  = \2  & \48 ,
  \188  = \234  | \187 ,
  \191  = (~\20  & \34 ) | (\20  & ~\34 ),
  \192  = \116  | \115 ,
  \194  = (~\21  & \35 ) | (\21  & ~\35 ),
  \195  = \121  | \120 ,
  \197  = (~\22  & \36 ) | (\22  & ~\36 ),
  \198  = \126  | \125 ,
  \[31]  = \235 ,
  \[32]  = \119 ,
  \[33]  = \124 ,
  \[34]  = \129 ,
  \[35]  = \134 ,
  \200  = (~\23  & \37 ) | (\23  & ~\37 ),
  \201  = \131  | \130 ,
  \203  = (~\24  & \38 ) | (\24  & ~\38 ),
  \204  = \136  | \135 ,
  \206  = (~\25  & \39 ) | (\25  & ~\39 ),
  \207  = \141  | \140 ,
  \209  = (~\26  & \40 ) | (\26  & ~\40 ),
  \[36]  = \139 ,
  \210  = \146  | \145 ,
  \212  = (~\27  & \41 ) | (\27  & ~\41 ),
  \213  = \151  | \150 ,
  \215  = (~\28  & \42 ) | (\28  & ~\42 ),
  \216  = \156  | \155 ,
  \218  = (~\29  & \43 ) | (\29  & ~\43 ),
  \219  = \161  | \160 ,
  \[37]  = \144 ,
  \221  = (~\30  & \44 ) | (\30  & ~\44 ),
  \222  = \166  | \165 ,
  \224  = (~\31  & \45 ) | (\31  & ~\45 ),
  \225  = \171  | \170 ,
  \227  = (~\32  & \46 ) | (\32  & ~\46 ),
  \228  = \176  | \175 ,
  \[38]  = \149 ,
  \230  = (~\33  & \47 ) | (\33  & ~\47 ),
  \231  = \181  | \180 ,
  \233  = (~\2  & \48 ) | (\2  & ~\48 ),
  \234  = \186  | \185 ,
  \235  = \18  & \1 ,
  \237  = \17  & \1 ,
  \239  = \16  & \1 ,
  \[39]  = \154 ,
  \241  = \15  & \1 ,
  \243  = \14  & \1 ,
  \245  = \13  & \1 ,
  \247  = \12  & \1 ,
  \249  = \11  & \1 ,
  \251  = \10  & \1 ,
  \253  = \9  & \1 ,
  \255  = \8  & \1 ,
  \257  = \7  & \1 ,
  \259  = \6  & \1 ,
  \261  = \5  & \1 ,
  \263  = \4  & \1 ,
  \265  = \3  & \1 ,
  \[40]  = \159 ,
  \[41]  = \164 ,
  \[42]  = \169 ,
  \[43]  = \174 ,
  \[44]  = \179 ,
  \[45]  = \184 ,
  \[46]  = \118 ,
  \[47]  = \123 ,
  \[48]  = \128 ,
  \[49]  = \133 ,
  \50  = \114 ,
  \[50]  = \138 ,
  \[51]  = \143 ,
  \[52]  = \148 ,
  \[53]  = \153 ,
  \[54]  = \158 ,
  \[55]  = \163 ,
  \[56]  = \168 ,
  \[57]  = \173 ,
  \[58]  = \178 ;
always begin
  \2  = \[31] ;
  \20  = \[32] ;
  \21  = \[33] ;
  \22  = \[34] ;
  \23  = \[35] ;
  \24  = \[36] ;
  \25  = \[37] ;
  \26  = \[38] ;
  \27  = \[39] ;
  \28  = \[40] ;
  \29  = \[41] ;
  \30  = \[42] ;
  \31  = \[43] ;
  \32  = \[44] ;
  \33  = \[45] ;
  \34  = \[46] ;
  \35  = \[47] ;
  \36  = \[48] ;
  \37  = \[49] ;
  \38  = \[50] ;
  \39  = \[51] ;
  \40  = \[52] ;
  \41  = \[53] ;
  \42  = \[54] ;
  \43  = \[55] ;
  \44  = \[56] ;
  \45  = \[57] ;
  \46  = \[58] ;
  \47  = \[59] ;
  \48  = \[60] ;
end
initial begin
  \2  = 0;
  \20  = 0;
  \21  = 0;
  \22  = 0;
  \23  = 0;
  \24  = 0;
  \25  = 0;
  \26  = 0;
  \27  = 0;
  \28  = 0;
  \29  = 0;
  \30  = 0;
  \31  = 0;
  \32  = 0;
  \33  = 0;
  \34  = 0;
  \35  = 0;
  \36  = 0;
  \37  = 0;
  \38  = 0;
  \39  = 0;
  \40  = 0;
  \41  = 0;
  \42  = 0;
  \43  = 0;
  \44  = 0;
  \45  = 0;
  \46  = 0;
  \47  = 0;
  \48  = 0;
end
endmodule

