module GtCLK_NOT ( Z, A );

input A;

output Z;

GTECH_NOT Gtclk1 (.Z(Z), .A(A));

endmodule
