//NOTE: no-implementation module stub

module GTECH_NOR2 (
    output Z,
    input A,
    input B
);

endmodule
