// IWLS benchmark module "pcler8_cl" printed on Wed May 29 17:28:07 2002
module pcler8_cl(a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, \x , y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0);
input
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r,
  s,
  t,
  u,
  v,
  w,
  \x ,
  y,
  z,
  a0;
output
  k0,
  l0,
  m0,
  n0,
  o0,
  p0,
  q0,
  r0,
  b0,
  c0,
  d0,
  e0,
  f0,
  g0,
  h0,
  i0,
  j0;
wire
  \[13] ,
  \[14] ,
  \[15] ,
  \[16] ,
  \[17] ,
  \[18] ,
  \[19] ,
  \[0] ,
  a2,
  \[1] ,
  b2,
  \[2] ,
  \[3] ,
  \[4] ,
  \[5] ,
  \[6] ,
  \[7] ,
  \[8] ,
  \[10] ,
  \[9] ,
  \[11] ,
  \[12] ;
assign
  k0 = \[9] ,
  \[13]  = (~\[19]  & (~b2 & (a2 & w))) | ((~b2 & (a2 & \x )) | ((\[0]  & p) | \[5] )),
  l0 = \[10] ,
  \[14]  = (~b2 & (y & a2)) | ((b2 & (~y & a2)) | ((q & \[0] ) | \[6] )),
  m0 = \[11] ,
  \[15]  = (~\[18]  & (a2 & ~z)) | ((\[18]  & (a2 & z)) | ((\[0]  & r) | \[7] )),
  n0 = \[12] ,
  \[16]  = (~\[18]  & (a2 & (~\[0]  & z))) | ((a2 & (~\[0]  & a0)) | ((\[0]  & s) | \[8] )),
  o0 = \[13] ,
  \[17]  = ~u | ~t,
  p0 = \[14] ,
  \[18]  = ~b2 | ~y,
  q0 = \[15] ,
  \[19]  = \[17]  | ~v,
  r0 = \[16] ,
  \[0]  = ~\[18]  & (a2 & (a0 & z)),
  a2 = ~k & (j & ~i),
  \[1]  = i & a,
  b0 = \[0] ,
  b2 = ~\[19]  & (\x  & w),
  \[2]  = i & b,
  c0 = \[1] ,
  \[3]  = i & c,
  d0 = \[2] ,
  \[4]  = i & d,
  e0 = \[3] ,
  \[5]  = i & e,
  f0 = \[4] ,
  \[6]  = i & f,
  g0 = \[5] ,
  \[7]  = i & g,
  h0 = \[6] ,
  \[8]  = i & h,
  \[10]  = (~u & (t & a2)) | ((u & (~t & a2)) | ((m & \[0] ) | \[2] )),
  i0 = \[7] ,
  \[9]  = (a2 & ~t) | ((\[0]  & l) | \[1] ),
  \[11]  = (~\[17]  & (a2 & ~v)) | ((\[17]  & (a2 & v)) | ((\[0]  & n) | \[3] )),
  j0 = \[8] ,
  \[12]  = (~\[19]  & (a2 & ~w)) | ((\[19]  & (a2 & w)) | ((\[0]  & o) | \[4] ));
endmodule

