module top ( g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 );
input g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 ;
output g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 ;

wire n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , 
     n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
     n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , 
     n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , 
     n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , 
     n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , 
     n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
     n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , 
     n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , 
     n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , 
     n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
     n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
     n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
     n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
     n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
     n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
     n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
     n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
     n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
     n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
     n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
     n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
     n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , 
     n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , 
     n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , 
     n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , 
     n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , 
     n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , 
     n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , 
     n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , 
     n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , 
     n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , 
     n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , 
     n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , 
     n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , 
     n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , 
     n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , 
     n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , 
     n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , 
     n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 ;
buf ( n1 , g0 );
buf ( n2 , g1 );
buf ( n3 , g2 );
buf ( n4 , g3 );
buf ( n5 , g4 );
buf ( n6 , g5 );
buf ( n7 , g6 );
buf ( n8 , g7 );
buf ( n9 , g8 );
buf ( n10 , g9 );
buf ( n11 , g10 );
buf ( n12 , g11 );
buf ( n13 , g12 );
buf ( n14 , g13 );
buf ( n15 , g14 );
buf ( n16 , g15 );
buf ( n17 , g16 );
buf ( n18 , g17 );
buf ( n19 , g18 );
buf ( n20 , g19 );
buf ( n21 , g20 );
buf ( n22 , g21 );
buf ( n23 , g22 );
buf ( n24 , g23 );
buf ( n25 , g24 );
buf ( g25 , n26 );
buf ( g26 , n27 );
buf ( g27 , n28 );
buf ( g28 , n29 );
buf ( g29 , n30 );
buf ( g30 , n31 );
buf ( g31 , n32 );
buf ( g32 , n33 );
buf ( g33 , n34 );
buf ( g34 , n35 );
buf ( g35 , n36 );
buf ( g36 , n37 );
buf ( g37 , n38 );
buf ( g38 , n39 );
buf ( g39 , n40 );
buf ( g40 , n41 );
buf ( g41 , n42 );
buf ( g42 , n43 );
buf ( g43 , n44 );
buf ( g44 , n45 );
buf ( g45 , n46 );
buf ( g46 , n47 );
buf ( g47 , n48 );
buf ( g48 , n49 );
buf ( g49 , n50 );
buf ( g50 , n51 );
buf ( g51 , n52 );
buf ( g52 , n53 );
buf ( g53 , n54 );
buf ( g54 , n55 );
buf ( g55 , n56 );
buf ( g56 , n57 );
buf ( g57 , n58 );
buf ( g58 , n59 );
buf ( g59 , n60 );
buf ( g60 , n61 );
buf ( g61 , n62 );
buf ( g62 , n63 );
buf ( g63 , n64 );
buf ( n26 , n351 );
buf ( n27 , n382 );
buf ( n28 , n383 );
buf ( n29 , n378 );
buf ( n30 , n377 );
buf ( n31 , n394 );
buf ( n32 , n387 );
buf ( n33 , n288 );
buf ( n34 , n393 );
buf ( n35 , n304 );
buf ( n36 , n390 );
buf ( n37 , n85 );
buf ( n38 , n396 );
buf ( n39 , n304 );
buf ( n40 , n386 );
buf ( n41 , n395 );
buf ( n42 , n397 );
buf ( n43 , n175 );
buf ( n44 , n389 );
buf ( n45 , 1'b0 );
buf ( n46 , 1'b0 );
buf ( n47 , n398 );
buf ( n48 , n333 );
buf ( n49 , 1'b0 );
buf ( n50 , 1'b0 );
buf ( n51 , n398 );
buf ( n52 , n247 );
buf ( n53 , 1'b0 );
buf ( n54 , 1'b0 );
buf ( n55 , n398 );
buf ( n56 , n309 );
buf ( n57 , 1'b0 );
buf ( n58 , 1'b0 );
buf ( n59 , n398 );
buf ( n60 , n376 );
buf ( n61 , 1'b0 );
buf ( n62 , 1'b0 );
buf ( n63 , n398 );
buf ( n64 , n177 );
not ( n77 , n14 );
not ( n78 , n77 );
not ( n79 , n22 );
nor ( n80 , n25 , n24 );
nand ( n81 , n79 , n80 , n21 );
nor ( n82 , n78 , n81 );
nand ( n83 , n22 , n23 );
nand ( n84 , n21 , n25 );
nor ( n85 , n83 , n84 );
or ( n86 , n82 , n85 );
not ( n87 , n16 );
nand ( n88 , n86 , n87 );
not ( n89 , n24 );
nor ( n90 , n89 , n25 );
not ( n91 , n90 );
not ( n92 , n21 );
not ( n93 , n25 );
nand ( n94 , n92 , n93 , n17 );
nand ( n95 , n23 , n25 );
nand ( n96 , n94 , n95 );
nor ( n97 , n15 , n18 , n16 , n22 );
not ( n98 , n24 );
nand ( n99 , n98 , n25 );
nand ( n100 , n91 , n96 , n97 , n99 );
not ( n101 , n16 );
not ( n102 , n14 );
nor ( n103 , n102 , n18 );
nor ( n104 , n21 , n22 );
nor ( n105 , n24 , n25 );
nand ( n106 , n101 , n103 , n104 , n105 );
nand ( n107 , n88 , n100 , n106 );
not ( n108 , n25 );
nand ( n109 , n108 , n24 );
nand ( n110 , n109 , n83 );
nand ( n111 , n110 , n77 );
nor ( n112 , n23 , n24 );
not ( n113 , n112 );
not ( n114 , n22 );
nand ( n115 , n23 , n24 );
nand ( n116 , n113 , n114 , n115 , n25 );
and ( n117 , n111 , n116 );
nor ( n118 , n13 , n16 );
not ( n119 , n118 );
nor ( n120 , n117 , n119 );
nor ( n121 , n107 , n120 );
not ( n122 , n23 );
not ( n123 , n25 );
nand ( n124 , n123 , n12 );
nor ( n125 , n122 , n124 );
not ( n126 , n24 );
or ( n127 , n126 , n22 );
not ( n128 , n21 );
nand ( n129 , n8 , n24 );
nand ( n130 , n128 , n129 );
nand ( n131 , n127 , n130 );
nand ( n132 , n125 , n131 );
not ( n133 , n25 );
nand ( n134 , n21 , n22 );
nor ( n135 , n133 , n134 );
nor ( n136 , n134 , n14 );
nor ( n137 , n135 , n136 );
nand ( n138 , n12 , n22 );
nor ( n139 , n138 , n21 , n23 );
not ( n140 , n4 );
not ( n141 , n6 );
and ( n142 , n140 , n141 );
nor ( n143 , n4 , n5 );
nor ( n144 , n142 , n143 );
nand ( n145 , n139 , n90 , n144 );
nand ( n146 , n132 , n137 , n145 );
nand ( n147 , n146 , n118 );
and ( n148 , n24 , n19 );
not ( n149 , n24 );
not ( n150 , n21 );
nand ( n151 , n150 , n14 );
and ( n152 , n149 , n151 );
nor ( n153 , n148 , n152 );
not ( n154 , n23 );
nand ( n155 , n154 , n22 , n25 );
not ( n156 , n155 );
and ( n157 , n153 , n156 , n87 );
nor ( n158 , n83 , n12 );
and ( n159 , n158 , n118 , n25 );
nor ( n160 , n157 , n159 );
not ( n161 , n10 );
nor ( n162 , n161 , n24 );
nor ( n163 , n162 , n23 );
not ( n164 , n163 );
not ( n165 , n22 );
nand ( n166 , n165 , n12 );
nand ( n167 , n166 , n126 );
nor ( n168 , n22 , n25 );
nor ( n169 , n12 , n25 );
nor ( n170 , n168 , n169 );
nand ( n171 , n164 , n167 , n170 );
not ( n172 , n21 );
nor ( n173 , n172 , n22 );
not ( n174 , n173 );
nor ( n175 , n174 , n99 , n23 );
nand ( n176 , n171 , n87 , n175 );
nand ( n177 , n121 , n147 , n160 , n176 );
not ( n178 , n2 );
not ( n179 , n7 );
nand ( n180 , n178 , n179 , n3 , n9 );
not ( n181 , n180 );
not ( n182 , n99 );
not ( n183 , n166 );
nand ( n184 , n181 , n182 , n183 , n23 );
nand ( n185 , n22 , n169 );
not ( n186 , n185 );
not ( n187 , n112 );
and ( n188 , n186 , n187 );
not ( n189 , n23 );
nand ( n190 , n189 , n22 , n21 );
not ( n191 , n190 );
nor ( n192 , n188 , n191 );
not ( n193 , n21 );
nand ( n194 , n193 , n23 );
not ( n195 , n194 );
nand ( n196 , n99 , n129 , n12 );
nand ( n197 , n195 , n196 );
or ( n198 , n4 , n5 );
not ( n199 , n22 );
nor ( n200 , n199 , n23 );
nand ( n201 , n198 , n200 , n90 );
nand ( n202 , n184 , n192 , n197 , n201 );
not ( n203 , n13 );
nand ( n204 , n203 , n14 );
nor ( n205 , n204 , n16 );
nand ( n206 , n202 , n205 );
not ( n207 , n25 );
nand ( n208 , n23 , n24 );
nor ( n209 , n207 , n208 , n22 );
nor ( n210 , n21 , n24 );
nor ( n211 , n22 , n25 );
nand ( n212 , n210 , n211 );
not ( n213 , n212 );
nor ( n214 , n209 , n213 );
not ( n215 , n214 );
not ( n216 , n18 );
nor ( n217 , n216 , n16 );
and ( n218 , n215 , n217 );
nor ( n219 , n22 , n23 );
nand ( n220 , n219 , n24 );
not ( n221 , n220 );
nand ( n222 , n221 , n118 );
nand ( n223 , n2 , n3 , n7 , n9 );
nand ( n224 , n12 , n25 );
nor ( n225 , n223 , n224 );
not ( n226 , n21 );
nor ( n227 , n226 , n14 );
nor ( n228 , n225 , n227 );
nor ( n229 , n222 , n228 );
nor ( n230 , n218 , n229 );
not ( n231 , n84 );
and ( n232 , n183 , n231 , n112 );
and ( n233 , n232 , n87 , n10 );
not ( n234 , n84 );
not ( n235 , n13 );
and ( n236 , n234 , n235 );
nor ( n237 , n19 , n25 );
and ( n238 , n210 , n237 );
nor ( n239 , n236 , n238 );
not ( n240 , n200 );
nor ( n241 , n239 , n240 , n16 );
nor ( n242 , n233 , n241 );
and ( n243 , n156 , n153 , n87 );
nand ( n244 , n103 , n104 , n105 );
nor ( n245 , n244 , n16 );
nor ( n246 , n243 , n245 );
nand ( n247 , n206 , n230 , n242 , n246 );
not ( n248 , n194 );
not ( n249 , n203 );
and ( n250 , n248 , n249 );
not ( n251 , n22 );
nand ( n252 , n251 , n25 );
not ( n253 , n252 );
not ( n254 , n23 );
nor ( n255 , n254 , n203 , n24 );
and ( n256 , n253 , n255 );
nor ( n257 , n250 , n256 );
not ( n258 , n124 );
nand ( n259 , n258 , n191 , n14 );
nand ( n260 , n221 , n227 );
nand ( n261 , n221 , n13 );
nand ( n262 , n257 , n259 , n260 , n261 );
not ( n263 , n23 );
nand ( n264 , n263 , n173 );
not ( n265 , n24 );
nand ( n266 , n265 , n134 );
nor ( n267 , n203 , n25 );
nand ( n268 , n264 , n266 , n267 );
not ( n269 , n23 );
nand ( n270 , n269 , n22 , n21 );
not ( n271 , n270 );
not ( n272 , n203 );
and ( n273 , n271 , n272 );
and ( n274 , n156 , n227 );
nor ( n275 , n273 , n274 );
nand ( n276 , n268 , n275 );
nor ( n277 , n262 , n276 );
not ( n278 , n6 );
nand ( n279 , n4 , n5 );
nand ( n280 , n278 , n279 , n14 , n12 );
nor ( n281 , n201 , n280 );
not ( n282 , n14 );
not ( n283 , n81 );
not ( n284 , n283 );
or ( n285 , n282 , n284 );
not ( n286 , n11 );
nand ( n287 , n286 , n21 , n22 );
nor ( n288 , n287 , n95 );
not ( n289 , n288 );
nand ( n290 , n285 , n289 );
nor ( n291 , n281 , n232 , n290 );
not ( n292 , n12 );
not ( n293 , n22 );
or ( n294 , n292 , n293 );
nand ( n295 , n21 , n24 );
nand ( n296 , n294 , n295 );
and ( n297 , n296 , n25 );
nand ( n298 , n12 , n24 );
nand ( n299 , n298 , n23 );
nor ( n300 , n297 , n299 );
not ( n301 , n135 );
and ( n302 , n300 , n301 , n14 );
not ( n303 , n209 );
not ( n304 , n303 );
nor ( n305 , n15 , n18 , n17 );
and ( n306 , n304 , n305 );
nor ( n307 , n302 , n306 );
and ( n308 , n277 , n291 , n307 );
nor ( n309 , n308 , n16 );
not ( n310 , n24 );
not ( n311 , n305 );
or ( n312 , n310 , n311 );
nand ( n313 , n312 , n21 );
and ( n314 , n313 , n253 );
nand ( n315 , n180 , n114 );
not ( n316 , n124 );
nor ( n317 , n316 , n204 );
and ( n318 , n315 , n317 );
not ( n319 , n24 );
nand ( n320 , n319 , n23 );
nor ( n321 , n318 , n320 );
nor ( n322 , n314 , n321 );
and ( n323 , n171 , n21 );
not ( n324 , n168 );
not ( n325 , n23 );
nand ( n326 , n325 , n93 , n143 );
nand ( n327 , n324 , n326 , n194 );
not ( n328 , n298 );
and ( n329 , n327 , n328 );
nor ( n330 , n323 , n329 );
nand ( n331 , n110 , n204 );
and ( n332 , n322 , n330 , n331 );
nor ( n333 , n332 , n16 );
not ( n334 , n325 );
not ( n335 , n173 );
or ( n336 , n334 , n335 );
nand ( n337 , n336 , n266 );
or ( n338 , n337 , n25 );
not ( n339 , n252 );
not ( n340 , n320 );
and ( n341 , n339 , n340 );
not ( n342 , n194 );
nor ( n343 , n341 , n342 );
nand ( n344 , n338 , n343 );
nand ( n345 , n220 , n270 );
nor ( n346 , n344 , n345 );
or ( n347 , n346 , n203 );
and ( n348 , n344 , n77 );
not ( n349 , n244 );
nor ( n350 , n348 , n349 );
nand ( n351 , n347 , n350 );
not ( n352 , n305 );
nor ( n353 , n352 , n303 );
not ( n354 , n19 );
nand ( n355 , n354 , n24 );
nor ( n356 , n155 , n355 );
or ( n357 , n353 , n356 , n288 );
nand ( n358 , n357 , n87 );
not ( n359 , n134 );
nand ( n360 , n359 , n125 );
nand ( n361 , n158 , n24 );
not ( n362 , n224 );
nand ( n363 , n362 , n342 );
nand ( n364 , n360 , n361 , n363 );
not ( n365 , n12 );
not ( n366 , n223 );
not ( n367 , n366 );
or ( n368 , n365 , n367 );
nand ( n369 , n368 , n221 );
not ( n370 , n83 );
nand ( n371 , n370 , n8 );
nand ( n372 , n371 , n90 );
nand ( n373 , n369 , n372 );
or ( n374 , n364 , n373 );
nand ( n375 , n374 , n205 );
nand ( n376 , n358 , n375 );
not ( n377 , n346 );
nor ( n378 , n214 , n216 );
or ( n379 , n5 , n6 );
not ( n380 , n204 );
nand ( n381 , n379 , n380 );
nor ( n382 , n145 , n381 );
nor ( n383 , n228 , n220 , n13 );
not ( n384 , n10 );
not ( n385 , n232 );
nor ( n386 , n384 , n385 );
not ( n387 , n360 );
nand ( n388 , n216 , n15 );
nor ( n389 , n212 , n388 , n14 );
and ( n390 , n85 , n11 );
nand ( n391 , n112 , n168 );
nand ( n392 , n14 , n21 );
nor ( n393 , n391 , n392 );
nor ( n394 , n190 , n124 );
not ( n395 , n391 );
nor ( n396 , n252 , n21 );
not ( n397 , n385 );
and ( n398 , n1 , n20 );
endmodule
