// IWLS benchmark module "i2" printed on Wed May 29 16:38:44 2002
module i2(\V62(1) , \V30(31) , \V30(29) , \V30(27) , \V30(25) , \V30(23) , \V30(21) , \V30(19) , \V30(17) , \V30(15) , \V30(13) , \V30(11) , \V30(9) , \V30(7) , \V30(5) , \V30(3) , \V30(2) , \V30(4) , \V30(6) , \V30(8) , \V30(10) , \V30(12) , \V30(14) , \V30(16) , \V30(18) , \V30(20) , \V30(22) , \V30(24) , \V30(26) , \V30(28) , \V30(30) , \V62(0) , \V64(0) , \V62(31) , \V62(29) , \V62(27) , \V62(25) , \V62(23) , \V62(21) , \V62(19) , \V62(17) , \V62(15) , \V62(13) , \V62(11) , \V62(9) , \V62(7) , \V62(5) , \V62(3) , \V62(2) , \V62(4) , \V62(6) , \V62(8) , \V62(10) , \V62(12) , \V62(14) , \V62(16) , \V62(18) , \V62(20) , \V62(22) , \V62(24) , \V62(26) , \V62(28) , \V62(30) , \V63(0) , \V126(1) , \V94(31) , \V94(29) , \V94(27) , \V94(25) , \V94(23) , \V94(21) , \V94(19) , \V94(17) , \V94(15) , \V94(13) , \V94(11) , \V94(9) , \V94(7) , \V94(5) , \V94(3) , \V94(2) , \V94(4) , \V94(6) , \V94(8) , \V94(10) , \V94(12) , \V94(14) , \V94(16) , \V94(18) , \V94(20) , \V94(22) , \V94(24) , \V94(26) , \V94(28) , \V94(30) , \V126(0) , \V128(0) , \V126(31) , \V126(29) , \V126(27) , \V126(25) , \V126(23) , \V126(21) , \V126(19) , \V126(17) , \V126(15) , \V126(13) , \V126(11) , \V126(9) , \V126(7) , \V126(5) , \V126(3) , \V126(2) , \V126(4) , \V126(6) , \V126(8) , \V126(10) , \V126(12) , \V126(14) , \V126(16) , \V126(18) , \V126(20) , \V126(22) , \V126(24) , \V126(26) , \V126(28) , \V126(30) , \V127(0) , \V201(0) , \V129(0) , \V201(1) , \V130(0) , \V176(1) , \V144(31) , \V144(29) , \V144(27) , \V144(25) , \V144(23) , \V144(21) , \V144(19) , \V144(18) , \V144(20) , \V144(22) , \V144(24) , \V144(26) , \V144(28) , \V144(30) , \V176(0) , \V176(17) , \V176(15) , \V176(13) , \V176(11) , \V176(9) , \V176(7) , \V176(5) , \V176(3) , \V176(2) , \V176(4) , \V176(6) , \V176(8) , \V176(10) , \V176(12) , \V176(14) , \V176(16) , \V178(1) , \V176(31) , \V176(29) , \V176(27) , \V176(25) , \V176(23) , \V176(21) , \V176(19) , \V176(18) , \V176(20) , \V176(22) , \V176(24) , \V176(26) , \V176(28) , \V176(30) , \V178(0) , \V201(3) , \V201(2) , \V188(25) , \V188(23) , \V188(22) , \V188(24) , \V188(29) , \V188(27) , \V188(26) , \V188(28) , \V190(1) , \V188(31) , \V188(30) , \V190(0) , \V201(5) , \V201(4) , \V201(7) , \V191(31) , \V201(6) , \V193(0) , \V193(1) , \V202(0) );
input
  \V126(17) ,
  \V144(21) ,
  \V30(29) ,
  \V126(1) ,
  \V126(16) ,
  \V144(20) ,
  \V30(28) ,
  \V126(0) ,
  \V126(19) ,
  \V144(23) ,
  \V126(18) ,
  \V144(22) ,
  \V62(13) ,
  \V144(25) ,
  \V62(12) ,
  \V191(31) ,
  \V144(24) ,
  \V62(15) ,
  \V94(31) ,
  \V62(14) ,
  \V126(7) ,
  \V94(30) ,
  \V126(6) ,
  \V144(19) ,
  \V30(31) ,
  \V201(3) ,
  \V126(9) ,
  \V144(18) ,
  \V62(11) ,
  \V30(30) ,
  \V201(2) ,
  \V126(8) ,
  \V126(11) ,
  \V62(10) ,
  \V201(5) ,
  \V126(10) ,
  \V201(4) ,
  \V126(13) ,
  \V176(31) ,
  \V126(12) ,
  \V176(30) ,
  \V94(2) ,
  \V126(15) ,
  \V63(0) ,
  \V201(1) ,
  \V94(3) ,
  \V126(14) ,
  \V62(17) ,
  \V201(0) ,
  \V94(4) ,
  \V193(1) ,
  \V62(16) ,
  \V94(5) ,
  \V193(0) ,
  \V62(19) ,
  \V94(6) ,
  \V62(18) ,
  \V176(3) ,
  \V94(7) ,
  \V62(23) ,
  \V176(2) ,
  \V94(8) ,
  \V129(0) ,
  \V62(22) ,
  \V176(5) ,
  \V201(7) ,
  \V94(9) ,
  \V62(25) ,
  \V176(4) ,
  \V201(6) ,
  \V62(24) ,
  \V176(27) ,
  \V176(26) ,
  \V176(1) ,
  \V176(29) ,
  \V62(21) ,
  \V176(0) ,
  \V176(28) ,
  \V62(20) ,
  \V188(31) ,
  \V176(7) ,
  \V62(0) ,
  \V188(30) ,
  \V62(27) ,
  \V176(6) ,
  \V62(1) ,
  \V62(26) ,
  \V176(9) ,
  \V176(21) ,
  \V62(2) ,
  \V62(29) ,
  \V176(8) ,
  \V176(20) ,
  \V62(3) ,
  \V62(28) ,
  \V176(23) ,
  \V62(4) ,
  \V176(22) ,
  \V62(5) ,
  \V94(13) ,
  \V128(0) ,
  \V176(25) ,
  \V62(6) ,
  \V94(12) ,
  \V176(24) ,
  \V62(7) ,
  \V94(15) ,
  \V30(13) ,
  \V130(0) ,
  \V176(17) ,
  \V62(8) ,
  \V94(14) ,
  \V30(12) ,
  \V176(16) ,
  \V62(9) ,
  \V188(27) ,
  \V30(15) ,
  \V176(19) ,
  \V188(26) ,
  \V62(31) ,
  \V30(14) ,
  \V126(31) ,
  \V176(18) ,
  \V94(11) ,
  \V188(29) ,
  \V62(30) ,
  \V126(30) ,
  \V94(10) ,
  \V188(28) ,
  \V30(11) ,
  \V30(10) ,
  \V144(31) ,
  \V94(17) ,
  \V176(11) ,
  \V144(30) ,
  \V94(16) ,
  \V176(10) ,
  \V94(19) ,
  \V30(17) ,
  \V176(13) ,
  \V94(18) ,
  \V30(16) ,
  \V176(12) ,
  \V126(27) ,
  \V94(23) ,
  \V188(23) ,
  \V30(2) ,
  \V30(19) ,
  \V176(15) ,
  \V126(26) ,
  \V94(22) ,
  \V188(22) ,
  \V30(3) ,
  \V127(0) ,
  \V30(18) ,
  \V176(14) ,
  \V126(29) ,
  \V94(25) ,
  \V188(25) ,
  \V30(4) ,
  \V30(23) ,
  \V126(28) ,
  \V94(24) ,
  \V188(24) ,
  \V30(5) ,
  \V30(22) ,
  \V30(6) ,
  \V30(25) ,
  \V30(7) ,
  \V30(24) ,
  \V144(27) ,
  \V94(21) ,
  \V30(8) ,
  \V144(26) ,
  \V94(20) ,
  \V30(9) ,
  \V178(1) ,
  \V144(29) ,
  \V178(0) ,
  \V30(21) ,
  \V144(28) ,
  \V30(20) ,
  \V126(21) ,
  \V126(3) ,
  \V126(20) ,
  \V126(2) ,
  \V126(23) ,
  \V94(27) ,
  \V126(5) ,
  \V126(22) ,
  \V94(26) ,
  \V64(0) ,
  \V126(4) ,
  \V126(25) ,
  \V94(29) ,
  \V190(1) ,
  \V30(27) ,
  \V126(24) ,
  \V94(28) ,
  \V190(0) ,
  \V30(26) ;
output
  \V202(0) ;
wire
  \V206(0) ,
  \V216(0) ,
  \[0] ,
  \V205(0) ,
  \V215(0) ,
  V207,
  V208,
  V209,
  V210,
  V211,
  V212,
  V213,
  V217,
  V218,
  V219,
  V220,
  V221,
  V222,
  V226,
  V227,
  V228,
  V229,
  \V225(0) ,
  V230,
  V231,
  V232,
  V233,
  V234,
  V235,
  V236,
  V237,
  \V204(0) ,
  \V214(0) ,
  \V224(0) ,
  \V203(0) ,
  \V223(0) ;
assign
  \V206(0)  = \V127(0)  | (\V126(30)  | (\V126(28)  | (\V126(26)  | (\V126(24)  | (\V126(22)  | (\V126(20)  | (\V126(18)  | (\V126(16)  | (\V126(14)  | (\V126(12)  | (\V126(10)  | (\V126(8)  | (\V126(6)  | (\V126(4)  | (\V126(2)  | (\V126(3)  | (\V126(5)  | (\V126(7)  | (\V126(9)  | (\V126(11)  | (\V126(13)  | (\V126(15)  | (\V126(17)  | (\V126(19)  | (\V126(21)  | (\V126(23)  | (\V126(25)  | (\V126(27)  | (\V126(29)  | (\V126(31)  | \V128(0) )))))))))))))))))))))))))))))),
  \V216(0)  = \V178(0)  | (\V176(30)  | (\V176(28)  | (\V176(26)  | (\V176(24)  | (\V176(22)  | (\V176(20)  | (\V176(18)  | (\V176(19)  | (\V176(21)  | (\V176(23)  | (\V176(25)  | (\V176(27)  | (\V176(29)  | (\V176(31)  | \V178(1) )))))))))))))),
  \[0]  = V235 | (V236 | (V232 | (V229 | (V230 | (V226 | (V220 | (V221 | (V217 | (V212 | (V210 | (V208 | (V209 | (V211 | (V213 | (V219 | (V218 | (V222 | (V228 | (V227 | (V231 | (V234 | (V233 | V237)))))))))))))))))))))),
  \V205(0)  = \V126(0)  | (\V94(30)  | (\V94(28)  | (\V94(26)  | (\V94(24)  | (\V94(22)  | (\V94(20)  | (\V94(18)  | (\V94(16)  | (\V94(14)  | (\V94(12)  | (\V94(10)  | (\V94(8)  | (\V94(6)  | (\V94(4)  | (\V94(2)  | (\V94(3)  | (\V94(5)  | (\V94(7)  | (\V94(9)  | (\V94(11)  | (\V94(13)  | (\V94(15)  | (\V94(17)  | (\V94(19)  | (\V94(21)  | (\V94(23)  | (\V94(25)  | (\V94(27)  | (\V94(29)  | (\V94(31)  | \V126(1) )))))))))))))))))))))))))))))),
  \V215(0)  = \V176(16)  | (\V176(14)  | (\V176(12)  | (\V176(10)  | (\V176(8)  | (\V176(6)  | (\V176(4)  | (\V176(2)  | (\V176(3)  | (\V176(5)  | (\V176(7)  | (\V176(9)  | (\V176(11)  | (\V176(13)  | (\V176(15)  | \V176(17) )))))))))))))),
  V207 = ~\V201(0) ,
  V208 = \V129(0)  & V207,
  V209 = V207 & (\V203(0)  & \V201(1) ),
  V210 = V207 & (\V204(0)  & \V201(1) ),
  V211 = \V130(0)  & \V201(0) ,
  V212 = \V201(0)  & (\V205(0)  & \V201(1) ),
  V213 = \V201(0)  & (\V206(0)  & \V201(1) ),
  V217 = \V201(2)  & (\V214(0)  & \V201(3) ),
  V218 = \V215(0)  & \V201(2) ,
  V219 = V218 & \V201(3) ,
  V220 = \V216(0)  & \V201(2) ,
  V221 = V220 & \V201(3) ,
  V222 = \V216(0)  & \V201(3) ,
  V226 = \V201(4)  & (\V223(0)  & \V201(5) ),
  V227 = \V224(0)  & \V201(4) ,
  V228 = V227 & \V201(5) ,
  V229 = \V225(0)  & \V201(4) ,
  \V225(0)  = \V190(0)  | (\V188(30)  | (\V188(31)  | \V190(1) )),
  V230 = V229 & \V201(5) ,
  V231 = \V225(0)  & \V201(5) ,
  V232 = \V201(6)  & (\V191(31)  & \V201(7) ),
  V233 = \V193(0)  & \V201(6) ,
  V234 = V233 & \V201(7) ,
  V235 = \V193(1)  & \V201(6) ,
  V236 = V235 & \V201(7) ,
  V237 = \V193(1)  & \V201(7) ,
  \V204(0)  = \V63(0)  | (\V62(30)  | (\V62(28)  | (\V62(26)  | (\V62(24)  | (\V62(22)  | (\V62(20)  | (\V62(18)  | (\V62(16)  | (\V62(14)  | (\V62(12)  | (\V62(10)  | (\V62(8)  | (\V62(6)  | (\V62(4)  | (\V62(2)  | (\V62(3)  | (\V62(5)  | (\V62(7)  | (\V62(9)  | (\V62(11)  | (\V62(13)  | (\V62(15)  | (\V62(17)  | (\V62(19)  | (\V62(21)  | (\V62(23)  | (\V62(25)  | (\V62(27)  | (\V62(29)  | (\V62(31)  | \V64(0) )))))))))))))))))))))))))))))),
  \V214(0)  = \V176(0)  | (\V144(30)  | (\V144(28)  | (\V144(26)  | (\V144(24)  | (\V144(22)  | (\V144(20)  | (\V144(18)  | (\V144(19)  | (\V144(21)  | (\V144(23)  | (\V144(25)  | (\V144(27)  | (\V144(29)  | (\V144(31)  | \V176(1) )))))))))))))),
  \V224(0)  = \V188(28)  | (\V188(26)  | (\V188(27)  | \V188(29) )),
  \V203(0)  = \V62(0)  | (\V30(30)  | (\V30(28)  | (\V30(26)  | (\V30(24)  | (\V30(22)  | (\V30(20)  | (\V30(18)  | (\V30(16)  | (\V30(14)  | (\V30(12)  | (\V30(10)  | (\V30(8)  | (\V30(6)  | (\V30(4)  | (\V30(2)  | (\V30(3)  | (\V30(5)  | (\V30(7)  | (\V30(9)  | (\V30(11)  | (\V30(13)  | (\V30(15)  | (\V30(17)  | (\V30(19)  | (\V30(21)  | (\V30(23)  | (\V30(25)  | (\V30(27)  | (\V30(29)  | (\V30(31)  | \V62(1) )))))))))))))))))))))))))))))),
  \V223(0)  = \V188(24)  | (\V188(22)  | (\V188(23)  | \V188(25) )),
  \V202(0)  = \[0] ;
endmodule

