// IWLS benchmark module "MinMax30" printed on Wed May 29 22:06:08 2002
module MinMax30(\1 , \2 , \3 , \4 , \5 , \6 , \7 , \8 , \9 , \10 , \11 , \12 , \13 , \14 , \15 , \16 , \17 , \18 , \19 , \20 , \21 , \22 , \23 , \24 , \25 , \26 , \27 , \28 , \29 , \30 , \31 , \32 , \33 , \124 , \125 , \126 , \127 , \128 , \129 , \130 , \131 , \132 , \133 , \134 , \135 , \136 , \137 , \138 , \139 , \140 , \141 , \142 , \143 , \144 , \145 , \146 , \147 , \148 , \149 , \150 , \151 , \152 , \153 );
input
  \1 ,
  \2 ,
  \3 ,
  \4 ,
  \5 ,
  \6 ,
  \7 ,
  \8 ,
  \9 ,
  \10 ,
  \11 ,
  \12 ,
  \13 ,
  \14 ,
  \15 ,
  \16 ,
  \17 ,
  \18 ,
  \19 ,
  \20 ,
  \21 ,
  \22 ,
  \23 ,
  \24 ,
  \25 ,
  \26 ,
  \27 ,
  \28 ,
  \29 ,
  \30 ,
  \31 ,
  \32 ,
  \33 ;
output
  \124 ,
  \125 ,
  \126 ,
  \127 ,
  \128 ,
  \129 ,
  \130 ,
  \131 ,
  \132 ,
  \133 ,
  \134 ,
  \135 ,
  \136 ,
  \137 ,
  \138 ,
  \139 ,
  \140 ,
  \141 ,
  \142 ,
  \143 ,
  \144 ,
  \145 ,
  \146 ,
  \147 ,
  \148 ,
  \149 ,
  \150 ,
  \151 ,
  \152 ,
  \153 ;
reg
  \34 ,
  \35 ,
  \36 ,
  \37 ,
  \38 ,
  \39 ,
  \40 ,
  \41 ,
  \42 ,
  \43 ,
  \44 ,
  \45 ,
  \46 ,
  \47 ,
  \48 ,
  \49 ,
  \50 ,
  \51 ,
  \52 ,
  \53 ,
  \54 ,
  \55 ,
  \56 ,
  \57 ,
  \58 ,
  \59 ,
  \60 ,
  \61 ,
  \62 ,
  \63 ,
  \64 ,
  \65 ,
  \66 ,
  \67 ,
  \68 ,
  \69 ,
  \70 ,
  \71 ,
  \72 ,
  \73 ,
  \74 ,
  \75 ,
  \76 ,
  \77 ,
  \78 ,
  \79 ,
  \80 ,
  \81 ,
  \82 ,
  \83 ,
  \84 ,
  \85 ,
  \86 ,
  \87 ,
  \88 ,
  \89 ,
  \90 ,
  \91 ,
  \92 ,
  \93 ,
  \94 ,
  \95 ,
  \96 ,
  \97 ,
  \98 ,
  \99 ,
  \100 ,
  \101 ,
  \102 ,
  \103 ,
  \104 ,
  \105 ,
  \106 ,
  \107 ,
  \108 ,
  \109 ,
  \110 ,
  \111 ,
  \112 ,
  \113 ,
  \114 ,
  \115 ,
  \116 ,
  \117 ,
  \118 ,
  \119 ,
  \120 ,
  \121 ,
  \122 ,
  \123 ;
wire
  \1180 ,
  \1181 ,
  \1182 ,
  \1184 ,
  \1185 ,
  \1186 ,
  \1187 ,
  \1188 ,
  \1189 ,
  \[189] ,
  \1190 ,
  \1192 ,
  \1193 ,
  \1194 ,
  \1195 ,
  \1196 ,
  \1197 ,
  \1198 ,
  \[190] ,
  \1200 ,
  \1201 ,
  \1202 ,
  \1203 ,
  \1204 ,
  \1205 ,
  \1206 ,
  \1208 ,
  \1209 ,
  \[191] ,
  \1210 ,
  \1211 ,
  \1212 ,
  \1213 ,
  \1214 ,
  \1216 ,
  \1217 ,
  \1218 ,
  \1219 ,
  \[192] ,
  \1220 ,
  \1221 ,
  \1222 ,
  \1224 ,
  \1225 ,
  \1226 ,
  \1227 ,
  \1228 ,
  \1229 ,
  \[193] ,
  \1230 ,
  \1232 ,
  \1233 ,
  \1234 ,
  \1235 ,
  \1236 ,
  \1237 ,
  \1238 ,
  \[194] ,
  \1240 ,
  \1241 ,
  \1242 ,
  \1243 ,
  \1244 ,
  \1245 ,
  \1246 ,
  \1248 ,
  \1249 ,
  \[195] ,
  \1250 ,
  \1251 ,
  \1252 ,
  \1253 ,
  \1254 ,
  \1256 ,
  \1257 ,
  \1258 ,
  \1259 ,
  \[196] ,
  \1260 ,
  \1261 ,
  \1262 ,
  \1264 ,
  \1265 ,
  \1266 ,
  \1267 ,
  \1268 ,
  \1269 ,
  \[197] ,
  \1270 ,
  \1272 ,
  \1273 ,
  \1274 ,
  \1275 ,
  \1276 ,
  \1277 ,
  \1278 ,
  \[198] ,
  \1280 ,
  \1281 ,
  \1282 ,
  \1283 ,
  \1284 ,
  \1285 ,
  \1286 ,
  \1288 ,
  \1289 ,
  \[199] ,
  \1290 ,
  \1291 ,
  \1292 ,
  \1293 ,
  \1294 ,
  \1296 ,
  \1297 ,
  \1298 ,
  \1299 ,
  \1300 ,
  \1301 ,
  \1302 ,
  \1304 ,
  \1305 ,
  \1306 ,
  \1307 ,
  \1308 ,
  \1309 ,
  \1310 ,
  \1312 ,
  \1313 ,
  \1314 ,
  \1315 ,
  \1316 ,
  \1317 ,
  \1318 ,
  \1320 ,
  \1321 ,
  \1322 ,
  \1323 ,
  \1324 ,
  \1325 ,
  \1326 ,
  \1328 ,
  \1329 ,
  \1330 ,
  \1331 ,
  \1332 ,
  \1333 ,
  \1334 ,
  \1336 ,
  \1337 ,
  \1338 ,
  \1339 ,
  \1340 ,
  \1341 ,
  \1342 ,
  \1344 ,
  \1345 ,
  \1346 ,
  \1347 ,
  \1348 ,
  \1349 ,
  \1350 ,
  \1352 ,
  \1353 ,
  \1354 ,
  \1355 ,
  \1356 ,
  \1357 ,
  \1358 ,
  \1360 ,
  \1361 ,
  \1362 ,
  \1363 ,
  \1364 ,
  \1365 ,
  \1366 ,
  \1368 ,
  \1371 ,
  \1373 ,
  \1376 ,
  \1378 ,
  \1381 ,
  \1383 ,
  \1386 ,
  \1388 ,
  \1391 ,
  \1393 ,
  \1396 ,
  \1398 ,
  \1401 ,
  \1403 ,
  \1406 ,
  \1408 ,
  \1411 ,
  \1413 ,
  \1416 ,
  \1418 ,
  \1421 ,
  \1423 ,
  \1426 ,
  \1428 ,
  \1431 ,
  \1433 ,
  \1436 ,
  \1438 ,
  \1441 ,
  \1443 ,
  \1446 ,
  \1448 ,
  \1451 ,
  \1453 ,
  \1456 ,
  \1458 ,
  \1461 ,
  \1463 ,
  \1466 ,
  \1468 ,
  \1471 ,
  \1473 ,
  \1476 ,
  \1478 ,
  \1481 ,
  \1483 ,
  \1486 ,
  \1488 ,
  \1491 ,
  \1493 ,
  \1496 ,
  \1498 ,
  \1501 ,
  \1503 ,
  \1506 ,
  \1508 ,
  \1511 ,
  \1513 ,
  \1516 ,
  \1518 ,
  \1520 ,
  \1521 ,
  \1523 ,
  \1524 ,
  \1526 ,
  \1528 ,
  \1529 ,
  \1531 ,
  \1532 ,
  \1534 ,
  \1536 ,
  \1537 ,
  \1539 ,
  \1540 ,
  \1542 ,
  \1544 ,
  \1545 ,
  \1547 ,
  \1548 ,
  \1550 ,
  \1552 ,
  \1553 ,
  \1555 ,
  \1556 ,
  \1558 ,
  \1560 ,
  \1561 ,
  \1563 ,
  \1564 ,
  \1566 ,
  \1568 ,
  \1569 ,
  \1571 ,
  \1572 ,
  \1574 ,
  \1576 ,
  \1577 ,
  \1579 ,
  \1580 ,
  \1582 ,
  \1584 ,
  \1585 ,
  \1587 ,
  \1588 ,
  \1590 ,
  \1592 ,
  \1593 ,
  \1595 ,
  \1596 ,
  \1598 ,
  \1600 ,
  \1601 ,
  \1603 ,
  \1604 ,
  \1606 ,
  \1608 ,
  \1609 ,
  \1611 ,
  \1612 ,
  \1614 ,
  \1616 ,
  \1617 ,
  \1619 ,
  \1620 ,
  \1622 ,
  \1624 ,
  \1625 ,
  \1627 ,
  \1628 ,
  \1630 ,
  \1632 ,
  \1633 ,
  \1635 ,
  \1636 ,
  \1638 ,
  \1640 ,
  \1641 ,
  \1643 ,
  \1644 ,
  \1646 ,
  \1648 ,
  \1649 ,
  \1651 ,
  \1652 ,
  \1654 ,
  \1656 ,
  \1657 ,
  \1659 ,
  \1660 ,
  \1662 ,
  \1664 ,
  \1665 ,
  \1667 ,
  \1668 ,
  \1670 ,
  \1672 ,
  \1673 ,
  \1675 ,
  \1676 ,
  \1678 ,
  \1680 ,
  \1681 ,
  \1683 ,
  \1684 ,
  \1686 ,
  \1688 ,
  \1689 ,
  \1691 ,
  \1692 ,
  \1694 ,
  \1696 ,
  \1697 ,
  \1699 ,
  \1700 ,
  \1702 ,
  \1704 ,
  \1705 ,
  \1707 ,
  \1708 ,
  \1710 ,
  \1712 ,
  \1713 ,
  \1715 ,
  \1716 ,
  \1718 ,
  \1720 ,
  \1721 ,
  \1723 ,
  \1724 ,
  \1726 ,
  \1728 ,
  \1729 ,
  \1731 ,
  \1732 ,
  \1734 ,
  \1736 ,
  \1737 ,
  \1739 ,
  \1740 ,
  \1742 ,
  \1744 ,
  \1745 ,
  \1747 ,
  \1748 ,
  \1750 ,
  \1752 ,
  \1753 ,
  \1755 ,
  \1756 ,
  \1758 ,
  \1761 ,
  \1764 ,
  \1766 ,
  \1769 ,
  \1772 ,
  \1774 ,
  \1777 ,
  \1780 ,
  \1782 ,
  \1785 ,
  \1788 ,
  \1790 ,
  \1793 ,
  \1796 ,
  \1798 ,
  \1801 ,
  \1804 ,
  \1806 ,
  \1809 ,
  \1812 ,
  \1814 ,
  \1817 ,
  \1820 ,
  \1822 ,
  \1825 ,
  \1828 ,
  \1830 ,
  \1833 ,
  \1836 ,
  \1838 ,
  \1841 ,
  \1844 ,
  \1846 ,
  \1849 ,
  \1852 ,
  \1854 ,
  \1857 ,
  \1860 ,
  \1862 ,
  \1865 ,
  \1868 ,
  \1870 ,
  \1873 ,
  \1876 ,
  \1878 ,
  \1881 ,
  \1884 ,
  \1886 ,
  \1889 ,
  \1892 ,
  \1894 ,
  \1897 ,
  \[200] ,
  \1900 ,
  \1902 ,
  \1905 ,
  \1908 ,
  \[201] ,
  \1910 ,
  \1913 ,
  \1916 ,
  \1918 ,
  \[202] ,
  \1921 ,
  \1924 ,
  \1926 ,
  \1929 ,
  \[203] ,
  \1932 ,
  \1934 ,
  \1937 ,
  \[204] ,
  \1940 ,
  \1942 ,
  \1945 ,
  \1948 ,
  \[205] ,
  \1950 ,
  \1953 ,
  \1956 ,
  \1958 ,
  \[206] ,
  \1961 ,
  \1964 ,
  \1966 ,
  \1969 ,
  \[207] ,
  \1972 ,
  \1974 ,
  \1977 ,
  \[208] ,
  \1980 ,
  \1982 ,
  \1985 ,
  \1988 ,
  \[209] ,
  \1990 ,
  \1993 ,
  \1996 ,
  \1998 ,
  \1999 ,
  \2000 ,
  \2001 ,
  \2002 ,
  \2003 ,
  \2004 ,
  \2005 ,
  \2006 ,
  \2007 ,
  \2008 ,
  \2009 ,
  \2010 ,
  \2011 ,
  \2012 ,
  \2013 ,
  \2014 ,
  \2015 ,
  \2016 ,
  \2017 ,
  \2018 ,
  \2019 ,
  \2020 ,
  \2021 ,
  \2022 ,
  \2023 ,
  \2024 ,
  \2025 ,
  \2026 ,
  \2027 ,
  \2028 ,
  \2029 ,
  \2030 ,
  \2031 ,
  \2032 ,
  \2033 ,
  \2034 ,
  \2035 ,
  \2036 ,
  \2037 ,
  \2038 ,
  \2039 ,
  \2040 ,
  \2041 ,
  \2042 ,
  \2043 ,
  \2044 ,
  \2045 ,
  \2046 ,
  \2047 ,
  \2048 ,
  \2049 ,
  \2050 ,
  \2051 ,
  \2052 ,
  \2053 ,
  \2054 ,
  \2055 ,
  \2056 ,
  \2057 ,
  \2058 ,
  \2059 ,
  \2060 ,
  \2061 ,
  \2062 ,
  \2063 ,
  \2064 ,
  \2065 ,
  \2066 ,
  \2067 ,
  \2068 ,
  \2069 ,
  \2070 ,
  \2071 ,
  \2072 ,
  \2073 ,
  \2074 ,
  \2075 ,
  \2076 ,
  \2077 ,
  \2078 ,
  \2079 ,
  \2080 ,
  \2081 ,
  \2082 ,
  \2083 ,
  \2084 ,
  \2085 ,
  \2086 ,
  \2087 ,
  \2088 ,
  \2089 ,
  \2090 ,
  \2091 ,
  \2092 ,
  \2093 ,
  \2094 ,
  \2095 ,
  \2096 ,
  \2097 ,
  \2098 ,
  \2099 ,
  \2100 ,
  \2101 ,
  \2102 ,
  \2103 ,
  \2104 ,
  \2105 ,
  \2106 ,
  \2107 ,
  \2108 ,
  \2109 ,
  \2110 ,
  \2111 ,
  \2112 ,
  \2113 ,
  \2114 ,
  \2115 ,
  \2116 ,
  \2117 ,
  \2118 ,
  \2119 ,
  \2120 ,
  \2121 ,
  \2122 ,
  \2123 ,
  \2124 ,
  \2125 ,
  \2126 ,
  \2127 ,
  \2128 ,
  \2129 ,
  \2130 ,
  \2131 ,
  \2132 ,
  \2133 ,
  \2134 ,
  \2135 ,
  \2136 ,
  \2137 ,
  \2138 ,
  \2139 ,
  \2140 ,
  \2141 ,
  \2142 ,
  \2143 ,
  \2144 ,
  \2145 ,
  \2146 ,
  \2147 ,
  \2148 ,
  \2149 ,
  \2150 ,
  \2151 ,
  \2152 ,
  \2153 ,
  \2154 ,
  \2155 ,
  \2156 ,
  \2157 ,
  \2158 ,
  \2159 ,
  \2160 ,
  \2161 ,
  \2162 ,
  \2163 ,
  \2164 ,
  \2165 ,
  \2166 ,
  \2167 ,
  \2168 ,
  \2169 ,
  \2170 ,
  \2171 ,
  \2172 ,
  \2173 ,
  \2174 ,
  \2175 ,
  \2176 ,
  \2177 ,
  \2178 ,
  \2179 ,
  \2180 ,
  \2181 ,
  \2182 ,
  \2183 ,
  \2184 ,
  \2185 ,
  \2186 ,
  \2187 ,
  \2188 ,
  \2189 ,
  \2190 ,
  \2191 ,
  \2192 ,
  \2193 ,
  \2194 ,
  \2195 ,
  \2196 ,
  \2197 ,
  \2198 ,
  \2199 ,
  \2200 ,
  \2201 ,
  \2202 ,
  \2203 ,
  \2204 ,
  \2205 ,
  \2206 ,
  \2207 ,
  \2208 ,
  \2209 ,
  \2210 ,
  \2211 ,
  \2212 ,
  \2213 ,
  \2214 ,
  \2215 ,
  \2216 ,
  \2217 ,
  \2218 ,
  \2219 ,
  \2220 ,
  \2221 ,
  \2222 ,
  \2223 ,
  \2224 ,
  \2225 ,
  \2226 ,
  \2227 ,
  \2228 ,
  \2229 ,
  \2230 ,
  \2231 ,
  \2232 ,
  \2233 ,
  \2234 ,
  \2235 ,
  \2236 ,
  \2237 ,
  \2238 ,
  \2239 ,
  \2240 ,
  \2241 ,
  \2242 ,
  \2243 ,
  \2244 ,
  \2245 ,
  \2246 ,
  \2247 ,
  \2248 ,
  \2249 ,
  \2250 ,
  \2251 ,
  \2252 ,
  \2253 ,
  \2254 ,
  \2255 ,
  \2256 ,
  \2257 ,
  \2258 ,
  \2259 ,
  \2260 ,
  \2261 ,
  \2262 ,
  \2263 ,
  \2264 ,
  \2265 ,
  \2266 ,
  \2267 ,
  \2268 ,
  \2269 ,
  \2270 ,
  \2271 ,
  \2272 ,
  \2273 ,
  \2274 ,
  \2275 ,
  \2276 ,
  \2277 ,
  \2278 ,
  \2279 ,
  \2280 ,
  \2281 ,
  \2282 ,
  \2283 ,
  \2284 ,
  \2285 ,
  \2286 ,
  \2287 ,
  \2288 ,
  \2289 ,
  \2290 ,
  \2291 ,
  \2292 ,
  \2293 ,
  \2294 ,
  \2295 ,
  \2296 ,
  \2297 ,
  \2299 ,
  \2301 ,
  \2302 ,
  \2303 ,
  \2304 ,
  \2305 ,
  \2306 ,
  \2307 ,
  \2308 ,
  \2309 ,
  \2310 ,
  \2311 ,
  \2312 ,
  \2313 ,
  \2314 ,
  \2315 ,
  \2316 ,
  \2317 ,
  \2318 ,
  \2319 ,
  \2320 ,
  \2321 ,
  \2322 ,
  \2323 ,
  \2324 ,
  \2325 ,
  \2326 ,
  \2327 ,
  \2328 ,
  \2329 ,
  \2330 ,
  \2331 ,
  \2332 ,
  \2333 ,
  \2334 ,
  \2335 ,
  \2336 ,
  \2337 ,
  \2338 ,
  \2339 ,
  \2340 ,
  \2341 ,
  \2342 ,
  \2343 ,
  \2344 ,
  \2345 ,
  \2346 ,
  \2347 ,
  \2348 ,
  \2349 ,
  \2350 ,
  \2351 ,
  \2352 ,
  \2353 ,
  \2354 ,
  \2355 ,
  \2356 ,
  \2357 ,
  \2358 ,
  \2359 ,
  \2360 ,
  \2361 ,
  \2362 ,
  \2363 ,
  \2364 ,
  \2365 ,
  \2366 ,
  \2367 ,
  \2368 ,
  \2369 ,
  \2370 ,
  \2371 ,
  \2372 ,
  \2373 ,
  \2374 ,
  \2375 ,
  \2376 ,
  \2377 ,
  \2378 ,
  \2379 ,
  \2380 ,
  \2381 ,
  \2382 ,
  \2383 ,
  \2384 ,
  \2385 ,
  \2386 ,
  \2387 ,
  \2388 ,
  \2389 ,
  \2391 ,
  \2393 ,
  \2394 ,
  \2395 ,
  \2396 ,
  \2397 ,
  \2398 ,
  \2399 ,
  \2400 ,
  \2401 ,
  \2402 ,
  \2403 ,
  \2404 ,
  \2405 ,
  \2406 ,
  \2407 ,
  \2408 ,
  \2409 ,
  \2410 ,
  \2411 ,
  \2412 ,
  \2413 ,
  \2414 ,
  \2415 ,
  \2416 ,
  \2417 ,
  \2418 ,
  \2419 ,
  \2420 ,
  \2421 ,
  \2422 ,
  \2423 ,
  \2424 ,
  \2425 ,
  \2426 ,
  \2427 ,
  \2428 ,
  \2429 ,
  \2430 ,
  \2431 ,
  \2432 ,
  \2433 ,
  \2434 ,
  \2435 ,
  \2436 ,
  \2437 ,
  \2438 ,
  \2439 ,
  \2440 ,
  \2441 ,
  \2442 ,
  \2443 ,
  \2444 ,
  \2445 ,
  \2446 ,
  \2447 ,
  \2448 ,
  \2449 ,
  \2450 ,
  \2451 ,
  \2452 ,
  \2453 ,
  \2454 ,
  \2455 ,
  \2456 ,
  \2457 ,
  \2458 ,
  \2459 ,
  \2460 ,
  \2461 ,
  \2462 ,
  \2463 ,
  \2464 ,
  \2465 ,
  \2466 ,
  \2467 ,
  \2468 ,
  \2469 ,
  \2470 ,
  \2471 ,
  \2472 ,
  \2473 ,
  \2474 ,
  \2475 ,
  \2476 ,
  \2477 ,
  \2478 ,
  \2479 ,
  \2480 ,
  \2481 ,
  \184 ,
  \185 ,
  \186 ,
  \187 ,
  \188 ,
  \189 ,
  \190 ,
  \191 ,
  \192 ,
  \193 ,
  \194 ,
  \195 ,
  \196 ,
  \197 ,
  \198 ,
  \199 ,
  \200 ,
  \201 ,
  \202 ,
  \203 ,
  \204 ,
  \205 ,
  \206 ,
  \207 ,
  \208 ,
  \209 ,
  \210 ,
  \211 ,
  \212 ,
  \213 ,
  \251 ,
  \253 ,
  \255 ,
  \257 ,
  \259 ,
  \261 ,
  \263 ,
  \265 ,
  \267 ,
  \269 ,
  \271 ,
  \273 ,
  \275 ,
  \277 ,
  \279 ,
  \281 ,
  \283 ,
  \285 ,
  \287 ,
  \289 ,
  \291 ,
  \293 ,
  \295 ,
  \297 ,
  \299 ,
  \301 ,
  \303 ,
  \305 ,
  \307 ,
  \309 ,
  \313 ,
  \315 ,
  \317 ,
  \319 ,
  \321 ,
  \323 ,
  \325 ,
  \327 ,
  \329 ,
  \331 ,
  \333 ,
  \335 ,
  \337 ,
  \339 ,
  \341 ,
  \343 ,
  \345 ,
  \347 ,
  \349 ,
  \351 ,
  \353 ,
  \355 ,
  \357 ,
  \359 ,
  \361 ,
  \363 ,
  \365 ,
  \367 ,
  \369 ,
  \371 ,
  \[120] ,
  \[121] ,
  \[122] ,
  \[123] ,
  \[124] ,
  \[125] ,
  \[126] ,
  \[127] ,
  \[128] ,
  \[129] ,
  \[130] ,
  \[131] ,
  \[132] ,
  \[133] ,
  \[134] ,
  \[135] ,
  \[136] ,
  \[137] ,
  \[138] ,
  \[139] ,
  \[140] ,
  \[141] ,
  \[142] ,
  \[143] ,
  \[144] ,
  \[145] ,
  \[146] ,
  \[147] ,
  \[148] ,
  \[149] ,
  \[150] ,
  \[151] ,
  \[152] ,
  \[153] ,
  \[154] ,
  \[155] ,
  \[156] ,
  \[157] ,
  \[158] ,
  \[159] ,
  \[160] ,
  \[161] ,
  \[162] ,
  \[163] ,
  \[164] ,
  \[165] ,
  \[166] ,
  \[167] ,
  \[168] ,
  \[169] ,
  \916 ,
  \917 ,
  \918 ,
  \919 ,
  \920 ,
  \921 ,
  \922 ,
  \923 ,
  \924 ,
  \925 ,
  \926 ,
  \927 ,
  \928 ,
  \929 ,
  \930 ,
  \931 ,
  \932 ,
  \933 ,
  \934 ,
  \935 ,
  \936 ,
  \937 ,
  \938 ,
  \939 ,
  \940 ,
  \941 ,
  \942 ,
  \943 ,
  \944 ,
  \945 ,
  \[170] ,
  \[171] ,
  \[172] ,
  \[173] ,
  \1036 ,
  \1037 ,
  \1039 ,
  \[174] ,
  \1040 ,
  \1041 ,
  \1042 ,
  \1043 ,
  \1044 ,
  \1045 ,
  \1046 ,
  \1047 ,
  \1048 ,
  \1049 ,
  \[175] ,
  \1050 ,
  \1051 ,
  \1052 ,
  \1053 ,
  \1054 ,
  \1055 ,
  \1056 ,
  \1057 ,
  \1058 ,
  \1059 ,
  \[176] ,
  \1060 ,
  \1061 ,
  \1062 ,
  \1063 ,
  \1064 ,
  \1065 ,
  \1066 ,
  \1067 ,
  \1068 ,
  \1069 ,
  \[177] ,
  \1070 ,
  \1071 ,
  \1072 ,
  \1073 ,
  \1074 ,
  \1075 ,
  \1076 ,
  \1077 ,
  \1078 ,
  \1079 ,
  \[178] ,
  \1080 ,
  \1081 ,
  \1082 ,
  \1083 ,
  \1084 ,
  \1085 ,
  \1086 ,
  \1087 ,
  \1088 ,
  \1089 ,
  \[179] ,
  \1090 ,
  \1091 ,
  \1092 ,
  \1093 ,
  \1094 ,
  \1095 ,
  \1096 ,
  \1097 ,
  \1098 ,
  \1099 ,
  \[180] ,
  \1100 ,
  \1101 ,
  \1102 ,
  \1103 ,
  \1104 ,
  \1105 ,
  \1106 ,
  \1107 ,
  \1108 ,
  \1109 ,
  \[181] ,
  \1110 ,
  \1111 ,
  \1112 ,
  \1113 ,
  \1114 ,
  \1115 ,
  \1116 ,
  \1117 ,
  \1118 ,
  \1119 ,
  \[182] ,
  \1120 ,
  \1121 ,
  \1122 ,
  \1123 ,
  \1124 ,
  \1125 ,
  \1126 ,
  \1127 ,
  \1128 ,
  \1129 ,
  \[183] ,
  \1130 ,
  \1131 ,
  \1132 ,
  \1133 ,
  \1134 ,
  \1136 ,
  \1137 ,
  \1138 ,
  \1139 ,
  \[184] ,
  \1140 ,
  \1141 ,
  \1142 ,
  \1144 ,
  \1145 ,
  \1146 ,
  \1147 ,
  \1148 ,
  \1149 ,
  \[185] ,
  \1150 ,
  \1152 ,
  \1153 ,
  \1154 ,
  \1155 ,
  \1156 ,
  \1157 ,
  \1158 ,
  \[186] ,
  \1160 ,
  \1161 ,
  \1162 ,
  \1163 ,
  \1164 ,
  \1165 ,
  \1166 ,
  \1168 ,
  \1169 ,
  \[187] ,
  \1170 ,
  \1171 ,
  \1172 ,
  \1173 ,
  \1174 ,
  \1176 ,
  \1177 ,
  \1178 ,
  \1179 ,
  \[188] ;
assign
  \1180  = \40  & ~\2 ,
  \1181  = \1180  | \1179 ,
  \1182  = \1181  & ~\1 ,
  \1184  = \924  & ~\3 ,
  \1185  = \11  & \3 ,
  \1186  = \1185  | \1184 ,
  \1187  = \1186  & \2 ,
  \1188  = \41  & ~\2 ,
  \1189  = \1188  | \1187 ,
  \[189]  = \1836 ,
  \1190  = \1189  & ~\1 ,
  \1192  = \925  & ~\3 ,
  \1193  = \12  & \3 ,
  \1194  = \1193  | \1192 ,
  \1195  = \1194  & \2 ,
  \1196  = \42  & ~\2 ,
  \1197  = \1196  | \1195 ,
  \1198  = \1197  & ~\1 ,
  \[190]  = \1844 ,
  \1200  = \926  & ~\3 ,
  \1201  = \13  & \3 ,
  \1202  = \1201  | \1200 ,
  \1203  = \1202  & \2 ,
  \1204  = \43  & ~\2 ,
  \1205  = \1204  | \1203 ,
  \1206  = \1205  & ~\1 ,
  \1208  = \927  & ~\3 ,
  \1209  = \14  & \3 ,
  \[191]  = \1852 ,
  \1210  = \1209  | \1208 ,
  \1211  = \1210  & \2 ,
  \1212  = \44  & ~\2 ,
  \1213  = \1212  | \1211 ,
  \1214  = \1213  & ~\1 ,
  \1216  = \928  & ~\3 ,
  \1217  = \15  & \3 ,
  \1218  = \1217  | \1216 ,
  \1219  = \1218  & \2 ,
  \[192]  = \1860 ,
  \1220  = \45  & ~\2 ,
  \1221  = \1220  | \1219 ,
  \1222  = \1221  & ~\1 ,
  \1224  = \929  & ~\3 ,
  \1225  = \16  & \3 ,
  \1226  = \1225  | \1224 ,
  \1227  = \1226  & \2 ,
  \1228  = \46  & ~\2 ,
  \1229  = \1228  | \1227 ,
  \[193]  = \1868 ,
  \1230  = \1229  & ~\1 ,
  \1232  = \930  & ~\3 ,
  \1233  = \17  & \3 ,
  \1234  = \1233  | \1232 ,
  \1235  = \1234  & \2 ,
  \1236  = \47  & ~\2 ,
  \1237  = \1236  | \1235 ,
  \1238  = \1237  & ~\1 ,
  \[194]  = \1876 ,
  \1240  = \931  & ~\3 ,
  \1241  = \18  & \3 ,
  \1242  = \1241  | \1240 ,
  \1243  = \1242  & \2 ,
  \1244  = \48  & ~\2 ,
  \1245  = \1244  | \1243 ,
  \1246  = \1245  & ~\1 ,
  \1248  = \932  & ~\3 ,
  \1249  = \19  & \3 ,
  \[195]  = \1884 ,
  \1250  = \1249  | \1248 ,
  \1251  = \1250  & \2 ,
  \1252  = \49  & ~\2 ,
  \1253  = \1252  | \1251 ,
  \1254  = \1253  & ~\1 ,
  \1256  = \933  & ~\3 ,
  \1257  = \20  & \3 ,
  \1258  = \1257  | \1256 ,
  \1259  = \1258  & \2 ,
  \[196]  = \1892 ,
  \1260  = \50  & ~\2 ,
  \1261  = \1260  | \1259 ,
  \1262  = \1261  & ~\1 ,
  \1264  = \934  & ~\3 ,
  \1265  = \21  & \3 ,
  \1266  = \1265  | \1264 ,
  \1267  = \1266  & \2 ,
  \1268  = \51  & ~\2 ,
  \1269  = \1268  | \1267 ,
  \[197]  = \1900 ,
  \1270  = \1269  & ~\1 ,
  \1272  = \935  & ~\3 ,
  \1273  = \22  & \3 ,
  \1274  = \1273  | \1272 ,
  \1275  = \1274  & \2 ,
  \1276  = \52  & ~\2 ,
  \1277  = \1276  | \1275 ,
  \1278  = \1277  & ~\1 ,
  \[198]  = \1908 ,
  \1280  = \936  & ~\3 ,
  \1281  = \23  & \3 ,
  \1282  = \1281  | \1280 ,
  \1283  = \1282  & \2 ,
  \1284  = \53  & ~\2 ,
  \1285  = \1284  | \1283 ,
  \1286  = \1285  & ~\1 ,
  \1288  = \937  & ~\3 ,
  \1289  = \24  & \3 ,
  \[199]  = \1916 ,
  \1290  = \1289  | \1288 ,
  \1291  = \1290  & \2 ,
  \1292  = \54  & ~\2 ,
  \1293  = \1292  | \1291 ,
  \1294  = \1293  & ~\1 ,
  \1296  = \938  & ~\3 ,
  \1297  = \25  & \3 ,
  \1298  = \1297  | \1296 ,
  \1299  = \1298  & \2 ,
  \1300  = \55  & ~\2 ,
  \1301  = \1300  | \1299 ,
  \1302  = \1301  & ~\1 ,
  \1304  = \939  & ~\3 ,
  \1305  = \26  & \3 ,
  \1306  = \1305  | \1304 ,
  \1307  = \1306  & \2 ,
  \1308  = \56  & ~\2 ,
  \1309  = \1308  | \1307 ,
  \1310  = \1309  & ~\1 ,
  \1312  = \940  & ~\3 ,
  \1313  = \27  & \3 ,
  \1314  = \1313  | \1312 ,
  \1315  = \1314  & \2 ,
  \1316  = \57  & ~\2 ,
  \1317  = \1316  | \1315 ,
  \1318  = \1317  & ~\1 ,
  \1320  = \941  & ~\3 ,
  \1321  = \28  & \3 ,
  \1322  = \1321  | \1320 ,
  \1323  = \1322  & \2 ,
  \1324  = \58  & ~\2 ,
  \1325  = \1324  | \1323 ,
  \1326  = \1325  & ~\1 ,
  \1328  = \942  & ~\3 ,
  \1329  = \29  & \3 ,
  \1330  = \1329  | \1328 ,
  \1331  = \1330  & \2 ,
  \1332  = \59  & ~\2 ,
  \1333  = \1332  | \1331 ,
  \1334  = \1333  & ~\1 ,
  \1336  = \943  & ~\3 ,
  \1337  = \30  & \3 ,
  \1338  = \1337  | \1336 ,
  \1339  = \1338  & \2 ,
  \1340  = \60  & ~\2 ,
  \1341  = \1340  | \1339 ,
  \1342  = \1341  & ~\1 ,
  \1344  = \944  & ~\3 ,
  \1345  = \31  & \3 ,
  \1346  = \1345  | \1344 ,
  \1347  = \1346  & \2 ,
  \1348  = \61  & ~\2 ,
  \1349  = \1348  | \1347 ,
  \1350  = \1349  & ~\1 ,
  \1352  = \945  & ~\3 ,
  \1353  = \32  & \3 ,
  \1354  = \1353  | \1352 ,
  \1355  = \1354  & \2 ,
  \1356  = \62  & ~\2 ,
  \1357  = \1356  | \1355 ,
  \1358  = \1357  & ~\1 ,
  \1360  = \916  & ~\3 ,
  \1361  = \33  & \3 ,
  \1362  = \1361  | \1360 ,
  \1363  = \1362  & \2 ,
  \1364  = \63  & ~\2 ,
  \1365  = \1364  | \1363 ,
  \1366  = \1365  & ~\1 ,
  \1368  = \4  & \2 ,
  \1371  = \1368  & ~\1 ,
  \1373  = \5  & \2 ,
  \1376  = \1373  & ~\1 ,
  \1378  = \6  & \2 ,
  \1381  = \1378  & ~\1 ,
  \1383  = \7  & \2 ,
  \1386  = \1383  & ~\1 ,
  \1388  = \8  & \2 ,
  \1391  = \1388  & ~\1 ,
  \1393  = \9  & \2 ,
  \1396  = \1393  & ~\1 ,
  \1398  = \10  & \2 ,
  \1401  = \1398  & ~\1 ,
  \1403  = \11  & \2 ,
  \1406  = \1403  & ~\1 ,
  \1408  = \12  & \2 ,
  \1411  = \1408  & ~\1 ,
  \1413  = \13  & \2 ,
  \1416  = \1413  & ~\1 ,
  \1418  = \14  & \2 ,
  \1421  = \1418  & ~\1 ,
  \1423  = \15  & \2 ,
  \1426  = \1423  & ~\1 ,
  \1428  = \16  & \2 ,
  \1431  = \1428  & ~\1 ,
  \1433  = \17  & \2 ,
  \1436  = \1433  & ~\1 ,
  \1438  = \18  & \2 ,
  \1441  = \1438  & ~\1 ,
  \1443  = \19  & \2 ,
  \1446  = \1443  & ~\1 ,
  \1448  = \20  & \2 ,
  \1451  = \1448  & ~\1 ,
  \1453  = \21  & \2 ,
  \1456  = \1453  & ~\1 ,
  \1458  = \22  & \2 ,
  \1461  = \1458  & ~\1 ,
  \1463  = \23  & \2 ,
  \1466  = \1463  & ~\1 ,
  \1468  = \24  & \2 ,
  \1471  = \1468  & ~\1 ,
  \1473  = \25  & \2 ,
  \1476  = \1473  & ~\1 ,
  \1478  = \26  & \2 ,
  \1481  = \1478  & ~\1 ,
  \1483  = \27  & \2 ,
  \1486  = \1483  & ~\1 ,
  \1488  = \28  & \2 ,
  \1491  = \1488  & ~\1 ,
  \1493  = \29  & \2 ,
  \1496  = \1493  & ~\1 ,
  \1498  = \30  & \2 ,
  \1501  = \1498  & ~\1 ,
  \1503  = \31  & \2 ,
  \1506  = \1503  & ~\1 ,
  \1508  = \32  & \2 ,
  \1511  = \1508  & ~\1 ,
  \1513  = \33  & \2 ,
  \1516  = \1513  & ~\1 ,
  \1518  = \1040  & ~\3 ,
  \1520  = \1518  | \3 ,
  \1521  = \1520  & \2 ,
  \1523  = \1521  | ~\2 ,
  \1524  = \1523  & ~\1 ,
  \1526  = \1043  & ~\3 ,
  \1528  = \1526  | \3 ,
  \1529  = \1528  & \2 ,
  \1531  = \1529  | ~\2 ,
  \1532  = \1531  & ~\1 ,
  \1534  = \1046  & ~\3 ,
  \1536  = \1534  | \3 ,
  \1537  = \1536  & \2 ,
  \1539  = \1537  | ~\2 ,
  \1540  = \1539  & ~\1 ,
  \1542  = \1049  & ~\3 ,
  \1544  = \1542  | \3 ,
  \1545  = \1544  & \2 ,
  \1547  = \1545  | ~\2 ,
  \1548  = \1547  & ~\1 ,
  \1550  = \1052  & ~\3 ,
  \1552  = \1550  | \3 ,
  \1553  = \1552  & \2 ,
  \1555  = \1553  | ~\2 ,
  \1556  = \1555  & ~\1 ,
  \1558  = \1055  & ~\3 ,
  \1560  = \1558  | \3 ,
  \1561  = \1560  & \2 ,
  \1563  = \1561  | ~\2 ,
  \1564  = \1563  & ~\1 ,
  \1566  = \1058  & ~\3 ,
  \1568  = \1566  | \3 ,
  \1569  = \1568  & \2 ,
  \1571  = \1569  | ~\2 ,
  \1572  = \1571  & ~\1 ,
  \1574  = \1061  & ~\3 ,
  \1576  = \1574  | \3 ,
  \1577  = \1576  & \2 ,
  \1579  = \1577  | ~\2 ,
  \1580  = \1579  & ~\1 ,
  \1582  = \1064  & ~\3 ,
  \1584  = \1582  | \3 ,
  \1585  = \1584  & \2 ,
  \1587  = \1585  | ~\2 ,
  \1588  = \1587  & ~\1 ,
  \1590  = \1067  & ~\3 ,
  \1592  = \1590  | \3 ,
  \1593  = \1592  & \2 ,
  \1595  = \1593  | ~\2 ,
  \1596  = \1595  & ~\1 ,
  \1598  = \1070  & ~\3 ,
  \1600  = \1598  | \3 ,
  \1601  = \1600  & \2 ,
  \1603  = \1601  | ~\2 ,
  \1604  = \1603  & ~\1 ,
  \1606  = \1073  & ~\3 ,
  \1608  = \1606  | \3 ,
  \1609  = \1608  & \2 ,
  \1611  = \1609  | ~\2 ,
  \1612  = \1611  & ~\1 ,
  \1614  = \1076  & ~\3 ,
  \1616  = \1614  | \3 ,
  \1617  = \1616  & \2 ,
  \1619  = \1617  | ~\2 ,
  \1620  = \1619  & ~\1 ,
  \1622  = \1079  & ~\3 ,
  \1624  = \1622  | \3 ,
  \1625  = \1624  & \2 ,
  \1627  = \1625  | ~\2 ,
  \1628  = \1627  & ~\1 ,
  \1630  = \1082  & ~\3 ,
  \1632  = \1630  | \3 ,
  \1633  = \1632  & \2 ,
  \1635  = \1633  | ~\2 ,
  \1636  = \1635  & ~\1 ,
  \1638  = \1085  & ~\3 ,
  \1640  = \1638  | \3 ,
  \1641  = \1640  & \2 ,
  \1643  = \1641  | ~\2 ,
  \1644  = \1643  & ~\1 ,
  \1646  = \1088  & ~\3 ,
  \1648  = \1646  | \3 ,
  \1649  = \1648  & \2 ,
  \1651  = \1649  | ~\2 ,
  \1652  = \1651  & ~\1 ,
  \1654  = \1091  & ~\3 ,
  \1656  = \1654  | \3 ,
  \1657  = \1656  & \2 ,
  \1659  = \1657  | ~\2 ,
  \1660  = \1659  & ~\1 ,
  \1662  = \1094  & ~\3 ,
  \1664  = \1662  | \3 ,
  \1665  = \1664  & \2 ,
  \1667  = \1665  | ~\2 ,
  \1668  = \1667  & ~\1 ,
  \1670  = \1097  & ~\3 ,
  \1672  = \1670  | \3 ,
  \1673  = \1672  & \2 ,
  \1675  = \1673  | ~\2 ,
  \1676  = \1675  & ~\1 ,
  \1678  = \1100  & ~\3 ,
  \1680  = \1678  | \3 ,
  \1681  = \1680  & \2 ,
  \1683  = \1681  | ~\2 ,
  \1684  = \1683  & ~\1 ,
  \1686  = \1103  & ~\3 ,
  \1688  = \1686  | \3 ,
  \1689  = \1688  & \2 ,
  \1691  = \1689  | ~\2 ,
  \1692  = \1691  & ~\1 ,
  \1694  = \1106  & ~\3 ,
  \1696  = \1694  | \3 ,
  \1697  = \1696  & \2 ,
  \1699  = \1697  | ~\2 ,
  \1700  = \1699  & ~\1 ,
  \1702  = \1109  & ~\3 ,
  \1704  = \1702  | \3 ,
  \1705  = \1704  & \2 ,
  \1707  = \1705  | ~\2 ,
  \1708  = \1707  & ~\1 ,
  \1710  = \1112  & ~\3 ,
  \1712  = \1710  | \3 ,
  \1713  = \1712  & \2 ,
  \1715  = \1713  | ~\2 ,
  \1716  = \1715  & ~\1 ,
  \1718  = \1115  & ~\3 ,
  \1720  = \1718  | \3 ,
  \1721  = \1720  & \2 ,
  \1723  = \1721  | ~\2 ,
  \1724  = \1723  & ~\1 ,
  \1726  = \1118  & ~\3 ,
  \1728  = \1726  | \3 ,
  \1729  = \1728  & \2 ,
  \1731  = \1729  | ~\2 ,
  \1732  = \1731  & ~\1 ,
  \1734  = \1121  & ~\3 ,
  \1736  = \1734  | \3 ,
  \1737  = \1736  & \2 ,
  \1739  = \1737  | ~\2 ,
  \1740  = \1739  & ~\1 ,
  \1742  = \1124  & ~\3 ,
  \1744  = \1742  | \3 ,
  \1745  = \1744  & \2 ,
  \1747  = \1745  | ~\2 ,
  \1748  = \1747  & ~\1 ,
  \1750  = \1127  & ~\3 ,
  \1752  = \1750  | \3 ,
  \1753  = \1752  & \2 ,
  \1755  = \1753  | ~\2 ,
  \1756  = \1755  & ~\1 ,
  \1758  = \1039  & ~\3 ,
  \1761  = \1758  & \2 ,
  \1764  = \1761  & ~\1 ,
  \1766  = \1042  & ~\3 ,
  \1769  = \1766  & \2 ,
  \1772  = \1769  & ~\1 ,
  \1774  = \1045  & ~\3 ,
  \1777  = \1774  & \2 ,
  \1780  = \1777  & ~\1 ,
  \1782  = \1048  & ~\3 ,
  \1785  = \1782  & \2 ,
  \1788  = \1785  & ~\1 ,
  \1790  = \1051  & ~\3 ,
  \1793  = \1790  & \2 ,
  \1796  = \1793  & ~\1 ,
  \1798  = \1054  & ~\3 ,
  \1801  = \1798  & \2 ,
  \1804  = \1801  & ~\1 ,
  \1806  = \1057  & ~\3 ,
  \1809  = \1806  & \2 ,
  \1812  = \1809  & ~\1 ,
  \1814  = \1060  & ~\3 ,
  \1817  = \1814  & \2 ,
  \1820  = \1817  & ~\1 ,
  \1822  = \1063  & ~\3 ,
  \1825  = \1822  & \2 ,
  \1828  = \1825  & ~\1 ,
  \1830  = \1066  & ~\3 ,
  \1833  = \1830  & \2 ,
  \1836  = \1833  & ~\1 ,
  \1838  = \1069  & ~\3 ,
  \1841  = \1838  & \2 ,
  \1844  = \1841  & ~\1 ,
  \1846  = \1072  & ~\3 ,
  \1849  = \1846  & \2 ,
  \1852  = \1849  & ~\1 ,
  \1854  = \1075  & ~\3 ,
  \1857  = \1854  & \2 ,
  \1860  = \1857  & ~\1 ,
  \1862  = \1078  & ~\3 ,
  \1865  = \1862  & \2 ,
  \1868  = \1865  & ~\1 ,
  \1870  = \1081  & ~\3 ,
  \1873  = \1870  & \2 ,
  \1876  = \1873  & ~\1 ,
  \1878  = \1084  & ~\3 ,
  \1881  = \1878  & \2 ,
  \1884  = \1881  & ~\1 ,
  \1886  = \1087  & ~\3 ,
  \1889  = \1886  & \2 ,
  \1892  = \1889  & ~\1 ,
  \1894  = \1090  & ~\3 ,
  \1897  = \1894  & \2 ,
  \[200]  = \1924 ,
  \1900  = \1897  & ~\1 ,
  \1902  = \1093  & ~\3 ,
  \1905  = \1902  & \2 ,
  \1908  = \1905  & ~\1 ,
  \[201]  = \1932 ,
  \1910  = \1096  & ~\3 ,
  \1913  = \1910  & \2 ,
  \1916  = \1913  & ~\1 ,
  \1918  = \1099  & ~\3 ,
  \[202]  = \1940 ,
  \1921  = \1918  & \2 ,
  \1924  = \1921  & ~\1 ,
  \1926  = \1102  & ~\3 ,
  \1929  = \1926  & \2 ,
  \[203]  = \1948 ,
  \1932  = \1929  & ~\1 ,
  \1934  = \1105  & ~\3 ,
  \1937  = \1934  & \2 ,
  \[204]  = \1956 ,
  \1940  = \1937  & ~\1 ,
  \1942  = \1108  & ~\3 ,
  \1945  = \1942  & \2 ,
  \1948  = \1945  & ~\1 ,
  \[205]  = \1964 ,
  \1950  = \1111  & ~\3 ,
  \1953  = \1950  & \2 ,
  \1956  = \1953  & ~\1 ,
  \1958  = \1114  & ~\3 ,
  \[206]  = \1972 ,
  \1961  = \1958  & \2 ,
  \1964  = \1961  & ~\1 ,
  \1966  = \1117  & ~\3 ,
  \1969  = \1966  & \2 ,
  \[207]  = \1980 ,
  \1972  = \1969  & ~\1 ,
  \1974  = \1120  & ~\3 ,
  \1977  = \1974  & \2 ,
  \[208]  = \1988 ,
  \1980  = \1977  & ~\1 ,
  \1982  = \1123  & ~\3 ,
  \1985  = \1982  & \2 ,
  \1988  = \1985  & ~\1 ,
  \[209]  = \1996 ,
  \1990  = \1126  & ~\3 ,
  \1993  = \1990  & \2 ,
  \1996  = \1993  & ~\1 ,
  \1998  = \1037  & \93 ,
  \1999  = ~\1037  & \33 ,
  \2000  = \1999  | \1998 ,
  \2001  = ~\3  & \2 ,
  \2002  = \2001  & ~\1 ,
  \2003  = ~\1036  & \123 ,
  \2004  = \1036  & \33 ,
  \2005  = \2004  | \2003 ,
  \2006  = ~\3  & \2 ,
  \2007  = \2006  & ~\1 ,
  \2008  = \1037  & \92 ,
  \2009  = ~\1037  & \32 ,
  \2010  = \2009  | \2008 ,
  \2011  = ~\3  & \2 ,
  \2012  = \2011  & ~\1 ,
  \2013  = ~\1036  & \122 ,
  \2014  = \1036  & \32 ,
  \2015  = \2014  | \2013 ,
  \2016  = ~\3  & \2 ,
  \2017  = \2016  & ~\1 ,
  \2018  = \1037  & \91 ,
  \2019  = ~\1037  & \31 ,
  \2020  = \2019  | \2018 ,
  \2021  = ~\3  & \2 ,
  \2022  = \2021  & ~\1 ,
  \2023  = ~\1036  & \121 ,
  \2024  = \1036  & \31 ,
  \2025  = \2024  | \2023 ,
  \2026  = ~\3  & \2 ,
  \2027  = \2026  & ~\1 ,
  \2028  = \1037  & \90 ,
  \2029  = ~\1037  & \30 ,
  \2030  = \2029  | \2028 ,
  \2031  = ~\3  & \2 ,
  \2032  = \2031  & ~\1 ,
  \2033  = ~\1036  & \120 ,
  \2034  = \1036  & \30 ,
  \2035  = \2034  | \2033 ,
  \2036  = ~\3  & \2 ,
  \2037  = \2036  & ~\1 ,
  \2038  = \1037  & \89 ,
  \2039  = ~\1037  & \29 ,
  \2040  = \2039  | \2038 ,
  \2041  = ~\3  & \2 ,
  \2042  = \2041  & ~\1 ,
  \2043  = ~\1036  & \119 ,
  \2044  = \1036  & \29 ,
  \2045  = \2044  | \2043 ,
  \2046  = ~\3  & \2 ,
  \2047  = \2046  & ~\1 ,
  \2048  = \1037  & \88 ,
  \2049  = ~\1037  & \28 ,
  \2050  = \2049  | \2048 ,
  \2051  = ~\3  & \2 ,
  \2052  = \2051  & ~\1 ,
  \2053  = ~\1036  & \118 ,
  \2054  = \1036  & \28 ,
  \2055  = \2054  | \2053 ,
  \2056  = ~\3  & \2 ,
  \2057  = \2056  & ~\1 ,
  \2058  = \1037  & \87 ,
  \2059  = ~\1037  & \27 ,
  \2060  = \2059  | \2058 ,
  \2061  = ~\3  & \2 ,
  \2062  = \2061  & ~\1 ,
  \2063  = ~\1036  & \117 ,
  \2064  = \1036  & \27 ,
  \2065  = \2064  | \2063 ,
  \2066  = ~\3  & \2 ,
  \2067  = \2066  & ~\1 ,
  \2068  = \1037  & \86 ,
  \2069  = ~\1037  & \26 ,
  \2070  = \2069  | \2068 ,
  \2071  = ~\3  & \2 ,
  \2072  = \2071  & ~\1 ,
  \2073  = ~\1036  & \116 ,
  \2074  = \1036  & \26 ,
  \2075  = \2074  | \2073 ,
  \2076  = ~\3  & \2 ,
  \2077  = \2076  & ~\1 ,
  \2078  = \1037  & \85 ,
  \2079  = ~\1037  & \25 ,
  \2080  = \2079  | \2078 ,
  \2081  = ~\3  & \2 ,
  \2082  = \2081  & ~\1 ,
  \2083  = ~\1036  & \115 ,
  \2084  = \1036  & \25 ,
  \2085  = \2084  | \2083 ,
  \2086  = ~\3  & \2 ,
  \2087  = \2086  & ~\1 ,
  \2088  = \1037  & \84 ,
  \2089  = ~\1037  & \24 ,
  \2090  = \2089  | \2088 ,
  \2091  = ~\3  & \2 ,
  \2092  = \2091  & ~\1 ,
  \2093  = ~\1036  & \114 ,
  \2094  = \1036  & \24 ,
  \2095  = \2094  | \2093 ,
  \2096  = ~\3  & \2 ,
  \2097  = \2096  & ~\1 ,
  \2098  = \1037  & \83 ,
  \2099  = ~\1037  & \23 ,
  \2100  = \2099  | \2098 ,
  \2101  = ~\3  & \2 ,
  \2102  = \2101  & ~\1 ,
  \2103  = ~\1036  & \113 ,
  \2104  = \1036  & \23 ,
  \2105  = \2104  | \2103 ,
  \2106  = ~\3  & \2 ,
  \2107  = \2106  & ~\1 ,
  \2108  = \1037  & \82 ,
  \2109  = ~\1037  & \22 ,
  \2110  = \2109  | \2108 ,
  \2111  = ~\3  & \2 ,
  \2112  = \2111  & ~\1 ,
  \2113  = ~\1036  & \112 ,
  \2114  = \1036  & \22 ,
  \2115  = \2114  | \2113 ,
  \2116  = ~\3  & \2 ,
  \2117  = \2116  & ~\1 ,
  \2118  = \1037  & \81 ,
  \2119  = ~\1037  & \21 ,
  \2120  = \2119  | \2118 ,
  \2121  = ~\3  & \2 ,
  \2122  = \2121  & ~\1 ,
  \2123  = ~\1036  & \111 ,
  \2124  = \1036  & \21 ,
  \2125  = \2124  | \2123 ,
  \2126  = ~\3  & \2 ,
  \2127  = \2126  & ~\1 ,
  \2128  = \1037  & \80 ,
  \2129  = ~\1037  & \20 ,
  \2130  = \2129  | \2128 ,
  \2131  = ~\3  & \2 ,
  \2132  = \2131  & ~\1 ,
  \2133  = ~\1036  & \110 ,
  \2134  = \1036  & \20 ,
  \2135  = \2134  | \2133 ,
  \2136  = ~\3  & \2 ,
  \2137  = \2136  & ~\1 ,
  \2138  = \1037  & \79 ,
  \2139  = ~\1037  & \19 ,
  \2140  = \2139  | \2138 ,
  \2141  = ~\3  & \2 ,
  \2142  = \2141  & ~\1 ,
  \2143  = ~\1036  & \109 ,
  \2144  = \1036  & \19 ,
  \2145  = \2144  | \2143 ,
  \2146  = ~\3  & \2 ,
  \2147  = \2146  & ~\1 ,
  \2148  = \1037  & \78 ,
  \2149  = ~\1037  & \18 ,
  \2150  = \2149  | \2148 ,
  \2151  = ~\3  & \2 ,
  \2152  = \2151  & ~\1 ,
  \2153  = ~\1036  & \108 ,
  \2154  = \1036  & \18 ,
  \2155  = \2154  | \2153 ,
  \2156  = ~\3  & \2 ,
  \2157  = \2156  & ~\1 ,
  \2158  = \1037  & \77 ,
  \2159  = ~\1037  & \17 ,
  \2160  = \2159  | \2158 ,
  \2161  = ~\3  & \2 ,
  \2162  = \2161  & ~\1 ,
  \2163  = ~\1036  & \107 ,
  \2164  = \1036  & \17 ,
  \2165  = \2164  | \2163 ,
  \2166  = ~\3  & \2 ,
  \2167  = \2166  & ~\1 ,
  \2168  = \1037  & \76 ,
  \2169  = ~\1037  & \16 ,
  \2170  = \2169  | \2168 ,
  \2171  = ~\3  & \2 ,
  \2172  = \2171  & ~\1 ,
  \2173  = ~\1036  & \106 ,
  \2174  = \1036  & \16 ,
  \2175  = \2174  | \2173 ,
  \2176  = ~\3  & \2 ,
  \2177  = \2176  & ~\1 ,
  \2178  = \1037  & \75 ,
  \2179  = ~\1037  & \15 ,
  \2180  = \2179  | \2178 ,
  \2181  = ~\3  & \2 ,
  \2182  = \2181  & ~\1 ,
  \2183  = ~\1036  & \105 ,
  \2184  = \1036  & \15 ,
  \2185  = \2184  | \2183 ,
  \2186  = ~\3  & \2 ,
  \2187  = \2186  & ~\1 ,
  \2188  = \1037  & \74 ,
  \2189  = ~\1037  & \14 ,
  \2190  = \2189  | \2188 ,
  \2191  = ~\3  & \2 ,
  \2192  = \2191  & ~\1 ,
  \2193  = ~\1036  & \104 ,
  \2194  = \1036  & \14 ,
  \2195  = \2194  | \2193 ,
  \2196  = ~\3  & \2 ,
  \2197  = \2196  & ~\1 ,
  \2198  = \1037  & \73 ,
  \2199  = ~\1037  & \13 ,
  \2200  = \2199  | \2198 ,
  \2201  = ~\3  & \2 ,
  \2202  = \2201  & ~\1 ,
  \2203  = ~\1036  & \103 ,
  \2204  = \1036  & \13 ,
  \2205  = \2204  | \2203 ,
  \2206  = ~\3  & \2 ,
  \2207  = \2206  & ~\1 ,
  \2208  = \1037  & \72 ,
  \2209  = ~\1037  & \12 ,
  \2210  = \2209  | \2208 ,
  \2211  = ~\3  & \2 ,
  \2212  = \2211  & ~\1 ,
  \2213  = ~\1036  & \102 ,
  \2214  = \1036  & \12 ,
  \2215  = \2214  | \2213 ,
  \2216  = ~\3  & \2 ,
  \2217  = \2216  & ~\1 ,
  \2218  = \1037  & \71 ,
  \2219  = ~\1037  & \11 ,
  \2220  = \2219  | \2218 ,
  \2221  = ~\3  & \2 ,
  \2222  = \2221  & ~\1 ,
  \2223  = ~\1036  & \101 ,
  \2224  = \1036  & \11 ,
  \2225  = \2224  | \2223 ,
  \2226  = ~\3  & \2 ,
  \2227  = \2226  & ~\1 ,
  \2228  = \1037  & \70 ,
  \2229  = ~\1037  & \10 ,
  \2230  = \2229  | \2228 ,
  \2231  = ~\3  & \2 ,
  \2232  = \2231  & ~\1 ,
  \2233  = ~\1036  & \100 ,
  \2234  = \1036  & \10 ,
  \2235  = \2234  | \2233 ,
  \2236  = ~\3  & \2 ,
  \2237  = \2236  & ~\1 ,
  \2238  = \1037  & \69 ,
  \2239  = ~\1037  & \9 ,
  \2240  = \2239  | \2238 ,
  \2241  = ~\3  & \2 ,
  \2242  = \2241  & ~\1 ,
  \2243  = ~\1036  & \99 ,
  \2244  = \1036  & \9 ,
  \2245  = \2244  | \2243 ,
  \2246  = ~\3  & \2 ,
  \2247  = \2246  & ~\1 ,
  \2248  = \1037  & \68 ,
  \2249  = ~\1037  & \8 ,
  \2250  = \2249  | \2248 ,
  \2251  = ~\3  & \2 ,
  \2252  = \2251  & ~\1 ,
  \2253  = ~\1036  & \98 ,
  \2254  = \1036  & \8 ,
  \2255  = \2254  | \2253 ,
  \2256  = ~\3  & \2 ,
  \2257  = \2256  & ~\1 ,
  \2258  = \1037  & \67 ,
  \2259  = ~\1037  & \7 ,
  \2260  = \2259  | \2258 ,
  \2261  = ~\3  & \2 ,
  \2262  = \2261  & ~\1 ,
  \2263  = ~\1036  & \97 ,
  \2264  = \1036  & \7 ,
  \2265  = \2264  | \2263 ,
  \2266  = ~\3  & \2 ,
  \2267  = \2266  & ~\1 ,
  \2268  = \1037  & \66 ,
  \2269  = ~\1037  & \6 ,
  \2270  = \2269  | \2268 ,
  \2271  = ~\3  & \2 ,
  \2272  = \2271  & ~\1 ,
  \2273  = ~\1036  & \96 ,
  \2274  = \1036  & \6 ,
  \2275  = \2274  | \2273 ,
  \2276  = ~\3  & \2 ,
  \2277  = \2276  & ~\1 ,
  \2278  = \1037  & \65 ,
  \2279  = ~\1037  & \5 ,
  \2280  = \2279  | \2278 ,
  \2281  = ~\3  & \2 ,
  \2282  = \2281  & ~\1 ,
  \2283  = ~\1036  & \95 ,
  \2284  = \1036  & \5 ,
  \2285  = \2284  | \2283 ,
  \2286  = ~\3  & \2 ,
  \2287  = \2286  & ~\1 ,
  \2288  = \1037  & \64 ,
  \2289  = ~\1037  & \4 ,
  \2290  = \2289  | \2288 ,
  \2291  = ~\3  & \2 ,
  \2292  = \2291  & ~\1 ,
  \2293  = ~\1036  & \94 ,
  \2294  = \1036  & \4 ,
  \2295  = \2294  | \2293 ,
  \2296  = ~\3  & \2 ,
  \2297  = \2296  & ~\1 ,
  \2299  = \371  & \4 ,
  \2301  = \2299  & ~\369 ,
  \2302  = \369  & \5 ,
  \2303  = \2302  | \2301 ,
  \2304  = \2303  & ~\367 ,
  \2305  = \367  & \6 ,
  \2306  = \2305  | \2304 ,
  \2307  = \2306  & ~\365 ,
  \2308  = \365  & \7 ,
  \2309  = \2308  | \2307 ,
  \2310  = \2309  & ~\363 ,
  \2311  = \363  & \8 ,
  \2312  = \2311  | \2310 ,
  \2313  = \2312  & ~\361 ,
  \2314  = \361  & \9 ,
  \2315  = \2314  | \2313 ,
  \2316  = \2315  & ~\359 ,
  \2317  = \359  & \10 ,
  \2318  = \2317  | \2316 ,
  \2319  = \2318  & ~\357 ,
  \2320  = \357  & \11 ,
  \2321  = \2320  | \2319 ,
  \2322  = \2321  & ~\355 ,
  \2323  = \355  & \12 ,
  \2324  = \2323  | \2322 ,
  \2325  = \2324  & ~\353 ,
  \2326  = \353  & \13 ,
  \2327  = \2326  | \2325 ,
  \2328  = \2327  & ~\351 ,
  \2329  = \351  & \14 ,
  \2330  = \2329  | \2328 ,
  \2331  = \2330  & ~\349 ,
  \2332  = \349  & \15 ,
  \2333  = \2332  | \2331 ,
  \2334  = \2333  & ~\347 ,
  \2335  = \347  & \16 ,
  \2336  = \2335  | \2334 ,
  \2337  = \2336  & ~\345 ,
  \2338  = \345  & \17 ,
  \2339  = \2338  | \2337 ,
  \2340  = \2339  & ~\343 ,
  \2341  = \343  & \18 ,
  \2342  = \2341  | \2340 ,
  \2343  = \2342  & ~\341 ,
  \2344  = \341  & \19 ,
  \2345  = \2344  | \2343 ,
  \2346  = \2345  & ~\339 ,
  \2347  = \339  & \20 ,
  \2348  = \2347  | \2346 ,
  \2349  = \2348  & ~\337 ,
  \2350  = \337  & \21 ,
  \2351  = \2350  | \2349 ,
  \2352  = \2351  & ~\335 ,
  \2353  = \335  & \22 ,
  \2354  = \2353  | \2352 ,
  \2355  = \2354  & ~\333 ,
  \2356  = \333  & \23 ,
  \2357  = \2356  | \2355 ,
  \2358  = \2357  & ~\331 ,
  \2359  = \331  & \24 ,
  \2360  = \2359  | \2358 ,
  \2361  = \2360  & ~\329 ,
  \2362  = \329  & \25 ,
  \2363  = \2362  | \2361 ,
  \2364  = \2363  & ~\327 ,
  \2365  = \327  & \26 ,
  \2366  = \2365  | \2364 ,
  \2367  = \2366  & ~\325 ,
  \2368  = \325  & \27 ,
  \2369  = \2368  | \2367 ,
  \2370  = \2369  & ~\323 ,
  \2371  = \323  & \28 ,
  \2372  = \2371  | \2370 ,
  \2373  = \2372  & ~\321 ,
  \2374  = \321  & \29 ,
  \2375  = \2374  | \2373 ,
  \2376  = \2375  & ~\319 ,
  \2377  = \319  & \30 ,
  \2378  = \2377  | \2376 ,
  \2379  = \2378  & ~\317 ,
  \2380  = \317  & \31 ,
  \2381  = \2380  | \2379 ,
  \2382  = \2381  & ~\315 ,
  \2383  = \315  & \32 ,
  \2384  = \2383  | \2382 ,
  \2385  = \2384  & ~\313 ,
  \2386  = \313  & \33 ,
  \2387  = \2386  | \2385 ,
  \2388  = ~\3  & \2 ,
  \2389  = \2388  & ~\1 ,
  \2391  = \309  & \4 ,
  \2393  = \2391  & ~\307 ,
  \2394  = \307  & \5 ,
  \2395  = \2394  | \2393 ,
  \2396  = \2395  & ~\305 ,
  \2397  = \305  & \6 ,
  \2398  = \2397  | \2396 ,
  \2399  = \2398  & ~\303 ,
  \2400  = \303  & \7 ,
  \2401  = \2400  | \2399 ,
  \2402  = \2401  & ~\301 ,
  \2403  = \301  & \8 ,
  \2404  = \2403  | \2402 ,
  \2405  = \2404  & ~\299 ,
  \2406  = \299  & \9 ,
  \2407  = \2406  | \2405 ,
  \2408  = \2407  & ~\297 ,
  \2409  = \297  & \10 ,
  \2410  = \2409  | \2408 ,
  \2411  = \2410  & ~\295 ,
  \2412  = \295  & \11 ,
  \2413  = \2412  | \2411 ,
  \2414  = \2413  & ~\293 ,
  \2415  = \293  & \12 ,
  \2416  = \2415  | \2414 ,
  \2417  = \2416  & ~\291 ,
  \2418  = \291  & \13 ,
  \2419  = \2418  | \2417 ,
  \2420  = \2419  & ~\289 ,
  \2421  = \289  & \14 ,
  \2422  = \2421  | \2420 ,
  \2423  = \2422  & ~\287 ,
  \2424  = \287  & \15 ,
  \2425  = \2424  | \2423 ,
  \2426  = \2425  & ~\285 ,
  \2427  = \285  & \16 ,
  \2428  = \2427  | \2426 ,
  \2429  = \2428  & ~\283 ,
  \2430  = \283  & \17 ,
  \2431  = \2430  | \2429 ,
  \2432  = \2431  & ~\281 ,
  \2433  = \281  & \18 ,
  \2434  = \2433  | \2432 ,
  \2435  = \2434  & ~\279 ,
  \2436  = \279  & \19 ,
  \2437  = \2436  | \2435 ,
  \2438  = \2437  & ~\277 ,
  \2439  = \277  & \20 ,
  \2440  = \2439  | \2438 ,
  \2441  = \2440  & ~\275 ,
  \2442  = \275  & \21 ,
  \2443  = \2442  | \2441 ,
  \2444  = \2443  & ~\273 ,
  \2445  = \273  & \22 ,
  \2446  = \2445  | \2444 ,
  \2447  = \2446  & ~\271 ,
  \2448  = \271  & \23 ,
  \2449  = \2448  | \2447 ,
  \2450  = \2449  & ~\269 ,
  \2451  = \269  & \24 ,
  \2452  = \2451  | \2450 ,
  \2453  = \2452  & ~\267 ,
  \2454  = \267  & \25 ,
  \2455  = \2454  | \2453 ,
  \2456  = \2455  & ~\265 ,
  \2457  = \265  & \26 ,
  \2458  = \2457  | \2456 ,
  \2459  = \2458  & ~\263 ,
  \2460  = \263  & \27 ,
  \2461  = \2460  | \2459 ,
  \2462  = \2461  & ~\261 ,
  \2463  = \261  & \28 ,
  \2464  = \2463  | \2462 ,
  \2465  = \2464  & ~\259 ,
  \2466  = \259  & \29 ,
  \2467  = \2466  | \2465 ,
  \2468  = \2467  & ~\257 ,
  \2469  = \257  & \30 ,
  \2470  = \2469  | \2468 ,
  \2471  = \2470  & ~\255 ,
  \2472  = \255  & \31 ,
  \2473  = \2472  | \2471 ,
  \2474  = \2473  & ~\253 ,
  \2475  = \253  & \32 ,
  \2476  = \2475  | \2474 ,
  \2477  = \2476  & ~\251 ,
  \2478  = \251  & \33 ,
  \2479  = \2478  | \2477 ,
  \2480  = ~\3  & \2 ,
  \2481  = \2480  & ~\1 ,
  \124  = \1134 ,
  \125  = \1142 ,
  \126  = \1150 ,
  \127  = \1158 ,
  \128  = \1166 ,
  \129  = \1174 ,
  \130  = \1182 ,
  \131  = \1190 ,
  \132  = \1198 ,
  \133  = \1206 ,
  \134  = \1214 ,
  \135  = \1222 ,
  \136  = \1230 ,
  \137  = \1238 ,
  \138  = \1246 ,
  \139  = \1254 ,
  \140  = \1262 ,
  \141  = \1270 ,
  \142  = \1278 ,
  \143  = \1286 ,
  \144  = \1294 ,
  \145  = \1302 ,
  \146  = \1310 ,
  \147  = \1318 ,
  \148  = \1326 ,
  \149  = \1334 ,
  \150  = \1342 ,
  \151  = \1350 ,
  \152  = \1358 ,
  \153  = \1366 ,
  \184  = \1524  | \1 ,
  \185  = \1532  | \1 ,
  \186  = \1540  | \1 ,
  \187  = \1548  | \1 ,
  \188  = \1556  | \1 ,
  \189  = \1564  | \1 ,
  \190  = \1572  | \1 ,
  \191  = \1580  | \1 ,
  \192  = \1588  | \1 ,
  \193  = \1596  | \1 ,
  \194  = \1604  | \1 ,
  \195  = \1612  | \1 ,
  \196  = \1620  | \1 ,
  \197  = \1628  | \1 ,
  \198  = \1636  | \1 ,
  \199  = \1644  | \1 ,
  \200  = \1652  | \1 ,
  \201  = \1660  | \1 ,
  \202  = \1668  | \1 ,
  \203  = \1676  | \1 ,
  \204  = \1684  | \1 ,
  \205  = \1692  | \1 ,
  \206  = \1700  | \1 ,
  \207  = \1708  | \1 ,
  \208  = \1716  | \1 ,
  \209  = \1724  | \1 ,
  \210  = \1732  | \1 ,
  \211  = \1740  | \1 ,
  \212  = \1748  | \1 ,
  \213  = \1756  | \1 ,
  \251  = (~\33  & \123 ) | (\33  & ~\123 ),
  \253  = (~\32  & \122 ) | (\32  & ~\122 ),
  \255  = (~\31  & \121 ) | (\31  & ~\121 ),
  \257  = (~\30  & \120 ) | (\30  & ~\120 ),
  \259  = (~\29  & \119 ) | (\29  & ~\119 ),
  \261  = (~\28  & \118 ) | (\28  & ~\118 ),
  \263  = (~\27  & \117 ) | (\27  & ~\117 ),
  \265  = (~\26  & \116 ) | (\26  & ~\116 ),
  \267  = (~\25  & \115 ) | (\25  & ~\115 ),
  \269  = (~\24  & \114 ) | (\24  & ~\114 ),
  \271  = (~\23  & \113 ) | (\23  & ~\113 ),
  \273  = (~\22  & \112 ) | (\22  & ~\112 ),
  \275  = (~\21  & \111 ) | (\21  & ~\111 ),
  \277  = (~\20  & \110 ) | (\20  & ~\110 ),
  \279  = (~\19  & \109 ) | (\19  & ~\109 ),
  \281  = (~\18  & \108 ) | (\18  & ~\108 ),
  \283  = (~\17  & \107 ) | (\17  & ~\107 ),
  \285  = (~\16  & \106 ) | (\16  & ~\106 ),
  \287  = (~\15  & \105 ) | (\15  & ~\105 ),
  \289  = (~\14  & \104 ) | (\14  & ~\104 ),
  \291  = (~\13  & \103 ) | (\13  & ~\103 ),
  \293  = (~\12  & \102 ) | (\12  & ~\102 ),
  \295  = (~\11  & \101 ) | (\11  & ~\101 ),
  \297  = (~\10  & \100 ) | (\10  & ~\100 ),
  \299  = (~\9  & \99 ) | (\9  & ~\99 ),
  \301  = (~\8  & \98 ) | (\8  & ~\98 ),
  \303  = (~\7  & \97 ) | (\7  & ~\97 ),
  \305  = (~\6  & \96 ) | (\6  & ~\96 ),
  \307  = (~\5  & \95 ) | (\5  & ~\95 ),
  \309  = (~\4  & \94 ) | (\4  & ~\94 ),
  \313  = (~\33  & \93 ) | (\33  & ~\93 ),
  \315  = (~\32  & \92 ) | (\32  & ~\92 ),
  \317  = (~\31  & \91 ) | (\31  & ~\91 ),
  \319  = (~\30  & \90 ) | (\30  & ~\90 ),
  \321  = (~\29  & \89 ) | (\29  & ~\89 ),
  \323  = (~\28  & \88 ) | (\28  & ~\88 ),
  \325  = (~\27  & \87 ) | (\27  & ~\87 ),
  \327  = (~\26  & \86 ) | (\26  & ~\86 ),
  \329  = (~\25  & \85 ) | (\25  & ~\85 ),
  \331  = (~\24  & \84 ) | (\24  & ~\84 ),
  \333  = (~\23  & \83 ) | (\23  & ~\83 ),
  \335  = (~\22  & \82 ) | (\22  & ~\82 ),
  \337  = (~\21  & \81 ) | (\21  & ~\81 ),
  \339  = (~\20  & \80 ) | (\20  & ~\80 ),
  \341  = (~\19  & \79 ) | (\19  & ~\79 ),
  \343  = (~\18  & \78 ) | (\18  & ~\78 ),
  \345  = (~\17  & \77 ) | (\17  & ~\77 ),
  \347  = (~\16  & \76 ) | (\16  & ~\76 ),
  \349  = (~\15  & \75 ) | (\15  & ~\75 ),
  \351  = (~\14  & \74 ) | (\14  & ~\74 ),
  \353  = (~\13  & \73 ) | (\13  & ~\73 ),
  \355  = (~\12  & \72 ) | (\12  & ~\72 ),
  \357  = (~\11  & \71 ) | (\11  & ~\71 ),
  \359  = (~\10  & \70 ) | (\10  & ~\70 ),
  \361  = (~\9  & \69 ) | (\9  & ~\69 ),
  \363  = (~\8  & \68 ) | (\8  & ~\68 ),
  \365  = (~\7  & \67 ) | (\7  & ~\67 ),
  \367  = (~\6  & \66 ) | (\6  & ~\66 ),
  \369  = (~\5  & \65 ) | (\5  & ~\65 ),
  \371  = (~\4  & \64 ) | (\4  & ~\64 ),
  \[120]  = \1371 ,
  \[121]  = \1376 ,
  \[122]  = \1381 ,
  \[123]  = \1386 ,
  \[124]  = \1391 ,
  \[125]  = \1396 ,
  \[126]  = \1401 ,
  \[127]  = \1406 ,
  \[128]  = \1411 ,
  \[129]  = \1416 ,
  \[130]  = \1421 ,
  \[131]  = \1426 ,
  \[132]  = \1431 ,
  \[133]  = \1436 ,
  \[134]  = \1441 ,
  \[135]  = \1446 ,
  \[136]  = \1451 ,
  \[137]  = \1456 ,
  \[138]  = \1461 ,
  \[139]  = \1466 ,
  \[140]  = \1471 ,
  \[141]  = \1476 ,
  \[142]  = \1481 ,
  \[143]  = \1486 ,
  \[144]  = \1491 ,
  \[145]  = \1496 ,
  \[146]  = \1501 ,
  \[147]  = \1506 ,
  \[148]  = \1511 ,
  \[149]  = \1516 ,
  \[150]  = \184 ,
  \[151]  = \185 ,
  \[152]  = \186 ,
  \[153]  = \187 ,
  \[154]  = \188 ,
  \[155]  = \189 ,
  \[156]  = \190 ,
  \[157]  = \191 ,
  \[158]  = \192 ,
  \[159]  = \193 ,
  \[160]  = \194 ,
  \[161]  = \195 ,
  \[162]  = \196 ,
  \[163]  = \197 ,
  \[164]  = \198 ,
  \[165]  = \199 ,
  \[166]  = \200 ,
  \[167]  = \201 ,
  \[168]  = \202 ,
  \[169]  = \203 ,
  \916  = (\1127  & \1126 ) | ((\1127  & \1125 ) | (\1126  & \1125 )),
  \917  = (~\1043  & (~\1042  & \1041 )) | ((~\1043  & (\1042  & ~\1041 )) | ((\1043  & (~\1042  & ~\1041 )) | (\1043  & (\1042  & \1041 )))),
  \918  = (~\1046  & (~\1045  & \1044 )) | ((~\1046  & (\1045  & ~\1044 )) | ((\1046  & (~\1045  & ~\1044 )) | (\1046  & (\1045  & \1044 )))),
  \919  = (~\1049  & (~\1048  & \1047 )) | ((~\1049  & (\1048  & ~\1047 )) | ((\1049  & (~\1048  & ~\1047 )) | (\1049  & (\1048  & \1047 )))),
  \920  = (~\1052  & (~\1051  & \1050 )) | ((~\1052  & (\1051  & ~\1050 )) | ((\1052  & (~\1051  & ~\1050 )) | (\1052  & (\1051  & \1050 )))),
  \921  = (~\1055  & (~\1054  & \1053 )) | ((~\1055  & (\1054  & ~\1053 )) | ((\1055  & (~\1054  & ~\1053 )) | (\1055  & (\1054  & \1053 )))),
  \922  = (~\1058  & (~\1057  & \1056 )) | ((~\1058  & (\1057  & ~\1056 )) | ((\1058  & (~\1057  & ~\1056 )) | (\1058  & (\1057  & \1056 )))),
  \923  = (~\1061  & (~\1060  & \1059 )) | ((~\1061  & (\1060  & ~\1059 )) | ((\1061  & (~\1060  & ~\1059 )) | (\1061  & (\1060  & \1059 )))),
  \924  = (~\1064  & (~\1063  & \1062 )) | ((~\1064  & (\1063  & ~\1062 )) | ((\1064  & (~\1063  & ~\1062 )) | (\1064  & (\1063  & \1062 )))),
  \925  = (~\1067  & (~\1066  & \1065 )) | ((~\1067  & (\1066  & ~\1065 )) | ((\1067  & (~\1066  & ~\1065 )) | (\1067  & (\1066  & \1065 )))),
  \926  = (~\1070  & (~\1069  & \1068 )) | ((~\1070  & (\1069  & ~\1068 )) | ((\1070  & (~\1069  & ~\1068 )) | (\1070  & (\1069  & \1068 )))),
  \927  = (~\1073  & (~\1072  & \1071 )) | ((~\1073  & (\1072  & ~\1071 )) | ((\1073  & (~\1072  & ~\1071 )) | (\1073  & (\1072  & \1071 )))),
  \928  = (~\1076  & (~\1075  & \1074 )) | ((~\1076  & (\1075  & ~\1074 )) | ((\1076  & (~\1075  & ~\1074 )) | (\1076  & (\1075  & \1074 )))),
  \929  = (~\1079  & (~\1078  & \1077 )) | ((~\1079  & (\1078  & ~\1077 )) | ((\1079  & (~\1078  & ~\1077 )) | (\1079  & (\1078  & \1077 )))),
  \930  = (~\1082  & (~\1081  & \1080 )) | ((~\1082  & (\1081  & ~\1080 )) | ((\1082  & (~\1081  & ~\1080 )) | (\1082  & (\1081  & \1080 )))),
  \931  = (~\1085  & (~\1084  & \1083 )) | ((~\1085  & (\1084  & ~\1083 )) | ((\1085  & (~\1084  & ~\1083 )) | (\1085  & (\1084  & \1083 )))),
  \932  = (~\1088  & (~\1087  & \1086 )) | ((~\1088  & (\1087  & ~\1086 )) | ((\1088  & (~\1087  & ~\1086 )) | (\1088  & (\1087  & \1086 )))),
  \933  = (~\1091  & (~\1090  & \1089 )) | ((~\1091  & (\1090  & ~\1089 )) | ((\1091  & (~\1090  & ~\1089 )) | (\1091  & (\1090  & \1089 )))),
  \934  = (~\1094  & (~\1093  & \1092 )) | ((~\1094  & (\1093  & ~\1092 )) | ((\1094  & (~\1093  & ~\1092 )) | (\1094  & (\1093  & \1092 )))),
  \935  = (~\1097  & (~\1096  & \1095 )) | ((~\1097  & (\1096  & ~\1095 )) | ((\1097  & (~\1096  & ~\1095 )) | (\1097  & (\1096  & \1095 )))),
  \936  = (~\1100  & (~\1099  & \1098 )) | ((~\1100  & (\1099  & ~\1098 )) | ((\1100  & (~\1099  & ~\1098 )) | (\1100  & (\1099  & \1098 )))),
  \937  = (~\1103  & (~\1102  & \1101 )) | ((~\1103  & (\1102  & ~\1101 )) | ((\1103  & (~\1102  & ~\1101 )) | (\1103  & (\1102  & \1101 )))),
  \938  = (~\1106  & (~\1105  & \1104 )) | ((~\1106  & (\1105  & ~\1104 )) | ((\1106  & (~\1105  & ~\1104 )) | (\1106  & (\1105  & \1104 )))),
  \939  = (~\1109  & (~\1108  & \1107 )) | ((~\1109  & (\1108  & ~\1107 )) | ((\1109  & (~\1108  & ~\1107 )) | (\1109  & (\1108  & \1107 )))),
  \940  = (~\1112  & (~\1111  & \1110 )) | ((~\1112  & (\1111  & ~\1110 )) | ((\1112  & (~\1111  & ~\1110 )) | (\1112  & (\1111  & \1110 )))),
  \941  = (~\1115  & (~\1114  & \1113 )) | ((~\1115  & (\1114  & ~\1113 )) | ((\1115  & (~\1114  & ~\1113 )) | (\1115  & (\1114  & \1113 )))),
  \942  = (~\1118  & (~\1117  & \1116 )) | ((~\1118  & (\1117  & ~\1116 )) | ((\1118  & (~\1117  & ~\1116 )) | (\1118  & (\1117  & \1116 )))),
  \943  = (~\1121  & (~\1120  & \1119 )) | ((~\1121  & (\1120  & ~\1119 )) | ((\1121  & (~\1120  & ~\1119 )) | (\1121  & (\1120  & \1119 )))),
  \944  = (~\1124  & (~\1123  & \1122 )) | ((~\1124  & (\1123  & ~\1122 )) | ((\1124  & (~\1123  & ~\1122 )) | (\1124  & (\1123  & \1122 )))),
  \945  = (~\1127  & (~\1126  & \1125 )) | ((~\1127  & (\1126  & ~\1125 )) | ((\1127  & (~\1126  & ~\1125 )) | (\1127  & (\1126  & \1125 )))),
  \[170]  = \204 ,
  \[171]  = \205 ,
  \[172]  = \206 ,
  \[173]  = \207 ,
  \1036  = \2481  & \2479 ,
  \1037  = \2389  & \2387 ,
  \1039  = \2297  & \2295 ,
  \[174]  = \208 ,
  \1040  = \2292  & \2290 ,
  \1041  = \1040  & \1039 ,
  \1042  = \2287  & \2285 ,
  \1043  = \2282  & \2280 ,
  \1044  = (\1043  & \1042 ) | ((\1043  & \1041 ) | (\1042  & \1041 )),
  \1045  = \2277  & \2275 ,
  \1046  = \2272  & \2270 ,
  \1047  = (\1046  & \1045 ) | ((\1046  & \1044 ) | (\1045  & \1044 )),
  \1048  = \2267  & \2265 ,
  \1049  = \2262  & \2260 ,
  \[175]  = \209 ,
  \1050  = (\1049  & \1048 ) | ((\1049  & \1047 ) | (\1048  & \1047 )),
  \1051  = \2257  & \2255 ,
  \1052  = \2252  & \2250 ,
  \1053  = (\1052  & \1051 ) | ((\1052  & \1050 ) | (\1051  & \1050 )),
  \1054  = \2247  & \2245 ,
  \1055  = \2242  & \2240 ,
  \1056  = (\1055  & \1054 ) | ((\1055  & \1053 ) | (\1054  & \1053 )),
  \1057  = \2237  & \2235 ,
  \1058  = \2232  & \2230 ,
  \1059  = (\1058  & \1057 ) | ((\1058  & \1056 ) | (\1057  & \1056 )),
  \[176]  = \210 ,
  \1060  = \2227  & \2225 ,
  \1061  = \2222  & \2220 ,
  \1062  = (\1061  & \1060 ) | ((\1061  & \1059 ) | (\1060  & \1059 )),
  \1063  = \2217  & \2215 ,
  \1064  = \2212  & \2210 ,
  \1065  = (\1064  & \1063 ) | ((\1064  & \1062 ) | (\1063  & \1062 )),
  \1066  = \2207  & \2205 ,
  \1067  = \2202  & \2200 ,
  \1068  = (\1067  & \1066 ) | ((\1067  & \1065 ) | (\1066  & \1065 )),
  \1069  = \2197  & \2195 ,
  \[177]  = \211 ,
  \1070  = \2192  & \2190 ,
  \1071  = (\1070  & \1069 ) | ((\1070  & \1068 ) | (\1069  & \1068 )),
  \1072  = \2187  & \2185 ,
  \1073  = \2182  & \2180 ,
  \1074  = (\1073  & \1072 ) | ((\1073  & \1071 ) | (\1072  & \1071 )),
  \1075  = \2177  & \2175 ,
  \1076  = \2172  & \2170 ,
  \1077  = (\1076  & \1075 ) | ((\1076  & \1074 ) | (\1075  & \1074 )),
  \1078  = \2167  & \2165 ,
  \1079  = \2162  & \2160 ,
  \[178]  = \212 ,
  \1080  = (\1079  & \1078 ) | ((\1079  & \1077 ) | (\1078  & \1077 )),
  \1081  = \2157  & \2155 ,
  \1082  = \2152  & \2150 ,
  \1083  = (\1082  & \1081 ) | ((\1082  & \1080 ) | (\1081  & \1080 )),
  \1084  = \2147  & \2145 ,
  \1085  = \2142  & \2140 ,
  \1086  = (\1085  & \1084 ) | ((\1085  & \1083 ) | (\1084  & \1083 )),
  \1087  = \2137  & \2135 ,
  \1088  = \2132  & \2130 ,
  \1089  = (\1088  & \1087 ) | ((\1088  & \1086 ) | (\1087  & \1086 )),
  \[179]  = \213 ,
  \1090  = \2127  & \2125 ,
  \1091  = \2122  & \2120 ,
  \1092  = (\1091  & \1090 ) | ((\1091  & \1089 ) | (\1090  & \1089 )),
  \1093  = \2117  & \2115 ,
  \1094  = \2112  & \2110 ,
  \1095  = (\1094  & \1093 ) | ((\1094  & \1092 ) | (\1093  & \1092 )),
  \1096  = \2107  & \2105 ,
  \1097  = \2102  & \2100 ,
  \1098  = (\1097  & \1096 ) | ((\1097  & \1095 ) | (\1096  & \1095 )),
  \1099  = \2097  & \2095 ,
  \[180]  = \1764 ,
  \1100  = \2092  & \2090 ,
  \1101  = (\1100  & \1099 ) | ((\1100  & \1098 ) | (\1099  & \1098 )),
  \1102  = \2087  & \2085 ,
  \1103  = \2082  & \2080 ,
  \1104  = (\1103  & \1102 ) | ((\1103  & \1101 ) | (\1102  & \1101 )),
  \1105  = \2077  & \2075 ,
  \1106  = \2072  & \2070 ,
  \1107  = (\1106  & \1105 ) | ((\1106  & \1104 ) | (\1105  & \1104 )),
  \1108  = \2067  & \2065 ,
  \1109  = \2062  & \2060 ,
  \[181]  = \1772 ,
  \1110  = (\1109  & \1108 ) | ((\1109  & \1107 ) | (\1108  & \1107 )),
  \1111  = \2057  & \2055 ,
  \1112  = \2052  & \2050 ,
  \1113  = (\1112  & \1111 ) | ((\1112  & \1110 ) | (\1111  & \1110 )),
  \1114  = \2047  & \2045 ,
  \1115  = \2042  & \2040 ,
  \1116  = (\1115  & \1114 ) | ((\1115  & \1113 ) | (\1114  & \1113 )),
  \1117  = \2037  & \2035 ,
  \1118  = \2032  & \2030 ,
  \1119  = (\1118  & \1117 ) | ((\1118  & \1116 ) | (\1117  & \1116 )),
  \[182]  = \1780 ,
  \1120  = \2027  & \2025 ,
  \1121  = \2022  & \2020 ,
  \1122  = (\1121  & \1120 ) | ((\1121  & \1119 ) | (\1120  & \1119 )),
  \1123  = \2017  & \2015 ,
  \1124  = \2012  & \2010 ,
  \1125  = (\1124  & \1123 ) | ((\1124  & \1122 ) | (\1123  & \1122 )),
  \1126  = \2007  & \2005 ,
  \1127  = \2002  & \2000 ,
  \1128  = \917  & ~\3 ,
  \1129  = \4  & \3 ,
  \[183]  = \1788 ,
  \1130  = \1129  | \1128 ,
  \1131  = \1130  & \2 ,
  \1132  = \34  & ~\2 ,
  \1133  = \1132  | \1131 ,
  \1134  = \1133  & ~\1 ,
  \1136  = \918  & ~\3 ,
  \1137  = \5  & \3 ,
  \1138  = \1137  | \1136 ,
  \1139  = \1138  & \2 ,
  \[184]  = \1796 ,
  \1140  = \35  & ~\2 ,
  \1141  = \1140  | \1139 ,
  \1142  = \1141  & ~\1 ,
  \1144  = \919  & ~\3 ,
  \1145  = \6  & \3 ,
  \1146  = \1145  | \1144 ,
  \1147  = \1146  & \2 ,
  \1148  = \36  & ~\2 ,
  \1149  = \1148  | \1147 ,
  \[185]  = \1804 ,
  \1150  = \1149  & ~\1 ,
  \1152  = \920  & ~\3 ,
  \1153  = \7  & \3 ,
  \1154  = \1153  | \1152 ,
  \1155  = \1154  & \2 ,
  \1156  = \37  & ~\2 ,
  \1157  = \1156  | \1155 ,
  \1158  = \1157  & ~\1 ,
  \[186]  = \1812 ,
  \1160  = \921  & ~\3 ,
  \1161  = \8  & \3 ,
  \1162  = \1161  | \1160 ,
  \1163  = \1162  & \2 ,
  \1164  = \38  & ~\2 ,
  \1165  = \1164  | \1163 ,
  \1166  = \1165  & ~\1 ,
  \1168  = \922  & ~\3 ,
  \1169  = \9  & \3 ,
  \[187]  = \1820 ,
  \1170  = \1169  | \1168 ,
  \1171  = \1170  & \2 ,
  \1172  = \39  & ~\2 ,
  \1173  = \1172  | \1171 ,
  \1174  = \1173  & ~\1 ,
  \1176  = \923  & ~\3 ,
  \1177  = \10  & \3 ,
  \1178  = \1177  | \1176 ,
  \1179  = \1178  & \2 ,
  \[188]  = \1828 ;
always begin
  \34  = \[120] ;
  \35  = \[121] ;
  \36  = \[122] ;
  \37  = \[123] ;
  \38  = \[124] ;
  \39  = \[125] ;
  \40  = \[126] ;
  \41  = \[127] ;
  \42  = \[128] ;
  \43  = \[129] ;
  \44  = \[130] ;
  \45  = \[131] ;
  \46  = \[132] ;
  \47  = \[133] ;
  \48  = \[134] ;
  \49  = \[135] ;
  \50  = \[136] ;
  \51  = \[137] ;
  \52  = \[138] ;
  \53  = \[139] ;
  \54  = \[140] ;
  \55  = \[141] ;
  \56  = \[142] ;
  \57  = \[143] ;
  \58  = \[144] ;
  \59  = \[145] ;
  \60  = \[146] ;
  \61  = \[147] ;
  \62  = \[148] ;
  \63  = \[149] ;
  \64  = \[150] ;
  \65  = \[151] ;
  \66  = \[152] ;
  \67  = \[153] ;
  \68  = \[154] ;
  \69  = \[155] ;
  \70  = \[156] ;
  \71  = \[157] ;
  \72  = \[158] ;
  \73  = \[159] ;
  \74  = \[160] ;
  \75  = \[161] ;
  \76  = \[162] ;
  \77  = \[163] ;
  \78  = \[164] ;
  \79  = \[165] ;
  \80  = \[166] ;
  \81  = \[167] ;
  \82  = \[168] ;
  \83  = \[169] ;
  \84  = \[170] ;
  \85  = \[171] ;
  \86  = \[172] ;
  \87  = \[173] ;
  \88  = \[174] ;
  \89  = \[175] ;
  \90  = \[176] ;
  \91  = \[177] ;
  \92  = \[178] ;
  \93  = \[179] ;
  \94  = \[180] ;
  \95  = \[181] ;
  \96  = \[182] ;
  \97  = \[183] ;
  \98  = \[184] ;
  \99  = \[185] ;
  \100  = \[186] ;
  \101  = \[187] ;
  \102  = \[188] ;
  \103  = \[189] ;
  \104  = \[190] ;
  \105  = \[191] ;
  \106  = \[192] ;
  \107  = \[193] ;
  \108  = \[194] ;
  \109  = \[195] ;
  \110  = \[196] ;
  \111  = \[197] ;
  \112  = \[198] ;
  \113  = \[199] ;
  \114  = \[200] ;
  \115  = \[201] ;
  \116  = \[202] ;
  \117  = \[203] ;
  \118  = \[204] ;
  \119  = \[205] ;
  \120  = \[206] ;
  \121  = \[207] ;
  \122  = \[208] ;
  \123  = \[209] ;
end
initial begin
  \64  = 1;
  \65  = 1;
  \66  = 1;
  \67  = 1;
  \68  = 1;
  \69  = 1;
  \70  = 1;
  \71  = 1;
  \72  = 1;
  \73  = 1;
  \74  = 1;
  \75  = 1;
  \76  = 1;
  \77  = 1;
  \78  = 1;
  \79  = 1;
  \80  = 1;
  \81  = 1;
  \82  = 1;
  \83  = 1;
  \84  = 1;
  \85  = 1;
  \86  = 1;
  \87  = 1;
  \88  = 1;
  \89  = 1;
  \90  = 1;
  \91  = 1;
  \92  = 1;
  \93  = 1;
  \94  = 0;
  \95  = 0;
  \96  = 0;
  \97  = 0;
  \98  = 0;
  \99  = 0;
  \100  = 0;
  \101  = 0;
  \102  = 0;
  \103  = 0;
  \104  = 0;
  \105  = 0;
  \106  = 0;
  \107  = 0;
  \108  = 0;
  \109  = 0;
  \110  = 0;
  \111  = 0;
  \112  = 0;
  \113  = 0;
  \114  = 0;
  \115  = 0;
  \116  = 0;
  \117  = 0;
  \118  = 0;
  \119  = 0;
  \120  = 0;
  \121  = 0;
  \122  = 0;
  \123  = 0;
end
endmodule

