//NOTE: no-implementation module stub

module GtCLK_OR2 (
    output Z,
    input A,
    input B
);

endmodule
