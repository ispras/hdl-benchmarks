module test ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , 
 n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , 
 n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , 
 n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , 
 n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , 
 n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , 
 n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , 
 n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , 
 n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , 
 n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , 
 n181 , n182 , n183 , n184 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 ;
output n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , 
 n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , 
 n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , 
 n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , 
 n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , 
 n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , 
 n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , 
 n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , 
 n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , 
 n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , 
 n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , 
 n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , 
 n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 ;
wire n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , 
 n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , 
 n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , 
 n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , 
 n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , 
 n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , 
 n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , 
 n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , 
 n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , 
 n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , 
 n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , 
 n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , 
 n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , 
 n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , 
 n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , 
 n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , 
 n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , 
 n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , 
 n551 , n552 , n553 , n554 , n40212 , n40213 , n40214 , n40215 , n40216 , n40217 , 
 n40218 , n40219 , n40220 , n40221 , n40222 , n40223 , n40224 , n40225 , n40226 , n40227 , 
 n40228 , n40229 , n40230 , n40231 , n40232 , n40233 , n40234 , n40235 , n40236 , n40237 , 
 n40238 , n40239 , n40240 , n40241 , n40242 , n40243 , n40244 , n40245 , n40246 , n40247 , 
 n40248 , n40249 , n40250 , n40251 , n40252 , n40253 , n40254 , n40255 , n40256 , n40257 , 
 n40258 , n40259 , n40260 , n40261 , n40262 , n40263 , n40264 , n40265 , n40266 , n40267 , 
 n40268 , n40269 , n40270 , n40271 , n40272 , n40273 , n40274 , n40275 , n40276 , n40277 , 
 n40278 , n40279 , n40280 , n40281 , n40282 , n40283 , n40284 , n40285 , n40286 , n40287 , 
 n40288 , n40289 , n40290 , n40291 , n40292 , n40293 , n40294 , n40295 , n40296 , n40297 , 
 n40298 , n40299 , n40300 , n40301 , n40302 , n40303 , n40304 , n40305 , n40306 , n40307 , 
 n40308 , n40309 , n40310 , n40311 , n40312 , n40313 , n40314 , n40315 , n40316 , n40317 , 
 n40318 , n40319 , n40320 , n40321 , n40322 , n40323 , n40324 , n40325 , n40326 , n40327 , 
 n40328 , n40329 , n40330 , n40331 , n40332 , n40333 , n40334 , n40335 , n40336 , n40337 , 
 n40338 , n40339 , n40340 , n40341 , n40342 , n40343 , n40344 , n40345 , n40346 , n40347 , 
 n40348 , n40349 , n40350 , n40351 , n40352 , n40353 , n40354 , n40355 , n40356 , n40357 , 
 n40358 , n40359 , n40360 , n40361 , n40362 , n40363 , n40364 , n40365 , n40366 , n40367 , 
 n40368 , n40369 , n40370 , n40371 , n40372 , n40373 , n40374 , n40375 , n40376 , n40377 , 
 n40378 , n40379 , n40380 , n40381 , n40382 , n40383 , n40384 , n40385 , n40386 , n40387 , 
 n40388 , n40389 , n40390 , n40391 , n40392 , n40393 , n40394 , n40395 , n40396 , n40397 , 
 n40398 , n40399 , n40400 , n40401 , n40402 , n40403 , n40404 , n40405 , n40406 , n40407 , 
 n40408 , n40409 , n40410 , n40411 , n40412 , n40413 , n40414 , n40415 , n40416 , n40417 , 
 n40418 , n40419 , n40420 , n40421 , n40422 , n40423 , n40424 , n40425 , n40426 , n40427 , 
 n40428 , n40429 , n40430 , n40431 , n40432 , n40433 , n40434 , n40435 , n40436 , n40437 , 
 n40438 , n40439 , n40440 , n40441 , n40442 , n40443 , n40444 , n40445 , n40446 , n40447 , 
 n40448 , n40449 , n40450 , n40451 , n40452 , n40453 , n40454 , n40455 , n40456 , n40457 , 
 n40458 , n40459 , n40460 , n40461 , n40462 , n40463 , n40464 , n40465 , n40466 , n40467 , 
 n40468 , n40469 , n40470 , n40471 , n40472 , n40473 , n40474 , n40475 , n40476 , n40477 , 
 n40478 , n40479 , n40480 , n40481 , n40482 , n40483 , n40484 , n40485 , n40486 , n40487 , 
 n40488 , n40489 , n40490 , n40491 , n40492 , n40493 , n40494 , n40495 , n40496 , n40497 , 
 n40498 , n40499 , n40500 , n40501 , n40502 , n40503 , n40504 , n40505 , n40506 , n40507 , 
 n40508 , n40509 , n40510 , n40511 , n40512 , n40513 , n40514 , n40515 , n40516 , n40517 , 
 n40518 , n40519 , n40520 , n40521 , n40522 , n40523 , n40524 , n40525 , n40526 , n40527 , 
 n40528 , n40529 , n40530 , n40531 , n40532 , n40533 , n40534 , n40535 , n40536 , n40537 , 
 n40538 , n40539 , n40540 , n40541 , n40542 , n40543 , n40544 , n40545 , n40546 , n40547 , 
 n40548 , n40549 , n40550 , n40551 , n40552 , n40553 , n40554 , n40555 , n40556 , n40557 , 
 n40558 , n40559 , n40560 , n40561 , n40562 , n40563 , n40564 , n40565 , n40566 , n40567 , 
 n40568 , n40569 , n40570 , n40571 , n40572 , n40573 , n40574 , n40575 , n40576 , n40577 , 
 n40578 , n40579 , n40580 , n40581 , n40582 , n40583 , n40584 , n40585 , n40586 , n40587 , 
 n40588 , n40589 , n40590 , n40591 , n40592 , n40593 , n40594 , n40595 , n40596 , n40597 , 
 n40598 , n40599 , n40600 , n40601 , n40602 , n40603 , n40604 , n40605 , n40606 , n40607 , 
 n40608 , n40609 , n40610 , n40611 , n40612 , n40613 , n40614 , n40615 , n40616 , n40617 , 
 n40618 , n40619 , n40620 , n40621 , n40622 , n40623 , n40624 , n40625 , n40626 , n40627 , 
 n40628 , n40629 , n40630 , n40631 , n40632 , n40633 , n40634 , n40635 , n40636 , n40637 , 
 n40638 , n40639 , n40640 , n40641 , n40642 , n40643 , n40644 , n40645 , n40646 , n40647 , 
 n40648 , n40649 , n40650 , n40651 , n40652 , n40653 , n40654 , n40655 , n40656 , n40657 , 
 n40658 , n40659 , n40660 , n40661 , n40662 , n40663 , n40664 , n40665 , n40666 , n40667 , 
 n40668 , n40669 , n40670 , n40671 , n40672 , n40673 , n40674 , n40675 , n40676 , n40677 , 
 n40678 , n40679 , n40680 , n40681 , n40682 , n40683 , n40684 , n40685 , n40686 , n40687 , 
 n40688 , n40689 , n40690 , n40691 , n40692 , n40693 , n40694 , n40695 , n40696 , n40697 , 
 n40698 , n40699 , n40700 , n40701 , n40702 , n40703 , n40704 , n40705 , n40706 , n40707 , 
 n40708 , n40709 , n40710 , n40711 , n40712 , n40713 , n40714 , n40715 , n40716 , n40717 , 
 n40718 , n40719 , n40720 , n40721 , n40722 , n40723 , n40724 , n40725 , n40726 , n40727 , 
 n40728 , n40729 , n40730 , n40731 , n40732 , n40733 , n40734 , n40735 , n40736 , n40737 , 
 n40738 , n40739 , n40740 , n40741 , n40742 , n40743 , n40744 , n40745 , n40746 , n40747 , 
 n40748 , n40749 , n40750 , n40751 , n40752 , n40753 , n40754 , n40755 , n40756 , n40757 , 
 n40758 , n40759 , n40760 , n40761 , n40762 , n40763 , n40764 , n40765 , n40766 , n40767 , 
 n40768 , n40769 , n40770 , n40771 , n40772 , n40773 , n40774 , n40775 , n40776 , n40777 , 
 n40778 , n40779 , n40780 , n40781 , n40782 , n40783 , n40784 , n40785 , n40786 , n40787 , 
 n40788 , n40789 , n40790 , n40791 , n40792 , n40793 , n40794 , n40795 , n40796 , n40797 , 
 n40798 , n40799 , n40800 , n40801 , n40802 , n40803 , n40804 , n40805 , n40806 , n40807 , 
 n40808 , n40809 , n40810 , n40811 , n40812 , n40813 , n40814 , n40815 , n40816 , n40817 , 
 n40818 , n40819 , n40820 , n40821 , n40822 , n40823 , n40824 , n40825 , n40826 , n40827 , 
 n40828 , n40829 , n40830 , n40831 , n40832 , n40833 , n40834 , n40835 , n40836 , n40837 , 
 n40838 , n40839 , n40840 , n40841 , n40842 , n40843 , n40844 , n40845 , n40846 , n40847 , 
 n40848 , n40849 , n40850 , n40851 , n40852 , n40853 , n40854 , n40855 , n40856 , n40857 , 
 n40858 , n40859 , n40860 , n40861 , n40862 , n40863 , n40864 , n40865 , n40866 , n40867 , 
 n40868 , n40869 , n40870 , n40871 , n40872 , n40873 , n40874 , n40875 , n40876 , n40877 , 
 n40878 , n40879 , n40880 , n40881 , n40882 , n40883 , n40884 , n40885 , n40886 , n40887 , 
 n40888 , n40889 , n40890 , n40891 , n40892 , n40893 , n40894 , n40895 , n40896 , n40897 , 
 n40898 , n40899 , n40900 , n40901 , n40902 , n40903 , n40904 , n40905 , n40906 , n40907 , 
 n40908 , n40909 , n40910 , n40911 , n40912 , n40913 , n40914 , n40915 , n40916 , n40917 , 
 n40918 , n40919 , n40920 , n40921 , n40922 , n40923 , n40924 , n40925 , n40926 , n40927 , 
 n40928 , n40929 , n40930 , n40931 , n40932 , n40933 , n40934 , n40935 , n40936 , n40937 , 
 n40938 , n40939 , n40940 , n40941 , n40942 , n40943 , n40944 , n40945 , n40946 , n40947 , 
 n40948 , n40949 , n40950 , n40951 , n40952 , n40953 , n40954 , n40955 , n40956 , n40957 , 
 n40958 , n40959 , n40960 , n40961 , n40962 , n40963 , n40964 , n40965 , n40966 , n40967 , 
 n40968 , n40969 , n40970 , n40971 , n40972 , n40973 , n40974 , n40975 , n40976 , n40977 , 
 n40978 , n40979 , n40980 , n40981 , n40982 , n40983 , n40984 , n40985 , n40986 , n40987 , 
 n40988 , n40989 , n40990 , n40991 , n40992 , n40993 , n40994 , n40995 , n40996 , n40997 , 
 n40998 , n40999 , n41000 , n41001 , n41002 , n41003 , n41004 , n41005 , n41006 , n41007 , 
 n41008 , n41009 , n41010 , n41011 , n41012 , n41013 , n41014 , n41015 , n41016 , n41017 , 
 n41018 , n41019 , n41020 , n41021 , n41022 , n41023 , n41024 , n41025 , n41026 , n41027 , 
 n41028 , n41029 , n41030 , n41031 , n41032 , n41033 , n41034 , n41035 , n41036 , n41037 , 
 n41038 , n41039 , n41040 , n41041 , n41042 , n41043 , n41044 , n41045 , n41046 , n41047 , 
 n41048 , n41049 , n41050 , n41051 , n41052 , n41053 , n41054 , n41055 , n41056 , n41057 , 
 n41058 , n41059 , n41060 , n41061 , n41062 , n41063 , n41064 , n41065 , n41066 , n41067 , 
 n41068 , n41069 , n41070 , n41071 , n41072 , n41073 , n41074 , n41075 , n41076 , n41077 , 
 n41078 , n41079 , n41080 , n41081 , n41082 , n41083 , n41084 , n41085 , n41086 , n41087 , 
 n41088 , n41089 , n41090 , n41091 , n41092 , n41093 , n41094 , n41095 , n41096 , n41097 , 
 n41098 , n41099 , n41100 , n41101 , n41102 , n41103 , n41104 , n41105 , n41106 , n41107 , 
 n41108 , n41109 , n41110 , n41111 , n41112 , n41113 , n41114 , n41115 , n41116 , n41117 , 
 n41118 , n41119 , n41120 , n41121 , n41122 , n41123 , n41124 , n41125 , n41126 , n41127 , 
 n41128 , n41129 , n41130 , n41131 , n41132 , n41133 , n41134 , n41135 , n41136 , n41137 , 
 n41138 , n41139 , n41140 , n41141 , n41142 , n41143 , n41144 , n41145 , n41146 , n41147 , 
 n41148 , n41149 , n41150 , n41151 , n41152 , n41153 , n41154 , n41155 , n41156 , n41157 , 
 n41158 , n41159 , n41160 , n41161 , n41162 , n41163 , n41164 , n41165 , n41166 , n41167 , 
 n41168 , n41169 , n41170 , n41171 , n41172 , n41173 , n41174 , n41175 , n41176 , n41177 , 
 n41178 , n41179 , n41180 , n41181 , n41182 , n41183 , n41184 , n41185 , n41186 , n41187 , 
 n41188 , n41189 , n41190 , n41191 , n41192 , n41193 , n41194 , n41195 , n41196 , n41197 , 
 n41198 , n41199 , n41200 , n41201 , n41202 , n41203 , n41204 , n41205 , n41206 , n41207 , 
 n41208 , n41209 , n41210 , n41211 , n41212 , n41213 , n41214 , n41215 , n41216 , n41217 , 
 n41218 , n41219 , n41220 , n41221 , n41222 , n41223 , n41224 , n41225 , n41226 , n41227 , 
 n41228 , n41229 , n41230 , n41231 , n41232 , n41233 , n41234 , n41235 , n41236 , n41237 , 
 n41238 , n41239 , n41240 , n41241 , n41242 , n41243 , n41244 , n41245 , n41246 , n41247 , 
 n41248 , n41249 , n41250 , n41251 , n41252 , n41253 , n41254 , n41255 , n41256 , n41257 , 
 n41258 , n41259 , n41260 , n41261 , n41262 , n41263 , n41264 , n41265 , n41266 , n41267 , 
 n41268 , n41269 , n41270 , n41271 , n41272 , n41273 , n41274 , n41275 , n41276 , n41277 , 
 n41278 , n41279 , n41280 , n41281 , n41282 , n41283 , n41284 , n41285 , n41286 , n41287 , 
 n41288 , n41289 , n41290 , n41291 , n41292 , n41293 , n41294 , n41295 , n41296 , n41297 , 
 n41298 , n41299 , n41300 , n41301 , n41302 , n41303 , n41304 , n41305 , n41306 , n41307 , 
 n41308 , n41309 , n41310 , n41311 , n41312 , n41313 , n41314 , n41315 , n41316 , n41317 , 
 n41318 , n41319 , n41320 , n41321 , n41322 , n41323 , n41324 , n41325 , n41326 , n41327 , 
 n41328 , n41329 , n41330 , n41331 , n41332 , n41333 , n41334 , n41335 , n41336 , n41337 , 
 n41338 , n41339 , n41340 , n41341 , n41342 , n41343 , n41344 , n41345 , n41346 , n41347 , 
 n41348 , n41349 , n41350 , n41351 , n41352 , n41353 , n41354 , n41355 , n41356 , n41357 , 
 n41358 , n41359 , n41360 , n41361 , n41362 , n41363 , n41364 , n41365 , n41366 , n41367 , 
 n41368 , n41369 , n41370 , n41371 , n41372 , n41373 , n41374 , n41375 , n41376 , n41377 , 
 n41378 , n41379 , n41380 , n41381 , n41382 , n41383 , n41384 , n41385 , n41386 , n41387 , 
 n41388 , n41389 , n41390 , n41391 , n41392 , n41393 , n41394 , n41395 , n41396 , n41397 , 
 n41398 , n41399 , n41400 , n41401 , n41402 , n41403 , n41404 , n41405 , n41406 , n41407 , 
 n41408 , n41409 , n41410 , n41411 , n41412 , n41413 , n41414 , n41415 , n41416 , n41417 , 
 n41418 , n41419 , n41420 , n41421 , n41422 , n41423 , n41424 , n41425 , n41426 , n41427 , 
 n41428 , n41429 , n41430 , n41431 , n41432 , n41433 , n41434 , n41435 , n41436 , n41437 , 
 n41438 , n41439 , n41440 , n41441 , n41442 , n41443 , n41444 , n41445 , n41446 , n41447 , 
 n41448 , n41449 , n41450 , n41451 , n41452 , n41453 , n41454 , n41455 , n41456 , n41457 , 
 n41458 , n41459 , n41460 , n41461 , n41462 , n41463 , n41464 , n41465 , n41466 , n41467 , 
 n41468 , n41469 , n41470 , n41471 , n41472 , n41473 , n41474 , n41475 , n41476 , n41477 , 
 n41478 , n41479 , n41480 , n41481 , n41482 , n41483 , n41484 , n41485 , n41486 , n41487 , 
 n41488 , n41489 , n41490 , n41491 , n41492 , n41493 , n41494 , n41495 , n41496 , n41497 , 
 n41498 , n41499 , n41500 , n41501 , n41502 , n41503 , n41504 , n41505 , n41506 , n41507 , 
 n41508 , n41509 , n41510 , n41511 , n41512 , n41513 , n41514 , n41515 , n41516 , n41517 , 
 n41518 , n41519 , n41520 , n41521 , n41522 , n41523 , n41524 , n41525 , n41526 , n41527 , 
 n41528 , n41529 , n41530 , n41531 , n41532 , n41533 , n41534 , n41535 , n41536 , n41537 , 
 n41538 , n41539 , n41540 , n41541 , n41542 , n41543 , n41544 , n41545 , n41546 , n41547 , 
 n41548 , n41549 , n41550 , n41551 , n41552 , n41553 , n41554 , n41555 , n41556 , n41557 , 
 n41558 , n41559 , n41560 , n41561 , n41562 , n41563 , n41564 , n41565 , n41566 , n41567 , 
 n41568 , n41569 , n41570 , n41571 , n41572 , n41573 , n41574 , n41575 , n41576 , n41577 , 
 n41578 , n41579 , n41580 , n41581 , n41582 , n41583 , n41584 , n41585 , n41586 , n41587 , 
 n41588 , n41589 , n41590 , n41591 , n41592 , n41593 , n41594 , n41595 , n41596 , n41597 , 
 n41598 , n41599 , n41600 , n41601 , n41602 , n41603 , n41604 , n41605 , n41606 , n41607 , 
 n41608 , n41609 , n41610 , n41611 , n41612 , n41613 , n41614 , n41615 , n41616 , n41617 , 
 n41618 , n41619 , n41620 , n41621 , n41622 , n41623 , n41624 , n41625 , n41626 , n41627 , 
 n41628 , n41629 , n41630 , n41631 , n41632 , n41633 , n41634 , n41635 , n41636 , n41637 , 
 n41638 , n41639 , n41640 , n41641 , n41642 , n41643 , n41644 , n41645 , n41646 , n41647 , 
 n41648 , n41649 , n41650 , n41651 , n41652 , n41653 , n41654 , n41655 , n41656 , n41657 , 
 n41658 , n41659 , n41660 , n41661 , n41662 , n41663 , n41664 , n41665 , n41666 , n41667 , 
 n41668 , n41669 , n41670 , n41671 , n41672 , n41673 , n41674 , n41675 , n41676 , n41677 , 
 n41678 , n41679 , n41680 , n41681 , n41682 , n41683 , n41684 , n41685 , n41686 , n41687 , 
 n41688 , n41689 , n41690 , n41691 , n41692 , n41693 , n41694 , n41695 , n41696 , n41697 , 
 n41698 , n41699 , n41700 , n41701 , n41702 , n41703 , n41704 , n41705 , n41706 , n41707 , 
 n41708 , n41709 , n41710 , n41711 , n41712 , n41713 , n41714 , n41715 , n41716 , n41717 , 
 n41718 , n41719 , n41720 , n41721 , n41722 , n41723 , n41724 , n41725 , n41726 , n41727 , 
 n41728 , n41729 , n41730 , n41731 , n41732 , n41733 , n41734 , n41735 , n41736 , n41737 , 
 n41738 , n41739 , n41740 , n41741 , n41742 , n41743 , n41744 , n41745 , n41746 , n41747 , 
 n41748 , n41749 , n41750 , n41751 , n41752 , n41753 , n41754 , n41755 , n41756 , n41757 , 
 n41758 , n41759 , n41760 , n41761 , n41762 , n41763 , n41764 , n41765 , n41766 , n41767 , 
 n41768 , n41769 , n41770 , n41771 , n41772 , n41773 , n41774 , n41775 , n41776 , n41777 , 
 n41778 , n41779 , n41780 , n41781 , n41782 , n41783 , n41784 , n41785 , n41786 , n41787 , 
 n41788 , n41789 , n41790 , n41791 , n41792 , n41793 , n41794 , n41795 , n41796 , n41797 , 
 n41798 , n41799 , n41800 , n41801 , n41802 , n41803 , n41804 , n41805 , n41806 , n41807 , 
 n41808 , n41809 , n41810 , n41811 , n41812 , n41813 , n41814 , n41815 , n41816 , n41817 , 
 n41818 , n41819 , n41820 , n41821 , n41822 , n41823 , n41824 , n41825 , n41826 , n41827 , 
 n41828 , n41829 , n41830 , n41831 , n41832 , n41833 , n41834 , n41835 , n41836 , n41837 , 
 n41838 , n41839 , n41840 , n41841 , n41842 , n41843 , n41844 , n41845 , n41846 , n41847 , 
 n41848 , n41849 , n41850 , n41851 , n41852 , n41853 , n41854 , n41855 , n41856 , n41857 , 
 n41858 , n41859 , n41860 , n41861 , n41862 , n41863 , n41864 , n41865 , n41866 , n41867 , 
 n41868 , n41869 , n41870 , n41871 , n41872 , n41873 , n41874 , n41875 , n41876 , n41877 , 
 n41878 , n41879 , n41880 , n41881 , n41882 , n41883 , n41884 , n41885 , n41886 , n41887 , 
 n41888 , n41889 , n41890 , n41891 , n41892 , n41893 , n41894 , n41895 , n41896 , n41897 , 
 n41898 , n41899 , n41900 , n41901 , n41902 , n41903 , n41904 , n41905 , n41906 , n41907 , 
 n41908 , n41909 , n41910 , n41911 , n41912 , n41913 , n41914 , n41915 , n41916 , n41917 , 
 n41918 , n41919 , n41920 , n41921 , n41922 , n41923 , n41924 , n41925 , n41926 , n41927 , 
 n41928 , n41929 , n41930 , n41931 , n41932 , n41933 , n41934 , n41935 , n41936 , n41937 , 
 n41938 , n41939 , n41940 , n41941 , n41942 , n41943 , n41944 , n41945 , n41946 , n41947 , 
 n41948 , n41949 , n41950 , n41951 , n41952 , n41953 , n41954 , n41955 , n41956 , n41957 , 
 n41958 , n41959 , n41960 , n41961 , n41962 , n41963 , n41964 , n41965 , n41966 , n41967 , 
 n41968 , n41969 , n41970 , n41971 , n41972 , n41973 , n41974 , n41975 , n41976 , n41977 , 
 n41978 , n41979 , n41980 , n41981 , n41982 , n41983 , n41984 , n41985 , n41986 , n41987 , 
 n41988 , n41989 , n41990 , n41991 , n41992 , n41993 , n41994 , n41995 , n41996 , n41997 , 
 n41998 , n41999 , n42000 , n42001 , n42002 , n42003 , n42004 , n42005 , n42006 , n42007 , 
 n42008 , n42009 , n42010 , n42011 , n42012 , n42013 , n42014 , n42015 , n42016 , n42017 , 
 n42018 , n42019 , n42020 , n42021 , n42022 , n42023 , n42024 , n42025 , n42026 , n42027 , 
 n42028 , n42029 , n42030 , n42031 , n42032 , n42033 , n42034 , n42035 , n42036 , n42037 , 
 n42038 , n42039 , n42040 , n42041 , n42042 , n42043 , n42044 , n42045 , n42046 , n42047 , 
 n42048 , n42049 , n42050 , n42051 , n42052 , n42053 , n42054 , n42055 , n42056 , n42057 , 
 n42058 , n42059 , n42060 , n42061 , n42062 , n42063 , n42064 , n42065 , n42066 , n42067 , 
 n42068 , n42069 , n42070 , n42071 , n42072 , n42073 , n42074 , n42075 , n42076 , n42077 , 
 n42078 , n42079 , n42080 , n42081 , n42082 , n42083 , n42084 , n42085 , n42086 , n42087 , 
 n42088 , n42089 , n42090 , n42091 , n42092 , n42093 , n42094 , n42095 , n42096 , n42097 , 
 n42098 , n42099 , n42100 , n42101 , n42102 , n42103 , n42104 , n42105 , n42106 , n42107 , 
 n42108 , n42109 , n42110 , n42111 , n42112 , n42113 , n42114 , n42115 , n42116 , n42117 , 
 n42118 , n42119 , n42120 , n42121 , n42122 , n42123 , n42124 , n42125 , n42126 , n42127 , 
 n42128 , n42129 , n42130 , n42131 , n42132 , n42133 , n42134 , n42135 , n42136 , n42137 , 
 n42138 , n42139 , n42140 , n42141 , n42142 , n42143 , n42144 , n42145 , n42146 , n42147 , 
 n42148 , n42149 , n42150 , n42151 , n42152 , n42153 , n42154 , n42155 , n42156 , n42157 , 
 n42158 , n42159 , n42160 , n42161 , n42162 , n42163 , n42164 , n42165 , n42166 , n42167 , 
 n42168 , n42169 , n42170 , n42171 , n42172 , n42173 , n42174 , n42175 , n42176 , n42177 , 
 n42178 , n42179 , n42180 , n42181 , n42182 , n42183 , n42184 , n42185 , n42186 , n42187 , 
 n42188 , n42189 , n42190 , n42191 , n42192 , n42193 , n42194 , n42195 , n42196 , n42197 , 
 n42198 , n42199 , n42200 , n42201 , n42202 , n42203 , n42204 , n42205 , n42206 , n42207 , 
 n42208 , n42209 , n42210 , n42211 , n42212 , n42213 , n42214 , n42215 , n42216 , n42217 , 
 n42218 , n42219 , n42220 , n42221 , n42222 , n42223 , n42224 , n42225 , n42226 , n42227 , 
 n42228 , n42229 , n42230 , n42231 , n42232 , n42233 , n42234 , n42235 , n42236 , n42237 , 
 n42238 , n42239 , n42240 , n42241 , n42242 , n42243 , n42244 , n42245 , n42246 , n42247 , 
 n42248 , n42249 , n42250 , n42251 , n42252 , n42253 , n42254 , n42255 , n42256 , n42257 , 
 n42258 , n42259 , n42260 , n42261 , n42262 , n42263 , n42264 , n42265 , n42266 , n42267 , 
 n42268 , n42269 , n42270 , n42271 , n42272 , n42273 , n42274 , n42275 , n42276 , n42277 , 
 n42278 , n42279 , n42280 , n42281 , n42282 , n42283 , n42284 , n42285 , n42286 , n42287 , 
 n42288 , n42289 , n42290 , n42291 , n42292 , n42293 , n42294 , n42295 , n42296 , n42297 , 
 n42298 , n42299 , n42300 , n42301 , n42302 , n42303 , n42304 , n42305 , n42306 , n42307 , 
 n42308 , n42309 , n42310 , n42311 , n42312 , n42313 , n42314 , n42315 , n42316 , n42317 , 
 n42318 , n42319 , n42320 , n42321 , n42322 , n42323 , n42324 , n42325 , n42326 , n42327 , 
 n42328 , n42329 , n42330 , n42331 , n42332 , n42333 , n42334 , n42335 , n42336 , n42337 , 
 n42338 , n42339 , n42340 , n42341 , n42342 , n42343 , n42344 , n42345 , n42346 , n42347 , 
 n42348 , n42349 , n42350 , n42351 , n42352 , n42353 , n42354 , n42355 , n42356 , n42357 , 
 n42358 , n42359 , n42360 , n42361 , n42362 , n42363 , n42364 , n42365 , n42366 , n42367 , 
 n42368 , n42369 , n42370 , n42371 , n42372 , n42373 , n42374 , n42375 , n42376 , n42377 , 
 n42378 , n42379 , n42380 , n42381 , n42382 , n42383 , n42384 , n42385 , n42386 , n42387 , 
 n42388 , n42389 , n42390 , n42391 , n42392 , n42393 , n42394 , n42395 , n42396 , n42397 , 
 n42398 , n42399 , n42400 , n42401 , n42402 , n42403 , n42404 , n42405 , n42406 , n42407 , 
 n42408 , n42409 , n42410 , n42411 , n42412 , n42413 , n42414 , n42415 , n42416 , n42417 , 
 n42418 , n42419 , n42420 , n42421 , n42422 , n42423 , n42424 , n42425 , n42426 , n42427 , 
 n42428 , n42429 , n42430 , n42431 , n42432 , n42433 , n42434 , n42435 , n42436 , n42437 , 
 n42438 , n42439 , n42440 , n42441 , n42442 , n42443 , n42444 , n42445 , n42446 , n42447 , 
 n42448 , n42449 , n42450 , n42451 , n42452 , n42453 , n42454 , n42455 , n42456 , n42457 , 
 n42458 , n42459 , n42460 , n42461 , n42462 , n42463 , n42464 , n42465 , n42466 , n42467 , 
 n42468 , n42469 , n42470 , n42471 , n42472 , n42473 , n42474 , n42475 , n42476 , n42477 , 
 n42478 , n42479 , n42480 , n42481 , n42482 , n42483 , n42484 , n42485 , n42486 , n42487 , 
 n42488 , n42489 , n42490 , n42491 , n42492 , n42493 , n42494 , n42495 , n42496 , n42497 , 
 n42498 , n42499 , n42500 , n42501 , n42502 , n42503 , n42504 , n42505 , n42506 , n42507 , 
 n42508 , n42509 , n42510 , n42511 , n42512 , n42513 , n42514 , n42515 , n42516 , n42517 , 
 n42518 , n42519 , n42520 , n42521 , n42522 , n42523 , n42524 , n42525 , n42526 , n42527 , 
 n42528 , n42529 , n42530 , n42531 , n42532 , n42533 , n42534 , n42535 , n42536 , n42537 , 
 n42538 , n42539 , n42540 , n42541 , n42542 , n42543 , n42544 , n42545 , n42546 , n42547 , 
 n42548 , n42549 , n42550 , n42551 , n42552 , n42553 , n42554 , n42555 , n42556 , n42557 , 
 n42558 , n42559 , n42560 , n42561 , n42562 , n42563 , n42564 , n42565 , n42566 , n42567 , 
 n42568 , n42569 , n42570 , n42571 , n42572 , n42573 , n42574 , n42575 , n42576 , n42577 , 
 n42578 , n42579 , n42580 , n42581 , n42582 , n42583 , n42584 , n42585 , n42586 , n42587 , 
 n42588 , n42589 , n42590 , n42591 , n42592 , n42593 , n42594 , n42595 , n42596 , n42597 , 
 n42598 , n42599 , n42600 , n42601 , n42602 , n42603 , n42604 , n42605 , n42606 , n42607 , 
 n42608 , n42609 , n42610 , n42611 , n42612 , n42613 , n42614 , n42615 , n42616 , n42617 , 
 n42618 , n42619 , n42620 , n42621 , n42622 , n42623 , n42624 , n42625 , n42626 , n42627 , 
 n42628 , n42629 , n42630 , n42631 , n42632 , n42633 , n42634 , n42635 , n42636 , n42637 , 
 n42638 , n42639 , n42640 , n42641 , n42642 , n42643 , n42644 , n42645 , n42646 , n42647 , 
 n42648 , n42649 , n42650 , n42651 , n42652 , n42653 , n42654 , n42655 , n42656 , n42657 , 
 n42658 , n42659 , n42660 , n42661 , n42662 , n42663 , n42664 , n42665 , n42666 , n42667 , 
 n42668 , n42669 , n42670 , n42671 , n42672 , n42673 , n42674 , n42675 , n42676 , n42677 , 
 n42678 , n42679 , n42680 , n42681 , n42682 , n42683 , n42684 , n42685 , n42686 , n42687 , 
 n42688 , n42689 , n42690 , n42691 , n42692 , n42693 , n42694 , n42695 , n42696 , n42697 , 
 n42698 , n42699 , n42700 , n42701 , n42702 , n42703 , n42704 , n42705 , n42706 , n42707 , 
 n42708 , n42709 , n42710 , n42711 , n42712 , n42713 , n42714 , n42715 , n42716 , n42717 , 
 n42718 , n42719 , n42720 , n42721 , n42722 , n42723 , n42724 , n42725 , n42726 , n42727 , 
 n42728 , n42729 , n42730 , n42731 , n42732 , n42733 , n42734 , n42735 , n42736 , n42737 , 
 n42738 , n42739 , n42740 , n42741 , n42742 , n42743 , n42744 , n42745 , n42746 , n42747 , 
 n42748 , n42749 , n42750 , n42751 , n42752 , n42753 , n42754 , n42755 , n42756 , n42757 , 
 n42758 , n42759 , n42760 , n42761 , n42762 , n42763 , n42764 , n42765 , n42766 , n42767 , 
 n42768 , n42769 , n42770 , n42771 , n42772 , n42773 , n42774 , n42775 , n42776 , n42777 , 
 n42778 , n42779 , n42780 , n42781 , n42782 , n42783 , n42784 , n42785 , n42786 , n42787 , 
 n42788 , n42789 , n42790 , n42791 , n42792 , n42793 , n42794 , n42795 , n42796 , n42797 , 
 n42798 , n42799 , n42800 , n42801 , n42802 , n42803 , n42804 , n42805 , n42806 , n42807 , 
 n42808 , n42809 , n42810 , n42811 , n42812 , n42813 , n42814 , n42815 , n42816 , n42817 , 
 n42818 , n42819 , n42820 , n42821 , n42822 , n42823 , n42824 , n42825 , n42826 , n42827 , 
 n42828 , n42829 , n42830 , n42831 , n42832 , n42833 , n42834 , n42835 , n42836 , n42837 , 
 n42838 , n42839 , n42840 , n42841 , n42842 , n42843 , n42844 , n42845 , n42846 , n42847 , 
 n42848 , n42849 , n42850 , n42851 , n42852 , n42853 , n42854 , n42855 , n42856 , n42857 , 
 n42858 , n42859 , n42860 , n42861 , n42862 , n42863 , n42864 , n42865 , n42866 , n42867 , 
 n42868 , n42869 , n42870 , n42871 , n42872 , n42873 , n42874 , n42875 , n42876 , n42877 , 
 n42878 , n42879 , n42880 , n42881 , n42882 , n42883 , n42884 , n42885 , n42886 , n42887 , 
 n42888 , n42889 , n42890 , n42891 , n42892 , n42893 , n42894 , n42895 , n42896 , n42897 , 
 n42898 , n42899 , n42900 , n42901 , n42902 , n42903 , n42904 , n42905 , n42906 , n42907 , 
 n42908 , n42909 , n42910 , n42911 , n42912 , n42913 , n42914 , n42915 , n42916 , n42917 , 
 n42918 , n42919 , n42920 , n42921 , n42922 , n42923 , n42924 , n42925 , n42926 , n42927 , 
 n42928 , n42929 , n42930 , n42931 , n42932 , n42933 , n42934 , n42935 , n42936 , n42937 , 
 n42938 , n42939 , n42940 , n42941 , n42942 , n42943 , n42944 , n42945 , n42946 , n42947 , 
 n42948 , n42949 , n42950 , n42951 , n42952 , n42953 , n42954 , n42955 , n42956 , n42957 , 
 n42958 , n42959 , n42960 , n42961 , n42962 , n42963 , n42964 , n42965 , n42966 , n42967 , 
 n42968 , n42969 , n42970 , n42971 , n42972 , n42973 , n42974 , n42975 , n42976 , n42977 , 
 n42978 , n42979 , n42980 , n42981 , n42982 , n42983 , n42984 , n42985 , n42986 , n42987 , 
 n42988 , n42989 , n42990 , n42991 , n42992 , n42993 , n42994 , n42995 , n42996 , n42997 , 
 n42998 , n42999 , n43000 , n43001 , n43002 , n43003 , n43004 , n43005 , n43006 , n43007 , 
 n43008 , n43009 , n43010 , n43011 , n43012 , n43013 , n43014 , n43015 , n43016 , n43017 , 
 n43018 , n43019 , n43020 , n43021 , n43022 , n43023 , n43024 , n43025 , n43026 , n43027 , 
 n43028 , n43029 , n43030 , n43031 , n43032 , n43033 , n43034 , n43035 , n43036 , n43037 , 
 n43038 , n43039 , n43040 , n43041 , n43042 , n43043 , n43044 , n43045 , n43046 , n43047 , 
 n43048 , n43049 , n43050 , n43051 , n43052 , n43053 , n43054 , n43055 , n43056 , n43057 , 
 n43058 , n43059 , n43060 , n43061 , n43062 , n43063 , n43064 , n43065 , n43066 , n43067 , 
 n43068 , n43069 , n43070 , n43071 , n43072 , n43073 , n43074 , n43075 , n43076 , n43077 , 
 n43078 , n43079 , n43080 , n43081 , n43082 , n43083 , n43084 , n43085 , n43086 , n43087 , 
 n43088 , n43089 , n43090 , n43091 , n43092 , n43093 , n43094 , n43095 , n43096 , n43097 , 
 n43098 , n43099 , n43100 , n43101 , n43102 , n43103 , n43104 , n43105 , n43106 , n43107 , 
 n43108 , n43109 , n43110 , n43111 , n43112 , n43113 , n43114 , n43115 , n43116 , n43117 , 
 n43118 , n43119 , n43120 , n43121 , n43122 , n43123 , n43124 , n43125 , n43126 , n43127 , 
 n43128 , n43129 , n43130 , n43131 , n43132 , n43133 , n43134 , n43135 , n43136 , n43137 , 
 n43138 , n43139 , n43140 , n43141 , n43142 , n43143 , n43144 , n43145 , n43146 , n43147 , 
 n43148 , n43149 , n43150 , n43151 , n43152 , n43153 , n43154 , n43155 , n43156 , n43157 , 
 n43158 , n43159 , n43160 , n43161 , n43162 , n43163 , n43164 , n43165 , n43166 , n43167 , 
 n43168 , n43169 , n43170 , n43171 , n43172 , n43173 , n43174 , n43175 , n43176 , n43177 , 
 n43178 , n43179 , n43180 , n43181 , n43182 , n43183 , n43184 , n43185 , n43186 , n43187 , 
 n43188 , n43189 , n43190 , n43191 , n43192 , n43193 , n43194 , n43195 , n43196 , n43197 , 
 n43198 , n43199 , n43200 , n43201 , n43202 , n43203 , n43204 , n43205 , n43206 , n43207 , 
 n43208 , n43209 , n43210 , n43211 , n43212 , n43213 , n43214 , n43215 , n43216 , n43217 , 
 n43218 , n43219 , n43220 , n43221 , n43222 , n43223 , n43224 , n43225 , n43226 , n43227 , 
 n43228 , n43229 , n43230 , n43231 , n43232 , n43233 , n43234 , n43235 , n43236 , n43237 , 
 n43238 , n43239 , n43240 , n43241 , n43242 , n43243 , n43244 , n43245 , n43246 , n43247 , 
 n43248 , n43249 , n43250 , n43251 , n43252 , n43253 , n43254 , n43255 , n43256 , n43257 , 
 n43258 , n43259 , n43260 , n43261 , n43262 , n43263 , n43264 , n43265 , n43266 , n43267 , 
 n43268 , n43269 , n43270 , n43271 , n43272 , n43273 , n43274 , n43275 , n43276 , n43277 , 
 n43278 , n43279 , n43280 , n43281 , n43282 , n43283 , n43284 , n43285 , n43286 , n43287 , 
 n43288 , n43289 , n43290 , n43291 , n43292 , n43293 , n43294 , n43295 , n43296 , n43297 , 
 n43298 , n43299 , n43300 , n43301 , n43302 , n43303 , n43304 , n43305 , n43306 , n43307 , 
 n43308 , n43309 , n43310 , n43311 , n43312 , n43313 , n43314 , n43315 , n43316 , n43317 , 
 n43318 , n43319 , n43320 , n43321 , n43322 , n43323 , n43324 , n43325 , n43326 , n43327 , 
 n43328 , n43329 , n43330 , n43331 , n43332 , n43333 , n43334 , n43335 , n43336 , n43337 , 
 n43338 , n43339 , n43340 , n43341 , n43342 , n43343 , n43344 , n43345 , n43346 , n43347 , 
 n43348 , n43349 , n43350 , n43351 , n43352 , n43353 , n43354 , n43355 , n43356 , n43357 , 
 n43358 , n43359 , n43360 , n43361 , n43362 , n43363 , n43364 , n43365 , n43366 , n43367 , 
 n43368 , n43369 , n43370 , n43371 , n43372 , n43373 , n43374 , n43375 , n43376 , n43377 , 
 n43378 , n43379 , n43380 , n43381 , n43382 , n43383 , n43384 , n43385 , n43386 , n43387 , 
 n43388 , n43389 , n43390 , n43391 , n43392 , n43393 , n43394 , n43395 , n43396 , n43397 , 
 n43398 , n43399 , n43400 , n43401 , n43402 , n43403 , n43404 , n43405 , n43406 , n43407 , 
 n43408 , n43409 , n43410 , n43411 , n43412 , n43413 , n43414 , n43415 , n43416 , n43417 , 
 n43418 , n43419 , n43420 , n43421 , n43422 , n43423 , n43424 , n43425 , n43426 , n43427 , 
 n43428 , n43429 , n43430 , n43431 , n43432 , n43433 , n43434 , n43435 , n43436 , n43437 , 
 n43438 , n43439 , n43440 , n43441 , n43442 , n43443 , n43444 , n43445 , n43446 , n43447 , 
 n43448 , n43449 , n43450 , n43451 , n43452 , n43453 , n43454 , n43455 , n43456 , n43457 , 
 n43458 , n43459 , n43460 , n43461 , n43462 , n43463 , n43464 , n43465 , n43466 , n43467 , 
 n43468 , n43469 , n43470 , n43471 , n43472 , n43473 , n43474 , n43475 , n43476 , n43477 , 
 n43478 , n43479 , n43480 , n43481 , n43482 , n43483 , n43484 , n43485 , n43486 , n43487 , 
 n43488 , n43489 , n43490 , n43491 , n43492 , n43493 , n43494 , n43495 , n43496 , n43497 , 
 n43498 , n43499 , n43500 , n43501 , n43502 , n43503 , n43504 , n43505 , n43506 , n43507 , 
 n43508 , n43509 , n43510 , n43511 , n43512 , n43513 , n43514 , n43515 , n43516 , n43517 , 
 n43518 , n43519 , n43520 , n43521 , n43522 , n43523 , n43524 , n43525 , n43526 , n43527 , 
 n43528 , n43529 , n43530 , n43531 , n43532 , n43533 , n43534 , n43535 , n43536 , n43537 , 
 n43538 , n43539 , n43540 , n43541 , n43542 , n43543 , n43544 , n43545 , n43546 , n43547 , 
 n43548 , n43549 , n43550 , n43551 , n43552 , n43553 , n43554 , n43555 , n43556 , n43557 , 
 n43558 , n43559 , n43560 , n43561 , n43562 , n43563 , n43564 , n43565 , n43566 , n43567 , 
 n43568 , n43569 , n43570 , n43571 , n43572 , n43573 , n43574 , n43575 , n43576 , n43577 , 
 n43578 , n43579 , n43580 , n43581 , n43582 , n43583 , n43584 , n43585 , n43586 , n43587 , 
 n43588 , n43589 , n43590 , n43591 , n43592 , n43593 , n43594 , n43595 , n43596 , n43597 , 
 n43598 , n43599 , n43600 , n43601 , n43602 , n43603 , n43604 , n43605 , n43606 , n43607 , 
 n43608 , n43609 , n43610 , n43611 , n43612 , n43613 , n43614 , n43615 , n43616 , n43617 , 
 n43618 , n43619 , n43620 , n43621 , n43622 , n43623 , n43624 , n43625 , n43626 , n43627 , 
 n43628 , n43629 , n43630 , n43631 , n43632 , n43633 , n43634 , n43635 , n43636 , n43637 , 
 n43638 , n43639 , n43640 , n43641 , n43642 , n43643 , n43644 , n43645 , n43646 , n43647 , 
 n43648 , n43649 , n43650 , n43651 , n43652 , n43653 , n43654 , n43655 , n43656 , n43657 , 
 n43658 , n43659 , n43660 , n43661 , n43662 , n43663 , n43664 , n43665 , n43666 , n43667 , 
 n43668 , n43669 , n43670 , n43671 , n43672 , n43673 , n43674 , n43675 , n43676 , n43677 , 
 n43678 , n43679 , n43680 , n43681 , n43682 , n43683 , n43684 , n43685 , n43686 , n43687 , 
 n43688 , n43689 , n43690 , n43691 , n43692 , n43693 , n43694 , n43695 , n43696 , n43697 , 
 n43698 , n43699 , n43700 , n43701 , n43702 , n43703 , n43704 , n43705 , n43706 , n43707 , 
 n43708 , n43709 , n43710 , n43711 , n43712 , n43713 , n43714 , n43715 , n43716 , n43717 , 
 n43718 , n43719 , n43720 , n43721 , n43722 , n43723 , n43724 , n43725 , n43726 , n43727 , 
 n43728 , n43729 , n43730 , n43731 , n43732 , n43733 , n43734 , n43735 , n43736 , n43737 , 
 n43738 , n43739 , n43740 , n43741 , n43742 , n43743 , n43744 , n43745 , n43746 , n43747 , 
 n43748 , n43749 , n43750 , n43751 , n43752 , n43753 , n43754 , n43755 , n43756 , n43757 , 
 n43758 , n43759 , n43760 , n43761 , n43762 , n43763 , n43764 , n43765 , n43766 , n43767 , 
 n43768 , n43769 , n43770 , n43771 , n43772 , n43773 , n43774 , n43775 , n43776 , n43777 , 
 n43778 , n43779 , n43780 , n43781 , n43782 , n43783 , n43784 , n43785 , n43786 , n43787 , 
 n43788 , n43789 , n43790 , n43791 , n43792 , n43793 , n43794 , n43795 , n43796 , n43797 , 
 n43798 , n43799 , n43800 , n43801 , n43802 , n43803 , n43804 , n43805 , n43806 , n43807 , 
 n43808 , n43809 , n43810 , n43811 , n43812 , n43813 , n43814 , n43815 , n43816 , n43817 , 
 n43818 , n43819 , n43820 , n43821 , n43822 , n43823 , n43824 , n43825 , n43826 , n43827 , 
 n43828 , n43829 , n43830 , n43831 , n43832 , n43833 , n43834 , n43835 , n43836 , n43837 , 
 n43838 , n43839 , n43840 , n43841 , n43842 , n43843 , n43844 , n43845 , n43846 , n43847 , 
 n43848 , n43849 , n43850 , n43851 , n43852 , n43853 , n43854 , n43855 , n43856 , n43857 , 
 n43858 , n43859 , n43860 , n43861 , n43862 , n43863 , n43864 , n43865 , n43866 , n43867 , 
 n43868 , n43869 , n43870 , n43871 , n43872 , n43873 , n43874 , n43875 , n43876 , n43877 , 
 n43878 , n43879 , n43880 , n43881 , n43882 , n43883 , n43884 , n43885 , n43886 , n43887 , 
 n43888 , n43889 , n43890 , n43891 , n43892 , n43893 , n43894 , n43895 , n43896 , n43897 , 
 n43898 , n43899 , n43900 , n43901 , n43902 , n43903 , n43904 , n43905 , n43906 , n43907 , 
 n43908 , n43909 , n43910 , n43911 , n43912 , n43913 , n43914 , n43915 , n43916 , n43917 , 
 n43918 , n43919 , n43920 , n43921 , n43922 , n43923 , n43924 , n43925 , n43926 , n43927 , 
 n43928 , n43929 , n43930 , n43931 , n43932 , n43933 , n43934 , n43935 , n43936 , n43937 , 
 n43938 , n43939 , n43940 , n43941 , n43942 , n43943 , n43944 , n43945 , n43946 , n43947 , 
 n43948 , n43949 , n43950 , n43951 , n43952 , n43953 , n43954 , n43955 , n43956 , n43957 , 
 n43958 , n43959 , n43960 , n43961 , n43962 , n43963 , n43964 , n43965 , n43966 , n43967 , 
 n43968 , n43969 , n43970 , n43971 , n43972 , n43973 , n43974 , n43975 , n43976 , n43977 , 
 n43978 , n43979 , n43980 , n43981 , n43982 , n43983 , n43984 , n43985 , n43986 , n43987 , 
 n43988 , n43989 , n43990 , n43991 , n43992 , n43993 , n43994 , n43995 , n43996 , n43997 , 
 n43998 , n43999 , n44000 , n44001 , n44002 , n44003 , n44004 , n44005 , n44006 , n44007 , 
 n44008 , n44009 , n44010 , n44011 , n44012 , n44013 , n44014 , n44015 , n44016 , n44017 , 
 n44018 , n44019 , n44020 , n44021 , n44022 , n44023 , n44024 , n44025 , n44026 , n44027 , 
 n44028 , n44029 , n44030 , n44031 , n44032 , n44033 , n44034 , n44035 , n44036 , n44037 , 
 n44038 , n44039 , n44040 , n44041 , n44042 , n44043 , n44044 , n44045 , n44046 , n44047 , 
 n44048 , n44049 , n44050 , n44051 , n44052 , n44053 , n44054 , n44055 , n44056 , n44057 , 
 n44058 , n44059 , n44060 , n44061 , n44062 , n44063 , n44064 , n44065 , n44066 , n44067 , 
 n44068 , n44069 , n44070 , n44071 , n44072 , n44073 , n44074 , n44075 , n44076 , n44077 , 
 n44078 , n44079 , n44080 , n44081 , n44082 , n44083 , n44084 , n44085 , n44086 , n44087 , 
 n44088 , n44089 , n44090 , n44091 , n44092 , n44093 , n44094 , n44095 , n44096 , n44097 , 
 n44098 , n44099 , n44100 , n44101 , n44102 , n44103 , n44104 , n44105 , n44106 , n44107 , 
 n44108 , n44109 , n44110 , n44111 , n44112 , n44113 , n44114 , n44115 , n44116 , n44117 , 
 n44118 , n44119 , n44120 , n44121 , n44122 , n44123 , n44124 , n44125 , n44126 , n44127 , 
 n44128 , n44129 , n44130 , n44131 , n44132 , n44133 , n44134 , n44135 , n44136 , n44137 , 
 n44138 , n44139 , n44140 , n44141 , n44142 , n44143 , n44144 , n44145 , n44146 , n44147 , 
 n44148 , n44149 , n44150 , n44151 , n44152 , n44153 , n44154 , n44155 , n44156 , n44157 , 
 n44158 , n44159 , n44160 , n44161 , n44162 , n44163 , n44164 , n44165 , n44166 , n44167 , 
 n44168 , n44169 , n44170 , n44171 , n44172 , n44173 , n44174 , n44175 , n44176 , n44177 , 
 n44178 , n44179 , n44180 , n44181 , n44182 , n44183 , n44184 , n44185 , n44186 , n44187 , 
 n44188 , n44189 , n44190 , n44191 , n44192 , n44193 , n44194 , n44195 , n44196 , n44197 , 
 n44198 , n44199 , n44200 , n44201 , n44202 , n44203 , n44204 , n44205 , n44206 , n44207 , 
 n44208 , n44209 , n44210 , n44211 , n44212 , n44213 , n44214 , n44215 , n44216 , n44217 , 
 n44218 , n44219 , n44220 , n44221 , n44222 , n44223 , n44224 , n44225 , n44226 , n44227 , 
 n44228 , n44229 , n44230 , n44231 , n44232 , n44233 , n44234 , n44235 , n44236 , n44237 , 
 n44238 , n44239 , n44240 , n44241 , n44242 , n44243 , n44244 , n44245 , n44246 , n44247 , 
 n44248 , n44249 , n44250 , n44251 , n44252 , n44253 , n44254 , n44255 , n44256 , n44257 , 
 n44258 , n44259 , n44260 , n44261 , n44262 , n44263 , n44264 , n44265 , n44266 , n44267 , 
 n44268 , n44269 , n44270 , n44271 , n44272 , n44273 , n44274 , n44275 , n44276 , n44277 , 
 n44278 , n44279 , n44280 , n44281 , n44282 , n44283 , n44284 , n44285 , n44286 , n44287 , 
 n44288 , n44289 , n44290 , n44291 , n44292 , n44293 , n44294 , n44295 , n44296 , n44297 , 
 n44298 , n44299 , n44300 , n44301 , n44302 , n44303 , n44304 , n44305 , n44306 , n44307 , 
 n44308 , n44309 , n44310 , n44311 , n44312 , n44313 , n44314 , n44315 , n44316 , n44317 , 
 n44318 , n44319 , n44320 , n44321 , n44322 , n44323 , n44324 , n44325 , n44326 , n44327 , 
 n44328 , n44329 , n44330 , n44331 , n44332 , n44333 , n44334 , n44335 , n44336 , n44337 , 
 n44338 , n44339 , n44340 , n44341 , n44342 , n44343 , n44344 , n44345 , n44346 , n44347 , 
 n44348 , n44349 , n44350 , n44351 , n44352 , n44353 , n44354 , n44355 , n44356 , n44357 , 
 n44358 , n44359 , n44360 , n44361 , n44362 , n44363 , n44364 , n44365 , n44366 , n44367 , 
 n44368 , n44369 , n44370 , n44371 , n44372 , n44373 , n44374 , n44375 , n44376 , n44377 , 
 n44378 , n44379 , n44380 , n44381 , n44382 , n44383 , n44384 , n44385 , n44386 , n44387 , 
 n44388 , n44389 , n44390 , n44391 , n44392 , n44393 , n44394 , n44395 , n44396 , n44397 , 
 n44398 , n44399 , n44400 , n44401 , n44402 , n44403 , n44404 , n44405 , n44406 , n44407 , 
 n44408 , n44409 , n44410 , n44411 , n44412 , n44413 , n44414 , n44415 , n44416 , n44417 , 
 n44418 , n44419 , n44420 , n44421 , n44422 , n44423 , n44424 , n44425 , n44426 , n44427 , 
 n44428 , n44429 , n44430 , n44431 , n44432 , n44433 , n44434 , n44435 , n44436 , n44437 , 
 n44438 , n44439 , n44440 , n44441 , n44442 , n44443 , n44444 , n44445 , n44446 , n44447 , 
 n44448 , n44449 , n44450 , n44451 , n44452 , n44453 , n44454 , n44455 , n44456 , n44457 , 
 n44458 , n44459 , n44460 , n44461 , n44462 , n44463 , n44464 , n44465 , n44466 , n44467 , 
 n44468 , n44469 , n44470 , n44471 , n44472 , n44473 , n44474 , n44475 , n44476 , n44477 , 
 n44478 , n44479 , n44480 , n44481 , n44482 , n44483 , n44484 , n44485 , n44486 , n44487 , 
 n44488 , n44489 , n44490 , n44491 , n44492 , n44493 , n44494 , n44495 , n44496 , n44497 , 
 n44498 , n44499 , n44500 , n44501 , n44502 , n44503 , n44504 , n44505 , n44506 , n44507 , 
 n44508 , n44509 , n44510 , n44511 , n44512 , n44513 , n44514 , n44515 , n44516 , n44517 , 
 n44518 , n44519 , n44520 , n44521 , n44522 , n44523 , n44524 , n44525 , n44526 , n44527 , 
 n44528 , n44529 , n44530 , n44531 , n44532 , n44533 , n44534 , n44535 , n44536 , n44537 , 
 n44538 , n44539 , n44540 , n44541 , n44542 , n44543 , n44544 , n44545 , n44546 , n44547 , 
 n44548 , n44549 , n44550 , n44551 , n44552 , n44553 , n44554 , n44555 , n44556 , n44557 , 
 n44558 , n44559 , n44560 , n44561 , n44562 , n44563 , n44564 , n44565 , n44566 , n44567 , 
 n44568 , n44569 , n44570 , n44571 , n44572 , n44573 , n44574 , n44575 , n44576 , n44577 , 
 n44578 , n44579 , n44580 , n44581 , n44582 , n44583 , n44584 , n44585 , n44586 , n44587 , 
 n44588 , n44589 , n44590 , n44591 , n44592 , n44593 , n44594 , n44595 , n44596 , n44597 , 
 n44598 , n44599 , n44600 , n44601 , n44602 , n44603 , n44604 , n44605 , n44606 , n44607 , 
 n44608 , n44609 , n44610 , n44611 , n44612 , n44613 , n44614 , n44615 , n44616 , n44617 , 
 n44618 , n44619 , n44620 , n44621 , n44622 , n44623 , n44624 , n44625 , n44626 , n44627 , 
 n44628 , n44629 , n44630 , n44631 , n44632 , n44633 , n44634 , n44635 , n44636 , n44637 , 
 n44638 , n44639 , n44640 , n44641 , n44642 , n44643 , n44644 , n44645 , n44646 , n44647 , 
 n44648 , n44649 , n44650 , n44651 , n44652 , n44653 , n44654 , n44655 , n44656 , n44657 , 
 n44658 , n44659 , n44660 , n44661 , n44662 , n44663 , n44664 , n44665 , n44666 , n44667 , 
 n44668 , n44669 , n44670 , n44671 , n44672 , n44673 , n44674 , n44675 , n44676 , n44677 , 
 n44678 , n44679 , n44680 , n44681 , n44682 , n44683 , n44684 , n44685 , n44686 , n44687 , 
 n44688 , n44689 , n44690 , n44691 , n44692 , n44693 , n44694 , n44695 , n44696 , n44697 , 
 n44698 , n44699 , n44700 , n44701 , n44702 , n44703 , n44704 , n44705 , n44706 , n44707 , 
 n44708 , n44709 , n44710 , n44711 , n44712 , n44713 , n44714 , n44715 , n44716 , n44717 , 
 n44718 , n44719 , n44720 , n44721 , n44722 , n44723 , n44724 , n44725 , n44726 , n44727 , 
 n44728 , n44729 , n44730 , n44731 , n44732 , n44733 , n44734 , n44735 , n44736 , n44737 , 
 n44738 , n44739 , n44740 , n44741 , n44742 , n44743 , n44744 , n44745 , n44746 , n44747 , 
 n44748 , n44749 , n44750 , n44751 , n44752 , n44753 , n44754 , n44755 , n44756 , n44757 , 
 n44758 , n44759 , n44760 , n44761 , n44762 , n44763 , n44764 , n44765 , n44766 , n44767 , 
 n44768 , n44769 , n44770 , n44771 , n44772 , n44773 , n44774 , n44775 , n44776 , n44777 , 
 n44778 , n44779 , n44780 , n44781 , n44782 , n44783 , n44784 , n44785 , n44786 , n44787 , 
 n44788 , n44789 , n44790 , n44791 , n44792 , n44793 , n44794 , n44795 , n44796 , n44797 , 
 n44798 , n44799 , n44800 , n44801 , n44802 , n44803 , n44804 , n44805 , n44806 , n44807 , 
 n44808 , n44809 , n44810 , n44811 , n44812 , n44813 , n44814 , n44815 , n44816 , n44817 , 
 n44818 , n44819 , n44820 , n44821 , n44822 , n44823 , n44824 , n44825 , n44826 , n44827 , 
 n44828 , n44829 , n44830 , n44831 , n44832 , n44833 , n44834 , n44835 , n44836 , n44837 , 
 n44838 , n44839 , n44840 , n44841 , n44842 , n44843 , n44844 , n44845 , n44846 , n44847 , 
 n44848 , n44849 , n44850 , n44851 , n44852 , n44853 , n44854 , n44855 , n44856 , n44857 , 
 n44858 , n44859 , n44860 , n44861 , n44862 , n44863 , n44864 , n44865 , n44866 , n44867 , 
 n44868 , n44869 , n44870 , n44871 , n44872 , n44873 , n44874 , n44875 , n44876 , n44877 , 
 n44878 , n44879 , n44880 , n44881 , n44882 , n44883 , n44884 , n44885 , n44886 , n44887 , 
 n44888 , n44889 , n44890 , n44891 , n44892 , n44893 , n44894 , n44895 , n44896 , n44897 , 
 n44898 , n44899 , n44900 , n44901 , n44902 , n44903 , n44904 , n44905 , n44906 , n44907 , 
 n44908 , n44909 , n44910 , n44911 , n44912 , n44913 , n44914 , n44915 , n44916 , n44917 , 
 n44918 , n44919 , n44920 , n44921 , n44922 , n44923 , n44924 , n44925 , n44926 , n44927 , 
 n44928 , n44929 , n44930 , n44931 , n44932 , n44933 , n44934 , n44935 , n44936 , n44937 , 
 n44938 , n44939 , n44940 , n44941 , n44942 , n44943 , n44944 , n44945 , n44946 , n44947 , 
 n44948 , n44949 , n44950 , n44951 , n44952 , n44953 , n44954 , n44955 , n44956 , n44957 , 
 n44958 , n44959 , n44960 , n44961 , n44962 , n44963 , n44964 , n44965 , n44966 , n44967 , 
 n44968 , n44969 , n44970 , n44971 , n44972 , n44973 , n44974 , n44975 , n44976 , n44977 , 
 n44978 , n44979 , n44980 , n44981 , n44982 , n44983 , n44984 , n44985 , n44986 , n44987 , 
 n44988 , n44989 , n44990 , n44991 , n44992 , n44993 , n44994 , n44995 , n44996 , n44997 , 
 n44998 , n44999 , n45000 , n45001 , n45002 , n45003 , n45004 , n45005 , n45006 , n45007 , 
 n45008 , n45009 , n45010 , n45011 , n45012 , n45013 , n45014 , n45015 , n45016 , n45017 , 
 n45018 , n45019 , n45020 , n45021 , n45022 , n45023 , n45024 , n45025 , n45026 , n45027 , 
 n45028 , n45029 , n45030 , n45031 , n45032 , n45033 , n45034 , n45035 , n45036 , n45037 , 
 n45038 , n45039 , n45040 , n45041 , n45042 , n45043 , n45044 , n45045 , n45046 , n45047 , 
 n45048 , n45049 , n45050 , n45051 , n45052 , n45053 , n45054 , n45055 , n45056 , n45057 , 
 n45058 , n45059 , n45060 , n45061 , n45062 , n45063 , n45064 , n45065 , n45066 , n45067 , 
 n45068 , n45069 , n45070 , n45071 , n45072 , n45073 , n45074 , n45075 , n45076 , n45077 , 
 n45078 , n45079 , n45080 , n45081 , n45082 , n45083 , n45084 , n45085 , n45086 , n45087 , 
 n45088 , n45089 , n45090 , n45091 , n45092 , n45093 , n45094 , n45095 , n45096 , n45097 , 
 n45098 , n45099 , n45100 , n45101 , n45102 , n45103 , n45104 , n45105 , n45106 , n45107 , 
 n45108 , n45109 , n45110 , n45111 , n45112 , n45113 , n45114 , n45115 , n45116 , n45117 , 
 n45118 , n45119 , n45120 , n45121 , n45122 , n45123 , n45124 , n45125 , n45126 , n45127 , 
 n45128 , n45129 , n45130 , n45131 , n45132 , n45133 , n45134 , n45135 , n45136 , n45137 , 
 n45138 , n45139 , n45140 , n45141 , n45142 , n45143 , n45144 , n45145 , n45146 , n45147 , 
 n45148 , n45149 , n45150 , n45151 , n45152 , n45153 , n45154 , n45155 , n45156 , n45157 , 
 n45158 , n45159 , n45160 , n45161 , n45162 , n45163 , n45164 , n45165 , n45166 , n45167 , 
 n45168 , n45169 , n45170 , n45171 , n45172 , n45173 , n45174 , n45175 , n45176 , n45177 , 
 n45178 , n45179 , n45180 , n45181 , n45182 , n45183 , n45184 , n45185 , n45186 , n45187 , 
 n45188 , n45189 , n45190 , n45191 , n45192 , n45193 , n45194 , n45195 , n45196 , n45197 , 
 n45198 , n45199 , n45200 , n45201 , n45202 , n45203 , n45204 , n45205 , n45206 , n45207 , 
 n45208 , n45209 , n45210 , n45211 , n45212 , n45213 , n45214 , n45215 , n45216 , n45217 , 
 n45218 , n45219 , n45220 , n45221 , n45222 , n45223 , n45224 , n45225 , n45226 , n45227 , 
 n45228 , n45229 , n45230 , n45231 , n45232 , n45233 , n45234 , n45235 , n45236 , n45237 , 
 n45238 , n45239 , n45240 , n45241 , n45242 , n45243 , n45244 , n45245 , n45246 , n45247 , 
 n45248 , n45249 , n45250 , n45251 , n45252 , n45253 , n45254 , n45255 , n45256 , n45257 , 
 n45258 , n45259 , n45260 , n45261 , n45262 , n45263 , n45264 , n45265 , n45266 , n45267 , 
 n45268 , n45269 , n45270 , n45271 , n45272 , n45273 , n45274 , n45275 , n45276 , n45277 , 
 n45278 , n45279 , n45280 , n45281 , n45282 , n45283 , n45284 , n45285 , n45286 , n45287 , 
 n45288 , n45289 , n45290 , n45291 , n45292 , n45293 , n45294 , n45295 , n45296 , n45297 , 
 n45298 , n45299 , n45300 , n45301 , n45302 , n45303 , n45304 , n45305 , n45306 , n45307 , 
 n45308 , n45309 , n45310 , n45311 , n45312 , n45313 , n45314 , n45315 , n45316 , n45317 , 
 n45318 , n45319 , n45320 , n45321 , n45322 , n45323 , n45324 , n45325 , n45326 , n45327 , 
 n45328 , n45329 , n45330 , n45331 , n45332 , n45333 , n45334 , n45335 , n45336 , n45337 , 
 n45338 , n45339 , n45340 , n45341 , n45342 , n45343 , n45344 , n45345 , n45346 , n45347 , 
 n45348 , n45349 , n45350 , n45351 , n45352 , n45353 , n45354 , n45355 , n45356 , n45357 , 
 n45358 , n45359 , n45360 , n45361 , n45362 , n45363 , n45364 , n45365 , n45366 , n45367 , 
 n45368 , n45369 , n45370 , n45371 , n45372 , n45373 , n45374 , n45375 , n45376 , n45377 , 
 n45378 , n45379 , n45380 , n45381 , n45382 , n45383 , n45384 , n45385 , n45386 , n45387 , 
 n45388 , n45389 , n45390 , n45391 , n45392 , n45393 , n45394 , n45395 , n45396 , n45397 , 
 n45398 , n45399 , n45400 , n45401 , n45402 , n45403 , n45404 , n45405 , n45406 , n45407 , 
 n45408 , n45409 , n45410 , n45411 , n45412 , n45413 , n45414 , n45415 , n45416 , n45417 , 
 n45418 , n45419 , n45420 , n45421 , n45422 , n45423 , n45424 , n45425 , n45426 , n45427 , 
 n45428 , n45429 , n45430 , n45431 , n45432 , n45433 , n45434 , n45435 , n45436 , n45437 , 
 n45438 , n45439 , n45440 , n45441 , n45442 , n45443 , n45444 , n45445 , n45446 , n45447 , 
 n45448 , n45449 , n45450 , n45451 , n45452 , n45453 , n45454 , n45455 , n45456 , n45457 , 
 n45458 , n45459 , n45460 , n45461 , n45462 , n45463 , n45464 , n45465 , n45466 , n45467 , 
 n45468 , n45469 , n45470 , n45471 , n45472 , n45473 , n45474 , n45475 , n45476 , n45477 , 
 n45478 , n45479 , n45480 , n45481 , n45482 , n45483 , n45484 , n45485 , n45486 , n45487 , 
 n45488 , n45489 , n45490 , n45491 , n45492 , n45493 , n45494 , n45495 , n45496 , n45497 , 
 n45498 , n45499 , n45500 , n45501 , n45502 , n45503 , n45504 , n45505 , n45506 , n45507 , 
 n45508 , n45509 , n45510 , n45511 , n45512 , n45513 , n45514 , n45515 , n45516 , n45517 , 
 n45518 , n45519 , n45520 , n45521 , n45522 , n45523 , n45524 , n45525 , n45526 , n45527 , 
 n45528 , n45529 , n45530 , n45531 , n45532 , n45533 , n45534 , n45535 , n45536 , n45537 , 
 n45538 , n45539 , n45540 , n45541 , n45542 , n45543 , n45544 , n45545 , n45546 , n45547 , 
 n45548 , n45549 , n45550 , n45551 , n45552 , n45553 , n45554 , n45555 , n45556 , n45557 , 
 n45558 , n45559 , n45560 , n45561 , n45562 , n45563 , n45564 , n45565 , n45566 , n45567 , 
 n45568 , n45569 , n45570 , n45571 , n45572 , n45573 , n45574 , n45575 , n45576 , n45577 , 
 n45578 , n45579 , n45580 , n45581 , n45582 , n45583 , n45584 , n45585 , n45586 , n45587 , 
 n45588 , n45589 , n45590 , n45591 , n45592 , n45593 , n45594 , n45595 , n45596 , n45597 , 
 n45598 , n45599 , n45600 , n45601 , n45602 , n45603 , n45604 , n45605 , n45606 , n45607 , 
 n45608 , n45609 , n45610 , n45611 , n45612 , n45613 , n45614 , n45615 , n45616 , n45617 , 
 n45618 , n45619 , n45620 , n45621 , n45622 , n45623 , n45624 , n45625 , n45626 , n45627 , 
 n45628 , n45629 , n45630 , n45631 , n45632 , n45633 , n45634 , n45635 , n45636 , n45637 , 
 n45638 , n45639 , n45640 , n45641 , n45642 , n45643 , n45644 , n45645 , n45646 , n45647 , 
 n45648 , n45649 , n45650 , n45651 , n45652 , n45653 , n45654 , n45655 , n45656 , n45657 , 
 n45658 , n45659 , n45660 , n45661 , n45662 , n45663 , n45664 , n45665 , n45666 , n45667 , 
 n45668 , n45669 , n45670 , n45671 , n45672 , n45673 , n45674 , n45675 , n45676 , n45677 , 
 n45678 , n45679 , n45680 , n45681 , n45682 , n45683 , n45684 , n45685 , n45686 , n45687 , 
 n45688 , n45689 , n45690 , n45691 , n45692 , n45693 , n45694 , n45695 , n45696 , n45697 , 
 n45698 , n45699 , n45700 , n45701 , n45702 , n45703 , n45704 , n45705 , n45706 , n45707 , 
 n45708 , n45709 , n45710 , n45711 , n45712 , n45713 , n45714 , n45715 , n45716 , n45717 , 
 n45718 , n45719 , n45720 , n45721 , n45722 , n45723 , n45724 , n45725 , n45726 , n45727 , 
 n45728 , n45729 , n45730 , n45731 , n45732 , n45733 , n45734 , n45735 , n45736 , n45737 , 
 n45738 , n45739 , n45740 , n45741 , n45742 , n45743 , n45744 , n45745 , n45746 , n45747 , 
 n45748 , n45749 , n45750 , n45751 , n45752 , n45753 , n45754 , n45755 , n45756 , n45757 , 
 n45758 , n45759 , n45760 , n45761 , n45762 , n45763 , n45764 , n45765 , n45766 , n45767 , 
 n45768 , n45769 , n45770 , n45771 , n45772 , n45773 , n45774 , n45775 , n45776 , n45777 , 
 n45778 , n45779 , n45780 , n45781 , n45782 , n45783 , n45784 , n45785 , n45786 , n45787 , 
 n45788 , n45789 , n45790 , n45791 , n45792 , n45793 , n45794 , n45795 , n45796 , n45797 , 
 n45798 , n45799 , n45800 , n45801 , n45802 , n45803 , n45804 , n45805 , n45806 , n45807 , 
 n45808 , n45809 , n45810 , n45811 , n45812 , n45813 , n45814 , n45815 , n45816 , n45817 , 
 n45818 , n45819 , n45820 , n45821 , n45822 , n45823 , n45824 , n45825 , n45826 , n45827 , 
 n45828 , n45829 , n45830 , n45831 , n45832 , n45833 , n45834 , n45835 , n45836 , n45837 , 
 n45838 , n45839 , n45840 , n45841 , n45842 , n45843 , n45844 , n45845 , n45846 , n45847 , 
 n45848 , n45849 , n45850 , n45851 , n45852 , n45853 , n45854 , n45855 , n45856 , n45857 , 
 n45858 , n45859 , n45860 , n45861 , n45862 , n45863 , n45864 , n45865 , n45866 , n45867 , 
 n45868 , n45869 , n45870 , n45871 , n45872 , n45873 , n45874 , n45875 , n45876 , n45877 , 
 n45878 , n45879 , n45880 , n45881 , n45882 , n45883 , n45884 , n45885 , n45886 , n45887 , 
 n45888 , n45889 , n45890 , n45891 , n45892 , n45893 , n45894 , n45895 , n45896 , n45897 , 
 n45898 , n45899 , n45900 , n45901 , n45902 , n45903 , n45904 , n45905 , n45906 , n45907 , 
 n45908 , n45909 , n45910 , n45911 , n45912 , n45913 , n45914 , n45915 , n45916 , n45917 , 
 n45918 , n45919 , n45920 , n45921 , n45922 , n45923 , n45924 , n45925 , n45926 , n45927 , 
 n45928 , n45929 , n45930 , n45931 , n45932 , n45933 , n45934 , n45935 , n45936 , n45937 , 
 n45938 , n45939 , n45940 , n45941 , n45942 , n45943 , n45944 , n45945 , n45946 , n45947 , 
 n45948 , n45949 , n45950 , n45951 , n45952 , n45953 , n45954 , n45955 , n45956 , n45957 , 
 n45958 , n45959 , n45960 , n45961 , n45962 , n45963 , n45964 , n45965 , n45966 , n45967 , 
 n45968 , n45969 , n45970 , n45971 , n45972 , n45973 , n45974 , n45975 , n45976 , n45977 , 
 n45978 , n45979 , n45980 , n45981 , n45982 , n45983 , n45984 , n45985 , n45986 , n45987 , 
 n45988 , n45989 , n45990 , n45991 , n45992 , n45993 , n45994 , n45995 , n45996 , n45997 , 
 n45998 , n45999 , n46000 , n46001 , n46002 , n46003 , n46004 , n46005 , n46006 , n46007 , 
 n46008 , n46009 , n46010 , n46011 , n46012 , n46013 , n46014 , n46015 , n46016 , n46017 , 
 n46018 , n46019 , n46020 , n46021 , n46022 , n46023 , n46024 , n46025 , n46026 , n46027 , 
 n46028 , n46029 , n46030 , n46031 , n46032 , n46033 , n46034 , n46035 , n46036 , n46037 , 
 n46038 , n46039 , n46040 , n46041 , n46042 , n46043 , n46044 , n46045 , n46046 , n46047 , 
 n46048 , n46049 , n46050 , n46051 , n46052 , n46053 , n46054 , n46055 , n46056 , n46057 , 
 n46058 , n46059 , n46060 , n46061 , n46062 , n46063 , n46064 , n46065 , n46066 , n46067 , 
 n46068 , n46069 , n46070 , n46071 , n46072 , n46073 , n46074 , n46075 , n46076 , n46077 , 
 n46078 , n46079 , n46080 , n46081 , n46082 , n46083 , n46084 , n46085 , n46086 , n46087 , 
 n46088 , n46089 , n46090 , n46091 , n46092 , n46093 , n46094 , n46095 , n46096 , n46097 , 
 n46098 , n46099 , n46100 , n46101 , n46102 , n46103 , n46104 , n46105 , n46106 , n46107 , 
 n46108 , n46109 , n46110 , n46111 , n46112 , n46113 , n46114 , n46115 , n46116 , n46117 , 
 n46118 , n46119 , n46120 , n46121 , n46122 , n46123 , n46124 , n46125 , n46126 , n46127 , 
 n46128 , n46129 , n46130 , n46131 , n46132 , n46133 , n46134 , n46135 , n46136 , n46137 , 
 n46138 , n46139 , n46140 , n46141 , n46142 , n46143 , n46144 , n46145 , n46146 , n46147 , 
 n46148 , n46149 , n46150 , n46151 , n46152 , n46153 , n46154 , n46155 , n46156 , n46157 , 
 n46158 , n46159 , n46160 , n46161 , n46162 , n46163 , n46164 , n46165 , n46166 , n46167 , 
 n46168 , n46169 , n46170 , n46171 , n46172 , n46173 , n46174 , n46175 , n46176 , n46177 , 
 n46178 , n46179 , n46180 , n46181 , n46182 , n46183 , n46184 , n46185 , n46186 , n46187 , 
 n46188 , n46189 , n46190 , n46191 , n46192 , n46193 , n46194 , n46195 , n46196 , n46197 , 
 n46198 , n46199 , n46200 , n46201 , n46202 , n46203 , n46204 , n46205 , n46206 , n46207 , 
 n46208 , n46209 , n46210 , n46211 , n46212 , n46213 , n46214 , n46215 , n46216 , n46217 , 
 n46218 , n46219 , n46220 , n46221 , n46222 , n46223 , n46224 , n46225 , n46226 , n46227 , 
 n46228 , n46229 , n46230 , n46231 , n46232 , n46233 , n46234 , n46235 , n46236 , n46237 , 
 n46238 , n46239 , n46240 , n46241 , n46242 , n46243 , n46244 , n46245 , n46246 , n46247 , 
 n46248 , n46249 , n46250 , n46251 , n46252 , n46253 , n46254 , n46255 , n46256 , n46257 , 
 n46258 , n46259 , n46260 , n46261 , n46262 , n46263 , n46264 , n46265 , n46266 , n46267 , 
 n46268 , n46269 , n46270 , n46271 , n46272 , n46273 , n46274 , n46275 , n46276 , n46277 , 
 n46278 , n46279 , n46280 , n46281 , n46282 , n46283 , n46284 , n46285 , n46286 , n46287 , 
 n46288 , n46289 , n46290 , n46291 , n46292 , n46293 , n46294 , n46295 , n46296 , n46297 , 
 n46298 , n46299 , n46300 , n46301 , n46302 , n46303 , n46304 , n46305 , n46306 , n46307 , 
 n46308 , n46309 , n46310 , n46311 , n46312 , n46313 , n46314 , n46315 , n46316 , n46317 , 
 n46318 , n46319 , n46320 , n46321 , n46322 , n46323 , n46324 , n46325 , n46326 , n46327 , 
 n46328 , n46329 , n46330 , n46331 , n46332 , n46333 , n46334 , n46335 , n46336 , n46337 , 
 n46338 , n46339 , n46340 , n46341 , n46342 , n46343 , n46344 , n46345 , n46346 , n46347 , 
 n46348 , n46349 , n46350 , n46351 , n46352 , n46353 , n46354 , n46355 , n46356 , n46357 , 
 n46358 , n46359 , n46360 , n46361 , n46362 , n46363 , n46364 , n46365 , n46366 , n46367 , 
 n46368 , n556 , n557 , n46371 , n46372 , n46373 , n46374 , n562 , n46376 , n564 , 
 n565 , n566 , n567 , n568 , n46382 , n46383 , n46384 , n572 , n46386 , n46387 , 
 n575 , n46389 , n46390 , n578 , n46392 , n46393 , n581 , n46395 , n46396 , n46397 , 
 n46398 , n46399 , n587 , n46401 , n589 , n590 , n591 , n46405 , n593 , n594 , 
 n595 , n596 , n46410 , n598 , n599 , n46413 , n601 , n602 , n603 , n604 , 
 n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , 
 n615 , n616 , n617 , n618 , n619 , n620 , n46434 , n46435 , n623 , n46437 , 
 n46438 , n626 , n46440 , n46441 , n46442 , n630 , n46444 , n632 , n633 , n634 , 
 n635 , n636 , n637 , n638 , n639 , n640 , n641 , n46455 , n46456 , n644 , 
 n46458 , n46459 , n647 , n46461 , n46462 , n650 , n46464 , n46465 , n653 , n654 , 
 n655 , n656 , n657 , n46471 , n659 , n46473 , n46474 , n662 , n46476 , n664 , 
 n665 , n666 , n667 , n668 , n669 , n670 , n671 , n46485 , n673 , n674 , 
 n675 , n676 , n677 , n678 , n679 , n680 , n46494 , n46495 , n46496 , n46497 , 
 n46498 , n46499 , n46500 , n46501 , n46502 , n690 , n691 , n692 , n693 , n694 , 
 n695 , n696 , n46510 , n698 , n46512 , n700 , n701 , n46515 , n46516 , n704 , 
 n46518 , n706 , n46520 , n46521 , n709 , n46523 , n46524 , n712 , n46526 , n46527 , 
 n715 , n46529 , n717 , n46531 , n719 , n46533 , n46534 , n722 , n723 , n46537 , 
 n725 , n726 , n727 , n728 , n729 , n46543 , n46544 , n732 , n46546 , n46547 , 
 n735 , n46549 , n737 , n46551 , n46552 , n46553 , n46554 , n742 , n46556 , n46557 , 
 n745 , n46559 , n747 , n46561 , n749 , n46563 , n46564 , n752 , n46566 , n754 , 
 n755 , n756 , n757 , n758 , n46572 , n760 , n46574 , n46575 , n763 , n46577 , 
 n46578 , n766 , n46580 , n46581 , n769 , n46583 , n771 , n772 , n773 , n774 , 
 n775 , n776 , n46590 , n46591 , n779 , n46593 , n781 , n782 , n783 , n784 , 
 n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n46607 , 
 n795 , n46609 , n46610 , n798 , n799 , n800 , n46614 , n802 , n803 , n46617 , 
 n805 , n46619 , n807 , n808 , n809 , n810 , n811 , n46625 , n813 , n46627 , 
 n815 , n816 , n817 , n46631 , n46632 , n820 , n46634 , n46635 , n823 , n46637 , 
 n46638 , n826 , n46640 , n46641 , n829 , n46643 , n46644 , n832 , n46646 , n834 , 
 n835 , n836 , n837 , n46651 , n839 , n46653 , n46654 , n842 , n46656 , n46657 , 
 n845 , n846 , n46660 , n848 , n46662 , n850 , n46664 , n46665 , n853 , n46667 , 
 n46668 , n856 , n857 , n46671 , n859 , n860 , n861 , n862 , n863 , n864 , 
 n865 , n46679 , n46680 , n868 , n46682 , n870 , n871 , n872 , n873 , n874 , 
 n875 , n46689 , n877 , n46691 , n879 , n880 , n881 , n882 , n46696 , n884 , 
 n885 , n46699 , n887 , n888 , n46702 , n890 , n891 , n46705 , n893 , n46707 , 
 n46708 , n896 , n897 , n46711 , n46712 , n46713 , n901 , n46715 , n46716 , n904 , 
 n46718 , n46719 , n907 , n46721 , n46722 , n910 , n911 , n912 , n913 , n914 , 
 n46728 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , 
 n925 , n46739 , n927 , n46741 , n46742 , n930 , n46744 , n46745 , n933 , n46747 , 
 n46748 , n936 , n937 , n46751 , n46752 , n940 , n46754 , n46755 , n943 , n944 , 
 n46758 , n46759 , n947 , n46761 , n46762 , n46763 , n951 , n46765 , n953 , n954 , 
 n955 , n46769 , n957 , n958 , n46772 , n960 , n46774 , n46775 , n46776 , n964 , 
 n46778 , n46779 , n46780 , n968 , n46782 , n46783 , n971 , n46785 , n46786 , n974 , 
 n975 , n976 , n46790 , n46791 , n46792 , n46793 , n981 , n46795 , n46796 , n46797 , 
 n985 , n46799 , n987 , n988 , n989 , n990 , n991 , n46805 , n993 , n46807 , 
 n46808 , n46809 , n997 , n46811 , n999 , n46813 , n46814 , n1002 , n46816 , n46817 , 
 n1005 , n46819 , n1007 , n1008 , n46822 , n1010 , n46824 , n1012 , n1013 , n1014 , 
 n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n46835 , n1023 , n46837 , 
 n1025 , n46839 , n1027 , n46841 , n46842 , n1030 , n46844 , n46845 , n1033 , n46847 , 
 n46848 , n1036 , n46850 , n46851 , n46852 , n46853 , n1041 , n46855 , n46856 , n1044 , 
 n46858 , n46859 , n1047 , n1048 , n1049 , n1050 , n46864 , n46865 , n1053 , n46867 , 
 n46868 , n46869 , n46870 , n1058 , n46872 , n46873 , n1061 , n46875 , n46876 , n1064 , 
 n46878 , n46879 , n1067 , n46881 , n1069 , n46883 , n46884 , n1072 , n1073 , n1074 , 
 n46888 , n46889 , n46890 , n1078 , n1079 , n46893 , n46894 , n1082 , n46896 , n1084 , 
 n1085 , n1086 , n1087 , n46901 , n1089 , n46903 , n1091 , n46905 , n1093 , n1094 , 
 n46908 , n1096 , n1097 , n46911 , n46912 , n1100 , n1101 , n46915 , n46916 , n1104 , 
 n46918 , n1106 , n46920 , n46921 , n1109 , n46923 , n46924 , n1112 , n46926 , n1114 , 
 n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , 
 n1125 , n46939 , n46940 , n1128 , n46942 , n46943 , n1131 , n46945 , n1133 , n46947 , 
 n1135 , n1136 , n1137 , n1138 , n1139 , n46953 , n1141 , n46955 , n46956 , n1144 , 
 n1145 , n1146 , n46960 , n1148 , n1149 , n1150 , n46964 , n1152 , n46966 , n1154 , 
 n46968 , n46969 , n1157 , n46971 , n1159 , n1160 , n1161 , n46975 , n1163 , n1164 , 
 n1165 , n1166 , n46980 , n1168 , n46982 , n1170 , n1171 , n1172 , n1173 , n1174 , 
 n1175 , n1176 , n46990 , n1178 , n46992 , n46993 , n1181 , n1182 , n46996 , n46997 , 
 n46998 , n46999 , n1187 , n47001 , n47002 , n1190 , n1191 , n47005 , n1193 , n47007 , 
 n47008 , n47009 , n1197 , n47011 , n47012 , n47013 , n1201 , n1202 , n47016 , n1204 , 
 n47018 , n47019 , n1207 , n47021 , n47022 , n1210 , n1211 , n1212 , n1213 , n1214 , 
 n1215 , n1216 , n47030 , n47031 , n1219 , n47033 , n1221 , n47035 , n47036 , n47037 , 
 n47038 , n1226 , n1227 , n47041 , n47042 , n1230 , n1231 , n47045 , n47046 , n1234 , 
 n47048 , n47049 , n1237 , n47051 , n47052 , n1240 , n47054 , n1242 , n1243 , n47057 , 
 n1245 , n47059 , n47060 , n47061 , n1249 , n47063 , n47064 , n1252 , n47066 , n1254 , 
 n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , 
 n1265 , n1266 , n1267 , n47081 , n1269 , n1270 , n1271 , n1272 , n1273 , n47087 , 
 n47088 , n1276 , n47090 , n47091 , n47092 , n47093 , n1281 , n47095 , n1283 , n1284 , 
 n1285 , n1286 , n1287 , n47101 , n47102 , n1290 , n1291 , n1292 , n47106 , n47107 , 
 n1295 , n47109 , n1297 , n47111 , n1299 , n47113 , n1301 , n1302 , n47116 , n47117 , 
 n1305 , n47119 , n1307 , n47121 , n47122 , n1310 , n47124 , n1312 , n47126 , n47127 , 
 n47128 , n1316 , n47130 , n47131 , n1319 , n1320 , n47134 , n1322 , n47136 , n47137 , 
 n47138 , n1326 , n47140 , n1328 , n1329 , n47143 , n47144 , n1332 , n47146 , n47147 , 
 n1335 , n47149 , n1337 , n1338 , n47152 , n1340 , n47154 , n1342 , n1343 , n1344 , 
 n1345 , n47159 , n47160 , n1348 , n47162 , n47163 , n1351 , n47165 , n47166 , n1354 , 
 n1355 , n47169 , n47170 , n1358 , n47172 , n1360 , n47174 , n1362 , n1363 , n47177 , 
 n1365 , n47179 , n1367 , n1368 , n47182 , n47183 , n1371 , n47185 , n47186 , n1374 , 
 n47188 , n47189 , n47190 , n1378 , n47192 , n47193 , n1381 , n47195 , n47196 , n1384 , 
 n1385 , n1386 , n47200 , n1388 , n1389 , n47203 , n1391 , n47205 , n47206 , n1394 , 
 n47208 , n47209 , n1397 , n1398 , n1399 , n47213 , n47214 , n1402 , n47216 , n1404 , 
 n1405 , n47219 , n1407 , n47221 , n1409 , n1410 , n1411 , n1412 , n47226 , n47227 , 
 n47228 , n47229 , n47230 , n1418 , n47232 , n47233 , n1421 , n47235 , n1423 , n47237 , 
 n1425 , n1426 , n47240 , n1428 , n47242 , n1430 , n1431 , n1432 , n47246 , n1434 , 
 n47248 , n47249 , n47250 , n1438 , n47252 , n47253 , n1441 , n47255 , n47256 , n1444 , 
 n1445 , n1446 , n47260 , n47261 , n47262 , n47263 , n1451 , n47265 , n1453 , n1454 , 
 n47268 , n47269 , n1457 , n1458 , n47272 , n1460 , n47274 , n47275 , n1463 , n1464 , 
 n47278 , n47279 , n47280 , n1468 , n47282 , n47283 , n1471 , n47285 , n47286 , n1474 , 
 n47288 , n47289 , n1477 , n47291 , n47292 , n1480 , n47294 , n47295 , n47296 , n47297 , 
 n1485 , n1486 , n47300 , n1488 , n47302 , n1490 , n47304 , n47305 , n1493 , n47307 , 
 n47308 , n1496 , n47310 , n47311 , n1499 , n47313 , n1501 , n47315 , n47316 , n1504 , 
 n47318 , n47319 , n47320 , n1508 , n47322 , n1510 , n47324 , n1512 , n1513 , n47327 , 
 n47328 , n1516 , n47330 , n47331 , n1519 , n47333 , n47334 , n1522 , n1523 , n47337 , 
 n47338 , n1526 , n1527 , n47341 , n1529 , n1530 , n47344 , n47345 , n47346 , n1534 , 
 n47348 , n47349 , n1537 , n47351 , n47352 , n1540 , n1541 , n1542 , n1543 , n1544 , 
 n1545 , n47359 , n47360 , n47361 , n47362 , n1550 , n47364 , n47365 , n47366 , n1554 , 
 n47368 , n47369 , n1557 , n1558 , n47372 , n47373 , n1561 , n1562 , n47376 , n47377 , 
 n1565 , n1566 , n47380 , n1568 , n47382 , n47383 , n1571 , n47385 , n1573 , n1574 , 
 n1575 , n1576 , n47390 , n47391 , n47392 , n47393 , n47394 , n47395 , n1583 , n1584 , 
 n47398 , n47399 , n1587 , n47401 , n1589 , n47403 , n47404 , n1592 , n47406 , n47407 , 
 n1595 , n1596 , n47410 , n47411 , n1599 , n47413 , n1601 , n47415 , n47416 , n47417 , 
 n47418 , n1606 , n47420 , n47421 , n47422 , n1610 , n47424 , n47425 , n47426 , n47427 , 
 n47428 , n1616 , n1617 , n47431 , n1619 , n1620 , n1621 , n47435 , n1623 , n47437 , 
 n1625 , n1626 , n47440 , n47441 , n1629 , n47443 , n1631 , n47445 , n47446 , n1634 , 
 n47448 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , 
 n1645 , n47459 , n47460 , n47461 , n47462 , n1650 , n47464 , n47465 , n1653 , n47467 , 
 n1655 , n47469 , n1657 , n47471 , n1659 , n47473 , n47474 , n1662 , n47476 , n1664 , 
 n1665 , n47479 , n1667 , n47481 , n1669 , n47483 , n47484 , n1672 , n47486 , n47487 , 
 n47488 , n1676 , n47490 , n1678 , n47492 , n47493 , n47494 , n1682 , n47496 , n47497 , 
 n1685 , n47499 , n47500 , n1688 , n1689 , n1690 , n47504 , n47505 , n1693 , n47507 , 
 n1695 , n1696 , n47510 , n1698 , n47512 , n1700 , n1701 , n47515 , n47516 , n1704 , 
 n47518 , n47519 , n1707 , n47521 , n1709 , n1710 , n1711 , n47525 , n47526 , n47527 , 
 n1715 , n47529 , n47530 , n1718 , n47532 , n1720 , n47534 , n1722 , n1723 , n47537 , 
 n47538 , n1726 , n1727 , n47541 , n1729 , n1730 , n47544 , n47545 , n47546 , n1734 , 
 n47548 , n47549 , n1737 , n47551 , n47552 , n1740 , n47554 , n47555 , n1743 , n1744 , 
 n47558 , n47559 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , 
 n1755 , n47569 , n1757 , n47571 , n47572 , n47573 , n1761 , n47575 , n1763 , n47577 , 
 n47578 , n1766 , n47580 , n47581 , n1769 , n47583 , n1771 , n1772 , n1773 , n1774 , 
 n1775 , n1776 , n47590 , n47591 , n47592 , n47593 , n47594 , n1782 , n1783 , n47597 , 
 n47598 , n1786 , n47600 , n1788 , n1789 , n1790 , n47604 , n47605 , n47606 , n1794 , 
 n47608 , n47609 , n1797 , n47611 , n1799 , n47613 , n47614 , n1802 , n47616 , n47617 , 
 n1805 , n47619 , n47620 , n47621 , n1809 , n47623 , n47624 , n47625 , n47626 , n47627 , 
 n1815 , n1816 , n47630 , n47631 , n1819 , n47633 , n47634 , n1822 , n47636 , n1824 , 
 n47638 , n47639 , n1827 , n47641 , n1829 , n47643 , n1831 , n47645 , n1833 , n1834 , 
 n47648 , n47649 , n1837 , n1838 , n47652 , n1840 , n1841 , n47655 , n47656 , n47657 , 
 n47658 , n1846 , n47660 , n47661 , n1849 , n1850 , n47664 , n47665 , n1853 , n1854 , 
 n47668 , n47669 , n1857 , n47671 , n1859 , n47673 , n1861 , n47675 , n47676 , n1864 , 
 n1865 , n1866 , n1867 , n1868 , n47682 , n47683 , n1871 , n47685 , n47686 , n1874 , 
 n47688 , n1876 , n47690 , n47691 , n47692 , n1880 , n47694 , n47695 , n1883 , n47697 , 
 n47698 , n47699 , n1887 , n47701 , n1889 , n47703 , n1891 , n47705 , n1893 , n1894 , 
 n47708 , n47709 , n1897 , n47711 , n47712 , n1900 , n47714 , n47715 , n47716 , n1904 , 
 n47718 , n1906 , n1907 , n47721 , n47722 , n47723 , n47724 , n47725 , n47726 , n1914 , 
 n47728 , n1916 , n1917 , n47731 , n47732 , n1920 , n1921 , n47735 , n47736 , n1924 , 
 n47738 , n47739 , n47740 , n47741 , n47742 , n1930 , n47744 , n47745 , n1933 , n47747 , 
 n47748 , n1936 , n47750 , n47751 , n1939 , n47753 , n47754 , n1942 , n47756 , n47757 , 
 n1945 , n47759 , n1947 , n47761 , n1949 , n47763 , n1951 , n1952 , n1953 , n47767 , 
 n1955 , n47769 , n1957 , n1958 , n47772 , n1960 , n47774 , n47775 , n1963 , n47777 , 
 n47778 , n1966 , n47780 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , 
 n1975 , n47789 , n47790 , n1978 , n47792 , n1980 , n47794 , n1982 , n1983 , n47797 , 
 n1985 , n47799 , n1987 , n47801 , n1989 , n1990 , n47804 , n1992 , n47806 , n1994 , 
 n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n47815 , n2003 , n2004 , 
 n2005 , n2006 , n2007 , n2008 , n47822 , n47823 , n2011 , n2012 , n2013 , n47827 , 
 n2015 , n47829 , n47830 , n2018 , n47832 , n47833 , n2021 , n2022 , n47836 , n2024 , 
 n47838 , n47839 , n2027 , n47841 , n47842 , n2030 , n2031 , n2032 , n47846 , n2034 , 
 n47848 , n2036 , n47850 , n2038 , n2039 , n47853 , n2041 , n47855 , n47856 , n47857 , 
 n2045 , n47859 , n47860 , n2048 , n47862 , n2050 , n47864 , n2052 , n47866 , n47867 , 
 n2055 , n47869 , n2057 , n2058 , n2059 , n2060 , n2061 , n47875 , n47876 , n2064 , 
 n47878 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , 
 n47888 , n47889 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , 
 n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , 
 n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , 
 n2105 , n2106 , n2107 , n47921 , n47922 , n2110 , n2111 , n2112 , n2113 , n2114 , 
 n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , 
 n47938 , n2126 , n47940 , n2128 , n47942 , n47943 , n2131 , n47945 , n2133 , n2134 , 
 n47948 , n47949 , n2137 , n47951 , n47952 , n2140 , n47954 , n47955 , n47956 , n47957 , 
 n2145 , n47959 , n47960 , n47961 , n2149 , n47963 , n2151 , n47965 , n47966 , n2154 , 
 n47968 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , 
 n2165 , n2166 , n47980 , n2168 , n47982 , n2170 , n2171 , n47985 , n47986 , n47987 , 
 n47988 , n47989 , n2177 , n47991 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , 
 n2185 , n2186 , n48000 , n48001 , n2189 , n48003 , n2191 , n2192 , n2193 , n2194 , 
 n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n48017 , 
 n48018 , n2206 , n48020 , n48021 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , 
 n2215 , n2216 , n2217 , n48031 , n48032 , n2220 , n48034 , n48035 , n2223 , n48037 , 
 n48038 , n2226 , n2227 , n2228 , n2229 , n2230 , n48044 , n48045 , n2233 , n48047 , 
 n48048 , n48049 , n48050 , n2238 , n48052 , n48053 , n48054 , n48055 , n48056 , n2244 , 
 n48058 , n2246 , n2247 , n2248 , n2249 , n2250 , n48064 , n2252 , n48066 , n2254 , 
 n48068 , n2256 , n48070 , n48071 , n48072 , n2260 , n48074 , n2262 , n48076 , n48077 , 
 n2265 , n48079 , n48080 , n2268 , n2269 , n48083 , n48084 , n48085 , n48086 , n48087 , 
 n48088 , n2276 , n48090 , n48091 , n2279 , n48093 , n48094 , n2282 , n2283 , n48097 , 
 n48098 , n2286 , n48100 , n48101 , n2289 , n48103 , n48104 , n2292 , n2293 , n48107 , 
 n48108 , n2296 , n48110 , n48111 , n2299 , n48113 , n2301 , n2302 , n2303 , n2304 , 
 n2305 , n48119 , n48120 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , 
 n48128 , n48129 , n2317 , n48131 , n2319 , n48133 , n48134 , n48135 , n48136 , n2324 , 
 n48138 , n48139 , n2327 , n48141 , n48142 , n2330 , n48144 , n2332 , n2333 , n48147 , 
 n2335 , n2336 , n48150 , n48151 , n48152 , n48153 , n48154 , n48155 , n2343 , n48157 , 
 n2345 , n48159 , n48160 , n2348 , n48162 , n48163 , n2351 , n48165 , n48166 , n48167 , 
 n2355 , n48169 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n48176 , n2364 , 
 n48178 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n48185 , n48186 , n2374 , 
 n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , 
 n2385 , n48199 , n48200 , n2388 , n48202 , n2390 , n2391 , n2392 , n2393 , n2394 , 
 n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , 
 n48218 , n48219 , n48220 , n2408 , n48222 , n2410 , n2411 , n48225 , n48226 , n2414 , 
 n48228 , n48229 , n2417 , n48231 , n2419 , n2420 , n2421 , n2422 , n2423 , n48237 , 
 n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , 
 n2435 , n2436 , n2437 , n48251 , n48252 , n2440 , n2441 , n2442 , n2443 , n2444 , 
 n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , 
 n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , 
 n48278 , n2466 , n2467 , n2468 , n2469 , n48283 , n48284 , n48285 , n2473 , n48287 , 
 n48288 , n48289 , n2477 , n48291 , n2479 , n48293 , n2481 , n48295 , n48296 , n2484 , 
 n48298 , n2486 , n48300 , n2488 , n48302 , n48303 , n2491 , n2492 , n2493 , n2494 , 
 n2495 , n2496 , n2497 , n48311 , n48312 , n2500 , n48314 , n2502 , n2503 , n48317 , 
 n48318 , n2506 , n48320 , n48321 , n2509 , n48323 , n2511 , n2512 , n2513 , n2514 , 
 n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , 
 n2525 , n2526 , n2527 , n2528 , n48342 , n2530 , n2531 , n2532 , n48346 , n2534 , 
 n48348 , n48349 , n48350 , n48351 , n48352 , n2540 , n48354 , n48355 , n2543 , n2544 , 
 n2545 , n2546 , n48360 , n2548 , n48362 , n2550 , n48364 , n2552 , n2553 , n48367 , 
 n2555 , n48369 , n48370 , n48371 , n2559 , n48373 , n48374 , n2562 , n48376 , n2564 , 
 n2565 , n2566 , n2567 , n2568 , n48382 , n48383 , n2571 , n2572 , n2573 , n2574 , 
 n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n48396 , n2584 , 
 n48398 , n2586 , n2587 , n2588 , n2589 , n48403 , n2591 , n2592 , n2593 , n2594 , 
 n48408 , n48409 , n2597 , n48411 , n2599 , n2600 , n2601 , n48415 , n48416 , n2604 , 
 n2605 , n48419 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n48426 , n2614 , 
 n2615 , n2616 , n48430 , n2618 , n48432 , n2620 , n48434 , n48435 , n2623 , n48437 , 
 n48438 , n2626 , n48440 , n48441 , n2629 , n2630 , n2631 , n48445 , n2633 , n48447 , 
 n48448 , n48449 , n2637 , n48451 , n2639 , n48453 , n2641 , n48455 , n2643 , n48457 , 
 n48458 , n2646 , n48460 , n2648 , n2649 , n48463 , n2651 , n48465 , n2653 , n48467 , 
 n48468 , n2656 , n2657 , n2658 , n48472 , n48473 , n2661 , n48475 , n48476 , n2664 , 
 n2665 , n48479 , n2667 , n48481 , n48482 , n48483 , n48484 , n2672 , n48486 , n48487 , 
 n2675 , n2676 , n2677 , n48491 , n2679 , n48493 , n48494 , n2682 , n48496 , n2684 , 
 n48498 , n48499 , n2687 , n48501 , n48502 , n48503 , n2691 , n48505 , n2693 , n48507 , 
 n48508 , n2696 , n48510 , n2698 , n2699 , n2700 , n2701 , n2702 , n48516 , n48517 , 
 n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n48526 , n2714 , 
 n2715 , n48529 , n2717 , n2718 , n2719 , n2720 , n2721 , n48535 , n2723 , n48537 , 
 n48538 , n48539 , n2727 , n48541 , n48542 , n48543 , n48544 , n48545 , n48546 , n2734 , 
 n2735 , n2736 , n48550 , n48551 , n2739 , n2740 , n2741 , n48555 , n2743 , n2744 , 
 n2745 , n48559 , n2747 , n48561 , n2749 , n2750 , n48564 , n2752 , n48566 , n2754 , 
 n48568 , n2756 , n48570 , n48571 , n2759 , n48573 , n48574 , n2762 , n48576 , n48577 , 
 n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , 
 n2775 , n2776 , n2777 , n48591 , n48592 , n2780 , n48594 , n2782 , n2783 , n48597 , 
 n48598 , n2786 , n48600 , n2788 , n48602 , n2790 , n48604 , n2792 , n48606 , n2794 , 
 n2795 , n2796 , n2797 , n2798 , n2799 , n48613 , n2801 , n2802 , n2803 , n48617 , 
 n48618 , n2806 , n48620 , n48621 , n48622 , n48623 , n2811 , n2812 , n48626 , n48627 , 
 n2815 , n48629 , n2817 , n48631 , n48632 , n2820 , n48634 , n48635 , n48636 , n48637 , 
 n48638 , n2826 , n2827 , n48641 , n2829 , n48643 , n2831 , n2832 , n48646 , n48647 , 
 n2835 , n48649 , n2837 , n2838 , n48652 , n2840 , n2841 , n2842 , n48656 , n2844 , 
 n48658 , n2846 , n48660 , n2848 , n48662 , n48663 , n2851 , n2852 , n48666 , n2854 , 
 n48668 , n48669 , n48670 , n2858 , n2859 , n48673 , n48674 , n48675 , n2863 , n48677 , 
 n2865 , n2866 , n2867 , n48681 , n2869 , n48683 , n48684 , n48685 , n48686 , n48687 , 
 n2875 , n48689 , n48690 , n2878 , n48692 , n48693 , n48694 , n2882 , n48696 , n2884 , 
 n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , 
 n2895 , n2896 , n2897 , n2898 , n2899 , n48713 , n2901 , n48715 , n48716 , n2904 , 
 n48718 , n2906 , n2907 , n2908 , n2909 , n48723 , n2911 , n2912 , n48726 , n2914 , 
 n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , 
 n2925 , n2926 , n2927 , n2928 , n48742 , n2930 , n48744 , n2932 , n48746 , n2934 , 
 n2935 , n2936 , n48750 , n2938 , n48752 , n48753 , n2941 , n2942 , n2943 , n2944 , 
 n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n48766 , n2954 , 
 n48768 , n48769 , n48770 , n2958 , n48772 , n48773 , n2961 , n48775 , n2963 , n48777 , 
 n48778 , n2966 , n2967 , n48781 , n2969 , n48783 , n48784 , n48785 , n48786 , n2974 , 
 n48788 , n48789 , n2977 , n48791 , n48792 , n2980 , n48794 , n48795 , n2983 , n48797 , 
 n48798 , n2986 , n48800 , n2988 , n2989 , n2990 , n2991 , n48805 , n48806 , n48807 , 
 n2995 , n48809 , n48810 , n2998 , n48812 , n3000 , n3001 , n48815 , n3003 , n48817 , 
 n3005 , n48819 , n48820 , n3008 , n48822 , n48823 , n3011 , n48825 , n3013 , n3014 , 
 n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n48836 , n48837 , 
 n3025 , n48839 , n48840 , n3028 , n3029 , n3030 , n3031 , n48845 , n3033 , n48847 , 
 n3035 , n48849 , n3037 , n48851 , n3039 , n48853 , n3041 , n48855 , n48856 , n3044 , 
 n3045 , n48859 , n48860 , n3048 , n48862 , n48863 , n3051 , n48865 , n48866 , n3054 , 
 n48868 , n3056 , n3057 , n3058 , n48872 , n3060 , n48874 , n3062 , n3063 , n48877 , 
 n3065 , n3066 , n48880 , n48881 , n3069 , n48883 , n48884 , n3072 , n48886 , n48887 , 
 n3075 , n48889 , n48890 , n3078 , n3079 , n48893 , n48894 , n3082 , n3083 , n48897 , 
 n3085 , n3086 , n3087 , n48901 , n3089 , n48903 , n48904 , n3092 , n48906 , n3094 , 
 n3095 , n48909 , n3097 , n48911 , n48912 , n3100 , n48914 , n48915 , n48916 , n3104 , 
 n48918 , n3106 , n48920 , n48921 , n3109 , n48923 , n48924 , n3112 , n48926 , n3114 , 
 n3115 , n3116 , n3117 , n3118 , n48932 , n3120 , n48934 , n3122 , n48936 , n3124 , 
 n3125 , n3126 , n48940 , n48941 , n3129 , n48943 , n3131 , n3132 , n48946 , n48947 , 
 n48948 , n3136 , n48950 , n3138 , n3139 , n3140 , n3141 , n48955 , n48956 , n3144 , 
 n48958 , n48959 , n3147 , n48961 , n48962 , n48963 , n3151 , n48965 , n48966 , n48967 , 
 n3155 , n48969 , n3157 , n48971 , n48972 , n3160 , n48974 , n3162 , n48976 , n3164 , 
 n3165 , n48979 , n48980 , n3168 , n48982 , n48983 , n3171 , n48985 , n48986 , n3174 , 
 n48988 , n48989 , n3177 , n3178 , n48992 , n48993 , n3181 , n3182 , n48996 , n48997 , 
 n3185 , n48999 , n3187 , n3188 , n49002 , n49003 , n3191 , n49005 , n3193 , n3194 , 
 n3195 , n49009 , n3197 , n49011 , n3199 , n49013 , n3201 , n3202 , n3203 , n49017 , 
 n49018 , n3206 , n49020 , n3208 , n3209 , n3210 , n3211 , n49025 , n3213 , n49027 , 
 n3215 , n49029 , n3217 , n49031 , n3219 , n49033 , n3221 , n49035 , n3223 , n49037 , 
 n3225 , n3226 , n49040 , n3228 , n3229 , n3230 , n49044 , n3232 , n49046 , n49047 , 
 n3235 , n49049 , n49050 , n3238 , n49052 , n3240 , n3241 , n49055 , n3243 , n49057 , 
 n3245 , n3246 , n49060 , n3248 , n49062 , n3250 , n3251 , n3252 , n3253 , n3254 , 
 n3255 , n3256 , n3257 , n3258 , n3259 , n49073 , n49074 , n3262 , n49076 , n3264 , 
 n3265 , n3266 , n3267 , n3268 , n49082 , n49083 , n3271 , n49085 , n3273 , n3274 , 
 n49088 , n3276 , n49090 , n3278 , n3279 , n49093 , n3281 , n49095 , n3283 , n49097 , 
 n49098 , n49099 , n3287 , n49101 , n3289 , n3290 , n3291 , n49105 , n49106 , n3294 , 
 n49108 , n3296 , n49110 , n3298 , n49112 , n3300 , n3301 , n3302 , n3303 , n3304 , 
 n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n49125 , n3313 , n49127 , 
 n3315 , n49129 , n49130 , n49131 , n49132 , n3320 , n49134 , n3322 , n49136 , n3324 , 
 n49138 , n3326 , n49140 , n49141 , n3329 , n49143 , n3331 , n49145 , n3333 , n3334 , 
 n49148 , n3336 , n49150 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , 
 n49158 , n3346 , n49160 , n3348 , n3349 , n49163 , n49164 , n3352 , n3353 , n49167 , 
 n49168 , n49169 , n49170 , n3358 , n49172 , n49173 , n49174 , n49175 , n49176 , n49177 , 
 n3365 , n3366 , n49180 , n3368 , n49182 , n49183 , n3371 , n3372 , n49186 , n49187 , 
 n3375 , n49189 , n49190 , n3378 , n49192 , n3380 , n49194 , n3382 , n3383 , n3384 , 
 n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n49205 , n49206 , n3395 , 
 n49208 , n3397 , n3398 , n49211 , n3400 , n49213 , n49214 , n49215 , n3404 , n49217 , 
 n3406 , n49219 , n49220 , n3409 , n49222 , n49223 , n3414 , n3415 , n3416 , n3417 , 
 n49228 , n3419 , n3420 , n3421 , n3422 , n49233 , n49234 , n3425 , n49236 , n3427 , 
 n49238 , n3429 , n49240 , n49241 , n49242 , n49243 , n3438 , n49245 , n49246 , n3441 , 
 n49248 , n3443 , n49250 , n49251 , n3446 , n3447 , n49254 , n3449 , n49256 , n49257 , 
 n3452 , n49259 , n49260 , n49261 , n3457 , n49263 , n3459 , n3460 , n3461 , n3462 , 
 n49268 , n49269 , n3465 , n49271 , n3472 , n49273 , n3474 , n49275 , n3476 , n49277 , 
 n49278 , n3486 , n49280 , n3488 , n3489 , n3490 , n49284 , n49285 , n3493 , n49287 , 
 n3495 , n49289 , n49290 , n3500 , n49292 , n49293 , n3511 , n49295 , n49296 , n49297 , 
 n3515 , n49299 , n49300 , n3518 , n49302 , n3520 , n49304 , n3522 , n3523 , n49307 , 
 n3525 , n49309 , n3527 , n49311 , n49312 , n3530 , n49314 , n3532 , n3533 , n3534 , 
 n3536 , n49319 , n49320 , n3539 , n49322 , n3541 , n49324 , n3543 , n49326 , n49327 , 
 n49328 , n3547 , n49330 , n49331 , n3550 , n49333 , n3552 , n49335 , n49336 , n49337 , 
 n3556 , n49339 , n49340 , n49341 , n3560 , n49343 , n49344 , n3563 , n49346 , n49347 , 
 n3566 , n49349 , n3568 , n3569 , n3570 , n49353 , n49354 , n3573 , n49356 , n49357 , 
 n3576 , n49359 , n3578 , n49361 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , 
 n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n49377 , 
 n3598 , n3599 , n3600 , n49381 , n3602 , n49383 , n3604 , n49385 , n49386 , n3607 , 
 n49388 , n3609 , n3610 , n3611 , n3612 , n49393 , n3614 , n49395 , n3616 , n3617 , 
 n3618 , n3619 , n3620 , n49401 , n3622 , n49403 , n3624 , n49405 , n49406 , n49407 , 
 n3628 , n49409 , n49410 , n3631 , n49412 , n49413 , n3634 , n49415 , n49416 , n3637 , 
 n49418 , n49419 , n3640 , n49421 , n49422 , n3644 , n3645 , n3646 , n49426 , n3648 , 
 n3649 , n3650 , n3651 , n3652 , n49432 , n3654 , n49434 , n49435 , n3657 , n49437 , 
 n49438 , n3660 , n49440 , n49441 , n3663 , n3664 , n49444 , n49445 , n3667 , n49447 , 
 n49448 , n3670 , n49450 , n49451 , n49452 , n3674 , n49454 , n49455 , n49456 , n3678 , 
 n49458 , n49459 , n3681 , n49461 , n49462 , n49463 , n49464 , n3686 , n49466 , n49467 , 
 n3689 , n49469 , n49470 , n3692 , n49472 , n3696 , n3697 , n49475 , n3699 , n49477 , 
 n3701 , n3702 , n3703 , n49481 , n49482 , n49483 , n3707 , n49485 , n49486 , n3710 , 
 n3711 , n49489 , n3713 , n3714 , n49492 , n3716 , n49494 , n3718 , n49496 , n49497 , 
 n3721 , n49499 , n49500 , n3724 , n49502 , n49503 , n3727 , n49505 , n49506 , n3730 , 
 n3731 , n49509 , n3733 , n3734 , n49512 , n3736 , n3737 , n49515 , n3739 , n49517 , 
 n49518 , n3742 , n49520 , n3744 , n3745 , n3746 , n3747 , n3748 , n49526 , n3750 , 
 n49528 , n49529 , n3753 , n49531 , n49532 , n49533 , n3757 , n49535 , n3759 , n49537 , 
 n49538 , n3762 , n49540 , n49541 , n3765 , n49543 , n49544 , n3768 , n49546 , n3770 , 
 n49548 , n3772 , n49550 , n49551 , n3775 , n49553 , n49554 , n3778 , n49556 , n49557 , 
 n3781 , n49559 , n3783 , n49561 , n3785 , n3786 , n49564 , n3788 , n3789 , n49567 , 
 n49568 , n3792 , n3793 , n49571 , n49572 , n3796 , n49574 , n3798 , n3799 , n49577 , 
 n49578 , n3802 , n49580 , n3804 , n3805 , n3806 , n3807 , n3808 , n49586 , n3810 , 
 n49588 , n3812 , n3813 , n3814 , n3815 , n49593 , n3817 , n49595 , n3819 , n3820 , 
 n49598 , n3822 , n49600 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , 
 n3831 , n3832 , n3833 , n3834 , n3835 , n49613 , n49614 , n3838 , n3839 , n49617 , 
 n3841 , n3842 , n49620 , n3844 , n3845 , n3846 , n49624 , n3848 , n49626 , n3850 , 
 n3851 , n49629 , n3853 , n3854 , n3855 , n3856 , n49634 , n49635 , n3859 , n49637 , 
 n3861 , n49639 , n3863 , n49641 , n49642 , n3866 , n3867 , n3868 , n49646 , n3870 , 
 n49648 , n49649 , n49650 , n3874 , n49652 , n3876 , n49654 , n49655 , n3879 , n49657 , 
 n3881 , n3882 , n3883 , n49661 , n3886 , n49663 , n3888 , n49665 , n49666 , n3891 , 
 n49668 , n49669 , n49670 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n49677 , 
 n3902 , n49679 , n49680 , n3905 , n3906 , n3907 , n49684 , n3909 , n3910 , n49687 , 
 n49688 , n3913 , n49690 , n49691 , n49692 , n3917 , n49694 , n49695 , n49696 , n3921 , 
 n49698 , n49699 , n3924 , n49701 , n49702 , n3927 , n3928 , n49705 , n49706 , n3931 , 
 n3932 , n49709 , n49710 , n3935 , n3936 , n49713 , n49714 , n3939 , n49716 , n3941 , 
 n49718 , n3943 , n49720 , n3945 , n49722 , n49723 , n3948 , n49725 , n3950 , n49727 , 
 n49728 , n3953 , n3954 , n3955 , n49732 , n49733 , n3958 , n49735 , n49736 , n3961 , 
 n49738 , n49739 , n49740 , n3965 , n49742 , n3967 , n49744 , n49745 , n3970 , n49747 , 
 n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , 
 n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , 
 n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , 
 n4002 , n49779 , n4004 , n49781 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , 
 n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , 
 n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n49807 , 
 n49808 , n4033 , n49810 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , 
 n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , 
 n4052 , n4053 , n4054 , n49831 , n49832 , n4057 , n49834 , n49835 , n4060 , n4061 , 
 n4062 , n49839 , n49840 , n4065 , n4066 , n49843 , n4068 , n49845 , n4070 , n4071 , 
 n4072 , n4073 , n4074 , n4075 , n4076 , n49853 , n4078 , n4079 , n49856 , n49857 , 
 n4082 , n49859 , n49860 , n4085 , n49862 , n49863 , n4088 , n4089 , n49866 , n49867 , 
 n4092 , n49869 , n49870 , n4095 , n49872 , n49873 , n4098 , n4099 , n4100 , n4101 , 
 n4102 , n4103 , n49880 , n4105 , n49882 , n4107 , n4108 , n4109 , n4110 , n4111 , 
 n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , 
 n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n49907 , 
 n4132 , n49909 , n4134 , n49911 , n49912 , n4137 , n49914 , n49915 , n4140 , n49917 , 
 n49918 , n49919 , n4144 , n4146 , n49922 , n4148 , n49924 , n49925 , n49926 , n4152 , 
 n49928 , n49929 , n49930 , n49931 , n49932 , n49933 , n49934 , n4160 , n49936 , n49937 , 
 n49938 , n49939 , n49940 , n4166 , n49942 , n49943 , n49944 , n49945 , n49946 , n49947 , 
 n49948 , n4174 , n49950 , n4176 , n49952 , n4178 , n49954 , n4180 , n49956 , n4182 , 
 n49958 , n4186 , n49960 , n4188 , n49962 , n4190 , n49964 , n4192 , n49966 , n49967 , 
 n49968 , n4196 , n49970 , n4198 , n49972 , n4200 , n49974 , n4202 , n49976 , n4204 , 
 n49978 , n4206 , n49980 , n49981 , n49982 , n49983 , n49984 , n4212 , n49986 , n4214 , 
 n49988 , n4216 , n49990 , n4218 , n49992 , n4220 , n49994 , n4222 , n49996 , n4224 , 
 n49998 , n49999 , n50000 , n50001 , n50002 , n4230 , n50004 , n50005 , n50006 , n50007 , 
 n50008 , n4236 , n50010 , n50011 , n50012 , n50013 , n50014 , n50015 , n50016 , n4244 , 
 n50018 , n50019 , n50020 , n50021 , n50022 , n4250 , n50024 , n4252 , n50026 , n4254 , 
 n50028 , n50029 , n50030 , n50031 , n50032 , n50033 , n50034 , n4262 , n50036 , n50037 , 
 n4265 , n50039 , n50040 , n4268 , n50042 , n50043 , n50044 , n4272 , n4273 , n4274 , 
 n50048 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , 
 n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , 
 n4295 , n4296 , n4297 , n4298 , n4299 , n50073 , n4301 , n4302 , n4303 , n4304 , 
 n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n50087 , 
 n4315 , n4316 , n4317 , n50091 , n4319 , n50093 , n4321 , n4322 , n50096 , n50097 , 
 n4325 , n50099 , n4327 , n50101 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , 
 n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , 
 n4345 , n4346 , n4347 , n4348 , n4349 , n50123 , n4351 , n50125 , n50126 , n4354 , 
 n4355 , n50129 , n4357 , n4358 , n50132 , n50133 , n4361 , n50135 , n50136 , n4364 , 
 n4365 , n50139 , n4367 , n4368 , n4369 , n50143 , n4371 , n50145 , n50146 , n50147 , 
 n4375 , n50149 , n50150 , n4378 , n50152 , n50153 , n4381 , n50155 , n4383 , n4384 , 
 n50158 , n4386 , n4387 , n50161 , n50162 , n4390 , n50164 , n4392 , n4393 , n50167 , 
 n50168 , n4396 , n50170 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , 
 n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , 
 n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n50195 , n50196 , n4424 , 
 n50198 , n4426 , n4427 , n4428 , n4429 , n4430 , n50204 , n4432 , n50206 , n4434 , 
 n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , 
 n4445 , n50219 , n4447 , n4448 , n4449 , n4450 , n4451 , n50225 , n4453 , n4454 , 
 n50228 , n4456 , n4457 , n4458 , n50232 , n4460 , n50234 , n4462 , n50236 , n4464 , 
 n50238 , n50239 , n4467 , n4468 , n50242 , n50243 , n4471 , n4472 , n50246 , n50247 , 
 n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n50255 , n4483 , n4484 , 
 n50258 , n50259 , n4487 , n50261 , n50262 , n4490 , n50264 , n50265 , n4493 , n50267 , 
 n4495 , n50269 , n4497 , n4498 , n50272 , n4500 , n50274 , n4502 , n4503 , n4504 , 
 n4505 , n50279 , n4507 , n50281 , n50282 , n50283 , n4511 , n50285 , n50286 , n4514 , 
 n50288 , n50289 , n4517 , n4518 , n4519 , n50293 , n50294 , n4522 , n4523 , n4524 , 
 n50298 , n50299 , n4527 , n4528 , n50302 , n50303 , n50304 , n50305 , n4533 , n50307 , 
 n50308 , n50309 , n50310 , n4538 , n50312 , n50313 , n4541 , n50315 , n50316 , n4544 , 
 n50318 , n50319 , n4547 , n50321 , n50322 , n4550 , n4551 , n4552 , n4553 , n50327 , 
 n50328 , n4556 , n50330 , n4558 , n50332 , n4560 , n50334 , n50335 , n4563 , n50337 , 
 n50338 , n4566 , n50340 , n50341 , n4569 , n50343 , n50344 , n50345 , n4573 , n50347 , 
 n50348 , n4576 , n4577 , n50351 , n4579 , n50353 , n4581 , n4582 , n4583 , n4584 , 
 n4585 , n4586 , n4587 , n4588 , n50362 , n4590 , n50364 , n4592 , n4593 , n4594 , 
 n4595 , n50369 , n4597 , n50371 , n50372 , n4600 , n50374 , n50375 , n50376 , n50377 , 
 n4605 , n50379 , n50380 , n4608 , n50382 , n50383 , n4611 , n4612 , n4613 , n4614 , 
 n50388 , n50389 , n4617 , n50391 , n50392 , n4620 , n4621 , n4622 , n4623 , n4624 , 
 n50398 , n4626 , n4627 , n50401 , n50402 , n4630 , n4631 , n50405 , n4633 , n4634 , 
 n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n50417 , 
 n4645 , n50419 , n4647 , n4648 , n50422 , n50423 , n4651 , n50425 , n50426 , n4654 , 
 n50428 , n50429 , n4657 , n50431 , n4659 , n50433 , n4661 , n50435 , n50436 , n4664 , 
 n4665 , n50439 , n50440 , n4668 , n4669 , n50443 , n4671 , n4672 , n4673 , n4674 , 
 n50448 , n4676 , n4677 , n50451 , n4679 , n50453 , n50454 , n4682 , n50456 , n50457 , 
 n50458 , n4686 , n50460 , n4688 , n50462 , n4690 , n4691 , n4692 , n4693 , n50467 , 
 n4695 , n50469 , n4697 , n50471 , n4699 , n50473 , n4701 , n50475 , n50476 , n4704 , 
 n50478 , n4706 , n4707 , n50481 , n4709 , n50483 , n4711 , n50485 , n50486 , n4714 , 
 n50488 , n50489 , n4717 , n50491 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , 
 n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n50507 , 
 n4735 , n50509 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , 
 n4745 , n4746 , n4747 , n4748 , n50522 , n50523 , n50524 , n4752 , n50526 , n4754 , 
 n50528 , n50529 , n4757 , n50531 , n50532 , n4760 , n50534 , n50535 , n4763 , n50537 , 
 n50538 , n4766 , n50540 , n50541 , n50542 , n4770 , n50544 , n4772 , n4773 , n50547 , 
 n4775 , n50549 , n50550 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , 
 n50558 , n4786 , n4787 , n50561 , n50562 , n4790 , n50564 , n4792 , n50566 , n4794 , 
 n4795 , n50569 , n4797 , n50571 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , 
 n4805 , n50579 , n4807 , n50581 , n50582 , n4810 , n50584 , n50585 , n4813 , n50587 , 
 n50588 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , 
 n4825 , n4826 , n4827 , n50601 , n4829 , n50603 , n50604 , n4832 , n50606 , n50607 , 
 n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n50617 , 
 n50618 , n50619 , n4847 , n50621 , n50622 , n4850 , n50624 , n50625 , n4853 , n4854 , 
 n50628 , n4856 , n4857 , n50631 , n50632 , n4860 , n50634 , n50635 , n4863 , n50637 , 
 n50638 , n50639 , n4867 , n50641 , n4869 , n4870 , n4871 , n4872 , n50646 , n4874 , 
 n50648 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , 
 n4885 , n4886 , n4887 , n4888 , n50662 , n4890 , n50664 , n4892 , n4893 , n4894 , 
 n4895 , n4896 , n50670 , n4898 , n50672 , n50673 , n4901 , n4902 , n4903 , n4904 , 
 n4905 , n4906 , n4907 , n50681 , n4909 , n50683 , n50684 , n4912 , n50686 , n50687 , 
 n4915 , n4916 , n4917 , n4918 , n50692 , n50693 , n4921 , n50695 , n50696 , n4924 , 
 n50698 , n50699 , n50700 , n4928 , n50702 , n4930 , n50704 , n50705 , n4933 , n50707 , 
 n50708 , n50709 , n4937 , n50711 , n4939 , n50713 , n4941 , n50715 , n4943 , n50717 , 
 n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , 
 n4955 , n4956 , n50730 , n50731 , n4959 , n50733 , n50734 , n4962 , n50736 , n4964 , 
 n50738 , n4966 , n50740 , n50741 , n4969 , n4970 , n50744 , n4972 , n50746 , n50747 , 
 n4975 , n50749 , n4977 , n50751 , n4979 , n4980 , n4981 , n4982 , n4983 , n50757 , 
 n4985 , n50759 , n50760 , n50761 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , 
 n50768 , n4996 , n4997 , n50771 , n50772 , n5000 , n5001 , n50775 , n5003 , n5004 , 
 n50778 , n5006 , n5007 , n50781 , n5009 , n50783 , n50784 , n5012 , n50786 , n5014 , 
 n50788 , n50789 , n5017 , n5018 , n50792 , n5020 , n50794 , n50795 , n5023 , n5024 , 
 n50798 , n50799 , n5027 , n5028 , n50802 , n5030 , n50804 , n5032 , n5033 , n50807 , 
 n50808 , n5036 , n50810 , n50811 , n5039 , n50813 , n50814 , n50815 , n5043 , n50817 , 
 n50818 , n5046 , n50820 , n5048 , n50822 , n5050 , n50824 , n5052 , n50826 , n50827 , 
 n5055 , n5056 , n50830 , n50831 , n5059 , n50833 , n50834 , n5062 , n50836 , n5064 , 
 n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , 
 n5075 , n5076 , n5077 , n50851 , n5079 , n50853 , n5081 , n5082 , n50856 , n50857 , 
 n5085 , n50859 , n50860 , n5088 , n50862 , n5090 , n5091 , n5092 , n5093 , n5094 , 
 n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n50875 , n5103 , n5104 , 
 n5105 , n50879 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , 
 n5115 , n5116 , n5117 , n50891 , n50892 , n5120 , n50894 , n5122 , n5123 , n5124 , 
 n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n50906 , n5134 , 
 n50908 , n5136 , n50910 , n5138 , n50912 , n5140 , n50914 , n5142 , n50916 , n5144 , 
 n50918 , n5146 , n50920 , n5148 , n50922 , n5150 , n50924 , n5152 , n50926 , n5154 , 
 n50928 , n5156 , n50930 , n5158 , n50932 , n5160 , n50934 , n5162 , n50936 , n5164 , 
 n50938 , n50939 , n50940 , n50941 , n50942 , n5170 , n50944 , n5172 , n50946 , n50947 , 
 n50948 , n50949 , n5177 , n50951 , n50952 , n50953 , n50954 , n50955 , n50956 , n50957 , 
 n50958 , n50959 , n50960 , n50961 , n50962 , n50963 , n50964 , n50965 , n50966 , n50967 , 
 n50968 , n50969 , n50970 , n50971 , n50972 , n50973 , n50974 , n50975 , n50976 , n50977 , 
 n50978 , n50979 , n50980 , n50981 , n50982 , n50983 , n50984 , n50985 , n50986 , n50987 , 
 n50988 , n50989 , n50990 , n50991 , n50992 , n50993 , n50994 , n50995 , n50996 , n50997 , 
 n50998 , n50999 , n51000 , n51001 , n51002 , n51003 , n51004 , n51005 , n51006 , n51007 , 
 n51008 , n51009 , n51010 , n51011 , n51012 , n51013 , n51014 , n51015 , n51016 , n51017 , 
 n51018 , n51019 , n51020 , n51021 , n51022 , n51023 , n51024 , n51025 , n51026 , n51027 , 
 n51028 , n51029 , n51030 , n51031 , n51032 , n51033 , n51034 , n51035 , n51036 , n51037 , 
 n51038 , n51039 , n51040 , n51041 , n51042 , n51043 , n51044 , n51045 , n51046 , n51047 , 
 n51048 , n51049 , n51050 , n51051 , n51052 , n51053 , n51054 , n51055 , n51056 , n51057 , 
 n51058 , n51059 , n51060 , n51061 , n51062 , n51063 , n51064 , n51065 , n51066 , n51067 , 
 n51068 , n51069 , n51070 , n51071 , n51072 , n51073 , n51074 , n51075 , n51076 , n51077 , 
 n51078 , n51079 , n51080 , n51081 , n51082 , n51083 , n51084 , n51085 , n51086 , n51087 , 
 n51088 , n51089 , n51090 , n51091 , n51092 , n51093 , n51094 , n51095 , n51096 , n51097 , 
 n51098 , n51099 , n51100 , n51101 , n51102 , n51103 , n51104 , n51105 , n51106 , n51107 , 
 n51108 , n51109 , n51110 , n51111 , n51112 , n51113 , n51114 , n51115 , n51116 , n51117 , 
 n51118 , n51119 , n51120 , n51121 , n51122 , n51123 , n51124 , n51125 , n51126 , n51127 , 
 n51128 , n51129 , n51130 , n51131 , n51132 , n51133 , n51134 , n51135 , n51136 , n51137 , 
 n51138 , n51139 , n51140 , n51141 , n51142 , n51143 , n51144 , n51145 , n51146 , n51147 , 
 n51148 , n51149 , n51150 , n51151 , n51152 , n51153 , n51154 , n51155 , n51156 , n51157 , 
 n51158 , n51159 , n51160 , n51161 , n51162 , n51163 , n51164 , n51165 , n51166 , n51167 , 
 n51168 , n51169 , n51170 , n51171 , n51172 , n51173 , n51174 , n51175 , n51176 , n51177 , 
 n51178 , n51179 , n51180 , n51181 , n51182 , n51183 , n51184 , n51185 , n51186 , n51187 , 
 n51188 , n51189 , n51190 , n51191 , n51192 , n51193 , n51194 , n51195 , n51196 , n51197 , 
 n51198 , n51199 , n51200 , n51201 , n51202 , n51203 , n51204 , n51205 , n51206 , n51207 , 
 n51208 , n51209 , n51210 , n51211 , n51212 , n51213 , n51214 , n51215 , n51216 , n51217 , 
 n51218 , n51219 , n51220 , n51221 , n51222 , n51223 , n51224 , n51225 , n51226 , n51227 , 
 n51228 , n51229 , n51230 , n51231 , n51232 , n51233 , n51234 , n51235 , n51236 , n51237 , 
 n51238 , n51239 , n51240 , n51241 , n51242 , n51243 , n51244 , n51245 , n51246 , n51247 , 
 n51248 , n51249 , n51250 , n51251 , n51252 , n51253 , n51254 , n51255 , n51256 , n51257 , 
 n51258 , n51259 , n51260 , n51261 , n51262 , n51263 , n51264 , n51265 , n51266 , n51267 , 
 n51268 , n51269 , n51270 , n51271 , n51272 , n51273 , n51274 , n51275 , n51276 , n51277 , 
 n51278 , n51279 , n51280 , n51281 , n51282 , n51283 , n51284 , n51285 , n51286 , n51287 , 
 n51288 , n51289 , n51290 , n51291 , n51292 , n51293 , n51294 , n51295 , n51296 , n51297 , 
 n51298 , n51299 , n51300 , n51301 , n51302 , n51303 , n51304 , n51305 , n51306 , n51307 , 
 n51308 , n51309 , n51310 , n51311 , n51312 , n51313 , n51314 , n51315 , n51316 , n51317 , 
 n51318 , n51319 , n51320 , n51321 , n51322 , n51323 , n5199 , n51325 , n5201 , n5202 , 
 n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , 
 n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n51345 , n5221 , n51347 , 
 n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , 
 n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , 
 n5243 , n51369 , n5245 , n51371 , n5247 , n5248 , n51374 , n51375 , n5251 , n51377 , 
 n5253 , n51379 , n5255 , n51381 , n5257 , n5258 , n5259 , n5260 , n51386 , n5262 , 
 n5263 , n51389 , n51390 , n5266 , n51392 , n51393 , n5269 , n51395 , n5271 , n51397 , 
 n5273 , n51399 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , 
 n51408 , n51409 , n5285 , n51411 , n51412 , n5288 , n51414 , n51415 , n5291 , n51417 , 
 n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , 
 n5303 , n51429 , n51430 , n5306 , n51432 , n51433 , n5309 , n51435 , n5311 , n51437 , 
 n51438 , n5314 , n51440 , n5316 , n51442 , n5318 , n5319 , n5320 , n5321 , n5322 , 
 n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n51456 , n5332 , 
 n51458 , n5334 , n51460 , n51461 , n5337 , n51463 , n5339 , n5340 , n5341 , n5342 , 
 n5343 , n51469 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n51476 , n5352 , 
 n5353 , n51479 , n51480 , n5356 , n51482 , n51483 , n5359 , n51485 , n5361 , n5362 , 
 n51488 , n51489 , n51490 , n5366 , n5367 , n51493 , n5369 , n5370 , n51496 , n51497 , 
 n5373 , n51499 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n51506 , n5382 , 
 n51508 , n51509 , n51510 , n5386 , n51512 , n5388 , n5389 , n51515 , n51516 , n5392 , 
 n5393 , n51519 , n51520 , n5396 , n51522 , n5398 , n51524 , n5400 , n5401 , n51527 , 
 n5403 , n51529 , n5405 , n51531 , n51532 , n5408 , n5409 , n51535 , n51536 , n5412 , 
 n51538 , n51539 , n5415 , n51541 , n51542 , n51543 , n5419 , n51545 , n51546 , n5422 , 
 n51548 , n51549 , n5425 , n5426 , n5427 , n51553 , n51554 , n5430 , n51556 , n5432 , 
 n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , 
 n5443 , n5444 , n51570 , n5446 , n51572 , n5448 , n5449 , n51575 , n5451 , n51577 , 
 n5453 , n5454 , n51580 , n51581 , n5457 , n51583 , n5459 , n51585 , n51586 , n5462 , 
 n5463 , n51589 , n51590 , n5466 , n51592 , n5468 , n51594 , n51595 , n5471 , n5472 , 
 n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n51604 , n5480 , n5481 , n51607 , 
 n51608 , n5484 , n51610 , n51611 , n5487 , n51613 , n51614 , n5490 , n5491 , n51617 , 
 n51618 , n5494 , n51620 , n5496 , n5497 , n51623 , n5499 , n51625 , n51626 , n5502 , 
 n51628 , n5504 , n51630 , n5506 , n51632 , n51633 , n5509 , n51635 , n5511 , n5512 , 
 n51638 , n5514 , n51640 , n5516 , n51642 , n51643 , n5519 , n51645 , n51646 , n5522 , 
 n51648 , n51649 , n5525 , n51651 , n51652 , n5528 , n51654 , n51655 , n5531 , n51657 , 
 n51658 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n51665 , n5541 , n51667 , 
 n5543 , n51669 , n5545 , n51671 , n5547 , n51673 , n5549 , n51675 , n5551 , n5552 , 
 n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n51687 , 
 n51688 , n5564 , n51690 , n5566 , n51692 , n5568 , n5569 , n51695 , n51696 , n5572 , 
 n51698 , n51699 , n5575 , n51701 , n51702 , n5578 , n5579 , n51705 , n51706 , n5582 , 
 n51708 , n51709 , n5585 , n51711 , n51712 , n5588 , n51714 , n5590 , n5591 , n5592 , 
 n5593 , n5594 , n51720 , n5596 , n5597 , n5598 , n51724 , n51725 , n5601 , n51727 , 
 n51728 , n5604 , n51730 , n51731 , n5607 , n51733 , n51734 , n5610 , n51736 , n5612 , 
 n51738 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n51747 , 
 n5623 , n51749 , n51750 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , 
 n5633 , n5634 , n5635 , n51761 , n5637 , n51763 , n5639 , n51765 , n51766 , n5642 , 
 n51768 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n51777 , 
 n5653 , n5654 , n5655 , n5656 , n5657 , n51783 , n5659 , n51785 , n5661 , n51787 , 
 n5663 , n5664 , n5665 , n51791 , n51792 , n51793 , n5669 , n51795 , n51796 , n5672 , 
 n51798 , n51799 , n5675 , n5676 , n5677 , n51803 , n5679 , n5680 , n5681 , n5682 , 
 n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , 
 n5693 , n5694 , n5695 , n51821 , n51822 , n51823 , n51824 , n51825 , n51826 , n51827 , 
 n51828 , n51829 , n51830 , n5703 , n51832 , n5705 , n51834 , n5707 , n51836 , n51837 , 
 n51838 , n5711 , n51840 , n5713 , n51842 , n51843 , n51844 , n5717 , n51846 , n51847 , 
 n51848 , n51849 , n51850 , n51851 , n51852 , n51853 , n51854 , n51855 , n51856 , n51857 , 
 n51858 , n51859 , n51860 , n51861 , n51862 , n51863 , n51864 , n51865 , n51866 , n51867 , 
 n51868 , n51869 , n51870 , n51871 , n51872 , n51873 , n51874 , n51875 , n51876 , n51877 , 
 n51878 , n51879 , n51880 , n51881 , n51882 , n51883 , n51884 , n51885 , n51886 , n51887 , 
 n51888 , n51889 , n51890 , n51891 , n51892 , n51893 , n51894 , n51895 , n51896 , n51897 , 
 n51898 , n51899 , n51900 , n51901 , n51902 , n51903 , n51904 , n51905 , n51906 , n51907 , 
 n51908 , n51909 , n51910 , n51911 , n51912 , n51913 , n51914 , n51915 , n51916 , n51917 , 
 n51918 , n51919 , n51920 , n51921 , n51922 , n51923 , n51924 , n51925 , n5726 , n5727 , 
 n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n51935 , n5736 , n51937 , 
 n51938 , n5739 , n51940 , n51941 , n5742 , n51943 , n5744 , n5745 , n51946 , n51947 , 
 n5748 , n51949 , n5750 , n51951 , n51952 , n5753 , n51954 , n5755 , n5756 , n5757 , 
 n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , 
 n5768 , n5769 , n5770 , n51971 , n5772 , n51973 , n5774 , n5775 , n5776 , n51977 , 
 n51978 , n5779 , n5780 , n51981 , n5782 , n51983 , n5784 , n5785 , n51986 , n51987 , 
 n5788 , n51989 , n51990 , n5791 , n51992 , n5793 , n5794 , n5795 , n5796 , n5797 , 
 n51998 , n51999 , n5800 , n52001 , n5802 , n5803 , n5804 , n52005 , n5806 , n5807 , 
 n5808 , n52009 , n52010 , n5811 , n5812 , n5813 , n52014 , n52015 , n5816 , n5817 , 
 n52018 , n52019 , n5820 , n5821 , n52022 , n52023 , n5824 , n5825 , n5826 , n5827 , 
 n5828 , n5829 , n5830 , n52031 , n5832 , n5833 , n52034 , n5835 , n5836 , n5837 , 
 n52038 , n52039 , n52040 , n5841 , n52042 , n5843 , n5844 , n52045 , n52046 , n5847 , 
 n52048 , n52049 , n5850 , n52051 , n52052 , n5853 , n5854 , n5855 , n5856 , n52057 , 
 n5858 , n5859 , n52060 , n5861 , n5862 , n52063 , n52064 , n5865 , n52066 , n52067 , 
 n5868 , n52069 , n52070 , n52071 , n5872 , n52073 , n5874 , n5875 , n5876 , n5877 , 
 n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , 
 n5888 , n5889 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , 
 n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , 
 n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , 
 n52118 , n5922 , n5923 , n5924 , n52122 , n52123 , n5927 , n52125 , n52126 , n5930 , 
 n5931 , n52129 , n5933 , n52131 , n52132 , n5936 , n5937 , n52135 , n52136 , n5940 , 
 n5941 , n52139 , n52140 , n5944 , n52142 , n52143 , n5947 , n5948 , n5949 , n5950 , 
 n5951 , n5952 , n5953 , n52151 , n5955 , n52153 , n5957 , n5958 , n5959 , n5960 , 
 n5961 , n52159 , n5963 , n52161 , n5965 , n5966 , n52164 , n52165 , n5969 , n5970 , 
 n52168 , n5972 , n5973 , n52171 , n52172 , n52173 , n5977 , n52175 , n52176 , n5980 , 
 n52178 , n52179 , n5983 , n5984 , n5985 , n5986 , n5987 , n52185 , n5989 , n52187 , 
 n5991 , n52189 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n52196 , n52197 , 
 n6001 , n52199 , n6003 , n52201 , n52202 , n6006 , n52204 , n52205 , n6009 , n52207 , 
 n52208 , n6012 , n6013 , n6014 , n52212 , n6016 , n6017 , n52215 , n52216 , n6020 , 
 n6021 , n6022 , n52220 , n6024 , n52222 , n6026 , n6027 , n52225 , n6029 , n6030 , 
 n6031 , n6032 , n52230 , n52231 , n6035 , n52233 , n52234 , n52235 , n52236 , n6040 , 
 n52238 , n52239 , n6043 , n52241 , n52242 , n6046 , n52244 , n6048 , n52246 , n52247 , 
 n6051 , n52249 , n52250 , n52251 , n6055 , n52253 , n6057 , n52255 , n52256 , n6060 , 
 n52258 , n52259 , n52260 , n6064 , n52262 , n6066 , n6067 , n6068 , n6069 , n6070 , 
 n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n52274 , n52275 , n6079 , n52277 , 
 n6081 , n6082 , n6083 , n52281 , n6085 , n52283 , n6087 , n52285 , n52286 , n6090 , 
 n6091 , n52289 , n52290 , n6094 , n52292 , n52293 , n6097 , n52295 , n52296 , n52297 , 
 n6101 , n52299 , n6103 , n6104 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , 
 n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6124 , n6125 , n6126 , n6127 , 
 n6128 , n52319 , n6130 , n52321 , n6132 , n6133 , n52324 , n52325 , n6136 , n52327 , 
 n52328 , n6139 , n52330 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , 
 n6148 , n6149 , n6150 , n52341 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , 
 n52348 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n52356 , n6167 , 
 n52358 , n6169 , n52360 , n6171 , n52362 , n6173 , n6174 , n52365 , n52366 , n6177 , 
 n52368 , n52369 , n6180 , n52371 , n52372 , n6183 , n6184 , n52375 , n52376 , n6187 , 
 n52378 , n52379 , n6190 , n6191 , n52382 , n52383 , n6194 , n52385 , n52386 , n6197 , 
 n6198 , n52389 , n6200 , n52391 , n52392 , n6203 , n52394 , n52395 , n6206 , n6207 , 
 n6208 , n6209 , n6210 , n6211 , n6212 , n52403 , n6214 , n52405 , n52406 , n6217 , 
 n52408 , n52409 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , 
 n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n52426 , n6237 , 
 n6238 , n52429 , n52430 , n6241 , n6242 , n52433 , n52434 , n6245 , n6246 , n52437 , 
 n6248 , n52439 , n6250 , n6251 , n52442 , n52443 , n6254 , n52445 , n52446 , n6257 , 
 n52448 , n6259 , n6260 , n6261 , n6262 , n6263 , n52454 , n6265 , n52456 , n52457 , 
 n52458 , n6269 , n52460 , n6271 , n52462 , n52463 , n6274 , n52465 , n52466 , n6277 , 
 n6278 , n52469 , n52470 , n52471 , n6282 , n52473 , n52474 , n6285 , n52476 , n6287 , 
 n6288 , n52479 , n52480 , n6291 , n52482 , n6293 , n52484 , n52485 , n6296 , n52487 , 
 n52488 , n6299 , n6300 , n6301 , n52492 , n52493 , n6304 , n6305 , n6306 , n6307 , 
 n6308 , n6309 , n52500 , n6311 , n52502 , n6313 , n52504 , n6315 , n6316 , n52507 , 
 n52508 , n6319 , n52510 , n52511 , n6322 , n52513 , n52514 , n6325 , n52516 , n52517 , 
 n6328 , n52519 , n52520 , n6331 , n6332 , n52523 , n6334 , n52525 , n6336 , n6337 , 
 n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n52536 , n6347 , 
 n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n52547 , 
 n6358 , n6359 , n52550 , n6361 , n52552 , n6363 , n52554 , n6365 , n6366 , n6367 , 
 n52558 , n52559 , n6370 , n6371 , n52562 , n6373 , n6374 , n52565 , n52566 , n52567 , 
 n6378 , n52569 , n6380 , n6381 , n6382 , n6383 , n52574 , n52575 , n52576 , n6387 , 
 n52578 , n6389 , n52580 , n52581 , n6392 , n52583 , n6394 , n6395 , n52586 , n52587 , 
 n6398 , n52589 , n6400 , n52591 , n52592 , n6403 , n52594 , n52595 , n6406 , n52597 , 
 n52598 , n6409 , n52600 , n6411 , n52602 , n6413 , n6414 , n6415 , n6416 , n6417 , 
 n52608 , n52609 , n6420 , n52611 , n6422 , n6423 , n6424 , n52615 , n6426 , n52617 , 
 n52618 , n6429 , n6430 , n6431 , n52622 , n6433 , n6434 , n52625 , n52626 , n6437 , 
 n6438 , n6439 , n52630 , n6441 , n52632 , n6443 , n6444 , n52635 , n6446 , n52637 , 
 n52638 , n6449 , n6450 , n52641 , n6452 , n52643 , n6454 , n6455 , n52646 , n52647 , 
 n6458 , n6459 , n52650 , n52651 , n6462 , n52653 , n52654 , n6465 , n6466 , n6467 , 
 n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , 
 n6478 , n6479 , n6480 , n52671 , n52672 , n6483 , n52674 , n6485 , n6486 , n6487 , 
 n6488 , n6489 , n6490 , n6491 , n52682 , n6493 , n52684 , n6495 , n52686 , n6497 , 
 n6498 , n52689 , n6500 , n52691 , n6502 , n52693 , n52694 , n6505 , n52696 , n52697 , 
 n6508 , n6509 , n52700 , n52701 , n6512 , n6513 , n52704 , n6515 , n6516 , n52707 , 
 n52708 , n52709 , n6520 , n6521 , n52712 , n52713 , n6524 , n6525 , n6526 , n6527 , 
 n6528 , n52719 , n52720 , n6531 , n52722 , n52723 , n52724 , n52725 , n6536 , n52727 , 
 n52728 , n6539 , n52730 , n52731 , n6542 , n52733 , n6544 , n52735 , n52736 , n52737 , 
 n6548 , n52739 , n52740 , n6551 , n52742 , n52743 , n6554 , n52745 , n52746 , n52747 , 
 n6558 , n52749 , n52750 , n6561 , n6562 , n6563 , n52754 , n52755 , n6566 , n52757 , 
 n52758 , n6569 , n52760 , n6571 , n6572 , n6573 , n52764 , n6575 , n6576 , n52767 , 
 n52768 , n52769 , n6580 , n52771 , n52772 , n6583 , n6584 , n52775 , n52776 , n6587 , 
 n6588 , n52779 , n52780 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n52787 , 
 n6598 , n6599 , n6600 , n52791 , n52792 , n6603 , n6604 , n6605 , n52796 , n6607 , 
 n6608 , n52799 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , 
 n6618 , n6619 , n6620 , n6621 , n52812 , n6623 , n52814 , n6625 , n52816 , n6627 , 
 n6628 , n52819 , n6630 , n52821 , n6632 , n52823 , n52824 , n6635 , n52826 , n6637 , 
 n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , 
 n52838 , n52839 , n6650 , n52841 , n6652 , n52843 , n6654 , n6655 , n6656 , n6657 , 
 n6658 , n6659 , n6660 , n6661 , n52852 , n6663 , n52854 , n6665 , n6666 , n6667 , 
 n6668 , n6669 , n6670 , n52861 , n6672 , n6673 , n52864 , n6675 , n52866 , n6677 , 
 n52868 , n52869 , n6680 , n52871 , n52872 , n6683 , n6684 , n6685 , n52876 , n52877 , 
 n6688 , n52879 , n52880 , n6691 , n6692 , n52883 , n6694 , n6695 , n52886 , n52887 , 
 n6698 , n52889 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n52896 , n6707 , 
 n6708 , n6709 , n6710 , n52901 , n6712 , n52903 , n6714 , n52905 , n6716 , n52907 , 
 n52908 , n6719 , n6720 , n6721 , n52912 , n52913 , n6724 , n52915 , n52916 , n6727 , 
 n52918 , n52919 , n52920 , n6731 , n6732 , n52923 , n6734 , n52925 , n52926 , n6737 , 
 n6738 , n52929 , n6740 , n6741 , n6742 , n6743 , n6744 , n52935 , n6746 , n6747 , 
 n6748 , n6749 , n52940 , n6751 , n6752 , n6753 , n6754 , n6755 , n52946 , n6757 , 
 n52948 , n52949 , n6760 , n6761 , n52952 , n52953 , n6764 , n52955 , n52956 , n6767 , 
 n52958 , n6769 , n52960 , n6771 , n6772 , n6773 , n6774 , n52965 , n6776 , n52967 , 
 n52968 , n6779 , n52970 , n6781 , n6782 , n52973 , n52974 , n6785 , n52976 , n6787 , 
 n6788 , n52979 , n52980 , n6791 , n52982 , n6793 , n52984 , n6795 , n6796 , n52987 , 
 n6798 , n52989 , n6800 , n52991 , n6802 , n6803 , n6804 , n6805 , n52996 , n6807 , 
 n52998 , n6809 , n6810 , n53001 , n53002 , n6813 , n53004 , n6815 , n6816 , n6817 , 
 n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n53015 , n6826 , n6827 , 
 n6828 , n6829 , n6830 , n6831 , n6832 , n53023 , n6834 , n6835 , n6836 , n6837 , 
 n6838 , n53029 , n53030 , n6841 , n53032 , n6843 , n53034 , n6845 , n53036 , n6847 , 
 n53038 , n53039 , n53040 , n6851 , n53042 , n6853 , n53044 , n53045 , n6856 , n53047 , 
 n6858 , n6859 , n6860 , n53051 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , 
 n6868 , n6869 , n6870 , n53061 , n6872 , n53063 , n6874 , n6875 , n6876 , n6877 , 
 n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , 
 n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , 
 n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , 
 n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , 
 n6918 , n53109 , n6920 , n53111 , n53112 , n6923 , n6924 , n6925 , n6926 , n6927 , 
 n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , 
 n6938 , n6939 , n6940 , n6941 , n53132 , n6943 , n53134 , n53135 , n6946 , n53137 , 
 n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , 
 n6958 , n6959 , n53150 , n6961 , n6962 , n53153 , n6964 , n53155 , n6966 , n6967 , 
 n6968 , n53159 , n6970 , n53161 , n53162 , n6973 , n53164 , n6975 , n6976 , n6977 , 
 n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , 
 n6988 , n6989 , n53180 , n53181 , n6992 , n53183 , n53184 , n6995 , n53186 , n6997 , 
 n53188 , n6999 , n53190 , n7001 , n53192 , n7003 , n53194 , n53195 , n53196 , n7007 , 
 n53198 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , 
 n7018 , n53209 , n7020 , n53211 , n53212 , n53213 , n7024 , n53215 , n7026 , n7027 , 
 n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , 
 n7038 , n7039 , n7040 , n7041 , n7042 , n7044 , n53234 , n7046 , n53236 , n7048 , 
 n53238 , n7050 , n7051 , n7052 , n7053 , n53243 , n53244 , n7056 , n53246 , n7058 , 
 n53248 , n53249 , n53250 , n7062 , n53252 , n53253 , n7065 , n7066 , n53256 , n7068 , 
 n53258 , n7070 , n53260 , n7072 , n53262 , n53263 , n7075 , n53265 , n53266 , n7078 , 
 n7079 , n7080 , n7081 , n7082 , n7083 , n53273 , n7085 , n7086 , n53276 , n7088 , 
 n53278 , n7090 , n53280 , n7092 , n53282 , n7094 , n7095 , n7096 , n7097 , n53287 , 
 n7099 , n7100 , n7101 , n7102 , n53292 , n53293 , n53294 , n7106 , n53296 , n53297 , 
 n53298 , n7110 , n53300 , n53301 , n53302 , n7114 , n7115 , n7116 , n7117 , n53307 , 
 n53308 , n53309 , n7121 , n53311 , n53312 , n7124 , n7125 , n53315 , n53316 , n53317 , 
 n7129 , n7130 , n53320 , n7132 , n7133 , n53323 , n53324 , n53325 , n7137 , n7138 , 
 n53328 , n7140 , n7141 , n53331 , n53332 , n7144 , n53334 , n53335 , n7147 , n53337 , 
 n53338 , n7150 , n53340 , n7152 , n53342 , n53343 , n7155 , n53345 , n53346 , n7158 , 
 n7159 , n53349 , n53350 , n7162 , n7163 , n53353 , n53354 , n53355 , n7168 , n53357 , 
 n53358 , n7171 , n53360 , n7173 , n7174 , n7175 , n53364 , n53365 , n7178 , n53367 , 
 n53368 , n7181 , n53370 , n53371 , n7184 , n53373 , n53374 , n7187 , n7188 , n53377 , 
 n7190 , n53379 , n7192 , n7193 , n53382 , n7200 , n53384 , n7202 , n53386 , n7204 , 
 n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n53394 , n53395 , n7213 , n53397 , 
 n7215 , n53399 , n53400 , n53401 , n7219 , n53403 , n7221 , n53405 , n53406 , n7224 , 
 n53408 , n53409 , n7227 , n53411 , n53412 , n7230 , n7231 , n53415 , n7233 , n7234 , 
 n53418 , n53419 , n53420 , n53421 , n7239 , n53423 , n53424 , n53425 , n7243 , n53427 , 
 n53428 , n7246 , n53430 , n7248 , n53432 , n53433 , n7251 , n53435 , n7253 , n7254 , 
 n53438 , n53439 , n7257 , n7258 , n53442 , n53443 , n7261 , n7262 , n7263 , n53447 , 
 n53448 , n7266 , n7267 , n53451 , n53452 , n7270 , n53454 , n53455 , n7273 , n53457 , 
 n53458 , n7276 , n7277 , n53461 , n53462 , n7280 , n53464 , n53465 , n7283 , n53467 , 
 n53468 , n7286 , n53470 , n53471 , n7289 , n53473 , n53474 , n53475 , n53476 , n7294 , 
 n53478 , n7296 , n53480 , n53481 , n7299 , n53483 , n53484 , n7302 , n53486 , n7304 , 
 n53488 , n53489 , n53490 , n7308 , n53492 , n53493 , n7311 , n7312 , n53496 , n7314 , 
 n7315 , n53499 , n53500 , n7318 , n53502 , n7320 , n7321 , n53505 , n53506 , n7324 , 
 n7325 , n53509 , n53510 , n7328 , n7329 , n7330 , n53514 , n53515 , n53516 , n53517 , 
 n7335 , n53519 , n53520 , n7338 , n7339 , n53523 , n53524 , n53525 , n7343 , n53527 , 
 n7345 , n53529 , n53530 , n7348 , n53532 , n53533 , n7351 , n7352 , n53536 , n53537 , 
 n7355 , n53539 , n53540 , n7358 , n53542 , n53543 , n7361 , n53545 , n53546 , n7364 , 
 n53548 , n53549 , n7367 , n7368 , n7369 , n53553 , n53554 , n7372 , n53556 , n53557 , 
 n7375 , n7376 , n53560 , n7378 , n7379 , n53563 , n7381 , n53565 , n53566 , n7384 , 
 n53568 , n7386 , n7387 , n7388 , n53572 , n53573 , n7391 , n53575 , n53576 , n7394 , 
 n7395 , n7396 , n53580 , n53581 , n53582 , n7400 , n53584 , n7402 , n53586 , n7404 , 
 n53588 , n7406 , n7407 , n53591 , n7409 , n53593 , n7411 , n53595 , n7413 , n53597 , 
 n7415 , n7416 , n53600 , n7418 , n53602 , n7420 , n53604 , n53605 , n7423 , n53607 , 
 n53608 , n7426 , n53610 , n7428 , n53612 , n53613 , n53614 , n53615 , n7436 , n53617 , 
 n53618 , n7439 , n53620 , n53621 , n53622 , n7443 , n53624 , n53625 , n53626 , n53627 , 
 n7448 , n53629 , n7450 , n53631 , n7452 , n7453 , n7454 , n53635 , n7456 , n53637 , 
 n53638 , n7459 , n7460 , n53641 , n7462 , n53643 , n7464 , n53645 , n53646 , n53647 , 
 n53648 , n7469 , n53650 , n53651 , n7472 , n53653 , n53654 , n7475 , n53656 , n53657 , 
 n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n53665 , n7486 , n53667 , 
 n7488 , n7489 , n53670 , n53671 , n7492 , n53673 , n7494 , n7495 , n7496 , n53677 , 
 n7498 , n53679 , n7500 , n53681 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , 
 n7508 , n7509 , n7510 , n53691 , n7512 , n53693 , n7514 , n53695 , n7516 , n7517 , 
 n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , 
 n7528 , n7529 , n7530 , n7535 , n53712 , n53713 , n7538 , n53715 , n7540 , n7541 , 
 n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n53727 , 
 n53728 , n7581 , n53730 , n7583 , n7584 , n7585 , n7586 , n53735 , n53736 , n7589 , 
 n53738 , n7591 , n53740 , n53741 , n53742 , n7595 , n53744 , n53745 , n7598 , n7599 , 
 n7600 , n7601 , n7602 , n53751 , n7604 , n7605 , n7606 , n7607 , n53756 , n7609 , 
 n7610 , n7611 , n7612 , n53761 , n53762 , n7615 , n53764 , n53765 , n7618 , n7619 , 
 n7620 , n7621 , n7622 , n7623 , n7624 , n53773 , n7626 , n7627 , n7628 , n7629 , 
 n53778 , n53779 , n53780 , n7633 , n53782 , n53783 , n53784 , n7637 , n53786 , n53787 , 
 n53788 , n7641 , n7642 , n7643 , n7644 , n53793 , n53794 , n53795 , n7648 , n53797 , 
 n53798 , n53799 , n7652 , n53801 , n53802 , n53803 , n7656 , n53805 , n53806 , n7659 , 
 n53808 , n7661 , n53810 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , 
 n53818 , n7671 , n53820 , n7673 , n53822 , n7675 , n7676 , n53825 , n7678 , n53827 , 
 n53828 , n7681 , n53830 , n53831 , n7684 , n7685 , n7686 , n7687 , n53836 , n7689 , 
 n53838 , n53839 , n7692 , n53841 , n53842 , n7695 , n7696 , n7697 , n7698 , n7699 , 
 n7700 , n7701 , n7702 , n53851 , n7704 , n7705 , n7706 , n7707 , n53856 , n53857 , 
 n7710 , n53859 , n7712 , n53861 , n53862 , n7715 , n53864 , n53865 , n53866 , n53867 , 
 n7720 , n53869 , n7722 , n7723 , n53872 , n7725 , n53874 , n53875 , n7728 , n53877 , 
 n53878 , n7731 , n7732 , n7733 , n7734 , n53883 , n7736 , n53885 , n7738 , n53887 , 
 n7740 , n53889 , n7742 , n53891 , n53892 , n7745 , n7746 , n7747 , n53896 , n7749 , 
 n53898 , n53899 , n53900 , n53901 , n7754 , n7755 , n7756 , n7757 , n7758 , n53907 , 
 n7760 , n53909 , n53910 , n53911 , n53912 , n7765 , n7766 , n7767 , n7768 , n7769 , 
 n53918 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , 
 n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , 
 n7790 , n7791 , n7792 , n7793 , n53942 , n7795 , n7796 , n7797 , n7798 , n7799 , 
 n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n53954 , n7807 , n7808 , n7809 , 
 n7810 , n7811 , n53960 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , 
 n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7829 , n7830 , 
 n7850 , n7851 , n53980 , n53981 , n53982 , n7855 , n53984 , n7857 , n53986 , n7859 , 
 n53988 , n7861 , n53990 , n7863 , n53992 , n7865 , n53994 , n7867 , n53996 , n7869 , 
 n53998 , n7871 , n54000 , n7873 , n54002 , n54003 , n7877 , n54005 , n7879 , n54007 , 
 n7881 , n54009 , n54010 , n54011 , n54012 , n54013 , n54014 , n54015 , n54016 , n54017 , 
 n54018 , n54019 , n7893 , n54021 , n54022 , n54023 , n54024 , n7923 , n7924 , n7925 , 
 n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n54034 , n7933 , n54036 , n54037 , 
 n7936 , n54039 , n54040 , n7939 , n54042 , n7946 , n7957 , n54045 , n54046 , n54047 , 
 n7961 , n54049 , n54050 , n7964 , n54052 , n54053 , n54054 , n54055 , n7971 , n54057 , 
 n54058 , n54059 , n54060 , n54061 , n54062 , n54063 , n7979 , n54065 , n54066 , n54067 , 
 n7983 , n54069 , n54070 , n54071 , n54072 , n54073 , n54074 , n54075 , n54076 , n54077 , 
 n54078 , n54079 , n54080 , n54081 , n54082 , n54083 , n54084 , n54085 , n54086 , n54087 , 
 n54088 , n54089 , n54090 , n54091 , n54092 , n54093 , n54094 , n54095 , n54096 , n54097 , 
 n54098 , n54099 , n54100 , n54101 , n54102 , n54103 , n54104 , n54105 , n54106 , n54107 , 
 n54108 , n54109 , n54110 , n54111 , n54112 , n54113 , n54114 , n54115 , n54116 , n54117 , 
 n54118 , n54119 , n54120 , n54121 , n54122 , n54123 , n54124 , n54125 , n54126 , n54127 , 
 n54128 , n54129 , n54130 , n54131 , n54132 , n8056 , n54134 , n54135 , n54136 , n8060 , 
 n54138 , n54139 , n54140 , n8064 , n8065 , n54143 , n8067 , n8068 , n54146 , n8070 , 
 n54148 , n8072 , n54150 , n8074 , n8075 , n8079 , n8080 , n8081 , n54156 , n54157 , 
 n8084 , n54159 , n8086 , n8087 , n8088 , n8089 , n8093 , n8094 , n8095 , n8096 , 
 n8097 , n8098 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n54177 , 
 n8108 , n54179 , n8110 , n8112 , n8113 , n8114 , n8115 , n8116 , n8121 , n8122 , 
 n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , 
 n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , 
 n8143 , n8144 , n8145 , n8146 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , 
 n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , 
 n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , 
 n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , 
 n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , 
 n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8206 , n8207 , 
 n8208 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , 
 n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , 
 n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , 
 n8239 , n54299 , n54300 , n8242 , n54302 , C0n , C0 , C1n , C1 ;
buf ( n370 , n0 );
buf ( n371 , n1 );
buf ( n372 , n2 );
buf ( n373 , n3 );
buf ( n374 , n4 );
buf ( n375 , n5 );
buf ( n376 , n6 );
buf ( n377 , n7 );
buf ( n378 , n8 );
buf ( n379 , n9 );
buf ( n380 , n10 );
buf ( n381 , n11 );
buf ( n382 , n12 );
buf ( n383 , n13 );
buf ( n384 , n14 );
buf ( n385 , n15 );
buf ( n386 , n16 );
buf ( n387 , n17 );
buf ( n388 , n18 );
buf ( n389 , n19 );
buf ( n390 , n20 );
buf ( n391 , n21 );
buf ( n392 , n22 );
buf ( n393 , n23 );
buf ( n394 , n24 );
buf ( n395 , n25 );
buf ( n396 , n26 );
buf ( n397 , n27 );
buf ( n398 , n28 );
buf ( n399 , n29 );
buf ( n400 , n30 );
buf ( n401 , n31 );
buf ( n402 , n32 );
buf ( n403 , n33 );
buf ( n404 , n34 );
buf ( n405 , n35 );
buf ( n406 , n36 );
buf ( n407 , n37 );
buf ( n408 , n38 );
buf ( n409 , n39 );
buf ( n410 , n40 );
buf ( n411 , n41 );
buf ( n412 , n42 );
buf ( n413 , n43 );
buf ( n414 , n44 );
buf ( n415 , n45 );
buf ( n416 , n46 );
buf ( n417 , n47 );
buf ( n418 , n48 );
buf ( n419 , n49 );
buf ( n420 , n50 );
buf ( n421 , n51 );
buf ( n422 , n52 );
buf ( n423 , n53 );
buf ( n424 , n54 );
buf ( n425 , n55 );
buf ( n56 , n426 );
buf ( n57 , n427 );
buf ( n58 , n428 );
buf ( n59 , n429 );
buf ( n60 , n430 );
buf ( n61 , n431 );
buf ( n62 , n432 );
buf ( n63 , n433 );
buf ( n64 , n434 );
buf ( n65 , n435 );
buf ( n66 , n436 );
buf ( n67 , n437 );
buf ( n68 , n438 );
buf ( n69 , n439 );
buf ( n70 , n440 );
buf ( n71 , n441 );
buf ( n72 , n442 );
buf ( n73 , n443 );
buf ( n74 , n444 );
buf ( n75 , n445 );
buf ( n76 , n446 );
buf ( n77 , n447 );
buf ( n78 , n448 );
buf ( n79 , n449 );
buf ( n80 , n450 );
buf ( n81 , n451 );
buf ( n82 , n452 );
buf ( n83 , n453 );
buf ( n84 , n454 );
buf ( n85 , n455 );
buf ( n86 , n456 );
buf ( n87 , n457 );
buf ( n88 , n458 );
buf ( n89 , n459 );
buf ( n90 , n460 );
buf ( n91 , n461 );
buf ( n92 , n462 );
buf ( n93 , n463 );
buf ( n94 , n464 );
buf ( n95 , n465 );
buf ( n96 , n466 );
buf ( n97 , n467 );
buf ( n98 , n468 );
buf ( n99 , n469 );
buf ( n100 , n470 );
buf ( n101 , n471 );
buf ( n102 , n472 );
buf ( n103 , n473 );
buf ( n104 , n474 );
buf ( n105 , n475 );
buf ( n106 , n476 );
buf ( n107 , n477 );
buf ( n108 , n478 );
buf ( n109 , n479 );
buf ( n110 , n480 );
buf ( n111 , n481 );
buf ( n112 , n482 );
buf ( n113 , n483 );
buf ( n114 , n484 );
buf ( n115 , n485 );
buf ( n116 , n486 );
buf ( n117 , n487 );
buf ( n118 , n488 );
buf ( n119 , n489 );
buf ( n120 , n490 );
buf ( n121 , n491 );
buf ( n122 , n492 );
buf ( n123 , n493 );
buf ( n124 , n494 );
buf ( n125 , n495 );
buf ( n126 , n496 );
buf ( n127 , n497 );
buf ( n128 , n498 );
buf ( n129 , n499 );
buf ( n130 , n500 );
buf ( n131 , n501 );
buf ( n132 , n502 );
buf ( n133 , n503 );
buf ( n134 , n504 );
buf ( n135 , n505 );
buf ( n136 , n506 );
buf ( n137 , n507 );
buf ( n138 , n508 );
buf ( n139 , n509 );
buf ( n140 , n510 );
buf ( n141 , n511 );
buf ( n142 , n512 );
buf ( n143 , n513 );
buf ( n144 , n514 );
buf ( n145 , n515 );
buf ( n146 , n516 );
buf ( n147 , n517 );
buf ( n148 , n518 );
buf ( n149 , n519 );
buf ( n150 , n520 );
buf ( n151 , n521 );
buf ( n152 , n522 );
buf ( n153 , n523 );
buf ( n154 , n524 );
buf ( n155 , n525 );
buf ( n156 , n526 );
buf ( n157 , n527 );
buf ( n158 , n528 );
buf ( n159 , n529 );
buf ( n160 , n530 );
buf ( n161 , n531 );
buf ( n162 , n532 );
buf ( n163 , n533 );
buf ( n164 , n534 );
buf ( n165 , n535 );
buf ( n166 , n536 );
buf ( n167 , n537 );
buf ( n168 , n538 );
buf ( n169 , n539 );
buf ( n170 , n540 );
buf ( n171 , n541 );
buf ( n172 , n542 );
buf ( n173 , n543 );
buf ( n174 , n544 );
buf ( n175 , n545 );
buf ( n176 , n546 );
buf ( n177 , n547 );
buf ( n178 , n548 );
buf ( n179 , n549 );
buf ( n180 , n550 );
buf ( n181 , n551 );
buf ( n182 , n552 );
buf ( n183 , n553 );
buf ( n184 , n554 );
buf ( n426 , C0 );
buf ( n427 , C0 );
buf ( n428 , C0 );
buf ( n429 , C0 );
buf ( n430 , C0 );
buf ( n431 , C0 );
buf ( n432 , C0 );
buf ( n433 , C0 );
buf ( n434 , C0 );
buf ( n435 , C0 );
buf ( n436 , C0 );
buf ( n437 , C0 );
buf ( n438 , C0 );
buf ( n439 , C0 );
buf ( n440 , C0 );
buf ( n441 , C0 );
buf ( n442 , C0 );
buf ( n443 , C0 );
buf ( n444 , C0 );
buf ( n445 , C0 );
buf ( n446 , C0 );
buf ( n447 , C0 );
buf ( n448 , C0 );
buf ( n449 , C0 );
buf ( n450 , C0 );
buf ( n451 , C0 );
buf ( n452 , C0 );
buf ( n453 , C0 );
buf ( n454 , C0 );
buf ( n455 , C0 );
buf ( n456 , C0 );
buf ( n457 , C0 );
buf ( n458 , C0 );
buf ( n459 , C0 );
buf ( n460 , C0 );
buf ( n461 , C0 );
buf ( n462 , C0 );
buf ( n463 , C0 );
buf ( n464 , C0 );
buf ( n465 , C0 );
buf ( n466 , C0 );
buf ( n467 , C0 );
buf ( n468 , C0 );
buf ( n469 , C0 );
buf ( n470 , C0 );
buf ( n471 , C0 );
buf ( n472 , C0 );
buf ( n473 , C0 );
buf ( n474 , C0 );
buf ( n475 , C0 );
buf ( n476 , C0 );
buf ( n477 , C0 );
buf ( n478 , C0 );
buf ( n479 , C0 );
buf ( n480 , C0 );
buf ( n481 , C0 );
buf ( n482 , C0 );
buf ( n483 , C0 );
buf ( n484 , C0 );
buf ( n485 , C0 );
buf ( n486 , C0 );
buf ( n487 , C0 );
buf ( n488 , C0 );
buf ( n489 , C0 );
buf ( n490 , n8183 );
buf ( n491 , n8149 );
buf ( n492 , n8162 );
buf ( n493 , n8098 );
buf ( n494 , n8238 );
buf ( n495 , n8081 );
buf ( n496 , n53735 );
buf ( n497 , n8212 );
buf ( n498 , n8196 );
buf ( n499 , n8239 );
buf ( n500 , n8239 );
buf ( n501 , n8239 );
buf ( n502 , n8239 );
buf ( n503 , n8239 );
buf ( n504 , n8239 );
buf ( n505 , n8239 );
buf ( n506 , n8158 );
buf ( n507 , n8158 );
buf ( n508 , n8158 );
buf ( n509 , n8158 );
buf ( n510 , n8158 );
buf ( n511 , n8158 );
buf ( n512 , n8158 );
buf ( n513 , n8158 );
buf ( n514 , n8158 );
buf ( n515 , n8158 );
buf ( n516 , n8158 );
buf ( n517 , n8158 );
buf ( n518 , n8159 );
buf ( n519 , n8159 );
buf ( n520 , n8159 );
buf ( n521 , n8159 );
buf ( n522 , n8159 );
buf ( n523 , n8159 );
buf ( n524 , n8159 );
buf ( n525 , n8159 );
buf ( n526 , n8159 );
buf ( n527 , n8159 );
buf ( n528 , n8159 );
buf ( n529 , n8159 );
buf ( n530 , n53243 );
buf ( n531 , n8175 );
buf ( n532 , n8218 );
buf ( n533 , n53292 );
buf ( n534 , n53307 );
buf ( n535 , n53756 );
buf ( n536 , n53793 );
buf ( n537 , n8143 );
buf ( n538 , n53778 );
buf ( n539 , n53856 );
buf ( n540 , n54302 );
buf ( n541 , n53836 );
buf ( n542 , n8202 );
buf ( n543 , n8187 );
buf ( n544 , n53883 );
buf ( n545 , n53907 );
buf ( n546 , n53918 );
buf ( n547 , n54146 );
buf ( n548 , n54092 );
buf ( n549 , n54130 );
buf ( n550 , n54134 );
buf ( n551 , n8129 );
buf ( n552 , n54123 );
buf ( n553 , n54126 );
buf ( n554 , n8228 );
not ( n40212 , n370 );
nand ( n40213 , n370 , n374 );
not ( n40214 , n40213 );
nand ( n40215 , n371 , n373 );
not ( n40216 , n40215 );
or ( n40217 , n40214 , n40216 );
and ( n40218 , n370 , n375 );
xor ( n40219 , n372 , n40218 );
and ( n40220 , n372 , n373 );
and ( n40221 , n40219 , n40220 );
and ( n40222 , n372 , n40218 );
or ( n40223 , n40221 , n40222 );
nand ( n40224 , n40217 , n40223 );
nand ( n40225 , n370 , n373 );
nand ( n40226 , n371 , n372 );
xor ( n40227 , n40225 , n40226 );
not ( n40228 , n371 );
xor ( n40229 , n40227 , n40228 );
not ( n40230 , n40213 );
not ( n40231 , n40215 );
nand ( n40232 , n40230 , n40231 );
nand ( n40233 , n40224 , n40229 , n40232 );
nand ( n40234 , n40225 , n40226 );
nand ( n40235 , n40225 , n40228 );
nand ( n40236 , n40226 , n40228 );
nand ( n40237 , n40234 , n40235 , n40236 );
nand ( n40238 , n370 , n372 );
nand ( n40239 , n40237 , n40238 );
nand ( n40240 , n40233 , n40239 );
nor ( n40241 , n40212 , n40240 );
not ( n40242 , n40241 );
nand ( n40243 , n371 , n374 );
not ( n40244 , n40243 );
xor ( n40245 , n372 , n40218 );
xor ( n40246 , n40245 , n40220 );
not ( n40247 , n40246 );
not ( n40248 , n40247 );
or ( n40249 , n40244 , n40248 );
nand ( n40250 , n370 , n376 );
not ( n40251 , n40250 );
not ( n40252 , n40251 );
nand ( n40253 , n371 , n375 );
not ( n40254 , n40253 );
not ( n40255 , n40254 );
or ( n40256 , n40252 , n40255 );
not ( n40257 , n40253 );
not ( n40258 , n40250 );
or ( n40259 , n40257 , n40258 );
and ( n40260 , n372 , n374 );
nand ( n40261 , n40259 , n40260 );
nand ( n40262 , n40256 , n40261 );
nand ( n40263 , n40249 , n40262 );
not ( n40264 , n40243 );
nand ( n40265 , n40246 , n40264 );
and ( n40266 , n40263 , n40265 );
not ( n40267 , n40231 );
not ( n40268 , n40213 );
and ( n40269 , n40267 , n40268 );
and ( n40270 , n40213 , n40231 );
nor ( n40271 , n40269 , n40270 );
xor ( n40272 , n40223 , n40271 );
nand ( n40273 , n40266 , n40272 );
not ( n40274 , n40273 );
nand ( n40275 , n373 , n374 );
not ( n40276 , n40275 );
not ( n40277 , n370 );
not ( n40278 , n377 );
or ( n40279 , n40277 , n40278 );
nand ( n40280 , n371 , n376 );
nand ( n40281 , n40279 , n40280 );
not ( n40282 , n40281 );
and ( n40283 , n372 , n375 );
not ( n40284 , n40283 );
or ( n40285 , n40282 , n40284 );
nand ( n40286 , n371 , n376 , n370 , n377 );
nand ( n40287 , n40285 , n40286 );
nor ( n40288 , n40276 , n40287 );
nand ( n40289 , n372 , n374 );
nand ( n40290 , n371 , n375 );
nand ( n40291 , n370 , n376 );
and ( n40292 , n40290 , n40291 );
not ( n40293 , n40290 );
and ( n40294 , n40293 , n40251 );
nor ( n40295 , n40292 , n40294 );
xor ( n40296 , n40289 , n40295 );
or ( n40297 , n40288 , n40296 );
not ( n40298 , n40275 );
nand ( n40299 , n40298 , n40287 );
nand ( n40300 , n40297 , n40299 );
not ( n40301 , n40300 );
not ( n40302 , n40301 );
xor ( n40303 , n40264 , n40262 );
xnor ( n40304 , n40303 , n40246 );
not ( n40305 , n40304 );
or ( n40306 , n40302 , n40305 );
nand ( n40307 , n373 , n375 , n372 , n376 );
not ( n40308 , n40307 );
nand ( n40309 , n40275 , n373 );
not ( n40310 , n40309 );
and ( n40311 , n40308 , n40310 );
nand ( n40312 , n372 , n375 );
nand ( n40313 , n371 , n376 );
and ( n40314 , n40312 , n40313 );
not ( n40315 , n40312 );
not ( n40316 , n40280 );
and ( n40317 , n40315 , n40316 );
nor ( n40318 , n40314 , n40317 );
and ( n40319 , n370 , n377 );
xor ( n40320 , n40318 , n40319 );
nand ( n40321 , n40309 , n40307 );
and ( n40322 , n40320 , n40321 );
nor ( n40323 , n40311 , n40322 );
xor ( n40324 , n40275 , n40287 );
xnor ( n40325 , n40324 , n40296 );
nand ( n40326 , n40323 , n40325 );
nand ( n40327 , n40306 , n40326 );
not ( n40328 , n40327 );
not ( n40329 , n40328 );
not ( n40330 , n40320 );
not ( n40331 , n40307 );
not ( n40332 , n374 );
not ( n40333 , n373 );
or ( n40334 , n40332 , n40333 );
nand ( n40335 , n40334 , n373 );
not ( n40336 , n40335 );
or ( n40337 , n40331 , n40336 );
or ( n40338 , n40335 , n40307 );
nand ( n40339 , n40337 , n40338 );
not ( n40340 , n40339 );
and ( n40341 , n40330 , n40340 );
and ( n40342 , n40339 , n40320 );
nor ( n40343 , n40341 , n40342 );
nand ( n40344 , n374 , n375 );
nand ( n40345 , n371 , n377 );
xor ( n40346 , n40344 , n40345 );
nand ( n40347 , n373 , n375 );
nand ( n40348 , n376 , n372 );
xnor ( n40349 , n40347 , n40348 );
and ( n40350 , n40346 , n40349 );
and ( n40351 , n40344 , n40345 );
or ( n40352 , n40350 , n40351 );
nand ( n40353 , n40343 , n40352 );
not ( n40354 , n40353 );
xor ( n40355 , n40344 , n40345 );
xor ( n40356 , n40355 , n40349 );
nand ( n40357 , n372 , n377 );
not ( n40358 , n40357 );
nand ( n40359 , n373 , n376 );
not ( n40360 , n40359 );
and ( n40361 , n40358 , n40360 );
nand ( n40362 , n40357 , n40359 );
not ( n40363 , n375 );
and ( n40364 , n40363 , n374 );
and ( n40365 , n40362 , n40364 );
nor ( n40366 , n40361 , n40365 );
nand ( n40367 , n40356 , n40366 );
not ( n40368 , n40367 );
nand ( n40369 , n377 , n374 , n375 );
not ( n40370 , n40369 );
nand ( n40371 , n375 , n377 );
nand ( n40372 , n377 , n376 );
nor ( n40373 , n40371 , n40372 );
nand ( n40374 , n40370 , n40373 );
nand ( n40375 , n374 , n376 );
not ( n40376 , n40375 );
nand ( n40377 , n373 , n377 );
not ( n40378 , n40377 );
or ( n40379 , n40376 , n40378 );
nand ( n40380 , n374 , n376 );
nand ( n40381 , n373 , n377 );
or ( n40382 , n40380 , n40381 );
nand ( n40383 , n40379 , n40382 );
nand ( n40384 , n40383 , n40369 );
and ( n40385 , n374 , n377 );
nand ( n40386 , n375 , n376 );
nor ( n40387 , n40385 , n40386 );
and ( n40388 , n40384 , n40387 );
nor ( n40389 , n40369 , n40383 );
nor ( n40390 , n40388 , n40389 );
nand ( n40391 , n40374 , n40390 );
not ( n40392 , n40391 );
or ( n40393 , n40357 , n40359 );
not ( n40394 , n373 );
not ( n40395 , n376 );
or ( n40396 , n40394 , n40395 );
nand ( n40397 , n372 , n377 );
nand ( n40398 , n40396 , n40397 );
nand ( n40399 , n40393 , n40398 );
not ( n40400 , n40399 );
not ( n40401 , n40364 );
and ( n40402 , n40400 , n40401 );
and ( n40403 , n40364 , n40399 );
nor ( n40404 , n40402 , n40403 );
not ( n40405 , n40275 );
and ( n40406 , n377 , n376 );
nand ( n40407 , n40405 , n40406 );
nand ( n40408 , n40404 , n40407 );
not ( n40409 , n40408 );
or ( n40410 , n40392 , n40409 );
not ( n40411 , n40404 );
not ( n40412 , n40407 );
nand ( n40413 , n40411 , n40412 );
nand ( n40414 , n40410 , n40413 );
not ( n40415 , n40414 );
or ( n40416 , n40368 , n40415 );
or ( n40417 , n40356 , n40366 );
nand ( n40418 , n40416 , n40417 );
not ( n40419 , n40418 );
or ( n40420 , n40354 , n40419 );
not ( n40421 , n40343 );
not ( n40422 , n40352 );
nand ( n40423 , n40421 , n40422 );
nand ( n40424 , n40420 , n40423 );
not ( n40425 , n40424 );
or ( n40426 , n40329 , n40425 );
not ( n40427 , n40304 );
not ( n40428 , n40301 );
and ( n40429 , n40427 , n40428 );
nand ( n40430 , n40304 , n40301 );
nor ( n40431 , n40323 , n40325 );
and ( n40432 , n40430 , n40431 );
nor ( n40433 , n40429 , n40432 );
nand ( n40434 , n40426 , n40433 );
not ( n40435 , n40434 );
or ( n40436 , n40274 , n40435 );
nor ( n40437 , n40272 , n40266 );
not ( n40438 , n40437 );
nand ( n40439 , n40436 , n40438 );
not ( n40440 , n40439 );
or ( n40441 , n40242 , n40440 );
not ( n40442 , n40232 );
not ( n40443 , n40224 );
or ( n40444 , n40442 , n40443 );
not ( n40445 , n40229 );
nand ( n40446 , n40444 , n40445 );
not ( n40447 , n40239 );
or ( n40448 , n40446 , n40447 );
or ( n40449 , n40237 , n40238 );
nand ( n40450 , n40448 , n40449 );
or ( n40451 , n40450 , n371 );
nand ( n40452 , n40451 , n370 );
nand ( n40453 , n40441 , n40452 );
buf ( n40454 , n40453 );
and ( n40455 , n40372 , n376 );
buf ( n40456 , n40455 );
and ( n40457 , n40454 , n40456 );
buf ( n40458 , n40457 );
buf ( n40459 , n40458 );
buf ( n40460 , n40424 );
buf ( n40461 , n40460 );
not ( n40462 , n40431 );
buf ( n40463 , n40326 );
nand ( n40464 , n40462 , n40463 );
not ( n40465 , n40464 );
and ( n40466 , n40461 , n40465 );
not ( n40467 , n40461 );
and ( n40468 , n40467 , n40464 );
nor ( n40469 , n40466 , n40468 );
buf ( n40470 , n40469 );
buf ( n40471 , n40470 );
buf ( n40472 , n40471 );
buf ( n40473 , n40472 );
and ( n40474 , n40459 , n40473 );
not ( n40475 , n40459 );
buf ( n40476 , n40472 );
not ( n40477 , n40476 );
buf ( n40478 , n40477 );
buf ( n40479 , n40478 );
and ( n40480 , n40475 , n40479 );
nor ( n40481 , n40474 , n40480 );
buf ( n40482 , n40481 );
not ( n40483 , n40447 );
nand ( n40484 , n40483 , n40449 );
not ( n40485 , n40484 );
not ( n40486 , n40273 );
not ( n40487 , n40233 );
nor ( n40488 , n40486 , n40487 );
not ( n40489 , n40488 );
buf ( n40490 , n40434 );
not ( n40491 , n40490 );
or ( n40492 , n40489 , n40491 );
and ( n40493 , n40437 , n40233 );
not ( n40494 , n40446 );
nor ( n40495 , n40493 , n40494 );
nand ( n40496 , n40492 , n40495 );
not ( n40497 , n40496 );
or ( n40498 , n40485 , n40497 );
or ( n40499 , n40484 , n40496 );
nand ( n40500 , n40498 , n40499 );
buf ( n40501 , n40500 );
not ( n40502 , n40501 );
buf ( n40503 , n40502 );
buf ( n40504 , n40503 );
not ( n40505 , n40504 );
buf ( n40506 , n40505 );
and ( n40507 , n40371 , n40406 );
not ( n40508 , n40371 );
and ( n40509 , n40508 , n40372 );
or ( n40510 , n40507 , n40509 );
nand ( n40511 , n40506 , n40510 );
buf ( n40512 , n40511 );
nand ( n40513 , n40228 , n370 );
not ( n40514 , n40513 );
not ( n40515 , n40514 );
nor ( n40516 , n40486 , n40240 );
not ( n40517 , n40516 );
not ( n40518 , n40434 );
or ( n40519 , n40517 , n40518 );
not ( n40520 , n40438 );
not ( n40521 , n40240 );
and ( n40522 , n40520 , n40521 );
nor ( n40523 , n40522 , n40450 );
nand ( n40524 , n40519 , n40523 );
not ( n40525 , n40524 );
not ( n40526 , n40525 );
or ( n40527 , n40515 , n40526 );
nand ( n40528 , n40524 , n40513 );
nand ( n40529 , n40527 , n40528 );
buf ( n40530 , n40529 );
not ( n40531 , n40530 );
buf ( n40532 , n40531 );
buf ( n40533 , n40532 );
not ( n40534 , n40533 );
buf ( n40535 , n40534 );
buf ( n40536 , n40535 );
buf ( n40537 , n40455 );
and ( n40538 , n40536 , n40537 );
xor ( n40539 , n40356 , n40366 );
xor ( n40540 , n40539 , n40414 );
nand ( n40541 , n40469 , n40540 );
buf ( n40542 , n40541 );
not ( n40543 , n40542 );
buf ( n40544 , n40543 );
buf ( n40545 , n40544 );
nor ( n40546 , n40538 , n40545 );
buf ( n40547 , n40546 );
buf ( n40548 , n40547 );
or ( n40549 , n40512 , n40548 );
buf ( n40550 , n40535 );
buf ( n40551 , n40544 );
buf ( n40552 , n40455 );
nand ( n40553 , n40550 , n40551 , n40552 );
buf ( n40554 , n40553 );
buf ( n40555 , n40554 );
nand ( n40556 , n40549 , n40555 );
buf ( n40557 , n40556 );
buf ( n40558 , n40557 );
not ( n40559 , n40558 );
buf ( n40560 , n40559 );
xor ( n40561 , n40482 , n40560 );
not ( n40562 , n40487 );
nand ( n40563 , n40562 , n40446 );
xnor ( n40564 , n40439 , n40563 );
buf ( n40565 , n40564 );
not ( n40566 , n40387 );
nand ( n40567 , n374 , n377 );
xor ( n40568 , n40567 , n375 );
nand ( n40569 , n40568 , n40386 );
nand ( n40570 , n40566 , n40569 );
and ( n40571 , n40570 , n40373 );
not ( n40572 , n40570 );
not ( n40573 , n40373 );
and ( n40574 , n40572 , n40573 );
or ( n40575 , n40571 , n40574 );
nand ( n40576 , n40565 , n40575 );
buf ( n40577 , n40576 );
not ( n40578 , n40577 );
not ( n40579 , n40486 );
nand ( n40580 , n40579 , n40438 );
not ( n40581 , n40580 );
not ( n40582 , n40581 );
not ( n40583 , n40490 );
not ( n40584 , n40583 );
or ( n40585 , n40582 , n40584 );
nand ( n40586 , n40490 , n40580 );
nand ( n40587 , n40585 , n40586 );
buf ( n40588 , n40587 );
not ( n40589 , n40588 );
buf ( n40590 , n40589 );
buf ( n40591 , n40590 );
not ( n40592 , n40591 );
buf ( n40593 , n40592 );
not ( n40594 , n40569 );
not ( n40595 , n40373 );
or ( n40596 , n40594 , n40595 );
nand ( n40597 , n40596 , n40566 );
not ( n40598 , n40597 );
not ( n40599 , n40598 );
not ( n40600 , n40389 );
nand ( n40601 , n40600 , n40384 );
not ( n40602 , n40601 );
not ( n40603 , n40602 );
or ( n40604 , n40599 , n40603 );
nand ( n40605 , n40601 , n40597 );
nand ( n40606 , n40604 , n40605 );
nand ( n40607 , n40593 , n40606 );
buf ( n40608 , n40607 );
not ( n40609 , n40608 );
or ( n40610 , n40578 , n40609 );
not ( n40611 , n40463 );
not ( n40612 , n40460 );
or ( n40613 , n40611 , n40612 );
not ( n40614 , n40431 );
nand ( n40615 , n40613 , n40614 );
not ( n40616 , n40615 );
and ( n40617 , n40304 , n40300 );
not ( n40618 , n40304 );
and ( n40619 , n40618 , n40301 );
nor ( n40620 , n40617 , n40619 );
not ( n40621 , n40620 );
and ( n40622 , n40616 , n40621 );
and ( n40623 , n40615 , n40620 );
nor ( n40624 , n40622 , n40623 );
not ( n40625 , n40624 );
nand ( n40626 , n40413 , n40408 );
xnor ( n40627 , n40391 , n40626 );
buf ( n40628 , n40627 );
buf ( n40629 , n40628 );
buf ( n40630 , n40629 );
nand ( n40631 , n40625 , n40630 );
buf ( n40632 , n40631 );
not ( n40633 , n40632 );
buf ( n40634 , n40633 );
buf ( n40635 , n40634 );
nand ( n40636 , n40610 , n40635 );
buf ( n40637 , n40636 );
buf ( n40638 , n40637 );
not ( n40639 , n40576 );
not ( n40640 , n40607 );
nand ( n40641 , n40639 , n40640 );
buf ( n40642 , n40641 );
nand ( n40643 , n40638 , n40642 );
buf ( n40644 , n40643 );
xnor ( n40645 , n40561 , n40644 );
buf ( n40646 , n40645 );
not ( n40647 , n40576 );
and ( n40648 , n40631 , n40647 );
not ( n40649 , n40631 );
and ( n40650 , n40649 , n40576 );
nor ( n40651 , n40648 , n40650 );
xor ( n40652 , n40640 , n40651 );
buf ( n40653 , n40652 );
not ( n40654 , n40653 );
nand ( n40655 , n40535 , n40455 );
xor ( n40656 , n40541 , n40655 );
xnor ( n40657 , n40656 , n40511 );
not ( n40658 , n40657 );
buf ( n40659 , n40658 );
not ( n40660 , n40659 );
or ( n40661 , n40654 , n40660 );
buf ( n40662 , n40453 );
buf ( n40663 , n40662 );
buf ( n40664 , n40663 );
buf ( n40665 , n40664 );
buf ( n40666 , n377 );
nand ( n40667 , n40665 , n40666 );
buf ( n40668 , n40667 );
and ( n40669 , n40421 , n40422 );
not ( n40670 , n40421 );
and ( n40671 , n40670 , n40352 );
nor ( n40672 , n40669 , n40671 );
not ( n40673 , n40672 );
buf ( n40674 , n40418 );
not ( n40675 , n40674 );
not ( n40676 , n40675 );
or ( n40677 , n40673 , n40676 );
not ( n40678 , n40672 );
nand ( n40679 , n40678 , n40674 );
nand ( n40680 , n40677 , n40679 );
buf ( n40681 , n40680 );
buf ( n40682 , n40681 );
buf ( n40683 , n40682 );
and ( n40684 , n40668 , n40683 );
not ( n40685 , n40668 );
buf ( n40686 , n40683 );
not ( n40687 , n40686 );
buf ( n40688 , n40687 );
and ( n40689 , n40685 , n40688 );
nor ( n40690 , n40684 , n40689 );
and ( n40691 , n40680 , n40630 );
not ( n40692 , n40514 );
not ( n40693 , n40525 );
or ( n40694 , n40692 , n40693 );
nand ( n40695 , n40694 , n40528 );
buf ( n40696 , n40695 );
nand ( n40697 , n40691 , n377 , n40696 );
nand ( n40698 , n40690 , n40697 );
not ( n40699 , n40698 );
buf ( n40700 , n40625 );
not ( n40701 , n40700 );
buf ( n40702 , n40575 );
not ( n40703 , n40702 );
buf ( n40704 , n40703 );
buf ( n40705 , n40704 );
nor ( n40706 , n40701 , n40705 );
buf ( n40707 , n40706 );
buf ( n40708 , n40707 );
buf ( n40709 , n40593 );
buf ( n40710 , n40510 );
and ( n40711 , n40709 , n40710 );
buf ( n40712 , n40711 );
buf ( n40713 , n40712 );
buf ( n40714 , n40565 );
buf ( n40715 , n40455 );
and ( n40716 , n40714 , n40715 );
buf ( n40717 , n40716 );
buf ( n40718 , n40717 );
and ( n40719 , n40708 , n40713 );
or ( n40720 , C0 , n40719 );
buf ( n40721 , n40720 );
not ( n40722 , n40721 );
or ( n40723 , n40699 , n40722 );
not ( n40724 , n40690 );
not ( n40725 , n40697 );
nand ( n40726 , n40724 , n40725 );
nand ( n40727 , n40723 , n40726 );
buf ( n40728 , n40727 );
nand ( n40729 , n40661 , n40728 );
buf ( n40730 , n40729 );
buf ( n40731 , n40730 );
not ( n40732 , n40652 );
nand ( n40733 , n40732 , n40657 );
buf ( n40734 , n40733 );
nand ( n40735 , n40731 , n40734 );
buf ( n40736 , n40735 );
buf ( n40737 , n40736 );
buf ( n40738 , n40469 );
not ( n40739 , n40672 );
not ( n40740 , n40675 );
or ( n40741 , n40739 , n40740 );
nand ( n40742 , n40741 , n40679 );
buf ( n40743 , n40742 );
nand ( n40744 , n40738 , n40743 );
buf ( n40745 , n40744 );
and ( n40746 , n40625 , n40540 );
xor ( n40747 , n40745 , n40746 );
buf ( n40748 , n40606 );
buf ( n40749 , n40565 );
nand ( n40750 , n40748 , n40749 );
buf ( n40751 , n40750 );
xnor ( n40752 , n40747 , n40751 );
not ( n40753 , n40752 );
buf ( n40754 , n40500 );
buf ( n40755 , n40575 );
and ( n40756 , n40754 , n40755 );
buf ( n40757 , n40756 );
buf ( n40758 , n40590 );
not ( n40759 , n40758 );
buf ( n40760 , n40759 );
buf ( n40761 , n40760 );
buf ( n40762 , n40627 );
and ( n40763 , n40761 , n40762 );
buf ( n40764 , n40763 );
xor ( n40765 , n40757 , n40764 );
buf ( n40766 , n40695 );
buf ( n40767 , n40510 );
and ( n40768 , n40766 , n40767 );
buf ( n40769 , n40768 );
xor ( n40770 , n40765 , n40769 );
not ( n40771 , n40770 );
or ( n40772 , n40753 , n40771 );
or ( n40773 , n40770 , n40752 );
nand ( n40774 , n40772 , n40773 );
buf ( n40775 , n40742 );
buf ( n40776 , n40540 );
nand ( n40777 , n40775 , n40776 );
buf ( n40778 , n40777 );
buf ( n40779 , n40778 );
not ( n40780 , n40779 );
buf ( n40781 , n40625 );
buf ( n40782 , n40606 );
nand ( n40783 , n40781 , n40782 );
buf ( n40784 , n40783 );
buf ( n40785 , n40784 );
not ( n40786 , n40785 );
or ( n40787 , n40780 , n40786 );
buf ( n40788 , n40469 );
buf ( n40789 , n40630 );
and ( n40790 , n40788 , n40789 );
buf ( n40791 , n40790 );
buf ( n40792 , n40791 );
nand ( n40793 , n40787 , n40792 );
buf ( n40794 , n40793 );
buf ( n40795 , n40794 );
buf ( n40796 , n40784 );
not ( n40797 , n40796 );
buf ( n40798 , n40778 );
not ( n40799 , n40798 );
buf ( n40800 , n40799 );
buf ( n40801 , n40800 );
nand ( n40802 , n40797 , n40801 );
buf ( n40803 , n40802 );
buf ( n40804 , n40803 );
nand ( n40805 , n40795 , n40804 );
buf ( n40806 , n40805 );
buf ( n40807 , n40806 );
buf ( n40808 , n40664 );
buf ( n40809 , n40683 );
buf ( n40810 , n377 );
and ( n40811 , n40808 , n40809 , n40810 );
buf ( n40812 , n40811 );
buf ( n40813 , n40812 );
xor ( n40814 , n40807 , n40813 );
buf ( n40815 , n40565 );
buf ( n40816 , n40510 );
nand ( n40817 , n40815 , n40816 );
buf ( n40818 , n40817 );
buf ( n40819 , n40818 );
not ( n40820 , n40819 );
buf ( n40821 , n40820 );
buf ( n40822 , n40821 );
not ( n40823 , n40822 );
buf ( n40824 , n40593 );
buf ( n40825 , n40575 );
and ( n40826 , n40824 , n40825 );
buf ( n40827 , n40826 );
buf ( n40828 , n40827 );
not ( n40829 , n40828 );
or ( n40830 , n40823 , n40829 );
buf ( n40831 , n40455 );
not ( n40832 , n40831 );
buf ( n40833 , n40832 );
buf ( n40834 , C1 );
buf ( n40835 , n40834 );
nand ( n40836 , n40830 , n40835 );
buf ( n40837 , n40836 );
buf ( n40838 , n40837 );
and ( n40839 , n40814 , n40838 );
and ( n40840 , n40807 , n40813 );
or ( n40841 , n40839 , n40840 );
buf ( n40842 , n40841 );
xor ( n40843 , n40774 , n40842 );
buf ( n40844 , n40843 );
xor ( n40845 , n40646 , n40737 );
xor ( n40846 , n40845 , n40844 );
buf ( n40847 , n40846 );
xor ( n40848 , n40646 , n40737 );
and ( n40849 , n40848 , n40844 );
and ( n40850 , n40646 , n40737 );
or ( n40851 , n40849 , n40850 );
buf ( n40852 , n40851 );
and ( n40853 , n40472 , n40664 , n40455 );
not ( n40854 , n40745 );
nand ( n40855 , n40854 , n40746 );
not ( n40856 , n40855 );
not ( n40857 , n40751 );
or ( n40858 , n40856 , n40857 );
not ( n40859 , n40746 );
nand ( n40860 , n40859 , n40745 );
nand ( n40861 , n40858 , n40860 );
xor ( n40862 , n40853 , n40861 );
xor ( n40863 , n40757 , n40764 );
and ( n40864 , n40863 , n40769 );
and ( n40865 , n40757 , n40764 );
or ( n40866 , n40864 , n40865 );
xnor ( n40867 , n40862 , n40866 );
buf ( n40868 , n40867 );
not ( n40869 , n40770 );
nand ( n40870 , n40869 , n40752 );
buf ( n40871 , n40870 );
not ( n40872 , n40871 );
buf ( n40873 , n40842 );
not ( n40874 , n40873 );
or ( n40875 , n40872 , n40874 );
not ( n40876 , n40752 );
nand ( n40877 , n40876 , n40770 );
buf ( n40878 , n40877 );
nand ( n40879 , n40875 , n40878 );
buf ( n40880 , n40879 );
buf ( n40881 , n40880 );
not ( n40882 , n40482 );
nand ( n40883 , n40882 , n40560 );
not ( n40884 , n40883 );
not ( n40885 , n40644 );
or ( n40886 , n40884 , n40885 );
not ( n40887 , n40560 );
nand ( n40888 , n40887 , n40482 );
nand ( n40889 , n40886 , n40888 );
buf ( n40890 , n40760 );
buf ( n40891 , n40540 );
and ( n40892 , n40890 , n40891 );
buf ( n40893 , n40892 );
buf ( n40894 , n40529 );
buf ( n40895 , n40575 );
and ( n40896 , n40894 , n40895 );
buf ( n40897 , n40896 );
xor ( n40898 , n40893 , n40897 );
buf ( n40899 , n40500 );
buf ( n40900 , n40606 );
and ( n40901 , n40899 , n40900 );
buf ( n40902 , n40901 );
xor ( n40903 , n40898 , n40902 );
buf ( n40904 , n40903 );
buf ( n40905 , n40625 );
buf ( n40906 , n40742 );
and ( n40907 , n40905 , n40906 );
buf ( n40908 , n40907 );
buf ( n40909 , n40908 );
not ( n40910 , n40452 );
nand ( n40911 , n40439 , n40241 );
not ( n40912 , n40911 );
or ( n40913 , n40910 , n40912 );
nand ( n40914 , n40913 , n40510 );
not ( n40915 , n40914 );
buf ( n40916 , n40915 );
xor ( n40917 , n40909 , n40916 );
buf ( n40918 , n40565 );
buf ( n40919 , n40630 );
and ( n40920 , n40918 , n40919 );
buf ( n40921 , n40920 );
buf ( n40922 , n40921 );
xor ( n40923 , n40917 , n40922 );
buf ( n40924 , n40923 );
buf ( n40925 , n40924 );
not ( n40926 , n40925 );
buf ( n40927 , n40926 );
buf ( n40928 , n40927 );
and ( n40929 , n40904 , n40928 );
not ( n40930 , n40904 );
buf ( n40931 , n40924 );
and ( n40932 , n40930 , n40931 );
nor ( n40933 , n40929 , n40932 );
buf ( n40934 , n40933 );
xnor ( n40935 , n40889 , n40934 );
buf ( n40936 , n40935 );
xor ( n40937 , n40868 , n40881 );
xor ( n40938 , n40937 , n40936 );
buf ( n40939 , n40938 );
xor ( n40940 , n40868 , n40881 );
and ( n40941 , n40940 , n40936 );
and ( n40942 , n40868 , n40881 );
or ( n40943 , n40941 , n40942 );
buf ( n40944 , n40943 );
not ( n40945 , n40727 );
and ( n40946 , n40652 , n40658 );
not ( n40947 , n40652 );
and ( n40948 , n40947 , n40657 );
nor ( n40949 , n40946 , n40948 );
xor ( n40950 , n40945 , n40949 );
not ( n40951 , n40950 );
xor ( n40952 , n40807 , n40813 );
xor ( n40953 , n40952 , n40838 );
buf ( n40954 , n40953 );
buf ( n40955 , n40954 );
not ( n40956 , n40955 );
buf ( n40957 , n40956 );
not ( n40958 , n40957 );
and ( n40959 , n40951 , n40958 );
buf ( n40960 , n40950 );
buf ( n40961 , n40957 );
nand ( n40962 , n40960 , n40961 );
buf ( n40963 , n40962 );
buf ( n40964 , n40800 );
buf ( n40965 , n40784 );
xor ( n40966 , n40964 , n40965 );
buf ( n40967 , n40791 );
xor ( n40968 , n40966 , n40967 );
buf ( n40969 , n40968 );
buf ( n40970 , n40969 );
not ( n40971 , n40970 );
buf ( n40972 , n40827 );
buf ( n40973 , n40821 );
and ( n40974 , n40972 , n40973 );
not ( n40975 , n40972 );
buf ( n40976 , n40818 );
and ( n40977 , n40975 , n40976 );
nor ( n40978 , n40974 , n40977 );
buf ( n40979 , n40978 );
buf ( n40980 , n40506 );
buf ( n40981 , n40455 );
and ( n40982 , n40980 , n40981 );
buf ( n40983 , n40982 );
xnor ( n40984 , n40979 , n40983 );
buf ( n40985 , n40984 );
not ( n40986 , n40985 );
buf ( n40987 , n40986 );
buf ( n40988 , n40987 );
nand ( n40989 , n40971 , n40988 );
buf ( n40990 , n40989 );
buf ( n40991 , n40990 );
buf ( n40992 , n40969 );
not ( n40993 , n40992 );
buf ( n40994 , n40984 );
not ( n40995 , n40994 );
or ( n40996 , n40993 , n40995 );
buf ( n40997 , n40469 );
buf ( n40998 , n40997 );
buf ( n40999 , n40998 );
buf ( n41000 , n40999 );
buf ( n41001 , n40606 );
and ( n41002 , n41000 , n41001 );
buf ( n41003 , n41002 );
buf ( n41004 , n41003 );
buf ( n41005 , n40500 );
buf ( n41006 , n41005 );
buf ( n41007 , n41006 );
buf ( n41008 , n41007 );
not ( n41009 , n41008 );
buf ( n41010 , n40540 );
buf ( n41011 , n41010 );
buf ( n41012 , n41011 );
buf ( n41013 , n41012 );
buf ( n41014 , n377 );
nand ( n41015 , n41013 , n41014 );
buf ( n41016 , n41015 );
buf ( n41017 , n41016 );
nor ( n41018 , n41009 , n41017 );
buf ( n41019 , n41018 );
buf ( n41020 , n41019 );
xor ( n41021 , n41004 , n41020 );
nand ( n41022 , n377 , n40695 );
xnor ( n41023 , n41022 , n40691 );
buf ( n41024 , n41023 );
and ( n41025 , n41021 , n41024 );
and ( n41026 , n41004 , n41020 );
or ( n41027 , n41025 , n41026 );
buf ( n41028 , n41027 );
buf ( n41029 , n41028 );
nand ( n41030 , n40996 , n41029 );
buf ( n41031 , n41030 );
buf ( n41032 , n41031 );
nand ( n41033 , n40991 , n41032 );
buf ( n41034 , n41033 );
and ( n41035 , n40963 , n41034 );
nor ( n41036 , n40959 , n41035 );
buf ( n41037 , n41036 );
not ( n41038 , n41037 );
buf ( n41039 , n41038 );
xor ( n41040 , n40708 , n40713 );
xor ( n41041 , n41040 , n40718 );
buf ( n41042 , n41041 );
buf ( n41043 , n41042 );
buf ( n41044 , n40540 );
buf ( n41045 , n40627 );
and ( n41046 , n41044 , n41045 );
buf ( n41047 , n41046 );
buf ( n41048 , n41047 );
buf ( n41049 , n40625 );
buf ( n41050 , n40510 );
and ( n41051 , n41049 , n41050 );
buf ( n41052 , n41051 );
buf ( n41053 , n41052 );
xor ( n41054 , n41048 , n41053 );
buf ( n41055 , n40760 );
buf ( n41056 , n40455 );
and ( n41057 , n41055 , n41056 );
buf ( n41058 , n41057 );
buf ( n41059 , n41058 );
and ( n41060 , n41054 , n41059 );
and ( n41061 , n41048 , n41053 );
or ( n41062 , n41060 , n41061 );
buf ( n41063 , n41062 );
buf ( n41064 , n41063 );
xor ( n41065 , n41043 , n41064 );
buf ( n41066 , n40742 );
buf ( n41067 , n40606 );
and ( n41068 , n41066 , n41067 );
buf ( n41069 , n41068 );
buf ( n41070 , n41069 );
buf ( n41071 , n40999 );
not ( n41072 , n41071 );
buf ( n41073 , n40704 );
nor ( n41074 , n41072 , n41073 );
buf ( n41075 , n41074 );
buf ( n41076 , n41075 );
xor ( n41077 , n41070 , n41076 );
buf ( n41078 , n40565 );
buf ( n41079 , n41078 );
buf ( n41080 , n377 );
nand ( n41081 , n41079 , n41080 );
buf ( n41082 , n41081 );
buf ( n41083 , n41082 );
buf ( n41084 , n40540 );
buf ( n41085 , n40606 );
nand ( n41086 , n41084 , n41085 );
buf ( n41087 , n41086 );
buf ( n41088 , n41087 );
nor ( n41089 , n41083 , n41088 );
buf ( n41090 , n41089 );
buf ( n41091 , n41090 );
and ( n41092 , n41077 , n41091 );
and ( n41093 , n41070 , n41076 );
or ( n41094 , n41092 , n41093 );
buf ( n41095 , n41094 );
buf ( n41096 , n41095 );
and ( n41097 , n41065 , n41096 );
and ( n41098 , n41043 , n41064 );
or ( n41099 , n41097 , n41098 );
buf ( n41100 , n41099 );
buf ( n41101 , n41100 );
buf ( n41102 , n40725 );
not ( n41103 , n41102 );
buf ( n41104 , n40690 );
not ( n41105 , n41104 );
or ( n41106 , n41103 , n41105 );
buf ( n41107 , n40725 );
buf ( n41108 , n40690 );
or ( n41109 , n41107 , n41108 );
nand ( n41110 , n41106 , n41109 );
buf ( n41111 , n41110 );
xor ( n41112 , n40721 , n41111 );
buf ( n41113 , n41112 );
buf ( n41114 , n40969 );
buf ( n41115 , n40987 );
xor ( n41116 , n41114 , n41115 );
buf ( n41117 , n41028 );
xnor ( n41118 , n41116 , n41117 );
buf ( n41119 , n41118 );
buf ( n41120 , n41119 );
xor ( n41121 , n41101 , n41113 );
xor ( n41122 , n41121 , n41120 );
buf ( n41123 , n41122 );
xor ( n41124 , n41101 , n41113 );
and ( n41125 , n41124 , n41120 );
and ( n41126 , n41101 , n41113 );
or ( n41127 , n41125 , n41126 );
buf ( n41128 , n41127 );
buf ( n41129 , n40950 );
buf ( n41130 , n40950 );
not ( n41131 , n41130 );
buf ( n41132 , n41131 );
buf ( n41133 , n41132 );
buf ( n41134 , n41034 );
buf ( n41135 , n40954 );
and ( n41136 , n41134 , n41135 );
not ( n41137 , n41134 );
buf ( n41138 , n40957 );
and ( n41139 , n41137 , n41138 );
nor ( n41140 , n41136 , n41139 );
buf ( n41141 , n41140 );
buf ( n41142 , n41141 );
and ( n41143 , n41142 , n41133 );
not ( n41144 , n41142 );
and ( n41145 , n41144 , n41129 );
nor ( n41146 , n41143 , n41145 );
buf ( n41147 , n41146 );
buf ( n41148 , n41078 );
buf ( n41149 , n40664 );
buf ( n41150 , n40683 );
nand ( n41151 , n41149 , n41150 );
buf ( n41152 , n41151 );
buf ( n41153 , n41152 );
xor ( n41154 , n41148 , n41153 );
buf ( n41155 , n40593 );
buf ( n41156 , n41155 );
buf ( n41157 , n41156 );
buf ( n41158 , n41157 );
buf ( n41159 , n41078 );
and ( n41160 , n41158 , n41159 );
buf ( n41161 , n41160 );
buf ( n41162 , n41161 );
xnor ( n41163 , n41154 , n41162 );
buf ( n41164 , n41163 );
buf ( n41165 , n41164 );
buf ( n41166 , n40696 );
buf ( n41167 , n40472 );
and ( n41168 , n41166 , n41167 );
buf ( n41169 , n41168 );
buf ( n41170 , n41169 );
buf ( n41171 , n40506 );
buf ( n41172 , n40624 );
not ( n41173 , n41172 );
buf ( n41174 , n41173 );
and ( n41175 , n41171 , n41174 );
buf ( n41176 , n41175 );
buf ( n41177 , n41176 );
xor ( n41178 , n41170 , n41177 );
buf ( n41179 , n40664 );
buf ( n41180 , n41012 );
nand ( n41181 , n41179 , n41180 );
buf ( n41182 , n41181 );
buf ( n41183 , n41182 );
not ( n41184 , n41183 );
buf ( n41185 , n40565 );
buf ( n41186 , n41173 );
nand ( n41187 , n41185 , n41186 );
buf ( n41188 , n41187 );
buf ( n41189 , n41188 );
not ( n41190 , n41189 );
or ( n41191 , n41184 , n41190 );
buf ( n41192 , n40696 );
not ( n41193 , n41192 );
buf ( n41194 , n40688 );
nor ( n41195 , n41193 , n41194 );
buf ( n41196 , n41195 );
buf ( n41197 , n41196 );
nand ( n41198 , n41191 , n41197 );
buf ( n41199 , n41198 );
buf ( n41200 , n41199 );
or ( n41201 , n41182 , n41188 );
buf ( n41202 , n41201 );
nand ( n41203 , n41200 , n41202 );
buf ( n41204 , n41203 );
buf ( n41205 , n41204 );
xor ( n41206 , n41178 , n41205 );
buf ( n41207 , n41206 );
buf ( n41208 , n41207 );
buf ( n41209 , n40506 );
buf ( n41210 , n40683 );
and ( n41211 , n41209 , n41210 );
buf ( n41212 , n41211 );
not ( n41213 , n41212 );
buf ( n41214 , n40535 );
buf ( n41215 , n40540 );
nand ( n41216 , n41214 , n41215 );
buf ( n41217 , n41216 );
buf ( n41218 , n41217 );
buf ( n41219 , n40593 );
buf ( n41220 , n40625 );
and ( n41221 , n41219 , n41220 );
buf ( n41222 , n41221 );
buf ( n41223 , n41222 );
not ( n41224 , n41223 );
buf ( n41225 , n41224 );
buf ( n41226 , n41225 );
nand ( n41227 , n41218 , n41226 );
buf ( n41228 , n41227 );
not ( n41229 , n41228 );
or ( n41230 , n41213 , n41229 );
buf ( n41231 , n40696 );
buf ( n41232 , n41012 );
nand ( n41233 , n41231 , n41232 );
buf ( n41234 , n41233 );
not ( n41235 , n41234 );
nand ( n41236 , n41235 , n41222 );
nand ( n41237 , n41230 , n41236 );
not ( n41238 , n41237 );
buf ( n41239 , n40506 );
not ( n41240 , n41239 );
buf ( n41241 , n40478 );
nor ( n41242 , n41240 , n41241 );
buf ( n41243 , n41242 );
not ( n41244 , n41243 );
or ( n41245 , n41238 , n41244 );
buf ( n41246 , n41243 );
not ( n41247 , n41246 );
buf ( n41248 , n41247 );
not ( n41249 , n41248 );
buf ( n41250 , n41237 );
not ( n41251 , n41250 );
buf ( n41252 , n41251 );
not ( n41253 , n41252 );
or ( n41254 , n41249 , n41253 );
buf ( n41255 , n41157 );
not ( n41256 , n41255 );
buf ( n41257 , n40469 );
not ( n41258 , n41257 );
buf ( n41259 , n41258 );
buf ( n41260 , n41259 );
not ( n41261 , n41260 );
buf ( n41262 , n40565 );
nand ( n41263 , n41261 , n41262 );
buf ( n41264 , n41263 );
buf ( n41265 , n41264 );
not ( n41266 , n41265 );
buf ( n41267 , n41266 );
buf ( n41268 , n41267 );
not ( n41269 , n41268 );
or ( n41270 , n41256 , n41269 );
buf ( n41271 , n41264 );
not ( n41272 , n41271 );
buf ( n41273 , n40593 );
not ( n41274 , n41273 );
buf ( n41275 , n41274 );
buf ( n41276 , n41275 );
not ( n41277 , n41276 );
or ( n41278 , n41272 , n41277 );
buf ( n41279 , n40453 );
buf ( n41280 , n40630 );
and ( n41281 , n41279 , n41280 );
buf ( n41282 , n41281 );
buf ( n41283 , n41282 );
nand ( n41284 , n41278 , n41283 );
buf ( n41285 , n41284 );
buf ( n41286 , n41285 );
nand ( n41287 , n41270 , n41286 );
buf ( n41288 , n41287 );
nand ( n41289 , n41254 , n41288 );
nand ( n41290 , n41245 , n41289 );
buf ( n41291 , n41290 );
xor ( n41292 , n41165 , n41208 );
xor ( n41293 , n41292 , n41291 );
buf ( n41294 , n41293 );
xor ( n41295 , n41165 , n41208 );
and ( n41296 , n41295 , n41291 );
and ( n41297 , n41165 , n41208 );
or ( n41298 , n41296 , n41297 );
buf ( n41299 , n41298 );
xor ( n41300 , n41070 , n41076 );
xor ( n41301 , n41300 , n41091 );
buf ( n41302 , n41301 );
buf ( n41303 , n41302 );
buf ( n41304 , n40627 );
buf ( n41305 , n40606 );
and ( n41306 , n41304 , n41305 );
buf ( n41307 , n41306 );
buf ( n41308 , n41307 );
buf ( n41309 , n40680 );
not ( n41310 , n41309 );
buf ( n41311 , n40510 );
not ( n41312 , n41311 );
buf ( n41313 , n41312 );
buf ( n41314 , n41313 );
nor ( n41315 , n41310 , n41314 );
buf ( n41316 , n41315 );
buf ( n41317 , n41316 );
xor ( n41318 , n41308 , n41317 );
buf ( n41319 , n40999 );
not ( n41320 , n41319 );
buf ( n41321 , n40833 );
nor ( n41322 , n41320 , n41321 );
buf ( n41323 , n41322 );
buf ( n41324 , n41323 );
and ( n41325 , n41318 , n41324 );
and ( n41326 , n41308 , n41317 );
or ( n41327 , n41325 , n41326 );
buf ( n41328 , n41327 );
buf ( n41329 , n41328 );
xor ( n41330 , n41087 , n41082 );
buf ( n41331 , n41330 );
xor ( n41332 , n41329 , n41331 );
buf ( n41333 , n40630 );
buf ( n41334 , n377 );
not ( n41335 , n41334 );
buf ( n41336 , n41275 );
nor ( n41337 , n41335 , n41336 );
buf ( n41338 , n41337 );
buf ( n41339 , n41338 );
and ( n41340 , n41333 , n41339 );
buf ( n41341 , n41340 );
buf ( n41342 , n41341 );
and ( n41343 , n41332 , n41342 );
and ( n41344 , n41329 , n41331 );
or ( n41345 , n41343 , n41344 );
buf ( n41346 , n41345 );
buf ( n41347 , n41346 );
buf ( n41348 , n40680 );
buf ( n41349 , n40575 );
nand ( n41350 , n41348 , n41349 );
buf ( n41351 , n41350 );
buf ( n41352 , n41351 );
not ( n41353 , n41352 );
buf ( n41354 , n40625 );
buf ( n41355 , n40455 );
nand ( n41356 , n41354 , n41355 );
buf ( n41357 , n41356 );
buf ( n41358 , n41357 );
not ( n41359 , n41358 );
or ( n41360 , n41353 , n41359 );
buf ( n41361 , n40999 );
buf ( n41362 , n40510 );
and ( n41363 , n41361 , n41362 );
buf ( n41364 , n41363 );
buf ( n41365 , n41364 );
nand ( n41366 , n41360 , n41365 );
buf ( n41367 , n41366 );
buf ( n41368 , n41367 );
buf ( n41369 , n41351 );
not ( n41370 , n41369 );
buf ( n41371 , n41370 );
buf ( n41372 , C1 );
buf ( n41373 , n41372 );
nand ( n41374 , n41368 , n41373 );
buf ( n41375 , n41374 );
buf ( n41376 , n41375 );
xor ( n41377 , n41048 , n41053 );
xor ( n41378 , n41377 , n41059 );
buf ( n41379 , n41378 );
buf ( n41380 , n41379 );
xor ( n41381 , n41376 , n41380 );
buf ( n41382 , n41007 );
buf ( n41383 , n377 );
nand ( n41384 , n41382 , n41383 );
buf ( n41385 , n41384 );
xnor ( n41386 , n41012 , n41385 );
buf ( n41387 , n41386 );
xor ( n41388 , n41381 , n41387 );
buf ( n41389 , n41388 );
buf ( n41390 , n41389 );
xor ( n41391 , n41303 , n41347 );
xor ( n41392 , n41391 , n41390 );
buf ( n41393 , n41392 );
xor ( n41394 , n41303 , n41347 );
and ( n41395 , n41394 , n41390 );
and ( n41396 , n41303 , n41347 );
or ( n41397 , n41395 , n41396 );
buf ( n41398 , n41397 );
xnor ( n41399 , n41364 , n41371 );
buf ( n41400 , n41399 );
buf ( n41401 , n41357 );
and ( n41402 , n41400 , n41401 );
nor ( n41403 , n41402 , C0 );
buf ( n41404 , n41403 );
buf ( n41405 , n41404 );
buf ( n41406 , n41012 );
buf ( n41407 , n40575 );
and ( n41408 , n41406 , n41407 );
buf ( n41409 , n41408 );
buf ( n41410 , n41409 );
nand ( n41411 , n41173 , n377 );
buf ( n41412 , n41411 );
buf ( n41413 , n40630 );
buf ( n41414 , n40575 );
nand ( n41415 , n41413 , n41414 );
buf ( n41416 , n41415 );
buf ( n41417 , n41416 );
nor ( n41418 , n41412 , n41417 );
buf ( n41419 , n41418 );
buf ( n41420 , n41419 );
xor ( n41421 , n41410 , n41420 );
xor ( n41422 , n41333 , n41339 );
buf ( n41423 , n41422 );
buf ( n41424 , n41423 );
and ( n41425 , n41421 , n41424 );
and ( n41426 , n41410 , n41420 );
or ( n41427 , n41425 , n41426 );
buf ( n41428 , n41427 );
buf ( n41429 , n41428 );
xor ( n41430 , n41329 , n41331 );
xor ( n41431 , n41430 , n41342 );
buf ( n41432 , n41431 );
buf ( n41433 , n41432 );
xor ( n41434 , n41405 , n41429 );
xor ( n41435 , n41434 , n41433 );
buf ( n41436 , n41435 );
xor ( n41437 , n41405 , n41429 );
and ( n41438 , n41437 , n41433 );
and ( n41439 , n41405 , n41429 );
or ( n41440 , n41438 , n41439 );
buf ( n41441 , n41440 );
xor ( n41442 , n41043 , n41064 );
xor ( n41443 , n41442 , n41096 );
buf ( n41444 , n41443 );
buf ( n41445 , n41173 );
buf ( n41446 , n40472 );
and ( n41447 , n41445 , n41446 );
buf ( n41448 , n41447 );
buf ( n41449 , n41448 );
xor ( n41450 , n40893 , n40897 );
and ( n41451 , n41450 , n40902 );
and ( n41452 , n40893 , n40897 );
or ( n41453 , n41451 , n41452 );
buf ( n41454 , n41453 );
xor ( n41455 , n40909 , n40916 );
and ( n41456 , n41455 , n40922 );
and ( n41457 , n40909 , n40916 );
or ( n41458 , n41456 , n41457 );
buf ( n41459 , n41458 );
buf ( n41460 , n41459 );
xor ( n41461 , n41449 , n41454 );
xor ( n41462 , n41461 , n41460 );
buf ( n41463 , n41462 );
xor ( n41464 , n41449 , n41454 );
and ( n41465 , n41464 , n41460 );
and ( n41466 , n41449 , n41454 );
or ( n41467 , n41465 , n41466 );
buf ( n41468 , n41467 );
xor ( n41469 , n41308 , n41317 );
xor ( n41470 , n41469 , n41324 );
buf ( n41471 , n41470 );
buf ( n41472 , n41471 );
buf ( n41473 , n41012 );
buf ( n41474 , n40510 );
and ( n41475 , n41473 , n41474 );
buf ( n41476 , n41475 );
buf ( n41477 , n41476 );
buf ( n41478 , n40683 );
buf ( n41479 , n40455 );
and ( n41480 , n41478 , n41479 );
buf ( n41481 , n41480 );
buf ( n41482 , n41481 );
xor ( n41483 , n41477 , n41482 );
buf ( n41484 , n40472 );
buf ( n41485 , n377 );
nand ( n41486 , n41484 , n41485 );
buf ( n41487 , n41486 );
buf ( n41488 , n41487 );
buf ( n41489 , n40606 );
not ( n41490 , n41489 );
buf ( n41491 , n41490 );
buf ( n41492 , n41491 );
nor ( n41493 , n41488 , n41492 );
buf ( n41494 , n41493 );
buf ( n41495 , n41494 );
and ( n41496 , n41483 , n41495 );
or ( n41497 , n41496 , C0 );
buf ( n41498 , n41497 );
buf ( n41499 , n41498 );
xor ( n41500 , n41410 , n41420 );
xor ( n41501 , n41500 , n41424 );
buf ( n41502 , n41501 );
buf ( n41503 , n41502 );
xor ( n41504 , n41472 , n41499 );
xor ( n41505 , n41504 , n41503 );
buf ( n41506 , n41505 );
xor ( n41507 , n41472 , n41499 );
and ( n41508 , n41507 , n41503 );
and ( n41509 , n41472 , n41499 );
or ( n41510 , n41508 , n41509 );
buf ( n41511 , n41510 );
buf ( n41512 , n40506 );
not ( n41513 , n41512 );
buf ( n41514 , n41513 );
buf ( n41515 , n41514 );
not ( n41516 , n41078 );
buf ( n41517 , n41516 );
nor ( n41518 , n41515 , n41517 );
buf ( n41519 , n41518 );
buf ( n41520 , n41519 );
buf ( n41521 , n40664 );
buf ( n41522 , n40472 );
and ( n41523 , n41521 , n41522 );
buf ( n41524 , n41523 );
buf ( n41525 , n41524 );
buf ( n41526 , n40506 );
not ( n41527 , n41526 );
buf ( n41528 , n41275 );
nor ( n41529 , n41527 , n41528 );
buf ( n41530 , n41529 );
buf ( n41531 , n41530 );
xor ( n41532 , n41525 , n41531 );
buf ( n41533 , n40696 );
buf ( n41534 , n41173 );
and ( n41535 , n41533 , n41534 );
buf ( n41536 , n41535 );
buf ( n41537 , n41536 );
and ( n41538 , n41532 , n41537 );
and ( n41539 , n41525 , n41531 );
or ( n41540 , n41538 , n41539 );
buf ( n41541 , n41540 );
buf ( n41542 , n41541 );
buf ( n41543 , n40664 );
buf ( n41544 , n41173 );
and ( n41545 , n41543 , n41544 );
buf ( n41546 , n41545 );
buf ( n41547 , n41546 );
buf ( n41548 , n41514 );
not ( n41549 , n41548 );
buf ( n41550 , n41549 );
buf ( n41551 , n41550 );
xor ( n41552 , n41547 , n41551 );
buf ( n41553 , n40696 );
buf ( n41554 , n41157 );
and ( n41555 , n41553 , n41554 );
buf ( n41556 , n41555 );
buf ( n41557 , n41556 );
xor ( n41558 , n41552 , n41557 );
buf ( n41559 , n41558 );
buf ( n41560 , n41559 );
xor ( n41561 , n41520 , n41542 );
xor ( n41562 , n41561 , n41560 );
buf ( n41563 , n41562 );
xor ( n41564 , n41520 , n41542 );
and ( n41565 , n41564 , n41560 );
and ( n41566 , n41520 , n41542 );
or ( n41567 , n41565 , n41566 );
buf ( n41568 , n41567 );
buf ( n41569 , n41078 );
not ( n41570 , n41569 );
buf ( n41571 , n41152 );
not ( n41572 , n41571 );
buf ( n41573 , n41572 );
buf ( n41574 , n41573 );
not ( n41575 , n41574 );
or ( n41576 , n41570 , n41575 );
buf ( n41577 , n41161 );
not ( n41578 , n41577 );
buf ( n41579 , n41578 );
buf ( n41580 , n41579 );
nand ( n41581 , n41576 , n41580 );
buf ( n41582 , n41581 );
buf ( n41583 , n41582 );
xor ( n41584 , n41525 , n41531 );
xor ( n41585 , n41584 , n41537 );
buf ( n41586 , n41585 );
buf ( n41587 , n41586 );
xor ( n41588 , n41170 , n41177 );
and ( n41589 , n41588 , n41205 );
and ( n41590 , n41170 , n41177 );
or ( n41591 , n41589 , n41590 );
buf ( n41592 , n41591 );
buf ( n41593 , n41592 );
xor ( n41594 , n41583 , n41587 );
xor ( n41595 , n41594 , n41593 );
buf ( n41596 , n41595 );
xor ( n41597 , n41583 , n41587 );
and ( n41598 , n41597 , n41593 );
and ( n41599 , n41583 , n41587 );
or ( n41600 , n41598 , n41599 );
buf ( n41601 , n41600 );
buf ( n41602 , n40903 );
not ( n41603 , n41602 );
buf ( n41604 , n40927 );
nand ( n41605 , n41603 , n41604 );
buf ( n41606 , n41605 );
buf ( n41607 , n41606 );
buf ( n41608 , n40889 );
nand ( n41609 , n40924 , n40903 );
buf ( n41610 , n41609 );
not ( n41611 , n41607 );
not ( n41612 , n41608 );
or ( n41613 , n41611 , n41612 );
nand ( n41614 , n41613 , n41610 );
buf ( n41615 , n41614 );
xor ( n41616 , n41376 , n41380 );
and ( n41617 , n41616 , n41387 );
and ( n41618 , n41376 , n41380 );
or ( n41619 , n41617 , n41618 );
buf ( n41620 , n41619 );
buf ( n41621 , n41012 );
buf ( n41622 , n40455 );
nand ( n41623 , n41621 , n41622 );
buf ( n41624 , n41623 );
buf ( n41625 , n41624 );
buf ( n41626 , n40630 );
buf ( n41627 , n40510 );
nand ( n41628 , n41626 , n41627 );
buf ( n41629 , n41628 );
buf ( n41630 , n41629 );
nand ( n41631 , n41625 , n41630 );
buf ( n41632 , n41631 );
not ( n41633 , n41632 );
buf ( n41634 , n40606 );
buf ( n41635 , n40575 );
and ( n41636 , n41634 , n41635 );
buf ( n41637 , n41636 );
not ( n41638 , n41637 );
or ( n41639 , n41633 , n41638 );
nand ( n41640 , n41639 , C1 );
buf ( n41641 , n41640 );
xor ( n41642 , n41416 , n41411 );
buf ( n41643 , n41642 );
xor ( n41644 , n41477 , n41482 );
xor ( n41645 , n41644 , n41495 );
buf ( n41646 , n41645 );
buf ( n41647 , n41646 );
xor ( n41648 , n41641 , n41643 );
xor ( n41649 , n41648 , n41647 );
buf ( n41650 , n41649 );
xor ( n41651 , n41641 , n41643 );
and ( n41652 , n41651 , n41647 );
and ( n41653 , n41641 , n41643 );
or ( n41654 , n41652 , n41653 );
buf ( n41655 , n41654 );
xor ( n41656 , n41188 , n41182 );
xor ( n41657 , n41656 , n41196 );
buf ( n41658 , n41657 );
and ( n41659 , n41288 , n41243 );
not ( n41660 , n41288 );
or ( n41661 , n41514 , n40478 );
and ( n41662 , n41660 , n41661 );
nor ( n41663 , n41659 , n41662 );
buf ( n41664 , n41663 );
not ( n41665 , n41664 );
buf ( n41666 , n41252 );
not ( n41667 , n41666 );
and ( n41668 , n41665 , n41667 );
buf ( n41669 , n41252 );
buf ( n41670 , n41663 );
and ( n41671 , n41669 , n41670 );
nor ( n41672 , n41668 , n41671 );
buf ( n41673 , n41672 );
buf ( n41674 , n41673 );
nand ( n41675 , n41658 , n41674 );
buf ( n41676 , n41675 );
buf ( n41677 , n41624 );
not ( n41678 , n41677 );
buf ( n41679 , n41637 );
not ( n41680 , n41679 );
buf ( n41681 , n41629 );
not ( n41682 , n41681 );
or ( n41683 , n41680 , n41682 );
buf ( n41684 , n41629 );
buf ( n41685 , n41637 );
or ( n41686 , n41684 , n41685 );
nand ( n41687 , n41683 , n41686 );
buf ( n41688 , n41687 );
buf ( n41689 , n41688 );
not ( n41690 , n41689 );
or ( n41691 , n41678 , n41690 );
buf ( n41692 , n41688 );
buf ( n41693 , n41624 );
or ( n41694 , n41692 , n41693 );
nand ( n41695 , n41691 , n41694 );
buf ( n41696 , n41695 );
buf ( n41697 , n41696 );
buf ( n41698 , n40606 );
buf ( n41699 , n40510 );
and ( n41700 , n41698 , n41699 );
buf ( n41701 , n41700 );
buf ( n41702 , n41701 );
buf ( n41703 , n40683 );
buf ( n41704 , n377 );
and ( n41705 , n41703 , n41704 );
buf ( n41706 , n41705 );
buf ( n41707 , n41706 );
and ( n41708 , n41702 , n41707 );
buf ( n41709 , n41708 );
buf ( n41710 , n41709 );
buf ( n41711 , n41487 );
buf ( n41712 , n41491 );
and ( n41713 , n41711 , n41712 );
not ( n41714 , n41711 );
buf ( n41715 , n40606 );
and ( n41716 , n41714 , n41715 );
nor ( n41717 , n41713 , n41716 );
buf ( n41718 , n41717 );
buf ( n41719 , n41718 );
xor ( n41720 , n41697 , n41710 );
xor ( n41721 , n41720 , n41719 );
buf ( n41722 , n41721 );
xor ( n41723 , n41697 , n41710 );
and ( n41724 , n41723 , n41719 );
and ( n41725 , n41697 , n41710 );
or ( n41726 , n41724 , n41725 );
buf ( n41727 , n41726 );
buf ( n41728 , n402 );
buf ( n41729 , n40627 );
buf ( n41730 , n377 );
and ( n41731 , n41729 , n41730 );
buf ( n41732 , n41731 );
buf ( n41733 , n41732 );
and ( n41734 , n41728 , n41733 );
buf ( n41735 , n41734 );
buf ( n41736 , n41735 );
buf ( n41737 , n40606 );
buf ( n41738 , n40455 );
and ( n41739 , n41737 , n41738 );
buf ( n41740 , n41739 );
buf ( n41741 , n41740 );
buf ( n41742 , n40575 );
buf ( n41743 , n40575 );
buf ( n41744 , n40510 );
nand ( n41745 , n41743 , n41744 );
buf ( n41746 , n41745 );
buf ( n41747 , n41746 );
xor ( n41748 , n41742 , n41747 );
buf ( n41749 , n41016 );
xor ( n41750 , n41748 , n41749 );
buf ( n41751 , n41750 );
buf ( n41752 , n41751 );
xor ( n41753 , n41736 , n41741 );
xor ( n41754 , n41753 , n41752 );
buf ( n41755 , n41754 );
xor ( n41756 , n41736 , n41741 );
and ( n41757 , n41756 , n41752 );
or ( n41758 , n41757 , C0 );
buf ( n41759 , n41758 );
buf ( n41760 , n40630 );
buf ( n41761 , n40455 );
and ( n41762 , n41760 , n41761 );
buf ( n41763 , n41762 );
buf ( n41764 , n41763 );
buf ( n41765 , n41016 );
not ( n41766 , n41765 );
buf ( n41767 , n40575 );
nand ( n41768 , n41766 , n41767 );
buf ( n41769 , n41768 );
buf ( n41770 , n41769 );
buf ( n41771 , n41746 );
nand ( n41772 , n41770 , n41771 );
buf ( n41773 , n41772 );
buf ( n41774 , n41773 );
xor ( n41775 , n41702 , n41707 );
buf ( n41776 , n41775 );
buf ( n41777 , n41776 );
xor ( n41778 , n41764 , n41774 );
xor ( n41779 , n41778 , n41777 );
buf ( n41780 , n41779 );
xor ( n41781 , n41764 , n41774 );
and ( n41782 , n41781 , n41777 );
or ( n41783 , n41782 , C0 );
buf ( n41784 , n41783 );
buf ( n41785 , n40696 );
buf ( n41786 , n41078 );
and ( n41787 , n41785 , n41786 );
buf ( n41788 , n41787 );
buf ( n41789 , n41788 );
buf ( n41790 , n41157 );
buf ( n41791 , n40664 );
and ( n41792 , n41790 , n41791 );
buf ( n41793 , n41792 );
buf ( n41794 , n41793 );
xor ( n41795 , n41547 , n41551 );
and ( n41796 , n41795 , n41557 );
and ( n41797 , n41547 , n41551 );
or ( n41798 , n41796 , n41797 );
buf ( n41799 , n41798 );
buf ( n41800 , n41799 );
xor ( n41801 , n41789 , n41794 );
xor ( n41802 , n41801 , n41800 );
buf ( n41803 , n41802 );
xor ( n41804 , n41789 , n41794 );
and ( n41805 , n41804 , n41800 );
and ( n41806 , n41789 , n41794 );
or ( n41807 , n41805 , n41806 );
buf ( n41808 , n41807 );
xor ( n41809 , n41004 , n41020 );
xor ( n41810 , n41809 , n41024 );
buf ( n41811 , n41810 );
buf ( n41812 , n40453 );
buf ( n41813 , n40606 );
and ( n41814 , n41812 , n41813 );
buf ( n41815 , n41814 );
buf ( n41816 , n41815 );
buf ( n41817 , n40593 );
buf ( n41818 , n40999 );
and ( n41819 , n41817 , n41818 );
buf ( n41820 , n41819 );
buf ( n41821 , n41820 );
xor ( n41822 , n41816 , n41821 );
buf ( n41823 , n40565 );
buf ( n41824 , n40680 );
and ( n41825 , n41823 , n41824 );
buf ( n41826 , n41825 );
buf ( n41827 , n41826 );
xor ( n41828 , n41822 , n41827 );
buf ( n41829 , n41828 );
buf ( n41830 , n41829 );
not ( n41831 , n41830 );
buf ( n41832 , n41831 );
buf ( n41833 , n41832 );
buf ( n41834 , n41173 );
buf ( n41835 , n40453 );
buf ( n41836 , n40575 );
and ( n41837 , n41835 , n41836 );
buf ( n41838 , n41837 );
buf ( n41839 , n41838 );
xor ( n41840 , n41834 , n41839 );
buf ( n41841 , n40565 );
buf ( n41842 , n40540 );
and ( n41843 , n41841 , n41842 );
buf ( n41844 , n41843 );
buf ( n41845 , n41844 );
and ( n41846 , n41840 , n41845 );
and ( n41847 , n41834 , n41839 );
or ( n41848 , n41846 , n41847 );
buf ( n41849 , n41848 );
buf ( n41850 , n41849 );
buf ( n41851 , n41832 );
buf ( n41852 , n41849 );
not ( n41853 , n41833 );
not ( n41854 , n41850 );
and ( n41855 , n41853 , n41854 );
and ( n41856 , n41851 , n41852 );
nor ( n41857 , n41855 , n41856 );
buf ( n41858 , n41857 );
buf ( n41859 , n41657 );
not ( n41860 , n41859 );
buf ( n41861 , n41860 );
and ( n41862 , n40760 , n40742 );
buf ( n41863 , n41862 );
buf ( n41864 , n40529 );
buf ( n41865 , n40606 );
and ( n41866 , n41864 , n41865 );
buf ( n41867 , n41866 );
buf ( n41868 , n41867 );
buf ( n41869 , n40506 );
buf ( n41870 , n40630 );
and ( n41871 , n41869 , n41870 );
buf ( n41872 , n41871 );
buf ( n41873 , n41872 );
xor ( n41874 , n41863 , n41868 );
xor ( n41875 , n41874 , n41873 );
buf ( n41876 , n41875 );
xor ( n41877 , n41863 , n41868 );
and ( n41878 , n41877 , n41873 );
and ( n41879 , n41863 , n41868 );
or ( n41880 , n41878 , n41879 );
buf ( n41881 , n41880 );
buf ( n41882 , n41832 );
buf ( n41883 , n41849 );
not ( n41884 , n41883 );
buf ( n41885 , n41884 );
buf ( n41886 , n41885 );
nand ( n41887 , n41882 , n41886 );
buf ( n41888 , n41887 );
xor ( n41889 , n41816 , n41821 );
and ( n41890 , n41889 , n41827 );
and ( n41891 , n41816 , n41821 );
or ( n41892 , n41890 , n41891 );
buf ( n41893 , n41892 );
buf ( n41894 , n40696 );
buf ( n41895 , n41516 );
not ( n41896 , n41895 );
buf ( n41897 , n40664 );
nand ( n41898 , n41896 , n41897 );
buf ( n41899 , n41898 );
buf ( n41900 , n41899 );
not ( n41901 , n41900 );
buf ( n41902 , n41901 );
buf ( n41903 , n41902 );
buf ( n41904 , n41550 );
buf ( n41905 , n40696 );
nand ( n41906 , n41904 , n41905 );
buf ( n41907 , n41906 );
buf ( n41908 , n41907 );
not ( n41909 , n41894 );
not ( n41910 , n41903 );
or ( n41911 , n41909 , n41910 );
nand ( n41912 , n41911 , n41908 );
buf ( n41913 , n41912 );
xor ( n41914 , n41728 , n41733 );
buf ( n41915 , n41914 );
buf ( n41916 , n404 );
buf ( n41917 , n40575 );
buf ( n41918 , n377 );
and ( n41919 , n41917 , n41918 );
buf ( n41920 , n41919 );
buf ( n41921 , n41920 );
xor ( n41922 , n41916 , n41921 );
buf ( n41923 , n41922 );
and ( n41924 , n41916 , n41921 );
buf ( n41925 , n41924 );
buf ( n41926 , n405 );
buf ( n41927 , n40455 );
xor ( n41928 , n41926 , n41927 );
buf ( n41929 , n41928 );
and ( n41930 , n41926 , n41927 );
buf ( n41931 , n41930 );
buf ( n41932 , n403 );
buf ( n41933 , n40510 );
xor ( n41934 , n41932 , n41933 );
buf ( n41935 , n41934 );
and ( n41936 , n41932 , n41933 );
buf ( n41937 , n41936 );
buf ( n41938 , n41222 );
buf ( n41939 , n41217 );
buf ( n41940 , n41234 );
buf ( n41941 , n41222 );
not ( n41942 , n41938 );
not ( n41943 , n41939 );
or ( n41944 , n41942 , n41943 );
or ( n41945 , n41940 , n41941 );
nand ( n41946 , n41944 , n41945 );
buf ( n41947 , n41946 );
buf ( n41948 , n41550 );
buf ( n41949 , n40664 );
and ( n41950 , n41948 , n41949 );
buf ( n41951 , n41950 );
buf ( n41952 , n40606 );
buf ( n41953 , n377 );
and ( n41954 , n41952 , n41953 );
buf ( n41955 , n41954 );
buf ( n41956 , n40696 );
buf ( n41957 , n40630 );
and ( n41958 , n41956 , n41957 );
buf ( n41959 , n41958 );
buf ( n41960 , n41550 );
buf ( n41961 , n41012 );
and ( n41962 , n41960 , n41961 );
buf ( n41963 , n41962 );
buf ( n41964 , n41832 );
buf ( n41965 , n41885 );
or ( n41966 , n41964 , n41965 );
buf ( n41967 , n41966 );
buf ( n41968 , n41157 );
buf ( n41969 , n41282 );
buf ( n41970 , n41267 );
xor ( n41971 , n41968 , n41969 );
xor ( n41972 , n41971 , n41970 );
buf ( n41973 , n41972 );
buf ( n41974 , n377 );
buf ( n41975 , n41313 );
not ( n41976 , n41974 );
nor ( n41977 , n41976 , n41975 );
buf ( n41978 , n41977 );
not ( n41979 , n41959 );
xor ( n41980 , n41979 , n41963 );
xnor ( n41981 , n41980 , n41881 );
not ( n41982 , n40853 );
nand ( n41983 , n41982 , n40861 );
not ( n41984 , n41983 );
not ( n41985 , n40866 );
or ( n41986 , n41984 , n41985 );
not ( n41987 , n40861 );
nand ( n41988 , n41987 , n40853 );
nand ( n41989 , n41986 , n41988 );
not ( n41990 , n41989 );
xor ( n41991 , n41834 , n41839 );
xor ( n41992 , n41991 , n41845 );
buf ( n41993 , n41992 );
not ( n41994 , n41993 );
not ( n41995 , n41876 );
nand ( n41996 , n41994 , n41995 );
not ( n41997 , n41996 );
or ( n41998 , n41990 , n41997 );
not ( n41999 , n41995 );
nand ( n42000 , n41999 , n41993 );
nand ( n42001 , n41998 , n42000 );
xor ( n42002 , n41981 , n42001 );
not ( n42003 , n41858 );
not ( n42004 , n42003 );
not ( n42005 , n41468 );
not ( n42006 , n42005 );
or ( n42007 , n42004 , n42006 );
nand ( n42008 , n41468 , n41858 );
nand ( n42009 , n42007 , n42008 );
xor ( n42010 , n42002 , n42009 );
buf ( n42011 , n42010 );
not ( n42012 , n41615 );
not ( n42013 , n41463 );
nand ( n42014 , n42012 , n42013 );
not ( n42015 , n42014 );
xor ( n42016 , n41994 , n41999 );
xnor ( n42017 , n42016 , n41989 );
not ( n42018 , n42017 );
or ( n42019 , n42015 , n42018 );
nand ( n42020 , n41615 , n41463 );
nand ( n42021 , n42019 , n42020 );
buf ( n42022 , n42021 );
nor ( n42023 , n42011 , n42022 );
buf ( n42024 , n42023 );
buf ( n42025 , n42024 );
not ( n42026 , n42025 );
not ( n42027 , n41861 );
not ( n42028 , n41673 );
not ( n42029 , n42028 );
or ( n42030 , n42027 , n42029 );
nand ( n42031 , n42030 , n41676 );
xor ( n42032 , n41893 , n41973 );
xor ( n42033 , n41947 , n41212 );
and ( n42034 , n42032 , n42033 );
and ( n42035 , n41893 , n41973 );
or ( n42036 , n42034 , n42035 );
xor ( n42037 , n42031 , n42036 );
not ( n42038 , n41959 );
not ( n42039 , n41963 );
or ( n42040 , n42038 , n42039 );
not ( n42041 , n41979 );
not ( n42042 , n41963 );
not ( n42043 , n42042 );
or ( n42044 , n42041 , n42043 );
nand ( n42045 , n42044 , n41881 );
nand ( n42046 , n42040 , n42045 );
xor ( n42047 , n41893 , n41973 );
xor ( n42048 , n42047 , n42033 );
xor ( n42049 , n42046 , n42048 );
not ( n42050 , n41888 );
not ( n42051 , n41468 );
or ( n42052 , n42050 , n42051 );
nand ( n42053 , n42052 , n41967 );
and ( n42054 , n42049 , n42053 );
and ( n42055 , n42046 , n42048 );
or ( n42056 , n42054 , n42055 );
nor ( n42057 , n42037 , n42056 );
buf ( n42058 , n42057 );
not ( n42059 , n42058 );
not ( n42060 , n40944 );
not ( n42061 , n41463 );
not ( n42062 , n42012 );
or ( n42063 , n42061 , n42062 );
nand ( n42064 , n41615 , n42013 );
nand ( n42065 , n42063 , n42064 );
and ( n42066 , n42065 , n42017 );
not ( n42067 , n42065 );
not ( n42068 , n42017 );
and ( n42069 , n42067 , n42068 );
nor ( n42070 , n42066 , n42069 );
not ( n42071 , n42070 );
nand ( n42072 , n42060 , n42071 );
buf ( n42073 , n42072 );
xor ( n42074 , n42046 , n42048 );
xor ( n42075 , n42074 , n42053 );
buf ( n42076 , n42075 );
not ( n42077 , n42076 );
buf ( n42078 , n41981 );
or ( n42079 , n42009 , n42078 );
buf ( n42080 , n42001 );
and ( n42081 , n42079 , n42080 );
and ( n42082 , n42009 , n42078 );
nor ( n42083 , n42081 , n42082 );
buf ( n42084 , n42083 );
nand ( n42085 , n42077 , n42084 );
buf ( n42086 , n42085 );
buf ( n42087 , n42086 );
nand ( n42088 , n42026 , n42059 , n42073 , n42087 );
buf ( n42089 , n42088 );
buf ( n42090 , n42089 );
buf ( n42091 , n41299 );
not ( n42092 , n42091 );
buf ( n42093 , n42092 );
buf ( n42094 , n42093 );
buf ( n42095 , n41596 );
not ( n42096 , n42095 );
buf ( n42097 , n42096 );
buf ( n42098 , n42097 );
or ( n42099 , n42094 , n42098 );
buf ( n42100 , n42099 );
not ( n42101 , n42100 );
not ( n42102 , n42028 );
not ( n42103 , n41657 );
or ( n42104 , n42102 , n42103 );
not ( n42105 , n41861 );
not ( n42106 , n41673 );
or ( n42107 , n42105 , n42106 );
nand ( n42108 , n42107 , n42036 );
nand ( n42109 , n42104 , n42108 );
buf ( n42110 , n42109 );
buf ( n42111 , n41294 );
nand ( n42112 , n42110 , n42111 );
buf ( n42113 , n42112 );
buf ( n42114 , n42113 );
not ( n42115 , n42114 );
buf ( n42116 , n42093 );
buf ( n42117 , n42097 );
nand ( n42118 , n42116 , n42117 );
buf ( n42119 , n42118 );
buf ( n42120 , n42119 );
nand ( n42121 , n42115 , n42120 );
buf ( n42122 , n42121 );
not ( n42123 , n42122 );
or ( n42124 , n42101 , n42123 );
or ( n42125 , n41803 , n41568 );
not ( n42126 , n41563 );
not ( n42127 , n41601 );
nand ( n42128 , n42126 , n42127 );
nand ( n42129 , n42125 , n42128 );
not ( n42130 , n42129 );
nand ( n42131 , n42124 , n42130 );
buf ( n42132 , n42131 );
nand ( n42133 , n41601 , n41563 );
not ( n42134 , n42125 );
or ( n42135 , n42133 , n42134 );
nand ( n42136 , n41803 , n41568 );
nand ( n42137 , n42135 , n42136 );
buf ( n42138 , n42137 );
xor ( n42139 , n41907 , n40696 );
xor ( n42140 , n42139 , n41899 );
nand ( n42141 , n41808 , n42140 );
buf ( n42142 , n42141 );
buf ( n42143 , n41913 );
buf ( n42144 , n41951 );
nor ( n42145 , n42143 , n42144 );
buf ( n42146 , n42145 );
buf ( n42147 , n42146 );
or ( n42148 , n42142 , n42147 );
buf ( n42149 , n41913 );
buf ( n42150 , n41951 );
nand ( n42151 , n42149 , n42150 );
buf ( n42152 , n42151 );
buf ( n42153 , n42152 );
nand ( n42154 , n42148 , n42153 );
buf ( n42155 , n42154 );
buf ( n42156 , n42155 );
nor ( n42157 , n42138 , n42156 );
buf ( n42158 , n42157 );
buf ( n42159 , n42158 );
nand ( n42160 , n42090 , n42132 , n42159 );
buf ( n42161 , n42160 );
buf ( n42162 , n42161 );
buf ( n42163 , n40852 );
not ( n42164 , n42163 );
buf ( n42165 , n40939 );
not ( n42166 , n42165 );
and ( n42167 , n42164 , n42166 );
buf ( n42168 , n40847 );
not ( n42169 , n42168 );
buf ( n42170 , n42169 );
buf ( n42171 , n42170 );
buf ( n42172 , n41039 );
not ( n42173 , n42172 );
buf ( n42174 , n42173 );
buf ( n42175 , n42174 );
and ( n42176 , n42171 , n42175 );
nor ( n42177 , n42167 , n42176 );
buf ( n42178 , n42177 );
buf ( n42179 , n41147 );
buf ( n42180 , n41128 );
nor ( n42181 , n42179 , n42180 );
buf ( n42182 , n42181 );
buf ( n42183 , n42182 );
buf ( n42184 , n41123 );
xor ( n42185 , n41811 , n41620 );
and ( n42186 , n42185 , n41444 );
and ( n42187 , n41811 , n41620 );
or ( n42188 , n42186 , n42187 );
buf ( n42189 , n42188 );
nor ( n42190 , n42184 , n42189 );
buf ( n42191 , n42190 );
buf ( n42192 , n42191 );
nor ( n42193 , n42183 , n42192 );
buf ( n42194 , n42193 );
nand ( n42195 , n42178 , n42194 );
nand ( n42196 , n42195 , n42131 , n42158 );
buf ( n42197 , n42196 );
buf ( n42198 , n42155 );
not ( n42199 , n42198 );
buf ( n42200 , n42146 );
not ( n42201 , n42200 );
buf ( n42202 , n41808 );
buf ( n42203 , n42140 );
or ( n42204 , n42202 , n42203 );
buf ( n42205 , n42204 );
buf ( n42206 , n42205 );
nand ( n42207 , n42201 , n42206 );
buf ( n42208 , n42207 );
buf ( n42209 , n42208 );
nand ( n42210 , n42199 , n42209 );
buf ( n42211 , n42210 );
buf ( n42212 , n42211 );
and ( n42213 , n42162 , n42197 , n42212 );
buf ( n42214 , n42213 );
buf ( n42215 , n42214 );
not ( n42216 , n41398 );
xor ( n42217 , n41811 , n41620 );
xor ( n42218 , n42217 , n41444 );
not ( n42219 , n42218 );
and ( n42220 , n42216 , n42219 );
nor ( n42221 , n41393 , n41441 );
nor ( n42222 , n42220 , n42221 );
not ( n42223 , n42222 );
buf ( n42224 , n41436 );
buf ( n42225 , n41511 );
nor ( n42226 , n42224 , n42225 );
buf ( n42227 , n42226 );
buf ( n42228 , n41506 );
buf ( n42229 , n41655 );
nand ( n42230 , n42228 , n42229 );
buf ( n42231 , n42230 );
or ( n42232 , n42227 , n42231 );
buf ( n42233 , n41436 );
buf ( n42234 , n41511 );
nand ( n42235 , n42233 , n42234 );
buf ( n42236 , n42235 );
nand ( n42237 , n42232 , n42236 );
not ( n42238 , n42237 );
or ( n42239 , n42223 , n42238 );
not ( n42240 , n42218 );
not ( n42241 , n41398 );
nand ( n42242 , n42240 , n42241 );
and ( n42243 , n41393 , n41441 );
and ( n42244 , n42242 , n42243 );
buf ( n42245 , n42218 );
buf ( n42246 , n41398 );
and ( n42247 , n42245 , n42246 );
buf ( n42248 , n42247 );
nor ( n42249 , n42244 , n42248 );
nand ( n42250 , n42239 , n42249 );
buf ( n42251 , n42250 );
buf ( n42252 , n42158 );
not ( n42253 , n42252 );
buf ( n42254 , n42253 );
buf ( n42255 , n42254 );
nor ( n42256 , n42251 , n42255 );
buf ( n42257 , n42256 );
buf ( n42258 , n42257 );
not ( n42259 , n42227 );
not ( n42260 , n42259 );
buf ( n42261 , n41506 );
buf ( n42262 , n41655 );
nor ( n42263 , n42261 , n42262 );
buf ( n42264 , n42263 );
buf ( n42265 , n42264 );
nor ( n42266 , n42260 , n42265 );
buf ( n42267 , n41780 );
buf ( n42268 , n41759 );
nor ( n42269 , n42267 , n42268 );
buf ( n42270 , n42269 );
buf ( n42271 , n42270 );
buf ( n42272 , n41755 );
and ( n42273 , n41937 , n41915 );
buf ( n42274 , n42273 );
nand ( n42275 , n42272 , n42274 );
buf ( n42276 , n42275 );
buf ( n42277 , n42276 );
or ( n42278 , n42271 , n42277 );
buf ( n42279 , n41780 );
buf ( n42280 , n41759 );
nand ( n42281 , n42279 , n42280 );
buf ( n42282 , n42281 );
buf ( n42283 , n42282 );
nand ( n42284 , n42278 , n42283 );
buf ( n42285 , n42284 );
not ( n42286 , n42285 );
buf ( n42287 , n41650 );
buf ( n42288 , n41727 );
nor ( n42289 , n42287 , n42288 );
buf ( n42290 , n42289 );
buf ( n42291 , n42290 );
buf ( n42292 , n41722 );
buf ( n42293 , n41784 );
nor ( n42294 , n42292 , n42293 );
buf ( n42295 , n42294 );
buf ( n42296 , n42295 );
nor ( n42297 , n42291 , n42296 );
buf ( n42298 , n42297 );
not ( n42299 , n42298 );
or ( n42300 , n42286 , n42299 );
buf ( n42301 , n42290 );
not ( n42302 , n42301 );
buf ( n42303 , n42302 );
buf ( n42304 , n42303 );
buf ( n42305 , n41784 );
buf ( n42306 , n41722 );
and ( n42307 , n42305 , n42306 );
buf ( n42308 , n42307 );
buf ( n42309 , n42308 );
and ( n42310 , n42304 , n42309 );
buf ( n42311 , n41650 );
buf ( n42312 , n41727 );
and ( n42313 , n42311 , n42312 );
nor ( n42314 , n42310 , n42313 );
buf ( n42315 , n42314 );
nand ( n42316 , n42300 , n42315 );
nand ( n42317 , n42222 , n42266 , n42316 );
buf ( n42318 , n42317 );
buf ( n42319 , n42131 );
nor ( n42320 , n42227 , n42265 );
not ( n42321 , n42295 );
or ( n42322 , n41755 , n42273 );
or ( n42323 , n41780 , n41759 );
xor ( n42324 , n41935 , n41955 );
buf ( n42325 , n42324 );
not ( n42326 , n42325 );
buf ( n42327 , n41925 );
not ( n42328 , n42327 );
and ( n42329 , n42326 , n42328 );
xor ( n42330 , n41937 , n41915 );
buf ( n42331 , n42330 );
and ( n42332 , n41935 , n41955 );
buf ( n42333 , n42332 );
nor ( n42334 , n42331 , n42333 );
buf ( n42335 , n42334 );
buf ( n42336 , n42335 );
nor ( n42337 , n42329 , n42336 );
buf ( n42338 , n42337 );
buf ( n42339 , n42338 );
buf ( n42340 , n41923 );
buf ( n42341 , n41931 );
nor ( n42342 , n42340 , n42341 );
buf ( n42343 , n42342 );
buf ( n42344 , n42343 );
buf ( n42345 , n406 );
not ( n42346 , n42345 );
and ( n42347 , C1 , n42346 );
buf ( n42348 , n407 );
buf ( n42349 , n408 );
buf ( n42350 , n377 );
buf ( n42351 , n409 );
nand ( n42352 , n42348 , n42349 , n42350 , n42351 );
buf ( n42353 , n42352 );
buf ( n42354 , n42353 );
nor ( n42355 , n42347 , n42354 );
buf ( n42356 , n42355 );
buf ( n42357 , n42356 );
nor ( n42358 , C0 , n42357 );
buf ( n42359 , n42358 );
buf ( n42360 , n42359 );
buf ( n42361 , n41978 );
buf ( n42362 , n41929 );
nor ( n42363 , n42361 , n42362 );
buf ( n42364 , n42363 );
buf ( n42365 , n42364 );
nor ( n42366 , n42344 , n42360 , n42365 );
buf ( n42367 , n42366 );
buf ( n42368 , n42367 );
nand ( n42369 , n42339 , n42368 );
buf ( n42370 , n42369 );
buf ( n42371 , n42370 );
buf ( n42372 , n42343 );
not ( n42373 , n42372 );
buf ( n42374 , n42373 );
buf ( n42375 , n42374 );
buf ( n42376 , n41978 );
buf ( n42377 , n41929 );
and ( n42378 , n42375 , n42376 , n42377 );
buf ( n42379 , n41923 );
buf ( n42380 , n41931 );
and ( n42381 , n42379 , n42380 );
nor ( n42382 , n42378 , n42381 );
buf ( n42383 , n42382 );
buf ( n42384 , n42383 );
not ( n42385 , n42384 );
buf ( n42386 , n42338 );
nand ( n42387 , n42385 , n42386 );
buf ( n42388 , n42387 );
buf ( n42389 , n42388 );
buf ( n42390 , n42335 );
not ( n42391 , n42390 );
buf ( n42392 , n42391 );
buf ( n42393 , n42392 );
buf ( n42394 , n42324 );
buf ( n42395 , n41925 );
and ( n42396 , n42393 , n42394 , n42395 );
buf ( n42397 , n42330 );
buf ( n42398 , n42332 );
and ( n42399 , n42397 , n42398 );
nor ( n42400 , n42396 , n42399 );
buf ( n42401 , n42400 );
buf ( n42402 , n42401 );
nand ( n42403 , n42371 , n42389 , n42402 );
buf ( n42404 , n42403 );
nand ( n42405 , n42322 , n42323 , n42404 );
nor ( n42406 , n42405 , n42290 );
nand ( n42407 , n42321 , n42406 );
nor ( n42408 , n42221 , n42407 );
nand ( n42409 , n42320 , n42408 , n42242 );
buf ( n42410 , n42409 );
nand ( n42411 , n42258 , n42318 , n42319 , n42410 );
buf ( n42412 , n42411 );
buf ( n42413 , n42412 );
buf ( n42414 , n42131 );
buf ( n42415 , n42109 );
buf ( n42416 , n41294 );
or ( n42417 , n42415 , n42416 );
buf ( n42418 , n42417 );
buf ( n42419 , n42418 );
buf ( n42420 , n42119 );
nand ( n42421 , n42419 , n42420 );
buf ( n42422 , n42421 );
buf ( n42423 , n42422 );
buf ( n42424 , n42129 );
nor ( n42425 , n42423 , n42424 );
buf ( n42426 , n42425 );
buf ( n42427 , n42426 );
buf ( n42428 , n42254 );
nor ( n42429 , n42427 , n42428 );
buf ( n42430 , n42429 );
buf ( n42431 , n42430 );
nand ( n42432 , n42414 , n42431 );
buf ( n42433 , n42432 );
buf ( n42434 , n42433 );
and ( n42435 , n42413 , n42434 );
buf ( n42436 , n42435 );
buf ( n42437 , n42436 );
nand ( n42438 , n42215 , n42437 );
buf ( n42439 , n42438 );
not ( n42440 , n42250 );
and ( n42441 , n42266 , n42408 , n42242 );
not ( n42442 , n42137 );
nand ( n42443 , n42442 , n42141 );
nor ( n42444 , n42441 , n42443 );
nand ( n42445 , n42131 , n42440 , n42317 , n42444 );
buf ( n42446 , n42445 );
buf ( n42447 , n42122 );
not ( n42448 , n42447 );
buf ( n42449 , n42448 );
buf ( n42450 , n42449 );
not ( n42451 , n42450 );
buf ( n42452 , n42136 );
buf ( n42453 , n42141 );
and ( n42454 , n42452 , n42453 );
buf ( n42455 , n42454 );
buf ( n42456 , n42455 );
buf ( n42457 , n42100 );
buf ( n42458 , n42133 );
nand ( n42459 , n42456 , n42457 , n42458 );
buf ( n42460 , n42459 );
buf ( n42461 , n42460 );
not ( n42462 , n42461 );
and ( n42463 , n42451 , n42462 );
buf ( n42464 , n42129 );
buf ( n42465 , n42455 );
and ( n42466 , n42464 , n42465 );
nor ( n42467 , n42463 , n42466 );
buf ( n42468 , n42467 );
buf ( n42469 , n42468 );
not ( n42470 , n42469 );
buf ( n42471 , n42426 );
not ( n42472 , n42471 );
and ( n42473 , n42470 , n42472 );
buf ( n42474 , n42024 );
not ( n42475 , n42474 );
buf ( n42476 , n42057 );
not ( n42477 , n42476 );
buf ( n42478 , n42072 );
buf ( n42479 , n42086 );
nand ( n42480 , n42475 , n42477 , n42478 , n42479 );
buf ( n42481 , n42480 );
buf ( n42482 , n42481 );
buf ( n42483 , n42468 );
not ( n42484 , n42483 );
buf ( n42485 , n42484 );
buf ( n42486 , n42485 );
and ( n42487 , n42482 , n42486 );
nor ( n42488 , n42473 , n42487 );
buf ( n42489 , n42488 );
buf ( n42490 , n42489 );
and ( n42491 , n42485 , n42195 );
buf ( n42492 , n42205 );
not ( n42493 , n42492 );
buf ( n42494 , n42493 );
nor ( n42495 , n42491 , n42494 );
buf ( n42496 , n42495 );
nand ( n42497 , n42446 , n42490 , n42496 );
buf ( n42498 , n42497 );
buf ( n42499 , n42418 );
buf ( n42500 , n42089 );
not ( n42501 , n42500 );
buf ( n42502 , n42501 );
not ( n42503 , n42502 );
buf ( n42504 , n41147 );
buf ( n42505 , n41128 );
nand ( n42506 , n42504 , n42505 );
buf ( n42507 , n42506 );
nand ( n42508 , n41123 , n42188 );
and ( n42509 , n42507 , n42508 );
nor ( n42510 , n42509 , n42182 );
buf ( n42511 , n42510 );
not ( n42512 , n42511 );
buf ( n42513 , n42178 );
not ( n42514 , n42513 );
or ( n42515 , n42512 , n42514 );
buf ( n42516 , n40852 );
not ( n42517 , n42516 );
buf ( n42518 , n40939 );
not ( n42519 , n42518 );
buf ( n42520 , n42519 );
buf ( n42521 , n42520 );
nand ( n42522 , n42517 , n42521 );
buf ( n42523 , n42522 );
buf ( n42524 , n42523 );
buf ( n42525 , n40847 );
buf ( n42526 , n41039 );
and ( n42527 , n42525 , n42526 );
buf ( n42528 , n42527 );
buf ( n42529 , n42528 );
and ( n42530 , n42524 , n42529 );
buf ( n42531 , n42520 );
not ( n42532 , n42531 );
buf ( n42533 , n42532 );
buf ( n42534 , n42533 );
buf ( n42535 , n40852 );
and ( n42536 , n42534 , n42535 );
nor ( n42537 , n42530 , n42536 );
buf ( n42538 , n42537 );
buf ( n42539 , n42538 );
nand ( n42540 , n42515 , n42539 );
buf ( n42541 , n42540 );
not ( n42542 , n42541 );
or ( n42543 , n42503 , n42542 );
buf ( n42544 , n42057 );
not ( n42545 , n42544 );
buf ( n42546 , n42545 );
nand ( n42547 , n42546 , n42086 );
not ( n42548 , n42547 );
not ( n42549 , n42024 );
buf ( n42550 , n40944 );
not ( n42551 , n42550 );
buf ( n42552 , n42070 );
not ( n42553 , n42552 );
or ( n42554 , n42551 , n42553 );
buf ( n42555 , n42010 );
buf ( n42556 , n42021 );
nand ( n42557 , n42555 , n42556 );
buf ( n42558 , n42557 );
buf ( n42559 , n42558 );
nand ( n42560 , n42554 , n42559 );
buf ( n42561 , n42560 );
nand ( n42562 , n42549 , n42561 );
not ( n42563 , n42562 );
and ( n42564 , n42548 , n42563 );
not ( n42565 , n42057 );
not ( n42566 , n42565 );
and ( n42567 , n42079 , n42080 );
nor ( n42568 , n42567 , n42082 );
not ( n42569 , n42075 );
nor ( n42570 , n42568 , n42569 );
not ( n42571 , n42570 );
or ( n42572 , n42566 , n42571 );
nand ( n42573 , n42037 , n42056 );
nand ( n42574 , n42572 , n42573 );
nor ( n42575 , n42564 , n42574 );
nand ( n42576 , n42543 , n42575 );
buf ( n42577 , n42576 );
nand ( n42578 , n42499 , n42577 );
buf ( n42579 , n42578 );
buf ( n42580 , n42579 );
nand ( n42581 , n42440 , n42409 , n42317 );
buf ( n42582 , n42581 );
buf ( n42583 , n42582 );
buf ( n42584 , n42178 );
not ( n42585 , n42584 );
buf ( n42586 , n42182 );
buf ( n42587 , n42191 );
or ( n42588 , n42586 , n42587 );
buf ( n42589 , n42588 );
buf ( n42590 , n42589 );
nor ( n42591 , n42585 , n42590 );
buf ( n42592 , n42591 );
and ( n42593 , n42502 , n42592 );
buf ( n42594 , n42593 );
buf ( n42595 , n42418 );
nand ( n42596 , n42583 , n42594 , n42595 );
buf ( n42597 , n42596 );
buf ( n42598 , n42597 );
buf ( n42599 , n42113 );
nand ( n42600 , n42580 , n42598 , n42599 );
buf ( n42601 , n42600 );
buf ( n42602 , n42582 );
not ( n42603 , n42072 );
buf ( n42604 , n42024 );
nor ( n42605 , n42603 , n42604 );
not ( n42606 , n42605 );
nor ( n42607 , n42606 , n42195 );
buf ( n42608 , n42607 );
nand ( n42609 , n42602 , n42608 );
buf ( n42610 , n42609 );
buf ( n42611 , C1 );
buf ( n42612 , n42426 );
not ( n42613 , n42612 );
buf ( n42614 , n42613 );
buf ( n42615 , n42614 );
buf ( n42616 , n42208 );
not ( n42617 , n42616 );
buf ( n42618 , n40664 );
nand ( n42619 , n42617 , n42618 );
buf ( n42620 , n42619 );
buf ( n42621 , n42620 );
nor ( n42622 , n42615 , n42621 );
buf ( n42623 , n42622 );
buf ( n42624 , C1 );
buf ( n42625 , n42576 );
not ( n42626 , n42422 );
buf ( n42627 , n42626 );
nand ( n42628 , n42625 , n42627 );
buf ( n42629 , n42628 );
buf ( n42630 , n42576 );
buf ( n42631 , n42426 );
nand ( n42632 , n42630 , n42631 );
buf ( n42633 , n42632 );
not ( n42634 , n42502 );
not ( n42635 , n42541 );
or ( n42636 , n42634 , n42635 );
nand ( n42637 , n42636 , n42575 );
buf ( n42638 , n42637 );
buf ( n42639 , n42623 );
nand ( n42640 , n42638 , n42639 );
buf ( n42641 , n42640 );
buf ( n42642 , n42576 );
not ( n42643 , n42642 );
buf ( n42644 , n42643 );
not ( n42645 , n42604 );
not ( n42646 , n42072 );
not ( n42647 , n42086 );
nor ( n42648 , n42646 , n42647 );
nand ( n42649 , n42645 , n42648 );
not ( n42650 , n42649 );
buf ( n42651 , n42650 );
buf ( n42652 , n42541 );
or ( n42653 , n42647 , n42562 );
not ( n42654 , n42570 );
nand ( n42655 , n42653 , n42654 );
buf ( n42656 , n42655 );
and ( n42657 , n42651 , n42652 );
nor ( n42658 , n42657 , n42656 );
buf ( n42659 , n42658 );
buf ( n42660 , n42137 );
not ( n42661 , n42660 );
buf ( n42662 , n42131 );
nand ( n42663 , n42661 , n42662 );
buf ( n42664 , n42663 );
buf ( n42665 , n42664 );
buf ( n42666 , n42620 );
not ( n42667 , n42666 );
buf ( n42668 , n42667 );
buf ( n42669 , n42668 );
buf ( n42670 , n40664 );
not ( n42671 , n42670 );
buf ( n42672 , n42155 );
not ( n42673 , n42672 );
or ( n42674 , n42671 , n42673 );
nand ( n42675 , n40696 , n40664 );
buf ( n42676 , n42675 );
nand ( n42677 , n42674 , n42676 );
buf ( n42678 , n42677 );
buf ( n42679 , n42678 );
and ( n42680 , n42665 , n42669 );
nor ( n42681 , n42680 , n42679 );
buf ( n42682 , n42681 );
buf ( n42683 , n42614 );
buf ( n42684 , n42208 );
nor ( n42685 , n42683 , n42684 );
buf ( n42686 , n42685 );
buf ( n42687 , n42614 );
buf ( n42688 , n42494 );
nor ( n42689 , n42687 , n42688 );
buf ( n42690 , n42689 );
not ( n42691 , n42647 );
nand ( n42692 , n42691 , n42654 );
buf ( n42693 , n42692 );
not ( n42694 , n42693 );
buf ( n42695 , n42694 );
buf ( n42696 , n42119 );
buf ( n42697 , n42100 );
nand ( n42698 , n42696 , n42697 );
buf ( n42699 , n42698 );
buf ( n42700 , n42601 );
buf ( n42701 , n42699 );
xnor ( n42702 , n42700 , n42701 );
buf ( n42703 , n42702 );
buf ( n42704 , n409 );
buf ( n42705 , n415 );
and ( n42706 , n42704 , n42705 );
buf ( n42707 , n42706 );
buf ( n42708 , n42707 );
buf ( n42709 , n407 );
buf ( n42710 , n417 );
and ( n42711 , n42709 , n42710 );
buf ( n42712 , n42711 );
buf ( n42713 , n42712 );
buf ( n42714 , n408 );
buf ( n42715 , n416 );
and ( n42716 , n42714 , n42715 );
buf ( n42717 , n42716 );
buf ( n42718 , n42717 );
xor ( n42719 , n42708 , n42713 );
xor ( n42720 , n42719 , n42718 );
buf ( n42721 , n42720 );
xor ( n42722 , n42708 , n42713 );
and ( n42723 , n42722 , n42718 );
and ( n42724 , n42708 , n42713 );
or ( n42725 , n42723 , n42724 );
buf ( n42726 , n42725 );
buf ( n42727 , n391 );
buf ( n42728 , n393 );
and ( n42729 , n42727 , n42728 );
buf ( n42730 , n42729 );
buf ( n42731 , n42730 );
buf ( n42732 , n392 );
buf ( n42733 , n393 );
nand ( n42734 , n42732 , n42733 );
buf ( n42735 , n42734 );
buf ( n42736 , n42735 );
buf ( n42737 , n409 );
buf ( n42738 , n416 );
nand ( n42739 , n42737 , n42738 );
buf ( n42740 , n42739 );
buf ( n42741 , n42740 );
nor ( n42742 , n42736 , n42741 );
buf ( n42743 , n42742 );
buf ( n42744 , n42743 );
buf ( n42745 , C0 );
xor ( n42746 , n42731 , n42744 );
xor ( n42747 , n42746 , n42745 );
buf ( n42748 , n42747 );
and ( n42749 , n42731 , n42744 );
or ( n42750 , C0 , n42749 );
buf ( n42751 , n42750 );
buf ( n42752 , n408 );
buf ( n42753 , n415 );
and ( n42754 , n42752 , n42753 );
buf ( n42755 , n42754 );
buf ( n42756 , n42755 );
buf ( n42757 , n407 );
buf ( n42758 , n416 );
and ( n42759 , n42757 , n42758 );
buf ( n42760 , n42759 );
buf ( n42761 , n42760 );
buf ( n42762 , n406 );
buf ( n42763 , n417 );
and ( n42764 , n42762 , n42763 );
buf ( n42765 , n42764 );
buf ( n42766 , n42765 );
xor ( n42767 , n42756 , n42761 );
xor ( n42768 , n42767 , n42766 );
buf ( n42769 , n42768 );
xor ( n42770 , n42756 , n42761 );
and ( n42771 , n42770 , n42766 );
and ( n42772 , n42756 , n42761 );
or ( n42773 , n42771 , n42772 );
buf ( n42774 , n42773 );
not ( n42775 , n392 );
nand ( n42776 , n42775 , n391 , n393 );
not ( n42777 , n391 );
nand ( n42778 , n42777 , n392 , n393 );
nand ( n42779 , n42776 , n42778 );
buf ( n42780 , n42779 );
buf ( n42781 , n409 );
buf ( n42782 , n414 );
nand ( n42783 , n42781 , n42782 );
buf ( n42784 , n42783 );
buf ( n42785 , n390 );
buf ( n42786 , n393 );
nand ( n42787 , n42785 , n42786 );
buf ( n42788 , n42787 );
xor ( n42789 , n42784 , n42788 );
buf ( n42790 , n42789 );
not ( n42791 , n392 );
nor ( n42792 , n42791 , n393 );
buf ( n42793 , n42792 );
xor ( n42794 , n42780 , n42790 );
xor ( n42795 , n42794 , n42793 );
buf ( n42796 , n42795 );
xor ( n42797 , n42780 , n42790 );
and ( n42798 , n42797 , n42793 );
and ( n42799 , n42780 , n42790 );
or ( n42800 , n42798 , n42799 );
buf ( n42801 , n42800 );
buf ( n42802 , n42726 );
buf ( n42803 , n42769 );
buf ( n42804 , n42751 );
xor ( n42805 , n42802 , n42803 );
xor ( n42806 , n42805 , n42804 );
buf ( n42807 , n42806 );
xor ( n42808 , n42802 , n42803 );
and ( n42809 , n42808 , n42804 );
and ( n42810 , n42802 , n42803 );
or ( n42811 , n42809 , n42810 );
buf ( n42812 , n42811 );
buf ( n42813 , n407 );
buf ( n42814 , n415 );
and ( n42815 , n42813 , n42814 );
buf ( n42816 , n42815 );
buf ( n42817 , n42816 );
buf ( n42818 , n409 );
buf ( n42819 , n413 );
and ( n42820 , n42818 , n42819 );
buf ( n42821 , n42820 );
buf ( n42822 , n42821 );
buf ( n42823 , n406 );
buf ( n42824 , n416 );
and ( n42825 , n42823 , n42824 );
buf ( n42826 , n42825 );
buf ( n42827 , n42826 );
xor ( n42828 , n42817 , n42822 );
xor ( n42829 , n42828 , n42827 );
buf ( n42830 , n42829 );
xor ( n42831 , n42817 , n42822 );
and ( n42832 , n42831 , n42827 );
and ( n42833 , n42817 , n42822 );
or ( n42834 , n42832 , n42833 );
buf ( n42835 , n42834 );
buf ( n42836 , n405 );
buf ( n42837 , n417 );
and ( n42838 , n42836 , n42837 );
buf ( n42839 , n42838 );
buf ( n42840 , n42839 );
buf ( n42841 , n408 );
buf ( n42842 , n414 );
and ( n42843 , n42841 , n42842 );
buf ( n42844 , n42843 );
buf ( n42845 , n42844 );
buf ( n42846 , n389 );
buf ( n42847 , n393 );
and ( n42848 , n42846 , n42847 );
buf ( n42849 , n42848 );
buf ( n42850 , n42849 );
xor ( n42851 , n42845 , n42850 );
buf ( n42852 , n42851 );
buf ( n42853 , n42852 );
buf ( n42854 , n42792 );
buf ( n42855 , n391 );
and ( n42856 , n42854 , n42855 );
buf ( n42857 , n42856 );
buf ( n42858 , n42857 );
xor ( n42859 , n42840 , n42853 );
xor ( n42860 , n42859 , n42858 );
buf ( n42861 , n42860 );
xor ( n42862 , n42840 , n42853 );
and ( n42863 , n42862 , n42858 );
and ( n42864 , n42840 , n42853 );
or ( n42865 , n42863 , n42864 );
buf ( n42866 , n42865 );
buf ( n42867 , n42788 );
buf ( n42868 , n42784 );
nor ( n42869 , n42867 , n42868 );
buf ( n42870 , n42869 );
buf ( n42871 , n42870 );
buf ( n42872 , n42779 );
buf ( n42873 , n392 );
and ( n42874 , n42872 , n42873 );
buf ( n42875 , n42874 );
buf ( n42876 , n42875 );
buf ( n42877 , n42774 );
xor ( n42878 , n42871 , n42876 );
xor ( n42879 , n42878 , n42877 );
buf ( n42880 , n42879 );
xor ( n42881 , n42871 , n42876 );
and ( n42882 , n42881 , n42877 );
and ( n42883 , n42871 , n42876 );
or ( n42884 , n42882 , n42883 );
buf ( n42885 , n42884 );
buf ( n42886 , n42830 );
buf ( n42887 , n42801 );
buf ( n42888 , n42861 );
xor ( n42889 , n42886 , n42887 );
xor ( n42890 , n42889 , n42888 );
buf ( n42891 , n42890 );
xor ( n42892 , n42886 , n42887 );
and ( n42893 , n42892 , n42888 );
and ( n42894 , n42886 , n42887 );
or ( n42895 , n42893 , n42894 );
buf ( n42896 , n42895 );
nand ( n42897 , n392 , n391 );
not ( n42898 , n42897 );
nand ( n42899 , n390 , n393 );
and ( n42900 , n42899 , n42777 );
not ( n42901 , n42899 );
and ( n42902 , n42901 , n391 );
or ( n42903 , n42900 , n42902 );
not ( n42904 , n42903 );
or ( n42905 , n42898 , n42904 );
and ( n42906 , n391 , n392 );
nand ( n42907 , n42906 , n42899 );
nand ( n42908 , n42905 , n42907 );
nand ( n42909 , n392 , n393 , n391 );
and ( n42910 , n42908 , n42909 );
not ( n42911 , n42908 );
not ( n42912 , n42909 );
and ( n42913 , n42911 , n42912 );
nor ( n42914 , n42910 , n42913 );
buf ( n42915 , n42914 );
buf ( n42916 , n42915 );
buf ( n42917 , n393 );
and ( n42918 , n42916 , n42917 );
buf ( n42919 , n42918 );
buf ( n42920 , n42919 );
buf ( n42921 , n42880 );
buf ( n42922 , n42812 );
xor ( n42923 , n42920 , n42921 );
xor ( n42924 , n42923 , n42922 );
buf ( n42925 , n42924 );
xor ( n42926 , n42920 , n42921 );
and ( n42927 , n42926 , n42922 );
and ( n42928 , n42920 , n42921 );
or ( n42929 , n42927 , n42928 );
buf ( n42930 , n42929 );
buf ( n42931 , n407 );
buf ( n42932 , n414 );
and ( n42933 , n42931 , n42932 );
buf ( n42934 , n42933 );
buf ( n42935 , n42934 );
buf ( n42936 , n408 );
buf ( n42937 , n413 );
and ( n42938 , n42936 , n42937 );
buf ( n42939 , n42938 );
buf ( n42940 , n42939 );
buf ( n42941 , n409 );
buf ( n42942 , n412 );
and ( n42943 , n42941 , n42942 );
buf ( n42944 , n42943 );
buf ( n42945 , n42944 );
xor ( n42946 , n42935 , n42940 );
xor ( n42947 , n42946 , n42945 );
buf ( n42948 , n42947 );
xor ( n42949 , n42935 , n42940 );
and ( n42950 , n42949 , n42945 );
and ( n42951 , n42935 , n42940 );
or ( n42952 , n42950 , n42951 );
buf ( n42953 , n42952 );
buf ( n42954 , n388 );
buf ( n42955 , n393 );
and ( n42956 , n42954 , n42955 );
buf ( n42957 , n42956 );
buf ( n42958 , n42957 );
buf ( n42959 , n404 );
buf ( n42960 , n417 );
and ( n42961 , n42959 , n42960 );
buf ( n42962 , n42961 );
buf ( n42963 , n42962 );
buf ( n42964 , n42792 );
buf ( n42965 , n390 );
and ( n42966 , n42964 , n42965 );
buf ( n42967 , n42966 );
buf ( n42968 , n42967 );
xor ( n42969 , n42958 , n42963 );
xor ( n42970 , n42969 , n42968 );
buf ( n42971 , n42970 );
xor ( n42972 , n42958 , n42963 );
and ( n42973 , n42972 , n42968 );
and ( n42974 , n42958 , n42963 );
or ( n42975 , n42973 , n42974 );
buf ( n42976 , n42975 );
buf ( n42977 , n405 );
buf ( n42978 , n416 );
and ( n42979 , n42977 , n42978 );
buf ( n42980 , n42979 );
buf ( n42981 , n42980 );
buf ( n42982 , n406 );
buf ( n42983 , n415 );
and ( n42984 , n42982 , n42983 );
buf ( n42985 , n42984 );
buf ( n42986 , n42985 );
xor ( n42987 , n42981 , n42986 );
buf ( n42988 , n42987 );
buf ( n42989 , n42988 );
buf ( n42990 , n42779 );
buf ( n42991 , n391 );
and ( n42992 , n42990 , n42991 );
buf ( n42993 , n42992 );
buf ( n42994 , n42993 );
and ( n42995 , n42845 , n42850 );
buf ( n42996 , n42995 );
buf ( n42997 , n42996 );
xor ( n42998 , n42989 , n42994 );
xor ( n42999 , n42998 , n42997 );
buf ( n43000 , n42999 );
xor ( n43001 , n42989 , n42994 );
and ( n43002 , n43001 , n42997 );
and ( n43003 , n42989 , n42994 );
or ( n43004 , n43002 , n43003 );
buf ( n43005 , n43004 );
buf ( n43006 , n42835 );
buf ( n43007 , n42948 );
buf ( n43008 , n42971 );
xor ( n43009 , n43006 , n43007 );
xor ( n43010 , n43009 , n43008 );
buf ( n43011 , n43010 );
xor ( n43012 , n43006 , n43007 );
and ( n43013 , n43012 , n43008 );
and ( n43014 , n43006 , n43007 );
or ( n43015 , n43013 , n43014 );
buf ( n43016 , n43015 );
buf ( n43017 , n42866 );
buf ( n43018 , n42885 );
buf ( n43019 , n43000 );
xor ( n43020 , n43017 , n43018 );
xor ( n43021 , n43020 , n43019 );
buf ( n43022 , n43021 );
xor ( n43023 , n43017 , n43018 );
and ( n43024 , n43023 , n43019 );
and ( n43025 , n43017 , n43018 );
or ( n43026 , n43024 , n43025 );
buf ( n43027 , n43026 );
buf ( n43028 , n42915 );
buf ( n43029 , n392 );
and ( n43030 , n43028 , n43029 );
buf ( n43031 , n43030 );
buf ( n43032 , n43031 );
nand ( n43033 , n392 , n390 );
nand ( n43034 , n393 , n389 );
or ( n43035 , n43033 , n43034 );
not ( n43036 , n393 );
not ( n43037 , n389 );
or ( n43038 , n43036 , n43037 );
nand ( n43039 , n392 , n390 );
nand ( n43040 , n43038 , n43039 );
nand ( n43041 , n43035 , n43040 );
buf ( n43042 , n43041 );
nand ( n43043 , n393 , n390 , n391 );
or ( n43044 , n43042 , n43043 );
nand ( n43045 , n43041 , n43043 );
buf ( n43046 , n43045 );
nand ( n43047 , n43044 , n43046 );
nand ( n43048 , n393 , n392 , n391 );
nand ( n43049 , n43048 , n42907 );
not ( n43050 , n43049 );
and ( n43051 , n43047 , n43050 );
not ( n43052 , n43047 );
and ( n43053 , n43052 , n43049 );
nor ( n43054 , n43051 , n43053 );
buf ( n43055 , n43054 );
buf ( n43056 , n393 );
and ( n43057 , n43055 , n43056 );
buf ( n43058 , n43057 );
buf ( n43059 , n43058 );
buf ( n43060 , n43011 );
xor ( n43061 , n43032 , n43059 );
xor ( n43062 , n43061 , n43060 );
buf ( n43063 , n43062 );
xor ( n43064 , n43032 , n43059 );
and ( n43065 , n43064 , n43060 );
and ( n43066 , n43032 , n43059 );
or ( n43067 , n43065 , n43066 );
buf ( n43068 , n43067 );
buf ( n43069 , n42896 );
buf ( n43070 , n43022 );
buf ( n43071 , n43063 );
xor ( n43072 , n43069 , n43070 );
xor ( n43073 , n43072 , n43071 );
buf ( n43074 , n43073 );
xor ( n43075 , n43069 , n43070 );
and ( n43076 , n43075 , n43071 );
and ( n43077 , n43069 , n43070 );
or ( n43078 , n43076 , n43077 );
buf ( n43079 , n43078 );
buf ( n43080 , n409 );
buf ( n43081 , n411 );
and ( n43082 , n43080 , n43081 );
buf ( n43083 , n43082 );
buf ( n43084 , n43083 );
buf ( n43085 , n387 );
buf ( n43086 , n393 );
and ( n43087 , n43085 , n43086 );
buf ( n43088 , n43087 );
buf ( n43089 , n43088 );
buf ( n43090 , n405 );
buf ( n43091 , n415 );
and ( n43092 , n43090 , n43091 );
buf ( n43093 , n43092 );
buf ( n43094 , n43093 );
xor ( n43095 , n43084 , n43089 );
xor ( n43096 , n43095 , n43094 );
buf ( n43097 , n43096 );
xor ( n43098 , n43084 , n43089 );
and ( n43099 , n43098 , n43094 );
and ( n43100 , n43084 , n43089 );
or ( n43101 , n43099 , n43100 );
buf ( n43102 , n43101 );
buf ( n43103 , n407 );
buf ( n43104 , n413 );
and ( n43105 , n43103 , n43104 );
buf ( n43106 , n43105 );
buf ( n43107 , n43106 );
buf ( n43108 , n408 );
buf ( n43109 , n412 );
and ( n43110 , n43108 , n43109 );
buf ( n43111 , n43110 );
buf ( n43112 , n43111 );
buf ( n43113 , n406 );
buf ( n43114 , n414 );
and ( n43115 , n43113 , n43114 );
buf ( n43116 , n43115 );
buf ( n43117 , n43116 );
xor ( n43118 , n43107 , n43112 );
xor ( n43119 , n43118 , n43117 );
buf ( n43120 , n43119 );
xor ( n43121 , n43107 , n43112 );
and ( n43122 , n43121 , n43117 );
and ( n43123 , n43107 , n43112 );
or ( n43124 , n43122 , n43123 );
buf ( n43125 , n43124 );
buf ( n43126 , n42779 );
buf ( n43127 , n390 );
and ( n43128 , n43126 , n43127 );
buf ( n43129 , n43128 );
buf ( n43130 , n43129 );
buf ( n43131 , n403 );
buf ( n43132 , n417 );
and ( n43133 , n43131 , n43132 );
buf ( n43134 , n43133 );
buf ( n43135 , n43134 );
buf ( n43136 , n404 );
buf ( n43137 , n416 );
and ( n43138 , n43136 , n43137 );
buf ( n43139 , n43138 );
buf ( n43140 , n43139 );
xor ( n43141 , n43135 , n43140 );
buf ( n43142 , n43141 );
buf ( n43143 , n43142 );
buf ( n43144 , n42792 );
buf ( n43145 , n389 );
and ( n43146 , n43144 , n43145 );
buf ( n43147 , n43146 );
buf ( n43148 , n43147 );
xor ( n43149 , n43130 , n43143 );
xor ( n43150 , n43149 , n43148 );
buf ( n43151 , n43150 );
xor ( n43152 , n43130 , n43143 );
and ( n43153 , n43152 , n43148 );
and ( n43154 , n43130 , n43143 );
or ( n43155 , n43153 , n43154 );
buf ( n43156 , n43155 );
and ( n43157 , n42981 , n42986 );
buf ( n43158 , n43157 );
buf ( n43159 , n43158 );
buf ( n43160 , n42953 );
buf ( n43161 , n43097 );
xor ( n43162 , n43159 , n43160 );
xor ( n43163 , n43162 , n43161 );
buf ( n43164 , n43163 );
xor ( n43165 , n43159 , n43160 );
and ( n43166 , n43165 , n43161 );
and ( n43167 , n43159 , n43160 );
or ( n43168 , n43166 , n43167 );
buf ( n43169 , n43168 );
buf ( n43170 , n43120 );
buf ( n43171 , n42976 );
buf ( n43172 , n43005 );
xor ( n43173 , n43170 , n43171 );
xor ( n43174 , n43173 , n43172 );
buf ( n43175 , n43174 );
xor ( n43176 , n43170 , n43171 );
and ( n43177 , n43176 , n43172 );
and ( n43178 , n43170 , n43171 );
or ( n43179 , n43177 , n43178 );
buf ( n43180 , n43179 );
buf ( n43181 , n42914 );
buf ( n43182 , n391 );
and ( n43183 , n43181 , n43182 );
buf ( n43184 , n43183 );
buf ( n43185 , n43184 );
buf ( n43186 , n43151 );
not ( n43187 , n43054 );
buf ( n43188 , n392 );
not ( n43189 , n43188 );
buf ( n43190 , n43189 );
nor ( n43191 , n43187 , n43190 );
buf ( n43192 , n43191 );
xor ( n43193 , n43185 , n43186 );
xor ( n43194 , n43193 , n43192 );
buf ( n43195 , n43194 );
xor ( n43196 , n43185 , n43186 );
and ( n43197 , n43196 , n43192 );
and ( n43198 , n43185 , n43186 );
or ( n43199 , n43197 , n43198 );
buf ( n43200 , n43199 );
buf ( n43201 , n43164 );
nand ( n43202 , n389 , n392 , n390 , n393 );
nand ( n43203 , n388 , n393 );
not ( n43204 , n43203 );
and ( n43205 , n389 , n392 );
xor ( n43206 , n43204 , n43205 );
not ( n43207 , n390 );
nor ( n43208 , n43207 , n391 );
xor ( n43209 , n43206 , n43208 );
xor ( n43210 , n43202 , n43209 );
not ( n43211 , n42907 );
not ( n43212 , n43211 );
not ( n43213 , n43045 );
or ( n43214 , n43212 , n43213 );
not ( n43215 , n43041 );
not ( n43216 , n43043 );
and ( n43217 , n43215 , n43216 );
not ( n43218 , n43048 );
and ( n43219 , n43045 , n43218 );
nor ( n43220 , n43217 , n43219 );
nand ( n43221 , n43214 , n43220 );
xnor ( n43222 , n43210 , n43221 );
buf ( n43223 , n43222 );
buf ( n43224 , n393 );
and ( n43225 , n43223 , n43224 );
buf ( n43226 , n43225 );
buf ( n43227 , n43226 );
buf ( n43228 , n43016 );
xor ( n43229 , n43201 , n43227 );
xor ( n43230 , n43229 , n43228 );
buf ( n43231 , n43230 );
xor ( n43232 , n43201 , n43227 );
and ( n43233 , n43232 , n43228 );
and ( n43234 , n43201 , n43227 );
or ( n43235 , n43233 , n43234 );
buf ( n43236 , n43235 );
buf ( n43237 , n43027 );
buf ( n43238 , n43175 );
buf ( n43239 , n43195 );
xor ( n43240 , n43237 , n43238 );
xor ( n43241 , n43240 , n43239 );
buf ( n43242 , n43241 );
xor ( n43243 , n43237 , n43238 );
and ( n43244 , n43243 , n43239 );
and ( n43245 , n43237 , n43238 );
or ( n43246 , n43244 , n43245 );
buf ( n43247 , n43246 );
buf ( n43248 , n43068 );
buf ( n43249 , n43231 );
buf ( n43250 , n43242 );
xor ( n43251 , n43248 , n43249 );
xor ( n43252 , n43251 , n43250 );
buf ( n43253 , n43252 );
xor ( n43254 , n43248 , n43249 );
and ( n43255 , n43254 , n43250 );
and ( n43256 , n43248 , n43249 );
or ( n43257 , n43255 , n43256 );
buf ( n43258 , n43257 );
buf ( n43259 , n406 );
buf ( n43260 , n413 );
and ( n43261 , n43259 , n43260 );
buf ( n43262 , n43261 );
buf ( n43263 , n43262 );
buf ( n43264 , n403 );
buf ( n43265 , n416 );
and ( n43266 , n43264 , n43265 );
buf ( n43267 , n43266 );
buf ( n43268 , n43267 );
buf ( n43269 , n404 );
buf ( n43270 , n415 );
and ( n43271 , n43269 , n43270 );
buf ( n43272 , n43271 );
buf ( n43273 , n43272 );
xor ( n43274 , n43263 , n43268 );
xor ( n43275 , n43274 , n43273 );
buf ( n43276 , n43275 );
xor ( n43277 , n43263 , n43268 );
and ( n43278 , n43277 , n43273 );
and ( n43279 , n43263 , n43268 );
or ( n43280 , n43278 , n43279 );
buf ( n43281 , n43280 );
buf ( n43282 , n409 );
buf ( n43283 , n410 );
and ( n43284 , n43282 , n43283 );
buf ( n43285 , n43284 );
buf ( n43286 , n43285 );
and ( n43287 , n405 , n414 );
buf ( n43288 , n43287 );
buf ( n43289 , n407 );
buf ( n43290 , n412 );
and ( n43291 , n43289 , n43290 );
buf ( n43292 , n43291 );
buf ( n43293 , n43292 );
xor ( n43294 , n43286 , n43288 );
xor ( n43295 , n43294 , n43293 );
buf ( n43296 , n43295 );
xor ( n43297 , n43286 , n43288 );
and ( n43298 , n43297 , n43293 );
and ( n43299 , n43286 , n43288 );
or ( n43300 , n43298 , n43299 );
buf ( n43301 , n43300 );
buf ( n43302 , n43247 );
buf ( n43303 , n43200 );
not ( n43304 , n43202 );
not ( n43305 , n43304 );
not ( n43306 , n43209 );
not ( n43307 , n43306 );
not ( n43308 , n43307 );
or ( n43309 , n43305 , n43308 );
not ( n43310 , n43202 );
not ( n43311 , n43306 );
or ( n43312 , n43310 , n43311 );
nand ( n43313 , n43312 , n43221 );
nand ( n43314 , n43309 , n43313 );
not ( n43315 , n43314 );
nand ( n43316 , n389 , n391 );
not ( n43317 , n43316 );
and ( n43318 , n388 , n392 );
xor ( n43319 , n43317 , n43318 );
xor ( n43320 , n43088 , n43319 );
and ( n43321 , n390 , n391 );
xor ( n43322 , n43320 , n43321 );
not ( n43323 , n43322 );
xor ( n43324 , n43204 , n43205 );
and ( n43325 , n43324 , n43208 );
and ( n43326 , n43204 , n43205 );
or ( n43327 , n43325 , n43326 );
and ( n43328 , n43323 , n43327 );
nand ( n43329 , n43315 , n43328 );
not ( n43330 , n43304 );
not ( n43331 , n43209 );
or ( n43332 , n43330 , n43331 );
or ( n43333 , n43209 , n43304 );
nand ( n43334 , n43333 , n43221 );
nand ( n43335 , n43332 , n43334 );
not ( n43336 , n43335 );
not ( n43337 , n43327 );
and ( n43338 , n43322 , n43337 );
nand ( n43339 , n43336 , n43338 );
nand ( n43340 , n43322 , n43327 );
not ( n43341 , n43340 );
nand ( n43342 , n43323 , n43337 );
not ( n43343 , n43342 );
or ( n43344 , n43341 , n43343 );
nand ( n43345 , n43344 , n43314 );
nand ( n43346 , n43329 , n43339 , n43345 );
buf ( n43347 , n43346 );
buf ( n43348 , n393 );
and ( n43349 , n43347 , n43348 );
buf ( n43350 , n43349 );
buf ( n43351 , n43350 );
xor ( n43352 , n43303 , n43351 );
buf ( n43353 , n43156 );
buf ( n43354 , n42915 );
buf ( n43355 , n390 );
and ( n43356 , n43354 , n43355 );
buf ( n43357 , n43356 );
buf ( n43358 , n43357 );
xor ( n43359 , n43353 , n43358 );
buf ( n43360 , n42792 );
buf ( n43361 , n388 );
and ( n43362 , n43360 , n43361 );
buf ( n43363 , n43362 );
buf ( n43364 , n43363 );
not ( n43365 , n42779 );
not ( n43366 , n389 );
nor ( n43367 , n43365 , n43366 );
buf ( n43368 , n43367 );
xor ( n43369 , n43364 , n43368 );
buf ( n43370 , n43102 );
xor ( n43371 , n43369 , n43370 );
buf ( n43372 , n43371 );
buf ( n43373 , n43372 );
xor ( n43374 , n43359 , n43373 );
buf ( n43375 , n43374 );
buf ( n43376 , n43375 );
xor ( n43377 , n43352 , n43376 );
buf ( n43378 , n43377 );
buf ( n43379 , n43378 );
buf ( n43380 , n43236 );
buf ( n43381 , n408 );
buf ( n43382 , n411 );
and ( n43383 , n43381 , n43382 );
buf ( n43384 , n43383 );
buf ( n43385 , n43384 );
buf ( n43386 , n402 );
buf ( n43387 , n417 );
nand ( n43388 , n43386 , n43387 );
buf ( n43389 , n43388 );
buf ( n43390 , n386 );
buf ( n43391 , n393 );
nand ( n43392 , n43390 , n43391 );
buf ( n43393 , n43392 );
xor ( n43394 , n43389 , n43393 );
buf ( n43395 , n43394 );
xor ( n43396 , n43385 , n43395 );
and ( n43397 , n43135 , n43140 );
buf ( n43398 , n43397 );
buf ( n43399 , n43398 );
xor ( n43400 , n43396 , n43399 );
buf ( n43401 , n43400 );
buf ( n43402 , n43401 );
buf ( n43403 , n43054 );
buf ( n43404 , n391 );
and ( n43405 , n43403 , n43404 );
buf ( n43406 , n43405 );
buf ( n43407 , n43406 );
xor ( n43408 , n43402 , n43407 );
buf ( n43409 , n43169 );
xor ( n43410 , n43408 , n43409 );
buf ( n43411 , n43410 );
buf ( n43412 , n43411 );
xor ( n43413 , n43380 , n43412 );
buf ( n43414 , n43180 );
buf ( n43415 , n43222 );
buf ( n43416 , n392 );
and ( n43417 , n43415 , n43416 );
buf ( n43418 , n43417 );
buf ( n43419 , n43418 );
xor ( n43420 , n43414 , n43419 );
buf ( n43421 , n43125 );
buf ( n43422 , n43296 );
xor ( n43423 , n43421 , n43422 );
buf ( n43424 , n43276 );
xor ( n43425 , n43423 , n43424 );
buf ( n43426 , n43425 );
buf ( n43427 , n43426 );
xor ( n43428 , n43420 , n43427 );
buf ( n43429 , n43428 );
buf ( n43430 , n43429 );
xor ( n43431 , n43413 , n43430 );
buf ( n43432 , n43431 );
buf ( n43433 , n43432 );
xor ( n43434 , n43302 , n43379 );
xor ( n43435 , n43434 , n43433 );
buf ( n43436 , n43435 );
xor ( n43437 , n43302 , n43379 );
and ( n43438 , n43437 , n43433 );
and ( n43439 , n43302 , n43379 );
or ( n43440 , n43438 , n43439 );
buf ( n43441 , n43440 );
xor ( n43442 , n43385 , n43395 );
and ( n43443 , n43442 , n43399 );
and ( n43444 , n43385 , n43395 );
or ( n43445 , n43443 , n43444 );
buf ( n43446 , n43445 );
xor ( n43447 , n43364 , n43368 );
and ( n43448 , n43447 , n43370 );
or ( n43449 , n43448 , C0 );
buf ( n43450 , n43449 );
xor ( n43451 , n43421 , n43422 );
and ( n43452 , n43451 , n43424 );
and ( n43453 , n43421 , n43422 );
or ( n43454 , n43452 , n43453 );
buf ( n43455 , n43454 );
xor ( n43456 , n43353 , n43358 );
and ( n43457 , n43456 , n43373 );
and ( n43458 , n43353 , n43358 );
or ( n43459 , n43457 , n43458 );
buf ( n43460 , n43459 );
xor ( n43461 , n43402 , n43407 );
and ( n43462 , n43461 , n43409 );
and ( n43463 , n43402 , n43407 );
or ( n43464 , n43462 , n43463 );
buf ( n43465 , n43464 );
xor ( n43466 , n43414 , n43419 );
and ( n43467 , n43466 , n43427 );
and ( n43468 , n43414 , n43419 );
or ( n43469 , n43467 , n43468 );
buf ( n43470 , n43469 );
xor ( n43471 , n43303 , n43351 );
and ( n43472 , n43471 , n43376 );
and ( n43473 , n43303 , n43351 );
or ( n43474 , n43472 , n43473 );
buf ( n43475 , n43474 );
xor ( n43476 , n43380 , n43412 );
and ( n43477 , n43476 , n43430 );
and ( n43478 , n43380 , n43412 );
or ( n43479 , n43477 , n43478 );
buf ( n43480 , n43479 );
buf ( n43481 , n408 );
buf ( n43482 , n410 );
and ( n43483 , n43481 , n43482 );
buf ( n43484 , n43483 );
buf ( n43485 , n43484 );
buf ( n43486 , n403 );
buf ( n43487 , n415 );
and ( n43488 , n43486 , n43487 );
buf ( n43489 , n43488 );
buf ( n43490 , n43489 );
buf ( n43491 , n404 );
buf ( n43492 , n414 );
and ( n43493 , n43491 , n43492 );
buf ( n43494 , n43493 );
buf ( n43495 , n43494 );
xor ( n43496 , n43485 , n43490 );
xor ( n43497 , n43496 , n43495 );
buf ( n43498 , n43497 );
xor ( n43499 , n43485 , n43490 );
and ( n43500 , n43499 , n43495 );
and ( n43501 , n43485 , n43490 );
or ( n43502 , n43500 , n43501 );
buf ( n43503 , n43502 );
buf ( n43504 , n402 );
buf ( n43505 , n416 );
and ( n43506 , n43504 , n43505 );
buf ( n43507 , n43506 );
buf ( n43508 , n43507 );
buf ( n43509 , n407 );
buf ( n43510 , n411 );
and ( n43511 , n43509 , n43510 );
buf ( n43512 , n43511 );
buf ( n43513 , n43512 );
buf ( n43514 , n405 );
buf ( n43515 , n413 );
and ( n43516 , n43514 , n43515 );
buf ( n43517 , n43516 );
buf ( n43518 , n43517 );
xor ( n43519 , n43508 , n43513 );
xor ( n43520 , n43519 , n43518 );
buf ( n43521 , n43520 );
xor ( n43522 , n43508 , n43513 );
and ( n43523 , n43522 , n43518 );
and ( n43524 , n43508 , n43513 );
or ( n43525 , n43523 , n43524 );
buf ( n43526 , n43525 );
buf ( n43527 , n43521 );
buf ( n43528 , n43498 );
xor ( n43529 , n43527 , n43528 );
buf ( n43530 , n43446 );
xor ( n43531 , n43529 , n43530 );
buf ( n43532 , n43531 );
buf ( n43533 , n43532 );
buf ( n43534 , n43222 );
buf ( n43535 , n391 );
and ( n43536 , n43534 , n43535 );
buf ( n43537 , n43536 );
buf ( n43538 , n43537 );
xor ( n43539 , n43533 , n43538 );
buf ( n43540 , n43460 );
xor ( n43541 , n43539 , n43540 );
buf ( n43542 , n43541 );
buf ( n43543 , n43542 );
buf ( n43544 , n43475 );
buf ( n43545 , n43346 );
buf ( n43546 , n392 );
and ( n43547 , n43545 , n43546 );
buf ( n43548 , n43547 );
buf ( n43549 , n43548 );
buf ( n43550 , n43465 );
xor ( n43551 , n43549 , n43550 );
buf ( n43552 , n406 );
buf ( n43553 , n412 );
and ( n43554 , n43552 , n43553 );
buf ( n43555 , n43554 );
buf ( n43556 , n43555 );
buf ( n43557 , n43393 );
buf ( n43558 , n43389 );
nor ( n43559 , n43557 , n43558 );
buf ( n43560 , n43559 );
buf ( n43561 , n43560 );
xor ( n43562 , n43556 , n43561 );
buf ( n43563 , n42779 );
not ( n43564 , n43563 );
buf ( n43565 , n388 );
not ( n43566 , n43565 );
buf ( n43567 , n43566 );
buf ( n43568 , n43567 );
nor ( n43569 , n43564 , n43568 );
buf ( n43570 , n43569 );
buf ( n43571 , n43570 );
xor ( n43572 , n43562 , n43571 );
buf ( n43573 , n43572 );
buf ( n43574 , n43573 );
buf ( n43575 , n43450 );
xor ( n43576 , n43574 , n43575 );
not ( n43577 , n42915 );
buf ( n43578 , n43577 );
buf ( n43579 , n43366 );
nor ( n43580 , n43578 , n43579 );
buf ( n43581 , n43580 );
buf ( n43582 , n43581 );
xor ( n43583 , n43576 , n43582 );
buf ( n43584 , n43583 );
buf ( n43585 , n43584 );
xor ( n43586 , n43551 , n43585 );
buf ( n43587 , n43586 );
buf ( n43588 , n43587 );
xor ( n43589 , n43543 , n43544 );
xor ( n43590 , n43589 , n43588 );
buf ( n43591 , n43590 );
xor ( n43592 , n43543 , n43544 );
and ( n43593 , n43592 , n43588 );
and ( n43594 , n43543 , n43544 );
or ( n43595 , n43593 , n43594 );
buf ( n43596 , n43595 );
xor ( n43597 , n43088 , n43319 );
and ( n43598 , n43597 , n43321 );
and ( n43599 , n43088 , n43319 );
or ( n43600 , n43598 , n43599 );
and ( n43601 , n389 , n390 );
xor ( n43602 , n389 , n43601 );
and ( n43603 , n43317 , n43318 );
xor ( n43604 , n43602 , n43603 );
nand ( n43605 , n387 , n392 );
not ( n43606 , n43605 );
and ( n43607 , n386 , n393 );
xor ( n43608 , n43606 , n43607 );
and ( n43609 , n388 , n391 );
xor ( n43610 , n43608 , n43609 );
xor ( n43611 , n43604 , n43610 );
not ( n43612 , n43611 );
xor ( n43613 , n43600 , n43612 );
not ( n43614 , n43342 );
not ( n43615 , n43335 );
or ( n43616 , n43614 , n43615 );
buf ( n43617 , n43340 );
nand ( n43618 , n43616 , n43617 );
xnor ( n43619 , n43613 , n43618 );
buf ( n43620 , n43619 );
buf ( n43621 , n43620 );
buf ( n43622 , n393 );
and ( n43623 , n43621 , n43622 );
buf ( n43624 , n43623 );
buf ( n43625 , n43624 );
buf ( n43626 , n43455 );
buf ( n43627 , n43054 );
buf ( n43628 , n390 );
and ( n43629 , n43627 , n43628 );
buf ( n43630 , n43629 );
buf ( n43631 , n43630 );
xor ( n43632 , n43626 , n43631 );
buf ( n43633 , n42792 );
buf ( n43634 , n387 );
and ( n43635 , n43633 , n43634 );
buf ( n43636 , n43635 );
buf ( n43637 , n43636 );
buf ( n43638 , n43281 );
xor ( n43639 , n43637 , n43638 );
buf ( n43640 , n43301 );
xor ( n43641 , n43639 , n43640 );
buf ( n43642 , n43641 );
buf ( n43643 , n43642 );
xor ( n43644 , n43632 , n43643 );
buf ( n43645 , n43644 );
buf ( n43646 , n43645 );
xor ( n43647 , n43625 , n43646 );
buf ( n43648 , n43470 );
xor ( n43649 , n43647 , n43648 );
buf ( n43650 , n43649 );
buf ( n43651 , n43650 );
buf ( n43652 , n43480 );
buf ( n43653 , n43591 );
xor ( n43654 , n43651 , n43652 );
xor ( n43655 , n43654 , n43653 );
buf ( n43656 , n43655 );
xor ( n43657 , n43651 , n43652 );
and ( n43658 , n43657 , n43653 );
and ( n43659 , n43651 , n43652 );
or ( n43660 , n43658 , n43659 );
buf ( n43661 , n43660 );
xor ( n43662 , n43556 , n43561 );
and ( n43663 , n43662 , n43571 );
and ( n43664 , n43556 , n43561 );
or ( n43665 , n43663 , n43664 );
buf ( n43666 , n43665 );
xor ( n43667 , n43637 , n43638 );
and ( n43668 , n43667 , n43640 );
and ( n43669 , n43637 , n43638 );
or ( n43670 , n43668 , n43669 );
buf ( n43671 , n43670 );
xor ( n43672 , n43527 , n43528 );
and ( n43673 , n43672 , n43530 );
and ( n43674 , n43527 , n43528 );
or ( n43675 , n43673 , n43674 );
buf ( n43676 , n43675 );
xor ( n43677 , n43574 , n43575 );
and ( n43678 , n43677 , n43582 );
and ( n43679 , n43574 , n43575 );
or ( n43680 , n43678 , n43679 );
buf ( n43681 , n43680 );
xor ( n43682 , n43626 , n43631 );
and ( n43683 , n43682 , n43643 );
and ( n43684 , n43626 , n43631 );
or ( n43685 , n43683 , n43684 );
buf ( n43686 , n43685 );
xor ( n43687 , n43533 , n43538 );
and ( n43688 , n43687 , n43540 );
and ( n43689 , n43533 , n43538 );
or ( n43690 , n43688 , n43689 );
buf ( n43691 , n43690 );
xor ( n43692 , n43549 , n43550 );
and ( n43693 , n43692 , n43585 );
and ( n43694 , n43549 , n43550 );
or ( n43695 , n43693 , n43694 );
buf ( n43696 , n43695 );
xor ( n43697 , n43625 , n43646 );
and ( n43698 , n43697 , n43648 );
and ( n43699 , n43625 , n43646 );
or ( n43700 , n43698 , n43699 );
buf ( n43701 , n43700 );
buf ( n43702 , n402 );
buf ( n43703 , n415 );
and ( n43704 , n43702 , n43703 );
buf ( n43705 , n43704 );
buf ( n43706 , n43705 );
buf ( n43707 , n403 );
buf ( n43708 , n414 );
and ( n43709 , n43707 , n43708 );
buf ( n43710 , n43709 );
buf ( n43711 , n43710 );
buf ( n43712 , n406 );
buf ( n43713 , n411 );
and ( n43714 , n43712 , n43713 );
buf ( n43715 , n43714 );
buf ( n43716 , n43715 );
xor ( n43717 , n43706 , n43711 );
xor ( n43718 , n43717 , n43716 );
buf ( n43719 , n43718 );
xor ( n43720 , n43706 , n43711 );
and ( n43721 , n43720 , n43716 );
and ( n43722 , n43706 , n43711 );
or ( n43723 , n43721 , n43722 );
buf ( n43724 , n43723 );
buf ( n43725 , n404 );
buf ( n43726 , n413 );
and ( n43727 , n43725 , n43726 );
buf ( n43728 , n43727 );
buf ( n43729 , n43728 );
buf ( n43730 , n405 );
buf ( n43731 , n412 );
and ( n43732 , n43730 , n43731 );
buf ( n43733 , n43732 );
buf ( n43734 , n43733 );
buf ( n43735 , n407 );
buf ( n43736 , n410 );
and ( n43737 , n43735 , n43736 );
buf ( n43738 , n43737 );
buf ( n43739 , n43738 );
xor ( n43740 , n43729 , n43734 );
xor ( n43741 , n43740 , n43739 );
buf ( n43742 , n43741 );
xor ( n43743 , n43729 , n43734 );
and ( n43744 , n43743 , n43739 );
and ( n43745 , n43729 , n43734 );
or ( n43746 , n43744 , n43745 );
buf ( n43747 , n43746 );
buf ( n43748 , n43701 );
buf ( n43749 , n43686 );
buf ( n43750 , n43346 );
buf ( n43751 , n391 );
and ( n43752 , n43750 , n43751 );
buf ( n43753 , n43752 );
buf ( n43754 , n43753 );
xor ( n43755 , n43749 , n43754 );
buf ( n43756 , n43666 );
buf ( n43757 , n42792 );
buf ( n43758 , n386 );
and ( n43759 , n43757 , n43758 );
buf ( n43760 , n43759 );
buf ( n43761 , n43760 );
buf ( n43762 , n42779 );
buf ( n43763 , n387 );
and ( n43764 , n43762 , n43763 );
buf ( n43765 , n43764 );
buf ( n43766 , n43765 );
xor ( n43767 , n43761 , n43766 );
buf ( n43768 , n43526 );
xor ( n43769 , n43767 , n43768 );
buf ( n43770 , n43769 );
buf ( n43771 , n43770 );
xor ( n43772 , n43756 , n43771 );
buf ( n43773 , n43577 );
buf ( n43774 , n43567 );
nor ( n43775 , n43773 , n43774 );
buf ( n43776 , n43775 );
buf ( n43777 , n43776 );
xor ( n43778 , n43772 , n43777 );
buf ( n43779 , n43778 );
buf ( n43780 , n43779 );
xor ( n43781 , n43755 , n43780 );
buf ( n43782 , n43781 );
buf ( n43783 , n43782 );
buf ( n43784 , n43620 );
buf ( n43785 , n392 );
and ( n43786 , n43784 , n43785 );
buf ( n43787 , n43786 );
buf ( n43788 , n43787 );
buf ( n43789 , n43671 );
buf ( n43790 , n43054 );
buf ( n43791 , n389 );
and ( n43792 , n43790 , n43791 );
buf ( n43793 , n43792 );
buf ( n43794 , n43793 );
xor ( n43795 , n43789 , n43794 );
buf ( n43796 , n43676 );
xor ( n43797 , n43795 , n43796 );
buf ( n43798 , n43797 );
buf ( n43799 , n43798 );
xor ( n43800 , n43788 , n43799 );
not ( n43801 , n43611 );
not ( n43802 , n43600 );
nand ( n43803 , n43801 , n43802 );
not ( n43804 , n43803 );
not ( n43805 , n43618 );
or ( n43806 , n43804 , n43805 );
nand ( n43807 , n43611 , n43600 );
nand ( n43808 , n43806 , n43807 );
buf ( n43809 , n43808 );
and ( n43810 , n389 , n43601 );
xor ( n43811 , n43606 , n43607 );
and ( n43812 , n43811 , n43609 );
and ( n43813 , n43606 , n43607 );
or ( n43814 , n43812 , n43813 );
xor ( n43815 , n43810 , n43814 );
and ( n43816 , n388 , n390 );
and ( n43817 , n387 , n391 );
xor ( n43818 , n43816 , n43817 );
and ( n43819 , n386 , n392 );
xor ( n43820 , n43818 , n43819 );
xor ( n43821 , n43815 , n43820 );
not ( n43822 , n43821 );
xor ( n43823 , n43602 , n43603 );
and ( n43824 , n43823 , n43610 );
and ( n43825 , n43602 , n43603 );
or ( n43826 , n43824 , n43825 );
not ( n43827 , n43826 );
nand ( n43828 , n43822 , n43827 );
nand ( n43829 , n43821 , n43826 );
nand ( n43830 , n43828 , n43829 );
not ( n43831 , n43830 );
and ( n43832 , n43809 , n43831 );
not ( n43833 , n43809 );
and ( n43834 , n43833 , n43830 );
nor ( n43835 , n43832 , n43834 );
buf ( n43836 , n43835 );
buf ( n43837 , n43836 );
buf ( n43838 , n43837 );
buf ( n43839 , n43838 );
buf ( n43840 , n393 );
and ( n43841 , n43839 , n43840 );
buf ( n43842 , n43841 );
buf ( n43843 , n43842 );
xor ( n43844 , n43800 , n43843 );
buf ( n43845 , n43844 );
buf ( n43846 , n43845 );
xor ( n43847 , n43748 , n43783 );
xor ( n43848 , n43847 , n43846 );
buf ( n43849 , n43848 );
xor ( n43850 , n43748 , n43783 );
and ( n43851 , n43850 , n43846 );
and ( n43852 , n43748 , n43783 );
or ( n43853 , n43851 , n43852 );
buf ( n43854 , n43853 );
buf ( n43855 , n43691 );
buf ( n43856 , n43503 );
buf ( n43857 , n43742 );
xor ( n43858 , n43856 , n43857 );
buf ( n43859 , n43719 );
xor ( n43860 , n43858 , n43859 );
buf ( n43861 , n43860 );
buf ( n43862 , n43861 );
buf ( n43863 , n43222 );
buf ( n43864 , n390 );
and ( n43865 , n43863 , n43864 );
buf ( n43866 , n43865 );
buf ( n43867 , n43866 );
xor ( n43868 , n43862 , n43867 );
buf ( n43869 , n43681 );
xor ( n43870 , n43868 , n43869 );
buf ( n43871 , n43870 );
buf ( n43872 , n43871 );
xor ( n43873 , n43855 , n43872 );
buf ( n43874 , n43696 );
xor ( n43875 , n43873 , n43874 );
buf ( n43876 , n43875 );
buf ( n43877 , n43876 );
buf ( n43878 , n43596 );
buf ( n43879 , n43849 );
xor ( n43880 , n43877 , n43878 );
xor ( n43881 , n43880 , n43879 );
buf ( n43882 , n43881 );
xor ( n43883 , n43877 , n43878 );
and ( n43884 , n43883 , n43879 );
and ( n43885 , n43877 , n43878 );
or ( n43886 , n43884 , n43885 );
buf ( n43887 , n43886 );
xor ( n43888 , n43761 , n43766 );
and ( n43889 , n43888 , n43768 );
or ( n43890 , n43889 , C0 );
buf ( n43891 , n43890 );
xor ( n43892 , n43856 , n43857 );
and ( n43893 , n43892 , n43859 );
and ( n43894 , n43856 , n43857 );
or ( n43895 , n43893 , n43894 );
buf ( n43896 , n43895 );
xor ( n43897 , n43756 , n43771 );
and ( n43898 , n43897 , n43777 );
and ( n43899 , n43756 , n43771 );
or ( n43900 , n43898 , n43899 );
buf ( n43901 , n43900 );
xor ( n43902 , n43789 , n43794 );
and ( n43903 , n43902 , n43796 );
and ( n43904 , n43789 , n43794 );
or ( n43905 , n43903 , n43904 );
buf ( n43906 , n43905 );
xor ( n43907 , n43862 , n43867 );
and ( n43908 , n43907 , n43869 );
and ( n43909 , n43862 , n43867 );
or ( n43910 , n43908 , n43909 );
buf ( n43911 , n43910 );
xor ( n43912 , n43749 , n43754 );
and ( n43913 , n43912 , n43780 );
and ( n43914 , n43749 , n43754 );
or ( n43915 , n43913 , n43914 );
buf ( n43916 , n43915 );
xor ( n43917 , n43788 , n43799 );
and ( n43918 , n43917 , n43843 );
and ( n43919 , n43788 , n43799 );
or ( n43920 , n43918 , n43919 );
buf ( n43921 , n43920 );
xor ( n43922 , n43855 , n43872 );
and ( n43923 , n43922 , n43874 );
and ( n43924 , n43855 , n43872 );
or ( n43925 , n43923 , n43924 );
buf ( n43926 , n43925 );
buf ( n43927 , n406 );
buf ( n43928 , n410 );
and ( n43929 , n43927 , n43928 );
buf ( n43930 , n43929 );
buf ( n43931 , n43930 );
buf ( n43932 , n404 );
buf ( n43933 , n412 );
and ( n43934 , n43932 , n43933 );
buf ( n43935 , n43934 );
buf ( n43936 , n43935 );
buf ( n43937 , n405 );
buf ( n43938 , n411 );
and ( n43939 , n43937 , n43938 );
buf ( n43940 , n43939 );
buf ( n43941 , n43940 );
xor ( n43942 , n43931 , n43936 );
xor ( n43943 , n43942 , n43941 );
buf ( n43944 , n43943 );
xor ( n43945 , n43931 , n43936 );
and ( n43946 , n43945 , n43941 );
and ( n43947 , n43931 , n43936 );
or ( n43948 , n43946 , n43947 );
buf ( n43949 , n43948 );
buf ( n43950 , n42779 );
buf ( n43951 , n386 );
and ( n43952 , n43950 , n43951 );
buf ( n43953 , n43952 );
buf ( n43954 , n43953 );
buf ( n43955 , n402 );
buf ( n43956 , n414 );
and ( n43957 , n43955 , n43956 );
buf ( n43958 , n43957 );
buf ( n43959 , n43958 );
buf ( n43960 , n403 );
buf ( n43961 , n413 );
and ( n43962 , n43960 , n43961 );
buf ( n43963 , n43962 );
buf ( n43964 , n43963 );
xor ( n43965 , n43959 , n43964 );
buf ( n43966 , n43965 );
buf ( n43967 , n43966 );
buf ( n43968 , n43747 );
xor ( n43969 , n43954 , n43967 );
xor ( n43970 , n43969 , n43968 );
buf ( n43971 , n43970 );
xor ( n43972 , n43954 , n43967 );
and ( n43973 , n43972 , n43968 );
and ( n43974 , n43954 , n43967 );
or ( n43975 , n43973 , n43974 );
buf ( n43976 , n43975 );
buf ( n43977 , n43916 );
buf ( n43978 , n43901 );
buf ( n43979 , n42914 );
not ( n43980 , n43979 );
buf ( n43981 , n387 );
not ( n43982 , n43981 );
buf ( n43983 , n43982 );
buf ( n43984 , n43983 );
nor ( n43985 , n43980 , n43984 );
buf ( n43986 , n43985 );
buf ( n43987 , n43986 );
buf ( n43988 , n43971 );
xor ( n43989 , n43987 , n43988 );
buf ( n43990 , n43896 );
xor ( n43991 , n43989 , n43990 );
buf ( n43992 , n43991 );
buf ( n43993 , n43992 );
xor ( n43994 , n43978 , n43993 );
not ( n43995 , n390 );
buf ( n43996 , n43346 );
not ( n43997 , n43996 );
buf ( n43998 , n43997 );
nor ( n43999 , n43995 , n43998 );
buf ( n44000 , n43999 );
xor ( n44001 , n43994 , n44000 );
buf ( n44002 , n44001 );
buf ( n44003 , n44002 );
xor ( n44004 , n43977 , n44003 );
buf ( n44005 , n43921 );
xor ( n44006 , n44004 , n44005 );
buf ( n44007 , n44006 );
buf ( n44008 , n44007 );
buf ( n44009 , n43854 );
buf ( n44010 , n43619 );
buf ( n44011 , n391 );
and ( n44012 , n44010 , n44011 );
buf ( n44013 , n44012 );
buf ( n44014 , n44013 );
buf ( n44015 , n43906 );
xor ( n44016 , n44014 , n44015 );
buf ( n44017 , n43911 );
xor ( n44018 , n44016 , n44017 );
buf ( n44019 , n44018 );
buf ( n44020 , n44019 );
buf ( n44021 , n43838 );
buf ( n44022 , n392 );
and ( n44023 , n44021 , n44022 );
buf ( n44024 , n44023 );
buf ( n44025 , n44024 );
buf ( n44026 , n43054 );
buf ( n44027 , n388 );
and ( n44028 , n44026 , n44027 );
buf ( n44029 , n44028 );
buf ( n44030 , n44029 );
buf ( n44031 , n43222 );
buf ( n44032 , n389 );
and ( n44033 , n44031 , n44032 );
buf ( n44034 , n44033 );
buf ( n44035 , n44034 );
xor ( n44036 , n44030 , n44035 );
buf ( n44037 , n43724 );
buf ( n44038 , n43944 );
xor ( n44039 , n44037 , n44038 );
buf ( n44040 , n43891 );
xor ( n44041 , n44039 , n44040 );
buf ( n44042 , n44041 );
buf ( n44043 , n44042 );
xor ( n44044 , n44036 , n44043 );
buf ( n44045 , n44044 );
buf ( n44046 , n44045 );
xor ( n44047 , n44025 , n44046 );
not ( n44048 , n43828 );
not ( n44049 , n43809 );
or ( n44050 , n44048 , n44049 );
nand ( n44051 , n44050 , n43829 );
xor ( n44052 , n43810 , n43814 );
and ( n44053 , n44052 , n43820 );
and ( n44054 , n43810 , n43814 );
or ( n44055 , n44053 , n44054 );
and ( n44056 , n387 , n390 );
xor ( n44057 , n43816 , n43817 );
and ( n44058 , n44057 , n43819 );
and ( n44059 , n43816 , n43817 );
or ( n44060 , n44058 , n44059 );
xor ( n44061 , n44056 , n44060 );
and ( n44062 , n388 , n389 );
xor ( n44063 , n388 , n44062 );
and ( n44064 , n386 , n391 );
xor ( n44065 , n44063 , n44064 );
xor ( n44066 , n44061 , n44065 );
buf ( n44067 , n44066 );
xor ( n44068 , n44055 , n44067 );
buf ( n44069 , n44068 );
and ( n44070 , n44051 , n44069 );
not ( n44071 , n44051 );
not ( n44072 , n44068 );
and ( n44073 , n44071 , n44072 );
nor ( n44074 , n44070 , n44073 );
buf ( n44075 , n44074 );
buf ( n44076 , n393 );
and ( n44077 , n44075 , n44076 );
buf ( n44078 , n44077 );
buf ( n44079 , n44078 );
xor ( n44080 , n44047 , n44079 );
buf ( n44081 , n44080 );
buf ( n44082 , n44081 );
xor ( n44083 , n44020 , n44082 );
buf ( n44084 , n43926 );
xor ( n44085 , n44083 , n44084 );
buf ( n44086 , n44085 );
buf ( n44087 , n44086 );
xor ( n44088 , n44008 , n44009 );
xor ( n44089 , n44088 , n44087 );
buf ( n44090 , n44089 );
xor ( n44091 , n44008 , n44009 );
and ( n44092 , n44091 , n44087 );
and ( n44093 , n44008 , n44009 );
or ( n44094 , n44092 , n44093 );
buf ( n44095 , n44094 );
xor ( n44096 , n44037 , n44038 );
and ( n44097 , n44096 , n44040 );
and ( n44098 , n44037 , n44038 );
or ( n44099 , n44097 , n44098 );
buf ( n44100 , n44099 );
xor ( n44101 , n43987 , n43988 );
and ( n44102 , n44101 , n43990 );
and ( n44103 , n43987 , n43988 );
or ( n44104 , n44102 , n44103 );
buf ( n44105 , n44104 );
xor ( n44106 , n44030 , n44035 );
and ( n44107 , n44106 , n44043 );
and ( n44108 , n44030 , n44035 );
or ( n44109 , n44107 , n44108 );
buf ( n44110 , n44109 );
xor ( n44111 , n43978 , n43993 );
and ( n44112 , n44111 , n44000 );
and ( n44113 , n43978 , n43993 );
or ( n44114 , n44112 , n44113 );
buf ( n44115 , n44114 );
xor ( n44116 , n44014 , n44015 );
and ( n44117 , n44116 , n44017 );
and ( n44118 , n44014 , n44015 );
or ( n44119 , n44117 , n44118 );
buf ( n44120 , n44119 );
xor ( n44121 , n44025 , n44046 );
and ( n44122 , n44121 , n44079 );
and ( n44123 , n44025 , n44046 );
or ( n44124 , n44122 , n44123 );
buf ( n44125 , n44124 );
xor ( n44126 , n43977 , n44003 );
and ( n44127 , n44126 , n44005 );
and ( n44128 , n43977 , n44003 );
or ( n44129 , n44127 , n44128 );
buf ( n44130 , n44129 );
xor ( n44131 , n44020 , n44082 );
and ( n44132 , n44131 , n44084 );
and ( n44133 , n44020 , n44082 );
or ( n44134 , n44132 , n44133 );
buf ( n44135 , n44134 );
buf ( n44136 , n402 );
buf ( n44137 , n413 );
and ( n44138 , n44136 , n44137 );
buf ( n44139 , n44138 );
buf ( n44140 , n44139 );
buf ( n44141 , n403 );
buf ( n44142 , n412 );
and ( n44143 , n44141 , n44142 );
buf ( n44144 , n44143 );
buf ( n44145 , n44144 );
buf ( n44146 , n404 );
buf ( n44147 , n411 );
and ( n44148 , n44146 , n44147 );
buf ( n44149 , n44148 );
buf ( n44150 , n44149 );
xor ( n44151 , n44140 , n44145 );
xor ( n44152 , n44151 , n44150 );
buf ( n44153 , n44152 );
xor ( n44154 , n44140 , n44145 );
and ( n44155 , n44154 , n44150 );
and ( n44156 , n44140 , n44145 );
or ( n44157 , n44155 , n44156 );
buf ( n44158 , n44157 );
buf ( n44159 , n405 );
buf ( n44160 , n410 );
and ( n44161 , n44159 , n44160 );
buf ( n44162 , n44161 );
buf ( n44163 , n44162 );
and ( n44164 , n43959 , n43964 );
buf ( n44165 , n44164 );
buf ( n44166 , n44165 );
buf ( n44167 , n43949 );
xor ( n44168 , n44163 , n44166 );
xor ( n44169 , n44168 , n44167 );
buf ( n44170 , n44169 );
xor ( n44171 , n44163 , n44166 );
and ( n44172 , n44171 , n44167 );
and ( n44173 , n44163 , n44166 );
or ( n44174 , n44172 , n44173 );
buf ( n44175 , n44174 );
buf ( n44176 , n44120 );
buf ( n44177 , n44105 );
buf ( n44178 , n42914 );
buf ( n44179 , n386 );
and ( n44180 , n44178 , n44179 );
buf ( n44181 , n44180 );
buf ( n44182 , n44181 );
buf ( n44183 , n43054 );
buf ( n44184 , n387 );
and ( n44185 , n44183 , n44184 );
buf ( n44186 , n44185 );
buf ( n44187 , n44186 );
xor ( n44188 , n44182 , n44187 );
buf ( n44189 , n43222 );
buf ( n44190 , n388 );
and ( n44191 , n44189 , n44190 );
buf ( n44192 , n44191 );
buf ( n44193 , n44192 );
xor ( n44194 , n44188 , n44193 );
buf ( n44195 , n44194 );
buf ( n44196 , n44195 );
xor ( n44197 , n44177 , n44196 );
and ( n44198 , n390 , n43619 );
buf ( n44199 , n44198 );
xor ( n44200 , n44197 , n44199 );
buf ( n44201 , n44200 );
buf ( n44202 , n44201 );
xor ( n44203 , n44176 , n44202 );
buf ( n44204 , n44125 );
xor ( n44205 , n44203 , n44204 );
buf ( n44206 , n44205 );
buf ( n44207 , n44206 );
buf ( n44208 , n44135 );
buf ( n44209 , n44110 );
buf ( n44210 , n43838 );
buf ( n44211 , n391 );
and ( n44212 , n44210 , n44211 );
buf ( n44213 , n44212 );
buf ( n44214 , n44213 );
xor ( n44215 , n44209 , n44214 );
buf ( n44216 , n44074 );
buf ( n44217 , n392 );
and ( n44218 , n44216 , n44217 );
buf ( n44219 , n44218 );
buf ( n44220 , n44219 );
xor ( n44221 , n44215 , n44220 );
buf ( n44222 , n44221 );
buf ( n44223 , n44222 );
buf ( n44224 , n44115 );
not ( n44225 , n43821 );
not ( n44226 , n43826 );
and ( n44227 , n44225 , n44226 );
nor ( n44228 , n44066 , n44055 );
nor ( n44229 , n44227 , n44228 );
not ( n44230 , n44229 );
not ( n44231 , n43808 );
or ( n44232 , n44230 , n44231 );
not ( n44233 , n44066 );
not ( n44234 , n44055 );
nand ( n44235 , n44233 , n44234 );
not ( n44236 , n43821 );
nor ( n44237 , n44236 , n43827 );
and ( n44238 , n44235 , n44237 );
nor ( n44239 , n44233 , n44234 );
nor ( n44240 , n44238 , n44239 );
nand ( n44241 , n44232 , n44240 );
buf ( n44242 , n44241 );
and ( n44243 , n387 , n389 );
and ( n44244 , n386 , n390 );
xor ( n44245 , n44243 , n44244 );
xor ( n44246 , n388 , n44062 );
and ( n44247 , n44246 , n44064 );
and ( n44248 , n388 , n44062 );
or ( n44249 , n44247 , n44248 );
xor ( n44250 , n44245 , n44249 );
xor ( n44251 , n44056 , n44060 );
and ( n44252 , n44251 , n44065 );
and ( n44253 , n44056 , n44060 );
or ( n44254 , n44252 , n44253 );
not ( n44255 , n44254 );
and ( n44256 , n44250 , n44255 );
not ( n44257 , n44250 );
and ( n44258 , n44257 , n44254 );
nor ( n44259 , n44256 , n44258 );
not ( n44260 , n44259 );
and ( n44261 , n44242 , n44260 );
not ( n44262 , n44242 );
and ( n44263 , n44262 , n44259 );
nor ( n44264 , n44261 , n44263 );
buf ( n44265 , n44264 );
buf ( n44266 , n393 );
and ( n44267 , n44265 , n44266 );
buf ( n44268 , n44267 );
buf ( n44269 , n44268 );
xor ( n44270 , n44224 , n44269 );
buf ( n44271 , n44100 );
buf ( n44272 , n44153 );
buf ( n44273 , n43976 );
xor ( n44274 , n44272 , n44273 );
buf ( n44275 , n44170 );
xor ( n44276 , n44274 , n44275 );
buf ( n44277 , n44276 );
buf ( n44278 , n44277 );
xor ( n44279 , n44271 , n44278 );
buf ( n44280 , n43998 );
buf ( n44281 , n43366 );
nor ( n44282 , n44280 , n44281 );
buf ( n44283 , n44282 );
buf ( n44284 , n44283 );
xor ( n44285 , n44279 , n44284 );
buf ( n44286 , n44285 );
buf ( n44287 , n44286 );
xor ( n44288 , n44270 , n44287 );
buf ( n44289 , n44288 );
buf ( n44290 , n44289 );
xor ( n44291 , n44223 , n44290 );
buf ( n44292 , n44130 );
xor ( n44293 , n44291 , n44292 );
buf ( n44294 , n44293 );
buf ( n44295 , n44294 );
xor ( n44296 , n44207 , n44208 );
xor ( n44297 , n44296 , n44295 );
buf ( n44298 , n44297 );
xor ( n44299 , n44207 , n44208 );
and ( n44300 , n44299 , n44295 );
and ( n44301 , n44207 , n44208 );
or ( n44302 , n44300 , n44301 );
buf ( n44303 , n44302 );
xor ( n44304 , n44272 , n44273 );
and ( n44305 , n44304 , n44275 );
and ( n44306 , n44272 , n44273 );
or ( n44307 , n44305 , n44306 );
buf ( n44308 , n44307 );
xor ( n44309 , n44182 , n44187 );
and ( n44310 , n44309 , n44193 );
and ( n44311 , n44182 , n44187 );
or ( n44312 , n44310 , n44311 );
buf ( n44313 , n44312 );
xor ( n44314 , n44271 , n44278 );
and ( n44315 , n44314 , n44284 );
and ( n44316 , n44271 , n44278 );
or ( n44317 , n44315 , n44316 );
buf ( n44318 , n44317 );
xor ( n44319 , n44177 , n44196 );
and ( n44320 , n44319 , n44199 );
and ( n44321 , n44177 , n44196 );
or ( n44322 , n44320 , n44321 );
buf ( n44323 , n44322 );
xor ( n44324 , n44209 , n44214 );
and ( n44325 , n44324 , n44220 );
and ( n44326 , n44209 , n44214 );
or ( n44327 , n44325 , n44326 );
buf ( n44328 , n44327 );
xor ( n44329 , n44224 , n44269 );
and ( n44330 , n44329 , n44287 );
and ( n44331 , n44224 , n44269 );
or ( n44332 , n44330 , n44331 );
buf ( n44333 , n44332 );
xor ( n44334 , n44176 , n44202 );
and ( n44335 , n44334 , n44204 );
and ( n44336 , n44176 , n44202 );
or ( n44337 , n44335 , n44336 );
buf ( n44338 , n44337 );
xor ( n44339 , n44223 , n44290 );
and ( n44340 , n44339 , n44292 );
and ( n44341 , n44223 , n44290 );
or ( n44342 , n44340 , n44341 );
buf ( n44343 , n44342 );
buf ( n44344 , n402 );
buf ( n44345 , n412 );
and ( n44346 , n44344 , n44345 );
buf ( n44347 , n44346 );
buf ( n44348 , n44347 );
buf ( n44349 , n403 );
buf ( n44350 , n411 );
and ( n44351 , n44349 , n44350 );
buf ( n44352 , n44351 );
buf ( n44353 , n44352 );
buf ( n44354 , n404 );
buf ( n44355 , n410 );
and ( n44356 , n44354 , n44355 );
buf ( n44357 , n44356 );
buf ( n44358 , n44357 );
xor ( n44359 , n44348 , n44353 );
xor ( n44360 , n44359 , n44358 );
buf ( n44361 , n44360 );
xor ( n44362 , n44348 , n44353 );
and ( n44363 , n44362 , n44358 );
and ( n44364 , n44348 , n44353 );
or ( n44365 , n44363 , n44364 );
buf ( n44366 , n44365 );
buf ( n44367 , n44158 );
buf ( n44368 , n44361 );
buf ( n44369 , n44175 );
xor ( n44370 , n44367 , n44368 );
xor ( n44371 , n44370 , n44369 );
buf ( n44372 , n44371 );
xor ( n44373 , n44367 , n44368 );
and ( n44374 , n44373 , n44369 );
and ( n44375 , n44367 , n44368 );
or ( n44376 , n44374 , n44375 );
buf ( n44377 , n44376 );
buf ( n44378 , n43054 );
buf ( n44379 , n386 );
and ( n44380 , n44378 , n44379 );
buf ( n44381 , n44380 );
buf ( n44382 , n44381 );
buf ( n44383 , n43222 );
buf ( n44384 , n387 );
and ( n44385 , n44383 , n44384 );
buf ( n44386 , n44385 );
buf ( n44387 , n44386 );
buf ( n44388 , n44308 );
xor ( n44389 , n44382 , n44387 );
xor ( n44390 , n44389 , n44388 );
buf ( n44391 , n44390 );
xor ( n44392 , n44382 , n44387 );
and ( n44393 , n44392 , n44388 );
and ( n44394 , n44382 , n44387 );
or ( n44395 , n44393 , n44394 );
buf ( n44396 , n44395 );
buf ( n44397 , n44372 );
buf ( n44398 , n43346 );
buf ( n44399 , n388 );
and ( n44400 , n44398 , n44399 );
buf ( n44401 , n44400 );
buf ( n44402 , n44401 );
buf ( n44403 , n44313 );
xor ( n44404 , n44397 , n44402 );
xor ( n44405 , n44404 , n44403 );
buf ( n44406 , n44405 );
xor ( n44407 , n44397 , n44402 );
and ( n44408 , n44407 , n44403 );
and ( n44409 , n44397 , n44402 );
or ( n44410 , n44408 , n44409 );
buf ( n44411 , n44410 );
and ( n44412 , n43620 , n389 );
buf ( n44413 , n44412 );
buf ( n44414 , n44391 );
buf ( n44415 , n43838 );
buf ( n44416 , n390 );
and ( n44417 , n44415 , n44416 );
buf ( n44418 , n44417 );
buf ( n44419 , n44418 );
xor ( n44420 , n44413 , n44414 );
xor ( n44421 , n44420 , n44419 );
buf ( n44422 , n44421 );
xor ( n44423 , n44413 , n44414 );
and ( n44424 , n44423 , n44419 );
and ( n44425 , n44413 , n44414 );
or ( n44426 , n44424 , n44425 );
buf ( n44427 , n44426 );
buf ( n44428 , n44318 );
and ( n44429 , n44074 , n391 );
buf ( n44430 , n44429 );
buf ( n44431 , n44406 );
xor ( n44432 , n44428 , n44430 );
xor ( n44433 , n44432 , n44431 );
buf ( n44434 , n44433 );
xor ( n44435 , n44428 , n44430 );
and ( n44436 , n44435 , n44431 );
and ( n44437 , n44428 , n44430 );
or ( n44438 , n44436 , n44437 );
buf ( n44439 , n44438 );
buf ( n44440 , n44323 );
not ( n44441 , n44250 );
nand ( n44442 , n44441 , n44255 );
not ( n44443 , n44442 );
not ( n44444 , n44241 );
or ( n44445 , n44443 , n44444 );
nand ( n44446 , n44250 , n44254 );
buf ( n44447 , n44446 );
nand ( n44448 , n44445 , n44447 );
and ( n44449 , n387 , n388 );
xor ( n44450 , n387 , n44449 );
and ( n44451 , n386 , n389 );
xor ( n44452 , n44450 , n44451 );
not ( n44453 , n44452 );
xor ( n44454 , n44243 , n44244 );
and ( n44455 , n44454 , n44249 );
and ( n44456 , n44243 , n44244 );
or ( n44457 , n44455 , n44456 );
not ( n44458 , n44457 );
or ( n44459 , n44453 , n44458 );
or ( n44460 , n44452 , n44457 );
nand ( n44461 , n44459 , n44460 );
not ( n44462 , n44461 );
and ( n44463 , n44448 , n44462 );
not ( n44464 , n44448 );
buf ( n44465 , n44461 );
and ( n44466 , n44464 , n44465 );
nor ( n44467 , n44463 , n44466 );
buf ( n44468 , n44467 );
buf ( n44469 , n44468 );
buf ( n44470 , n44469 );
buf ( n44471 , n44470 );
buf ( n44472 , n393 );
nand ( n44473 , n44471 , n44472 );
buf ( n44474 , n44473 );
buf ( n44475 , n44474 );
not ( n44476 , n44475 );
buf ( n44477 , n44476 );
buf ( n44478 , n44477 );
buf ( n44479 , n44264 );
not ( n44480 , n44479 );
buf ( n44481 , n43190 );
nor ( n44482 , n44480 , n44481 );
buf ( n44483 , n44482 );
buf ( n44484 , n44483 );
xor ( n44485 , n44440 , n44478 );
xor ( n44486 , n44485 , n44484 );
buf ( n44487 , n44486 );
xor ( n44488 , n44440 , n44478 );
and ( n44489 , n44488 , n44484 );
and ( n44490 , n44440 , n44478 );
or ( n44491 , n44489 , n44490 );
buf ( n44492 , n44491 );
buf ( n44493 , n44422 );
buf ( n44494 , n44328 );
buf ( n44495 , n44333 );
xor ( n44496 , n44493 , n44494 );
xor ( n44497 , n44496 , n44495 );
buf ( n44498 , n44497 );
xor ( n44499 , n44493 , n44494 );
and ( n44500 , n44499 , n44495 );
and ( n44501 , n44493 , n44494 );
or ( n44502 , n44500 , n44501 );
buf ( n44503 , n44502 );
buf ( n44504 , n44434 );
buf ( n44505 , n44487 );
buf ( n44506 , n44338 );
xor ( n44507 , n44504 , n44505 );
xor ( n44508 , n44507 , n44506 );
buf ( n44509 , n44508 );
xor ( n44510 , n44504 , n44505 );
and ( n44511 , n44510 , n44506 );
and ( n44512 , n44504 , n44505 );
or ( n44513 , n44511 , n44512 );
buf ( n44514 , n44513 );
buf ( n44515 , n44498 );
buf ( n44516 , n44343 );
buf ( n44517 , n44509 );
xor ( n44518 , n44515 , n44516 );
xor ( n44519 , n44518 , n44517 );
buf ( n44520 , n44519 );
xor ( n44521 , n44515 , n44516 );
and ( n44522 , n44521 , n44517 );
and ( n44523 , n44515 , n44516 );
or ( n44524 , n44522 , n44523 );
buf ( n44525 , n44524 );
buf ( n44526 , n402 );
buf ( n44527 , n411 );
and ( n44528 , n44526 , n44527 );
buf ( n44529 , n44528 );
buf ( n44530 , n44529 );
buf ( n44531 , n403 );
buf ( n44532 , n410 );
and ( n44533 , n44531 , n44532 );
buf ( n44534 , n44533 );
buf ( n44535 , n44534 );
buf ( n44536 , n44366 );
xor ( n44537 , n44530 , n44535 );
xor ( n44538 , n44537 , n44536 );
buf ( n44539 , n44538 );
xor ( n44540 , n44530 , n44535 );
and ( n44541 , n44540 , n44536 );
and ( n44542 , n44530 , n44535 );
or ( n44543 , n44541 , n44542 );
buf ( n44544 , n44543 );
buf ( n44545 , n44539 );
buf ( n44546 , n43222 );
buf ( n44547 , n386 );
and ( n44548 , n44546 , n44547 );
buf ( n44549 , n44548 );
buf ( n44550 , n44549 );
buf ( n44551 , n44377 );
xor ( n44552 , n44545 , n44550 );
xor ( n44553 , n44552 , n44551 );
buf ( n44554 , n44553 );
xor ( n44555 , n44545 , n44550 );
and ( n44556 , n44555 , n44551 );
and ( n44557 , n44545 , n44550 );
or ( n44558 , n44556 , n44557 );
buf ( n44559 , n44558 );
buf ( n44560 , n43346 );
buf ( n44561 , n387 );
and ( n44562 , n44560 , n44561 );
buf ( n44563 , n44562 );
buf ( n44564 , n44563 );
and ( n44565 , n43620 , n388 );
buf ( n44566 , n44565 );
buf ( n44567 , n44396 );
xor ( n44568 , n44564 , n44566 );
xor ( n44569 , n44568 , n44567 );
buf ( n44570 , n44569 );
xor ( n44571 , n44564 , n44566 );
and ( n44572 , n44571 , n44567 );
and ( n44573 , n44564 , n44566 );
or ( n44574 , n44572 , n44573 );
buf ( n44575 , n44574 );
buf ( n44576 , n43835 );
buf ( n44577 , n389 );
and ( n44578 , n44576 , n44577 );
buf ( n44579 , n44578 );
buf ( n44580 , n44579 );
buf ( n44581 , n44554 );
and ( n44582 , n44051 , n44069 );
not ( n44583 , n44051 );
and ( n44584 , n44583 , n44072 );
nor ( n44585 , n44582 , n44584 );
buf ( n44586 , n44585 );
buf ( n44587 , n390 );
and ( n44588 , n44586 , n44587 );
buf ( n44589 , n44588 );
buf ( n44590 , n44589 );
xor ( n44591 , n44580 , n44581 );
xor ( n44592 , n44591 , n44590 );
buf ( n44593 , n44592 );
xor ( n44594 , n44580 , n44581 );
and ( n44595 , n44594 , n44590 );
and ( n44596 , n44580 , n44581 );
or ( n44597 , n44595 , n44596 );
buf ( n44598 , n44597 );
buf ( n44599 , n44467 );
buf ( n44600 , n392 );
and ( n44601 , n44599 , n44600 );
buf ( n44602 , n44601 );
buf ( n44603 , n44602 );
buf ( n44604 , n44264 );
buf ( n44605 , n391 );
and ( n44606 , n44604 , n44605 );
buf ( n44607 , n44606 );
buf ( n44608 , n44607 );
buf ( n44609 , n44411 );
xor ( n44610 , n44603 , n44608 );
xor ( n44611 , n44610 , n44609 );
buf ( n44612 , n44611 );
xor ( n44613 , n44603 , n44608 );
and ( n44614 , n44613 , n44609 );
and ( n44615 , n44603 , n44608 );
or ( n44616 , n44614 , n44615 );
buf ( n44617 , n44616 );
buf ( n44618 , n44570 );
buf ( n44619 , n44427 );
not ( n44620 , n44460 );
not ( n44621 , n44442 );
not ( n44622 , n44241 );
or ( n44623 , n44621 , n44622 );
nand ( n44624 , n44623 , n44446 );
not ( n44625 , n44624 );
or ( n44626 , n44620 , n44625 );
nand ( n44627 , n44457 , n44452 );
nand ( n44628 , n44626 , n44627 );
xor ( n44629 , n387 , n44449 );
and ( n44630 , n44629 , n44451 );
and ( n44631 , n387 , n44449 );
or ( n44632 , n44630 , n44631 );
and ( n44633 , n386 , n388 );
nor ( n44634 , n44632 , n44633 );
not ( n44635 , n44634 );
nand ( n44636 , n44632 , n44633 );
nand ( n44637 , n44635 , n44636 );
not ( n44638 , n44637 );
and ( n44639 , n44628 , n44638 );
not ( n44640 , n44628 );
and ( n44641 , n44640 , n44637 );
nor ( n44642 , n44639 , n44641 );
buf ( n44643 , n44642 );
buf ( n44644 , n393 );
and ( n44645 , n44643 , n44644 );
buf ( n44646 , n44645 );
buf ( n44647 , n44646 );
xor ( n44648 , n44618 , n44619 );
xor ( n44649 , n44648 , n44647 );
buf ( n44650 , n44649 );
xor ( n44651 , n44618 , n44619 );
and ( n44652 , n44651 , n44647 );
and ( n44653 , n44618 , n44619 );
or ( n44654 , n44652 , n44653 );
buf ( n44655 , n44654 );
buf ( n44656 , n44593 );
buf ( n44657 , n44492 );
buf ( n44658 , n44439 );
xor ( n44659 , n44656 , n44657 );
xor ( n44660 , n44659 , n44658 );
buf ( n44661 , n44660 );
xor ( n44662 , n44656 , n44657 );
and ( n44663 , n44662 , n44658 );
and ( n44664 , n44656 , n44657 );
or ( n44665 , n44663 , n44664 );
buf ( n44666 , n44665 );
buf ( n44667 , n44612 );
buf ( n44668 , n44650 );
buf ( n44669 , n44503 );
xor ( n44670 , n44667 , n44668 );
xor ( n44671 , n44670 , n44669 );
buf ( n44672 , n44671 );
xor ( n44673 , n44667 , n44668 );
and ( n44674 , n44673 , n44669 );
and ( n44675 , n44667 , n44668 );
or ( n44676 , n44674 , n44675 );
buf ( n44677 , n44676 );
buf ( n44678 , n44661 );
buf ( n44679 , n44514 );
buf ( n44680 , n44672 );
xor ( n44681 , n44678 , n44679 );
xor ( n44682 , n44681 , n44680 );
buf ( n44683 , n44682 );
xor ( n44684 , n44678 , n44679 );
and ( n44685 , n44684 , n44680 );
and ( n44686 , n44678 , n44679 );
or ( n44687 , n44685 , n44686 );
buf ( n44688 , n44687 );
buf ( n44689 , n402 );
buf ( n44690 , n410 );
and ( n44691 , n44689 , n44690 );
buf ( n44692 , n44691 );
buf ( n44693 , n44692 );
buf ( n44694 , n44544 );
buf ( n44695 , n386 );
not ( n44696 , n44695 );
buf ( n44697 , n43998 );
nor ( n44698 , n44696 , n44697 );
buf ( n44699 , n44698 );
buf ( n44700 , n44699 );
xor ( n44701 , n44693 , n44694 );
xor ( n44702 , n44701 , n44700 );
buf ( n44703 , n44702 );
xor ( n44704 , n44693 , n44694 );
and ( n44705 , n44704 , n44700 );
and ( n44706 , n44693 , n44694 );
or ( n44707 , n44705 , n44706 );
buf ( n44708 , n44707 );
buf ( n44709 , n43619 );
not ( n44710 , n44709 );
buf ( n44711 , n43983 );
nor ( n44712 , n44710 , n44711 );
buf ( n44713 , n44712 );
buf ( n44714 , n44713 );
buf ( n44715 , n43835 );
buf ( n44716 , n388 );
and ( n44717 , n44715 , n44716 );
buf ( n44718 , n44717 );
buf ( n44719 , n44718 );
buf ( n44720 , n44559 );
xor ( n44721 , n44714 , n44719 );
xor ( n44722 , n44721 , n44720 );
buf ( n44723 , n44722 );
xor ( n44724 , n44714 , n44719 );
and ( n44725 , n44724 , n44720 );
and ( n44726 , n44714 , n44719 );
or ( n44727 , n44725 , n44726 );
buf ( n44728 , n44727 );
buf ( n44729 , n44703 );
buf ( n44730 , n44074 );
buf ( n44731 , n389 );
and ( n44732 , n44730 , n44731 );
buf ( n44733 , n44732 );
buf ( n44734 , n44733 );
and ( n44735 , n44242 , n44260 );
not ( n44736 , n44242 );
and ( n44737 , n44736 , n44259 );
nor ( n44738 , n44735 , n44737 );
buf ( n44739 , n44738 );
buf ( n44740 , n390 );
and ( n44741 , n44739 , n44740 );
buf ( n44742 , n44741 );
buf ( n44743 , n44742 );
xor ( n44744 , n44729 , n44734 );
xor ( n44745 , n44744 , n44743 );
buf ( n44746 , n44745 );
xor ( n44747 , n44729 , n44734 );
and ( n44748 , n44747 , n44743 );
and ( n44749 , n44729 , n44734 );
or ( n44750 , n44748 , n44749 );
buf ( n44751 , n44750 );
buf ( n44752 , n44467 );
buf ( n44753 , n391 );
and ( n44754 , n44752 , n44753 );
buf ( n44755 , n44754 );
buf ( n44756 , n44755 );
not ( n44757 , n393 );
and ( n44758 , n43983 , n386 );
nor ( n44759 , n44757 , n44758 );
not ( n44760 , n44759 );
not ( n44761 , n44452 );
not ( n44762 , n44457 );
and ( n44763 , n44761 , n44762 );
nor ( n44764 , n44763 , n44634 );
not ( n44765 , n44764 );
not ( n44766 , n44624 );
or ( n44767 , n44765 , n44766 );
not ( n44768 , n44627 );
not ( n44769 , n44634 );
and ( n44770 , n44768 , n44769 );
not ( n44771 , n44636 );
nor ( n44772 , n44770 , n44771 );
nand ( n44773 , n44767 , n44772 );
not ( n44774 , n44773 );
or ( n44775 , n44760 , n44774 );
nand ( n44776 , n44624 , n44764 );
and ( n44777 , n44758 , n393 );
nand ( n44778 , n44776 , n44772 , n44777 );
nand ( n44779 , n44775 , n44778 );
buf ( n44780 , n44779 );
buf ( n44781 , n44575 );
xor ( n44782 , n44756 , n44780 );
xor ( n44783 , n44782 , n44781 );
buf ( n44784 , n44783 );
xor ( n44785 , n44756 , n44780 );
and ( n44786 , n44785 , n44781 );
and ( n44787 , n44756 , n44780 );
or ( n44788 , n44786 , n44787 );
buf ( n44789 , n44788 );
buf ( n44790 , n44598 );
and ( n44791 , n44642 , n392 );
buf ( n44792 , n44791 );
buf ( n44793 , n44723 );
xor ( n44794 , n44790 , n44792 );
xor ( n44795 , n44794 , n44793 );
buf ( n44796 , n44795 );
xor ( n44797 , n44790 , n44792 );
and ( n44798 , n44797 , n44793 );
and ( n44799 , n44790 , n44792 );
or ( n44800 , n44798 , n44799 );
buf ( n44801 , n44800 );
buf ( n44802 , n44617 );
buf ( n44803 , n44746 );
buf ( n44804 , n44655 );
xor ( n44805 , n44802 , n44803 );
xor ( n44806 , n44805 , n44804 );
buf ( n44807 , n44806 );
xor ( n44808 , n44802 , n44803 );
and ( n44809 , n44808 , n44804 );
and ( n44810 , n44802 , n44803 );
or ( n44811 , n44809 , n44810 );
buf ( n44812 , n44811 );
buf ( n44813 , n44784 );
buf ( n44814 , n44796 );
buf ( n44815 , n44666 );
xor ( n44816 , n44813 , n44814 );
xor ( n44817 , n44816 , n44815 );
buf ( n44818 , n44817 );
xor ( n44819 , n44813 , n44814 );
and ( n44820 , n44819 , n44815 );
and ( n44821 , n44813 , n44814 );
or ( n44822 , n44820 , n44821 );
buf ( n44823 , n44822 );
buf ( n44824 , n44807 );
buf ( n44825 , n44677 );
buf ( n44826 , n44818 );
xor ( n44827 , n44824 , n44825 );
xor ( n44828 , n44827 , n44826 );
buf ( n44829 , n44828 );
xor ( n44830 , n44824 , n44825 );
and ( n44831 , n44830 , n44826 );
and ( n44832 , n44824 , n44825 );
or ( n44833 , n44831 , n44832 );
buf ( n44834 , n44833 );
and ( n44835 , n386 , n43620 );
buf ( n44836 , n44835 );
buf ( n44837 , n43838 );
buf ( n44838 , n387 );
and ( n44839 , n44837 , n44838 );
buf ( n44840 , n44839 );
buf ( n44841 , n44840 );
buf ( n44842 , n44585 );
buf ( n44843 , n388 );
and ( n44844 , n44842 , n44843 );
buf ( n44845 , n44844 );
buf ( n44846 , n44845 );
xor ( n44847 , n44836 , n44841 );
xor ( n44848 , n44847 , n44846 );
buf ( n44849 , n44848 );
xor ( n44850 , n44836 , n44841 );
and ( n44851 , n44850 , n44846 );
and ( n44852 , n44836 , n44841 );
or ( n44853 , n44851 , n44852 );
buf ( n44854 , n44853 );
buf ( n44855 , n44708 );
buf ( n44856 , n44470 );
buf ( n44857 , n390 );
nand ( n44858 , n44856 , n44857 );
buf ( n44859 , n44858 );
buf ( n44860 , n44859 );
not ( n44861 , n44860 );
buf ( n44862 , n44861 );
buf ( n44863 , n44862 );
buf ( n44864 , n44264 );
buf ( n44865 , n389 );
and ( n44866 , n44864 , n44865 );
buf ( n44867 , n44866 );
buf ( n44868 , n44867 );
xor ( n44869 , n44855 , n44863 );
xor ( n44870 , n44869 , n44868 );
buf ( n44871 , n44870 );
xor ( n44872 , n44855 , n44863 );
and ( n44873 , n44872 , n44868 );
and ( n44874 , n44855 , n44863 );
or ( n44875 , n44873 , n44874 );
buf ( n44876 , n44875 );
and ( n44877 , n44764 , n386 );
not ( n44878 , n44877 );
not ( n44879 , n44448 );
or ( n44880 , n44878 , n44879 );
not ( n44881 , n43983 );
not ( n44882 , n44772 );
or ( n44883 , n44881 , n44882 );
nand ( n44884 , n44883 , n386 );
nand ( n44885 , n44880 , n44884 );
buf ( n44886 , n44885 );
buf ( n44887 , n393 );
and ( n44888 , n44886 , n44887 );
buf ( n44889 , n44888 );
buf ( n44890 , n44889 );
buf ( n44891 , n44728 );
xnor ( n44892 , n44773 , n44758 );
nor ( n44893 , n44892 , n43190 );
buf ( n44894 , n44893 );
xor ( n44895 , n44890 , n44891 );
xor ( n44896 , n44895 , n44894 );
buf ( n44897 , n44896 );
xor ( n44898 , n44890 , n44891 );
and ( n44899 , n44898 , n44894 );
and ( n44900 , n44890 , n44891 );
or ( n44901 , n44899 , n44900 );
buf ( n44902 , n44901 );
buf ( n44903 , n44849 );
buf ( n44904 , n44642 );
buf ( n44905 , n391 );
and ( n44906 , n44904 , n44905 );
buf ( n44907 , n44906 );
buf ( n44908 , n44907 );
buf ( n44909 , n44751 );
xor ( n44910 , n44903 , n44908 );
xor ( n44911 , n44910 , n44909 );
buf ( n44912 , n44911 );
xor ( n44913 , n44903 , n44908 );
and ( n44914 , n44913 , n44909 );
and ( n44915 , n44903 , n44908 );
or ( n44916 , n44914 , n44915 );
buf ( n44917 , n44916 );
buf ( n44918 , n44789 );
buf ( n44919 , n44871 );
buf ( n44920 , n44897 );
xor ( n44921 , n44918 , n44919 );
xor ( n44922 , n44921 , n44920 );
buf ( n44923 , n44922 );
xor ( n44924 , n44918 , n44919 );
and ( n44925 , n44924 , n44920 );
and ( n44926 , n44918 , n44919 );
or ( n44927 , n44925 , n44926 );
buf ( n44928 , n44927 );
buf ( n44929 , n44801 );
buf ( n44930 , n44912 );
buf ( n44931 , n44812 );
xor ( n44932 , n44929 , n44930 );
xor ( n44933 , n44932 , n44931 );
buf ( n44934 , n44933 );
xor ( n44935 , n44929 , n44930 );
and ( n44936 , n44935 , n44931 );
and ( n44937 , n44929 , n44930 );
or ( n44938 , n44936 , n44937 );
buf ( n44939 , n44938 );
buf ( n44940 , n44923 );
buf ( n44941 , n44823 );
buf ( n44942 , n44934 );
xor ( n44943 , n44940 , n44941 );
xor ( n44944 , n44943 , n44942 );
buf ( n44945 , n44944 );
xor ( n44946 , n44940 , n44941 );
and ( n44947 , n44946 , n44942 );
and ( n44948 , n44940 , n44941 );
or ( n44949 , n44947 , n44948 );
buf ( n44950 , n44949 );
buf ( n44951 , n43838 );
buf ( n44952 , n386 );
and ( n44953 , n44951 , n44952 );
buf ( n44954 , n44953 );
buf ( n44955 , n44954 );
buf ( n44956 , n44585 );
buf ( n44957 , n387 );
and ( n44958 , n44956 , n44957 );
buf ( n44959 , n44958 );
buf ( n44960 , n44959 );
buf ( n44961 , n44885 );
buf ( n44962 , n392 );
and ( n44963 , n44961 , n44962 );
buf ( n44964 , n44963 );
buf ( n44965 , n44964 );
xor ( n44966 , n44955 , n44960 );
xor ( n44967 , n44966 , n44965 );
buf ( n44968 , n44967 );
xor ( n44969 , n44955 , n44960 );
and ( n44970 , n44969 , n44965 );
and ( n44971 , n44955 , n44960 );
or ( n44972 , n44970 , n44971 );
buf ( n44973 , n44972 );
buf ( n44974 , n44470 );
buf ( n44975 , n389 );
and ( n44976 , n44974 , n44975 );
buf ( n44977 , n44976 );
buf ( n44978 , n44977 );
buf ( n44979 , n44738 );
buf ( n44980 , n388 );
and ( n44981 , n44979 , n44980 );
buf ( n44982 , n44981 );
buf ( n44983 , n44982 );
not ( n44984 , n44758 );
not ( n44985 , n44773 );
not ( n44986 , n44985 );
or ( n44987 , n44984 , n44986 );
or ( n44988 , n44985 , n44758 );
nand ( n44989 , n44987 , n44988 );
buf ( n44990 , n44989 );
buf ( n44991 , n391 );
and ( n44992 , n44990 , n44991 );
buf ( n44993 , n44992 );
buf ( n44994 , n44993 );
xor ( n44995 , n44978 , n44983 );
xor ( n44996 , n44995 , n44994 );
buf ( n44997 , n44996 );
xor ( n44998 , n44978 , n44983 );
and ( n44999 , n44998 , n44994 );
and ( n45000 , n44978 , n44983 );
or ( n45001 , n44999 , n45000 );
buf ( n45002 , n45001 );
and ( n45003 , n44642 , n390 );
buf ( n45004 , n45003 );
buf ( n45005 , n44854 );
buf ( n45006 , n44876 );
xor ( n45007 , n45004 , n45005 );
xor ( n45008 , n45007 , n45006 );
buf ( n45009 , n45008 );
xor ( n45010 , n45004 , n45005 );
and ( n45011 , n45010 , n45006 );
and ( n45012 , n45004 , n45005 );
or ( n45013 , n45011 , n45012 );
buf ( n45014 , n45013 );
buf ( n45015 , n44968 );
buf ( n45016 , n44902 );
buf ( n45017 , n44997 );
xor ( n45018 , n45015 , n45016 );
xor ( n45019 , n45018 , n45017 );
buf ( n45020 , n45019 );
xor ( n45021 , n45015 , n45016 );
and ( n45022 , n45021 , n45017 );
and ( n45023 , n45015 , n45016 );
or ( n45024 , n45022 , n45023 );
buf ( n45025 , n45024 );
buf ( n45026 , n45009 );
buf ( n45027 , n44917 );
buf ( n45028 , n44928 );
xor ( n45029 , n45026 , n45027 );
xor ( n45030 , n45029 , n45028 );
buf ( n45031 , n45030 );
xor ( n45032 , n45026 , n45027 );
and ( n45033 , n45032 , n45028 );
and ( n45034 , n45026 , n45027 );
or ( n45035 , n45033 , n45034 );
buf ( n45036 , n45035 );
buf ( n45037 , n45020 );
buf ( n45038 , n45031 );
buf ( n45039 , n44939 );
xor ( n45040 , n45037 , n45038 );
xor ( n45041 , n45040 , n45039 );
buf ( n45042 , n45041 );
xor ( n45043 , n45037 , n45038 );
and ( n45044 , n45043 , n45039 );
and ( n45045 , n45037 , n45038 );
or ( n45046 , n45044 , n45045 );
buf ( n45047 , n45046 );
buf ( n45048 , n44074 );
buf ( n45049 , n386 );
and ( n45050 , n45048 , n45049 );
buf ( n45051 , n45050 );
buf ( n45052 , n45051 );
buf ( n45053 , n44470 );
buf ( n45054 , n45053 );
buf ( n45055 , n45054 );
buf ( n45056 , n45055 );
buf ( n45057 , n388 );
nand ( n45058 , n45056 , n45057 );
buf ( n45059 , n45058 );
buf ( n45060 , n45059 );
not ( n45061 , n45060 );
buf ( n45062 , n45061 );
buf ( n45063 , n45062 );
buf ( n45064 , n44738 );
not ( n45065 , n45064 );
buf ( n45066 , n43983 );
nor ( n45067 , n45065 , n45066 );
buf ( n45068 , n45067 );
buf ( n45069 , n45068 );
xor ( n45070 , n45052 , n45063 );
xor ( n45071 , n45070 , n45069 );
buf ( n45072 , n45071 );
xor ( n45073 , n45052 , n45063 );
and ( n45074 , n45073 , n45069 );
and ( n45075 , n45052 , n45063 );
or ( n45076 , n45074 , n45075 );
buf ( n45077 , n45076 );
buf ( n45078 , n44885 );
buf ( n45079 , n45078 );
buf ( n45080 , n45079 );
buf ( n45081 , n45080 );
buf ( n45082 , n391 );
and ( n45083 , n45081 , n45082 );
buf ( n45084 , n45083 );
buf ( n45085 , n45084 );
and ( n45086 , n44989 , n390 );
buf ( n45087 , n45086 );
buf ( n45088 , n44642 );
buf ( n45089 , n389 );
and ( n45090 , n45088 , n45089 );
buf ( n45091 , n45090 );
buf ( n45092 , n45091 );
xor ( n45093 , n45085 , n45087 );
xor ( n45094 , n45093 , n45092 );
buf ( n45095 , n45094 );
xor ( n45096 , n45085 , n45087 );
and ( n45097 , n45096 , n45092 );
and ( n45098 , n45085 , n45087 );
or ( n45099 , n45097 , n45098 );
buf ( n45100 , n45099 );
buf ( n45101 , n44973 );
buf ( n45102 , n45002 );
buf ( n45103 , n45072 );
xor ( n45104 , n45101 , n45102 );
xor ( n45105 , n45104 , n45103 );
buf ( n45106 , n45105 );
xor ( n45107 , n45101 , n45102 );
and ( n45108 , n45107 , n45103 );
and ( n45109 , n45101 , n45102 );
or ( n45110 , n45108 , n45109 );
buf ( n45111 , n45110 );
buf ( n45112 , n45095 );
buf ( n45113 , n45014 );
buf ( n45114 , n45025 );
xor ( n45115 , n45112 , n45113 );
xor ( n45116 , n45115 , n45114 );
buf ( n45117 , n45116 );
xor ( n45118 , n45112 , n45113 );
and ( n45119 , n45118 , n45114 );
and ( n45120 , n45112 , n45113 );
or ( n45121 , n45119 , n45120 );
buf ( n45122 , n45121 );
buf ( n45123 , n45106 );
buf ( n45124 , n45117 );
buf ( n45125 , n45036 );
xor ( n45126 , n45123 , n45124 );
xor ( n45127 , n45126 , n45125 );
buf ( n45128 , n45127 );
xor ( n45129 , n45123 , n45124 );
and ( n45130 , n45129 , n45125 );
and ( n45131 , n45123 , n45124 );
or ( n45132 , n45130 , n45131 );
buf ( n45133 , n45132 );
buf ( n45134 , n45080 );
buf ( n45135 , n390 );
and ( n45136 , n45134 , n45135 );
buf ( n45137 , n45136 );
buf ( n45138 , n45137 );
buf ( n45139 , n44738 );
buf ( n45140 , n386 );
and ( n45141 , n45139 , n45140 );
buf ( n45142 , n45141 );
buf ( n45143 , n45142 );
buf ( n45144 , n45055 );
buf ( n45145 , n387 );
and ( n45146 , n45144 , n45145 );
buf ( n45147 , n45146 );
buf ( n45148 , n45147 );
xor ( n45149 , n45138 , n45143 );
xor ( n45150 , n45149 , n45148 );
buf ( n45151 , n45150 );
xor ( n45152 , n45138 , n45143 );
and ( n45153 , n45152 , n45148 );
and ( n45154 , n45138 , n45143 );
or ( n45155 , n45153 , n45154 );
buf ( n45156 , n45155 );
buf ( n45157 , n44989 );
buf ( n45158 , n389 );
and ( n45159 , n45157 , n45158 );
buf ( n45160 , n45159 );
buf ( n45161 , n45160 );
and ( n45162 , n44642 , n388 );
buf ( n45163 , n45162 );
buf ( n45164 , n45077 );
xor ( n45165 , n45161 , n45163 );
xor ( n45166 , n45165 , n45164 );
buf ( n45167 , n45166 );
xor ( n45168 , n45161 , n45163 );
and ( n45169 , n45168 , n45164 );
and ( n45170 , n45161 , n45163 );
or ( n45171 , n45169 , n45170 );
buf ( n45172 , n45171 );
buf ( n45173 , n45151 );
buf ( n45174 , n45100 );
buf ( n45175 , n45167 );
xor ( n45176 , n45173 , n45174 );
xor ( n45177 , n45176 , n45175 );
buf ( n45178 , n45177 );
xor ( n45179 , n45173 , n45174 );
and ( n45180 , n45179 , n45175 );
and ( n45181 , n45173 , n45174 );
or ( n45182 , n45180 , n45181 );
buf ( n45183 , n45182 );
buf ( n45184 , n45111 );
buf ( n45185 , n45178 );
buf ( n45186 , n45122 );
xor ( n45187 , n45184 , n45185 );
xor ( n45188 , n45187 , n45186 );
buf ( n45189 , n45188 );
xor ( n45190 , n45184 , n45185 );
and ( n45191 , n45190 , n45186 );
and ( n45192 , n45184 , n45185 );
or ( n45193 , n45191 , n45192 );
buf ( n45194 , n45193 );
buf ( n45195 , n45080 );
buf ( n45196 , n389 );
and ( n45197 , n45195 , n45196 );
buf ( n45198 , n45197 );
buf ( n45199 , n45198 );
buf ( n45200 , n45055 );
buf ( n45201 , n386 );
and ( n45202 , n45200 , n45201 );
buf ( n45203 , n45202 );
buf ( n45204 , n45203 );
buf ( n45205 , n44989 );
buf ( n45206 , n388 );
and ( n45207 , n45205 , n45206 );
buf ( n45208 , n45207 );
buf ( n45209 , n45208 );
xor ( n45210 , n45199 , n45204 );
xor ( n45211 , n45210 , n45209 );
buf ( n45212 , n45211 );
xor ( n45213 , n45199 , n45204 );
and ( n45214 , n45213 , n45209 );
and ( n45215 , n45199 , n45204 );
or ( n45216 , n45214 , n45215 );
buf ( n45217 , n45216 );
buf ( n45218 , n44642 );
buf ( n45219 , n387 );
and ( n45220 , n45218 , n45219 );
buf ( n45221 , n45220 );
buf ( n45222 , n45221 );
buf ( n45223 , n45156 );
buf ( n45224 , n45212 );
xor ( n45225 , n45222 , n45223 );
xor ( n45226 , n45225 , n45224 );
buf ( n45227 , n45226 );
xor ( n45228 , n45222 , n45223 );
and ( n45229 , n45228 , n45224 );
and ( n45230 , n45222 , n45223 );
or ( n45231 , n45229 , n45230 );
buf ( n45232 , n45231 );
buf ( n45233 , n45172 );
buf ( n45234 , n45227 );
buf ( n45235 , n45183 );
xor ( n45236 , n45233 , n45234 );
xor ( n45237 , n45236 , n45235 );
buf ( n45238 , n45237 );
xor ( n45239 , n45233 , n45234 );
and ( n45240 , n45239 , n45235 );
and ( n45241 , n45233 , n45234 );
or ( n45242 , n45240 , n45241 );
buf ( n45243 , n45242 );
buf ( n45244 , n45080 );
buf ( n45245 , n388 );
and ( n45246 , n45244 , n45245 );
buf ( n45247 , n45246 );
buf ( n45248 , n45247 );
buf ( n45249 , n44989 );
buf ( n45250 , n387 );
and ( n45251 , n45249 , n45250 );
buf ( n45252 , n45251 );
buf ( n45253 , n45252 );
buf ( n45254 , n44642 );
buf ( n45255 , n386 );
and ( n45256 , n45254 , n45255 );
buf ( n45257 , n45256 );
buf ( n45258 , n45257 );
xor ( n45259 , n45248 , n45253 );
xor ( n45260 , n45259 , n45258 );
buf ( n45261 , n45260 );
and ( n45262 , n45248 , n45253 );
or ( n45263 , C0 , n45262 );
buf ( n45264 , n45263 );
buf ( n45265 , n45217 );
buf ( n45266 , n45261 );
buf ( n45267 , n45232 );
xor ( n45268 , n45265 , n45266 );
xor ( n45269 , n45268 , n45267 );
buf ( n45270 , n45269 );
xor ( n45271 , n45265 , n45266 );
and ( n45272 , n45271 , n45267 );
and ( n45273 , n45265 , n45266 );
or ( n45274 , n45272 , n45273 );
buf ( n45275 , n45274 );
buf ( n45276 , n45080 );
buf ( n45277 , n387 );
and ( n45278 , n45276 , n45277 );
buf ( n45279 , n45278 );
buf ( n45280 , n45279 );
buf ( n45281 , n44989 );
buf ( n45282 , n386 );
and ( n45283 , n45281 , n45282 );
buf ( n45284 , n45283 );
buf ( n45285 , n45284 );
buf ( n45286 , n45264 );
xor ( n45287 , n45280 , n45285 );
xor ( n45288 , n45287 , n45286 );
buf ( n45289 , n45288 );
and ( n45290 , n45280 , n45285 );
or ( n45291 , C0 , n45290 );
buf ( n45292 , n45291 );
not ( n45293 , n45047 );
not ( n45294 , n45293 );
not ( n45295 , n45128 );
not ( n45296 , n45295 );
or ( n45297 , n45294 , n45296 );
not ( n45298 , n45128 );
not ( n45299 , n45047 );
or ( n45300 , n45298 , n45299 );
nand ( n45301 , n45042 , n44950 );
nand ( n45302 , n45300 , n45301 );
nand ( n45303 , n45297 , n45302 );
not ( n45304 , n45303 );
not ( n45305 , n45133 );
not ( n45306 , n45189 );
nand ( n45307 , n45305 , n45306 );
not ( n45308 , n45194 );
not ( n45309 , n45238 );
nand ( n45310 , n45308 , n45309 );
and ( n45311 , n45307 , n45310 );
and ( n45312 , n45304 , n45311 );
not ( n45313 , n45194 );
nand ( n45314 , n45313 , n45309 );
not ( n45315 , n45314 );
nand ( n45316 , n45189 , n45133 );
not ( n45317 , n45316 );
not ( n45318 , n45317 );
or ( n45319 , n45315 , n45318 );
not ( n45320 , n45309 );
nand ( n45321 , n45320 , n45194 );
nand ( n45322 , n45319 , n45321 );
nor ( n45323 , n45312 , n45322 );
buf ( n45324 , n45323 );
not ( n45325 , n45324 );
buf ( n45326 , n45325 );
not ( n45327 , n45293 );
not ( n45328 , n45295 );
or ( n45329 , n45327 , n45328 );
buf ( n45330 , n45042 );
not ( n45331 , n45330 );
buf ( n45332 , n45331 );
buf ( n45333 , n44950 );
not ( n45334 , n45333 );
buf ( n45335 , n45334 );
nand ( n45336 , n45332 , n45335 );
nand ( n45337 , n45329 , n45336 );
not ( n45338 , n45337 );
buf ( n45339 , n45338 );
buf ( n45340 , n45311 );
or ( n45341 , n45270 , n45243 );
buf ( n45342 , n45275 );
buf ( n45343 , n45289 );
or ( n45344 , n45342 , n45343 );
buf ( n45345 , n45344 );
nand ( n45346 , n45341 , n45345 );
not ( n45347 , n45292 );
buf ( n45348 , n45080 );
buf ( n45349 , n386 );
nand ( n45350 , n45348 , n45349 );
buf ( n45351 , n45350 );
nand ( n45352 , n45347 , n45351 );
not ( n45353 , n45352 );
nor ( n45354 , n45346 , n45353 );
buf ( n45355 , n45354 );
and ( n45356 , n45339 , n45340 , n45355 );
buf ( n45357 , n45356 );
buf ( n45358 , n45332 );
not ( n45359 , n45358 );
buf ( n45360 , n44950 );
nand ( n45361 , n45359 , n45360 );
buf ( n45362 , n45361 );
buf ( n45363 , n45362 );
buf ( n45364 , n45336 );
and ( n45365 , n45363 , n45364 );
buf ( n45366 , n45365 );
buf ( n45367 , n45362 );
not ( n45368 , n45367 );
buf ( n45369 , n45368 );
nand ( n45370 , n44834 , n44945 );
buf ( n45371 , n45370 );
not ( n45372 , n45371 );
buf ( n45373 , n45372 );
buf ( n45374 , n44683 );
buf ( n45375 , n44525 );
nand ( n45376 , n45374 , n45375 );
buf ( n45377 , n45376 );
buf ( n45378 , n44520 );
not ( n45379 , n45378 );
buf ( n45380 , n45379 );
or ( n45381 , n44298 , n44095 );
buf ( n45382 , n45381 );
nand ( n45383 , n44298 , n44095 );
buf ( n45384 , n45383 );
buf ( n45385 , n45384 );
nand ( n45386 , n45382 , n45385 );
buf ( n45387 , n45386 );
not ( n45388 , n43079 );
not ( n45389 , n43253 );
or ( n45390 , n45388 , n45389 );
not ( n45391 , n42925 );
not ( n45392 , n42807 );
buf ( n45393 , n42735 );
buf ( n45394 , n42740 );
xnor ( n45395 , n45393 , n45394 );
buf ( n45396 , n45395 );
buf ( n45397 , n45396 );
buf ( n45398 , n393 );
buf ( n45399 , n409 );
nand ( n45400 , n45398 , n45399 );
buf ( n45401 , n45400 );
buf ( n45402 , n45401 );
not ( n45403 , n45402 );
buf ( n45404 , n408 );
nand ( n45405 , n45403 , n45404 );
buf ( n45406 , n45405 );
buf ( n45407 , n45406 );
nand ( n45408 , n45397 , n45407 );
buf ( n45409 , n45408 );
buf ( n45410 , n45409 );
buf ( n45411 , n408 );
not ( n45412 , n45411 );
buf ( n45413 , n45401 );
nand ( n45414 , n45412 , n45413 );
buf ( n45415 , n45414 );
buf ( n45416 , n45415 );
buf ( n45417 , n417 );
and ( n45418 , n45410 , n45416 , n45417 );
buf ( n45419 , n45418 );
buf ( n45420 , n45419 );
not ( n45421 , n45420 );
buf ( n45422 , n42748 );
not ( n45423 , n45422 );
or ( n45424 , n45421 , n45423 );
buf ( n45425 , n42721 );
not ( n45426 , n45425 );
buf ( n45427 , n45426 );
buf ( n45428 , n45427 );
nand ( n45429 , n45424 , n45428 );
buf ( n45430 , n45429 );
buf ( n45431 , n42748 );
buf ( n45432 , n45419 );
or ( n45433 , n45431 , n45432 );
buf ( n45434 , n45433 );
and ( n45435 , n42796 , n45430 , n45434 );
not ( n45436 , n45435 );
and ( n45437 , n45392 , n45436 );
buf ( n45438 , n45430 );
buf ( n45439 , n45434 );
and ( n45440 , n45438 , n45439 );
buf ( n45441 , n42796 );
nor ( n45442 , n45440 , n45441 );
buf ( n45443 , n45442 );
nor ( n45444 , n45437 , n45443 );
nand ( n45445 , n45444 , n42891 );
nand ( n45446 , n45391 , n45445 );
or ( n45447 , n45444 , n42891 );
and ( n45448 , n45446 , n45447 , n42930 );
or ( n45449 , n45448 , n43074 );
not ( n45450 , n42930 );
nand ( n45451 , n45446 , n45447 );
nand ( n45452 , n45450 , n45451 );
nand ( n45453 , n45449 , n45452 );
nand ( n45454 , n45390 , n45453 );
buf ( n45455 , n45454 );
buf ( n45456 , n43253 );
buf ( n45457 , n43079 );
or ( n45458 , n45456 , n45457 );
buf ( n45459 , n45458 );
buf ( n45460 , n45459 );
buf ( n45461 , n43258 );
and ( n45462 , n45455 , n45460 );
nor ( n45463 , n45462 , n45461 );
buf ( n45464 , n45463 );
buf ( n45465 , n45275 );
buf ( n45466 , n45289 );
nand ( n45467 , n45465 , n45466 );
buf ( n45468 , n45467 );
buf ( n45469 , n45468 );
not ( n45470 , n45469 );
buf ( n45471 , n45470 );
buf ( n45472 , n45292 );
not ( n45473 , n45472 );
buf ( n45474 , n45473 );
buf ( n45475 , n45474 );
buf ( n45476 , n45351 );
nor ( n45477 , n45475 , n45476 );
buf ( n45478 , n45477 );
nand ( n45479 , n45341 , n45307 , n45310 );
buf ( n45480 , n45479 );
buf ( n45481 , n45338 );
not ( n45482 , n45480 );
nand ( n45483 , n45482 , n45481 );
buf ( n45484 , n45483 );
buf ( n45485 , n45293 );
buf ( n45486 , n45295 );
or ( n45487 , n45485 , n45486 );
buf ( n45488 , n45487 );
xnor ( n45489 , n413 , n412 );
buf ( n45490 , n411 );
buf ( n45491 , n412 );
xor ( n45492 , n45490 , n45491 );
buf ( n45493 , n45492 );
and ( n45494 , n45489 , n45493 );
buf ( n45495 , n45494 );
not ( n45496 , n45495 );
buf ( n45497 , n45496 );
nand ( n45498 , n45497 , n45489 );
not ( n45499 , n411 );
and ( n45500 , n421 , n425 );
buf ( n45501 , n422 );
buf ( n45502 , n423 );
or ( n45503 , n45501 , n45502 );
buf ( n45504 , n373 );
not ( n45505 , n45504 );
buf ( n45506 , n45505 );
buf ( n45507 , n45506 );
nand ( n45508 , n45503 , n45507 );
buf ( n45509 , n45508 );
nand ( n45510 , n422 , n423 );
nand ( n45511 , n45509 , n45510 );
xor ( n45512 , n45500 , n45511 );
buf ( n45513 , n372 );
not ( n45514 , n45513 );
buf ( n45515 , n421 );
not ( n45516 , n45515 );
and ( n45517 , n45514 , n45516 );
buf ( n45518 , n372 );
buf ( n45519 , n421 );
and ( n45520 , n45518 , n45519 );
nor ( n45521 , n45517 , n45520 );
buf ( n45522 , n45521 );
nand ( n45523 , n424 , n422 );
and ( n45524 , n45522 , n45523 );
not ( n45525 , n45522 );
not ( n45526 , n45523 );
and ( n45527 , n45525 , n45526 );
nor ( n45528 , n45524 , n45527 );
xor ( n45529 , n45512 , n45528 );
buf ( n45530 , n422 );
buf ( n45531 , n425 );
nand ( n45532 , n45530 , n45531 );
buf ( n45533 , n45532 );
buf ( n45534 , n45533 );
not ( n45535 , n45534 );
buf ( n45536 , n424 );
buf ( n45537 , n423 );
nand ( n45538 , n45536 , n45537 );
buf ( n45539 , n45538 );
buf ( n45540 , n45539 );
not ( n45541 , n45540 );
or ( n45542 , n45535 , n45541 );
buf ( n45543 , n424 );
buf ( n45544 , n423 );
nor ( n45545 , n45543 , n45544 );
buf ( n45546 , n45545 );
buf ( n45547 , n45546 );
buf ( n45548 , n374 );
or ( n45549 , n45547 , n45548 );
buf ( n45550 , n45539 );
nand ( n45551 , n45549 , n45550 );
buf ( n45552 , n45551 );
buf ( n45553 , n45552 );
nand ( n45554 , n45542 , n45553 );
buf ( n45555 , n45554 );
buf ( n45556 , n45555 );
not ( n45557 , n45556 );
buf ( n45558 , n45557 );
nor ( n45559 , n45529 , n45558 );
buf ( n45560 , n45559 );
buf ( n45561 , n424 );
buf ( n45562 , n423 );
and ( n45563 , n45561 , n45562 );
buf ( n45564 , n45563 );
buf ( n45565 , n45564 );
buf ( n45566 , n45533 );
and ( n45567 , n45565 , n45566 );
not ( n45568 , n45565 );
buf ( n45569 , n45533 );
not ( n45570 , n45569 );
buf ( n45571 , n45570 );
buf ( n45572 , n45571 );
and ( n45573 , n45568 , n45572 );
nor ( n45574 , n45567 , n45573 );
buf ( n45575 , n45574 );
xnor ( n45576 , n45575 , n45552 );
buf ( n45577 , n45576 );
xor ( n45578 , n423 , n373 );
xnor ( n45579 , n45578 , n422 );
buf ( n45580 , n45579 );
nor ( n45581 , n45577 , n45580 );
buf ( n45582 , n45581 );
buf ( n45583 , n45582 );
nor ( n45584 , n45560 , n45583 );
buf ( n45585 , n45584 );
buf ( n45586 , n45585 );
xor ( n45587 , n45500 , n45511 );
and ( n45588 , n45587 , n45528 );
and ( n45589 , n45500 , n45511 );
or ( n45590 , n45588 , n45589 );
not ( n45591 , n45590 );
not ( n45592 , n421 );
nand ( n45593 , n45592 , n372 );
not ( n45594 , n45593 );
and ( n45595 , n422 , n424 );
not ( n45596 , n45595 );
or ( n45597 , n45594 , n45596 );
not ( n45598 , n372 );
nand ( n45599 , n45598 , n421 );
nand ( n45600 , n45597 , n45599 );
not ( n45601 , n45600 );
xor ( n45602 , n371 , n420 );
and ( n45603 , n45602 , n422 );
not ( n45604 , n45602 );
not ( n45605 , n422 );
and ( n45606 , n45604 , n45605 );
nor ( n45607 , n45603 , n45606 );
not ( n45608 , n45607 );
not ( n45609 , n45608 );
or ( n45610 , n45601 , n45609 );
or ( n45611 , n45600 , n45608 );
nand ( n45612 , n45610 , n45611 );
not ( n45613 , n45612 );
and ( n45614 , n422 , n423 );
buf ( n45615 , n420 );
buf ( n45616 , n425 );
and ( n45617 , n45615 , n45616 );
buf ( n45618 , n45617 );
nand ( n45619 , n424 , n421 );
and ( n45620 , n45618 , n45619 );
not ( n45621 , n45618 );
not ( n45622 , n45619 );
and ( n45623 , n45621 , n45622 );
or ( n45624 , n45620 , n45623 );
xor ( n45625 , n45614 , n45624 );
not ( n45626 , n45625 );
or ( n45627 , n45613 , n45626 );
or ( n45628 , n45612 , n45625 );
nand ( n45629 , n45627 , n45628 );
not ( n45630 , n45629 );
nand ( n45631 , n45591 , n45630 );
buf ( n45632 , n45631 );
not ( n45633 , n425 );
nand ( n45634 , n45633 , n419 );
and ( n45635 , n45634 , n370 );
not ( n45636 , n45634 );
not ( n45637 , n370 );
and ( n45638 , n45636 , n45637 );
nor ( n45639 , n45635 , n45638 );
buf ( n45640 , n45639 );
not ( n45641 , n45614 );
not ( n45642 , n45622 );
or ( n45643 , n45641 , n45642 );
not ( n45644 , n45510 );
not ( n45645 , n45619 );
or ( n45646 , n45644 , n45645 );
nand ( n45647 , n45646 , n45618 );
nand ( n45648 , n45643 , n45647 );
buf ( n45649 , n45648 );
xor ( n45650 , n45640 , n45649 );
buf ( n45651 , n424 );
buf ( n45652 , n420 );
nand ( n45653 , n45651 , n45652 );
buf ( n45654 , n45653 );
buf ( n45655 , n45654 );
not ( n45656 , n45655 );
buf ( n45657 , n45656 );
buf ( n45658 , n45657 );
buf ( n45659 , n421 );
buf ( n45660 , n423 );
and ( n45661 , n45659 , n45660 );
buf ( n45662 , n45661 );
buf ( n45663 , n45662 );
xor ( n45664 , n45658 , n45663 );
buf ( n45665 , n420 );
buf ( n45666 , n422 );
nor ( n45667 , n45665 , n45666 );
buf ( n45668 , n45667 );
buf ( n45669 , n45668 );
buf ( n45670 , n371 );
or ( n45671 , n45669 , n45670 );
buf ( n45672 , n420 );
buf ( n45673 , n422 );
nand ( n45674 , n45672 , n45673 );
buf ( n45675 , n45674 );
buf ( n45676 , n45675 );
nand ( n45677 , n45671 , n45676 );
buf ( n45678 , n45677 );
buf ( n45679 , n45678 );
xor ( n45680 , n45664 , n45679 );
buf ( n45681 , n45680 );
buf ( n45682 , n45681 );
xor ( n45683 , n45650 , n45682 );
buf ( n45684 , n45683 );
buf ( n45685 , n45684 );
not ( n45686 , n45685 );
buf ( n45687 , n45600 );
not ( n45688 , n45687 );
buf ( n45689 , n45607 );
buf ( n45690 , n45689 );
nand ( n45691 , n45688 , n45690 );
buf ( n45692 , n45691 );
and ( n45693 , n45625 , n45692 );
not ( n45694 , n45600 );
nor ( n45695 , n45694 , n45689 );
nor ( n45696 , n45693 , n45695 );
buf ( n45697 , n45696 );
nand ( n45698 , n45686 , n45697 );
buf ( n45699 , n45698 );
buf ( n45700 , n45699 );
xor ( n45701 , n424 , n374 );
not ( n45702 , n423 );
xor ( n45703 , n45701 , n45702 );
buf ( n45704 , n45703 );
buf ( n45705 , n423 );
buf ( n45706 , n425 );
and ( n45707 , n45705 , n45706 );
buf ( n45708 , n45707 );
buf ( n45709 , n45708 );
or ( n45710 , n45704 , n45709 );
not ( n45711 , n376 );
not ( n45712 , n377 );
and ( n45713 , n45711 , n45712 );
nor ( n45714 , n45713 , n425 );
buf ( n45715 , n45714 );
and ( n45716 , n424 , n425 );
nor ( n45717 , n45716 , n40363 );
buf ( n45718 , n45717 );
nor ( n45719 , n45715 , n45718 );
buf ( n45720 , n45719 );
buf ( n45721 , n45720 );
nand ( n45722 , n45710 , n45721 );
buf ( n45723 , n45722 );
buf ( n45724 , n45703 );
buf ( n45725 , n45708 );
nand ( n45726 , n45724 , n45725 );
buf ( n45727 , n45726 );
nand ( n45728 , n45723 , n45727 );
buf ( n45729 , n45728 );
nand ( n45730 , n45586 , n45632 , n45700 , n45729 );
buf ( n45731 , n45730 );
buf ( n45732 , n45629 );
buf ( n45733 , n45590 );
nor ( n45734 , n45732 , n45733 );
buf ( n45735 , n45734 );
buf ( n45736 , n45735 );
buf ( n45737 , n45559 );
nor ( n45738 , n45736 , n45737 );
buf ( n45739 , n45738 );
buf ( n45740 , n45739 );
buf ( n45741 , n45699 );
nand ( n45742 , n45529 , n45558 );
buf ( n45743 , n45742 );
nand ( n45744 , n45576 , n45579 );
buf ( n45745 , n45744 );
nand ( n45746 , n45743 , n45745 );
buf ( n45747 , n45746 );
buf ( n45748 , n45747 );
nand ( n45749 , n45740 , n45741 , n45748 );
buf ( n45750 , n45749 );
buf ( n45751 , n45684 );
not ( n45752 , n45751 );
buf ( n45753 , n45696 );
nand ( n45754 , n45752 , n45753 );
buf ( n45755 , n45754 );
buf ( n45756 , n45755 );
buf ( n45757 , n45629 );
buf ( n45758 , n45590 );
and ( n45759 , n45757 , n45758 );
buf ( n45760 , n45759 );
buf ( n45761 , n45760 );
nand ( n45762 , n45756 , n45761 );
buf ( n45763 , n45762 );
buf ( n45764 , n45696 );
not ( n45765 , n45764 );
buf ( n45766 , n45684 );
buf ( n45767 , n45766 );
buf ( n45768 , n45767 );
buf ( n45769 , n45768 );
nand ( n45770 , n45765 , n45769 );
buf ( n45771 , n45770 );
nand ( n45772 , n45731 , n45750 , n45763 , n45771 );
buf ( n45773 , n45772 );
buf ( n45774 , n419 );
not ( n45775 , n45774 );
buf ( n45776 , n418 );
buf ( n45777 , n420 );
nand ( n45778 , n45776 , n45777 );
buf ( n45779 , n45778 );
buf ( n45780 , n45779 );
nand ( n45781 , n45775 , n45780 );
buf ( n45782 , n45781 );
buf ( n45783 , n419 );
not ( n45784 , n45783 );
buf ( n45785 , n418 );
nand ( n45786 , n45784 , n45785 );
buf ( n45787 , n45786 );
or ( n45788 , n45782 , n45787 );
not ( n45789 , n45788 );
buf ( n45790 , n418 );
buf ( n45791 , n422 );
nand ( n45792 , n45790 , n45791 );
buf ( n45793 , n45792 );
buf ( n45794 , n419 );
buf ( n45795 , n421 );
nand ( n45796 , n45794 , n45795 );
buf ( n45797 , n45796 );
nand ( n45798 , n45793 , n45797 );
buf ( n45799 , n45798 );
not ( n45800 , n45799 );
buf ( n45801 , n419 );
not ( n45802 , n45801 );
buf ( n45803 , n420 );
nor ( n45804 , n45802 , n45803 );
buf ( n45805 , n45804 );
buf ( n45806 , n45805 );
not ( n45807 , n45806 );
buf ( n45808 , n45807 );
buf ( n45809 , n45808 );
not ( n45810 , n45809 );
or ( n45811 , n45800 , n45810 );
buf ( n45812 , n418 );
buf ( n45813 , n421 );
nand ( n45814 , n45812 , n45813 );
buf ( n45815 , n45814 );
buf ( n45816 , n45815 );
nand ( n45817 , n45811 , n45816 );
buf ( n45818 , n45817 );
buf ( n45819 , n45818 );
buf ( n45820 , n419 );
not ( n45821 , n45820 );
buf ( n45822 , n45779 );
nor ( n45823 , n45821 , n45822 );
buf ( n45824 , n45823 );
buf ( n45825 , n45824 );
not ( n45826 , n45825 );
buf ( n45827 , n45782 );
nand ( n45828 , n45826 , n45827 );
buf ( n45829 , n45828 );
buf ( n45830 , n45829 );
nor ( n45831 , n45819 , n45830 );
buf ( n45832 , n45831 );
not ( n45833 , n45832 );
not ( n45834 , n420 );
buf ( n45835 , n418 );
buf ( n45836 , n423 );
nand ( n45837 , n45835 , n45836 );
buf ( n45838 , n45837 );
nand ( n45839 , n45834 , n45838 );
not ( n45840 , n45797 );
not ( n45841 , n45793 );
or ( n45842 , n45840 , n45841 );
buf ( n45843 , n419 );
buf ( n45844 , n422 );
nand ( n45845 , n45843 , n45844 );
buf ( n45846 , n45845 );
not ( n45847 , n45846 );
not ( n45848 , n45815 );
nand ( n45849 , n45847 , n45848 );
nand ( n45850 , n45842 , n45849 );
xor ( n45851 , n45839 , n45850 );
buf ( n45852 , n420 );
buf ( n45853 , n421 );
nand ( n45854 , n45852 , n45853 );
buf ( n45855 , n45854 );
buf ( n45856 , n45855 );
buf ( n45857 , n45846 );
nand ( n45858 , n45856 , n45857 );
buf ( n45859 , n45858 );
buf ( n45860 , n45675 );
buf ( n45861 , n419 );
buf ( n45862 , n423 );
nand ( n45863 , n45861 , n45862 );
buf ( n45864 , n45863 );
buf ( n45865 , n45864 );
nand ( n45866 , n45860 , n45865 );
buf ( n45867 , n45866 );
and ( n45868 , n45859 , n45867 );
and ( n45869 , n45851 , n45868 );
and ( n45870 , n45839 , n45850 );
or ( n45871 , n45869 , n45870 );
xor ( n45872 , n45848 , n45805 );
xnor ( n45873 , n45872 , n45798 );
or ( n45874 , n45871 , n45873 );
nand ( n45875 , n45833 , n45874 );
nor ( n45876 , n45789 , n45875 );
xor ( n45877 , n45658 , n45663 );
and ( n45878 , n45877 , n45679 );
and ( n45879 , n45658 , n45663 );
or ( n45880 , n45878 , n45879 );
buf ( n45881 , n45880 );
buf ( n45882 , n45881 );
nand ( n45883 , n421 , n422 );
nand ( n45884 , n420 , n423 );
xor ( n45885 , n45883 , n45884 );
nand ( n45886 , n424 , n419 );
xnor ( n45887 , n45885 , n45886 );
buf ( n45888 , n45887 );
xor ( n45889 , n45882 , n45888 );
buf ( n45890 , n425 );
buf ( n45891 , n418 );
nand ( n45892 , n45890 , n45891 );
buf ( n45893 , n45892 );
buf ( n45894 , n45893 );
not ( n45895 , n45894 );
buf ( n45896 , n45895 );
buf ( n45897 , n45896 );
buf ( n45898 , n418 );
buf ( n45899 , n421 );
xnor ( n45900 , n45898 , n45899 );
buf ( n45901 , n45900 );
buf ( n45902 , n45901 );
xor ( n45903 , n45897 , n45902 );
not ( n45904 , n419 );
not ( n45905 , n45637 );
or ( n45906 , n45904 , n45905 );
nand ( n45907 , n419 , n425 );
nand ( n45908 , n45906 , n45907 );
buf ( n45909 , n45908 );
xor ( n45910 , n45903 , n45909 );
buf ( n45911 , n45910 );
buf ( n45912 , n45911 );
and ( n45913 , n45889 , n45912 );
and ( n45914 , n45882 , n45888 );
or ( n45915 , n45913 , n45914 );
buf ( n45916 , n45915 );
buf ( n45917 , n45916 );
not ( n45918 , n45917 );
or ( n45919 , n45864 , n45675 );
nand ( n45920 , n45919 , n45867 );
xor ( n45921 , n45897 , n45902 );
and ( n45922 , n45921 , n45909 );
and ( n45923 , n45897 , n45902 );
or ( n45924 , n45922 , n45923 );
buf ( n45925 , n45924 );
xor ( n45926 , n45920 , n45925 );
and ( n45927 , n424 , n419 );
not ( n45928 , n45927 );
not ( n45929 , n420 );
not ( n45930 , n423 );
or ( n45931 , n45929 , n45930 );
nand ( n45932 , n421 , n422 );
nand ( n45933 , n45931 , n45932 );
not ( n45934 , n45933 );
or ( n45935 , n45928 , n45934 );
nand ( n45936 , n421 , n422 , n420 , n423 );
nand ( n45937 , n45935 , n45936 );
buf ( n45938 , n418 );
not ( n45939 , n45938 );
buf ( n45940 , n421 );
not ( n45941 , n45940 );
and ( n45942 , n45939 , n45941 );
buf ( n45943 , n424 );
buf ( n45944 , n418 );
and ( n45945 , n45943 , n45944 );
nor ( n45946 , n45942 , n45945 );
buf ( n45947 , n45946 );
and ( n45948 , n45937 , n45947 );
not ( n45949 , n45937 );
not ( n45950 , n45947 );
and ( n45951 , n45949 , n45950 );
nor ( n45952 , n45948 , n45951 );
xor ( n45953 , n45926 , n45952 );
buf ( n45954 , n45953 );
not ( n45955 , n45954 );
and ( n45956 , n45918 , n45955 );
xor ( n45957 , n45640 , n45649 );
and ( n45958 , n45957 , n45682 );
and ( n45959 , n45640 , n45649 );
or ( n45960 , n45958 , n45959 );
buf ( n45961 , n45960 );
xor ( n45962 , n45882 , n45888 );
xor ( n45963 , n45962 , n45912 );
buf ( n45964 , n45963 );
nor ( n45965 , n45961 , n45964 );
buf ( n45966 , n45965 );
nor ( n45967 , n45956 , n45966 );
buf ( n45968 , n45967 );
buf ( n45969 , n45968 );
buf ( n45970 , n423 );
not ( n45971 , n45970 );
buf ( n45972 , n45779 );
not ( n45973 , n45972 );
buf ( n45974 , n45973 );
buf ( n45975 , n45974 );
not ( n45976 , n45975 );
or ( n45977 , n45971 , n45976 );
buf ( n45978 , n45839 );
nand ( n45979 , n45977 , n45978 );
buf ( n45980 , n45979 );
buf ( n45981 , n45980 );
not ( n45982 , n45855 );
not ( n45983 , n45847 );
or ( n45984 , n45982 , n45983 );
nand ( n45985 , n419 , n422 );
nand ( n45986 , n45985 , n420 , n421 );
nand ( n45987 , n45984 , n45986 );
xor ( n45988 , n45987 , n45867 );
buf ( n45989 , n45988 );
xor ( n45990 , n45981 , n45989 );
buf ( n45991 , n421 );
not ( n45992 , n45991 );
buf ( n45993 , n45937 );
not ( n45994 , n45993 );
or ( n45995 , n45992 , n45994 );
buf ( n45996 , n424 );
buf ( n45997 , n418 );
nand ( n45998 , n45996 , n45997 );
buf ( n45999 , n45998 );
buf ( n46000 , n45999 );
nand ( n46001 , n45995 , n46000 );
buf ( n46002 , n46001 );
buf ( n46003 , n46002 );
xor ( n46004 , n45990 , n46003 );
buf ( n46005 , n46004 );
buf ( n46006 , n45952 );
not ( n46007 , n46006 );
buf ( n46008 , n46007 );
not ( n46009 , n46008 );
buf ( n46010 , n45920 );
not ( n46011 , n46010 );
buf ( n46012 , n46011 );
not ( n46013 , n46012 );
and ( n46014 , n46009 , n46013 );
buf ( n46015 , n46008 );
buf ( n46016 , n46012 );
nand ( n46017 , n46015 , n46016 );
buf ( n46018 , n46017 );
buf ( n46019 , n45925 );
buf ( n46020 , n46019 );
buf ( n46021 , n46020 );
and ( n46022 , n46018 , n46021 );
nor ( n46023 , n46014 , n46022 );
buf ( n46024 , n46023 );
not ( n46025 , n46024 );
buf ( n46026 , n46025 );
nor ( n46027 , n46005 , n46026 );
xor ( n46028 , n45981 , n45989 );
and ( n46029 , n46028 , n46003 );
and ( n46030 , n45981 , n45989 );
or ( n46031 , n46029 , n46030 );
buf ( n46032 , n46031 );
xor ( n46033 , n45839 , n45850 );
xor ( n46034 , n46033 , n45868 );
nor ( n46035 , n46032 , n46034 );
nor ( n46036 , n46027 , n46035 );
buf ( n46037 , n46036 );
nand ( n46038 , n45773 , n45876 , n45969 , n46037 );
buf ( n46039 , n46038 );
not ( n46040 , n46036 );
or ( n46041 , n45916 , n45953 );
nand ( n46042 , n45964 , n45961 );
not ( n46043 , n46042 );
nand ( n46044 , n46041 , n46043 );
nand ( n46045 , n45916 , n45953 );
nand ( n46046 , n46044 , n46045 );
not ( n46047 , n46046 );
or ( n46048 , n46040 , n46047 );
nand ( n46049 , n46032 , n46034 );
not ( n46050 , n46049 );
nand ( n46051 , n46005 , n46026 );
nor ( n46052 , n46035 , n46051 );
nor ( n46053 , n46050 , n46052 );
nand ( n46054 , n46048 , n46053 );
nand ( n46055 , n46054 , n45876 );
buf ( n46056 , n46055 );
buf ( n46057 , n45871 );
buf ( n46058 , n45873 );
nand ( n46059 , n46057 , n46058 );
buf ( n46060 , n46059 );
buf ( n46061 , n46060 );
buf ( n46062 , n45832 );
or ( n46063 , n46061 , n46062 );
buf ( n46064 , n45818 );
buf ( n46065 , n45829 );
nand ( n46066 , n46064 , n46065 );
buf ( n46067 , n46066 );
buf ( n46068 , n46067 );
nand ( n46069 , n46063 , n46068 );
buf ( n46070 , n46069 );
and ( n46071 , n46070 , n45788 );
buf ( n46072 , n46071 );
buf ( n46073 , n418 );
not ( n46074 , n46073 );
buf ( n46075 , n45782 );
buf ( n46076 , n45787 );
nand ( n46077 , n46075 , n46076 );
buf ( n46078 , n46077 );
buf ( n46079 , n46078 );
nand ( n46080 , n46074 , n46079 );
buf ( n46081 , n46080 );
buf ( n46082 , n46081 );
nor ( n46083 , n46072 , n46082 );
buf ( n46084 , n46083 );
buf ( n46085 , n46084 );
nand ( n46086 , n46039 , n46056 , n46085 );
buf ( n46087 , n46086 );
buf ( n46088 , n46087 );
not ( n46089 , n46088 );
buf ( n46090 , n46089 );
buf ( n46091 , n46090 );
not ( n46092 , n46091 );
buf ( n46093 , n46092 );
not ( n46094 , n46093 );
or ( n46095 , n45499 , n46094 );
buf ( n46096 , n411 );
not ( n46097 , n46096 );
buf ( n46098 , n46090 );
nand ( n46099 , n46097 , n46098 );
buf ( n46100 , n46099 );
nand ( n46101 , n46095 , n46100 );
nand ( n46102 , n45498 , n46101 );
not ( n46103 , n46102 );
buf ( n46104 , n46090 );
not ( n46105 , n46104 );
buf ( n46106 , n416 );
not ( n46107 , n46106 );
buf ( n46108 , n46107 );
buf ( n46109 , n46108 );
buf ( n46110 , n415 );
and ( n46111 , n46109 , n46110 );
buf ( n46112 , n46111 );
buf ( n46113 , n46112 );
nand ( n46114 , n46105 , n46113 );
buf ( n46115 , n46114 );
buf ( n46116 , n415 );
not ( n46117 , n46116 );
buf ( n46118 , n46087 );
not ( n46119 , n46118 );
or ( n46120 , n46117 , n46119 );
buf ( n46121 , n46090 );
buf ( n46122 , n415 );
not ( n46123 , n46122 );
buf ( n46124 , n46123 );
buf ( n46125 , n46124 );
nand ( n46126 , n46121 , n46125 );
buf ( n46127 , n46126 );
buf ( n46128 , n46127 );
nand ( n46129 , n46120 , n46128 );
buf ( n46130 , n46129 );
buf ( n46131 , n46130 );
buf ( n46132 , n416 );
nand ( n46133 , n46131 , n46132 );
buf ( n46134 , n46133 );
nand ( n46135 , n46115 , n46134 );
not ( n46136 , n46135 );
or ( n46137 , n46103 , n46136 );
buf ( n46138 , n46134 );
buf ( n46139 , n46115 );
nand ( n46140 , n46138 , n46139 );
buf ( n46141 , n46140 );
buf ( n46142 , n46141 );
not ( n46143 , n46142 );
and ( n46144 , n46101 , n45498 );
buf ( n46145 , n46144 );
nand ( n46146 , n46143 , n46145 );
buf ( n46147 , n46146 );
nand ( n46148 , n46137 , n46147 );
not ( n46149 , n413 );
not ( n46150 , n46093 );
or ( n46151 , n46149 , n46150 );
buf ( n46152 , n46090 );
not ( n46153 , n413 );
buf ( n46154 , n46153 );
nand ( n46155 , n46152 , n46154 );
buf ( n46156 , n46155 );
nand ( n46157 , n46151 , n46156 );
buf ( n46158 , n46153 );
buf ( n46159 , n414 );
not ( n46160 , n46159 );
buf ( n46161 , n46160 );
buf ( n46162 , n46161 );
and ( n46163 , n46158 , n46162 );
buf ( n46164 , n413 );
buf ( n46165 , n414 );
and ( n46166 , n46164 , n46165 );
nor ( n46167 , n46163 , n46166 );
buf ( n46168 , n46167 );
not ( n46169 , n415 );
not ( n46170 , n414 );
or ( n46171 , n46169 , n46170 );
buf ( n46172 , n46124 );
buf ( n46173 , n46161 );
nand ( n46174 , n46172 , n46173 );
buf ( n46175 , n46174 );
nand ( n46176 , n46171 , n46175 );
and ( n46177 , n46168 , n46176 );
buf ( n46178 , n46177 );
not ( n46179 , n46178 );
buf ( n46180 , n46179 );
nand ( n46181 , n46180 , n46176 );
nand ( n46182 , n46157 , n46181 );
buf ( n46183 , n46182 );
buf ( n46184 , n46090 );
xor ( n46185 , n410 , n411 );
buf ( n46186 , n46185 );
nand ( n46187 , n46184 , n46186 );
buf ( n46188 , n46187 );
not ( n46189 , n46188 );
buf ( n46190 , n46185 );
not ( n46191 , n46190 );
buf ( n46192 , n46191 );
buf ( n46193 , n46192 );
buf ( n46194 , n410 );
and ( n46195 , n46193 , n46194 );
buf ( n46196 , n46195 );
and ( n46197 , n46196 , n46090 );
nor ( n46198 , n46189 , n46197 );
buf ( n46199 , n46198 );
nand ( n46200 , n46183 , n46199 );
and ( n46201 , n46148 , n46200 );
not ( n46202 , n46148 );
not ( n46203 , n46200 );
and ( n46204 , n46202 , n46203 );
nor ( n46205 , n46201 , n46204 );
not ( n46206 , n46205 );
not ( n46207 , n46182 );
not ( n46208 , n46198 );
nor ( n46209 , n46207 , n46208 );
not ( n46210 , n46209 );
not ( n46211 , n46176 );
not ( n46212 , n46180 );
or ( n46213 , n46211 , n46212 );
nand ( n46214 , n46213 , n46157 );
buf ( n46215 , n46214 );
not ( n46216 , n46215 );
buf ( n46217 , n46216 );
buf ( n46218 , n46217 );
buf ( n46219 , n46208 );
nand ( n46220 , n46218 , n46219 );
buf ( n46221 , n46220 );
nand ( n46222 , n46210 , n46221 );
not ( n46223 , n46222 );
nand ( n46224 , n46206 , n46223 );
not ( n46225 , n46224 );
buf ( n46226 , n46102 );
buf ( n46227 , n46209 );
nand ( n46228 , n46226 , n46227 );
buf ( n46229 , n46228 );
not ( n46230 , n46229 );
buf ( n46231 , n46135 );
not ( n46232 , n46231 );
or ( n46233 , n46230 , n46232 );
not ( n46234 , n46209 );
buf ( n46235 , n46234 );
buf ( n46236 , n46144 );
buf ( n46237 , n46236 );
buf ( n46238 , n46237 );
buf ( n46239 , n46238 );
nand ( n46240 , n46235 , n46239 );
buf ( n46241 , n46240 );
nand ( n46242 , n46233 , n46241 );
not ( n46243 , n46242 );
or ( n46244 , n46225 , n46243 );
nand ( n46245 , n46205 , n46222 );
nand ( n46246 , n46244 , n46245 );
buf ( n46247 , n46246 );
not ( n46248 , n46247 );
buf ( n46249 , n46248 );
buf ( n46250 , n46242 );
not ( n46251 , n46250 );
not ( n46252 , n46206 );
not ( n46253 , n46222 );
or ( n46254 , n46252 , n46253 );
nand ( n46255 , n46205 , n46223 );
nand ( n46256 , n46254 , n46255 );
not ( n46257 , n46256 );
buf ( n46258 , n46257 );
not ( n46259 , n46258 );
or ( n46260 , n46251 , n46259 );
buf ( n46261 , n46256 );
buf ( n46262 , n46242 );
not ( n46263 , n46262 );
buf ( n46264 , n46263 );
buf ( n46265 , n46264 );
nand ( n46266 , n46261 , n46265 );
buf ( n46267 , n46266 );
buf ( n46268 , n46267 );
nand ( n46269 , n46260 , n46268 );
buf ( n46270 , n46269 );
buf ( n46271 , n376 );
buf ( n46272 , n382 );
nand ( n46273 , n46271 , n46272 );
buf ( n46274 , n46273 );
nand ( n46275 , n374 , n380 );
or ( n46276 , n46274 , n46275 );
nand ( n46277 , n377 , n379 );
not ( n46278 , n46277 );
nand ( n46279 , n375 , n381 );
not ( n46280 , n46279 );
or ( n46281 , n46278 , n46280 );
or ( n46282 , n46277 , n46279 );
nand ( n46283 , n372 , n384 );
nand ( n46284 , n46282 , n46283 );
nand ( n46285 , n46281 , n46284 );
xor ( n46286 , n46276 , n46285 );
buf ( n46287 , n374 );
buf ( n46288 , n381 );
nand ( n46289 , n46287 , n46288 );
buf ( n46290 , n46289 );
buf ( n46291 , n373 );
buf ( n46292 , n382 );
nand ( n46293 , n46291 , n46292 );
buf ( n46294 , n46293 );
buf ( n46295 , n370 );
buf ( n46296 , n385 );
nand ( n46297 , n46295 , n46296 );
buf ( n46298 , n46297 );
nand ( n46299 , n46290 , n46294 , n46298 );
not ( n46300 , n46290 );
not ( n46301 , n46298 );
nand ( n46302 , n46300 , n46294 , n46301 );
not ( n46303 , n46294 );
nand ( n46304 , n46303 , n46298 , n46300 );
nand ( n46305 , n46301 , n46303 , n46290 );
nand ( n46306 , n46299 , n46302 , n46304 , n46305 );
xor ( n46307 , n46286 , n46306 );
buf ( n46308 , n46276 );
buf ( n46309 , n376 );
buf ( n46310 , n380 );
nand ( n46311 , n46309 , n46310 );
buf ( n46312 , n46311 );
buf ( n46313 , n46312 );
buf ( n46314 , n374 );
buf ( n46315 , n382 );
nand ( n46316 , n46314 , n46315 );
buf ( n46317 , n46316 );
buf ( n46318 , n46317 );
nand ( n46319 , n46313 , n46318 );
buf ( n46320 , n46319 );
buf ( n46321 , n46320 );
nand ( n46322 , n46308 , n46321 );
buf ( n46323 , n46322 );
not ( n46324 , n46323 );
nand ( n46325 , n375 , n381 );
xor ( n46326 , n46325 , n46277 );
xor ( n46327 , n46326 , n46283 );
buf ( n46328 , n372 );
buf ( n46329 , n385 );
nand ( n46330 , n46328 , n46329 );
buf ( n46331 , n46330 );
not ( n46332 , n46331 );
buf ( n46333 , n376 );
buf ( n46334 , n381 );
nand ( n46335 , n46333 , n46334 );
buf ( n46336 , n46335 );
not ( n46337 , n46336 );
or ( n46338 , n46332 , n46337 );
not ( n46339 , n46331 );
not ( n46340 , n46339 );
not ( n46341 , n46336 );
not ( n46342 , n46341 );
or ( n46343 , n46340 , n46342 );
nand ( n46344 , n374 , n383 );
nand ( n46345 , n46343 , n46344 );
nand ( n46346 , n46338 , n46345 );
or ( n46347 , n46327 , n46346 );
not ( n46348 , n46347 );
or ( n46349 , n46324 , n46348 );
nand ( n46350 , n46327 , n46346 );
nand ( n46351 , n46349 , n46350 );
xor ( n46352 , n46307 , n46351 );
buf ( n46353 , n372 );
buf ( n46354 , n383 );
nand ( n46355 , n46353 , n46354 );
buf ( n46356 , n46355 );
not ( n46357 , n46356 );
buf ( n46358 , n371 );
buf ( n46359 , n384 );
nand ( n46360 , n46358 , n46359 );
buf ( n46361 , n46360 );
not ( n46362 , n46361 );
or ( n46363 , n46357 , n46362 );
nand ( n46364 , n371 , n383 );
not ( n46365 , n46364 );
nand ( n46366 , n46365 , n372 , n384 );
nand ( n46367 , n46363 , n46366 );
nand ( n46368 , n376 , n379 );
nand ( n556 , n377 , n378 );
xor ( n557 , n46368 , n556 );
buf ( n46371 , n375 );
buf ( n46372 , n380 );
nand ( n46373 , n46371 , n46372 );
buf ( n46374 , n46373 );
not ( n562 , n46374 );
and ( n46376 , n557 , n562 );
not ( n564 , n557 );
and ( n565 , n564 , n46374 );
or ( n566 , n46376 , n565 );
xor ( n567 , n46367 , n566 );
nand ( n568 , n377 , n380 );
buf ( n46382 , n568 );
buf ( n46383 , n373 );
buf ( n46384 , n383 );
nand ( n572 , n46383 , n46384 );
buf ( n46386 , n572 );
buf ( n46387 , n46386 );
or ( n575 , n46382 , n46387 );
buf ( n46389 , n371 );
buf ( n46390 , n385 );
nand ( n578 , n46389 , n46390 );
buf ( n46392 , n578 );
buf ( n46393 , n46392 );
nand ( n581 , n575 , n46393 );
buf ( n46395 , n581 );
buf ( n46396 , n568 );
buf ( n46397 , n46386 );
nand ( n46398 , n46396 , n46397 );
buf ( n46399 , n46398 );
nand ( n587 , n46395 , n46399 );
xor ( n46401 , n567 , n587 );
and ( n589 , n46352 , n46401 );
and ( n590 , n46307 , n46351 );
or ( n591 , n589 , n590 );
buf ( n46405 , n591 );
xor ( n593 , n46367 , n566 );
and ( n594 , n593 , n587 );
and ( n595 , n46367 , n566 );
or ( n596 , n594 , n595 );
nand ( n46410 , n46290 , n46294 );
not ( n598 , n46300 );
not ( n599 , n46303 );
or ( n46413 , n598 , n599 );
nand ( n601 , n46413 , n46298 );
nand ( n602 , n46410 , n601 );
nand ( n603 , n371 , n383 );
xor ( n604 , n603 , n46275 );
nand ( n605 , n376 , n378 );
xor ( n606 , n604 , n605 );
not ( n607 , n606 );
not ( n608 , n46366 );
nand ( n609 , n607 , n608 );
nand ( n610 , n606 , n46366 );
nand ( n611 , n609 , n610 );
and ( n612 , n602 , n611 );
not ( n613 , n602 );
and ( n614 , n606 , n46366 );
not ( n615 , n606 );
and ( n616 , n615 , n608 );
nor ( n617 , n614 , n616 );
and ( n618 , n613 , n617 );
or ( n619 , n612 , n618 );
xor ( n620 , n596 , n619 );
buf ( n46434 , n372 );
buf ( n46435 , n382 );
nand ( n623 , n46434 , n46435 );
buf ( n46437 , n623 );
buf ( n46438 , n46437 );
not ( n626 , n46438 );
buf ( n46440 , n626 );
buf ( n46441 , n370 );
buf ( n46442 , n384 );
nand ( n630 , n46441 , n46442 );
buf ( n46444 , n630 );
xor ( n632 , n46440 , n46444 );
nand ( n633 , n376 , n379 );
not ( n634 , n633 );
not ( n635 , n634 );
not ( n636 , n562 );
or ( n637 , n635 , n636 );
nand ( n638 , n637 , n556 );
nand ( n639 , n46374 , n633 );
nand ( n640 , n638 , n639 );
xnor ( n641 , n632 , n640 );
buf ( n46455 , n373 );
buf ( n46456 , n381 );
nand ( n644 , n46455 , n46456 );
buf ( n46458 , n644 );
buf ( n46459 , n46458 );
not ( n647 , n46459 );
buf ( n46461 , n375 );
buf ( n46462 , n379 );
nand ( n650 , n46461 , n46462 );
buf ( n46464 , n650 );
buf ( n46465 , n46464 );
not ( n653 , n46465 );
or ( n654 , n647 , n653 );
nand ( n655 , n373 , n379 );
not ( n656 , n655 );
nand ( n657 , n656 , n375 , n381 );
buf ( n46471 , n657 );
nand ( n659 , n654 , n46471 );
buf ( n46473 , n659 );
buf ( n46474 , n46473 );
not ( n662 , n46474 );
buf ( n46476 , n662 );
xor ( n664 , n641 , n46476 );
xor ( n665 , n46276 , n46285 );
and ( n666 , n665 , n46306 );
and ( n667 , n46276 , n46285 );
or ( n668 , n666 , n667 );
not ( n669 , n668 );
xor ( n670 , n664 , n669 );
xor ( n671 , n620 , n670 );
buf ( n46485 , n671 );
xor ( n673 , n46405 , n46485 );
not ( n674 , n46185 );
nand ( n675 , n45630 , n45591 );
not ( n676 , n45744 );
not ( n677 , n45529 );
nand ( n678 , n677 , n45555 );
nand ( n679 , n676 , n678 );
nand ( n680 , n679 , n45742 );
nand ( n46494 , n675 , n680 );
buf ( n46495 , n675 );
buf ( n46496 , n45585 );
buf ( n46497 , n45728 );
nand ( n46498 , n46495 , n46496 , n46497 );
buf ( n46499 , n46498 );
buf ( n46500 , n45760 );
not ( n46501 , n46500 );
buf ( n46502 , n46501 );
nand ( n690 , n46494 , n46499 , n46502 );
nand ( n691 , n45755 , n45771 );
and ( n692 , n690 , n691 );
not ( n693 , n690 );
not ( n694 , n691 );
and ( n695 , n693 , n694 );
nor ( n696 , n692 , n695 );
buf ( n46510 , n696 );
not ( n698 , n46510 );
buf ( n46512 , n698 );
not ( n700 , n46512 );
or ( n701 , n674 , n700 );
buf ( n46515 , n675 );
buf ( n46516 , n46502 );
and ( n704 , n46515 , n46516 );
buf ( n46518 , n704 );
not ( n706 , n680 );
buf ( n46520 , n45585 );
buf ( n46521 , n45728 );
nand ( n709 , n46520 , n46521 );
buf ( n46523 , n709 );
nand ( n46524 , n706 , n46523 );
xor ( n712 , n46518 , n46524 );
buf ( n46526 , n712 );
buf ( n46527 , n46196 );
nand ( n715 , n46526 , n46527 );
buf ( n46529 , n715 );
nand ( n717 , n701 , n46529 );
buf ( n46531 , n717 );
xor ( n719 , n673 , n46531 );
buf ( n46533 , n719 );
buf ( n46534 , n46533 );
xor ( n722 , n46307 , n46351 );
xor ( n723 , n722 , n46401 );
buf ( n46537 , n723 );
not ( n725 , n46537 );
xor ( n726 , n46386 , n46392 );
not ( n727 , n568 );
xor ( n728 , n726 , n727 );
not ( n729 , n728 );
buf ( n46543 , n375 );
buf ( n46544 , n382 );
nand ( n732 , n46543 , n46544 );
buf ( n46546 , n732 );
buf ( n46547 , n46546 );
not ( n735 , n46547 );
buf ( n46549 , n568 );
nand ( n737 , n735 , n46549 );
buf ( n46551 , n737 );
buf ( n46552 , n46551 );
buf ( n46553 , n373 );
buf ( n46554 , n384 );
nand ( n742 , n46553 , n46554 );
buf ( n46556 , n742 );
buf ( n46557 , n46556 );
and ( n745 , n46552 , n46557 );
buf ( n46559 , n46546 );
not ( n747 , n46559 );
buf ( n46561 , n568 );
nor ( n749 , n747 , n46561 );
buf ( n46563 , n749 );
buf ( n46564 , n46563 );
nor ( n752 , n745 , n46564 );
buf ( n46566 , n752 );
not ( n754 , n46566 );
and ( n755 , n729 , n754 );
xor ( n756 , n46344 , n46339 );
xnor ( n757 , n756 , n46336 );
not ( n758 , n757 );
buf ( n46572 , n46294 );
not ( n760 , n46572 );
buf ( n46574 , n376 );
buf ( n46575 , n385 );
nand ( n763 , n46574 , n46575 );
buf ( n46577 , n763 );
buf ( n46578 , n46577 );
not ( n766 , n46578 );
buf ( n46580 , n766 );
buf ( n46581 , n46580 );
nand ( n769 , n760 , n46581 );
buf ( n46583 , n769 );
not ( n771 , n46583 );
nand ( n772 , n374 , n384 );
not ( n773 , n772 );
nand ( n774 , n377 , n381 );
not ( n775 , n774 );
or ( n776 , n773 , n775 );
buf ( n46590 , n375 );
buf ( n46591 , n383 );
nand ( n779 , n46590 , n46591 );
buf ( n46593 , n779 );
not ( n781 , n46593 );
nor ( n782 , n772 , n774 );
or ( n783 , n781 , n782 );
nand ( n784 , n776 , n783 );
not ( n785 , n784 );
nand ( n786 , n771 , n785 );
not ( n787 , n786 );
or ( n788 , n758 , n787 );
nand ( n789 , n46583 , n784 );
nand ( n790 , n788 , n789 );
nand ( n791 , n46566 , n728 );
and ( n792 , n790 , n791 );
nor ( n793 , n755 , n792 );
buf ( n46607 , n793 );
nand ( n795 , n725 , n46607 );
buf ( n46609 , n795 );
buf ( n46610 , n46609 );
not ( n798 , n46610 );
xor ( n799 , n46327 , n46346 );
xor ( n800 , n799 , n46323 );
buf ( n46614 , n800 );
not ( n802 , n46614 );
not ( n803 , n45728 );
buf ( n46617 , n45582 );
not ( n805 , n46617 );
buf ( n46619 , n805 );
not ( n807 , n46619 );
or ( n808 , n803 , n807 );
nand ( n809 , n808 , n45744 );
not ( n810 , n809 );
nor ( n811 , n45529 , n45558 );
not ( n46625 , n811 );
nand ( n813 , n46625 , n45742 );
not ( n46627 , n813 );
or ( n815 , n810 , n46627 );
or ( n816 , n809 , n813 );
nand ( n817 , n815 , n816 );
buf ( n46631 , n817 );
buf ( n46632 , n46185 );
nand ( n820 , n46631 , n46632 );
buf ( n46634 , n820 );
buf ( n46635 , n46634 );
not ( n823 , n46635 );
buf ( n46637 , n823 );
buf ( n46638 , n46637 );
not ( n826 , n46638 );
or ( n46640 , n802 , n826 );
buf ( n46641 , n800 );
not ( n829 , n46641 );
buf ( n46643 , n829 );
buf ( n46644 , n46643 );
not ( n832 , n46644 );
buf ( n46646 , n46634 );
not ( n834 , n46646 );
or ( n835 , n832 , n834 );
xor ( n836 , n46566 , n728 );
xor ( n837 , n836 , n790 );
buf ( n46651 , n837 );
nand ( n839 , n835 , n46651 );
buf ( n46653 , n839 );
buf ( n46654 , n46653 );
nand ( n842 , n46640 , n46654 );
buf ( n46656 , n842 );
buf ( n46657 , n46656 );
not ( n845 , n46657 );
or ( n846 , n798 , n845 );
buf ( n46660 , n723 );
not ( n848 , n793 );
buf ( n46662 , n848 );
nand ( n850 , n46660 , n46662 );
buf ( n46664 , n850 );
buf ( n46665 , n46664 );
nand ( n853 , n846 , n46665 );
buf ( n46667 , n853 );
buf ( n46668 , n46667 );
xor ( n856 , n46534 , n46668 );
not ( n857 , n45489 );
buf ( n46671 , n857 );
not ( n859 , n46671 );
or ( n860 , n45964 , n45961 );
not ( n861 , n860 );
not ( n862 , n45772 );
or ( n863 , n861 , n862 );
nand ( n864 , n45964 , n45961 );
nand ( n865 , n863 , n864 );
buf ( n46679 , n45916 );
buf ( n46680 , n45953 );
or ( n868 , n46679 , n46680 );
buf ( n46682 , n868 );
nand ( n870 , n46682 , n46045 );
not ( n871 , n870 );
and ( n872 , n865 , n871 );
not ( n873 , n865 );
and ( n874 , n873 , n870 );
nor ( n875 , n872 , n874 );
buf ( n46689 , n875 );
not ( n877 , n46689 );
buf ( n46691 , n877 );
and ( n879 , n411 , n46691 );
not ( n880 , n411 );
and ( n881 , n880 , n875 );
or ( n882 , n879 , n881 );
buf ( n46696 , n882 );
not ( n884 , n46696 );
or ( n885 , n859 , n884 );
buf ( n46699 , n411 );
and ( n887 , n860 , n864 );
xor ( n888 , n887 , n45773 );
buf ( n46702 , n888 );
and ( n890 , n46699 , n46702 );
not ( n891 , n46699 );
buf ( n46705 , n888 );
not ( n893 , n46705 );
buf ( n46707 , n893 );
buf ( n46708 , n46707 );
and ( n896 , n891 , n46708 );
nor ( n897 , n890 , n896 );
buf ( n46711 , n897 );
buf ( n46712 , n46711 );
buf ( n46713 , n45494 );
nand ( n901 , n46712 , n46713 );
buf ( n46715 , n901 );
buf ( n46716 , n46715 );
nand ( n904 , n885 , n46716 );
buf ( n46718 , n904 );
buf ( n46719 , n46718 );
xor ( n907 , n856 , n46719 );
buf ( n46721 , n907 );
buf ( n46722 , n46721 );
xor ( n910 , n46556 , n46546 );
and ( n911 , n910 , n727 );
not ( n912 , n910 );
and ( n913 , n912 , n568 );
nor ( n914 , n911 , n913 );
buf ( n46728 , n914 );
not ( n916 , n785 );
not ( n917 , n46583 );
or ( n918 , n916 , n917 );
nand ( n919 , n771 , n784 );
nand ( n920 , n918 , n919 );
and ( n921 , n920 , n757 );
not ( n922 , n920 );
not ( n923 , n757 );
and ( n924 , n922 , n923 );
nor ( n925 , n921 , n924 );
buf ( n46739 , n925 );
xor ( n927 , n46728 , n46739 );
buf ( n46741 , n374 );
buf ( n46742 , n385 );
nand ( n930 , n46741 , n46742 );
buf ( n46744 , n930 );
buf ( n46745 , n46744 );
not ( n933 , n46745 );
buf ( n46747 , n933 );
buf ( n46748 , n46747 );
not ( n936 , n46748 );
xor ( n937 , n774 , n46593 );
buf ( n46751 , n937 );
buf ( n46752 , n772 );
xnor ( n940 , n46751 , n46752 );
buf ( n46754 , n940 );
buf ( n46755 , n46754 );
not ( n943 , n46755 );
or ( n944 , n936 , n943 );
buf ( n46758 , n377 );
buf ( n46759 , n382 );
nand ( n947 , n46758 , n46759 );
buf ( n46761 , n947 );
buf ( n46762 , n375 );
buf ( n46763 , n384 );
nand ( n951 , n46762 , n46763 );
buf ( n46765 , n951 );
xor ( n953 , n46761 , n46765 );
nand ( n954 , n376 , n383 );
and ( n955 , n953 , n954 );
and ( n46769 , n46761 , n46765 );
nor ( n957 , n955 , n46769 );
not ( n958 , n957 );
buf ( n46772 , n958 );
nand ( n960 , n944 , n46772 );
buf ( n46774 , n960 );
buf ( n46775 , n46774 );
buf ( n46776 , n46754 );
not ( n964 , n46776 );
buf ( n46778 , n964 );
buf ( n46779 , n46778 );
buf ( n46780 , n46744 );
nand ( n968 , n46779 , n46780 );
buf ( n46782 , n968 );
buf ( n46783 , n46782 );
nand ( n971 , n46775 , n46783 );
buf ( n46785 , n971 );
buf ( n46786 , n46785 );
and ( n974 , n927 , n46786 );
and ( n975 , n46728 , n46739 );
or ( n976 , n974 , n975 );
buf ( n46790 , n976 );
buf ( n46791 , n46790 );
buf ( n46792 , n46765 );
buf ( n46793 , n46577 );
nor ( n981 , n46792 , n46793 );
buf ( n46795 , n981 );
buf ( n46796 , n46795 );
buf ( n46797 , n46744 );
nand ( n985 , n46796 , n46797 );
buf ( n46799 , n985 );
not ( n987 , n46799 );
xor ( n988 , n46761 , n46765 );
xor ( n989 , n988 , n954 );
not ( n990 , n989 );
or ( n991 , n987 , n990 );
buf ( n46805 , n46795 );
not ( n993 , n46805 );
buf ( n46807 , n993 );
buf ( n46808 , n46807 );
buf ( n46809 , n46747 );
nand ( n997 , n46808 , n46809 );
buf ( n46811 , n997 );
nand ( n999 , n991 , n46811 );
buf ( n46813 , n373 );
buf ( n46814 , n385 );
nand ( n1002 , n46813 , n46814 );
buf ( n46816 , n1002 );
buf ( n46817 , n46816 );
not ( n1005 , n46817 );
buf ( n46819 , n46274 );
not ( n1007 , n46819 );
or ( n1008 , n1005 , n1007 );
buf ( n46822 , n46583 );
nand ( n1010 , n1008 , n46822 );
buf ( n46824 , n1010 );
and ( n1012 , n999 , n46824 );
not ( n1013 , n46747 );
not ( n1014 , n957 );
or ( n1015 , n1013 , n1014 );
nand ( n1016 , n958 , n46744 );
nand ( n1017 , n1015 , n1016 );
xnor ( n1018 , n1017 , n46778 );
or ( n1019 , n1012 , n1018 );
or ( n1020 , n999 , n46824 );
nand ( n1021 , n1019 , n1020 );
buf ( n46835 , n1021 );
not ( n1023 , n46835 );
buf ( n46837 , n412 );
not ( n1025 , n46837 );
buf ( n46839 , n46153 );
nand ( n1027 , n1025 , n46839 );
buf ( n46841 , n1027 );
buf ( n46842 , n46841 );
not ( n1030 , n46842 );
buf ( n46844 , n817 );
not ( n46845 , n46844 );
or ( n1033 , n1030 , n46845 );
buf ( n46847 , n412 );
buf ( n46848 , n413 );
and ( n1036 , n46847 , n46848 );
buf ( n46850 , n411 );
not ( n46851 , n46850 );
buf ( n46852 , n46851 );
buf ( n46853 , n46852 );
nor ( n1041 , n1036 , n46853 );
buf ( n46855 , n1041 );
buf ( n46856 , n46855 );
nand ( n1044 , n1033 , n46856 );
buf ( n46858 , n1044 );
buf ( n46859 , n46858 );
not ( n1047 , n46859 );
or ( n1048 , n1023 , n1047 );
xor ( n1049 , n46728 , n46739 );
xor ( n1050 , n1049 , n46786 );
buf ( n46864 , n1050 );
buf ( n46865 , n46864 );
nand ( n1053 , n1048 , n46865 );
buf ( n46867 , n1053 );
buf ( n46868 , n46867 );
buf ( n46869 , n46858 );
buf ( n46870 , n1021 );
or ( n1058 , n46869 , n46870 );
buf ( n46872 , n1058 );
buf ( n46873 , n46872 );
nand ( n1061 , n46868 , n46873 );
buf ( n46875 , n1061 );
buf ( n46876 , n46875 );
xor ( n1064 , n46791 , n46876 );
buf ( n46878 , n800 );
buf ( n46879 , n837 );
xor ( n1067 , n46878 , n46879 );
buf ( n46881 , n46634 );
xnor ( n1069 , n1067 , n46881 );
buf ( n46883 , n1069 );
buf ( n46884 , n46883 );
and ( n1072 , n1064 , n46884 );
and ( n1073 , n46791 , n46876 );
or ( n1074 , n1072 , n1073 );
buf ( n46888 , n1074 );
buf ( n46889 , n46888 );
buf ( n46890 , n46177 );
not ( n1078 , n46890 );
xnor ( n1079 , n46153 , n875 );
buf ( n46893 , n1079 );
not ( n46894 , n46893 );
or ( n1082 , n1078 , n46894 );
buf ( n46896 , n46153 );
not ( n1084 , n46896 );
not ( n1085 , n45772 );
not ( n1086 , n45968 );
or ( n1087 , n1085 , n1086 );
buf ( n46901 , n46046 );
not ( n1089 , n46901 );
buf ( n46903 , n1089 );
nand ( n1091 , n1087 , n46903 );
not ( n46905 , n46051 );
nor ( n1093 , n46027 , n46905 );
xor ( n1094 , n1091 , n1093 );
buf ( n46908 , n1094 );
not ( n1096 , n46908 );
or ( n1097 , n1084 , n1096 );
buf ( n46911 , n1094 );
buf ( n46912 , n46153 );
or ( n1100 , n46911 , n46912 );
nand ( n1101 , n1097 , n1100 );
buf ( n46915 , n1101 );
buf ( n46916 , n46915 );
not ( n1104 , n46176 );
buf ( n46918 , n1104 );
nand ( n1106 , n46916 , n46918 );
buf ( n46920 , n1106 );
buf ( n46921 , n46920 );
nand ( n1109 , n1082 , n46921 );
buf ( n46923 , n1109 );
buf ( n46924 , n46923 );
xor ( n1112 , n46889 , n46924 );
buf ( n46926 , n415 );
not ( n1114 , n46926 );
not ( n1115 , n46035 );
nand ( n1116 , n1115 , n46049 );
not ( n1117 , n1116 );
not ( n1118 , n45968 );
not ( n1119 , n46023 );
nor ( n1120 , n1119 , n46005 );
nor ( n1121 , n1118 , n1120 );
not ( n1122 , n1121 );
not ( n1123 , n45773 );
or ( n1124 , n1122 , n1123 );
nand ( n1125 , n46044 , n46045 );
buf ( n46939 , n1125 );
buf ( n46940 , n46027 );
not ( n1128 , n46940 );
buf ( n46942 , n1128 );
buf ( n46943 , n46942 );
and ( n1131 , n46939 , n46943 );
buf ( n46945 , n46905 );
nor ( n1133 , n1131 , n46945 );
buf ( n46947 , n1133 );
nand ( n1135 , n1124 , n46947 );
not ( n1136 , n1135 );
or ( n1137 , n1117 , n1136 );
or ( n1138 , n1116 , n1135 );
nand ( n1139 , n1137 , n1138 );
buf ( n46953 , n1139 );
not ( n1141 , n46953 );
buf ( n46955 , n1141 );
buf ( n46956 , n46955 );
not ( n1144 , n46956 );
or ( n1145 , n1114 , n1144 );
and ( n1146 , n1135 , n1116 );
not ( n46960 , n1135 );
not ( n1148 , n1116 );
and ( n1149 , n46960 , n1148 );
nor ( n1150 , n1146 , n1149 );
buf ( n46964 , n1150 );
not ( n1152 , n46964 );
buf ( n46966 , n46124 );
nand ( n1154 , n1152 , n46966 );
buf ( n46968 , n1154 );
buf ( n46969 , n46968 );
nand ( n1157 , n1145 , n46969 );
buf ( n46971 , n1157 );
not ( n1159 , n46971 );
not ( n1160 , n46112 );
or ( n1161 , n1159 , n1160 );
buf ( n46975 , n415 );
and ( n1163 , n45968 , n46036 );
not ( n1164 , n1163 );
not ( n1165 , n45773 );
or ( n1166 , n1164 , n1165 );
buf ( n46980 , n46054 );
not ( n1168 , n46980 );
buf ( n46982 , n1168 );
nand ( n1170 , n1166 , n46982 );
nand ( n1171 , n45874 , n46060 );
not ( n1172 , n1171 );
and ( n1173 , n1170 , n1172 );
not ( n1174 , n1170 );
and ( n1175 , n1174 , n1171 );
nor ( n1176 , n1173 , n1175 );
buf ( n46990 , n1176 );
not ( n1178 , n46990 );
buf ( n46992 , n1178 );
buf ( n46993 , n46992 );
and ( n1181 , n46975 , n46993 );
not ( n1182 , n46975 );
buf ( n46996 , n1176 );
not ( n46997 , n46996 );
buf ( n46998 , n46997 );
buf ( n46999 , n46998 );
not ( n1187 , n46999 );
buf ( n47001 , n1187 );
buf ( n47002 , n47001 );
and ( n1190 , n1182 , n47002 );
nor ( n1191 , n1181 , n1190 );
buf ( n47005 , n1191 );
or ( n1193 , n47005 , n46108 );
nand ( n47007 , n1161 , n1193 );
buf ( n47008 , n47007 );
and ( n47009 , n1112 , n47008 );
and ( n1197 , n46889 , n46924 );
or ( n47011 , n47009 , n1197 );
buf ( n47012 , n47011 );
buf ( n47013 , n47012 );
and ( n1201 , n46722 , n47013 );
not ( n1202 , n46722 );
buf ( n47016 , n47012 );
not ( n1204 , n47016 );
buf ( n47018 , n1204 );
buf ( n47019 , n47018 );
and ( n1207 , n1202 , n47019 );
nor ( n47021 , n1201 , n1207 );
buf ( n47022 , n47021 );
not ( n1210 , n1104 );
and ( n1211 , n413 , n1150 );
not ( n1212 , n413 );
and ( n1213 , n1212 , n1139 );
or ( n1214 , n1211 , n1213 );
not ( n1215 , n1214 );
or ( n1216 , n1210 , n1215 );
buf ( n47030 , n46915 );
buf ( n47031 , n46177 );
nand ( n1219 , n47030 , n47031 );
buf ( n47033 , n1219 );
nand ( n1221 , n1216 , n47033 );
buf ( n47035 , n1221 );
buf ( n47036 , n857 );
not ( n47037 , n47036 );
buf ( n47038 , n46711 );
not ( n1226 , n47038 );
or ( n1227 , n47037 , n1226 );
and ( n47041 , n411 , n696 );
not ( n47042 , n411 );
and ( n1230 , n47042 , n46512 );
or ( n1231 , n47041 , n1230 );
buf ( n47045 , n1231 );
buf ( n47046 , n45494 );
nand ( n1234 , n47045 , n47046 );
buf ( n47048 , n1234 );
buf ( n47049 , n47048 );
nand ( n1237 , n1227 , n47049 );
buf ( n47051 , n1237 );
buf ( n47052 , n46185 );
not ( n1240 , n47052 );
buf ( n47054 , n712 );
not ( n1242 , n47054 );
or ( n1243 , n1240 , n1242 );
buf ( n47057 , n817 );
buf ( n1245 , n47057 );
buf ( n47059 , n1245 );
buf ( n47060 , n47059 );
buf ( n47061 , n46196 );
nand ( n1249 , n47060 , n47061 );
buf ( n47063 , n1249 );
buf ( n47064 , n47063 );
nand ( n1252 , n1243 , n47064 );
buf ( n47066 , n1252 );
or ( n1254 , n47051 , n47066 );
and ( n1255 , n723 , n793 );
not ( n1256 , n723 );
and ( n1257 , n1256 , n848 );
nor ( n1258 , n1255 , n1257 );
buf ( n1259 , n1258 );
not ( n1260 , n46656 );
and ( n1261 , n1259 , n1260 );
not ( n1262 , n1259 );
and ( n1263 , n1262 , n46656 );
nor ( n1264 , n1261 , n1263 );
nand ( n1265 , n1254 , n1264 );
nand ( n1266 , n47051 , n47066 );
nand ( n1267 , n1265 , n1266 );
buf ( n47081 , n1267 );
xor ( n1269 , n47035 , n47081 );
not ( n1270 , n416 );
not ( n1271 , n46067 );
nor ( n1272 , n1271 , n45832 );
not ( n1273 , n1272 );
buf ( n47087 , n46054 );
buf ( n47088 , n45874 );
nand ( n1276 , n47087 , n47088 );
buf ( n47090 , n1276 );
buf ( n47091 , n1163 );
buf ( n47092 , n45773 );
buf ( n47093 , n45874 );
nand ( n1281 , n47091 , n47092 , n47093 );
buf ( n47095 , n1281 );
nand ( n1283 , n47090 , n47095 , n46060 );
not ( n1284 , n1283 );
not ( n1285 , n1284 );
or ( n1286 , n1273 , n1285 );
not ( n1287 , n1272 );
nand ( n47101 , n1283 , n1287 );
nand ( n47102 , n1286 , n47101 );
xor ( n1290 , n415 , n47102 );
not ( n1291 , n1290 );
or ( n1292 , n1270 , n1291 );
not ( n47106 , n47005 );
nand ( n47107 , n47106 , n46112 );
nand ( n1295 , n1292 , n47107 );
buf ( n47109 , n1295 );
xnor ( n1297 , n1269 , n47109 );
buf ( n47111 , n1297 );
xor ( n1299 , n47022 , n47111 );
buf ( n47113 , n1299 );
xor ( n1301 , n46889 , n46924 );
xor ( n1302 , n1301 , n47008 );
buf ( n47116 , n1302 );
buf ( n47117 , n47116 );
not ( n1305 , n47117 );
buf ( n47119 , n1305 );
not ( n1307 , n47119 );
buf ( n47121 , n1258 );
buf ( n47122 , n47066 );
xor ( n1310 , n47121 , n47122 );
buf ( n47124 , n46656 );
xor ( n1312 , n1310 , n47124 );
buf ( n47126 , n1312 );
buf ( n47127 , n47126 );
buf ( n47128 , n47051 );
not ( n1316 , n47128 );
buf ( n47130 , n1316 );
buf ( n47131 , n47130 );
and ( n1319 , n47127 , n47131 );
not ( n1320 , n47127 );
buf ( n47134 , n47051 );
and ( n1322 , n1320 , n47134 );
nor ( n47136 , n1319 , n1322 );
buf ( n47137 , n47136 );
buf ( n47138 , n47137 );
not ( n1326 , n47138 );
buf ( n47140 , n1326 );
not ( n1328 , n47140 );
and ( n1329 , n1307 , n1328 );
buf ( n47143 , n47119 );
buf ( n47144 , n47140 );
nand ( n1332 , n47143 , n47144 );
buf ( n47146 , n1332 );
buf ( n47147 , n857 );
not ( n1335 , n47147 );
buf ( n47149 , n1231 );
not ( n1337 , n47149 );
or ( n1338 , n1335 , n1337 );
buf ( n47152 , n712 );
not ( n1340 , n47152 );
buf ( n47154 , n1340 );
and ( n1342 , n411 , n47154 );
not ( n1343 , n411 );
and ( n1344 , n1343 , n712 );
or ( n1345 , n1342 , n1344 );
buf ( n47159 , n1345 );
buf ( n47160 , n45494 );
nand ( n1348 , n47159 , n47160 );
buf ( n47162 , n1348 );
buf ( n47163 , n47162 );
nand ( n1351 , n1338 , n47163 );
buf ( n47165 , n1351 );
buf ( n47166 , n47165 );
xor ( n1354 , n46791 , n46876 );
xor ( n1355 , n1354 , n46884 );
buf ( n47169 , n1355 );
buf ( n47170 , n47169 );
xor ( n1358 , n47166 , n47170 );
buf ( n47172 , n1104 );
not ( n1360 , n47172 );
buf ( n47174 , n1079 );
not ( n1362 , n47174 );
or ( n1363 , n1360 , n1362 );
buf ( n47177 , n413 );
not ( n1365 , n47177 );
buf ( n47179 , n46707 );
not ( n1367 , n47179 );
or ( n1368 , n1365 , n1367 );
buf ( n47182 , n888 );
buf ( n47183 , n46153 );
nand ( n1371 , n47182 , n47183 );
buf ( n47185 , n1371 );
buf ( n47186 , n47185 );
nand ( n1374 , n1368 , n47186 );
buf ( n47188 , n1374 );
buf ( n47189 , n47188 );
buf ( n47190 , n46177 );
nand ( n1378 , n47189 , n47190 );
buf ( n47192 , n1378 );
buf ( n47193 , n47192 );
nand ( n1381 , n1363 , n47193 );
buf ( n47195 , n1381 );
buf ( n47196 , n47195 );
and ( n1384 , n1358 , n47196 );
and ( n1385 , n47166 , n47170 );
or ( n1386 , n1384 , n1385 );
buf ( n47200 , n1386 );
and ( n1388 , n47146 , n47200 );
nor ( n1389 , n1329 , n1388 );
buf ( n47203 , n1389 );
nand ( n1391 , n47113 , n47203 );
buf ( n47205 , n1391 );
buf ( n47206 , n47205 );
buf ( n1394 , n47206 );
buf ( n47208 , n1394 );
buf ( n47209 , n47208 );
not ( n1397 , n47209 );
xor ( n1398 , n46858 , n1021 );
xor ( n1399 , n1398 , n46864 );
buf ( n47213 , n1399 );
buf ( n47214 , n857 );
not ( n1402 , n47214 );
buf ( n47216 , n1345 );
not ( n1404 , n47216 );
or ( n1405 , n1402 , n1404 );
buf ( n47219 , n47059 );
not ( n1407 , n47219 );
buf ( n47221 , n1407 );
and ( n1409 , n411 , n47221 );
not ( n1410 , n411 );
and ( n1411 , n1410 , n47059 );
or ( n1412 , n1409 , n1411 );
buf ( n47226 , n1412 );
buf ( n47227 , n45494 );
nand ( n47228 , n47226 , n47227 );
buf ( n47229 , n47228 );
buf ( n47230 , n47229 );
nand ( n1418 , n1405 , n47230 );
buf ( n47232 , n1418 );
buf ( n47233 , n47232 );
xor ( n1421 , n47213 , n47233 );
buf ( n47235 , n1104 );
not ( n1423 , n47235 );
buf ( n47237 , n47188 );
not ( n1425 , n47237 );
or ( n1426 , n1423 , n1425 );
buf ( n47240 , n413 );
not ( n1428 , n47240 );
buf ( n47242 , n696 );
not ( n1430 , n47242 );
or ( n1431 , n1428 , n1430 );
nand ( n1432 , n46512 , n46153 );
buf ( n47246 , n1432 );
nand ( n1434 , n1431 , n47246 );
buf ( n47248 , n1434 );
buf ( n47249 , n47248 );
buf ( n47250 , n46177 );
nand ( n1438 , n47249 , n47250 );
buf ( n47252 , n1438 );
buf ( n47253 , n47252 );
nand ( n1441 , n1426 , n47253 );
buf ( n47255 , n1441 );
buf ( n47256 , n47255 );
and ( n1444 , n1421 , n47256 );
and ( n1445 , n47213 , n47233 );
or ( n1446 , n1444 , n1445 );
buf ( n47260 , n1446 );
buf ( n47261 , n47260 );
not ( n47262 , n47261 );
buf ( n47263 , n416 );
not ( n1451 , n47263 );
buf ( n47265 , n46971 );
not ( n1453 , n47265 );
or ( n1454 , n1451 , n1453 );
buf ( n47268 , n415 );
buf ( n47269 , n1094 );
and ( n1457 , n47268 , n47269 );
not ( n1458 , n47268 );
buf ( n47272 , n1094 );
not ( n1460 , n47272 );
buf ( n47274 , n1460 );
buf ( n47275 , n47274 );
and ( n1463 , n1458 , n47275 );
nor ( n1464 , n1457 , n1463 );
buf ( n47278 , n1464 );
buf ( n47279 , n47278 );
buf ( n47280 , n46112 );
nand ( n1468 , n47279 , n47280 );
buf ( n47282 , n1468 );
buf ( n47283 , n47282 );
nand ( n1471 , n1454 , n47283 );
buf ( n47285 , n1471 );
buf ( n47286 , n47285 );
not ( n1474 , n47286 );
buf ( n47288 , n1474 );
buf ( n47289 , n47288 );
nand ( n1477 , n47262 , n47289 );
buf ( n47291 , n1477 );
buf ( n47292 , n47291 );
not ( n1480 , n47292 );
xor ( n47294 , n47166 , n47170 );
xor ( n47295 , n47294 , n47196 );
buf ( n47296 , n47295 );
buf ( n47297 , n47296 );
not ( n1485 , n47297 );
or ( n1486 , n1480 , n1485 );
buf ( n47300 , n47288 );
not ( n1488 , n47300 );
buf ( n47302 , n47260 );
nand ( n1490 , n1488 , n47302 );
buf ( n47304 , n1490 );
buf ( n47305 , n47304 );
nand ( n1493 , n1486 , n47305 );
buf ( n47307 , n1493 );
buf ( n47308 , n47307 );
not ( n1496 , n47308 );
buf ( n47310 , n47137 );
buf ( n47311 , n47200 );
xor ( n1499 , n47310 , n47311 );
buf ( n47313 , n47116 );
xnor ( n1501 , n1499 , n47313 );
buf ( n47315 , n1501 );
buf ( n47316 , n47315 );
nand ( n1504 , n1496 , n47316 );
buf ( n47318 , n1504 );
buf ( n47319 , n47318 );
buf ( n47320 , n416 );
not ( n1508 , n47320 );
buf ( n47322 , n415 );
not ( n1510 , n47322 );
buf ( n47324 , n46691 );
not ( n1512 , n47324 );
or ( n1513 , n1510 , n1512 );
buf ( n47327 , n46124 );
buf ( n47328 , n875 );
nand ( n1516 , n47327 , n47328 );
buf ( n47330 , n1516 );
buf ( n47331 , n47330 );
nand ( n1519 , n1513 , n47331 );
buf ( n47333 , n1519 );
buf ( n47334 , n47333 );
not ( n1522 , n47334 );
or ( n1523 , n1508 , n1522 );
buf ( n47337 , n415 );
buf ( n47338 , n888 );
and ( n1526 , n47337 , n47338 );
not ( n1527 , n47337 );
buf ( n47341 , n46707 );
and ( n1529 , n1527 , n47341 );
nor ( n1530 , n1526 , n1529 );
buf ( n47344 , n1530 );
buf ( n47345 , n47344 );
buf ( n47346 , n46112 );
nand ( n1534 , n47345 , n47346 );
buf ( n47348 , n1534 );
buf ( n47349 , n47348 );
nand ( n1537 , n1523 , n47349 );
buf ( n47351 , n1537 );
buf ( n47352 , n47351 );
xor ( n1540 , n712 , n46153 );
not ( n1541 , n1540 );
not ( n1542 , n46180 );
and ( n1543 , n1541 , n1542 );
and ( n1544 , n47248 , n1104 );
nor ( n1545 , n1543 , n1544 );
buf ( n47359 , n1545 );
not ( n47360 , n47359 );
buf ( n47361 , n47360 );
buf ( n47362 , n47361 );
nor ( n1550 , n47352 , n47362 );
buf ( n47364 , n1550 );
buf ( n47365 , n47364 );
buf ( n47366 , n1018 );
not ( n1554 , n47366 );
buf ( n47368 , n999 );
buf ( n47369 , n46824 );
not ( n1557 , n47369 );
xor ( n1558 , n47368 , n1557 );
buf ( n47372 , n1558 );
buf ( n47373 , n47372 );
not ( n1561 , n47373 );
or ( n1562 , n1554 , n1561 );
buf ( n47376 , n47372 );
buf ( n47377 , n1018 );
or ( n1565 , n47376 , n47377 );
nand ( n1566 , n1562 , n1565 );
buf ( n47380 , n1566 );
not ( n1568 , n47380 );
buf ( n47382 , n47059 );
buf ( n47383 , n857 );
nand ( n1571 , n47382 , n47383 );
buf ( n47385 , n1571 );
not ( n1573 , n47385 );
and ( n1574 , n1568 , n1573 );
and ( n1575 , n47380 , n47385 );
nor ( n1576 , n1574 , n1575 );
buf ( n47390 , n989 );
buf ( n47391 , n46807 );
buf ( n47392 , n46747 );
and ( n47393 , n47391 , n47392 );
not ( n47394 , n47391 );
buf ( n47395 , n46744 );
and ( n1583 , n47394 , n47395 );
nor ( n1584 , n47393 , n1583 );
buf ( n47398 , n1584 );
buf ( n47399 , n47398 );
xnor ( n1587 , n47390 , n47399 );
buf ( n47401 , n1587 );
not ( n1589 , n47401 );
buf ( n47403 , n375 );
buf ( n47404 , n385 );
and ( n1592 , n47403 , n47404 );
buf ( n47406 , n376 );
buf ( n47407 , n384 );
and ( n1595 , n47406 , n47407 );
nor ( n1596 , n1592 , n1595 );
buf ( n47410 , n1596 );
buf ( n47411 , n47410 );
not ( n1599 , n47411 );
buf ( n47413 , n46807 );
nand ( n1601 , n1599 , n47413 );
buf ( n47415 , n1601 );
buf ( n47416 , n47415 );
buf ( n47417 , n377 );
buf ( n47418 , n383 );
nand ( n1606 , n47417 , n47418 );
buf ( n47420 , n1606 );
buf ( n47421 , n47420 );
buf ( n47422 , n46577 );
or ( n1610 , n47421 , n47422 );
buf ( n47424 , n1610 );
buf ( n47425 , n47424 );
and ( n47426 , n47416 , n47425 );
buf ( n47427 , n47420 );
buf ( n47428 , n46577 );
and ( n1616 , n47427 , n47428 );
nor ( n1617 , n47426 , n1616 );
buf ( n47431 , n1617 );
not ( n1619 , n47431 );
nand ( n1620 , n1589 , n1619 );
not ( n1621 , n1620 );
buf ( n47435 , n46175 );
not ( n1623 , n47435 );
buf ( n47437 , n817 );
not ( n1625 , n47437 );
or ( n1626 , n1623 , n1625 );
buf ( n47440 , n414 );
buf ( n47441 , n415 );
and ( n1629 , n47440 , n47441 );
buf ( n47443 , n46153 );
nor ( n1631 , n1629 , n47443 );
buf ( n47445 , n1631 );
buf ( n47446 , n47445 );
nand ( n1634 , n1626 , n47446 );
buf ( n47448 , n1634 );
not ( n1636 , n47448 );
or ( n1637 , n1621 , n1636 );
nand ( n1638 , n47401 , n47431 );
nand ( n1639 , n1637 , n1638 );
and ( n1640 , n1576 , n1639 );
not ( n1641 , n1576 );
not ( n1642 , n1639 );
and ( n1643 , n1641 , n1642 );
nor ( n1644 , n1640 , n1643 );
not ( n1645 , n1644 );
buf ( n47459 , n1645 );
or ( n47460 , n47365 , n47459 );
buf ( n47461 , n47351 );
buf ( n47462 , n47361 );
nand ( n1650 , n47461 , n47462 );
buf ( n47464 , n1650 );
buf ( n47465 , n47464 );
nand ( n1653 , n47460 , n47465 );
buf ( n47467 , n1653 );
not ( n1655 , n47467 );
buf ( n47469 , n47380 );
not ( n1657 , n47469 );
buf ( n47471 , n47385 );
nand ( n1659 , n1657 , n47471 );
buf ( n47473 , n1659 );
buf ( n47474 , n47473 );
not ( n1662 , n47474 );
buf ( n47476 , n1642 );
not ( n1664 , n47476 );
or ( n1665 , n1662 , n1664 );
buf ( n47479 , n47385 );
not ( n1667 , n47479 );
buf ( n47481 , n47380 );
nand ( n1669 , n1667 , n47481 );
buf ( n47483 , n1669 );
buf ( n47484 , n47483 );
nand ( n1672 , n1665 , n47484 );
buf ( n47486 , n1672 );
buf ( n47487 , n47486 );
buf ( n47488 , n46112 );
not ( n1676 , n47488 );
buf ( n47490 , n47333 );
not ( n1678 , n47490 );
or ( n47492 , n1676 , n1678 );
buf ( n47493 , n47278 );
buf ( n47494 , n416 );
nand ( n1682 , n47493 , n47494 );
buf ( n47496 , n1682 );
buf ( n47497 , n47496 );
nand ( n1685 , n47492 , n47497 );
buf ( n47499 , n1685 );
buf ( n47500 , n47499 );
xor ( n1688 , n47487 , n47500 );
xor ( n1689 , n47213 , n47233 );
xor ( n1690 , n1689 , n47256 );
buf ( n47504 , n1690 );
buf ( n47505 , n47504 );
xnor ( n1693 , n1688 , n47505 );
buf ( n47507 , n1693 );
nand ( n1695 , n1655 , n47507 );
not ( n1696 , n1695 );
buf ( n47510 , n413 );
not ( n1698 , n47510 );
buf ( n47512 , n47221 );
not ( n1700 , n47512 );
or ( n1701 , n1698 , n1700 );
buf ( n47515 , n47059 );
buf ( n47516 , n46153 );
nand ( n1704 , n47515 , n47516 );
buf ( n47518 , n1704 );
buf ( n47519 , n47518 );
nand ( n1707 , n1701 , n47519 );
buf ( n47521 , n1707 );
not ( n1709 , n47521 );
not ( n1710 , n46177 );
or ( n1711 , n1709 , n1710 );
or ( n47525 , n1540 , n46176 );
nand ( n47526 , n1711 , n47525 );
buf ( n47527 , n47526 );
not ( n1715 , n47527 );
buf ( n47529 , n1715 );
buf ( n47530 , n47529 );
not ( n1718 , n47530 );
buf ( n47532 , n416 );
not ( n1720 , n47532 );
buf ( n47534 , n47344 );
not ( n1722 , n47534 );
or ( n1723 , n1720 , n1722 );
buf ( n47537 , n415 );
buf ( n47538 , n46512 );
and ( n1726 , n47537 , n47538 );
not ( n1727 , n47537 );
buf ( n47541 , n696 );
and ( n1729 , n1727 , n47541 );
nor ( n1730 , n1726 , n1729 );
buf ( n47544 , n1730 );
buf ( n47545 , n47544 );
buf ( n47546 , n46112 );
nand ( n1734 , n47545 , n47546 );
buf ( n47548 , n1734 );
buf ( n47549 , n47548 );
nand ( n1737 , n1723 , n47549 );
buf ( n47551 , n1737 );
buf ( n47552 , n47551 );
not ( n1740 , n47552 );
buf ( n47554 , n1740 );
buf ( n47555 , n47554 );
not ( n1743 , n47555 );
or ( n1744 , n1718 , n1743 );
not ( n47558 , n47448 );
not ( n47559 , n1619 );
not ( n1747 , n47401 );
or ( n1748 , n47559 , n1747 );
nand ( n1749 , n1589 , n47431 );
nand ( n1750 , n1748 , n1749 );
and ( n1751 , n47558 , n1750 );
not ( n1752 , n47558 );
not ( n1753 , n1750 );
and ( n1754 , n1752 , n1753 );
nor ( n1755 , n1751 , n1754 );
buf ( n47569 , n1755 );
nand ( n1757 , n1744 , n47569 );
buf ( n47571 , n1757 );
buf ( n47572 , n47571 );
buf ( n47573 , n47554 );
not ( n1761 , n47573 );
buf ( n47575 , n47526 );
nand ( n1763 , n1761 , n47575 );
buf ( n47577 , n1763 );
buf ( n47578 , n47577 );
nand ( n1766 , n47572 , n47578 );
buf ( n47580 , n1766 );
buf ( n47581 , n47580 );
not ( n1769 , n47581 );
buf ( n47583 , n47351 );
not ( n1771 , n47583 );
not ( n1772 , n1545 );
not ( n1773 , n1645 );
or ( n1774 , n1772 , n1773 );
or ( n1775 , n1645 , n1545 );
nand ( n1776 , n1774 , n1775 );
buf ( n47590 , n1776 );
not ( n47591 , n47590 );
and ( n47592 , n1771 , n47591 );
buf ( n47593 , n47351 );
buf ( n47594 , n1776 );
and ( n1782 , n47593 , n47594 );
nor ( n1783 , n47592 , n1782 );
buf ( n47597 , n1783 );
buf ( n47598 , n47597 );
nand ( n1786 , n1769 , n47598 );
buf ( n47600 , n1786 );
not ( n1788 , n47600 );
xor ( n1789 , n1755 , n47526 );
xnor ( n1790 , n1789 , n47554 );
buf ( n47604 , n1790 );
buf ( n47605 , n377 );
buf ( n47606 , n384 );
nand ( n1794 , n47605 , n47606 );
buf ( n47608 , n1794 );
buf ( n47609 , n47608 );
not ( n1797 , n47609 );
buf ( n47611 , n46577 );
nand ( n1799 , n1797 , n47611 );
buf ( n47613 , n1799 );
buf ( n47614 , n47613 );
not ( n1802 , n47614 );
buf ( n47616 , n47059 );
buf ( n47617 , n416 );
nand ( n1805 , n47616 , n47617 );
buf ( n47619 , n1805 );
buf ( n47620 , n47619 );
buf ( n47621 , n415 );
nand ( n1809 , n47620 , n47621 );
buf ( n47623 , n1809 );
buf ( n47624 , n47623 );
not ( n47625 , n47624 );
buf ( n47626 , n47625 );
buf ( n47627 , n47626 );
not ( n1815 , n47627 );
or ( n1816 , n1802 , n1815 );
buf ( n47630 , n46580 );
buf ( n47631 , n47608 );
nand ( n1819 , n47630 , n47631 );
buf ( n47633 , n1819 );
buf ( n47634 , n47633 );
nand ( n1822 , n1816 , n47634 );
buf ( n47636 , n1822 );
not ( n1824 , n47636 );
buf ( n47638 , n47059 );
buf ( n47639 , n1104 );
nand ( n1827 , n47638 , n47639 );
buf ( n47641 , n1827 );
or ( n1829 , n1824 , n47641 );
buf ( n47643 , n47641 );
not ( n1831 , n47643 );
buf ( n47645 , n1824 );
not ( n1833 , n47645 );
or ( n1834 , n1831 , n1833 );
buf ( n47648 , n47420 );
buf ( n47649 , n46577 );
and ( n1837 , n47648 , n47649 );
not ( n1838 , n47648 );
buf ( n47652 , n46580 );
and ( n1840 , n1838 , n47652 );
nor ( n1841 , n1837 , n1840 );
buf ( n47655 , n1841 );
buf ( n47656 , n47655 );
not ( n47657 , n47656 );
buf ( n47658 , n47415 );
not ( n1846 , n47658 );
buf ( n47660 , n1846 );
buf ( n47661 , n47660 );
not ( n1849 , n47661 );
or ( n1850 , n47657 , n1849 );
buf ( n47664 , n47660 );
buf ( n47665 , n47655 );
or ( n1853 , n47664 , n47665 );
nand ( n1854 , n1850 , n1853 );
buf ( n47668 , n1854 );
buf ( n47669 , n47668 );
nand ( n1857 , n1834 , n47669 );
buf ( n47671 , n1857 );
nand ( n1859 , n1829 , n47671 );
buf ( n47673 , n1859 );
nor ( n1861 , n47604 , n47673 );
buf ( n47675 , n1861 );
buf ( n47676 , n47675 );
xor ( n1864 , n47668 , n47641 );
and ( n1865 , n1864 , n47636 );
not ( n1866 , n1864 );
and ( n1867 , n1866 , n1824 );
nor ( n1868 , n1865 , n1867 );
buf ( n47682 , n47544 );
buf ( n47683 , n416 );
nand ( n1871 , n47682 , n47683 );
buf ( n47685 , n1871 );
buf ( n47686 , n415 );
not ( n1874 , n47686 );
buf ( n47688 , n47154 );
not ( n1876 , n47688 );
or ( n47690 , n1874 , n1876 );
buf ( n47691 , n712 );
buf ( n47692 , n46124 );
nand ( n1880 , n47691 , n47692 );
buf ( n47694 , n1880 );
buf ( n47695 , n47694 );
nand ( n1883 , n47690 , n47695 );
buf ( n47697 , n1883 );
buf ( n47698 , n47697 );
buf ( n47699 , n46112 );
nand ( n1887 , n47698 , n47699 );
buf ( n47701 , n1887 );
nand ( n1889 , n1868 , n47685 , n47701 );
buf ( n47703 , n416 );
not ( n1891 , n47703 );
buf ( n47705 , n47697 );
not ( n1893 , n47705 );
or ( n1894 , n1891 , n1893 );
buf ( n47708 , n47221 );
buf ( n47709 , n46112 );
nand ( n1897 , n47708 , n47709 );
buf ( n47711 , n1897 );
buf ( n47712 , n47711 );
nand ( n1900 , n1894 , n47712 );
buf ( n47714 , n1900 );
buf ( n47715 , n47714 );
buf ( n47716 , n47608 );
not ( n1904 , n47716 );
buf ( n47718 , n46577 );
not ( n1906 , n47718 );
and ( n1907 , n1904 , n1906 );
buf ( n47721 , n47608 );
buf ( n47722 , n46577 );
and ( n47723 , n47721 , n47722 );
nor ( n47724 , n1907 , n47723 );
buf ( n47725 , n47724 );
buf ( n47726 , n47725 );
not ( n1914 , n47726 );
buf ( n47728 , n47626 );
not ( n1916 , n47728 );
or ( n1917 , n1914 , n1916 );
buf ( n47731 , n47626 );
buf ( n47732 , n47725 );
or ( n1920 , n47731 , n47732 );
nand ( n1921 , n1917 , n1920 );
buf ( n47735 , n1921 );
buf ( n47736 , n47735 );
nor ( n1924 , n47715 , n47736 );
buf ( n47738 , n1924 );
buf ( n47739 , n47738 );
buf ( n47740 , n47619 );
buf ( n47741 , n377 );
buf ( n47742 , n385 );
and ( n1930 , n47741 , n47742 );
buf ( n47744 , n1930 );
buf ( n47745 , n47744 );
nand ( n1933 , n47740 , n47745 );
buf ( n47747 , n1933 );
buf ( n47748 , n47747 );
not ( n1936 , n47748 );
buf ( n47750 , n1936 );
buf ( n47751 , n47750 );
or ( n1939 , n47739 , n47751 );
buf ( n47753 , n47714 );
buf ( n47754 , n47735 );
nand ( n1942 , n47753 , n47754 );
buf ( n47756 , n1942 );
buf ( n47757 , n47756 );
nand ( n1945 , n1939 , n47757 );
buf ( n47759 , n1945 );
and ( n1947 , n1889 , n47759 );
buf ( n47761 , n1868 );
not ( n1949 , n47761 );
buf ( n47763 , n1949 );
and ( n1951 , n47544 , n416 );
and ( n1952 , n47697 , n46112 );
nor ( n1953 , n1951 , n1952 );
buf ( n47767 , n1953 );
not ( n1955 , n47767 );
buf ( n47769 , n1955 );
and ( n1957 , n47763 , n47769 );
nor ( n1958 , n1947 , n1957 );
buf ( n47772 , n1958 );
or ( n1960 , n47676 , n47772 );
buf ( n47774 , n1790 );
buf ( n47775 , n1859 );
nand ( n1963 , n47774 , n47775 );
buf ( n47777 , n1963 );
buf ( n47778 , n47777 );
nand ( n1966 , n1960 , n47778 );
buf ( n47780 , n1966 );
not ( n1968 , n47780 );
or ( n1969 , n1788 , n1968 );
not ( n1970 , n47597 );
nand ( n1971 , n1970 , n47580 );
nand ( n1972 , n1969 , n1971 );
not ( n1973 , n1972 );
or ( n1974 , n1696 , n1973 );
not ( n1975 , n47507 );
buf ( n47789 , n47364 );
buf ( n47790 , n1645 );
or ( n1978 , n47789 , n47790 );
buf ( n47792 , n47464 );
nand ( n1980 , n1978 , n47792 );
buf ( n47794 , n1980 );
nand ( n1982 , n1975 , n47794 );
nand ( n1983 , n1974 , n1982 );
buf ( n47797 , n1983 );
not ( n1985 , n47486 );
buf ( n47799 , n46112 );
not ( n1987 , n47799 );
buf ( n47801 , n47333 );
not ( n1989 , n47801 );
or ( n1990 , n1987 , n1989 );
buf ( n47804 , n47496 );
nand ( n1992 , n1990 , n47804 );
buf ( n47806 , n1992 );
not ( n1994 , n47806 );
nand ( n1995 , n1985 , n1994 );
not ( n1996 , n1995 );
not ( n1997 , n47504 );
or ( n1998 , n1996 , n1997 );
not ( n1999 , n1994 );
nand ( n2000 , n1999 , n47486 );
nand ( n2001 , n1998 , n2000 );
buf ( n47815 , n2001 );
not ( n2003 , n47815 );
not ( n2004 , n47288 );
and ( n2005 , n47260 , n2004 );
not ( n2006 , n47260 );
and ( n2007 , n2006 , n47288 );
nor ( n2008 , n2005 , n2007 );
not ( n47822 , n47296 );
and ( n47823 , n2008 , n47822 );
not ( n2011 , n2008 );
and ( n2012 , n2011 , n47296 );
nor ( n2013 , n47823 , n2012 );
buf ( n47827 , n2013 );
nand ( n2015 , n2003 , n47827 );
buf ( n47829 , n2015 );
buf ( n47830 , n47829 );
nand ( n2018 , n47797 , n47830 );
buf ( n47832 , n2018 );
buf ( n47833 , n47832 );
not ( n2021 , n2013 );
nand ( n2022 , n2021 , n2001 );
buf ( n47836 , n2022 );
nand ( n2024 , n47833 , n47836 );
buf ( n47838 , n2024 );
buf ( n47839 , n47838 );
and ( n2027 , n47319 , n47839 );
buf ( n47841 , n2027 );
buf ( n47842 , n47841 );
not ( n2030 , n47842 );
or ( n2031 , n1397 , n2030 );
not ( n2032 , n47205 );
buf ( n47846 , n47307 );
not ( n2034 , n47846 );
buf ( n47848 , n47315 );
nor ( n2036 , n2034 , n47848 );
buf ( n47850 , n2036 );
not ( n2038 , n47850 );
or ( n2039 , n2032 , n2038 );
buf ( n47853 , n1299 );
not ( n2041 , n47853 );
buf ( n47855 , n2041 );
buf ( n47856 , n47855 );
buf ( n47857 , n1389 );
not ( n2045 , n47857 );
buf ( n47859 , n2045 );
buf ( n47860 , n47859 );
nand ( n2048 , n47856 , n47860 );
buf ( n47862 , n2048 );
nand ( n2050 , n2039 , n47862 );
buf ( n47864 , n2050 );
not ( n2052 , n47864 );
buf ( n47866 , n2052 );
buf ( n47867 , n47866 );
nand ( n2055 , n2031 , n47867 );
buf ( n47869 , n2055 );
not ( n2057 , n47869 );
not ( n2058 , n46177 );
not ( n2059 , n413 );
not ( n2060 , n46998 );
or ( n2061 , n2059 , n2060 );
buf ( n47875 , n46153 );
buf ( n47876 , n1176 );
nand ( n2064 , n47875 , n47876 );
buf ( n47878 , n2064 );
nand ( n2066 , n2061 , n47878 );
not ( n2067 , n2066 );
or ( n2068 , n2058 , n2067 );
xnor ( n2069 , n1272 , n413 );
and ( n2070 , n2069 , n1283 );
not ( n2071 , n2069 );
and ( n2072 , n2071 , n1284 );
or ( n2073 , n2070 , n2072 );
nand ( n2074 , n2073 , n1104 );
nand ( n47888 , n2068 , n2074 );
not ( n47889 , n47888 );
xor ( n2077 , n596 , n619 );
and ( n2078 , n2077 , n670 );
and ( n2079 , n596 , n619 );
or ( n2080 , n2078 , n2079 );
not ( n2081 , n2080 );
nand ( n2082 , n381 , n372 );
not ( n2083 , n2082 );
nand ( n2084 , n373 , n380 );
nand ( n2085 , n383 , n370 );
nor ( n2086 , n2083 , n2084 , n2085 );
not ( n2087 , n2086 );
nand ( n2088 , n381 , n372 );
nand ( n2089 , n2084 , n2088 , n2085 );
not ( n2090 , n2085 );
nand ( n2091 , n2090 , n2083 , n2084 );
not ( n2092 , n2084 );
not ( n2093 , n2088 );
nand ( n2094 , n2092 , n2093 , n2085 );
nand ( n2095 , n2087 , n2089 , n2091 , n2094 );
not ( n2096 , n2095 );
not ( n2097 , n657 );
not ( n2098 , n603 );
nand ( n2099 , n374 , n380 );
not ( n2100 , n2099 );
or ( n2101 , n2098 , n2100 );
or ( n2102 , n2099 , n46364 );
nand ( n2103 , n2102 , n605 );
nand ( n2104 , n2101 , n2103 );
and ( n2105 , n2097 , n2104 );
and ( n2106 , n2096 , n2105 );
not ( n2107 , n2096 );
nor ( n47921 , n657 , n2104 );
and ( n47922 , n2107 , n47921 );
nor ( n2110 , n2106 , n47922 );
nand ( n2111 , n2095 , n2104 );
or ( n2112 , n2111 , n2097 );
not ( n2113 , n2104 );
nand ( n2114 , n2113 , n2096 , n657 );
and ( n2115 , n2110 , n2112 , n2114 );
not ( n2116 , n46476 );
not ( n2117 , n641 );
not ( n2118 , n2117 );
or ( n2119 , n2116 , n2118 );
nand ( n2120 , n2119 , n668 );
not ( n2121 , n46476 );
nand ( n2122 , n2121 , n641 );
nand ( n2123 , n2120 , n2122 );
xor ( n2124 , n2115 , n2123 );
buf ( n47938 , n46444 );
not ( n2126 , n47938 );
buf ( n47940 , n46440 );
nand ( n2128 , n2126 , n47940 );
buf ( n47942 , n2128 );
buf ( n47943 , n47942 );
not ( n2131 , n47943 );
buf ( n47945 , n640 );
not ( n2133 , n47945 );
or ( n2134 , n2131 , n2133 );
buf ( n47948 , n46437 );
buf ( n47949 , n46444 );
nand ( n2137 , n47948 , n47949 );
buf ( n47951 , n2137 );
buf ( n47952 , n47951 );
nand ( n2140 , n2134 , n47952 );
buf ( n47954 , n2140 );
not ( n47955 , n47954 );
buf ( n47956 , n374 );
buf ( n47957 , n379 );
nand ( n2145 , n47956 , n47957 );
buf ( n47959 , n2145 );
buf ( n47960 , n375 );
buf ( n47961 , n378 );
nand ( n2149 , n47960 , n47961 );
buf ( n47963 , n2149 );
xor ( n2151 , n47959 , n47963 );
buf ( n47965 , n371 );
buf ( n47966 , n382 );
nand ( n2154 , n47965 , n47966 );
buf ( n47968 , n2154 );
xnor ( n2156 , n2151 , n47968 );
xor ( n2157 , n47955 , n2156 );
not ( n2158 , n602 );
not ( n2159 , n609 );
or ( n2160 , n2158 , n2159 );
nand ( n2161 , n2160 , n610 );
xor ( n2162 , n2157 , n2161 );
xnor ( n2163 , n2124 , n2162 );
not ( n2164 , n2163 );
nand ( n2165 , n2081 , n2164 );
not ( n2166 , n2165 );
buf ( n47980 , n46185 );
not ( n2168 , n47980 );
buf ( n47982 , n888 );
not ( n2170 , n47982 );
or ( n2171 , n2168 , n2170 );
buf ( n47985 , n46512 );
buf ( n47986 , n46196 );
nand ( n47987 , n47985 , n47986 );
buf ( n47988 , n47987 );
buf ( n47989 , n47988 );
nand ( n2177 , n2171 , n47989 );
buf ( n47991 , n2177 );
not ( n2179 , n47991 );
or ( n2180 , n2166 , n2179 );
nand ( n2181 , n2163 , n2080 );
nand ( n2182 , n2180 , n2181 );
not ( n2183 , n2182 );
not ( n2184 , n46185 );
not ( n2185 , n875 );
or ( n2186 , n2184 , n2185 );
buf ( n48000 , n888 );
buf ( n48001 , n46196 );
nand ( n2189 , n48000 , n48001 );
buf ( n48003 , n2189 );
nand ( n2191 , n2186 , n48003 );
not ( n2192 , n2191 );
not ( n2193 , n2192 );
and ( n2194 , n2183 , n2193 );
and ( n2195 , n2182 , n2192 );
nor ( n2196 , n2194 , n2195 );
not ( n2197 , n2196 );
or ( n2198 , n47889 , n2197 );
or ( n2199 , n47888 , n2196 );
nand ( n2200 , n2198 , n2199 );
not ( n2201 , n2200 );
xor ( n2202 , n2080 , n2164 );
xnor ( n2203 , n2202 , n47991 );
buf ( n48017 , n2203 );
buf ( n48018 , n46112 );
not ( n2206 , n48018 );
buf ( n48020 , n1290 );
not ( n48021 , n48020 );
or ( n2209 , n2206 , n48021 );
nand ( n2210 , n45788 , n46078 );
xor ( n2211 , n2210 , n415 );
not ( n2212 , n45875 );
nand ( n2213 , n45773 , n1163 , n2212 );
nand ( n2214 , n2212 , n46054 );
not ( n2215 , n46070 );
nand ( n2216 , n2213 , n2214 , n2215 );
xnor ( n2217 , n2211 , n2216 );
buf ( n48031 , n2217 );
buf ( n48032 , n416 );
nand ( n2220 , n48031 , n48032 );
buf ( n48034 , n2220 );
buf ( n48035 , n48034 );
nand ( n2223 , n2209 , n48035 );
buf ( n48037 , n2223 );
buf ( n48038 , n48037 );
or ( n2226 , n48017 , n48038 );
xor ( n2227 , n46534 , n46668 );
and ( n2228 , n2227 , n46719 );
and ( n2229 , n46534 , n46668 );
or ( n2230 , n2228 , n2229 );
buf ( n48044 , n2230 );
buf ( n48045 , n48044 );
nand ( n2233 , n2226 , n48045 );
buf ( n48047 , n2233 );
buf ( n48048 , n48047 );
buf ( n48049 , n48037 );
buf ( n48050 , n2203 );
nand ( n2238 , n48049 , n48050 );
buf ( n48052 , n2238 );
buf ( n48053 , n48052 );
nand ( n48054 , n48048 , n48053 );
buf ( n48055 , n48054 );
buf ( n48056 , n48055 );
not ( n2244 , n48056 );
buf ( n48058 , n2244 );
not ( n2246 , n48058 );
or ( n2247 , n2201 , n2246 );
not ( n2248 , n2200 );
nand ( n2249 , n48055 , n2248 );
nand ( n2250 , n2247 , n2249 );
buf ( n48064 , n416 );
not ( n2252 , n48064 );
buf ( n48066 , n415 );
not ( n2254 , n48066 );
buf ( n48068 , n418 );
not ( n2256 , n48068 );
buf ( n48070 , n46055 );
buf ( n48071 , n46038 );
buf ( n48072 , n46078 );
not ( n2260 , n48072 );
buf ( n48074 , n46071 );
nor ( n2262 , n2260 , n48074 );
buf ( n48076 , n2262 );
buf ( n48077 , n48076 );
nand ( n2265 , n48070 , n48071 , n48077 );
buf ( n48079 , n2265 );
buf ( n48080 , n48079 );
not ( n2268 , n48080 );
or ( n2269 , n2256 , n2268 );
buf ( n48083 , n46055 );
buf ( n48084 , n46084 );
buf ( n48085 , n46038 );
nand ( n48086 , n48083 , n48084 , n48085 );
buf ( n48087 , n48086 );
buf ( n48088 , n48087 );
nand ( n2276 , n2269 , n48088 );
buf ( n48090 , n2276 );
buf ( n48091 , n48090 );
not ( n2279 , n48091 );
buf ( n48093 , n2279 );
buf ( n48094 , n48093 );
not ( n2282 , n48094 );
or ( n2283 , n2254 , n2282 );
buf ( n48097 , n48090 );
buf ( n48098 , n46124 );
nand ( n2286 , n48097 , n48098 );
buf ( n48100 , n2286 );
buf ( n48101 , n48100 );
nand ( n2289 , n2283 , n48101 );
buf ( n48103 , n2289 );
buf ( n48104 , n48103 );
not ( n2292 , n48104 );
or ( n2293 , n2252 , n2292 );
buf ( n48107 , n2217 );
buf ( n48108 , n46112 );
nand ( n2296 , n48107 , n48108 );
buf ( n48110 , n2296 );
buf ( n48111 , n48110 );
nand ( n2299 , n2293 , n48111 );
buf ( n48113 , n2299 );
not ( n2301 , n2115 );
not ( n2302 , n2123 );
not ( n2303 , n2302 );
or ( n2304 , n2301 , n2303 );
nand ( n2305 , n2304 , n2162 );
or ( n48119 , n2302 , n2115 );
nand ( n48120 , n2305 , n48119 );
not ( n2308 , n47955 );
not ( n2309 , n2156 );
or ( n2310 , n2308 , n2309 );
nand ( n2311 , n2310 , n2161 );
not ( n2312 , n2156 );
nand ( n2313 , n2312 , n47954 );
nand ( n2314 , n2311 , n2313 );
buf ( n48128 , n47968 );
buf ( n48129 , n47959 );
or ( n2317 , n48128 , n48129 );
buf ( n48131 , n47963 );
nand ( n2319 , n2317 , n48131 );
buf ( n48133 , n2319 );
buf ( n48134 , n48133 );
buf ( n48135 , n47959 );
buf ( n48136 , n47968 );
nand ( n2324 , n48135 , n48136 );
buf ( n48138 , n2324 );
buf ( n48139 , n48138 );
nand ( n2327 , n48134 , n48139 );
buf ( n48141 , n2327 );
buf ( n48142 , n48141 );
nand ( n2330 , n370 , n382 );
buf ( n48144 , n2330 );
not ( n2332 , n48144 );
and ( n2333 , n373 , n379 );
buf ( n48147 , n2333 );
not ( n2335 , n48147 );
or ( n2336 , n2332 , n2335 );
buf ( n48150 , n2330 );
buf ( n48151 , n2333 );
or ( n48152 , n48150 , n48151 );
nand ( n48153 , n2336 , n48152 );
buf ( n48154 , n48153 );
buf ( n48155 , n48154 );
nand ( n2343 , n371 , n381 );
buf ( n48157 , n2343 );
xor ( n2345 , n48155 , n48157 );
buf ( n48159 , n2345 );
buf ( n48160 , n48159 );
xor ( n2348 , n48142 , n48160 );
buf ( n48162 , n372 );
buf ( n48163 , n380 );
nand ( n2351 , n48162 , n48163 );
buf ( n48165 , n2351 );
buf ( n48166 , n374 );
buf ( n48167 , n378 );
nand ( n2355 , n48166 , n48167 );
buf ( n48169 , n2355 );
xor ( n2357 , n48165 , n48169 );
or ( n2358 , n2082 , n2085 );
nand ( n2359 , n2358 , n2084 );
nand ( n2360 , n2088 , n2085 );
nand ( n2361 , n2359 , n2360 );
xor ( n2362 , n2357 , n2361 );
buf ( n48176 , n2362 );
xor ( n2364 , n2348 , n48176 );
buf ( n48178 , n2364 );
not ( n2366 , n48178 );
or ( n2367 , n2095 , n2104 );
nand ( n2368 , n2367 , n657 );
nand ( n2369 , n2368 , n2111 );
or ( n2370 , n2314 , n2366 , n2369 );
nand ( n2371 , n2366 , n2369 );
or ( n48185 , n2371 , n2314 );
nand ( n48186 , n2370 , n48185 );
not ( n2374 , n48186 );
not ( n2375 , n2369 );
nand ( n2376 , n2375 , n2366 );
not ( n2377 , n2376 );
and ( n2378 , n2377 , n2314 );
and ( n2379 , n48178 , n2369 );
and ( n2380 , n2379 , n2314 );
nor ( n2381 , n2378 , n2380 );
nand ( n2382 , n2374 , n2381 );
xor ( n2383 , n48120 , n2382 );
not ( n2384 , n2383 );
not ( n2385 , n2384 );
buf ( n48199 , n411 );
buf ( n48200 , n1094 );
xor ( n2388 , n48199 , n48200 );
buf ( n48202 , n2388 );
not ( n2390 , n48202 );
not ( n2391 , n2390 );
not ( n2392 , n45497 );
and ( n2393 , n2391 , n2392 );
not ( n2394 , n411 );
not ( n2395 , n1150 );
or ( n2396 , n2394 , n2395 );
nand ( n2397 , n1139 , n46852 );
nand ( n2398 , n2396 , n2397 );
and ( n2399 , n2398 , n857 );
nor ( n2400 , n2393 , n2399 );
not ( n2401 , n2400 );
not ( n2402 , n2401 );
or ( n2403 , n2385 , n2402 );
nand ( n2404 , n2400 , n2383 );
nand ( n48218 , n2403 , n2404 );
xor ( n48219 , n48113 , n48218 );
buf ( n48220 , n45494 );
not ( n2408 , n48220 );
buf ( n48222 , n882 );
not ( n2410 , n48222 );
or ( n2411 , n2408 , n2410 );
buf ( n48225 , n48202 );
buf ( n48226 , n857 );
nand ( n2414 , n48225 , n48226 );
buf ( n48228 , n2414 );
buf ( n48229 , n48228 );
nand ( n2417 , n2411 , n48229 );
buf ( n48231 , n2417 );
not ( n2419 , n48231 );
xor ( n2420 , n46405 , n46485 );
and ( n2421 , n2420 , n46531 );
and ( n2422 , n46405 , n46485 );
or ( n2423 , n2421 , n2422 );
buf ( n48237 , n2423 );
not ( n2425 , n48237 );
nand ( n2426 , n2419 , n2425 );
not ( n2427 , n2426 );
not ( n2428 , n1104 );
not ( n2429 , n2066 );
or ( n2430 , n2428 , n2429 );
nand ( n2431 , n1214 , n46177 );
nand ( n2432 , n2430 , n2431 );
not ( n2433 , n2432 );
or ( n2434 , n2427 , n2433 );
nand ( n2435 , n48237 , n48231 );
nand ( n2436 , n2434 , n2435 );
xor ( n2437 , n48219 , n2436 );
not ( n48251 , n2437 );
and ( n48252 , n2250 , n48251 );
not ( n2440 , n2250 );
and ( n2441 , n2440 , n2437 );
nor ( n2442 , n48252 , n2441 );
not ( n2443 , n1221 );
not ( n2444 , n1295 );
or ( n2445 , n2443 , n2444 );
not ( n2446 , n1266 );
not ( n2447 , n1265 );
or ( n2448 , n2446 , n2447 );
or ( n2449 , n1295 , n1221 );
nand ( n2450 , n2448 , n2449 );
nand ( n2451 , n2445 , n2450 );
not ( n2452 , n2451 );
xor ( n2453 , n2425 , n48231 );
xnor ( n2454 , n2453 , n2432 );
buf ( n2455 , n2454 );
not ( n2456 , n2455 );
or ( n2457 , n2452 , n2456 );
or ( n2458 , n2455 , n2451 );
xor ( n2459 , n2203 , n48037 );
xor ( n2460 , n2459 , n48044 );
nand ( n2461 , n2458 , n2460 );
nand ( n2462 , n2457 , n2461 );
not ( n2463 , n2462 );
nand ( n2464 , n2442 , n2463 );
buf ( n48278 , n2464 );
not ( n2466 , n48278 );
xor ( n2467 , n2454 , n2451 );
xnor ( n2468 , n2467 , n2460 );
not ( n2469 , n2468 );
buf ( n48283 , n47018 );
not ( n48284 , n48283 );
buf ( n48285 , n46721 );
nor ( n2473 , n48284 , n48285 );
buf ( n48287 , n2473 );
buf ( n48288 , n48287 );
buf ( n48289 , n47111 );
or ( n2477 , n48288 , n48289 );
buf ( n48291 , n47018 );
not ( n2479 , n48291 );
buf ( n48293 , n46721 );
nand ( n2481 , n2479 , n48293 );
buf ( n48295 , n2481 );
buf ( n48296 , n48295 );
nand ( n2484 , n2477 , n48296 );
buf ( n48298 , n2484 );
nor ( n2486 , n2469 , n48298 );
buf ( n48300 , n2486 );
nor ( n2488 , n2466 , n48300 );
buf ( n48302 , n2488 );
buf ( n48303 , n48302 );
not ( n2491 , n45494 );
not ( n2492 , n2398 );
or ( n2493 , n2491 , n2492 );
xor ( n2494 , n1171 , n411 );
xnor ( n2495 , n2494 , n1170 );
nand ( n2496 , n857 , n2495 );
nand ( n2497 , n2493 , n2496 );
buf ( n48311 , n2497 );
buf ( n48312 , n46112 );
not ( n2500 , n48312 );
buf ( n48314 , n48103 );
not ( n2502 , n48314 );
or ( n2503 , n2500 , n2502 );
buf ( n48317 , n46134 );
buf ( n48318 , n48317 );
nand ( n2506 , n2503 , n48318 );
buf ( n48320 , n2506 );
buf ( n48321 , n48320 );
xor ( n2509 , n48311 , n48321 );
buf ( n48323 , n1104 );
not ( n2511 , n48323 );
not ( n2512 , n2210 );
not ( n2513 , n46153 );
and ( n2514 , n2512 , n2513 );
not ( n2515 , n2512 );
not ( n2516 , n413 );
and ( n2517 , n2515 , n2516 );
or ( n2518 , n2514 , n2517 );
and ( n2519 , n2216 , n2518 );
not ( n2520 , n2216 );
not ( n2521 , n46153 );
and ( n2522 , n2210 , n2521 );
not ( n2523 , n2210 );
not ( n2524 , n413 );
and ( n2525 , n2523 , n2524 );
or ( n2526 , n2522 , n2525 );
and ( n2527 , n2520 , n2526 );
or ( n2528 , n2519 , n2527 );
buf ( n48342 , n2528 );
not ( n2530 , n48342 );
or ( n2531 , n2511 , n2530 );
nand ( n2532 , n2073 , n46177 );
buf ( n48346 , n2532 );
nand ( n2534 , n2531 , n48346 );
buf ( n48348 , n2534 );
buf ( n48349 , n48348 );
not ( n48350 , n48349 );
buf ( n48351 , n48350 );
buf ( n48352 , n48351 );
xnor ( n2540 , n2509 , n48352 );
buf ( n48354 , n2540 );
buf ( n48355 , n48354 );
xor ( n2543 , n48113 , n48218 );
and ( n2544 , n2543 , n2436 );
and ( n2545 , n48113 , n48218 );
or ( n2546 , n2544 , n2545 );
buf ( n48360 , n2546 );
xor ( n2548 , n48355 , n48360 );
buf ( n48362 , n46196 );
not ( n2550 , n48362 );
buf ( n48364 , n875 );
not ( n2552 , n48364 );
or ( n2553 , n2550 , n2552 );
buf ( n48367 , n47274 );
not ( n2555 , n48367 );
buf ( n48369 , n2555 );
buf ( n48370 , n48369 );
buf ( n48371 , n46185 );
nand ( n2559 , n48370 , n48371 );
buf ( n48373 , n2559 );
buf ( n48374 , n48373 );
nand ( n2562 , n2553 , n48374 );
buf ( n48376 , n2562 );
xor ( n2564 , n48165 , n48169 );
and ( n2565 , n2564 , n2361 );
and ( n2566 , n48165 , n48169 );
or ( n2567 , n2565 , n2566 );
nand ( n2568 , n371 , n380 );
nand ( n48382 , n370 , n382 );
not ( n48383 , n48382 );
not ( n2571 , n2343 );
or ( n2572 , n48383 , n2571 );
or ( n2573 , n2343 , n48382 );
nand ( n2574 , n2573 , n655 );
nand ( n2575 , n2572 , n2574 );
xor ( n2576 , n2568 , n2575 );
nand ( n2577 , n372 , n379 );
nand ( n2578 , n373 , n378 );
xor ( n2579 , n2577 , n2578 );
nand ( n2580 , n370 , n381 );
xor ( n2581 , n2579 , n2580 );
xor ( n2582 , n2576 , n2581 );
buf ( n48396 , n2582 );
not ( n2584 , n48396 );
buf ( n48398 , n2584 );
and ( n2586 , n2567 , n48398 );
not ( n2587 , n2567 );
and ( n2588 , n2587 , n2582 );
or ( n2589 , n2586 , n2588 );
buf ( n48403 , n2589 );
xor ( n2591 , n48142 , n48160 );
and ( n2592 , n2591 , n48176 );
and ( n2593 , n48142 , n48160 );
or ( n2594 , n2592 , n2593 );
buf ( n48408 , n2594 );
buf ( n48409 , n48408 );
xnor ( n2597 , n48403 , n48409 );
buf ( n48411 , n2597 );
not ( n2599 , n2314 );
not ( n2600 , n2376 );
or ( n2601 , n2599 , n2600 );
not ( n48415 , n2379 );
nand ( n48416 , n2601 , n48415 );
xnor ( n2604 , n48411 , n48416 );
xnor ( n2605 , n48376 , n2604 );
buf ( n48419 , n2605 );
or ( n2607 , n48120 , n2382 );
not ( n2608 , n2607 );
not ( n2609 , n2401 );
or ( n2610 , n2608 , n2609 );
nand ( n2611 , n48120 , n2382 );
nand ( n2612 , n2610 , n2611 );
buf ( n48426 , n2612 );
xor ( n2614 , n48419 , n48426 );
or ( n2615 , n2191 , n47888 );
nand ( n2616 , n2615 , n2182 );
buf ( n48430 , n2616 );
nand ( n2618 , n2191 , n47888 );
buf ( n48432 , n2618 );
nand ( n2620 , n48430 , n48432 );
buf ( n48434 , n2620 );
buf ( n48435 , n48434 );
xnor ( n2623 , n2614 , n48435 );
buf ( n48437 , n2623 );
buf ( n48438 , n48437 );
xnor ( n2626 , n2548 , n48438 );
buf ( n48440 , n2626 );
buf ( n48441 , n48440 );
not ( n2629 , n2248 );
not ( n2630 , n48251 );
or ( n2631 , n2629 , n2630 );
buf ( n48445 , n48055 );
buf ( n2633 , n48445 );
buf ( n48447 , n2633 );
nand ( n48448 , n2631 , n48447 );
buf ( n48449 , n48448 );
nand ( n2637 , n2437 , n2200 );
buf ( n48451 , n2637 );
nand ( n2639 , n48449 , n48451 );
buf ( n48453 , n2639 );
not ( n2641 , n48453 );
buf ( n48455 , n2641 );
nand ( n2643 , n48441 , n48455 );
buf ( n48457 , n2643 );
buf ( n48458 , n48457 );
and ( n2646 , n48303 , n48458 );
buf ( n48460 , n2646 );
not ( n2648 , n48460 );
or ( n2649 , n2057 , n2648 );
buf ( n48463 , n2442 );
not ( n2651 , n48463 );
buf ( n48465 , n2462 );
nand ( n2653 , n2651 , n48465 );
buf ( n48467 , n2653 );
buf ( n48468 , n48467 );
not ( n2656 , n48468 );
not ( n2657 , n48298 );
nor ( n2658 , n2468 , n2657 );
buf ( n48472 , n2658 );
buf ( n48473 , n2464 );
nand ( n2661 , n48472 , n48473 );
buf ( n48475 , n2661 );
buf ( n48476 , n48475 );
not ( n2664 , n48476 );
or ( n2665 , n2656 , n2664 );
buf ( n48479 , n48453 );
not ( n2667 , n48479 );
buf ( n48481 , n48440 );
nand ( n48482 , n2667 , n48481 );
buf ( n48483 , n48482 );
buf ( n48484 , n48483 );
nand ( n2672 , n2665 , n48484 );
buf ( n48486 , n2672 );
buf ( n48487 , n48486 );
not ( n2675 , n48440 );
buf ( n2676 , n48453 );
nand ( n2677 , n2675 , n2676 );
buf ( n48491 , n2677 );
nand ( n2679 , n48487 , n48491 );
buf ( n48493 , n2679 );
buf ( n48494 , n48493 );
not ( n2682 , n48494 );
buf ( n48496 , n2682 );
nand ( n2684 , n2649 , n48496 );
buf ( n48498 , n371 );
buf ( n48499 , n379 );
nand ( n2687 , n48498 , n48499 );
buf ( n48501 , n2687 );
buf ( n48502 , n370 );
buf ( n48503 , n380 );
nand ( n2691 , n48502 , n48503 );
buf ( n48505 , n2691 );
xor ( n2693 , n48501 , n48505 );
buf ( n48507 , n372 );
buf ( n48508 , n378 );
nand ( n2696 , n48507 , n48508 );
buf ( n48510 , n2696 );
xor ( n2698 , n2693 , n48510 );
xor ( n2699 , n2577 , n2578 );
and ( n2700 , n2699 , n2580 );
and ( n2701 , n2577 , n2578 );
or ( n2702 , n2700 , n2701 );
xor ( n48516 , n2568 , n2575 );
and ( n48517 , n48516 , n2581 );
and ( n2705 , n2568 , n2575 );
or ( n2706 , n48517 , n2705 );
xor ( n2707 , n2702 , n2706 );
xor ( n2708 , n2698 , n2707 );
not ( n2709 , n2708 );
not ( n2710 , n46955 );
nand ( n2711 , n2710 , n46185 );
not ( n2712 , n47274 );
nand ( n48526 , n2712 , n46196 );
nand ( n2714 , n2711 , n48526 );
not ( n2715 , n2714 );
or ( n48529 , n2709 , n2715 );
not ( n2717 , n2708 );
and ( n2718 , n48526 , n2717 );
not ( n2719 , n2718 );
not ( n2720 , n2711 );
or ( n2721 , n2719 , n2720 );
not ( n48535 , n2567 );
not ( n2723 , n2582 );
or ( n48537 , n48535 , n2723 );
buf ( n48538 , n48408 );
buf ( n48539 , n2567 );
not ( n2727 , n48539 );
buf ( n48541 , n48398 );
nand ( n48542 , n2727 , n48541 );
buf ( n48543 , n48542 );
buf ( n48544 , n48543 );
nand ( n48545 , n48538 , n48544 );
buf ( n48546 , n48545 );
nand ( n2734 , n48537 , n48546 );
nand ( n2735 , n2721 , n2734 );
nand ( n2736 , n48529 , n2735 );
buf ( n48550 , n2736 );
buf ( n48551 , n857 );
not ( n2739 , n48551 );
xor ( n2740 , n2512 , n2216 );
xor ( n2741 , n2740 , n411 );
buf ( n48555 , n2741 );
not ( n2743 , n48555 );
or ( n2744 , n2739 , n2743 );
not ( n2745 , n411 );
buf ( n48559 , n47102 );
not ( n2747 , n48559 );
buf ( n48561 , n2747 );
not ( n2749 , n48561 );
or ( n2750 , n2745 , n2749 );
buf ( n48564 , n411 );
not ( n2752 , n48564 );
buf ( n48566 , n47102 );
nand ( n2754 , n2752 , n48566 );
buf ( n48568 , n2754 );
nand ( n2756 , n2750 , n48568 );
buf ( n48570 , n2756 );
buf ( n48571 , n45494 );
nand ( n2759 , n48570 , n48571 );
buf ( n48573 , n2759 );
buf ( n48574 , n48573 );
nand ( n2762 , n2744 , n48574 );
buf ( n48576 , n2762 );
buf ( n48577 , n48576 );
xor ( n2765 , n48550 , n48577 );
not ( n2766 , n857 );
not ( n2767 , n2756 );
or ( n2768 , n2766 , n2767 );
nand ( n2769 , n2495 , n45494 );
nand ( n2770 , n2768 , n2769 );
not ( n2771 , n2770 );
not ( n2772 , n46135 );
and ( n2773 , n48090 , n46153 );
not ( n2774 , n48090 );
and ( n2775 , n2774 , n413 );
or ( n2776 , n2773 , n2775 );
nand ( n2777 , n2776 , n1104 );
buf ( n48591 , n2528 );
buf ( n48592 , n46177 );
nand ( n2780 , n48591 , n48592 );
buf ( n48594 , n2780 );
nand ( n2782 , n2772 , n2777 , n48594 );
not ( n2783 , n2782 );
or ( n48597 , n2771 , n2783 );
buf ( n48598 , n46231 );
nand ( n2786 , n2777 , n48594 );
buf ( n48600 , n2786 );
nand ( n2788 , n48598 , n48600 );
buf ( n48602 , n2788 );
nand ( n2790 , n48597 , n48602 );
buf ( n48604 , n2790 );
xor ( n2792 , n2765 , n48604 );
buf ( n48606 , n2792 );
not ( n2794 , n2734 );
not ( n2795 , n2708 );
and ( n2796 , n2794 , n2795 );
and ( n2797 , n2734 , n2708 );
nor ( n2798 , n2796 , n2797 );
not ( n2799 , n2798 );
not ( n48613 , n2714 );
or ( n2801 , n2799 , n48613 );
or ( n2802 , n2714 , n2798 );
nand ( n2803 , n2801 , n2802 );
buf ( n48617 , n2803 );
buf ( n48618 , n48411 );
not ( n2806 , n48618 );
buf ( n48620 , n2806 );
buf ( n48621 , n48620 );
not ( n48622 , n48621 );
buf ( n48623 , n48376 );
not ( n2811 , n48623 );
or ( n2812 , n48622 , n2811 );
buf ( n48626 , n48376 );
buf ( n48627 , n48620 );
or ( n2815 , n48626 , n48627 );
buf ( n48629 , n48416 );
nand ( n2817 , n2815 , n48629 );
buf ( n48631 , n2817 );
buf ( n48632 , n48631 );
nand ( n2820 , n2812 , n48632 );
buf ( n48634 , n2820 );
buf ( n48635 , n48634 );
not ( n48636 , n48635 );
buf ( n48637 , n48636 );
buf ( n48638 , n48637 );
xor ( n2826 , n48617 , n48638 );
not ( n2827 , n48351 );
buf ( n48641 , n48320 );
not ( n2829 , n48641 );
buf ( n48643 , n2829 );
not ( n2831 , n48643 );
and ( n2832 , n2827 , n2831 );
buf ( n48646 , n48351 );
buf ( n48647 , n48643 );
nand ( n2835 , n48646 , n48647 );
buf ( n48649 , n2835 );
and ( n2837 , n48649 , n2497 );
nor ( n2838 , n2832 , n2837 );
buf ( n48652 , n2838 );
and ( n2840 , n2826 , n48652 );
and ( n2841 , n48617 , n48638 );
or ( n2842 , n2840 , n2841 );
buf ( n48656 , n2842 );
xor ( n2844 , n48606 , n48656 );
buf ( n48658 , n46955 );
not ( n2846 , n48658 );
buf ( n48660 , n46196 );
not ( n2848 , n48660 );
buf ( n48662 , n2848 );
buf ( n48663 , n48662 );
not ( n2851 , n48663 );
and ( n2852 , n2846 , n2851 );
buf ( n48666 , n46992 );
not ( n2854 , n48666 );
buf ( n48668 , n2854 );
buf ( n48669 , n48668 );
buf ( n48670 , n46185 );
and ( n2858 , n48669 , n48670 );
nor ( n2859 , n2852 , n2858 );
buf ( n48673 , n2859 );
buf ( n48674 , n48673 );
buf ( n48675 , n46177 );
not ( n2863 , n48675 );
buf ( n48677 , n2776 );
not ( n2865 , n48677 );
or ( n2866 , n2863 , n2865 );
nand ( n2867 , n46157 , n1104 );
buf ( n48681 , n2867 );
nand ( n2869 , n2866 , n48681 );
buf ( n48683 , n2869 );
buf ( n48684 , n48683 );
not ( n48685 , n48684 );
buf ( n48686 , n48685 );
buf ( n48687 , n48686 );
xor ( n2875 , n48674 , n48687 );
buf ( n48689 , n371 );
buf ( n48690 , n378 );
nand ( n2878 , n48689 , n48690 );
buf ( n48692 , n2878 );
buf ( n48693 , n370 );
buf ( n48694 , n379 );
nand ( n2882 , n48693 , n48694 );
buf ( n48696 , n2882 );
xor ( n2884 , n48692 , n48696 );
xor ( n2885 , n48501 , n48505 );
and ( n2886 , n2885 , n48510 );
and ( n2887 , n48501 , n48505 );
or ( n2888 , n2886 , n2887 );
xor ( n2889 , n2884 , n2888 );
xor ( n2890 , n48501 , n48505 );
xor ( n2891 , n2890 , n48510 );
and ( n2892 , n2702 , n2891 );
xor ( n2893 , n48501 , n48505 );
xor ( n2894 , n2893 , n48510 );
and ( n2895 , n2706 , n2894 );
and ( n2896 , n2702 , n2706 );
or ( n2897 , n2892 , n2895 , n2896 );
xor ( n2898 , n2897 , n46141 );
xor ( n2899 , n2889 , n2898 );
buf ( n48713 , n2899 );
xnor ( n2901 , n2875 , n48713 );
buf ( n48715 , n2901 );
buf ( n48716 , n48715 );
not ( n2904 , n48716 );
buf ( n48718 , n2904 );
and ( n2906 , n2844 , n48718 );
not ( n2907 , n2844 );
and ( n2908 , n2907 , n48715 );
nor ( n2909 , n2906 , n2908 );
buf ( n48723 , n2909 );
xor ( n2911 , n48617 , n48638 );
xor ( n2912 , n2911 , n48652 );
buf ( n48726 , n2912 );
not ( n2914 , n48726 );
xor ( n2915 , n2770 , n2786 );
not ( n2916 , n46231 );
and ( n2917 , n2915 , n2916 );
not ( n2918 , n2915 );
and ( n2919 , n2918 , n46231 );
nor ( n2920 , n2917 , n2919 );
not ( n2921 , n2920 );
and ( n2922 , n2914 , n2921 );
nand ( n2923 , n48726 , n2920 );
not ( n2924 , n2612 );
nand ( n2925 , n2924 , n2605 );
not ( n2926 , n2925 );
not ( n2927 , n48434 );
or ( n2928 , n2926 , n2927 );
buf ( n48742 , n2605 );
not ( n2930 , n48742 );
buf ( n48744 , n2612 );
nand ( n2932 , n2930 , n48744 );
buf ( n48746 , n2932 );
nand ( n2934 , n2928 , n48746 );
and ( n2935 , n2923 , n2934 );
nor ( n2936 , n2922 , n2935 );
buf ( n48750 , n2936 );
nand ( n2938 , n48723 , n48750 );
buf ( n48752 , n2938 );
buf ( n48753 , n48752 );
not ( n2941 , n2920 );
not ( n2942 , n2941 );
not ( n2943 , n2934 );
not ( n2944 , n2943 );
or ( n2945 , n2942 , n2944 );
nand ( n2946 , n2920 , n2934 );
nand ( n2947 , n2945 , n2946 );
not ( n2948 , n48726 );
and ( n2949 , n2947 , n2948 );
not ( n2950 , n2947 );
and ( n2951 , n2950 , n48726 );
nor ( n2952 , n2949 , n2951 );
buf ( n48766 , n2952 );
not ( n2954 , n48766 );
buf ( n48768 , n2954 );
buf ( n48769 , n48768 );
buf ( n48770 , n48354 );
not ( n2958 , n48770 );
buf ( n48772 , n2958 );
buf ( n48773 , n48772 );
not ( n2961 , n48773 );
buf ( n48775 , n48437 );
not ( n2963 , n48775 );
buf ( n48777 , n2963 );
buf ( n48778 , n48777 );
not ( n2966 , n48778 );
or ( n2967 , n2961 , n2966 );
buf ( n48781 , n2546 );
nand ( n2969 , n2967 , n48781 );
buf ( n48783 , n2969 );
buf ( n48784 , n48783 );
buf ( n48785 , n48777 );
buf ( n48786 , n48772 );
or ( n2974 , n48785 , n48786 );
buf ( n48788 , n2974 );
buf ( n48789 , n48788 );
nand ( n2977 , n48784 , n48789 );
buf ( n48791 , n2977 );
buf ( n48792 , n48791 );
not ( n2980 , n48792 );
buf ( n48794 , n2980 );
buf ( n48795 , n48794 );
nand ( n2983 , n48769 , n48795 );
buf ( n48797 , n2983 );
buf ( n48798 , n48797 );
and ( n2986 , n48753 , n48798 );
buf ( n48800 , n2986 );
xor ( n2988 , n48550 , n48577 );
and ( n2989 , n2988 , n48604 );
and ( n2990 , n48550 , n48577 );
or ( n2991 , n2989 , n2990 );
buf ( n48805 , n2991 );
buf ( n48806 , n48686 );
buf ( n48807 , n48673 );
nand ( n2995 , n48806 , n48807 );
buf ( n48809 , n2995 );
buf ( n48810 , n48809 );
not ( n2998 , n48810 );
buf ( n48812 , n2899 );
not ( n3000 , n48812 );
or ( n3001 , n2998 , n3000 );
buf ( n48815 , n48673 );
not ( n3003 , n48815 );
buf ( n48817 , n48683 );
nand ( n3005 , n3003 , n48817 );
buf ( n48819 , n3005 );
buf ( n48820 , n48819 );
nand ( n3008 , n3001 , n48820 );
buf ( n48822 , n3008 );
buf ( n48823 , n48822 );
not ( n3011 , n48823 );
buf ( n48825 , n3011 );
xor ( n3013 , n48805 , n48825 );
xor ( n3014 , n48692 , n48696 );
xor ( n3015 , n3014 , n2888 );
and ( n3016 , n2897 , n3015 );
xor ( n3017 , n48692 , n48696 );
xor ( n3018 , n3017 , n2888 );
and ( n3019 , n46141 , n3018 );
and ( n3020 , n2897 , n46141 );
or ( n3021 , n3016 , n3019 , n3020 );
xor ( n3022 , n46217 , n3021 );
buf ( n48836 , n370 );
buf ( n48837 , n378 );
nand ( n3025 , n48836 , n48837 );
buf ( n48839 , n3025 );
buf ( n48840 , n48839 );
xor ( n3028 , n48692 , n48696 );
and ( n3029 , n3028 , n2888 );
and ( n3030 , n48692 , n48696 );
or ( n3031 , n3029 , n3030 );
buf ( n48845 , n3031 );
xor ( n3033 , n48840 , n48845 );
buf ( n48847 , n46141 );
xor ( n3035 , n3033 , n48847 );
buf ( n48849 , n3035 );
xor ( n3037 , n3022 , n48849 );
buf ( n48851 , n46185 );
not ( n3039 , n48851 );
buf ( n48853 , n48561 );
not ( n3041 , n48853 );
buf ( n48855 , n3041 );
buf ( n48856 , n48855 );
not ( n3044 , n48856 );
or ( n3045 , n3039 , n3044 );
buf ( n48859 , n48668 );
buf ( n48860 , n46196 );
nand ( n3048 , n48859 , n48860 );
buf ( n48862 , n3048 );
buf ( n48863 , n48862 );
nand ( n3051 , n3045 , n48863 );
buf ( n48865 , n3051 );
buf ( n48866 , n48865 );
not ( n3054 , n48866 );
buf ( n48868 , n857 );
not ( n3056 , n48868 );
and ( n3057 , n411 , n48093 );
not ( n3058 , n411 );
buf ( n48872 , n48093 );
not ( n3060 , n48872 );
buf ( n48874 , n3060 );
and ( n3062 , n3058 , n48874 );
or ( n3063 , n3057 , n3062 );
buf ( n48877 , n3063 );
not ( n3065 , n48877 );
or ( n3066 , n3056 , n3065 );
buf ( n48880 , n2741 );
buf ( n48881 , n45494 );
nand ( n3069 , n48880 , n48881 );
buf ( n48883 , n3069 );
buf ( n48884 , n48883 );
nand ( n3072 , n3066 , n48884 );
buf ( n48886 , n3072 );
buf ( n48887 , n48886 );
not ( n3075 , n48887 );
buf ( n48889 , n3075 );
buf ( n48890 , n48889 );
not ( n3078 , n48890 );
or ( n3079 , n3054 , n3078 );
buf ( n48893 , n48889 );
buf ( n48894 , n48865 );
or ( n3082 , n48893 , n48894 );
nand ( n3083 , n3079 , n3082 );
buf ( n48897 , n3083 );
xor ( n3085 , n3037 , n48897 );
xnor ( n3086 , n3013 , n3085 );
not ( n3087 , n3086 );
buf ( n48901 , n48606 );
not ( n3089 , n48901 );
buf ( n48903 , n3089 );
buf ( n48904 , n48903 );
not ( n3092 , n48904 );
buf ( n48906 , n48715 );
not ( n3094 , n48906 );
or ( n3095 , n3092 , n3094 );
buf ( n48909 , n48656 );
not ( n3097 , n48909 );
buf ( n48911 , n3097 );
buf ( n48912 , n48911 );
nand ( n3100 , n3095 , n48912 );
buf ( n48914 , n3100 );
buf ( n48915 , n48914 );
buf ( n48916 , n48903 );
not ( n3104 , n48916 );
buf ( n48918 , n48718 );
nand ( n3106 , n3104 , n48918 );
buf ( n48920 , n3106 );
buf ( n48921 , n48920 );
nand ( n3109 , n48915 , n48921 );
buf ( n48923 , n3109 );
buf ( n48924 , n48923 );
not ( n3112 , n48924 );
buf ( n48926 , n3112 );
nand ( n3114 , n3087 , n48926 );
xor ( n3115 , n46217 , n3021 );
and ( n3116 , n3115 , n48849 );
and ( n3117 , n46217 , n3021 );
or ( n3118 , n3116 , n3117 );
buf ( n48932 , n48865 );
not ( n3120 , n48932 );
buf ( n48934 , n48889 );
nand ( n3122 , n3120 , n48934 );
buf ( n48936 , n3122 );
not ( n3124 , n48936 );
not ( n3125 , n3037 );
or ( n3126 , n3124 , n3125 );
buf ( n48940 , n48886 );
buf ( n48941 , n48865 );
nand ( n3129 , n48940 , n48941 );
buf ( n48943 , n3129 );
nand ( n3131 , n3126 , n48943 );
xor ( n3132 , n3118 , n3131 );
buf ( n48946 , n46141 );
not ( n48947 , n48946 );
buf ( n48948 , n48947 );
xor ( n3136 , n46214 , n48948 );
buf ( n48950 , n3136 );
xor ( n3138 , n48840 , n48845 );
and ( n3139 , n3138 , n48847 );
and ( n3140 , n48840 , n48845 );
or ( n3141 , n3139 , n3140 );
buf ( n48955 , n3141 );
buf ( n48956 , n48955 );
xor ( n3144 , n48950 , n48956 );
buf ( n48958 , n3144 );
buf ( n48959 , n48958 );
not ( n3147 , n48959 );
buf ( n48961 , n3147 );
not ( n48962 , n48961 );
buf ( n48963 , n45494 );
not ( n3151 , n48963 );
buf ( n48965 , n3063 );
not ( n48966 , n48965 );
or ( n48967 , n3151 , n48966 );
nand ( n3155 , n46101 , n857 );
buf ( n48969 , n3155 );
nand ( n3157 , n48967 , n48969 );
buf ( n48971 , n3157 );
buf ( n48972 , n48971 );
not ( n3160 , n48972 );
buf ( n48974 , n46196 );
not ( n3162 , n48974 );
buf ( n48976 , n48855 );
not ( n3164 , n48976 );
or ( n3165 , n3162 , n3164 );
buf ( n48979 , n2740 );
buf ( n48980 , n46185 );
nand ( n3168 , n48979 , n48980 );
buf ( n48982 , n3168 );
buf ( n48983 , n48982 );
nand ( n3171 , n3165 , n48983 );
buf ( n48985 , n3171 );
buf ( n48986 , n48985 );
not ( n3174 , n48986 );
buf ( n48988 , n3174 );
buf ( n48989 , n48988 );
not ( n3177 , n48989 );
and ( n3178 , n3160 , n3177 );
buf ( n48992 , n48971 );
buf ( n48993 , n48988 );
and ( n3181 , n48992 , n48993 );
nor ( n3182 , n3178 , n3181 );
buf ( n48996 , n3182 );
buf ( n48997 , n48996 );
not ( n3185 , n48997 );
buf ( n48999 , n3185 );
not ( n3187 , n48999 );
or ( n3188 , n48962 , n3187 );
buf ( n49002 , n48958 );
buf ( n49003 , n48996 );
nand ( n3191 , n49002 , n49003 );
buf ( n49005 , n3191 );
nand ( n3193 , n3188 , n49005 );
xor ( n3194 , n3132 , n3193 );
not ( n3195 , n3194 );
buf ( n49009 , n48805 );
not ( n3197 , n49009 );
buf ( n49011 , n48825 );
nand ( n3199 , n3197 , n49011 );
buf ( n49013 , n3199 );
not ( n3201 , n49013 );
not ( n3202 , n3085 );
or ( n3203 , n3201 , n3202 );
buf ( n49017 , n48805 );
buf ( n49018 , n48822 );
nand ( n3206 , n49017 , n49018 );
buf ( n49020 , n3206 );
nand ( n3208 , n3203 , n49020 );
not ( n3209 , n3208 );
nand ( n3210 , n3195 , n3209 );
and ( n3211 , n2684 , n48800 , n3114 , n3210 );
buf ( n49025 , n48971 );
not ( n3213 , n49025 );
buf ( n49027 , n48988 );
nand ( n3215 , n3213 , n49027 );
buf ( n49029 , n3215 );
not ( n3217 , n49029 );
not ( n49031 , n48958 );
or ( n3219 , n3217 , n49031 );
buf ( n49033 , n48988 );
not ( n3221 , n49033 );
buf ( n49035 , n48971 );
nand ( n3223 , n3221 , n49035 );
buf ( n49037 , n3223 );
nand ( n3225 , n3219 , n49037 );
not ( n3226 , n3225 );
not ( n49040 , n3226 );
not ( n3228 , n49040 );
not ( n3229 , n46102 );
and ( n3230 , n46214 , n48948 );
buf ( n49044 , n3230 );
not ( n3232 , n49044 );
buf ( n49046 , n46231 );
buf ( n49047 , n46217 );
nand ( n3235 , n49046 , n49047 );
buf ( n49049 , n3235 );
buf ( n49050 , n49049 );
nand ( n3238 , n3232 , n49050 );
buf ( n49052 , n3238 );
xor ( n3240 , n3229 , n49052 );
not ( n3241 , n3230 );
buf ( n49055 , n3241 );
not ( n3243 , n49055 );
buf ( n49057 , n48955 );
not ( n3245 , n49057 );
or ( n3246 , n3243 , n3245 );
buf ( n49060 , n49049 );
nand ( n3248 , n3246 , n49060 );
buf ( n49062 , n3248 );
xnor ( n3250 , n3240 , n49062 );
not ( n3251 , n3250 );
not ( n3252 , n3251 );
or ( n3253 , n3228 , n3252 );
not ( n3254 , n3226 );
not ( n3255 , n3250 );
or ( n3256 , n3254 , n3255 );
not ( n3257 , n46185 );
not ( n3258 , n48874 );
or ( n3259 , n3257 , n3258 );
buf ( n49073 , n2740 );
buf ( n49074 , n46196 );
nand ( n3262 , n49073 , n49074 );
buf ( n49076 , n3262 );
nand ( n3264 , n3259 , n49076 );
nand ( n3265 , n3256 , n3264 );
nand ( n3266 , n3253 , n3265 );
or ( n3267 , n49062 , n46238 );
nand ( n3268 , n3267 , n49052 );
buf ( n49082 , n49062 );
buf ( n49083 , n46238 );
nand ( n3271 , n49082 , n49083 );
buf ( n49085 , n3271 );
nand ( n3273 , n3268 , n49085 );
not ( n3274 , n3273 );
buf ( n49088 , n46196 );
not ( n3276 , n49088 );
buf ( n49090 , n48874 );
not ( n3278 , n49090 );
or ( n3279 , n3276 , n3278 );
buf ( n49093 , n46188 );
nand ( n3281 , n3279 , n49093 );
buf ( n49095 , n3281 );
not ( n3283 , n49095 );
not ( n49097 , n3283 );
buf ( n49098 , n2916 );
buf ( n49099 , n3241 );
nand ( n3287 , n49098 , n49099 );
buf ( n49101 , n3287 );
not ( n3289 , n46214 );
not ( n3290 , n46144 );
or ( n3291 , n3289 , n3290 );
buf ( n49105 , n46207 );
buf ( n49106 , n46102 );
nand ( n3294 , n49105 , n49106 );
buf ( n49108 , n3294 );
nand ( n3296 , n3291 , n49108 );
buf ( n49110 , n3296 );
not ( n3298 , n49110 );
buf ( n49112 , n3298 );
xor ( n3300 , n49101 , n49112 );
not ( n3301 , n3300 );
or ( n3302 , n49097 , n3301 );
or ( n3303 , n3300 , n3283 );
nand ( n3304 , n3302 , n3303 );
not ( n3305 , n3304 );
or ( n3306 , n3274 , n3305 );
or ( n3307 , n3273 , n3304 );
nand ( n3308 , n3306 , n3307 );
nor ( n3309 , n3266 , n3308 );
not ( n3310 , n3309 );
not ( n3311 , n3273 );
buf ( n49125 , n49095 );
not ( n3313 , n49125 );
buf ( n49127 , n3300 );
nand ( n3315 , n3313 , n49127 );
buf ( n49129 , n3315 );
not ( n49130 , n49129 );
or ( n49131 , n3311 , n49130 );
buf ( n49132 , n3300 );
not ( n3320 , n49132 );
buf ( n49134 , n49095 );
nand ( n3322 , n3320 , n49134 );
buf ( n49136 , n3322 );
nand ( n3324 , n49131 , n49136 );
buf ( n49138 , n3324 );
not ( n3326 , n49138 );
not ( n49140 , n2916 );
buf ( n49141 , n46207 );
not ( n3329 , n49141 );
buf ( n49143 , n46102 );
nand ( n3331 , n3329 , n49143 );
buf ( n49145 , n3331 );
not ( n3333 , n49145 );
or ( n3334 , n49140 , n3333 );
buf ( n49148 , n49145 );
not ( n3336 , n49148 );
buf ( n49150 , n3336 );
nand ( n3338 , n46231 , n49150 );
nand ( n3339 , n3334 , n3338 );
not ( n3340 , n3296 );
and ( n3341 , n3339 , n3340 );
not ( n3342 , n3339 );
and ( n3343 , n3342 , n3296 );
nor ( n3344 , n3341 , n3343 );
buf ( n49158 , n3344 );
not ( n3346 , n49158 );
buf ( n49160 , n46199 );
not ( n3348 , n49160 );
and ( n3349 , n3346 , n3348 );
buf ( n49163 , n3344 );
buf ( n49164 , n46199 );
and ( n3352 , n49163 , n49164 );
nor ( n3353 , n3349 , n3352 );
buf ( n49167 , n3353 );
buf ( n49168 , n49167 );
buf ( n49169 , n2916 );
buf ( n49170 , n3296 );
nand ( n3358 , n49169 , n49170 );
buf ( n49172 , n3358 );
buf ( n49173 , n49172 );
buf ( n49174 , n3241 );
nand ( n49175 , n49173 , n49174 );
buf ( n49176 , n49175 );
buf ( n49177 , n49176 );
and ( n3365 , n49168 , n49177 );
not ( n3366 , n49168 );
buf ( n49180 , n49176 );
not ( n3368 , n49180 );
buf ( n49182 , n3368 );
buf ( n49183 , n49182 );
and ( n3371 , n3366 , n49183 );
nor ( n3372 , n3365 , n3371 );
buf ( n49186 , n3372 );
buf ( n49187 , n49186 );
not ( n3375 , n49187 );
buf ( n49189 , n3375 );
buf ( n49190 , n49189 );
nand ( n3378 , n3326 , n49190 );
buf ( n49192 , n3378 );
nand ( n3380 , n3310 , n49192 );
buf ( n49194 , n3380 );
not ( n3382 , n3193 );
not ( n3383 , n3118 );
or ( n3384 , n3382 , n3383 );
nor ( n3385 , n3193 , n3118 );
not ( n3386 , n3131 );
or ( n3387 , n3385 , n3386 );
nand ( n3388 , n3384 , n3387 );
xor ( n3389 , n3264 , n3225 );
xnor ( n3390 , n3389 , n3250 );
nor ( n3391 , n3388 , n3390 );
buf ( n49205 , n3391 );
buf ( n49206 , n46199 );
not ( n3395 , n49206 );
buf ( n49208 , n49176 );
not ( n3397 , n49208 );
or ( n3398 , n3395 , n3397 );
buf ( n49211 , n3344 );
nand ( n3400 , n3398 , n49211 );
buf ( n49213 , n3400 );
buf ( n49214 , n49213 );
buf ( n49215 , n49182 );
not ( n3404 , n46199 );
buf ( n49217 , n3404 );
nand ( n3406 , n49215 , n49217 );
buf ( n49219 , n3406 );
buf ( n49220 , n49219 );
nand ( n3409 , n49214 , n49220 );
buf ( n49222 , n3409 );
buf ( n49223 , n46223 );
and ( n3414 , n46148 , n49150 );
not ( n3415 , n46148 );
and ( n3416 , n3415 , n49145 );
or ( n3417 , n3414 , n3416 );
buf ( n49228 , n3417 );
xor ( n3419 , n49223 , n49228 );
not ( n3420 , n49172 );
not ( n3421 , n49145 );
or ( n3422 , n3420 , n3421 );
buf ( n49233 , n49112 );
buf ( n49234 , n46231 );
nand ( n3425 , n49233 , n49234 );
buf ( n49236 , n3425 );
nand ( n3427 , n3422 , n49236 );
buf ( n49238 , n3427 );
xor ( n3429 , n3419 , n49238 );
buf ( n49240 , n3429 );
buf ( n49241 , C1 );
buf ( n49242 , C0 );
buf ( n49243 , n49242 );
nand ( n3438 , n3417 , n46222 );
buf ( n49245 , n3438 );
buf ( n49246 , n46223 );
not ( n3441 , n49246 );
buf ( n49248 , n3417 );
not ( n3443 , n49248 );
buf ( n49250 , n3443 );
buf ( n49251 , n49250 );
not ( n3446 , n49251 );
or ( n3447 , n3441 , n3446 );
buf ( n49254 , n3427 );
nand ( n3449 , n3447 , n49254 );
buf ( n49256 , n3449 );
buf ( n49257 , n49256 );
nand ( n3452 , n49245 , n49257 );
buf ( n49259 , n3452 );
buf ( n49260 , n46231 );
buf ( n49261 , n46238 );
nor ( n3457 , n49260 , n49261 );
buf ( n49263 , n3457 );
or ( n3459 , n49263 , n49150 );
not ( n3460 , n3459 );
not ( n3461 , n46256 );
or ( n3462 , n3460 , n3461 );
buf ( n49268 , n46256 );
or ( n49269 , n49268 , n3459 );
nand ( n3465 , n3462 , n49269 );
buf ( n49271 , n46224 );
nor ( n3472 , n49263 , n49150 );
buf ( n49273 , n3472 );
nand ( n3474 , n49271 , n49273 );
buf ( n49275 , n3474 );
nand ( n3476 , n49275 , n46245 );
buf ( n49277 , C0 );
buf ( n49278 , n49277 );
nor ( n3486 , n49194 , n49205 , n49243 , n49278 );
buf ( n49280 , n3486 );
nand ( n3488 , n3211 , n49280 );
nand ( n3489 , n3390 , n3388 );
nand ( n3490 , n3266 , n3308 );
buf ( n49284 , n3324 );
buf ( n49285 , n49186 );
nand ( n3493 , n49284 , n49285 );
buf ( n49287 , n3493 );
nand ( n3495 , n3489 , n3490 , n49287 );
buf ( n49289 , n46270 );
buf ( n49290 , n3476 );
nand ( n3500 , n49289 , n49290 );
buf ( n49292 , n3500 );
buf ( n49293 , C1 );
and ( n3511 , n3495 , n49293 , n49241 );
buf ( n49295 , n3511 );
buf ( n49296 , n3380 );
buf ( n49297 , n49287 );
nand ( n3515 , n49296 , n49297 );
buf ( n49299 , n3515 );
buf ( n49300 , n49299 );
and ( n3518 , n49295 , n49300 );
buf ( n49302 , n49259 );
not ( n3520 , n49302 );
buf ( n49304 , n3465 );
not ( n3522 , n49304 );
or ( n3523 , n3520 , n3522 );
buf ( n49307 , n49240 );
not ( n3525 , n49307 );
buf ( n49309 , n49222 );
nand ( n3527 , n3525 , n49309 );
buf ( n49311 , n3527 );
buf ( n49312 , n49311 );
nand ( n3530 , n3523 , n49312 );
buf ( n49314 , n3530 );
not ( n3532 , n49314 );
nand ( n3533 , n3532 , n49292 );
not ( n3534 , n3533 );
or ( n3536 , n3534 , C0 );
buf ( n49319 , n46270 );
buf ( n49320 , n46246 );
nand ( n3539 , n49319 , n49320 );
buf ( n49322 , n3539 );
nand ( n3541 , n3536 , n49322 );
buf ( n49324 , n3541 );
nor ( n3543 , n3518 , n49324 );
buf ( n49326 , n3543 );
buf ( n49327 , n2952 );
buf ( n49328 , n48791 );
nand ( n3547 , n49327 , n49328 );
buf ( n49330 , n3547 );
buf ( n49331 , n49330 );
not ( n3550 , n49331 );
buf ( n49333 , n48752 );
nand ( n3552 , n3550 , n49333 );
buf ( n49335 , n3552 );
buf ( n49336 , n49335 );
buf ( n49337 , n2909 );
not ( n3556 , n49337 );
buf ( n49339 , n3556 );
buf ( n49340 , n49339 );
buf ( n49341 , n2936 );
not ( n3560 , n49341 );
buf ( n49343 , n3560 );
buf ( n49344 , n49343 );
nand ( n3563 , n49340 , n49344 );
buf ( n49346 , n3563 );
buf ( n49347 , n49346 );
nand ( n3566 , n49336 , n49347 );
buf ( n49349 , n3566 );
not ( n3568 , n49349 );
not ( n3569 , n3114 );
or ( n3570 , n3568 , n3569 );
buf ( n49353 , n3194 );
buf ( n49354 , n3208 );
nand ( n3573 , n49353 , n49354 );
buf ( n49356 , n3573 );
buf ( n49357 , n48926 );
not ( n3576 , n49357 );
buf ( n49359 , n3086 );
nand ( n3578 , n3576 , n49359 );
buf ( n49361 , n3578 );
nand ( n3580 , n49356 , n49361 );
not ( n3581 , n3580 );
nand ( n3582 , n3570 , n3581 );
not ( n3583 , n3324 );
not ( n3584 , n49186 );
and ( n3585 , n3583 , n3584 );
nor ( n3586 , n3585 , n49242 );
and ( n3587 , n3586 , n3210 );
not ( n3588 , n3391 );
and ( n3589 , n49293 , n3588 , n3310 );
nand ( n3590 , n3582 , n3587 , n3589 );
nand ( n3591 , n3488 , n49326 , n3590 );
not ( n3592 , n3591 );
not ( n3593 , n3592 );
or ( n3594 , C0 , n3593 );
buf ( n49377 , n49322 );
not ( n3598 , n49377 );
or ( n3599 , C0 , n3598 );
not ( n3600 , n49326 );
buf ( n49381 , n3600 );
nand ( n3602 , n3599 , n49381 );
buf ( n49383 , n3602 );
nand ( n3604 , n3594 , n49383 );
buf ( n49385 , n3604 );
buf ( n49386 , n381 );
not ( n3607 , n49386 );
buf ( n49388 , n3607 );
not ( n3609 , n380 );
and ( n3610 , n49388 , n3609 );
and ( n3611 , n380 , n381 );
nor ( n3612 , n3610 , n3611 );
buf ( n49393 , n382 );
not ( n3614 , n49393 );
buf ( n49395 , n3614 );
and ( n3616 , n381 , n49395 );
not ( n3617 , n381 );
and ( n3618 , n3617 , n382 );
nor ( n3619 , n3616 , n3618 );
and ( n3620 , n3612 , n3619 );
buf ( n49401 , n3620 );
not ( n3622 , n3619 );
buf ( n49403 , n3622 );
nor ( n3624 , n49401 , n49403 );
buf ( n49405 , n3624 );
buf ( n49406 , n49405 );
buf ( n49407 , n3609 );
or ( n3628 , n49406 , n49407 );
buf ( n49409 , n3628 );
buf ( n49410 , n49409 );
not ( n3631 , n49410 );
buf ( n49412 , n3631 );
buf ( n49413 , n49412 );
and ( n3634 , n49385 , n49413 );
buf ( n49415 , n3634 );
buf ( n49416 , n49415 );
buf ( n3637 , n49416 );
buf ( n49418 , n3637 );
buf ( n49419 , n49418 );
not ( n3640 , n49419 );
buf ( n49421 , n3640 );
buf ( n49422 , n49421 );
not ( n3644 , n3592 );
or ( n3645 , C0 , n3644 );
nand ( n3646 , n3645 , n49383 );
buf ( n49426 , n3646 );
and ( n3648 , n379 , n3609 );
not ( n3649 , n379 );
and ( n3650 , n3649 , n380 );
or ( n3651 , n3648 , n3650 );
not ( n3652 , n3651 );
buf ( n49432 , n3652 );
not ( n3654 , n378 );
buf ( n49434 , n3654 );
buf ( n49435 , n379 );
not ( n3657 , n49435 );
buf ( n49437 , n3657 );
buf ( n49438 , n49437 );
and ( n3660 , n49434 , n49438 );
buf ( n49440 , n378 );
buf ( n49441 , n379 );
and ( n3663 , n49440 , n49441 );
nor ( n3664 , n3660 , n3663 );
buf ( n49444 , n3664 );
buf ( n49445 , n49444 );
and ( n3667 , n49432 , n49445 );
buf ( n49447 , n3667 );
buf ( n49448 , n49447 );
not ( n3670 , n49448 );
buf ( n49450 , n3670 );
buf ( n49451 , n49450 );
buf ( n49452 , n3652 );
nand ( n3674 , n49451 , n49452 );
buf ( n49454 , n3674 );
buf ( n49455 , n49454 );
buf ( n49456 , n378 );
and ( n3678 , n49455 , n49456 );
buf ( n49458 , n3678 );
buf ( n49459 , n49458 );
nand ( n3681 , n49426 , n49459 );
buf ( n49461 , n3681 );
buf ( n49462 , n49461 );
buf ( n49463 , n49412 );
buf ( n49464 , n49458 );
nand ( n3686 , n49463 , n49464 );
buf ( n49466 , n3686 );
buf ( n49467 , n49466 );
and ( n3689 , n49422 , n49462 , n49467 );
buf ( n49469 , n3689 );
buf ( n49470 , n49469 );
not ( n3692 , n49470 );
buf ( n49472 , n3592 );
not ( n3696 , n49472 );
or ( n3697 , C0 , n3696 );
buf ( n49475 , n49383 );
nand ( n3699 , n3697 , n49475 );
buf ( n49477 , n3699 );
or ( n3701 , n49477 , n49412 );
nand ( n3702 , n3604 , n49412 );
nand ( n3703 , n3701 , n3702 );
buf ( n49481 , n3703 );
buf ( n49482 , n384 );
buf ( n49483 , n49458 );
not ( n3707 , n49483 );
buf ( n49485 , n3707 );
buf ( n49486 , n49485 );
and ( n3710 , n49482 , n49486 );
not ( n3711 , n49482 );
buf ( n49489 , n49458 );
and ( n3713 , n3711 , n49489 );
nor ( n3714 , n3710 , n3713 );
buf ( n49492 , n3714 );
xor ( n3716 , n383 , n384 );
buf ( n49494 , n3716 );
not ( n3718 , n49494 );
buf ( n49496 , n3718 );
buf ( n49497 , n49496 );
not ( n3721 , n49497 );
buf ( n49499 , n49395 );
buf ( n49500 , n383 );
not ( n3724 , n49500 );
buf ( n49502 , n3724 );
buf ( n49503 , n49502 );
and ( n3727 , n49499 , n49503 );
buf ( n49505 , n382 );
buf ( n49506 , n383 );
and ( n3730 , n49505 , n49506 );
nor ( n3731 , n3727 , n3730 );
buf ( n49509 , n3731 );
and ( n3733 , n49496 , n49509 );
not ( n3734 , n3733 );
buf ( n49512 , n3734 );
not ( n3736 , n49512 );
or ( n3737 , n3721 , n3736 );
buf ( n49515 , n382 );
nand ( n3739 , n3737 , n49515 );
buf ( n49517 , n3739 );
buf ( n49518 , n49517 );
not ( n3742 , n49518 );
buf ( n49520 , n3742 );
and ( n3744 , n49492 , n49520 );
not ( n3745 , n49492 );
and ( n3746 , n3745 , n49517 );
or ( n3747 , n3744 , n3746 );
not ( n3748 , n3747 );
buf ( n49526 , n3748 );
nand ( n3750 , n49481 , n49526 );
buf ( n49528 , n3750 );
buf ( n49529 , n49528 );
nand ( n3753 , n3692 , n49529 );
buf ( n49531 , n3753 );
buf ( n49532 , n49531 );
buf ( n49533 , n3748 );
not ( n3757 , n49533 );
buf ( n49535 , n3703 );
not ( n3759 , n49535 );
buf ( n49537 , n3759 );
buf ( n49538 , n49537 );
nand ( n3762 , n3757 , n49538 );
buf ( n49540 , n3762 );
buf ( n49541 , n49540 );
nand ( n3765 , n49532 , n49541 );
buf ( n49543 , n3765 );
buf ( n49544 , n49537 );
not ( n3768 , n49544 );
buf ( n49546 , n3768 );
not ( n3770 , n49546 );
buf ( n49548 , n49415 );
not ( n3772 , n49548 );
buf ( n49550 , n49520 );
buf ( n49551 , n384 );
and ( n3775 , n49550 , n49551 );
buf ( n49553 , n3775 );
buf ( n49554 , n49553 );
not ( n3778 , n49554 );
buf ( n49556 , n3778 );
buf ( n49557 , n384 );
not ( n3781 , n49557 );
buf ( n49559 , n49517 );
nand ( n3783 , n3781 , n49559 );
buf ( n49561 , n3783 );
nand ( n3785 , n49561 , n49458 );
and ( n3786 , n49556 , n3785 );
buf ( n49564 , n3786 );
not ( n3788 , n49564 );
and ( n3789 , n3772 , n3788 );
buf ( n49567 , n49415 );
buf ( n49568 , n3786 );
and ( n3792 , n49567 , n49568 );
nor ( n3793 , n3789 , n3792 );
buf ( n49571 , n3793 );
buf ( n49572 , n49571 );
not ( n3796 , n49572 );
buf ( n49574 , n3796 );
not ( n3798 , n49574 );
or ( n3799 , n3770 , n3798 );
buf ( n49577 , n49571 );
buf ( n49578 , n49537 );
nand ( n3802 , n49577 , n49578 );
buf ( n49580 , n3802 );
nand ( n3804 , n3799 , n49580 );
not ( n3805 , n3747 );
or ( n3806 , n3804 , n3805 );
nand ( n3807 , n3804 , n3748 );
nand ( n3808 , n3806 , n3807 );
buf ( n49586 , n3808 );
not ( n3810 , n49586 );
buf ( n49588 , n3810 );
and ( n3812 , n49543 , n49588 );
not ( n3813 , n49543 );
and ( n3814 , n3813 , n3808 );
or ( n3815 , n3812 , n3814 );
buf ( n49593 , n49561 );
not ( n3817 , n49593 );
buf ( n49595 , n49418 );
not ( n3819 , n49595 );
or ( n3820 , n3817 , n3819 );
buf ( n49598 , n49556 );
nand ( n3822 , n3820 , n49598 );
buf ( n49600 , n3822 );
not ( n3824 , n49469 );
not ( n3825 , n3824 );
and ( n3826 , n3747 , n49546 );
not ( n3827 , n3747 );
and ( n3828 , n3827 , n49537 );
or ( n3829 , n3826 , n3828 );
not ( n3830 , n3829 );
not ( n3831 , n3830 );
or ( n3832 , n3825 , n3831 );
nand ( n3833 , n3829 , n49469 );
nand ( n3834 , n3832 , n3833 );
xor ( n3835 , n49600 , n3834 );
buf ( n49613 , n384 );
buf ( n49614 , n49517 );
and ( n3838 , n49613 , n49614 );
not ( n3839 , n49613 );
buf ( n49617 , n49520 );
and ( n3841 , n3839 , n49617 );
nor ( n3842 , n3838 , n3841 );
buf ( n49620 , n3842 );
not ( n3844 , n49620 );
not ( n3845 , n49421 );
or ( n3846 , n3844 , n3845 );
buf ( n49624 , n49620 );
not ( n3848 , n49624 );
buf ( n49626 , n3848 );
nand ( n3850 , n49626 , n49418 );
nand ( n3851 , n3846 , n3850 );
buf ( n49629 , n3851 );
not ( n3853 , n49629 );
not ( n3854 , n49458 );
not ( n3855 , n3703 );
or ( n3856 , n3854 , n3855 );
buf ( n49634 , n49537 );
buf ( n49635 , n49485 );
nand ( n3859 , n49634 , n49635 );
buf ( n49637 , n3859 );
nand ( n3861 , n3856 , n49637 );
buf ( n49639 , n3861 );
not ( n3863 , n49639 );
buf ( n49641 , n3863 );
buf ( n49642 , n49641 );
not ( n3866 , n49642 );
or ( n3867 , n3853 , n3866 );
not ( n3868 , n3786 );
buf ( n49646 , n3868 );
nand ( n3870 , n3867 , n49646 );
buf ( n49648 , n3870 );
buf ( n49649 , n49648 );
buf ( n49650 , n3851 );
not ( n3874 , n49650 );
buf ( n49652 , n3861 );
nand ( n3876 , n3874 , n49652 );
buf ( n49654 , n3876 );
buf ( n49655 , n49654 );
nand ( n3879 , n49649 , n49655 );
buf ( n49657 , n3879 );
and ( n3881 , n3835 , n49657 );
and ( n3882 , n49600 , n3834 );
or ( n3883 , n3881 , n3882 );
buf ( n49661 , C0 );
nor ( n3886 , n3815 , n3883 );
buf ( n49663 , n3886 );
nor ( n3888 , n49661 , n49663 );
buf ( n49665 , n3888 );
buf ( n49666 , n49665 );
not ( n3891 , n49666 );
buf ( n49668 , n3891 );
buf ( n49669 , n49668 );
buf ( n49670 , n49665 );
xor ( n3895 , n49600 , n3834 );
xor ( n3896 , n3895 , n49657 );
not ( n3897 , n49528 );
not ( n3898 , n49553 );
or ( n3899 , n3897 , n3898 );
nand ( n3900 , n3899 , n49540 );
buf ( n49677 , n3900 );
not ( n3902 , n49677 );
buf ( n49679 , n3902 );
buf ( n49680 , n49679 );
not ( n3905 , n49680 );
xor ( n3906 , n3786 , n3861 );
xnor ( n3907 , n3906 , n3851 );
buf ( n49684 , n3907 );
not ( n3909 , n49684 );
or ( n3910 , n3905 , n3909 );
buf ( n49687 , n49626 );
buf ( n49688 , n49553 );
nor ( n3913 , n49687 , n49688 );
buf ( n49690 , n3913 );
buf ( n49691 , n49690 );
buf ( n49692 , n49409 );
or ( n3917 , n49691 , n49692 );
buf ( n49694 , n3917 );
buf ( n49695 , n49694 );
buf ( n49696 , n49626 );
not ( n3921 , n49696 );
buf ( n49698 , n49553 );
buf ( n49699 , n49409 );
and ( n3924 , n49698 , n49699 );
buf ( n49701 , n49556 );
buf ( n49702 , n49412 );
and ( n3927 , n49701 , n49702 );
nor ( n3928 , n3924 , n3927 );
buf ( n49705 , n3928 );
buf ( n49706 , n49705 );
not ( n3931 , n49706 );
or ( n3932 , n3921 , n3931 );
buf ( n49709 , n49705 );
buf ( n49710 , n49626 );
or ( n3935 , n49709 , n49710 );
nand ( n3936 , n3932 , n3935 );
buf ( n49713 , n3936 );
buf ( n49714 , n49713 );
not ( n3939 , n49714 );
buf ( n49716 , n49694 );
nand ( n3941 , n3939 , n49716 );
buf ( n49718 , n3941 );
nand ( n3943 , n49718 , n3646 );
buf ( n49720 , n3943 );
xor ( n3945 , n49695 , n49720 );
buf ( n49722 , n49553 );
buf ( n49723 , n3747 );
xor ( n3948 , n49722 , n49723 );
buf ( n49725 , n49537 );
xnor ( n3950 , n3948 , n49725 );
buf ( n49727 , n3950 );
buf ( n49728 , n49727 );
and ( n3953 , n3945 , n49728 );
and ( n3954 , n49695 , n49720 );
or ( n3955 , n3953 , n3954 );
buf ( n49732 , n3955 );
buf ( n49733 , n49732 );
not ( n3958 , n49733 );
buf ( n49735 , n3958 );
buf ( n49736 , n49735 );
nand ( n3961 , n3910 , n49736 );
buf ( n49738 , n3961 );
buf ( n49739 , n49738 );
buf ( n49740 , n3907 );
not ( n3965 , n49740 );
buf ( n49742 , n3900 );
nand ( n3967 , n3965 , n49742 );
buf ( n49744 , n3967 );
buf ( n49745 , n49744 );
nand ( n3970 , n49739 , n49745 );
buf ( n49747 , n3970 );
or ( n3972 , n3896 , n49747 );
not ( n3973 , n45352 );
not ( n3974 , n45346 );
not ( n3975 , n3974 );
not ( n3976 , n45326 );
or ( n3977 , n3975 , n3976 );
buf ( n3978 , n45270 );
and ( n3979 , n45345 , n3978 , n45243 );
nor ( n3980 , n3979 , n45471 );
buf ( n3981 , n3980 );
nand ( n3982 , n3977 , n3981 );
not ( n3983 , n3982 );
or ( n3984 , n3973 , n3983 );
not ( n3985 , n44688 );
not ( n3986 , n44829 );
or ( n3987 , n3985 , n3986 );
nand ( n3988 , n3987 , n45377 );
not ( n3989 , n3988 );
buf ( n3990 , n3989 );
not ( n3991 , n45380 );
not ( n3992 , n44303 );
not ( n3993 , n3992 );
or ( n3994 , n3991 , n3993 );
or ( n3995 , n44683 , n44525 );
nand ( n3996 , n3994 , n3995 );
not ( n3997 , n3996 );
not ( n3998 , n44303 );
not ( n3999 , n44520 );
or ( n4000 , n3998 , n3999 );
nand ( n4001 , n4000 , n45383 );
not ( n4002 , n4001 );
buf ( n49779 , n44095 );
not ( n4004 , n49779 );
buf ( n49781 , n4004 );
not ( n4006 , n49781 );
not ( n4007 , n44298 );
not ( n4008 , n4007 );
or ( n4009 , n4006 , n4008 );
nor ( n4010 , n44090 , n43887 );
and ( n4011 , n43656 , n43441 );
nor ( n4012 , n4011 , n43661 );
or ( n4013 , n43656 , n43441 );
not ( n4014 , n43253 );
not ( n4015 , n43079 );
and ( n4016 , n4014 , n4015 );
not ( n4017 , n43258 );
nor ( n4018 , n4016 , n4017 );
and ( n4019 , n45454 , n4018 );
nor ( n4020 , n4019 , n43436 );
nor ( n4021 , n4020 , n45464 );
nand ( n4022 , n4013 , n4021 );
nand ( n4023 , n4012 , n4022 );
and ( n4024 , n4023 , n43882 );
nand ( n4025 , n43656 , n43441 );
and ( n4026 , n4022 , n4025 );
not ( n4027 , n43661 );
nor ( n4028 , n4026 , n4027 );
nor ( n4029 , n4024 , n4028 );
or ( n4030 , n4010 , n4029 );
buf ( n49807 , n44090 );
buf ( n49808 , n43887 );
nand ( n4033 , n49807 , n49808 );
buf ( n49810 , n4033 );
nand ( n4035 , n4030 , n49810 );
nand ( n4036 , n4009 , n4035 );
nand ( n4037 , n4002 , n4036 );
nand ( n4038 , n3997 , n4037 );
buf ( n4039 , n4038 );
and ( n4040 , n3990 , n4039 );
not ( n4041 , n44945 );
not ( n4042 , n44834 );
and ( n4043 , n4041 , n4042 );
nor ( n4044 , n44688 , n44829 );
nor ( n4045 , n4043 , n4044 );
not ( n4046 , n4045 );
nor ( n4047 , n4040 , n4046 );
nor ( n4048 , n4047 , n45373 );
not ( n4049 , n4048 );
and ( n4050 , n45357 , n4049 );
nor ( n4051 , n4050 , n45478 );
nand ( n4052 , n3984 , n4051 );
not ( n4053 , n4052 );
not ( n4054 , n4053 );
buf ( n49831 , n4054 );
buf ( n49832 , n378 );
nand ( n4057 , n49831 , n49832 );
buf ( n49834 , n4057 );
buf ( n49835 , n49834 );
not ( n4060 , n49835 );
xor ( n4061 , n49695 , n49720 );
xor ( n4062 , n4061 , n49728 );
buf ( n49839 , n4062 );
buf ( n49840 , n49839 );
not ( n4065 , n49840 );
or ( n4066 , n4060 , n4065 );
buf ( n49843 , n49447 );
not ( n4068 , n49843 );
buf ( n49845 , n378 );
not ( n4070 , n49845 );
nand ( n4071 , n45351 , n45474 );
not ( n4072 , n4071 );
not ( n4073 , n3982 );
or ( n4074 , n4072 , n4073 );
nand ( n4075 , n4074 , n4051 );
not ( n4076 , n4075 );
buf ( n49853 , n4076 );
not ( n4078 , n49853 );
or ( n4079 , n4070 , n4078 );
buf ( n49856 , n4054 );
buf ( n49857 , n3654 );
nand ( n4082 , n49856 , n49857 );
buf ( n49859 , n4082 );
buf ( n49860 , n49859 );
nand ( n4085 , n4079 , n49860 );
buf ( n49862 , n4085 );
buf ( n49863 , n49862 );
not ( n4088 , n49863 );
or ( n4089 , n4068 , n4088 );
buf ( n49866 , n3651 );
buf ( n49867 , n378 );
nand ( n4092 , n49866 , n49867 );
buf ( n49869 , n4092 );
buf ( n49870 , n49869 );
nand ( n4095 , n4089 , n49870 );
buf ( n49872 , n4095 );
buf ( n49873 , n49872 );
not ( n4098 , n3974 );
nor ( n4099 , n45189 , n45133 );
not ( n4100 , n4099 );
not ( n4101 , n45128 );
nand ( n4102 , n4101 , n45293 );
nand ( n4103 , n4100 , n4102 , n45310 );
buf ( n49880 , n45336 );
not ( n4105 , n49880 );
buf ( n49882 , n4105 );
nor ( n4107 , n4103 , n49882 );
not ( n4108 , n4107 );
not ( n4109 , n3989 );
not ( n4110 , n3996 );
nand ( n4111 , n4110 , n4037 );
not ( n4112 , n4111 );
or ( n4113 , n4109 , n4112 );
nand ( n4114 , n4113 , n4045 );
buf ( n4115 , n45370 );
nand ( n4116 , n4114 , n4115 );
not ( n4117 , n4116 );
or ( n4118 , n4108 , n4117 );
nand ( n4119 , n4118 , n45323 );
not ( n4120 , n4119 );
or ( n4121 , n4098 , n4120 );
nand ( n4122 , n4121 , n3981 );
not ( n4123 , n45478 );
nand ( n4124 , n4123 , n45352 );
not ( n4125 , n4124 );
and ( n4126 , n4122 , n4125 );
not ( n4127 , n4122 );
and ( n4128 , n4127 , n4124 );
nor ( n4129 , n4126 , n4128 );
not ( n4130 , n4129 );
buf ( n49907 , n4130 );
not ( n4132 , n49907 );
buf ( n49909 , n378 );
nand ( n4134 , n4132 , n49909 );
buf ( n49911 , n4134 );
buf ( n49912 , n49911 );
not ( n4137 , n49912 );
buf ( n49914 , n4137 );
buf ( n49915 , n49914 );
or ( n4140 , n49873 , n49915 );
buf ( n49917 , n49718 );
buf ( n49918 , n3646 );
and ( n49919 , n49917 , n49918 );
not ( n4144 , n49917 );
not ( n4146 , n3592 );
or ( n49922 , C0 , n4146 );
nand ( n4148 , n49922 , n49383 );
not ( n49924 , n4148 );
buf ( n49925 , n49924 );
and ( n49926 , n4144 , n49925 );
nor ( n4152 , n49919 , n49926 );
buf ( n49928 , n4152 );
buf ( n49929 , n49928 );
nand ( n49930 , n4140 , n49929 );
buf ( n49931 , n49930 );
buf ( n49932 , n49931 );
buf ( n49933 , n49872 );
buf ( n49934 , n49914 );
nand ( n4160 , n49933 , n49934 );
buf ( n49936 , n4160 );
buf ( n49937 , n49936 );
nand ( n49938 , n49932 , n49937 );
buf ( n49939 , n49938 );
buf ( n49940 , n49939 );
nand ( n4166 , n4066 , n49940 );
buf ( n49942 , n4166 );
buf ( n49943 , n49834 );
not ( n49944 , n49943 );
buf ( n49945 , n49839 );
not ( n49946 , n49945 );
buf ( n49947 , n49946 );
buf ( n49948 , n49947 );
nand ( n4174 , n49944 , n49948 );
buf ( n49950 , n4174 );
nand ( n4176 , n49942 , n49950 );
not ( n49952 , n4176 );
not ( n4178 , n49679 );
not ( n49954 , n49735 );
or ( n4180 , n4178 , n49954 );
nand ( n49956 , n49732 , n3900 );
nand ( n4182 , n4180 , n49956 );
not ( n49958 , n4182 );
and ( n4186 , n49958 , n3907 );
nor ( n49960 , C0 , n4186 );
not ( n4188 , n49960 );
nand ( n49962 , n49952 , n4188 );
buf ( n4190 , n49962 );
and ( n49964 , n3972 , n4190 );
not ( n4192 , n49964 );
buf ( n49966 , n49626 );
buf ( n49967 , n378 );
buf ( n49968 , n45133 );
not ( n4196 , n49968 );
buf ( n49970 , n45189 );
buf ( n4198 , n49970 );
buf ( n49972 , n4198 );
not ( n4200 , n49972 );
and ( n49974 , n4196 , n4200 );
not ( n4202 , n4114 );
nand ( n49976 , n4202 , n45338 );
not ( n4204 , n45128 );
not ( n49978 , n45047 );
and ( n4206 , n4204 , n49978 );
buf ( n49980 , n44945 );
buf ( n49981 , n44834 );
nand ( n49982 , n49980 , n49981 );
buf ( n49983 , n49982 );
nor ( n49984 , n4206 , n49983 );
not ( n4212 , n49984 );
not ( n49986 , n45336 );
or ( n4214 , n4212 , n49986 );
nand ( n49988 , n4214 , n45303 );
nor ( n4216 , n49988 , n45317 );
and ( n49990 , n49976 , n4216 );
nor ( n4218 , n49974 , n49990 );
nand ( n49992 , n45321 , n45314 );
and ( n4220 , n4218 , n49992 );
not ( n49994 , n4218 );
not ( n4222 , n49992 );
and ( n49996 , n49994 , n4222 );
nor ( n4224 , n4220 , n49996 );
not ( n49998 , n4224 );
buf ( n49999 , n49998 );
and ( n50000 , n49967 , n49999 );
buf ( n50001 , n50000 );
buf ( n50002 , n50001 );
xor ( n4230 , n49966 , n50002 );
not ( n50004 , n3588 );
buf ( n50005 , n3211 );
not ( n50006 , n50005 );
buf ( n50007 , n50006 );
buf ( n50008 , n50007 );
not ( n4236 , n50008 );
buf ( n50010 , n4236 );
buf ( n50011 , n49349 );
buf ( n50012 , n3210 );
buf ( n50013 , n3114 );
and ( n50014 , n50011 , n50012 , n50013 );
buf ( n50015 , n50014 );
buf ( n50016 , n50015 );
not ( n4244 , n50016 );
buf ( n50018 , n3580 );
buf ( n50019 , n3210 );
nand ( n50020 , n50018 , n50019 );
buf ( n50021 , n50020 );
buf ( n50022 , n50021 );
nand ( n4250 , n4244 , n50022 );
buf ( n50024 , n4250 );
or ( n4252 , n50010 , n50024 );
not ( n50026 , n4252 );
or ( n4254 , n50004 , n50026 );
nand ( n50028 , n4254 , n3489 );
buf ( n50029 , n50028 );
buf ( n50030 , n3310 );
buf ( n50031 , n3490 );
nand ( n50032 , n50030 , n50031 );
buf ( n50033 , n50032 );
buf ( n50034 , n50033 );
not ( n4262 , n50034 );
buf ( n50036 , n4262 );
buf ( n50037 , n50036 );
and ( n4265 , n50029 , n50037 );
not ( n50039 , n50029 );
buf ( n50040 , n50033 );
and ( n4268 , n50039 , n50040 );
nor ( n50042 , n4265 , n4268 );
buf ( n50043 , n50042 );
buf ( n50044 , n50043 );
and ( n4272 , n4230 , n50044 );
and ( n4273 , n49966 , n50002 );
or ( n4274 , n4272 , n4273 );
buf ( n50048 , n4274 );
not ( n4276 , n3620 );
not ( n4277 , n380 );
not ( n4278 , n4076 );
or ( n4279 , n4277 , n4278 );
or ( n4280 , n4076 , n380 );
nand ( n4281 , n4279 , n4280 );
not ( n4282 , n4281 );
or ( n4283 , n4276 , n4282 );
nand ( n4284 , n3622 , n380 );
nand ( n4285 , n4283 , n4284 );
not ( n4286 , n4285 );
xor ( n4287 , n50048 , n4286 );
not ( n4288 , n3489 );
nor ( n4289 , n3391 , n4288 );
not ( n4290 , n4289 );
not ( n4291 , n4290 );
not ( n4292 , n4252 );
or ( n4293 , n4291 , n4292 );
not ( n4294 , n50010 );
not ( n4295 , n50024 );
nand ( n4296 , n4294 , n4295 , n4289 );
nand ( n4297 , n4293 , n4296 );
and ( n4298 , n384 , n4297 );
not ( n4299 , n4298 );
buf ( n50073 , n3620 );
not ( n4301 , n50073 );
not ( n4302 , n4122 );
not ( n4303 , n3609 );
nor ( n4304 , n4303 , n4124 );
nand ( n4305 , n4302 , n4304 );
and ( n4306 , n4124 , n380 );
nand ( n4307 , n4302 , n4306 );
and ( n4308 , n4124 , n3609 );
nand ( n4309 , n4308 , n4122 );
not ( n4310 , n380 );
nor ( n4311 , n4310 , n4124 );
nand ( n4312 , n4311 , n4122 );
nand ( n4313 , n4305 , n4307 , n4309 , n4312 );
buf ( n50087 , n4313 );
not ( n4315 , n50087 );
or ( n4316 , n4301 , n4315 );
nand ( n4317 , n4281 , n3622 );
buf ( n50091 , n4317 );
nand ( n4319 , n4316 , n50091 );
buf ( n50093 , n4319 );
not ( n4321 , n50093 );
or ( n4322 , n4299 , n4321 );
buf ( n50096 , n50093 );
buf ( n50097 , n4298 );
or ( n4325 , n50096 , n50097 );
buf ( n50099 , n3651 );
not ( n4327 , n50099 );
buf ( n50101 , n378 );
and ( n4329 , n45468 , n45345 );
not ( n4330 , n4329 );
or ( n4331 , n45484 , n4048 );
not ( n4332 , n45479 );
not ( n4333 , n45304 );
not ( n4334 , n4333 );
and ( n4335 , n4332 , n4334 );
not ( n4336 , n45243 );
not ( n4337 , n45270 );
or ( n4338 , n4336 , n4337 );
nand ( n4339 , n45322 , n45341 );
nand ( n4340 , n4338 , n4339 );
nor ( n4341 , n4335 , n4340 );
nand ( n4342 , n4331 , n4341 );
not ( n4343 , n4342 );
or ( n4344 , n4330 , n4343 );
or ( n4345 , n45484 , n4048 );
not ( n4346 , n4329 );
nand ( n4347 , n4345 , n4341 , n4346 );
nand ( n4348 , n4344 , n4347 );
not ( n4349 , n4348 );
buf ( n50123 , n4349 );
not ( n4351 , n50123 );
buf ( n50125 , n4351 );
buf ( n50126 , n50125 );
and ( n4354 , n50101 , n50126 );
not ( n4355 , n50101 );
buf ( n50129 , n4349 );
and ( n4357 , n4355 , n50129 );
nor ( n4358 , n4354 , n4357 );
buf ( n50132 , n4358 );
buf ( n50133 , n50132 );
not ( n4361 , n50133 );
buf ( n50135 , n4361 );
buf ( n50136 , n50135 );
not ( n4364 , n50136 );
or ( n4365 , n4327 , n4364 );
buf ( n50139 , n378 );
nand ( n4367 , n3978 , n45243 );
and ( n4368 , n4367 , n45341 );
xor ( n4369 , n4119 , n4368 );
buf ( n50143 , n4369 );
xor ( n4371 , n50139 , n50143 );
buf ( n50145 , n4371 );
buf ( n50146 , n50145 );
buf ( n50147 , n49447 );
nand ( n4375 , n50146 , n50147 );
buf ( n50149 , n4375 );
buf ( n50150 , n50149 );
nand ( n4378 , n4365 , n50150 );
buf ( n50152 , n4378 );
buf ( n50153 , n50152 );
nand ( n4381 , n4325 , n50153 );
buf ( n50155 , n4381 );
nand ( n4383 , n4322 , n50155 );
xnor ( n4384 , n4287 , n4383 );
buf ( n50158 , n4384 );
not ( n4386 , n45317 );
not ( n4387 , n4386 );
buf ( n50161 , n49968 );
buf ( n50162 , n49972 );
nor ( n4390 , n50161 , n50162 );
buf ( n50164 , n4390 );
nor ( n4392 , n4387 , n50164 );
not ( n4393 , n4392 );
buf ( n50167 , n44688 );
buf ( n50168 , n44829 );
nor ( n4396 , n50167 , n50168 );
buf ( n50170 , n4396 );
not ( n4398 , n50170 );
not ( n4399 , n4398 );
not ( n4400 , n3988 );
or ( n4401 , n4399 , n4400 );
not ( n4402 , n4044 );
nand ( n4403 , n4402 , n4037 , n4110 );
nand ( n4404 , n4401 , n4403 );
not ( n4405 , n4404 );
not ( n4406 , n44945 );
not ( n4407 , n44834 );
nand ( n4408 , n4406 , n4407 );
not ( n4409 , n4408 );
nor ( n4410 , n45337 , n4409 );
not ( n4411 , n4410 );
or ( n4412 , n4405 , n4411 );
not ( n4413 , n49988 );
nand ( n4414 , n4412 , n4413 );
not ( n4415 , n4414 );
not ( n4416 , n4415 );
or ( n4417 , n4393 , n4416 );
not ( n4418 , n50164 );
nand ( n4419 , n4418 , n4386 );
nand ( n4420 , n4419 , n4414 );
nand ( n4421 , n4417 , n4420 );
buf ( n50195 , n4421 );
buf ( n50196 , n378 );
nand ( n4424 , n50195 , n50196 );
buf ( n50198 , n4424 );
nand ( n4426 , n3210 , n49356 );
not ( n4427 , n4426 );
not ( n4428 , n48800 );
not ( n4429 , n2684 );
or ( n4430 , n4428 , n4429 );
buf ( n50204 , n49349 );
not ( n4432 , n50204 );
buf ( n50206 , n4432 );
nand ( n4434 , n4430 , n50206 );
not ( n4435 , n4434 );
not ( n4436 , n3114 );
or ( n4437 , n4435 , n4436 );
buf ( n4438 , n49361 );
nand ( n4439 , n4437 , n4438 );
not ( n4440 , n4439 );
or ( n4441 , n4427 , n4440 );
or ( n4442 , n4426 , n4439 );
nand ( n4443 , n4441 , n4442 );
nand ( n4444 , n4443 , n384 );
nand ( n4445 , n50198 , n4444 );
buf ( n50219 , n4445 );
not ( n4447 , n50219 );
not ( n4448 , n3651 );
not ( n4449 , n50145 );
or ( n4450 , n4448 , n4449 );
xor ( n4451 , n49967 , n49999 );
buf ( n50225 , n4451 );
nand ( n4453 , n50225 , n49447 );
nand ( n4454 , n4450 , n4453 );
buf ( n50228 , n4454 );
not ( n4456 , n50228 );
or ( n4457 , n4447 , n4456 );
not ( n4458 , n4444 );
buf ( n50232 , n50198 );
not ( n4460 , n50232 );
buf ( n50234 , n4460 );
nand ( n4462 , n4458 , n50234 );
buf ( n50236 , n4462 );
nand ( n4464 , n4457 , n50236 );
buf ( n50238 , n4464 );
buf ( n50239 , n50238 );
xor ( n4467 , n49966 , n50002 );
xor ( n4468 , n4467 , n50044 );
buf ( n50242 , n4468 );
buf ( n50243 , n50242 );
xor ( n4471 , n50239 , n50243 );
xor ( n4472 , n384 , n4297 );
buf ( n50246 , n4472 );
buf ( n50247 , n3733 );
not ( n4475 , n50247 );
not ( n4476 , n382 );
not ( n4477 , n4052 );
not ( n4478 , n4477 );
or ( n4479 , n4476 , n4478 );
or ( n4480 , n4053 , n382 );
nand ( n4481 , n4479 , n4480 );
buf ( n50255 , n4481 );
not ( n4483 , n50255 );
or ( n4484 , n4475 , n4483 );
buf ( n50258 , n3716 );
buf ( n50259 , n382 );
nand ( n4487 , n50258 , n50259 );
buf ( n50261 , n4487 );
buf ( n50262 , n50261 );
nand ( n4490 , n4484 , n50262 );
buf ( n50264 , n4490 );
buf ( n50265 , n50264 );
xor ( n4493 , n50246 , n50265 );
buf ( n50267 , n3622 );
not ( n4495 , n50267 );
buf ( n50269 , n4313 );
not ( n4497 , n50269 );
or ( n4498 , n4495 , n4497 );
buf ( n50272 , n380 );
not ( n4500 , n50272 );
buf ( n50274 , n50125 );
not ( n4502 , n50274 );
or ( n4503 , n4500 , n4502 );
not ( n4504 , n4348 );
nand ( n4505 , n4504 , n3609 );
buf ( n50279 , n4505 );
nand ( n4507 , n4503 , n50279 );
buf ( n50281 , n4507 );
buf ( n50282 , n50281 );
buf ( n50283 , n3620 );
nand ( n4511 , n50282 , n50283 );
buf ( n50285 , n4511 );
buf ( n50286 , n50285 );
nand ( n4514 , n4498 , n50286 );
buf ( n50288 , n4514 );
buf ( n50289 , n50288 );
and ( n4517 , n4493 , n50289 );
and ( n4518 , n50246 , n50265 );
or ( n4519 , n4517 , n4518 );
buf ( n50293 , n4519 );
buf ( n50294 , n50293 );
and ( n4522 , n4471 , n50294 );
and ( n4523 , n50239 , n50243 );
or ( n4524 , n4522 , n4523 );
buf ( n50298 , n4524 );
buf ( n50299 , n50298 );
or ( n4527 , n50158 , n50299 );
and ( n4528 , n50139 , n50143 );
buf ( n50302 , n4528 );
buf ( n50303 , n50302 );
buf ( n50304 , n49287 );
buf ( n50305 , n49192 );
nand ( n4533 , n50304 , n50305 );
buf ( n50307 , n4533 );
buf ( n50308 , n50307 );
buf ( n50309 , n50010 );
buf ( n50310 , n50015 );
or ( n4538 , n50309 , n50310 );
buf ( n50312 , n3588 );
buf ( n50313 , n3310 );
nand ( n4541 , n50312 , n50313 );
buf ( n50315 , n4541 );
buf ( n50316 , n50315 );
not ( n4544 , n50316 );
buf ( n50318 , n4544 );
buf ( n50319 , n50318 );
nand ( n4547 , n4538 , n50319 );
buf ( n50321 , n4547 );
buf ( n50322 , n50321 );
not ( n4550 , n50021 );
not ( n4551 , n50315 );
and ( n4552 , n4550 , n4551 );
nand ( n4553 , n3310 , n4288 );
buf ( n50327 , n4553 );
buf ( n50328 , n3490 );
nand ( n4556 , n50327 , n50328 );
buf ( n50330 , n4556 );
nor ( n4558 , n4552 , n50330 );
buf ( n50332 , n4558 );
nand ( n4560 , n50322 , n50332 );
buf ( n50334 , n4560 );
buf ( n50335 , n50334 );
or ( n4563 , n50308 , n50335 );
buf ( n50337 , n50334 );
buf ( n50338 , n50307 );
nand ( n4566 , n50337 , n50338 );
buf ( n50340 , n4566 );
buf ( n50341 , n50340 );
nand ( n4569 , n4563 , n50341 );
buf ( n50343 , n4569 );
buf ( n50344 , n50343 );
buf ( n50345 , n49690 );
xnor ( n4573 , n50344 , n50345 );
buf ( n50347 , n4573 );
buf ( n50348 , n50347 );
xor ( n4576 , n50303 , n50348 );
not ( n4577 , n3651 );
buf ( n50351 , n378 );
not ( n4579 , n50351 );
buf ( n50353 , n4130 );
not ( n4581 , n50353 );
or ( n4582 , n4579 , n4581 );
not ( n4583 , n4125 );
not ( n4584 , n4302 );
or ( n4585 , n4583 , n4584 );
nand ( n4586 , n4124 , n4122 );
nand ( n4587 , n4585 , n4586 );
nand ( n4588 , n4587 , n3654 );
buf ( n50362 , n4588 );
nand ( n4590 , n4582 , n50362 );
buf ( n50364 , n4590 );
not ( n4592 , n50364 );
or ( n4593 , n4577 , n4592 );
or ( n4594 , n50132 , n49450 );
nand ( n4595 , n4593 , n4594 );
buf ( n50369 , n4595 );
xor ( n4597 , n4576 , n50369 );
buf ( n50371 , n4597 );
buf ( n50372 , n50371 );
nand ( n4600 , n4527 , n50372 );
buf ( n50374 , n4600 );
buf ( n50375 , n50374 );
buf ( n50376 , n50298 );
buf ( n50377 , n4384 );
nand ( n4605 , n50376 , n50377 );
buf ( n50379 , n4605 );
buf ( n50380 , n50379 );
nand ( n4608 , n50375 , n50380 );
buf ( n50382 , n4608 );
buf ( n50383 , n50382 );
not ( n4611 , n50383 );
and ( n4612 , n4349 , n378 );
not ( n4613 , n4612 );
xor ( n4614 , n49713 , n4613 );
buf ( n50388 , n49311 );
buf ( n50389 , n49241 );
nand ( n4617 , n50388 , n50389 );
buf ( n50391 , n4617 );
buf ( n50392 , n50391 );
not ( n4620 , n50392 );
not ( n4621 , n49192 );
not ( n4622 , n50334 );
or ( n4623 , n4621 , n4622 );
nand ( n4624 , n4623 , n49287 );
buf ( n50398 , n4624 );
not ( n4626 , n50398 );
or ( n4627 , n4620 , n4626 );
buf ( n50401 , n4624 );
buf ( n50402 , n50391 );
or ( n4630 , n50401 , n50402 );
nand ( n4631 , n4627 , n4630 );
buf ( n50405 , n4631 );
xnor ( n4633 , n4614 , n50405 );
not ( n4634 , n4285 );
not ( n4635 , n50048 );
or ( n4636 , n4634 , n4635 );
not ( n4637 , n4286 );
not ( n4638 , n50048 );
not ( n4639 , n4638 );
or ( n4640 , n4637 , n4639 );
nand ( n4641 , n4640 , n4383 );
nand ( n4642 , n4636 , n4641 );
xor ( n4643 , n4633 , n4642 );
buf ( n50417 , n49447 );
not ( n4645 , n50417 );
buf ( n50419 , n50364 );
not ( n4647 , n50419 );
or ( n4648 , n4645 , n4647 );
buf ( n50422 , n49862 );
buf ( n50423 , n3651 );
nand ( n4651 , n50422 , n50423 );
buf ( n50425 , n4651 );
buf ( n50426 , n50425 );
nand ( n4654 , n4648 , n50426 );
buf ( n50428 , n4654 );
buf ( n50429 , n50428 );
not ( n4657 , n50429 );
buf ( n50431 , n49690 );
not ( n4659 , n50431 );
buf ( n50433 , n50343 );
nand ( n4661 , n4659 , n50433 );
buf ( n50435 , n4661 );
buf ( n50436 , n50435 );
not ( n4664 , n50436 );
and ( n4665 , n4657 , n4664 );
buf ( n50439 , n50428 );
buf ( n50440 , n50435 );
and ( n4668 , n50439 , n50440 );
nor ( n4669 , n4665 , n4668 );
buf ( n50443 , n4669 );
xor ( n4671 , n50303 , n50348 );
and ( n4672 , n4671 , n50369 );
and ( n4673 , n50303 , n50348 );
or ( n4674 , n4672 , n4673 );
buf ( n50448 , n4674 );
xor ( n4676 , n50443 , n50448 );
xnor ( n4677 , n4643 , n4676 );
buf ( n50451 , n4677 );
not ( n4679 , n50451 );
buf ( n50453 , n4679 );
buf ( n50454 , n50453 );
nand ( n4682 , n4611 , n50454 );
buf ( n50456 , n4682 );
buf ( n50457 , n49834 );
buf ( n50458 , n49947 );
xor ( n4686 , n50457 , n50458 );
buf ( n50460 , n49939 );
xor ( n4688 , n4686 , n50460 );
buf ( n50462 , n4688 );
or ( n4690 , n49713 , n50405 );
nand ( n4691 , n4690 , n4612 );
nand ( n4692 , n50405 , n49713 );
nand ( n4693 , n4691 , n4692 );
buf ( n50467 , n4693 );
not ( n4695 , n50467 );
buf ( n50469 , n4695 );
not ( n4697 , n50469 );
buf ( n50471 , n50428 );
not ( n4699 , n50471 );
buf ( n50473 , n50435 );
nand ( n4701 , n4699 , n50473 );
buf ( n50475 , n4701 );
buf ( n50476 , n50475 );
not ( n4704 , n50476 );
buf ( n50478 , n50448 );
not ( n4706 , n50478 );
or ( n4707 , n4704 , n4706 );
buf ( n50481 , n50435 );
not ( n4709 , n50481 );
buf ( n50483 , n50428 );
nand ( n4711 , n4709 , n50483 );
buf ( n50485 , n4711 );
buf ( n50486 , n50485 );
nand ( n4714 , n4707 , n50486 );
buf ( n50488 , n4714 );
buf ( n50489 , n50488 );
not ( n4717 , n50489 );
buf ( n50491 , n4717 );
not ( n4719 , n50491 );
or ( n4720 , n4697 , n4719 );
xor ( n4721 , n49928 , n49911 );
xor ( n4722 , n4721 , n49872 );
not ( n4723 , n4722 );
nand ( n4724 , n4720 , n4723 );
nand ( n4725 , n50488 , n4693 );
nand ( n4726 , n50462 , n4724 , n4725 );
nand ( n4727 , n50456 , n4726 );
not ( n4728 , n4722 );
not ( n4729 , n4693 );
or ( n4730 , n4728 , n4729 );
or ( n4731 , n4722 , n4693 );
nand ( n4732 , n4730 , n4731 );
xor ( n4733 , n50488 , n4732 );
buf ( n50507 , n4733 );
not ( n4735 , n50507 );
buf ( n50509 , n4735 );
not ( n4737 , n4676 );
not ( n4738 , n4737 );
not ( n4739 , n4633 );
not ( n4740 , n4642 );
nand ( n4741 , n4739 , n4740 );
not ( n4742 , n4741 );
or ( n4743 , n4738 , n4742 );
not ( n4744 , n4740 );
nand ( n4745 , n4744 , n4633 );
nand ( n4746 , n4743 , n4745 );
not ( n4747 , n4746 );
nand ( n4748 , n50509 , n4747 );
buf ( n50522 , n4748 );
buf ( n50523 , n4298 );
buf ( n50524 , n50152 );
xor ( n4752 , n50523 , n50524 );
buf ( n50526 , n50093 );
xnor ( n4754 , n4752 , n50526 );
buf ( n50528 , n4754 );
buf ( n50529 , n50528 );
not ( n4757 , n50529 );
buf ( n50531 , n4116 );
buf ( n50532 , n45366 );
xor ( n4760 , n50531 , n50532 );
buf ( n50534 , n4760 );
buf ( n50535 , n50534 );
not ( n4763 , n50535 );
buf ( n50537 , n4763 );
buf ( n50538 , n50537 );
not ( n4766 , n50538 );
buf ( n50540 , n4766 );
buf ( n50541 , n49361 );
buf ( n50542 , n3114 );
nand ( n4770 , n50541 , n50542 );
buf ( n50544 , n4770 );
xnor ( n4772 , n4434 , n50544 );
nand ( n4773 , n378 , n50540 , n4772 );
buf ( n50547 , n4773 );
not ( n4775 , n50547 );
buf ( n50549 , n4775 );
buf ( n50550 , n50549 );
not ( n4778 , n50550 );
and ( n4779 , n3733 , n382 );
and ( n4780 , n4130 , n4779 );
and ( n4781 , n4481 , n3716 );
nor ( n4782 , n4780 , n4781 );
nand ( n4783 , n4587 , n49395 , n3733 );
nand ( n4784 , n4782 , n4783 );
buf ( n50558 , n4784 );
not ( n4786 , n50558 );
or ( n4787 , n4778 , n4786 );
buf ( n50561 , n4784 );
buf ( n50562 , n50549 );
or ( n4790 , n50561 , n50562 );
buf ( n50564 , n3622 );
not ( n4792 , n50564 );
buf ( n50566 , n50281 );
not ( n4794 , n50566 );
or ( n4795 , n4792 , n4794 );
buf ( n50569 , n4369 );
not ( n4797 , n50569 );
buf ( n50571 , n4797 );
nand ( n4799 , n380 , n50571 );
not ( n4800 , n4799 );
not ( n4801 , n380 );
nand ( n4802 , n4801 , n4369 );
not ( n4803 , n4802 );
or ( n4804 , n4800 , n4803 );
nand ( n4805 , n4804 , n3620 );
buf ( n50579 , n4805 );
nand ( n4807 , n4795 , n50579 );
buf ( n50581 , n4807 );
buf ( n50582 , n50581 );
nand ( n4810 , n4790 , n50582 );
buf ( n50584 , n4810 );
buf ( n50585 , n50584 );
nand ( n4813 , n4787 , n50585 );
buf ( n50587 , n4813 );
buf ( n50588 , n50587 );
not ( n4816 , n50588 );
not ( n4817 , n4454 );
not ( n4818 , n4817 );
and ( n4819 , n4444 , n50234 );
not ( n4820 , n4444 );
and ( n4821 , n4820 , n50198 );
nor ( n4822 , n4819 , n4821 );
not ( n4823 , n4822 );
not ( n4824 , n4823 );
or ( n4825 , n4818 , n4824 );
nand ( n4826 , n4822 , n4454 );
nand ( n4827 , n4825 , n4826 );
buf ( n50601 , n4827 );
buf ( n4829 , n50601 );
buf ( n50603 , n4829 );
buf ( n50604 , n50603 );
not ( n4832 , n50604 );
buf ( n50606 , n4832 );
buf ( n50607 , n50606 );
and ( n4835 , n4408 , n45336 );
not ( n4836 , n4835 );
not ( n4837 , n4404 );
or ( n4838 , n4836 , n4837 );
not ( n4839 , n49882 );
not ( n4840 , n45370 );
and ( n4841 , n4839 , n4840 );
nor ( n4842 , n4841 , n45369 );
nand ( n4843 , n4838 , n4842 );
buf ( n50617 , n4843 );
buf ( n50618 , n4102 );
buf ( n50619 , n45488 );
nand ( n4847 , n50618 , n50619 );
buf ( n50621 , n4847 );
buf ( n50622 , n50621 );
not ( n4850 , n50622 );
buf ( n50624 , n4850 );
buf ( n50625 , n50624 );
and ( n4853 , n50617 , n50625 );
not ( n4854 , n50617 );
buf ( n50628 , n50621 );
and ( n4856 , n4854 , n50628 );
nor ( n4857 , n4853 , n4856 );
buf ( n50631 , n4857 );
buf ( n50632 , n50631 );
not ( n4860 , n50632 );
buf ( n50634 , n4860 );
buf ( n50635 , n50634 );
not ( n4863 , n50635 );
buf ( n50637 , n4863 );
buf ( n50638 , n50637 );
buf ( n50639 , n378 );
nand ( n4867 , n50638 , n50639 );
buf ( n50641 , n4867 );
xor ( n4869 , n384 , n4426 );
xor ( n4870 , n4869 , n4439 );
nand ( n4871 , n50641 , n4870 );
not ( n4872 , n4871 );
buf ( n50646 , n3651 );
not ( n4874 , n50646 );
buf ( n50648 , n50225 );
not ( n4876 , n50648 );
or ( n4877 , n4874 , n4876 );
and ( n4878 , n4419 , n3654 );
not ( n4879 , n4419 );
and ( n4880 , n4879 , n378 );
nor ( n4881 , n4878 , n4880 );
buf ( n4882 , n4415 );
not ( n4883 , n4882 );
and ( n4884 , n4881 , n4883 );
not ( n4885 , n4881 );
and ( n4886 , n4885 , n4882 );
nor ( n4887 , n4884 , n4886 );
nand ( n4888 , n4887 , n49447 );
buf ( n50662 , n4888 );
nand ( n4890 , n4877 , n50662 );
buf ( n50664 , n4890 );
not ( n4892 , n50664 );
or ( n4893 , n4872 , n4892 );
or ( n4894 , n4870 , n50641 );
nand ( n4895 , n4893 , n4894 );
not ( n4896 , n4895 );
buf ( n50670 , n4896 );
nand ( n4898 , n50607 , n50670 );
buf ( n50672 , n4898 );
buf ( n50673 , n50672 );
not ( n4901 , n50673 );
or ( n4902 , n4816 , n4901 );
not ( n4903 , n4871 );
not ( n4904 , n50664 );
or ( n4905 , n4903 , n4904 );
nand ( n4906 , n4905 , n4894 );
nand ( n4907 , n50603 , n4906 );
buf ( n50681 , n4907 );
nand ( n4909 , n4902 , n50681 );
buf ( n50683 , n4909 );
buf ( n50684 , n50683 );
not ( n4912 , n50684 );
buf ( n50686 , n4912 );
buf ( n50687 , n50686 );
not ( n4915 , n50687 );
or ( n4916 , n4757 , n4915 );
xor ( n4917 , n50239 , n50243 );
xor ( n4918 , n4917 , n50294 );
buf ( n50692 , n4918 );
buf ( n50693 , n50692 );
buf ( n4921 , n50693 );
buf ( n50695 , n4921 );
buf ( n50696 , n50695 );
nand ( n4924 , n4916 , n50696 );
buf ( n50698 , n4924 );
buf ( n50699 , n50698 );
buf ( n50700 , n50528 );
not ( n4928 , n50700 );
buf ( n50702 , n50683 );
nand ( n4930 , n4928 , n50702 );
buf ( n50704 , n4930 );
buf ( n50705 , n50704 );
and ( n4933 , n50699 , n50705 );
buf ( n50707 , n4933 );
buf ( n50708 , n50371 );
buf ( n50709 , n50298 );
xor ( n4937 , n50708 , n50709 );
buf ( n50711 , n4384 );
xnor ( n4939 , n4937 , n50711 );
buf ( n50713 , n4939 );
nand ( n4941 , n50707 , n50713 );
buf ( n50715 , n4941 );
nand ( n4943 , n50522 , n50715 );
buf ( n50717 , n4943 );
nor ( n4945 , n4727 , n50717 );
not ( n4946 , n4945 );
xor ( n4947 , n4773 , n50581 );
xnor ( n4948 , n4947 , n4784 );
nand ( n4949 , n4408 , n45370 );
not ( n4950 , n4949 );
not ( n4951 , n4950 );
not ( n4952 , n4404 );
not ( n4953 , n4952 );
or ( n4954 , n4951 , n4953 );
nand ( n4955 , n4404 , n4949 );
nand ( n4956 , n4954 , n4955 );
buf ( n50730 , n4956 );
buf ( n50731 , n378 );
and ( n4959 , n50730 , n50731 );
buf ( n50733 , n4959 );
buf ( n50734 , n50733 );
and ( n4962 , n49346 , n48752 );
buf ( n50736 , n48797 );
not ( n4964 , n50736 );
buf ( n50738 , n2684 );
buf ( n4966 , n50738 );
buf ( n50740 , n4966 );
buf ( n50741 , n50740 );
not ( n4969 , n50741 );
or ( n4970 , n4964 , n4969 );
buf ( n50744 , n49330 );
buf ( n4972 , n50744 );
buf ( n50746 , n4972 );
buf ( n50747 , n50746 );
nand ( n4975 , n4970 , n50747 );
buf ( n50749 , n4975 );
xor ( n4977 , n4962 , n50749 );
buf ( n50751 , n4977 );
xor ( n4979 , n50734 , n50751 );
and ( n4980 , n50746 , n48797 );
xor ( n4981 , n4980 , n50740 );
nand ( n4982 , n42624 , n42641 , n42682 );
and ( n4983 , n4981 , n4982 );
buf ( n50757 , n4983 );
xor ( n4985 , n4979 , n50757 );
buf ( n50759 , n4985 );
buf ( n50760 , n50759 );
buf ( n50761 , n3716 );
not ( n4989 , n50761 );
not ( n4990 , n382 );
not ( n4991 , n50125 );
or ( n4992 , n4990 , n4991 );
nand ( n4993 , n4349 , n49395 );
nand ( n4994 , n4992 , n4993 );
buf ( n50768 , n4994 );
not ( n4996 , n50768 );
or ( n4997 , n4989 , n4996 );
buf ( n50771 , n382 );
buf ( n50772 , n50571 );
and ( n5000 , n50771 , n50772 );
not ( n5001 , n50771 );
buf ( n50775 , n4369 );
and ( n5003 , n5001 , n50775 );
nor ( n5004 , n5000 , n5003 );
buf ( n50778 , n5004 );
not ( n5006 , n50778 );
nand ( n5007 , n5006 , n3733 );
buf ( n50781 , n5007 );
nand ( n5009 , n4997 , n50781 );
buf ( n50783 , n5009 );
buf ( n50784 , n50783 );
xor ( n5012 , n50760 , n50784 );
buf ( n50786 , n49447 );
not ( n5014 , n50786 );
buf ( n50788 , n378 );
buf ( n50789 , n4956 );
and ( n5017 , n50788 , n50789 );
not ( n5018 , n50788 );
buf ( n50792 , n4956 );
not ( n5020 , n50792 );
buf ( n50794 , n5020 );
buf ( n50795 , n50794 );
and ( n5023 , n5018 , n50795 );
nor ( n5024 , n5017 , n5023 );
buf ( n50798 , n5024 );
buf ( n50799 , n50798 );
not ( n5027 , n50799 );
or ( n5028 , n5014 , n5027 );
buf ( n50802 , n378 );
not ( n5030 , n50802 );
buf ( n50804 , n50537 );
not ( n5032 , n50804 );
or ( n5033 , n5030 , n5032 );
buf ( n50807 , n3654 );
buf ( n50808 , n50534 );
nand ( n5036 , n50807 , n50808 );
buf ( n50810 , n5036 );
buf ( n50811 , n50810 );
nand ( n5039 , n5033 , n50811 );
buf ( n50813 , n5039 );
buf ( n50814 , n50813 );
buf ( n50815 , n3651 );
nand ( n5043 , n50814 , n50815 );
buf ( n50817 , n5043 );
buf ( n50818 , n50817 );
nand ( n5046 , n5028 , n50818 );
buf ( n50820 , n5046 );
not ( n5048 , n50820 );
buf ( n50822 , n380 );
not ( n5050 , n50822 );
buf ( n50824 , n4421 );
not ( n5052 , n50824 );
buf ( n50826 , n5052 );
buf ( n50827 , n50826 );
not ( n5055 , n50827 );
or ( n5056 , n5050 , n5055 );
buf ( n50830 , n4421 );
buf ( n50831 , n3609 );
nand ( n5059 , n50830 , n50831 );
buf ( n50833 , n5059 );
buf ( n50834 , n50833 );
nand ( n5062 , n5056 , n50834 );
buf ( n50836 , n5062 );
nand ( n5064 , n50836 , n3622 );
not ( n5065 , n3609 );
and ( n5066 , n4843 , n50621 );
not ( n5067 , n4843 );
and ( n5068 , n5067 , n50624 );
nor ( n5069 , n5066 , n5068 );
not ( n5070 , n5069 );
not ( n5071 , n5070 );
or ( n5072 , n5065 , n5071 );
or ( n5073 , n3609 , n5070 );
nand ( n5074 , n5072 , n5073 );
nand ( n5075 , n5074 , n3620 );
nand ( n5076 , n5048 , n5064 , n5075 );
not ( n5077 , n5076 );
buf ( n50851 , n382 );
not ( n5079 , n50851 );
buf ( n50853 , n4224 );
not ( n5081 , n50853 );
or ( n5082 , n5079 , n5081 );
buf ( n50856 , n49998 );
buf ( n50857 , n49395 );
nand ( n5085 , n50856 , n50857 );
buf ( n50859 , n5085 );
buf ( n50860 , n50859 );
nand ( n5088 , n5082 , n50860 );
buf ( n50862 , n5088 );
not ( n5090 , n50862 );
not ( n5091 , n3733 );
or ( n5092 , n5090 , n5091 );
or ( n5093 , n50778 , n49496 );
nand ( n5094 , n5092 , n5093 );
not ( n5095 , n5094 );
or ( n5096 , n5077 , n5095 );
not ( n5097 , n5075 );
not ( n5098 , n5064 );
or ( n5099 , n5097 , n5098 );
nand ( n5100 , n5099 , n50820 );
nand ( n5101 , n5096 , n5100 );
buf ( n50875 , n5101 );
and ( n5103 , n5012 , n50875 );
and ( n5104 , n50760 , n50784 );
or ( n5105 , n5103 , n5104 );
buf ( n50879 , n5105 );
not ( n5107 , n50879 );
nand ( n5108 , n50540 , n378 );
not ( n5109 , n4772 );
and ( n5110 , n5108 , n5109 );
not ( n5111 , n5108 );
and ( n5112 , n5111 , n4772 );
nor ( n5113 , n5110 , n5112 );
not ( n5114 , n49447 );
not ( n5115 , n378 );
not ( n5116 , n5069 );
or ( n5117 , n5115 , n5116 );
buf ( n50891 , n50631 );
buf ( n50892 , n3654 );
nand ( n5120 , n50891 , n50892 );
buf ( n50894 , n5120 );
nand ( n5122 , n5117 , n50894 );
not ( n5123 , n5122 );
or ( n5124 , n5114 , n5123 );
nand ( n5125 , n4887 , n3651 );
nand ( n5126 , n5124 , n5125 );
xor ( n5127 , n5113 , n5126 );
xor ( n5128 , n49992 , n380 );
not ( n5129 , n49968 );
not ( n5130 , n49972 );
and ( n5131 , n5129 , n5130 );
and ( n5132 , n49976 , n4216 );
nor ( n50906 , n5131 , n5132 );
xnor ( n5134 , n5128 , n50906 );
not ( n50908 , n5134 );
not ( n5136 , n3620 );
or ( n50910 , n50908 , n5136 );
not ( n5138 , n4799 );
not ( n50912 , n4802 );
or ( n5140 , n5138 , n50912 );
nand ( n50914 , n5140 , n3622 );
nand ( n5142 , n50910 , n50914 );
xor ( n50916 , n5127 , n5142 );
not ( n5144 , n50916 );
not ( n50918 , n50836 );
not ( n5146 , n3620 );
or ( n50920 , n50918 , n5146 );
nand ( n5148 , n5134 , n3622 );
nand ( n50922 , n50920 , n5148 );
not ( n5150 , n50922 );
nand ( n50924 , n4038 , n45377 );
not ( n5152 , n50924 );
not ( n50926 , n50170 );
nand ( n5154 , n44829 , n44688 );
nand ( n50928 , n50926 , n5154 );
not ( n5156 , n50928 );
or ( n50930 , n5152 , n5156 );
not ( n5158 , n50924 );
not ( n50932 , n5154 );
nor ( n5160 , n50932 , n50170 );
nand ( n50934 , n5158 , n5160 );
nand ( n5162 , n50930 , n50934 );
and ( n50936 , n378 , n5162 );
not ( n5164 , n50936 );
not ( n50938 , n5164 );
buf ( n50939 , n2464 );
buf ( n50940 , n50939 );
buf ( n50941 , n50940 );
buf ( n50942 , n50941 );
not ( n5170 , n50942 );
buf ( n50944 , n2486 );
not ( n5172 , n50944 );
buf ( n50946 , n5172 );
buf ( n50947 , n50946 );
not ( n50948 , n50947 );
buf ( n50949 , n47869 );
not ( n5177 , n50949 );
or ( n50951 , n50948 , n5177 );
buf ( n50952 , n2658 );
not ( n50953 , n50952 );
buf ( n50954 , n50953 );
buf ( n50955 , n50954 );
nand ( n50956 , n50951 , n50955 );
buf ( n50957 , n50956 );
buf ( n50958 , n50957 );
not ( n50959 , n50958 );
or ( n50960 , n5170 , n50959 );
buf ( n50961 , n48467 );
not ( n50962 , n50961 );
buf ( n50963 , n50962 );
buf ( n50964 , n50963 );
not ( n50965 , n50964 );
buf ( n50966 , n50965 );
buf ( n50967 , n50966 );
nand ( n50968 , n50960 , n50967 );
buf ( n50969 , n50968 );
buf ( n50970 , n2677 );
buf ( n50971 , n48457 );
nand ( n50972 , n50970 , n50971 );
buf ( n50973 , n50972 );
not ( n50974 , n50973 );
and ( n50975 , n50969 , n50974 );
not ( n50976 , n50969 );
and ( n50977 , n50976 , n50973 );
nor ( n50978 , n50975 , n50977 );
nand ( n50979 , n45380 , n3992 );
not ( n50980 , n50979 );
not ( n50981 , n4001 );
or ( n50982 , n50980 , n50981 );
nand ( n50983 , n45381 , n4035 , n50979 );
nand ( n50984 , n50982 , n50983 );
not ( n50985 , n44525 );
not ( n50986 , n50985 );
not ( n50987 , n44683 );
not ( n50988 , n50987 );
or ( n50989 , n50986 , n50988 );
nand ( n50990 , n50989 , n45377 );
not ( n50991 , n50990 );
and ( n50992 , n50984 , n50991 );
not ( n50993 , n50984 );
not ( n50994 , n50985 );
not ( n50995 , n50987 );
or ( n50996 , n50994 , n50995 );
nand ( n50997 , n50996 , n45377 );
and ( n50998 , n50993 , n50997 );
nor ( n50999 , n50992 , n50998 );
nand ( n51000 , n50999 , n378 );
not ( n51001 , n51000 );
nand ( n51002 , n50978 , n51001 );
not ( n51003 , n51002 );
or ( n51004 , n50938 , n51003 );
xor ( n51005 , n4981 , n4982 );
nand ( n51006 , n51004 , n51005 );
not ( n51007 , n51002 );
nand ( n51008 , n51007 , n50936 );
nand ( n51009 , n51006 , n51008 );
not ( n51010 , n51009 );
not ( n51011 , n3651 );
not ( n51012 , n5122 );
or ( n51013 , n51011 , n51012 );
nand ( n51014 , n50813 , n49447 );
nand ( n51015 , n51013 , n51014 );
not ( n51016 , n51015 );
nand ( n51017 , n51010 , n51016 );
not ( n51018 , n51017 );
or ( n51019 , n5150 , n51018 );
nand ( n51020 , n51015 , n51009 );
nand ( n51021 , n51019 , n51020 );
buf ( n51022 , n51021 );
not ( n51023 , n51022 );
buf ( n51024 , n51023 );
nand ( n51025 , n5144 , n51024 );
not ( n51026 , n51025 );
or ( n51027 , n5107 , n51026 );
buf ( n51028 , n5144 );
not ( n51029 , n51028 );
buf ( n51030 , n51029 );
buf ( n51031 , n51030 );
buf ( n51032 , n51021 );
nand ( n51033 , n51031 , n51032 );
buf ( n51034 , n51033 );
nand ( n51035 , n51027 , n51034 );
xor ( n51036 , n4948 , n51035 );
xor ( n51037 , n5113 , n5126 );
and ( n51038 , n51037 , n5142 );
and ( n51039 , n5113 , n5126 );
or ( n51040 , n51038 , n51039 );
buf ( n51041 , n51040 );
not ( n51042 , n51041 );
buf ( n51043 , n50641 );
buf ( n51044 , n4870 );
xor ( n51045 , n51043 , n51044 );
buf ( n51046 , n50664 );
xnor ( n51047 , n51045 , n51046 );
buf ( n51048 , n51047 );
buf ( n51049 , n51048 );
not ( n51050 , n51049 );
or ( n51051 , n51042 , n51050 );
buf ( n51052 , n51048 );
buf ( n51053 , n51040 );
or ( n51054 , n51052 , n51053 );
nand ( n51055 , n51051 , n51054 );
buf ( n51056 , n51055 );
not ( n51057 , n3733 );
not ( n51058 , n4994 );
or ( n51059 , n51057 , n51058 );
xor ( n51060 , n4124 , n382 );
xnor ( n51061 , n51060 , n4122 );
nand ( n51062 , n51061 , n3716 );
nand ( n51063 , n51059 , n51062 );
not ( n51064 , n51063 );
not ( n51065 , n385 );
and ( n51066 , n51065 , n384 );
buf ( n51067 , n51066 );
not ( n51068 , n51067 );
buf ( n51069 , n4076 );
not ( n51070 , n51069 );
or ( n51071 , n51068 , n51070 );
buf ( n51072 , n384 );
buf ( n51073 , n385 );
nand ( n51074 , n51072 , n51073 );
buf ( n51075 , n51074 );
buf ( n51076 , n51075 );
nand ( n51077 , n51071 , n51076 );
buf ( n51078 , n51077 );
not ( n51079 , n51078 );
or ( n51080 , n51064 , n51079 );
buf ( n51081 , n51078 );
not ( n51082 , n51081 );
buf ( n51083 , n51082 );
nand ( n51084 , n3733 , n4994 );
and ( n51085 , n51083 , n51084 , n51062 );
xor ( n51086 , n50734 , n50751 );
and ( n51087 , n51086 , n50757 );
and ( n51088 , n50734 , n50751 );
or ( n51089 , n51087 , n51088 );
buf ( n51090 , n51089 );
buf ( n51091 , n51090 );
not ( n51092 , n51091 );
buf ( n51093 , n51092 );
or ( n51094 , n51085 , n51093 );
nand ( n51095 , n51080 , n51094 );
and ( n51096 , n51056 , n51095 );
not ( n51097 , n51056 );
not ( n51098 , n51095 );
and ( n51099 , n51097 , n51098 );
nor ( n51100 , n51096 , n51099 );
xor ( n51101 , n51036 , n51100 );
buf ( n51102 , n51101 );
not ( n51103 , n51102 );
buf ( n51104 , n51103 );
and ( n51105 , n51093 , n51083 );
not ( n51106 , n51093 );
and ( n51107 , n51106 , n51078 );
nor ( n51108 , n51105 , n51107 );
not ( n51109 , n51108 );
not ( n51110 , n51063 );
and ( n51111 , n51109 , n51110 );
and ( n51112 , n51108 , n51063 );
nor ( n51113 , n51111 , n51112 );
buf ( n51114 , n51066 );
not ( n51115 , n51114 );
and ( n51116 , n384 , n4130 );
not ( n51117 , n384 );
and ( n51118 , n51117 , n4129 );
or ( n51119 , n51116 , n51118 );
buf ( n51120 , n51119 );
not ( n51121 , n51120 );
or ( n51122 , n51115 , n51121 );
buf ( n51123 , n384 );
buf ( n51124 , n4054 );
and ( n51125 , n51123 , n51124 );
not ( n51126 , n51123 );
buf ( n51127 , n4076 );
and ( n51128 , n51126 , n51127 );
nor ( n51129 , n51125 , n51128 );
buf ( n51130 , n51129 );
buf ( n51131 , n51130 );
buf ( n51132 , n385 );
nand ( n51133 , n51131 , n51132 );
buf ( n51134 , n51133 );
buf ( n51135 , n51134 );
nand ( n51136 , n51122 , n51135 );
buf ( n51137 , n51136 );
not ( n51138 , n51137 );
and ( n51139 , n51015 , n51009 );
not ( n51140 , n51015 );
and ( n51141 , n51140 , n51010 );
nor ( n51142 , n51139 , n51141 );
not ( n51143 , n50922 );
and ( n51144 , n51142 , n51143 );
not ( n51145 , n51142 );
and ( n51146 , n51145 , n50922 );
nor ( n51147 , n51144 , n51146 );
buf ( n51148 , n51147 );
not ( n51149 , n51148 );
buf ( n51150 , n51149 );
not ( n51151 , n51150 );
or ( n51152 , n51138 , n51151 );
buf ( n51153 , n51150 );
buf ( n51154 , n51137 );
or ( n51155 , n51153 , n51154 );
xor ( n51156 , n5164 , n51007 );
xnor ( n51157 , n51156 , n51005 );
not ( n51158 , n51157 );
buf ( n51159 , n50963 );
not ( n51160 , n51159 );
buf ( n51161 , n50941 );
nand ( n51162 , n51160 , n51161 );
buf ( n51163 , n51162 );
xnor ( n51164 , n50957 , n51163 );
buf ( n51165 , n51164 );
nand ( n51166 , n4036 , n45384 );
not ( n51167 , n44303 );
not ( n51168 , n44520 );
or ( n51169 , n51167 , n51168 );
nand ( n51170 , n51169 , n50979 );
not ( n51171 , n51170 );
and ( n51172 , n51166 , n51171 );
not ( n51173 , n51166 );
and ( n51174 , n51173 , n51170 );
nor ( n51175 , n51172 , n51174 );
and ( n51176 , n51175 , n378 );
buf ( n51177 , n51176 );
and ( n51178 , n51165 , n51177 );
buf ( n51179 , n51178 );
buf ( n51180 , n51179 );
not ( n51181 , n51180 );
nand ( n51182 , n42675 , n40664 );
not ( n51183 , n51182 );
nand ( n51184 , n42637 , n42686 );
nand ( n51185 , n51184 , n42439 );
not ( n51186 , n51185 );
or ( n51187 , n51183 , n51186 );
not ( n51188 , n51182 );
nand ( n51189 , n51188 , n42439 , n51184 );
nand ( n51190 , n51187 , n51189 );
buf ( n51191 , n51190 );
not ( n51192 , n51191 );
or ( n51193 , n51181 , n51192 );
not ( n51194 , n51179 );
not ( n51195 , n51194 );
not ( n51196 , n51190 );
not ( n51197 , n51196 );
or ( n51198 , n51195 , n51197 );
buf ( n51199 , n50978 );
buf ( n51200 , n51000 );
and ( n51201 , n51199 , n51200 );
not ( n51202 , n51199 );
buf ( n51203 , n51001 );
and ( n51204 , n51202 , n51203 );
nor ( n51205 , n51201 , n51204 );
buf ( n51206 , n51205 );
buf ( n51207 , n51206 );
not ( n51208 , n51207 );
buf ( n51209 , n51208 );
nand ( n51210 , n51198 , n51209 );
buf ( n51211 , n51210 );
nand ( n51212 , n51193 , n51211 );
buf ( n51213 , n51212 );
buf ( n51214 , n51213 );
not ( n51215 , n51214 );
buf ( n51216 , n51215 );
nand ( n51217 , n51158 , n51216 );
not ( n51218 , n51217 );
not ( n51219 , n3651 );
not ( n51220 , n50798 );
or ( n51221 , n51219 , n51220 );
xor ( n51222 , n378 , n5162 );
buf ( n51223 , n51222 );
buf ( n51224 , n49447 );
nand ( n51225 , n51223 , n51224 );
buf ( n51226 , n51225 );
nand ( n51227 , n51221 , n51226 );
not ( n51228 , n51227 );
not ( n51229 , n51228 );
buf ( n51230 , n3651 );
not ( n51231 , n51230 );
buf ( n51232 , n51222 );
not ( n51233 , n51232 );
or ( n51234 , n51231 , n51233 );
xor ( n51235 , n378 , n50997 );
xnor ( n51236 , n51235 , n50984 );
buf ( n51237 , n51236 );
buf ( n51238 , n49447 );
nand ( n51239 , n51237 , n51238 );
buf ( n51240 , n51239 );
buf ( n51241 , n51240 );
nand ( n51242 , n51234 , n51241 );
buf ( n51243 , n51242 );
not ( n51244 , n51243 );
buf ( n51245 , n51176 );
buf ( n51246 , n51164 );
not ( n51247 , n51246 );
buf ( n51248 , n51247 );
buf ( n51249 , n51248 );
and ( n51250 , n51245 , n51249 );
not ( n51251 , n51245 );
buf ( n51252 , n51164 );
and ( n51253 , n51251 , n51252 );
nor ( n51254 , n51250 , n51253 );
buf ( n51255 , n51254 );
buf ( n51256 , n51255 );
xor ( n51257 , n43887 , n44090 );
not ( n51258 , n4028 );
nand ( n51259 , n4023 , n43882 );
nand ( n51260 , n51258 , n51259 );
xor ( n51261 , n51257 , n51260 );
buf ( n51262 , n51261 );
buf ( n51263 , n51262 );
buf ( n51264 , n51263 );
nand ( n51265 , n51264 , n378 );
not ( n51266 , n51265 );
not ( n51267 , n47862 );
nor ( n51268 , n51267 , n47841 );
not ( n51269 , n51268 );
buf ( n51270 , n47850 );
not ( n51271 , n51270 );
buf ( n51272 , n51271 );
and ( n51273 , n51272 , n47208 );
not ( n51274 , n51273 );
or ( n51275 , n51269 , n51274 );
not ( n51276 , n47841 );
not ( n51277 , n51276 );
not ( n51278 , n51272 );
or ( n51279 , n51277 , n51278 );
nand ( n51280 , n47208 , n47862 );
nand ( n51281 , n51279 , n51280 );
nand ( n51282 , n51275 , n51281 );
nand ( n51283 , n51266 , n51282 );
buf ( n51284 , n51283 );
not ( n51285 , n51284 );
buf ( n51286 , n50954 );
buf ( n51287 , n50946 );
nand ( n51288 , n51286 , n51287 );
buf ( n51289 , n51288 );
buf ( n51290 , n51289 );
not ( n51291 , n51290 );
buf ( n51292 , n47208 );
not ( n51293 , n51292 );
buf ( n51294 , n47841 );
not ( n51295 , n51294 );
or ( n51296 , n51293 , n51295 );
buf ( n51297 , n47866 );
nand ( n51298 , n51296 , n51297 );
buf ( n51299 , n51298 );
buf ( n51300 , n51299 );
not ( n51301 , n51300 );
or ( n51302 , n51291 , n51301 );
buf ( n51303 , n51299 );
buf ( n51304 , n51289 );
or ( n51305 , n51303 , n51304 );
buf ( n51306 , n51305 );
buf ( n51307 , n51306 );
nand ( n51308 , n51302 , n51307 );
buf ( n51309 , n51308 );
buf ( n51310 , n51309 );
nand ( n51311 , n51285 , n51310 );
buf ( n51312 , n51311 );
buf ( n51313 , n51312 );
nand ( n51314 , n51256 , n51313 );
buf ( n51315 , n51314 );
not ( n51316 , n51315 );
or ( n51317 , n51244 , n51316 );
buf ( n51318 , n51312 );
not ( n51319 , n51318 );
buf ( n51320 , n51255 );
not ( n51321 , n51320 );
buf ( n51322 , n51321 );
buf ( n51323 , n51322 );
nand ( n5199 , n51319 , n51323 );
buf ( n51325 , n5199 );
nand ( n5201 , n51317 , n51325 );
buf ( n5202 , n5201 );
or ( n5203 , n51229 , n5202 );
not ( n5204 , n3622 );
not ( n5205 , n5074 );
or ( n5206 , n5204 , n5205 );
and ( n5207 , n50534 , n3609 );
not ( n5208 , n50534 );
and ( n5209 , n5208 , n380 );
or ( n5210 , n5207 , n5209 );
nand ( n5211 , n5210 , n3620 );
nand ( n5212 , n5206 , n5211 );
nand ( n5213 , n5203 , n5212 );
nand ( n5214 , n5202 , n51229 );
nand ( n5215 , n5213 , n5214 );
not ( n5216 , n5215 );
or ( n5217 , n51218 , n5216 );
nand ( n5218 , n51213 , n51157 );
nand ( n5219 , n5217 , n5218 );
buf ( n51345 , n5219 );
nand ( n5221 , n51155 , n51345 );
buf ( n51347 , n5221 );
nand ( n5223 , n51152 , n51347 );
xor ( n5224 , n51113 , n5223 );
and ( n5225 , n50916 , n51021 );
not ( n5226 , n50916 );
and ( n5227 , n5226 , n51024 );
nor ( n5228 , n5225 , n5227 );
and ( n5229 , n50879 , n5228 );
not ( n5230 , n50879 );
not ( n5231 , n5228 );
and ( n5232 , n5230 , n5231 );
nor ( n5233 , n5229 , n5232 );
and ( n5234 , n5224 , n5233 );
and ( n5235 , n51113 , n5223 );
or ( n5236 , n5234 , n5235 );
not ( n5237 , n5236 );
nand ( n5238 , n51104 , n5237 );
xor ( n5239 , n51113 , n5223 );
xor ( n5240 , n5239 , n5233 );
not ( n5241 , n5240 );
not ( n5242 , n51147 );
not ( n5243 , n5242 );
buf ( n51369 , n51137 );
not ( n5245 , n51369 );
buf ( n51371 , n5245 );
not ( n5247 , n51371 );
or ( n5248 , n5243 , n5247 );
buf ( n51374 , n51137 );
buf ( n51375 , n51147 );
nand ( n5251 , n51374 , n51375 );
buf ( n51377 , n5251 );
nand ( n5253 , n5248 , n51377 );
buf ( n51379 , n5219 );
not ( n5255 , n51379 );
buf ( n51381 , n5255 );
and ( n5257 , n5253 , n51381 );
not ( n5258 , n5253 );
and ( n5259 , n5258 , n5219 );
nor ( n5260 , n5257 , n5259 );
buf ( n51386 , n5260 );
xor ( n5262 , n50760 , n50784 );
xor ( n5263 , n5262 , n50875 );
buf ( n51389 , n5263 );
buf ( n51390 , n51389 );
not ( n5266 , n51390 );
buf ( n51392 , n5266 );
buf ( n51393 , n51392 );
nand ( n5269 , n51386 , n51393 );
buf ( n51395 , n5269 );
not ( n5271 , n51395 );
buf ( n51397 , n385 );
not ( n5273 , n51397 );
buf ( n51399 , n51119 );
not ( n5275 , n51399 );
or ( n5276 , n5273 , n5275 );
not ( n5277 , n384 );
not ( n5278 , n50125 );
or ( n5279 , n5277 , n5278 );
not ( n5280 , n384 );
nand ( n5281 , n5280 , n4349 );
nand ( n5282 , n5279 , n5281 );
buf ( n51408 , n5282 );
buf ( n51409 , n51066 );
nand ( n5285 , n51408 , n51409 );
buf ( n51411 , n5285 );
buf ( n51412 , n51411 );
nand ( n5288 , n5276 , n51412 );
buf ( n51414 , n5288 );
buf ( n51415 , n3716 );
not ( n5291 , n51415 );
buf ( n51417 , n50862 );
not ( n5293 , n51417 );
or ( n5294 , n5291 , n5293 );
not ( n5295 , n49395 );
not ( n5296 , n4392 );
not ( n5297 , n4415 );
or ( n5298 , n5296 , n5297 );
nand ( n5299 , n5298 , n4420 );
not ( n5300 , n5299 );
or ( n5301 , n5295 , n5300 );
or ( n5302 , n49395 , n4421 );
nand ( n5303 , n5301 , n5302 );
buf ( n51429 , n5303 );
buf ( n51430 , n3733 );
nand ( n5306 , n51429 , n51430 );
buf ( n51432 , n5306 );
buf ( n51433 , n51432 );
nand ( n5309 , n5294 , n51433 );
buf ( n51435 , n5309 );
not ( n5311 , n51435 );
buf ( n51437 , n51179 );
buf ( n51438 , n51190 );
xor ( n5314 , n51437 , n51438 );
buf ( n51440 , n51206 );
xor ( n5316 , n5314 , n51440 );
buf ( n51442 , n5316 );
not ( n5318 , n51442 );
not ( n5319 , n5318 );
or ( n5320 , n5311 , n5319 );
not ( n5321 , n51442 );
not ( n5322 , n51432 );
and ( n5323 , n3716 , n50862 );
nor ( n5324 , n5322 , n5323 );
not ( n5325 , n5324 );
or ( n5326 , n5321 , n5325 );
not ( n5327 , n42637 );
not ( n5328 , n42690 );
or ( n5329 , n5327 , n5328 );
nand ( n5330 , n5329 , n42498 );
buf ( n51456 , n42146 );
not ( n5332 , n51456 );
buf ( n51458 , n42152 );
nand ( n5334 , n5332 , n51458 );
buf ( n51460 , n5334 );
buf ( n51461 , n51460 );
not ( n5337 , n51461 );
buf ( n51463 , n5337 );
and ( n5339 , n5330 , n51463 );
not ( n5340 , n5330 );
and ( n5341 , n5340 , n51460 );
nor ( n5342 , n5339 , n5341 );
not ( n5343 , n5342 );
buf ( n51469 , n3620 );
not ( n5345 , n51469 );
not ( n5346 , n3609 );
not ( n5347 , n4956 );
or ( n5348 , n5346 , n5347 );
nand ( n5349 , n380 , n50794 );
nand ( n5350 , n5348 , n5349 );
buf ( n51476 , n5350 );
not ( n5352 , n51476 );
or ( n5353 , n5345 , n5352 );
buf ( n51479 , n5210 );
buf ( n51480 , n3622 );
nand ( n5356 , n51479 , n51480 );
buf ( n51482 , n5356 );
buf ( n51483 , n51482 );
nand ( n5359 , n5353 , n51483 );
buf ( n51485 , n5359 );
not ( n5361 , n51485 );
or ( n5362 , n5343 , n5361 );
buf ( n51488 , n51485 );
buf ( n51489 , n5330 );
buf ( n51490 , n51463 );
and ( n5366 , n51489 , n51490 );
not ( n5367 , n51489 );
buf ( n51493 , n51460 );
and ( n5369 , n5367 , n51493 );
nor ( n5370 , n5366 , n5369 );
buf ( n51496 , n5370 );
buf ( n51497 , n51496 );
or ( n5373 , n51488 , n51497 );
buf ( n51499 , n378 );
not ( n5375 , n4035 );
and ( n5376 , n5375 , n45387 );
not ( n5377 , n5375 );
not ( n5378 , n45387 );
and ( n5379 , n5377 , n5378 );
nor ( n5380 , n5376 , n5379 );
buf ( n51506 , n5380 );
and ( n5382 , n51499 , n51506 );
buf ( n51508 , n5382 );
buf ( n51509 , n51508 );
buf ( n51510 , n51283 );
not ( n5386 , n51510 );
buf ( n51512 , n51309 );
not ( n5388 , n51512 );
or ( n5389 , n5386 , n5388 );
buf ( n51515 , n51309 );
buf ( n51516 , n51283 );
or ( n5392 , n51515 , n51516 );
nand ( n5393 , n5389 , n5392 );
buf ( n51519 , n5393 );
buf ( n51520 , n51519 );
xor ( n5396 , n51509 , n51520 );
buf ( n51522 , n3651 );
not ( n5398 , n51522 );
buf ( n51524 , n51236 );
not ( n5400 , n51524 );
or ( n5401 , n5398 , n5400 );
buf ( n51527 , n378 );
not ( n5403 , n51527 );
buf ( n51529 , n51175 );
not ( n5405 , n51529 );
buf ( n51531 , n5405 );
buf ( n51532 , n51531 );
not ( n5408 , n51532 );
or ( n5409 , n5403 , n5408 );
buf ( n51535 , n51175 );
buf ( n51536 , n3654 );
nand ( n5412 , n51535 , n51536 );
buf ( n51538 , n5412 );
buf ( n51539 , n51538 );
nand ( n5415 , n5409 , n51539 );
buf ( n51541 , n5415 );
buf ( n51542 , n51541 );
buf ( n51543 , n49447 );
nand ( n5419 , n51542 , n51543 );
buf ( n51545 , n5419 );
buf ( n51546 , n51545 );
nand ( n5422 , n5401 , n51546 );
buf ( n51548 , n5422 );
buf ( n51549 , n51548 );
and ( n5425 , n5396 , n51549 );
and ( n5426 , n51509 , n51520 );
or ( n5427 , n5425 , n5426 );
buf ( n51553 , n5427 );
buf ( n51554 , n51553 );
nand ( n5430 , n5373 , n51554 );
buf ( n51556 , n5430 );
nand ( n5432 , n5362 , n51556 );
nand ( n5433 , n5326 , n5432 );
nand ( n5434 , n5320 , n5433 );
xor ( n5435 , n51414 , n5434 );
nand ( n5436 , n5075 , n5064 );
xor ( n5437 , n5048 , n5436 );
xnor ( n5438 , n5437 , n5094 );
and ( n5439 , n5435 , n5438 );
and ( n5440 , n51414 , n5434 );
or ( n5441 , n5439 , n5440 );
not ( n5442 , n5441 );
or ( n5443 , n5271 , n5442 );
not ( n5444 , n51392 );
buf ( n51570 , n5260 );
not ( n5446 , n51570 );
buf ( n51572 , n5446 );
nand ( n5448 , n5444 , n51572 );
nand ( n5449 , n5443 , n5448 );
buf ( n51575 , n5449 );
not ( n5451 , n51575 );
buf ( n51577 , n5451 );
nand ( n5453 , n5241 , n51577 );
and ( n5454 , n5238 , n5453 );
buf ( n51580 , n50528 );
buf ( n51581 , n50692 );
xor ( n5457 , n51580 , n51581 );
buf ( n51583 , n50683 );
xor ( n5459 , n5457 , n51583 );
buf ( n51585 , n5459 );
buf ( n51586 , n51585 );
xor ( n5462 , n50246 , n50265 );
xor ( n5463 , n5462 , n50289 );
buf ( n51589 , n5463 );
buf ( n51590 , n51589 );
not ( n5466 , n51590 );
buf ( n51592 , n50587 );
not ( n5468 , n51592 );
buf ( n51594 , n5468 );
buf ( n51595 , n51594 );
not ( n5471 , n51595 );
not ( n5472 , n4906 );
and ( n5473 , n5472 , n4827 );
not ( n5474 , n5472 );
not ( n5475 , n4827 );
and ( n5476 , n5474 , n5475 );
nor ( n5477 , n5473 , n5476 );
not ( n5478 , n5477 );
buf ( n51604 , n5478 );
not ( n5480 , n51604 );
or ( n5481 , n5471 , n5480 );
buf ( n51607 , n50587 );
buf ( n51608 , n5477 );
nand ( n5484 , n51607 , n51608 );
buf ( n51610 , n5484 );
buf ( n51611 , n51610 );
nand ( n5487 , n5481 , n51611 );
buf ( n51613 , n5487 );
buf ( n51614 , n51613 );
not ( n5490 , n51614 );
or ( n5491 , n5466 , n5490 );
buf ( n51617 , n51589 );
buf ( n51618 , n51594 );
not ( n5494 , n51618 );
buf ( n51620 , n5478 );
not ( n5496 , n51620 );
or ( n5497 , n5494 , n5496 );
buf ( n51623 , n51610 );
nand ( n5499 , n5497 , n51623 );
buf ( n51625 , n5499 );
buf ( n51626 , n51625 );
or ( n5502 , n51617 , n51626 );
buf ( n51628 , n51040 );
not ( n5504 , n51628 );
buf ( n51630 , n51048 );
nand ( n5506 , n5504 , n51630 );
buf ( n51632 , n5506 );
buf ( n51633 , n51632 );
not ( n5509 , n51633 );
buf ( n51635 , n51095 );
not ( n5511 , n51635 );
or ( n5512 , n5509 , n5511 );
buf ( n51638 , n51048 );
not ( n5514 , n51638 );
buf ( n51640 , n51040 );
nand ( n5516 , n5514 , n51640 );
buf ( n51642 , n5516 );
buf ( n51643 , n51642 );
nand ( n5519 , n5512 , n51643 );
buf ( n51645 , n5519 );
buf ( n51646 , n51645 );
nand ( n5522 , n5502 , n51646 );
buf ( n51648 , n5522 );
buf ( n51649 , n51648 );
nand ( n5525 , n5491 , n51649 );
buf ( n51651 , n5525 );
buf ( n51652 , n51651 );
not ( n5528 , n51652 );
buf ( n51654 , n5528 );
buf ( n51655 , n51654 );
nand ( n5531 , n51586 , n51655 );
buf ( n51657 , n5531 );
buf ( n51658 , n51657 );
xor ( n5534 , n51589 , n51613 );
xnor ( n5535 , n5534 , n51645 );
xor ( n5536 , n4948 , n51035 );
and ( n5537 , n5536 , n51100 );
and ( n5538 , n4948 , n51035 );
or ( n5539 , n5537 , n5538 );
buf ( n51665 , n5539 );
not ( n5541 , n51665 );
buf ( n51667 , n5541 );
nand ( n5543 , n5535 , n51667 );
buf ( n51669 , n5543 );
and ( n5545 , n51658 , n51669 );
buf ( n51671 , n5545 );
nand ( n5547 , n5454 , n51671 );
buf ( n51673 , n5547 );
not ( n5549 , n51673 );
buf ( n51675 , n5549 );
not ( n5551 , n51322 );
not ( n5552 , n51312 );
not ( n5553 , n5552 );
and ( n5554 , n5551 , n5553 );
and ( n5555 , n51322 , n5552 );
nor ( n5556 , n5554 , n5555 );
and ( n5557 , n5556 , n51243 );
not ( n5558 , n5556 );
not ( n5559 , n51243 );
and ( n5560 , n5558 , n5559 );
nor ( n5561 , n5557 , n5560 );
buf ( n51687 , n5561 );
buf ( n51688 , n3733 );
not ( n5564 , n51688 );
buf ( n51690 , n382 );
not ( n5566 , n51690 );
buf ( n51692 , n50634 );
not ( n5568 , n51692 );
or ( n5569 , n5566 , n5568 );
buf ( n51695 , n50637 );
buf ( n51696 , n49395 );
nand ( n5572 , n51695 , n51696 );
buf ( n51698 , n5572 );
buf ( n51699 , n51698 );
nand ( n5575 , n5569 , n51699 );
buf ( n51701 , n5575 );
buf ( n51702 , n51701 );
not ( n5578 , n51702 );
or ( n5579 , n5564 , n5578 );
buf ( n51705 , n5303 );
buf ( n51706 , n3716 );
nand ( n5582 , n51705 , n51706 );
buf ( n51708 , n5582 );
buf ( n51709 , n51708 );
nand ( n5585 , n5579 , n51709 );
buf ( n51711 , n5585 );
buf ( n51712 , n51711 );
xor ( n5588 , n51687 , n51712 );
buf ( n51714 , n385 );
not ( n5590 , n51714 );
and ( n5591 , n384 , n50571 );
not ( n5592 , n384 );
and ( n5593 , n5592 , n4369 );
or ( n5594 , n5591 , n5593 );
buf ( n51720 , n5594 );
not ( n5596 , n51720 );
or ( n5597 , n5590 , n5596 );
xor ( n5598 , n384 , n49998 );
buf ( n51724 , n5598 );
buf ( n51725 , n51066 );
nand ( n5601 , n51724 , n51725 );
buf ( n51727 , n5601 );
buf ( n51728 , n51727 );
nand ( n5604 , n5597 , n51728 );
buf ( n51730 , n5604 );
buf ( n51731 , n51730 );
xnor ( n5607 , n5588 , n51731 );
buf ( n51733 , n5607 );
buf ( n51734 , n51733 );
not ( n5610 , n51734 );
buf ( n51736 , n385 );
not ( n5612 , n51736 );
buf ( n51738 , n5598 );
not ( n5614 , n51738 );
or ( n5615 , n5612 , n5614 );
and ( n5616 , n5299 , n384 );
not ( n5617 , n5299 );
not ( n5618 , n384 );
and ( n5619 , n5617 , n5618 );
nor ( n5620 , n5616 , n5619 );
nand ( n5621 , n51066 , n5620 );
buf ( n51747 , n5621 );
nand ( n5623 , n5615 , n51747 );
buf ( n51749 , n5623 );
buf ( n51750 , n51749 );
not ( n5626 , n42494 );
nand ( n5627 , n5626 , n42141 );
not ( n5628 , n5627 );
not ( n5629 , n42664 );
nand ( n5630 , n42611 , n42633 , n5629 );
not ( n5631 , n5630 );
or ( n5632 , n5628 , n5631 );
nor ( n5633 , n42664 , n5627 );
nand ( n5634 , n42611 , n42633 , n5633 );
nand ( n5635 , n5632 , n5634 );
buf ( n51761 , n47838 );
buf ( n5637 , n51761 );
buf ( n51763 , n5637 );
not ( n5639 , n51763 );
buf ( n51765 , n51272 );
buf ( n51766 , n47318 );
nand ( n5642 , n51765 , n51766 );
buf ( n51768 , n5642 );
not ( n5644 , n51768 );
not ( n5645 , n5644 );
or ( n5646 , n5639 , n5645 );
not ( n5647 , n51768 );
or ( n5648 , n51763 , n5647 );
nand ( n5649 , n5646 , n5648 );
not ( n5650 , n394 );
nor ( n5651 , n5649 , n5650 );
buf ( n51777 , n5651 );
not ( n5653 , n51265 );
not ( n5654 , n51282 );
or ( n5655 , n5653 , n5654 );
or ( n5656 , n51265 , n51282 );
nand ( n5657 , n5655 , n5656 );
buf ( n51783 , n5657 );
xor ( n5659 , n51777 , n51783 );
buf ( n51785 , n3651 );
not ( n5661 , n51785 );
buf ( n51787 , n51541 );
not ( n5663 , n51787 );
or ( n5664 , n5661 , n5663 );
xor ( n5665 , n51499 , n51506 );
buf ( n51791 , n5665 );
buf ( n51792 , n51791 );
buf ( n51793 , n49447 );
nand ( n5669 , n51792 , n51793 );
buf ( n51795 , n5669 );
buf ( n51796 , n51795 );
nand ( n5672 , n5664 , n51796 );
buf ( n51798 , n5672 );
buf ( n51799 , n51798 );
and ( n5675 , n5659 , n51799 );
and ( n5676 , n51777 , n51783 );
or ( n5677 , n5675 , n5676 );
buf ( n51803 , n5677 );
not ( n5679 , n51803 );
xor ( n5680 , n5635 , n5679 );
not ( n5681 , n3622 );
not ( n5682 , n5350 );
or ( n5683 , n5681 , n5682 );
not ( n5684 , n50924 );
not ( n5685 , n50928 );
or ( n5686 , n5684 , n5685 );
nand ( n5687 , n5686 , n50934 );
and ( n5688 , n5687 , n380 );
not ( n5689 , n5687 );
not ( n5690 , n380 );
and ( n5691 , n5689 , n5690 );
nor ( n5692 , n5688 , n5691 );
nand ( n5693 , n3620 , n5692 );
nand ( n5694 , n5683 , n5693 );
xnor ( n5695 , n5680 , n5694 );
buf ( n51821 , n5695 );
xor ( n51822 , n51750 , n51821 );
xor ( n51823 , n51777 , n51783 );
xor ( n51824 , n51823 , n51799 );
buf ( n51825 , n51824 );
buf ( n51826 , n51825 );
buf ( n51827 , n3651 );
not ( n51828 , n51827 );
buf ( n51829 , n51791 );
not ( n51830 , n51829 );
or ( n5703 , n51828 , n51830 );
buf ( n51832 , n378 );
not ( n5705 , n51832 );
buf ( n51834 , n51264 );
not ( n5707 , n51834 );
buf ( n51836 , n5707 );
buf ( n51837 , n51836 );
not ( n51838 , n51837 );
or ( n5711 , n5705 , n51838 );
buf ( n51840 , n51261 );
buf ( n5713 , n51840 );
buf ( n51842 , n5713 );
buf ( n51843 , n51842 );
buf ( n51844 , n3654 );
nand ( n5717 , n51843 , n51844 );
buf ( n51846 , n5717 );
buf ( n51847 , n51846 );
nand ( n51848 , n5711 , n51847 );
buf ( n51849 , n51848 );
buf ( n51850 , n51849 );
buf ( n51851 , n49447 );
nand ( n51852 , n51850 , n51851 );
buf ( n51853 , n51852 );
buf ( n51854 , n51853 );
nand ( n51855 , n5703 , n51854 );
buf ( n51856 , n51855 );
buf ( n51857 , n51856 );
buf ( n51858 , n47507 );
not ( n51859 , n51858 );
buf ( n51860 , n47467 );
nand ( n51861 , n51859 , n51860 );
buf ( n51862 , n51861 );
and ( n51863 , n51862 , n1695 );
buf ( n51864 , n1972 );
xor ( n51865 , n51863 , n51864 );
and ( n51866 , n396 , n51865 );
buf ( n51867 , n395 );
and ( n51868 , n2022 , n47829 );
buf ( n51869 , n1983 );
xor ( n51870 , n51868 , n51869 );
buf ( n51871 , n51870 );
xor ( n51872 , n51867 , n51871 );
buf ( n51873 , n51261 );
not ( n51874 , n51873 );
buf ( n51875 , n3652 );
nor ( n51876 , n51874 , n51875 );
buf ( n51877 , n51876 );
buf ( n51878 , n51877 );
xor ( n51879 , n51872 , n51878 );
buf ( n51880 , n51879 );
xor ( n51881 , n51866 , n51880 );
xor ( n51882 , n396 , n51865 );
not ( n51883 , n51882 );
buf ( n51884 , n398 );
not ( n51885 , n47769 );
not ( n51886 , n47763 );
or ( n51887 , n51885 , n51886 );
nand ( n51888 , n51887 , n1889 );
nand ( n51889 , n47759 , n399 );
and ( n51890 , n51888 , n51889 );
not ( n51891 , n51888 );
not ( n51892 , n47759 );
nand ( n51893 , n51892 , n399 );
and ( n51894 , n51891 , n51893 );
nor ( n51895 , n51890 , n51894 );
buf ( n51896 , n51895 );
xor ( n51897 , n51884 , n51896 );
buf ( n51898 , n47675 );
not ( n51899 , n51898 );
buf ( n51900 , n47777 );
nand ( n51901 , n51899 , n51900 );
buf ( n51902 , n51901 );
xor ( n51903 , n1958 , n51902 );
buf ( n51904 , n51903 );
and ( n51905 , n51897 , n51904 );
and ( n51906 , n51884 , n51896 );
or ( n51907 , n51905 , n51906 );
buf ( n51908 , n51907 );
and ( n51909 , n397 , n51908 );
not ( n51910 , n51909 );
nand ( n51911 , n51883 , n51910 );
not ( n51912 , n51911 );
buf ( n51913 , n49395 );
buf ( n51914 , n49388 );
nand ( n51915 , n51913 , n51914 );
buf ( n51916 , n51915 );
not ( n51917 , n51916 );
not ( n51918 , n51264 );
or ( n51919 , n51917 , n51918 );
buf ( n51920 , n381 );
buf ( n51921 , n382 );
and ( n51922 , n51920 , n51921 );
buf ( n51923 , n3609 );
nor ( n51924 , n51922 , n51923 );
buf ( n51925 , n51924 );
nand ( n5726 , n51919 , n51925 );
not ( n5727 , n5726 );
not ( n5728 , n5727 );
or ( n5729 , n51912 , n5728 );
nand ( n5730 , n51882 , n51909 );
nand ( n5731 , n5729 , n5730 );
and ( n5732 , n51881 , n5731 );
and ( n5733 , n51866 , n51880 );
or ( n5734 , n5732 , n5733 );
buf ( n51935 , n5734 );
xor ( n5736 , n51857 , n51935 );
buf ( n51937 , n3609 );
buf ( n51938 , n49437 );
nand ( n5739 , n51937 , n51938 );
buf ( n51940 , n5739 );
buf ( n51941 , n51940 );
not ( n5742 , n51941 );
buf ( n51943 , n51264 );
not ( n5744 , n51943 );
or ( n5745 , n5742 , n5744 );
buf ( n51946 , n379 );
buf ( n51947 , n380 );
and ( n5748 , n51946 , n51947 );
buf ( n51949 , n3654 );
nor ( n5750 , n5748 , n51949 );
buf ( n51951 , n5750 );
buf ( n51952 , n51951 );
nand ( n5753 , n5745 , n51952 );
buf ( n51954 , n5753 );
not ( n5755 , n5650 );
not ( n5756 , n51763 );
not ( n5757 , n5644 );
or ( n5758 , n5756 , n5757 );
or ( n5759 , n51763 , n5647 );
nand ( n5760 , n5758 , n5759 );
not ( n5761 , n5760 );
or ( n5762 , n5755 , n5761 );
or ( n5763 , n5649 , n5650 );
nand ( n5764 , n5762 , n5763 );
not ( n5765 , n5764 );
xor ( n5766 , n51954 , n5765 );
xor ( n5767 , n51867 , n51871 );
and ( n5768 , n5767 , n51878 );
and ( n5769 , n51867 , n51871 );
or ( n5770 , n5768 , n5769 );
buf ( n51971 , n5770 );
xnor ( n5772 , n5766 , n51971 );
buf ( n51973 , n5772 );
and ( n5774 , n5736 , n51973 );
and ( n5775 , n51857 , n51935 );
or ( n5776 , n5774 , n5775 );
buf ( n51977 , n5776 );
buf ( n51978 , n51977 );
xor ( n5779 , n51826 , n51978 );
not ( n5780 , n3716 );
buf ( n51981 , n382 );
not ( n5782 , n51981 );
buf ( n51983 , n50537 );
not ( n5784 , n51983 );
or ( n5785 , n5782 , n5784 );
buf ( n51986 , n50540 );
buf ( n51987 , n49395 );
nand ( n5788 , n51986 , n51987 );
buf ( n51989 , n5788 );
buf ( n51990 , n51989 );
nand ( n5791 , n5785 , n51990 );
buf ( n51992 , n5791 );
not ( n5793 , n51992 );
or ( n5794 , n5780 , n5793 );
not ( n5795 , n382 );
not ( n5796 , n50794 );
or ( n5797 , n5795 , n5796 );
buf ( n51998 , n4956 );
buf ( n51999 , n49395 );
nand ( n5800 , n51998 , n51999 );
buf ( n52001 , n5800 );
nand ( n5802 , n5797 , n52001 );
nand ( n5803 , n5802 , n3733 );
nand ( n5804 , n5794 , n5803 );
buf ( n52005 , n5804 );
and ( n5806 , n5779 , n52005 );
and ( n5807 , n51826 , n51978 );
or ( n5808 , n5806 , n5807 );
buf ( n52009 , n5808 );
buf ( n52010 , n52009 );
and ( n5811 , n51822 , n52010 );
and ( n5812 , n51750 , n51821 );
or ( n5813 , n5811 , n5812 );
buf ( n52014 , n5813 );
buf ( n52015 , n52014 );
not ( n5816 , n52015 );
or ( n5817 , n5610 , n5816 );
buf ( n52018 , n52014 );
buf ( n52019 , n51733 );
or ( n5820 , n52018 , n52019 );
nand ( n5821 , n5817 , n5820 );
buf ( n52022 , n5821 );
buf ( n52023 , n52022 );
not ( n5824 , n5635 );
not ( n5825 , n5824 );
not ( n5826 , n5679 );
or ( n5827 , n5825 , n5826 );
nand ( n5828 , n5827 , n5694 );
nand ( n5829 , n51803 , n5635 );
nand ( n5830 , n5828 , n5829 );
buf ( n52031 , n5830 );
xor ( n5832 , n5342 , n51553 );
xnor ( n5833 , n5832 , n51485 );
buf ( n52034 , n5833 );
xor ( n5835 , n52031 , n52034 );
xor ( n5836 , n51509 , n51520 );
xor ( n5837 , n5836 , n51549 );
buf ( n52038 , n5837 );
buf ( n52039 , n52038 );
buf ( n52040 , n3716 );
not ( n5841 , n52040 );
buf ( n52042 , n51701 );
not ( n5843 , n52042 );
or ( n5844 , n5841 , n5843 );
buf ( n52045 , n51992 );
buf ( n52046 , n3733 );
nand ( n5847 , n52045 , n52046 );
buf ( n52048 , n5847 );
buf ( n52049 , n52048 );
nand ( n5850 , n5844 , n52049 );
buf ( n52051 , n5850 );
buf ( n52052 , n52051 );
xor ( n5853 , n52039 , n52052 );
not ( n5854 , n3622 );
not ( n5855 , n5692 );
or ( n5856 , n5854 , n5855 );
buf ( n52057 , n380 );
not ( n5858 , n52057 );
not ( n5859 , n50999 );
buf ( n52060 , n5859 );
not ( n5861 , n52060 );
or ( n5862 , n5858 , n5861 );
buf ( n52063 , n50999 );
buf ( n52064 , n3609 );
nand ( n5865 , n52063 , n52064 );
buf ( n52066 , n5865 );
buf ( n52067 , n52066 );
nand ( n5868 , n5862 , n52067 );
buf ( n52069 , n5868 );
buf ( n52070 , n52069 );
buf ( n52071 , n3620 );
nand ( n5872 , n52070 , n52071 );
buf ( n52073 , n5872 );
nand ( n5874 , n5856 , n52073 );
not ( n5875 , n5874 );
not ( n5876 , n42136 );
nor ( n5877 , n5876 , n42134 );
not ( n5878 , n5877 );
not ( n5879 , n42562 );
nor ( n5880 , n5879 , n42574 );
not ( n5881 , n5880 );
nand ( n5882 , n42541 , n42605 );
not ( n5883 , n5882 );
or ( n5884 , n5881 , n5883 );
not ( n5885 , n42547 );
nor ( n5886 , n42574 , n5885 );
nand ( n5887 , n42626 , n42128 );
nor ( n5888 , n5886 , n5887 );
nand ( n5889 , n5884 , n5888 );
not ( n5893 , n42128 );
nand ( n5894 , n42122 , n42100 );
not ( n5895 , n5894 );
or ( n5896 , n5893 , n5895 );
nand ( n5897 , n5896 , n42133 );
nor ( n5898 , C0 , n5897 );
nand ( n5899 , n5889 , n5898 );
not ( n5900 , n5899 );
or ( n5901 , n5878 , n5900 );
not ( n5902 , n5877 );
nand ( n5903 , n5898 , n5889 , n5902 );
nand ( n5904 , n5901 , n5903 );
nand ( n5905 , n5875 , n5904 );
not ( n5906 , n5905 );
not ( n5907 , n5765 );
not ( n5908 , n51954 );
not ( n5909 , n5908 );
or ( n5910 , n5907 , n5909 );
not ( n5911 , n51954 );
not ( n5912 , n5764 );
or ( n5913 , n5911 , n5912 );
nand ( n5914 , n5913 , n51971 );
nand ( n5915 , n5910 , n5914 );
not ( n5916 , n5915 );
or ( n5917 , n5906 , n5916 );
not ( n5918 , n5904 );
nand ( n5919 , n5918 , n5874 );
nand ( n5920 , n5917 , n5919 );
buf ( n52118 , n5920 );
and ( n5922 , n5853 , n52118 );
and ( n5923 , n52039 , n52052 );
or ( n5924 , n5922 , n5923 );
buf ( n52122 , n5924 );
buf ( n52123 , n52122 );
xor ( n5927 , n5835 , n52123 );
buf ( n52125 , n5927 );
buf ( n52126 , n52125 );
and ( n5930 , n52023 , n52126 );
not ( n5931 , n52023 );
buf ( n52129 , n52125 );
not ( n5933 , n52129 );
buf ( n52131 , n5933 );
buf ( n52132 , n52131 );
and ( n5936 , n5931 , n52132 );
nor ( n5937 , n5930 , n5936 );
buf ( n52135 , n5937 );
buf ( n52136 , n52135 );
xor ( n5940 , n52039 , n52052 );
xor ( n5941 , n5940 , n52118 );
buf ( n52139 , n5941 );
buf ( n52140 , n52139 );
not ( n5944 , n52140 );
buf ( n52142 , n5944 );
buf ( n52143 , n52142 );
not ( n5947 , n52143 );
not ( n5948 , n385 );
not ( n5949 , n5620 );
or ( n5950 , n5948 , n5949 );
not ( n5951 , n384 );
not ( n5952 , n50634 );
or ( n5953 , n5951 , n5952 );
buf ( n52151 , n384 );
not ( n5955 , n52151 );
buf ( n52153 , n5955 );
nand ( n5957 , n5070 , n52153 );
nand ( n5958 , n5953 , n5957 );
nand ( n5959 , n5958 , n51066 );
nand ( n5960 , n5950 , n5959 );
not ( n5961 , n5960 );
buf ( n52159 , n3622 );
not ( n5963 , n52159 );
buf ( n52161 , n52069 );
not ( n5965 , n52161 );
or ( n5966 , n5963 , n5965 );
buf ( n52164 , n380 );
buf ( n52165 , n51175 );
and ( n5969 , n52164 , n52165 );
not ( n5970 , n52164 );
buf ( n52168 , n51531 );
and ( n5972 , n5970 , n52168 );
nor ( n5973 , n5969 , n5972 );
buf ( n52171 , n5973 );
buf ( n52172 , n52171 );
buf ( n52173 , n3620 );
nand ( n5977 , n52172 , n52173 );
buf ( n52175 , n5977 );
buf ( n52176 , n52175 );
nand ( n5980 , n5966 , n52176 );
buf ( n52178 , n5980 );
buf ( n52179 , n52178 );
nand ( n5983 , n42582 , n42626 , n42593 );
not ( n5984 , n5894 );
nand ( n5985 , n42629 , n5983 , n5984 );
nand ( n5986 , n42128 , n42133 );
xnor ( n5987 , n5985 , n5986 );
buf ( n52185 , n5987 );
xor ( n5989 , n52179 , n52185 );
buf ( n52187 , n3716 );
not ( n5991 , n52187 );
buf ( n52189 , n5802 );
not ( n5993 , n52189 );
or ( n5994 , n5991 , n5993 );
not ( n5995 , n382 );
not ( n5996 , n5687 );
not ( n5997 , n5996 );
or ( n5998 , n5995 , n5997 );
buf ( n52196 , n49395 );
buf ( n52197 , n5687 );
nand ( n6001 , n52196 , n52197 );
buf ( n52199 , n6001 );
nand ( n6003 , n5998 , n52199 );
buf ( n52201 , n6003 );
buf ( n52202 , n3733 );
nand ( n6006 , n52201 , n52202 );
buf ( n52204 , n6006 );
buf ( n52205 , n52204 );
nand ( n6009 , n5994 , n52205 );
buf ( n52207 , n6009 );
buf ( n52208 , n52207 );
and ( n6012 , n5989 , n52208 );
and ( n6013 , n52179 , n52185 );
or ( n6014 , n6012 , n6013 );
buf ( n52212 , n6014 );
not ( n6016 , n52212 );
or ( n6017 , n5961 , n6016 );
buf ( n52215 , n52212 );
buf ( n52216 , n5960 );
or ( n6020 , n52215 , n52216 );
xor ( n6021 , n5915 , n5904 );
xnor ( n6022 , n6021 , n5874 );
buf ( n52220 , n6022 );
nand ( n6024 , n6020 , n52220 );
buf ( n52222 , n6024 );
nand ( n6026 , n6017 , n52222 );
not ( n6027 , n6026 );
buf ( n52225 , n6027 );
not ( n6029 , n52225 );
or ( n6030 , n5947 , n6029 );
xor ( n6031 , n51750 , n51821 );
xor ( n6032 , n6031 , n52010 );
buf ( n52230 , n6032 );
buf ( n52231 , n52230 );
nand ( n6035 , n6030 , n52231 );
buf ( n52233 , n6035 );
buf ( n52234 , n52233 );
buf ( n52235 , n52142 );
buf ( n52236 , n6027 );
or ( n6040 , n52235 , n52236 );
buf ( n52238 , n6040 );
buf ( n52239 , n52238 );
and ( n6043 , n52234 , n52239 );
buf ( n52241 , n6043 );
buf ( n52242 , n52241 );
nand ( n6046 , n52136 , n52242 );
buf ( n52244 , n6046 );
not ( n6048 , n52244 );
buf ( n52246 , n51264 );
buf ( n52247 , n3622 );
and ( n6051 , n52246 , n52247 );
buf ( n52249 , n6051 );
buf ( n52250 , n1971 );
buf ( n52251 , n47580 );
not ( n6055 , n52251 );
buf ( n52253 , n47597 );
nand ( n6057 , n6055 , n52253 );
buf ( n52255 , n6057 );
buf ( n52256 , n52255 );
nand ( n6060 , n52250 , n52256 );
buf ( n52258 , n6060 );
buf ( n52259 , n52258 );
buf ( n52260 , n47780 );
xnor ( n6064 , n52259 , n52260 );
buf ( n52262 , n6064 );
xor ( n6066 , n397 , n51908 );
and ( n6067 , n52262 , n6066 );
not ( n6068 , n52262 );
not ( n6069 , n6066 );
and ( n6070 , n6068 , n6069 );
nor ( n6071 , n6067 , n6070 );
xor ( n6072 , n52249 , n6071 );
not ( n6073 , n3716 );
not ( n6074 , n382 );
not ( n6075 , n51531 );
or ( n6076 , n6074 , n6075 );
buf ( n52274 , n51175 );
buf ( n52275 , n49395 );
nand ( n6079 , n52274 , n52275 );
buf ( n52277 , n6079 );
nand ( n6081 , n6076 , n52277 );
not ( n6082 , n6081 );
or ( n6083 , n6073 , n6082 );
buf ( n52281 , n382 );
not ( n6085 , n52281 );
buf ( n52283 , n5380 );
not ( n6087 , n52283 );
buf ( n52285 , n6087 );
buf ( n52286 , n52285 );
not ( n6090 , n52286 );
or ( n6091 , n6085 , n6090 );
buf ( n52289 , n49395 );
buf ( n52290 , n5380 );
nand ( n6094 , n52289 , n52290 );
buf ( n52292 , n6094 );
buf ( n52293 , n52292 );
nand ( n6097 , n6091 , n52293 );
buf ( n52295 , n6097 );
buf ( n52296 , n52295 );
buf ( n52297 , n3733 );
nand ( n6101 , n52296 , n52297 );
buf ( n52299 , n6101 );
nand ( n6103 , n6083 , n52299 );
xor ( n6104 , n6072 , n6103 );
nand ( n6109 , C1 , n42659 );
nand ( n6110 , n42546 , n42573 );
not ( n6111 , n6110 );
and ( n6112 , n6109 , n6111 );
not ( n6113 , n6109 );
and ( n6114 , n6113 , n6110 );
nor ( n6115 , n6112 , n6114 );
and ( n6116 , n6104 , n6115 );
and ( n6117 , n6072 , n6103 );
or ( n6118 , n6116 , n6117 );
not ( n6119 , n6118 );
nand ( n6120 , n42418 , n42113 );
nand ( n6124 , C1 , n42644 );
or ( n6125 , n6120 , n6124 );
nand ( n6126 , n6124 , n6120 );
nand ( n6127 , n6125 , n6126 );
not ( n6128 , n6127 );
buf ( n52319 , n382 );
not ( n6130 , n52319 );
buf ( n52321 , n5859 );
not ( n6132 , n52321 );
or ( n6133 , n6130 , n6132 );
buf ( n52324 , n49395 );
buf ( n52325 , n50999 );
nand ( n6136 , n52324 , n52325 );
buf ( n52327 , n6136 );
buf ( n52328 , n52327 );
nand ( n6139 , n6133 , n52328 );
buf ( n52330 , n6139 );
and ( n6141 , n52330 , n3716 );
and ( n6142 , n6081 , n3733 );
nor ( n6143 , n6141 , n6142 );
nand ( n6144 , n6128 , n6143 );
not ( n6145 , n6144 );
or ( n6146 , n6119 , n6145 );
not ( n6147 , n6143 );
nand ( n6148 , n6147 , n6127 );
nand ( n6149 , n6146 , n6148 );
not ( n6150 , n6149 );
buf ( n52341 , n6150 );
not ( n6152 , n52341 );
not ( n6153 , n3716 );
not ( n6154 , n6003 );
or ( n6155 , n6153 , n6154 );
nand ( n6156 , n52330 , n3733 );
nand ( n6157 , n6155 , n6156 );
buf ( n52348 , n6157 );
not ( n6159 , n52262 );
nand ( n6160 , n6159 , n6069 );
not ( n6161 , n6160 );
not ( n6162 , n52249 );
or ( n6163 , n6161 , n6162 );
nand ( n6164 , n6066 , n52262 );
nand ( n6165 , n6163 , n6164 );
buf ( n52356 , n6165 );
not ( n6167 , n52356 );
buf ( n52358 , n3622 );
not ( n6169 , n52358 );
buf ( n52360 , n380 );
not ( n6171 , n52360 );
buf ( n52362 , n52285 );
not ( n6173 , n52362 );
or ( n6174 , n6171 , n6173 );
buf ( n52365 , n3609 );
buf ( n52366 , n5380 );
nand ( n6177 , n52365 , n52366 );
buf ( n52368 , n6177 );
buf ( n52369 , n52368 );
nand ( n6180 , n6174 , n52369 );
buf ( n52371 , n6180 );
buf ( n52372 , n52371 );
not ( n6183 , n52372 );
or ( n6184 , n6169 , n6183 );
buf ( n52375 , n51842 );
buf ( n52376 , n3609 );
nand ( n6187 , n52375 , n52376 );
buf ( n52378 , n6187 );
buf ( n52379 , n52378 );
not ( n6190 , n52379 );
not ( n6191 , n51842 );
buf ( n52382 , n6191 );
buf ( n52383 , n380 );
nand ( n6194 , n52382 , n52383 );
buf ( n52385 , n6194 );
buf ( n52386 , n52385 );
not ( n6197 , n52386 );
or ( n6198 , n6190 , n6197 );
buf ( n52389 , n3620 );
nand ( n6200 , n6198 , n52389 );
buf ( n52391 , n6200 );
buf ( n52392 , n52391 );
nand ( n6203 , n6184 , n52392 );
buf ( n52394 , n6203 );
buf ( n52395 , n52394 );
not ( n6206 , n52395 );
or ( n6207 , n6167 , n6206 );
or ( n6208 , n52394 , n6165 );
xor ( n6209 , n51882 , n51910 );
xnor ( n6210 , n6209 , n5726 );
not ( n6211 , n6210 );
nand ( n6212 , n6208 , n6211 );
buf ( n52403 , n6212 );
nand ( n6214 , n6207 , n52403 );
buf ( n52405 , n6214 );
buf ( n52406 , n52405 );
xnor ( n6217 , n52348 , n52406 );
buf ( n52408 , n6217 );
buf ( n52409 , n52408 );
not ( n6220 , n52409 );
not ( n6221 , n385 );
and ( n6222 , n384 , n50537 );
not ( n6223 , n384 );
and ( n6224 , n6223 , n50540 );
or ( n6225 , n6222 , n6224 );
not ( n6226 , n6225 );
or ( n6227 , n6221 , n6226 );
not ( n6228 , n384 );
not ( n6229 , n50794 );
or ( n6230 , n6228 , n6229 );
not ( n6231 , n384 );
nand ( n6232 , n6231 , n4956 );
nand ( n6233 , n6230 , n6232 );
nand ( n6234 , n6233 , n51066 );
nand ( n6235 , n6227 , n6234 );
buf ( n52426 , n6235 );
not ( n6237 , n52426 );
and ( n6238 , n6220 , n6237 );
buf ( n52429 , n6235 );
buf ( n52430 , n52408 );
and ( n6241 , n52429 , n52430 );
nor ( n6242 , n6238 , n6241 );
buf ( n52433 , n6242 );
buf ( n52434 , n52433 );
not ( n6245 , n52434 );
or ( n6246 , n6152 , n6245 );
buf ( n52437 , n3622 );
not ( n6248 , n52437 );
buf ( n52439 , n52171 );
not ( n6250 , n52439 );
or ( n6251 , n6248 , n6250 );
buf ( n52442 , n52371 );
buf ( n52443 , n3620 );
nand ( n6254 , n52442 , n52443 );
buf ( n52445 , n6254 );
buf ( n52446 , n52445 );
nand ( n6257 , n6251 , n52446 );
buf ( n52448 , n6257 );
xor ( n6259 , n51866 , n51880 );
xor ( n6260 , n6259 , n5731 );
xor ( n6261 , n52448 , n6260 );
xnor ( n6262 , n6261 , n42703 );
not ( n6263 , n6262 );
buf ( n52454 , n6263 );
nand ( n6265 , n6246 , n52454 );
buf ( n52456 , n6265 );
buf ( n52457 , n52456 );
buf ( n52458 , n52433 );
not ( n6269 , n52458 );
buf ( n52460 , n6149 );
nand ( n6271 , n6269 , n52460 );
buf ( n52462 , n6271 );
buf ( n52463 , n52462 );
nand ( n6274 , n52457 , n52463 );
buf ( n52465 , n6274 );
buf ( n52466 , n52465 );
xor ( n6277 , n52179 , n52185 );
xor ( n6278 , n6277 , n52208 );
buf ( n52469 , n6278 );
buf ( n52470 , n52469 );
buf ( n52471 , n6157 );
buf ( n6282 , n52471 );
buf ( n52473 , n6282 );
buf ( n52474 , n52473 );
not ( n6285 , n52474 );
buf ( n52476 , n6235 );
not ( n6287 , n52476 );
or ( n6288 , n6285 , n6287 );
buf ( n52479 , n6235 );
buf ( n52480 , n52473 );
or ( n6291 , n52479 , n52480 );
buf ( n52482 , n52405 );
nand ( n6293 , n6291 , n52482 );
buf ( n52484 , n6293 );
buf ( n52485 , n52484 );
nand ( n6296 , n6288 , n52485 );
buf ( n52487 , n6296 );
buf ( n52488 , n52487 );
xor ( n6299 , n52470 , n52488 );
xor ( n6300 , n51857 , n51935 );
xor ( n6301 , n6300 , n51973 );
buf ( n52492 , n6301 );
buf ( n52493 , n52492 );
not ( n6304 , n52448 );
not ( n6305 , n6260 );
or ( n6306 , n6304 , n6305 );
or ( n6307 , n52448 , n6260 );
nand ( n6308 , n6307 , n42703 );
nand ( n6309 , n6306 , n6308 );
buf ( n52500 , n6309 );
xor ( n6311 , n52493 , n52500 );
buf ( n52502 , n385 );
not ( n6313 , n52502 );
buf ( n52504 , n5958 );
not ( n6315 , n52504 );
or ( n6316 , n6313 , n6315 );
buf ( n52507 , n6225 );
buf ( n52508 , n51066 );
nand ( n6319 , n52507 , n52508 );
buf ( n52510 , n6319 );
buf ( n52511 , n52510 );
nand ( n6322 , n6316 , n52511 );
buf ( n52513 , n6322 );
buf ( n52514 , n52513 );
xor ( n6325 , n6311 , n52514 );
buf ( n52516 , n6325 );
buf ( n52517 , n52516 );
xor ( n6328 , n6299 , n52517 );
buf ( n52519 , n6328 );
buf ( n52520 , n52519 );
xor ( n6331 , n52466 , n52520 );
not ( n6332 , n6211 );
buf ( n52523 , n6165 );
not ( n6334 , n52523 );
buf ( n52525 , n6334 );
not ( n6336 , n52525 );
or ( n6337 , n6332 , n6336 );
nand ( n6338 , n6210 , n6165 );
nand ( n6339 , n6337 , n6338 );
not ( n6340 , n52394 );
and ( n6341 , n6339 , n6340 );
not ( n6342 , n6339 );
and ( n6343 , n6342 , n52394 );
nor ( n6344 , n6341 , n6343 );
not ( n6345 , n6344 );
buf ( n52536 , n6345 );
not ( n6347 , n52536 );
not ( n6348 , n385 );
not ( n6349 , n6233 );
or ( n6350 , n6348 , n6349 );
and ( n6351 , n384 , n5996 );
not ( n6352 , n384 );
and ( n6353 , n6352 , n5687 );
or ( n6354 , n6351 , n6353 );
nand ( n6355 , n6354 , n51066 );
nand ( n6356 , n6350 , n6355 );
buf ( n52547 , n6356 );
not ( n6358 , n52547 );
or ( n6359 , n6347 , n6358 );
buf ( n52550 , n6356 );
not ( n6361 , n52550 );
buf ( n52552 , n6344 );
nand ( n6363 , n6361 , n52552 );
buf ( n52554 , n6363 );
not ( n6365 , n385 );
not ( n6366 , n6354 );
or ( n6367 , n6365 , n6366 );
buf ( n52558 , n384 );
buf ( n52559 , n50999 );
and ( n6370 , n52558 , n52559 );
not ( n6371 , n52558 );
buf ( n52562 , n5859 );
and ( n6373 , n6371 , n52562 );
nor ( n6374 , n6370 , n6373 );
buf ( n52565 , n6374 );
buf ( n52566 , n52565 );
buf ( n52567 , n51066 );
nand ( n6378 , n52566 , n52567 );
buf ( n52569 , n6378 );
nand ( n6380 , n6367 , n52569 );
not ( n6381 , n6380 );
xor ( n6382 , n51884 , n51896 );
xor ( n6383 , n6382 , n51904 );
buf ( n52574 , n6383 );
buf ( n52575 , n52574 );
buf ( n52576 , n384 );
not ( n6387 , n52576 );
buf ( n52578 , n49502 );
nand ( n6389 , n6387 , n52578 );
buf ( n52580 , n6389 );
buf ( n52581 , n52580 );
not ( n6392 , n52581 );
buf ( n52583 , n51842 );
not ( n6394 , n52583 );
or ( n6395 , n6392 , n6394 );
buf ( n52586 , n383 );
buf ( n52587 , n384 );
and ( n6398 , n52586 , n52587 );
buf ( n52589 , n49395 );
nor ( n6400 , n6398 , n52589 );
buf ( n52591 , n6400 );
buf ( n52592 , n52591 );
nand ( n6403 , n6395 , n52592 );
buf ( n52594 , n6403 );
buf ( n52595 , n52594 );
not ( n6406 , n52595 );
buf ( n52597 , n6406 );
buf ( n52598 , n52597 );
xor ( n6409 , n52575 , n52598 );
buf ( n52600 , n3716 );
not ( n6411 , n52600 );
buf ( n52602 , n52295 );
not ( n6413 , n52602 );
or ( n6414 , n6411 , n6413 );
not ( n6415 , n51842 );
nand ( n6416 , n6415 , n382 );
not ( n6417 , n6416 );
buf ( n52608 , n51842 );
buf ( n52609 , n49395 );
nand ( n6420 , n52608 , n52609 );
buf ( n52611 , n6420 );
not ( n6422 , n52611 );
or ( n6423 , n6417 , n6422 );
nand ( n6424 , n6423 , n3733 );
buf ( n52615 , n6424 );
nand ( n6426 , n6414 , n52615 );
buf ( n52617 , n6426 );
buf ( n52618 , n52617 );
and ( n6429 , n6409 , n52618 );
and ( n6430 , n52575 , n52598 );
or ( n6431 , n6429 , n6430 );
buf ( n52622 , n6431 );
not ( n6433 , n52622 );
or ( n6434 , n6381 , n6433 );
buf ( n52625 , n52622 );
buf ( n52626 , n6380 );
or ( n6437 , n52625 , n52626 );
xor ( n6438 , n6072 , n6103 );
xor ( n6439 , n6438 , n6115 );
buf ( n52630 , n6439 );
nand ( n6441 , n6437 , n52630 );
buf ( n52632 , n6441 );
nand ( n6443 , n6434 , n52632 );
nand ( n6444 , n52554 , n6443 );
buf ( n52635 , n6444 );
nand ( n6446 , n6359 , n52635 );
buf ( n52637 , n6446 );
buf ( n52638 , n52637 );
not ( n6449 , n52638 );
xnor ( n6450 , n6262 , n6149 );
buf ( n52641 , n6450 );
not ( n6452 , n52641 );
buf ( n52643 , n52433 );
not ( n6454 , n52643 );
and ( n6455 , n6452 , n6454 );
buf ( n52646 , n6450 );
buf ( n52647 , n52433 );
and ( n6458 , n52646 , n52647 );
nor ( n6459 , n6455 , n6458 );
buf ( n52650 , n6459 );
buf ( n52651 , n52650 );
nand ( n6462 , n6449 , n52651 );
buf ( n52653 , n6462 );
buf ( n52654 , n52653 );
not ( n6465 , n52654 );
not ( n6466 , n6356 );
not ( n6467 , n6345 );
or ( n6468 , n6466 , n6467 );
not ( n6469 , n6356 );
nand ( n6470 , n6469 , n6344 );
nand ( n6471 , n6468 , n6470 );
not ( n6472 , n6471 );
not ( n6473 , n6443 );
or ( n6474 , n6472 , n6473 );
not ( n6475 , n6127 );
not ( n6476 , n6143 );
not ( n6477 , n6476 );
or ( n6478 , n6475 , n6477 );
or ( n6479 , n6127 , n6476 );
nand ( n6480 , n6478 , n6479 );
buf ( n52671 , n6480 );
buf ( n52672 , n6118 );
xor ( n6483 , n52671 , n52672 );
buf ( n52674 , n6483 );
nand ( n6485 , n6474 , n52674 );
not ( n6486 , n6485 );
not ( n6487 , n6443 );
not ( n6488 , n6471 );
nand ( n6489 , n6487 , n6488 );
nand ( n6490 , n6486 , n6489 );
not ( n6491 , n6490 );
buf ( n52682 , n51066 );
not ( n6493 , n52682 );
buf ( n52684 , n384 );
not ( n6495 , n52684 );
buf ( n52686 , n52285 );
not ( n6497 , n52686 );
or ( n6498 , n6495 , n6497 );
buf ( n52689 , n384 );
not ( n6500 , n52689 );
buf ( n52691 , n5380 );
nand ( n6502 , n6500 , n52691 );
buf ( n52693 , n6502 );
buf ( n52694 , n52693 );
nand ( n6505 , n6498 , n52694 );
buf ( n52696 , n6505 );
buf ( n52697 , n52696 );
not ( n6508 , n52697 );
or ( n6509 , n6493 , n6508 );
buf ( n52700 , n384 );
buf ( n52701 , n51531 );
and ( n6512 , n52700 , n52701 );
not ( n6513 , n52700 );
buf ( n52704 , n51175 );
and ( n6515 , n6513 , n52704 );
nor ( n6516 , n6512 , n6515 );
buf ( n52707 , n6516 );
buf ( n52708 , n52707 );
buf ( n52709 , n51065 );
or ( n6520 , n52708 , n52709 );
nand ( n6521 , n6509 , n6520 );
buf ( n52712 , n6521 );
buf ( n52713 , n52712 );
not ( n6524 , n47759 );
not ( n6525 , n51888 );
or ( n6526 , n6524 , n6525 );
or ( n6527 , n51888 , n47759 );
nand ( n6528 , n6526 , n6527 );
buf ( n52719 , n6528 );
buf ( n52720 , n399 );
xor ( n6531 , n52719 , n52720 );
buf ( n52722 , n6531 );
buf ( n52723 , n52722 );
buf ( n52724 , n51842 );
buf ( n52725 , n3716 );
and ( n6536 , n52724 , n52725 );
buf ( n52727 , n6536 );
buf ( n52728 , n52727 );
xor ( n6539 , n52723 , n52728 );
buf ( n52730 , n400 );
buf ( n52731 , n47738 );
not ( n6542 , n52731 );
buf ( n52733 , n47756 );
nand ( n6544 , n6542 , n52733 );
buf ( n52735 , n6544 );
buf ( n52736 , n52735 );
buf ( n52737 , n47750 );
xor ( n6548 , n52736 , n52737 );
buf ( n52739 , n6548 );
buf ( n52740 , n52739 );
xor ( n6551 , n52730 , n52740 );
buf ( n52742 , n51261 );
buf ( n52743 , n385 );
nand ( n6554 , n52742 , n52743 );
buf ( n52745 , n6554 );
buf ( n52746 , n52745 );
buf ( n52747 , n384 );
and ( n6558 , n52746 , n52747 );
buf ( n52749 , n6558 );
buf ( n52750 , n52749 );
and ( n6561 , n6551 , n52750 );
and ( n6562 , n52730 , n52740 );
or ( n6563 , n6561 , n6562 );
buf ( n52754 , n6563 );
buf ( n52755 , n52754 );
xor ( n6566 , n6539 , n52755 );
buf ( n52757 , n6566 );
buf ( n52758 , n52757 );
xor ( n6569 , n52713 , n52758 );
buf ( n52760 , n401 );
not ( n6571 , n52760 );
or ( n6572 , n47619 , n47744 );
nand ( n6573 , n6572 , n47747 );
buf ( n52764 , n6573 );
not ( n6575 , n52764 );
or ( n6576 , n6571 , n6575 );
buf ( n52767 , n52745 );
buf ( n52768 , n6573 );
buf ( n52769 , n401 );
nor ( n6580 , n52768 , n52769 );
buf ( n52771 , n6580 );
buf ( n52772 , n52771 );
or ( n6583 , n52767 , n52772 );
nand ( n6584 , n6576 , n6583 );
buf ( n52775 , n6584 );
buf ( n52776 , n52775 );
xor ( n6587 , n52730 , n52740 );
xor ( n6588 , n6587 , n52750 );
buf ( n52779 , n6588 );
buf ( n52780 , n52779 );
xor ( n6591 , n52776 , n52780 );
not ( n6592 , n385 );
not ( n6593 , n52696 );
or ( n6594 , n6592 , n6593 );
nand ( n6595 , n6191 , n51066 );
nand ( n6596 , n6594 , n6595 );
buf ( n52787 , n6596 );
and ( n6598 , n6591 , n52787 );
and ( n6599 , n52776 , n52780 );
or ( n6600 , n6598 , n6599 );
buf ( n52791 , n6600 );
buf ( n52792 , n52791 );
and ( n6603 , n6569 , n52792 );
and ( n6604 , n52713 , n52758 );
or ( n6605 , n6603 , n6604 );
buf ( n52796 , n6605 );
xor ( n6607 , n52575 , n52598 );
xor ( n6608 , n6607 , n52618 );
buf ( n52799 , n6608 );
nor ( n6610 , n52796 , n52799 );
not ( n6611 , n5879 );
and ( n6612 , n5882 , n6611 );
nand ( n6613 , n6612 , n42610 );
and ( n6614 , n6613 , n42695 );
not ( n6615 , n6613 );
and ( n6616 , n6615 , n42692 );
nor ( n6617 , n6614 , n6616 );
xor ( n6618 , n52723 , n52728 );
and ( n6619 , n6618 , n52755 );
and ( n6620 , n52723 , n52728 );
or ( n6621 , n6619 , n6620 );
buf ( n52812 , n6621 );
xor ( n6623 , n6617 , n52812 );
buf ( n52814 , n385 );
not ( n6625 , n52814 );
buf ( n52816 , n52565 );
not ( n6627 , n52816 );
or ( n6628 , n6625 , n6627 );
buf ( n52819 , n52707 );
not ( n6630 , n52819 );
buf ( n52821 , n51066 );
nand ( n6632 , n6630 , n52821 );
buf ( n52823 , n6632 );
buf ( n52824 , n52823 );
nand ( n6635 , n6628 , n52824 );
buf ( n52826 , n6635 );
xor ( n6637 , n6623 , n52826 );
not ( n6638 , n6637 );
or ( n6639 , n6610 , n6638 );
nand ( n6640 , n52796 , n52799 );
nand ( n6641 , n6639 , n6640 );
not ( n6642 , n6641 );
xor ( n6643 , n6617 , n52812 );
and ( n6644 , n6643 , n52826 );
and ( n6645 , n6617 , n52812 );
or ( n6646 , n6644 , n6645 );
not ( n6647 , n6646 );
buf ( n52838 , n52622 );
buf ( n52839 , n6380 );
xor ( n6650 , n52838 , n52839 );
buf ( n52841 , n6439 );
xnor ( n6652 , n6650 , n52841 );
buf ( n52843 , n6652 );
nand ( n6654 , n6647 , n52843 );
not ( n6655 , n6654 );
or ( n6656 , n6642 , n6655 );
not ( n6657 , n52843 );
nand ( n6658 , n6657 , n6646 );
nand ( n6659 , n6656 , n6658 );
not ( n6660 , n6659 );
or ( n6661 , n6491 , n6660 );
buf ( n52852 , n52674 );
not ( n6663 , n52852 );
buf ( n52854 , n6663 );
not ( n6665 , n6487 );
nand ( n6666 , n6665 , n6488 );
not ( n6667 , n6443 );
nand ( n6668 , n6667 , n6471 );
nand ( n6669 , n52854 , n6666 , n6668 );
nand ( n6670 , n6661 , n6669 );
buf ( n52861 , n6670 );
not ( n6672 , n52861 );
or ( n6673 , n6465 , n6672 );
buf ( n52864 , n52650 );
not ( n6675 , n52864 );
buf ( n52866 , n52637 );
nand ( n6677 , n6675 , n52866 );
buf ( n52868 , n6677 );
buf ( n52869 , n52868 );
nand ( n6680 , n6673 , n52869 );
buf ( n52871 , n6680 );
buf ( n52872 , n52871 );
and ( n6683 , n6331 , n52872 );
and ( n6684 , n52466 , n52520 );
or ( n6685 , n6683 , n6684 );
buf ( n52876 , n6685 );
buf ( n52877 , n52876 );
not ( n6688 , n52877 );
buf ( n52879 , n52139 );
buf ( n52880 , n6026 );
and ( n6691 , n52879 , n52880 );
not ( n6692 , n52879 );
buf ( n52883 , n6027 );
and ( n6694 , n6692 , n52883 );
nor ( n6695 , n6691 , n6694 );
buf ( n52886 , n6695 );
buf ( n52887 , n52230 );
not ( n6698 , n52887 );
buf ( n52889 , n6698 );
and ( n6700 , n52886 , n52889 );
not ( n6701 , n52886 );
and ( n6702 , n6701 , n52230 );
nor ( n6703 , n6700 , n6702 );
xor ( n6704 , n51826 , n51978 );
xor ( n6705 , n6704 , n52005 );
buf ( n52896 , n6705 );
xor ( n6707 , n52493 , n52500 );
and ( n6708 , n6707 , n52514 );
and ( n6709 , n52493 , n52500 );
or ( n6710 , n6708 , n6709 );
buf ( n52901 , n6710 );
xor ( n6712 , n52896 , n52901 );
buf ( n52903 , n6022 );
not ( n6714 , n52903 );
buf ( n52905 , n5960 );
not ( n6716 , n52905 );
buf ( n52907 , n6716 );
buf ( n52908 , n52907 );
not ( n6719 , n52908 );
or ( n6720 , n6714 , n6719 );
not ( n6721 , n6022 );
buf ( n52912 , n6721 );
buf ( n52913 , n5960 );
nand ( n6724 , n52912 , n52913 );
buf ( n52915 , n6724 );
buf ( n52916 , n52915 );
nand ( n6727 , n6720 , n52916 );
buf ( n52918 , n6727 );
buf ( n52919 , n52918 );
buf ( n52920 , n52212 );
and ( n6731 , n52919 , n52920 );
not ( n6732 , n52919 );
buf ( n52923 , n52212 );
not ( n6734 , n52923 );
buf ( n52925 , n6734 );
buf ( n52926 , n52925 );
and ( n6737 , n6732 , n52926 );
nor ( n6738 , n6731 , n6737 );
buf ( n52929 , n6738 );
and ( n6740 , n6712 , n52929 );
and ( n6741 , n52896 , n52901 );
or ( n6742 , n6740 , n6741 );
not ( n6743 , n6742 );
nand ( n6744 , n6703 , n6743 );
buf ( n52935 , n6744 );
xor ( n6746 , n52470 , n52488 );
and ( n6747 , n6746 , n52517 );
and ( n6748 , n52470 , n52488 );
or ( n6749 , n6747 , n6748 );
buf ( n52940 , n6749 );
not ( n6751 , n52940 );
xor ( n6752 , n52896 , n52901 );
xor ( n6753 , n6752 , n52929 );
not ( n6754 , n6753 );
nand ( n6755 , n6751 , n6754 );
buf ( n52946 , n6755 );
and ( n6757 , n52935 , n52946 );
buf ( n52948 , n6757 );
buf ( n52949 , n52948 );
not ( n6760 , n52949 );
or ( n6761 , n6688 , n6760 );
buf ( n52952 , n6753 );
buf ( n52953 , n52940 );
nand ( n6764 , n52952 , n52953 );
buf ( n52955 , n6764 );
buf ( n52956 , n52955 );
not ( n6767 , n52956 );
buf ( n52958 , n6744 );
nand ( n6769 , n6767 , n52958 );
buf ( n52960 , n6769 );
not ( n6771 , n6703 );
buf ( n6772 , n6742 );
nand ( n6773 , n6771 , n6772 );
nand ( n6774 , n52960 , n6773 );
buf ( n52965 , n6774 );
not ( n6776 , n52965 );
buf ( n52967 , n6776 );
buf ( n52968 , n52967 );
nand ( n6779 , n6761 , n52968 );
buf ( n52970 , n6779 );
not ( n6781 , n52970 );
or ( n6782 , n6048 , n6781 );
buf ( n52973 , n52135 );
buf ( n52974 , n52241 );
or ( n6785 , n52973 , n52974 );
buf ( n52976 , n6785 );
nand ( n6787 , n6782 , n52976 );
not ( n6788 , n6787 );
buf ( n52979 , n51389 );
buf ( n52980 , n5441 );
xor ( n6791 , n52979 , n52980 );
buf ( n52982 , n51572 );
xnor ( n6793 , n6791 , n52982 );
buf ( n52984 , n6793 );
xor ( n6795 , n51414 , n5434 );
xor ( n6796 , n6795 , n5438 );
buf ( n52987 , n6796 );
not ( n6798 , n52987 );
buf ( n52989 , n6798 );
not ( n6800 , n52989 );
buf ( n52991 , n5215 );
and ( n6802 , n51157 , n51213 );
not ( n6803 , n51157 );
and ( n6804 , n6803 , n51216 );
nor ( n6805 , n6802 , n6804 );
buf ( n52996 , n6805 );
xnor ( n6807 , n52991 , n52996 );
buf ( n52998 , n6807 );
not ( n6809 , n52998 );
and ( n6810 , n6800 , n6809 );
buf ( n53001 , n52989 );
buf ( n53002 , n52998 );
nand ( n6813 , n53001 , n53002 );
buf ( n53004 , n6813 );
and ( n6815 , n51228 , n5201 );
not ( n6816 , n51228 );
not ( n6817 , n5201 );
and ( n6818 , n6816 , n6817 );
nor ( n6819 , n6815 , n6818 );
and ( n6820 , n6819 , n5212 );
not ( n6821 , n6819 );
not ( n6822 , n5212 );
and ( n6823 , n6821 , n6822 );
nor ( n6824 , n6820 , n6823 );
buf ( n53015 , n6824 );
not ( n6826 , n53015 );
not ( n6827 , n51066 );
not ( n6828 , n5594 );
or ( n6829 , n6827 , n6828 );
nand ( n6830 , n5282 , n385 );
nand ( n6831 , n6829 , n6830 );
not ( n6832 , n6831 );
buf ( n53023 , n6832 );
not ( n6834 , n53023 );
or ( n6835 , n6826 , n6834 );
not ( n6836 , n51711 );
not ( n6837 , n51730 );
or ( n6838 , n6836 , n6837 );
buf ( n53029 , n51730 );
buf ( n53030 , n51711 );
or ( n6841 , n53029 , n53030 );
buf ( n53032 , n5561 );
nand ( n6843 , n6841 , n53032 );
buf ( n53034 , n6843 );
nand ( n6845 , n6838 , n53034 );
buf ( n53036 , n6845 );
nand ( n6847 , n6835 , n53036 );
buf ( n53038 , n6847 );
buf ( n53039 , n53038 );
buf ( n53040 , n6824 );
not ( n6851 , n53040 );
buf ( n53042 , n6831 );
nand ( n6853 , n6851 , n53042 );
buf ( n53044 , n6853 );
buf ( n53045 , n53044 );
nand ( n6856 , n53039 , n53045 );
buf ( n53047 , n6856 );
and ( n6858 , n53004 , n53047 );
nor ( n6859 , n6810 , n6858 );
nand ( n6860 , n52984 , n6859 );
buf ( n53051 , n6860 );
not ( n6862 , n5432 );
not ( n6863 , n5318 );
not ( n6864 , n51435 );
not ( n6865 , n6864 );
or ( n6866 , n6863 , n6865 );
nand ( n6867 , n51442 , n51435 );
nand ( n6868 , n6866 , n6867 );
xnor ( n6869 , n6862 , n6868 );
not ( n6870 , n6869 );
buf ( n53061 , n5830 );
not ( n6872 , n53061 );
buf ( n53063 , n6872 );
not ( n6874 , n53063 );
not ( n6875 , n5833 );
or ( n6876 , n6874 , n6875 );
nand ( n6877 , n6876 , n52122 );
not ( n6878 , n5833 );
nand ( n6879 , n6878 , n5830 );
nand ( n6880 , n6877 , n6879 );
not ( n6881 , n6880 );
or ( n6882 , n6870 , n6881 );
not ( n6883 , n6832 );
not ( n6884 , n6824 );
not ( n6885 , n6884 );
or ( n6886 , n6883 , n6885 );
nand ( n6887 , n6824 , n6831 );
nand ( n6888 , n6886 , n6887 );
and ( n6889 , n6888 , n6845 );
not ( n6890 , n6888 );
not ( n6891 , n6845 );
and ( n6892 , n6890 , n6891 );
nor ( n6893 , n6889 , n6892 );
not ( n6894 , n6893 );
not ( n6895 , n6862 );
not ( n6896 , n6868 );
not ( n6897 , n6896 );
or ( n6898 , n6895 , n6897 );
nand ( n6899 , n6868 , n5432 );
nand ( n6900 , n6898 , n6899 );
not ( n6901 , n6900 );
nor ( n6902 , n6901 , n6880 );
or ( n6903 , n6894 , n6902 );
nand ( n6904 , n6882 , n6903 );
not ( n6905 , n6904 );
not ( n6906 , n52998 );
not ( n6907 , n53047 );
not ( n6908 , n6907 );
or ( n6909 , n6906 , n6908 );
not ( n6910 , n52998 );
nand ( n6911 , n6910 , n53047 );
nand ( n6912 , n6909 , n6911 );
and ( n6913 , n6912 , n6796 );
not ( n6914 , n6912 );
not ( n6915 , n6796 );
and ( n6916 , n6914 , n6915 );
nor ( n6917 , n6913 , n6916 );
nand ( n6918 , n6905 , n6917 );
buf ( n53109 , n6918 );
not ( n6920 , n53109 );
buf ( n53111 , n6920 );
buf ( n53112 , n53111 );
and ( n6923 , n6880 , n6869 );
not ( n6924 , n6880 );
and ( n6925 , n6924 , n6900 );
nor ( n6926 , n6923 , n6925 );
and ( n6927 , n6926 , n6894 );
not ( n6928 , n6926 );
and ( n6929 , n6928 , n6893 );
nor ( n6930 , n6927 , n6929 );
not ( n6931 , n6930 );
not ( n6932 , n51733 );
not ( n6933 , n6932 );
not ( n6934 , n52131 );
or ( n6935 , n6933 , n6934 );
not ( n6936 , n51733 );
not ( n6937 , n52125 );
or ( n6938 , n6936 , n6937 );
nand ( n6939 , n6938 , n52014 );
nand ( n6940 , n6935 , n6939 );
nor ( n6941 , n6931 , n6940 );
buf ( n53132 , n6941 );
nor ( n6943 , n53112 , n53132 );
buf ( n53134 , n6943 );
buf ( n53135 , n53134 );
and ( n6946 , n53051 , n53135 );
buf ( n53137 , n6946 );
not ( n6948 , n53137 );
or ( n6949 , n6788 , n6948 );
not ( n6950 , n6860 );
not ( n6951 , n6932 );
not ( n6952 , n52131 );
or ( n6953 , n6951 , n6952 );
nand ( n6954 , n6953 , n6939 );
not ( n6955 , n6954 );
nor ( n6956 , n6955 , n6930 );
not ( n6957 , n6956 );
not ( n6958 , n6918 );
or ( n6959 , n6957 , n6958 );
buf ( n53150 , n6917 );
not ( n6961 , n53150 );
buf ( n6962 , n6904 );
buf ( n53153 , n6962 );
nand ( n6964 , n6961 , n53153 );
buf ( n53155 , n6964 );
nand ( n6966 , n6959 , n53155 );
not ( n6967 , n6966 );
or ( n6968 , n6950 , n6967 );
buf ( n53159 , n52984 );
not ( n6970 , n53159 );
buf ( n53161 , n6970 );
buf ( n53162 , n6859 );
not ( n6973 , n53162 );
buf ( n53164 , n6973 );
nand ( n6975 , n53161 , n53164 );
nand ( n6976 , n6968 , n6975 );
not ( n6977 , n6976 );
nand ( n6978 , n6949 , n6977 );
and ( n6979 , n51675 , n6978 );
not ( n6980 , n6979 );
or ( n6981 , n4946 , n6980 );
not ( n6982 , n50491 );
not ( n6983 , n50469 );
and ( n6984 , n6982 , n6983 );
and ( n6985 , n50491 , n50469 );
nor ( n6986 , n6985 , n4722 );
nor ( n6987 , n6984 , n6986 );
nor ( n6988 , n50462 , n6987 );
not ( n6989 , n6988 );
buf ( n53180 , n4677 );
buf ( n53181 , n50382 );
nand ( n6992 , n53180 , n53181 );
buf ( n53183 , n6992 );
buf ( n53184 , n53183 );
nand ( n6995 , n4733 , n4746 );
buf ( n53186 , n6995 );
and ( n6997 , n53184 , n53186 );
buf ( n53188 , n6997 );
not ( n6999 , n53188 );
buf ( n53190 , n50382 );
not ( n7001 , n53190 );
buf ( n53192 , n50453 );
nand ( n7003 , n7001 , n53192 );
buf ( n53194 , n7003 );
buf ( n53195 , n50713 );
buf ( n53196 , n50707 );
nor ( n7007 , n53195 , n53196 );
buf ( n53198 , n7007 );
nand ( n7009 , n53194 , n53198 );
not ( n7010 , n7009 );
or ( n7011 , n6999 , n7010 );
and ( n7012 , n4726 , n4748 );
nand ( n7013 , n7011 , n7012 );
nand ( n7014 , n6989 , n7013 );
nor ( n7015 , n51667 , n5535 );
not ( n7016 , n7015 );
not ( n7017 , n51657 );
or ( n7018 , n7016 , n7017 );
buf ( n53209 , n51585 );
not ( n7020 , n53209 );
buf ( n53211 , n7020 );
buf ( n53212 , n53211 );
buf ( n53213 , n51651 );
nand ( n7024 , n53212 , n53213 );
buf ( n53215 , n7024 );
nand ( n7026 , n7018 , n53215 );
not ( n7027 , n7026 );
nand ( n7028 , n5240 , n5449 );
nand ( n7029 , n51101 , n5236 );
nand ( n7030 , n7028 , n7029 );
nand ( n7031 , n7030 , n5238 , n5543 , n51657 );
nand ( n7032 , n7027 , n7031 );
nor ( n7033 , n4727 , n50717 );
nand ( n7034 , n7032 , n7033 );
not ( n7035 , n7034 );
nor ( n7036 , n7014 , n7035 );
nand ( n7037 , n6981 , n7036 );
not ( n7038 , n7037 );
or ( n7039 , n4192 , n7038 );
nor ( n7040 , n49747 , n3896 );
nand ( n7041 , n4176 , n49960 );
or ( n7042 , n7040 , n7041 );
nand ( n7044 , n7042 , C1 );
buf ( n53234 , n7044 );
not ( n7046 , n53234 );
buf ( n53236 , n7046 );
nand ( n7048 , n7039 , n53236 );
buf ( n53238 , n7048 );
and ( n7050 , n53238 , n49670 );
not ( n7051 , n53238 );
and ( n7052 , n7051 , n49669 );
nor ( n7053 , n7050 , n7052 );
buf ( n53243 , n7053 );
buf ( n53244 , n6988 );
not ( n7056 , n53244 );
buf ( n53246 , n4726 );
nand ( n7058 , n7056 , n53246 );
buf ( n53248 , n7058 );
buf ( n53249 , n53248 );
buf ( n53250 , n53248 );
not ( n7062 , n53250 );
buf ( n53252 , n7062 );
buf ( n53253 , n53252 );
buf ( n7065 , n4748 );
not ( n7066 , n7065 );
buf ( n53256 , n4941 );
not ( n7068 , n53256 );
buf ( n53258 , n50453 );
not ( n7070 , n53258 );
buf ( n53260 , n50382 );
nor ( n7072 , n7070 , n53260 );
buf ( n53262 , n7072 );
buf ( n53263 , n53262 );
nor ( n7075 , n7068 , n53263 );
buf ( n53265 , n7075 );
buf ( n53266 , n53265 );
not ( n7078 , n53266 );
not ( n7079 , n6978 );
not ( n7080 , n51675 );
or ( n7081 , n7079 , n7080 );
not ( n7082 , n7032 );
nand ( n7083 , n7081 , n7082 );
buf ( n53273 , n7083 );
not ( n7085 , n53273 );
or ( n7086 , n7078 , n7085 );
buf ( n53276 , n53183 );
buf ( n7088 , n53276 );
buf ( n53278 , n7088 );
and ( n7090 , n7009 , n53278 );
buf ( n53280 , n7090 );
nand ( n7092 , n7086 , n53280 );
buf ( n53282 , n7092 );
not ( n7094 , n53282 );
or ( n7095 , n7066 , n7094 );
buf ( n7096 , n6995 );
nand ( n7097 , n7095 , n7096 );
buf ( n53287 , n7097 );
and ( n7099 , n53287 , n53253 );
not ( n7100 , n53287 );
and ( n7101 , n7100 , n53249 );
nor ( n7102 , n7099 , n7101 );
buf ( n53292 , n7102 );
buf ( n53293 , n4748 );
buf ( n53294 , n7096 );
nand ( n7106 , n53293 , n53294 );
buf ( n53296 , n7106 );
buf ( n53297 , n53296 );
buf ( n53298 , n53296 );
not ( n7110 , n53298 );
buf ( n53300 , n7110 );
buf ( n53301 , n53300 );
buf ( n53302 , n53282 );
and ( n7114 , n53302 , n53301 );
not ( n7115 , n53302 );
and ( n7116 , n7115 , n53297 );
nor ( n7117 , n7114 , n7116 );
buf ( n53307 , n7117 );
buf ( n53308 , n49412 );
buf ( n53309 , n49520 );
and ( n7121 , n53308 , n53309 );
buf ( n53311 , n49409 );
buf ( n53312 , n49517 );
and ( n7124 , n53311 , n53312 );
nor ( n7125 , n7121 , n7124 );
buf ( n53315 , n7125 );
buf ( n53316 , n53315 );
buf ( n53317 , n49485 );
and ( n7129 , n53316 , n53317 );
not ( n7130 , n53316 );
buf ( n53320 , n49458 );
and ( n7132 , n7130 , n53320 );
or ( n7133 , n7129 , n7132 );
buf ( n53323 , n7133 );
buf ( n53324 , n53323 );
buf ( n53325 , n49412 );
and ( n7137 , n53324 , n53325 );
not ( n7138 , n53324 );
buf ( n53328 , n49409 );
and ( n7140 , n7138 , n53328 );
nor ( n7141 , n7137 , n7140 );
buf ( n53331 , n7141 );
buf ( n53332 , n53331 );
not ( n7144 , n53332 );
buf ( n53334 , n49412 );
buf ( n53335 , n49517 );
or ( n7147 , n53334 , n53335 );
buf ( n53337 , n49409 );
buf ( n53338 , n49520 );
or ( n7150 , n53337 , n53338 );
buf ( n53340 , n49458 );
nand ( n7152 , n7150 , n53340 );
buf ( n53342 , n7152 );
buf ( n53343 , n53342 );
nand ( n7155 , n7147 , n53343 );
buf ( n53345 , n7155 );
buf ( n53346 , n53345 );
not ( n7158 , n53346 );
and ( n7159 , n7144 , n7158 );
buf ( n53349 , n53331 );
buf ( n53350 , n53345 );
and ( n7162 , n53349 , n53350 );
nor ( n7163 , n7159 , n7162 );
buf ( n53353 , n7163 );
buf ( n53354 , n49924 );
buf ( n53355 , n49517 );
nand ( n7168 , n53354 , n53355 );
buf ( n53357 , n7168 );
buf ( n53358 , n53357 );
not ( n7171 , n53358 );
buf ( n53360 , n7171 );
not ( n7173 , n53360 );
not ( n7174 , n53323 );
and ( n7175 , n7173 , n7174 );
buf ( n53364 , n53323 );
buf ( n53365 , n53360 );
nand ( n7178 , n53364 , n53365 );
buf ( n53367 , n7178 );
buf ( n53368 , n5618 );
not ( n7181 , n53368 );
buf ( n53370 , n49409 );
buf ( n53371 , n49485 );
nand ( n7184 , n53370 , n53371 );
buf ( n53373 , n7184 );
buf ( n53374 , n53373 );
not ( n7187 , n53374 );
or ( n7188 , n7181 , n7187 );
buf ( n53377 , n49466 );
nand ( n7190 , n7188 , n53377 );
buf ( n53379 , n7190 );
and ( n7192 , n53367 , n53379 );
nor ( n7193 , n7175 , n7192 );
buf ( n53382 , n49415 );
not ( n7200 , n53382 );
buf ( n53384 , n3786 );
nand ( n7202 , n7200 , n53384 );
buf ( n53386 , n7202 );
not ( n7204 , n53386 );
not ( n7205 , n4148 );
not ( n7206 , n49520 );
or ( n7207 , n7205 , n7206 );
nand ( n7208 , n7207 , n53357 );
not ( n7209 , n7208 );
or ( n7210 , n7204 , n7209 );
buf ( n53394 , n49418 );
buf ( n53395 , n3868 );
nand ( n7213 , n53394 , n53395 );
buf ( n53397 , n7213 );
nand ( n7215 , n7210 , n53397 );
buf ( n53399 , n7215 );
buf ( n53400 , n53379 );
buf ( n53401 , n53323 );
xor ( n7219 , n53400 , n53401 );
buf ( n53403 , n53357 );
xnor ( n7221 , n7219 , n53403 );
buf ( n53405 , n7221 );
buf ( n53406 , n53405 );
or ( n7224 , n53399 , n53406 );
buf ( n53408 , n7224 );
buf ( n53409 , n53408 );
not ( n7227 , n53409 );
buf ( n53411 , n49492 );
buf ( n53412 , n49412 );
and ( n7230 , n53411 , n53412 );
not ( n7231 , n53411 );
buf ( n53415 , n49409 );
and ( n7233 , n7231 , n53415 );
nor ( n7234 , n7230 , n7233 );
buf ( n53418 , n7234 );
buf ( n53419 , n53418 );
buf ( n53420 , n53386 );
buf ( n53421 , n49537 );
nand ( n7239 , n53420 , n53421 );
buf ( n53423 , n7239 );
buf ( n53424 , n53423 );
buf ( n53425 , n53397 );
nand ( n7243 , n53424 , n53425 );
buf ( n53427 , n7243 );
buf ( n53428 , n53427 );
xor ( n7246 , n53419 , n53428 );
buf ( n53430 , n7208 );
not ( n7248 , n53430 );
buf ( n53432 , n7248 );
buf ( n53433 , n53432 );
not ( n7251 , n53433 );
buf ( n53435 , n49574 );
not ( n7253 , n53435 );
or ( n7254 , n7251 , n7253 );
buf ( n53438 , n49574 );
buf ( n53439 , n53432 );
or ( n7257 , n53438 , n53439 );
nand ( n7258 , n7254 , n7257 );
buf ( n53442 , n7258 );
buf ( n53443 , n53442 );
and ( n7261 , n7246 , n53443 );
and ( n7262 , n53419 , n53428 );
or ( n7263 , n7261 , n7262 );
buf ( n53447 , n7263 );
buf ( n53448 , n53447 );
not ( n7266 , n53448 );
or ( n7267 , n7227 , n7266 );
buf ( n53451 , n7215 );
buf ( n53452 , n53405 );
nand ( n7270 , n53451 , n53452 );
buf ( n53454 , n7270 );
buf ( n53455 , n53454 );
nand ( n7273 , n7267 , n53455 );
buf ( n53457 , n7273 );
buf ( n53458 , n53457 );
not ( n7276 , n53458 );
or ( n7277 , C0 , n7276 );
buf ( n53461 , n7193 );
buf ( n53462 , n53353 );
nor ( n7280 , n53461 , n53462 );
buf ( n53464 , n7280 );
buf ( n53465 , n53464 );
not ( n7283 , n53465 );
buf ( n53467 , n7283 );
buf ( n53468 , n53467 );
nand ( n7286 , n7277 , n53468 );
buf ( n53470 , n7286 );
buf ( n53471 , n46229 );
not ( n7289 , n53471 );
buf ( n53473 , n7289 );
buf ( n53474 , n53473 );
buf ( n53475 , n415 );
buf ( n53476 , n416 );
and ( n7294 , n53475 , n53476 );
buf ( n53478 , n46115 );
not ( n7296 , n53478 );
buf ( n53480 , n7296 );
buf ( n53481 , n53480 );
nor ( n7299 , n7294 , n53481 );
buf ( n53483 , n7299 );
buf ( n53484 , n53483 );
or ( n7302 , n53474 , n53484 );
buf ( n53486 , n46241 );
nand ( n7304 , n7302 , n53486 );
buf ( n53488 , n7304 );
buf ( n53489 , n53488 );
buf ( n53490 , n46234 );
xor ( n7308 , n53489 , n53490 );
buf ( n53492 , n3404 );
buf ( n53493 , n415 );
and ( n7311 , n53492 , n53493 );
not ( n7312 , n53492 );
buf ( n53496 , n46124 );
and ( n7314 , n7312 , n53496 );
nor ( n7315 , n7311 , n7314 );
buf ( n53499 , n7315 );
buf ( n53500 , n53499 );
not ( n7318 , n53500 );
buf ( n53502 , n3296 );
not ( n7320 , n53502 );
or ( n7321 , n7318 , n7320 );
buf ( n53505 , n3296 );
buf ( n53506 , n53499 );
or ( n7324 , n53505 , n53506 );
nand ( n7325 , n7321 , n7324 );
buf ( n53509 , n7325 );
buf ( n53510 , n53509 );
and ( n7328 , n7308 , n53510 );
and ( n7329 , n53489 , n53490 );
or ( n7330 , n7328 , n7329 );
buf ( n53514 , n7330 );
buf ( n53515 , n53514 );
buf ( n53516 , n49150 );
buf ( n53517 , n53499 );
or ( n7335 , n53516 , n53517 );
buf ( n53519 , n46102 );
buf ( n53520 , n46214 );
or ( n7338 , n53519 , n53520 );
nand ( n7339 , n7335 , n7338 );
buf ( n53523 , n7339 );
buf ( n53524 , n53523 );
buf ( n53525 , n46199 );
xor ( n7343 , n53524 , n53525 );
buf ( n53527 , n46238 );
not ( n7345 , n46157 );
buf ( n53529 , n7345 );
buf ( n53530 , n46180 );
or ( n7348 , n53529 , n53530 );
buf ( n53532 , n46176 );
buf ( n53533 , n46153 );
or ( n7351 , n53532 , n53533 );
nand ( n7352 , n7348 , n7351 );
buf ( n53536 , n7352 );
buf ( n53537 , n53536 );
xor ( n7355 , n53527 , n53537 );
buf ( n53539 , n46199 );
buf ( n53540 , n415 );
nor ( n7358 , n53539 , n53540 );
buf ( n53542 , n7358 );
buf ( n53543 , n53542 );
xor ( n7361 , n7355 , n53543 );
buf ( n53545 , n7361 );
buf ( n53546 , n53545 );
xor ( n7364 , n7343 , n53546 );
buf ( n53548 , n7364 );
buf ( n53549 , n53548 );
xor ( n7367 , n53515 , n53549 );
xor ( n7368 , n53489 , n53490 );
xor ( n7369 , n7368 , n53510 );
buf ( n53553 , n7369 );
buf ( n53554 , n53553 );
not ( n7372 , n53554 );
buf ( n53556 , n53483 );
buf ( n53557 , n46238 );
and ( n7375 , n53556 , n53557 );
not ( n7376 , n53556 );
buf ( n53560 , n46102 );
and ( n7378 , n7376 , n53560 );
nor ( n7379 , n7375 , n7378 );
buf ( n53563 , n7379 );
xor ( n7381 , n53563 , n46234 );
buf ( n53565 , n7381 );
buf ( n53566 , n46223 );
xor ( n7384 , n53565 , n53566 );
buf ( n53568 , n46264 );
and ( n7386 , n7384 , n53568 );
and ( n7387 , n53565 , n53566 );
or ( n7388 , n7386 , n7387 );
buf ( n53572 , n7388 );
buf ( n53573 , n53572 );
nand ( n7391 , n7372 , n53573 );
buf ( n53575 , n7391 );
buf ( n53576 , n53575 );
not ( n7394 , n53576 );
xor ( n7395 , n53565 , n53566 );
xor ( n7396 , n7395 , n53568 );
buf ( n53580 , n7396 );
buf ( n53581 , n53580 );
buf ( n53582 , n46249 );
nand ( n7400 , n53581 , n53582 );
buf ( n53584 , n7400 );
not ( n7402 , n53584 );
buf ( n53586 , n3591 );
buf ( n7404 , n53586 );
buf ( n53588 , n7404 );
not ( n7406 , n53588 );
or ( n7407 , n7402 , n7406 );
buf ( n53591 , n53580 );
not ( n7409 , n53591 );
buf ( n53593 , n46246 );
nand ( n7411 , n7409 , n53593 );
buf ( n53595 , n7411 );
nand ( n7413 , n7407 , n53595 );
buf ( n53597 , n7413 );
not ( n7415 , n53597 );
or ( n7416 , n7394 , n7415 );
buf ( n53600 , n53572 );
not ( n7418 , n53600 );
buf ( n53602 , n53553 );
nand ( n7420 , n7418 , n53602 );
buf ( n53604 , n7420 );
buf ( n53605 , n53604 );
nand ( n7423 , n7416 , n53605 );
buf ( n53607 , n7423 );
buf ( n53608 , n53607 );
xor ( n7426 , n7367 , n53608 );
buf ( n53610 , n7426 );
not ( n7428 , n53610 );
buf ( n53612 , C1 );
buf ( n53613 , n53612 );
buf ( n53614 , n53470 );
buf ( n53615 , n7428 );
nand ( n7436 , n53614 , n53615 );
buf ( n53617 , n7436 );
buf ( n53618 , n53617 );
nand ( n7439 , n53613 , n53618 );
buf ( n53620 , n7439 );
buf ( n53621 , n53620 );
buf ( n53622 , n53620 );
not ( n7443 , n53622 );
buf ( n53624 , n7443 );
buf ( n53625 , n53624 );
buf ( n53626 , n53604 );
buf ( n53627 , n53575 );
nand ( n7448 , n53626 , n53627 );
buf ( n53629 , n7448 );
xnor ( n7450 , n53629 , n7413 );
buf ( n53631 , n7450 );
not ( n7452 , n53631 );
xor ( n7453 , n53353 , n7193 );
xnor ( n7454 , n7453 , n53457 );
buf ( n53635 , n7454 );
nand ( n7456 , n7452 , n53635 );
buf ( n53637 , n7456 );
buf ( n53638 , n53637 );
and ( n7459 , n53595 , n53584 );
xor ( n7460 , n7459 , n53588 );
buf ( n53641 , n7460 );
not ( n7462 , n53641 );
buf ( n53643 , n53447 );
buf ( n7464 , n53643 );
buf ( n53645 , n7464 );
buf ( n53646 , n53645 );
buf ( n53647 , n7215 );
buf ( n53648 , n53405 );
xor ( n7469 , n53647 , n53648 );
buf ( n53650 , n7469 );
buf ( n53651 , n53650 );
xnor ( n7472 , n53646 , n53651 );
buf ( n53653 , n7472 );
buf ( n53654 , n53653 );
nand ( n7475 , n7462 , n53654 );
buf ( n53656 , n7475 );
buf ( n53657 , n53656 );
not ( n7478 , n49546 );
not ( n7479 , n49574 );
or ( n7480 , n7478 , n7479 );
nand ( n7481 , n7480 , n49580 );
not ( n7482 , n7481 );
nand ( n7483 , n7482 , n3748 );
not ( n7484 , n7483 );
buf ( n53665 , n53427 );
buf ( n7486 , n53665 );
buf ( n53667 , n7486 );
not ( n7488 , n53667 );
or ( n7489 , n7484 , n7488 );
buf ( n53670 , n7481 );
buf ( n53671 , n3747 );
nand ( n7492 , n53670 , n53671 );
buf ( n53673 , n7492 );
nand ( n7494 , n7489 , n53673 );
xor ( n7495 , n53419 , n53428 );
xor ( n7496 , n7495 , n53443 );
buf ( n53677 , n7496 );
or ( n7498 , n7494 , n53677 );
buf ( n53679 , n7498 );
and ( n7500 , n53638 , n53657 , n53679 );
buf ( n53681 , n7500 );
not ( n7502 , n53681 );
not ( n7503 , n7483 );
not ( n7504 , n49543 );
or ( n7505 , n7503 , n7504 );
nand ( n7506 , n7505 , n53673 );
not ( n7507 , n7506 );
not ( n7508 , n53667 );
not ( n7509 , n49588 );
or ( n7510 , n7508 , n7509 );
buf ( n53691 , n53667 );
not ( n7512 , n53691 );
buf ( n53693 , n3808 );
nand ( n7514 , n7512 , n53693 );
buf ( n53695 , n7514 );
nand ( n7516 , n7510 , n53695 );
not ( n7517 , n7516 );
and ( n7518 , n7507 , n7517 );
not ( n7519 , n3815 );
not ( n7520 , n3883 );
and ( n7521 , n7519 , n7520 );
nor ( n7522 , n7518 , n7521 );
and ( n7523 , n3972 , n7522 , n49962 );
not ( n7524 , n7523 );
nor ( n7525 , n7524 , n4727 );
nor ( n7526 , n5547 , n50717 );
nand ( n7527 , n6978 , n7525 , n7526 );
not ( n7528 , n7522 );
not ( n7529 , n7044 );
or ( n7530 , n7528 , n7529 );
nand ( n7535 , n7530 , C1 );
buf ( n53712 , n7535 );
buf ( n53713 , n6988 );
nor ( n7538 , n53712 , n53713 );
buf ( n53715 , n7538 );
nand ( n7540 , n7013 , n53715 );
or ( n7541 , n7035 , n7540 );
not ( n7542 , n7535 );
not ( n7543 , n7523 );
and ( n7544 , n7542 , n7543 );
nor ( n7545 , n7494 , n7516 );
nor ( n7546 , n7544 , n7545 );
nand ( n7547 , n7541 , n7546 );
nand ( n7548 , n7527 , n7547 );
not ( n7549 , n7548 );
or ( n7550 , n7502 , n7549 );
buf ( n53727 , C0 );
buf ( n53728 , C1 );
nand ( n7581 , n7550 , C1 );
buf ( n53730 , n7581 );
and ( n7583 , n53730 , n53625 );
not ( n7584 , n53730 );
and ( n7585 , n7584 , n53621 );
nor ( n7586 , n7583 , n7585 );
buf ( n53735 , n7586 );
buf ( n53736 , n53262 );
not ( n7589 , n53736 );
buf ( n53738 , n53278 );
nand ( n7591 , n7589 , n53738 );
buf ( n53740 , n7591 );
buf ( n53741 , n53740 );
buf ( n53742 , n53740 );
not ( n7595 , n53742 );
buf ( n53744 , n7595 );
buf ( n53745 , n53744 );
not ( n7598 , n4941 );
not ( n7599 , n7083 );
or ( n7600 , n7598 , n7599 );
not ( n7601 , n53198 );
nand ( n7602 , n7600 , n7601 );
buf ( n53751 , n7602 );
and ( n7604 , n53751 , n53745 );
not ( n7605 , n53751 );
and ( n7606 , n7605 , n53741 );
nor ( n7607 , n7604 , n7606 );
buf ( n53756 , n7607 );
buf ( n7609 , n7015 );
not ( n7610 , n7609 );
buf ( n7611 , n5543 );
nand ( n7612 , n7610 , n7611 );
buf ( n53761 , n7612 );
buf ( n53762 , n7612 );
not ( n7615 , n53762 );
buf ( n53764 , n7615 );
buf ( n53765 , n53764 );
not ( n7618 , n6978 );
not ( n7619 , n5454 );
or ( n7620 , n7618 , n7619 );
buf ( n7621 , n5238 );
buf ( n7622 , n7030 );
nand ( n7623 , n7621 , n7622 );
nand ( n7624 , n7620 , n7623 );
buf ( n53773 , n7624 );
and ( n7626 , n53773 , n53765 );
not ( n7627 , n53773 );
and ( n7628 , n7627 , n53761 );
nor ( n7629 , n7626 , n7628 );
buf ( n53778 , n7629 );
buf ( n53779 , n7601 );
buf ( n53780 , n4941 );
nand ( n7633 , n53779 , n53780 );
buf ( n53782 , n7633 );
buf ( n53783 , n53782 );
buf ( n53784 , n53782 );
not ( n7637 , n53784 );
buf ( n53786 , n7637 );
buf ( n53787 , n53786 );
buf ( n53788 , n7083 );
and ( n7641 , n53788 , n53787 );
not ( n7642 , n53788 );
and ( n7643 , n7642 , n53783 );
nor ( n7644 , n7641 , n7643 );
buf ( n53793 , n7644 );
buf ( n53794 , n6860 );
buf ( n53795 , n6975 );
nand ( n7648 , n53794 , n53795 );
buf ( n53797 , n7648 );
buf ( n53798 , n53797 );
buf ( n53799 , n53797 );
not ( n7652 , n53799 );
buf ( n53801 , n7652 );
buf ( n53802 , n53801 );
buf ( n53803 , n53111 );
not ( n7656 , n53803 );
buf ( n53805 , n7656 );
buf ( n53806 , n53805 );
not ( n7659 , n53806 );
buf ( n53808 , n6941 );
not ( n7661 , n53808 );
buf ( n53810 , n7661 );
not ( n7663 , n53810 );
not ( n7664 , n52244 );
not ( n7665 , n52970 );
or ( n7666 , n7664 , n7665 );
nand ( n7667 , n7666 , n52976 );
not ( n7668 , n7667 );
or ( n7669 , n7663 , n7668 );
buf ( n53818 , n6956 );
not ( n7671 , n53818 );
buf ( n53820 , n7671 );
nand ( n7673 , n7669 , n53820 );
buf ( n53822 , n7673 );
not ( n7675 , n53822 );
or ( n7676 , n7659 , n7675 );
buf ( n53825 , n53155 );
buf ( n7678 , n53825 );
buf ( n53827 , n7678 );
buf ( n53828 , n53827 );
nand ( n7681 , n7676 , n53828 );
buf ( n53830 , n7681 );
buf ( n53831 , n53830 );
and ( n7684 , n53831 , n53802 );
not ( n7685 , n53831 );
and ( n7686 , n7685 , n53798 );
nor ( n7687 , n7684 , n7686 );
buf ( n53836 , n7687 );
nand ( n7689 , n7621 , n7029 );
buf ( n53838 , n7689 );
buf ( n53839 , n7689 );
not ( n7692 , n53839 );
buf ( n53841 , n7692 );
buf ( n53842 , n53841 );
buf ( n7695 , n5453 );
buf ( n7696 , n7695 );
not ( n7697 , n7696 );
buf ( n7698 , n6978 );
not ( n7699 , n7698 );
or ( n7700 , n7697 , n7699 );
buf ( n7701 , n7028 );
nand ( n7702 , n7700 , n7701 );
buf ( n53851 , n7702 );
and ( n7704 , n53851 , n53842 );
not ( n7705 , n53851 );
and ( n7706 , n7705 , n53838 );
nor ( n7707 , n7704 , n7706 );
buf ( n53856 , n7707 );
buf ( n53857 , n52976 );
buf ( n7710 , n52244 );
buf ( n53859 , n7710 );
nand ( n7712 , n53857 , n53859 );
buf ( n53861 , n7712 );
buf ( n53862 , n53861 );
not ( n7715 , n53862 );
buf ( n53864 , n7715 );
buf ( n53865 , n53864 );
buf ( n53866 , n53861 );
buf ( n53867 , n52876 );
not ( n7720 , n53867 );
buf ( n53869 , n52948 );
not ( n7722 , n53869 );
or ( n7723 , n7720 , n7722 );
buf ( n53872 , n52967 );
nand ( n7725 , n7723 , n53872 );
buf ( n53874 , n7725 );
buf ( n53875 , n53874 );
not ( n7728 , n53875 );
buf ( n53877 , n7728 );
buf ( n53878 , n53877 );
and ( n7731 , n53878 , n53866 );
not ( n7732 , n53878 );
and ( n7733 , n7732 , n53865 );
nor ( n7734 , n7731 , n7733 );
buf ( n53883 , n7734 );
nand ( n7736 , n6773 , n6744 );
buf ( n53885 , n7736 );
buf ( n7738 , n6755 );
buf ( n53887 , n7738 );
not ( n7740 , n53887 );
buf ( n53889 , n52876 );
buf ( n7742 , n53889 );
buf ( n53891 , n7742 );
buf ( n53892 , n53891 );
not ( n7745 , n53892 );
or ( n7746 , n7740 , n7745 );
buf ( n7747 , n52955 );
buf ( n53896 , n7747 );
nand ( n7749 , n7746 , n53896 );
buf ( n53898 , n7749 );
buf ( n53899 , n53898 );
buf ( n53900 , n7736 );
buf ( n53901 , n53898 );
not ( n7754 , n53885 );
not ( n7755 , n53899 );
or ( n7756 , n7754 , n7755 );
or ( n7757 , n53900 , n53901 );
nand ( n7758 , n7756 , n7757 );
buf ( n53907 , n7758 );
nand ( n7760 , n7738 , n7747 );
buf ( n53909 , n7760 );
buf ( n53910 , n53891 );
buf ( n53911 , n53891 );
buf ( n53912 , n7760 );
not ( n7765 , n53909 );
not ( n7766 , n53910 );
or ( n7767 , n7765 , n7766 );
or ( n7768 , n53911 , n53912 );
nand ( n7769 , n7767 , n7768 );
buf ( n53918 , n7769 );
or ( n7771 , n45489 , n46852 );
not ( n7772 , n46101 );
or ( n7773 , n7772 , n45497 );
nand ( n7774 , n7771 , n7773 );
xor ( n7775 , n7774 , n46199 );
nand ( n7776 , n46181 , n413 );
xor ( n7777 , n3404 , n7776 );
and ( n7778 , n7777 , n46238 );
and ( n7779 , n3404 , n7776 );
or ( n7780 , n7778 , n7779 );
and ( n7781 , n7775 , n7780 );
and ( n7782 , n7774 , n46199 );
or ( n7783 , n7781 , n7782 );
nand ( n7784 , n45498 , n411 );
xnor ( n7785 , n7783 , n7784 );
not ( n7786 , n7785 );
xor ( n7787 , n3404 , n7776 );
xor ( n7788 , n7787 , n46238 );
xor ( n7789 , n7788 , n3404 );
xor ( n7790 , n53527 , n53537 );
and ( n7791 , n7790 , n53543 );
and ( n7792 , n53527 , n53537 );
or ( n7793 , n7791 , n7792 );
buf ( n53942 , n7793 );
and ( n7795 , n7789 , n53942 );
and ( n7796 , n7788 , n3404 );
or ( n7797 , n7795 , n7796 );
xor ( n7798 , n7774 , n46199 );
xor ( n7799 , n7798 , n7780 );
nor ( n7800 , n7797 , n7799 );
not ( n7801 , n7800 );
xor ( n7802 , n53515 , n53549 );
and ( n7803 , n7802 , n53608 );
and ( n7804 , n53515 , n53549 );
or ( n7805 , n7803 , n7804 );
buf ( n53954 , n7805 );
buf ( n7807 , n53954 );
xor ( n7808 , n53524 , n53525 );
and ( n7809 , n7808 , n53546 );
and ( n7810 , n53524 , n53525 );
or ( n7811 , n7809 , n7810 );
buf ( n53960 , n7811 );
not ( n7813 , n53960 );
xor ( n7814 , n7788 , n3404 );
xor ( n7815 , n7814 , n53942 );
not ( n7816 , n7815 );
nand ( n7817 , n7813 , n7816 );
nand ( n7818 , n7801 , n7807 , n7817 );
not ( n7819 , n7800 );
nand ( n7820 , n7819 , n53960 , n7815 );
nand ( n7821 , n7797 , n7799 );
nand ( n7822 , n7818 , n7820 , n7821 );
not ( n7823 , n7822 );
or ( n7824 , n7786 , n7823 );
or ( n7825 , n7822 , n7785 );
nand ( n7826 , n7824 , n7825 );
not ( n7827 , n7826 );
not ( n7829 , n53457 );
or ( n7830 , C0 , n7829 );
nor ( n7850 , C0 , n53464 );
nand ( n7851 , n7830 , n7850 );
nand ( n53980 , n7827 , n7851 );
buf ( n53981 , n53980 );
not ( n53982 , n7817 );
not ( n7855 , n7807 );
or ( n53984 , n53982 , n7855 );
nand ( n7857 , n53960 , n7815 );
nand ( n53986 , n53984 , n7857 );
not ( n7859 , n7799 );
nand ( n53988 , n7859 , n7797 );
nor ( n7861 , n53986 , n53988 );
not ( n53990 , n7797 );
nand ( n7863 , n53990 , n7799 );
nor ( n53992 , n53986 , n7863 );
nor ( n7865 , n7861 , n53992 );
not ( n53994 , n7821 );
or ( n7867 , n53994 , n7800 );
nand ( n53996 , n7867 , n53986 );
nand ( n7869 , n7865 , n53996 );
not ( n53998 , n7869 );
nand ( n7871 , n53998 , n7851 );
buf ( n54000 , n7871 );
nand ( n7873 , n53981 , n54000 );
buf ( n54002 , n7873 );
nand ( n54003 , n7807 , n53960 , n7815 );
not ( n7877 , n7817 );
nand ( n54005 , n7877 , n7807 );
not ( n7879 , n7807 );
nand ( n54007 , n7879 , n53960 , n7816 );
nand ( n7881 , n7879 , n7813 , n7815 );
nand ( n54009 , n54003 , n54005 , n54007 , n7881 );
buf ( n54010 , n54009 );
not ( n54011 , n54010 );
buf ( n54012 , n7851 );
nand ( n54013 , n54011 , n54012 );
buf ( n54014 , n54013 );
buf ( n54015 , n54014 );
buf ( n54016 , n53617 );
nand ( n54017 , n54015 , n54016 );
buf ( n54018 , n54017 );
buf ( n54019 , n54018 );
not ( n7893 , n54019 );
buf ( n54021 , n7893 );
not ( n54022 , n7851 );
buf ( n54023 , C1 );
buf ( n54024 , C1 );
or ( n7923 , n7783 , n7784 );
not ( n7924 , n7923 );
not ( n7925 , n7822 );
or ( n7926 , n7924 , n7925 );
nand ( n7927 , n7783 , n7784 );
nand ( n7928 , n7926 , n7927 );
not ( n7929 , n46197 );
and ( n7930 , n3404 , n7929 );
nor ( n7931 , n7928 , n7930 );
buf ( n54034 , n7931 );
not ( n7933 , n54034 );
buf ( n54036 , n7928 );
buf ( n54037 , n7930 );
nand ( n7936 , n54036 , n54037 );
buf ( n54039 , n7936 );
buf ( n54040 , n54039 );
nand ( n7939 , n7933 , n54040 );
buf ( n54042 , n7939 );
xnor ( n7946 , n7929 , n7931 );
or ( n7957 , n7946 , n54022 );
buf ( n54045 , n7957 );
buf ( n54046 , n54022 );
buf ( n54047 , n54042 );
or ( n7961 , n54046 , n54047 );
buf ( n54049 , n7961 );
buf ( n54050 , n54049 );
nand ( n7964 , n54045 , n54050 );
buf ( n54052 , n7964 );
buf ( n54053 , C1 );
buf ( n54054 , n53810 );
buf ( n54055 , n53820 );
nand ( n7971 , n54054 , n54055 );
buf ( n54057 , n7971 );
buf ( n54058 , n54057 );
not ( n54059 , n54058 );
buf ( n54060 , n54059 );
nor ( n54061 , n54002 , n54018 );
buf ( n54062 , n54061 );
buf ( n54063 , n53681 );
nand ( n7979 , n54062 , n54063 );
buf ( n54065 , n7979 );
buf ( n54066 , n54065 );
buf ( n54067 , n54052 );
nor ( n7983 , n54066 , n54067 );
buf ( n54069 , n7983 );
buf ( n54070 , n54065 );
not ( n54071 , n54070 );
buf ( n54072 , n54071 );
buf ( n54073 , C0 );
nor ( n54074 , C0 , n54073 );
buf ( n54075 , n54074 );
buf ( n54076 , n52868 );
buf ( n54077 , n52653 );
nand ( n54078 , n54076 , n54077 );
buf ( n54079 , n54078 );
buf ( n54080 , n54079 );
buf ( n54081 , n6670 );
buf ( n54082 , n54081 );
buf ( n54083 , n54082 );
buf ( n54084 , n54083 );
buf ( n54085 , n54083 );
buf ( n54086 , n54079 );
not ( n54087 , n54080 );
not ( n54088 , n54084 );
or ( n54089 , n54087 , n54088 );
or ( n54090 , n54085 , n54086 );
nand ( n54091 , n54089 , n54090 );
buf ( n54092 , n54091 );
buf ( n54093 , n54023 );
buf ( n54094 , n54014 );
nand ( n54095 , n54093 , n54094 );
buf ( n54096 , n54095 );
buf ( n54097 , n54096 );
not ( n54098 , n54097 );
buf ( n54099 , n54098 );
buf ( n54100 , n53980 );
buf ( n54101 , C1 );
nand ( n54102 , n54100 , n54101 );
buf ( n54103 , n54102 );
buf ( n54104 , n54103 );
not ( n54105 , n54104 );
buf ( n54106 , n54105 );
buf ( n54107 , C1 );
buf ( n54108 , n6669 );
buf ( n54109 , n6490 );
and ( n54110 , n54108 , n54109 );
buf ( n54111 , n54110 );
buf ( n54112 , n6658 );
buf ( n54113 , n6654 );
nand ( n54114 , n54112 , n54113 );
buf ( n54115 , n54114 );
buf ( n54116 , C1 );
buf ( n54117 , n7498 );
buf ( n54118 , C1 );
nand ( n54119 , n54117 , n54118 );
buf ( n54120 , n54119 );
xor ( n54121 , n52713 , n52758 );
xor ( n54122 , n54121 , n52792 );
buf ( n54123 , n54122 );
xor ( n54124 , n52776 , n52780 );
xor ( n54125 , n54124 , n52787 );
buf ( n54126 , n54125 );
buf ( n54127 , n54111 );
buf ( n54128 , n6659 );
xor ( n54129 , n54127 , n54128 );
buf ( n54130 , n54129 );
buf ( n54131 , n54115 );
buf ( n54132 , n6641 );
xnor ( n8056 , n54131 , n54132 );
buf ( n54134 , n8056 );
buf ( n54135 , n51657 );
buf ( n54136 , n53215 );
nand ( n8060 , n54135 , n54136 );
buf ( n54138 , n8060 );
buf ( n54139 , n7545 );
buf ( n54140 , C1 );
not ( n8064 , n54139 );
nand ( n8065 , n8064 , n54140 );
buf ( n54143 , n8065 );
xor ( n8067 , n52466 , n52520 );
xor ( n8068 , n8067 , n52872 );
buf ( n54146 , n8068 );
not ( n8070 , n54096 );
nand ( n54148 , n8070 , n53612 );
or ( n8072 , n7581 , n54148 );
not ( n54150 , n53617 );
nor ( n8074 , n54150 , n54099 );
nand ( n8075 , n7581 , n8074 );
nor ( n8079 , n54096 , C0 , n53617 );
nor ( n8080 , C0 , n8079 );
nand ( n8081 , n8072 , n8075 , n8080 );
buf ( n54156 , n53681 );
buf ( n54157 , n54021 );
and ( n8084 , n54156 , n54157 );
buf ( n54159 , n8084 );
and ( n8086 , n54159 , n7871 );
not ( n8087 , n8086 );
not ( n8088 , n7548 );
or ( n8089 , n8087 , n8088 );
nor ( n8093 , C0 , C0 );
nand ( n8094 , n8089 , n8093 );
and ( n8095 , n8094 , n54106 );
not ( n8096 , n8094 );
and ( n8097 , n8096 , n54103 );
nor ( n8098 , n8095 , n8097 );
and ( n8100 , n7957 , C1 );
not ( n8101 , n54072 );
not ( n8102 , n52244 );
not ( n8103 , n52970 );
or ( n8104 , n8102 , n8103 );
nand ( n8105 , n8104 , n52976 );
not ( n8106 , n8105 );
not ( n54177 , n53137 );
or ( n8108 , n8106 , n54177 );
nand ( n54179 , n8108 , n6977 );
and ( n8110 , n7526 , n54179 , n7525 );
nor ( n8112 , n8110 , C0 );
nand ( n8113 , n7547 , n8112 );
not ( n8114 , n8113 );
or ( n8115 , n8101 , n8114 );
nand ( n8116 , n8115 , n54024 );
not ( n8121 , n52799 );
nand ( n8122 , n6637 , n8121 );
or ( n8123 , n8122 , n52796 );
or ( n8124 , n6638 , n6640 );
and ( n8125 , n6638 , n52796 , n8121 );
not ( n8126 , n52796 );
and ( n8127 , n6638 , n8126 , n52799 );
nor ( n8128 , n8125 , n8127 );
nand ( n8129 , n8123 , n8124 , n8128 );
nand ( n8130 , n53728 , n53637 );
not ( n8131 , n8130 );
not ( n8132 , n54143 );
not ( n8133 , n7624 );
nor ( n8134 , n7609 , n54138 );
nand ( n8135 , n8133 , n8134 );
and ( n8136 , n7609 , n54138 );
not ( n8137 , n7609 );
nor ( n8138 , n54138 , n7611 );
and ( n8139 , n8137 , n8138 );
nor ( n8140 , n8136 , n8139 );
and ( n8141 , n7611 , n54138 );
nand ( n8142 , n8141 , n7624 );
nand ( n8143 , n8135 , n8140 , n8142 );
not ( n8144 , n8116 );
and ( n8145 , n8100 , n54107 );
nand ( n8146 , n8144 , n8145 );
nand ( n8149 , n8146 , C1 , C1 );
not ( n8150 , n53656 );
nor ( n8151 , n8150 , n8131 );
nor ( n8152 , n8130 , n53727 , n53656 );
not ( n8153 , n8113 );
and ( n8154 , n8153 , n8132 );
nor ( n8157 , n8154 , C0 );
not ( n8158 , n8157 );
not ( n8159 , n8157 );
or ( n8160 , n54022 , n54042 );
nand ( n8161 , n8160 , n54107 );
xnor ( n8162 , n8161 , n8116 );
and ( n8163 , n3972 , C1 );
not ( n8164 , n4190 );
not ( n8165 , n7037 );
or ( n8166 , n8164 , n8165 );
nand ( n8167 , n4176 , n49960 );
nand ( n8168 , n8166 , n8167 );
and ( n8169 , n8163 , n8168 );
not ( n8170 , n8163 );
and ( n8171 , n7037 , n4190 );
not ( n8172 , n8167 );
nor ( n8173 , n8171 , n8172 );
and ( n8174 , n8170 , n8173 );
nor ( n8175 , n8169 , n8174 );
not ( n8176 , n54069 );
not ( n8177 , n8113 );
or ( n8178 , n8176 , n8177 );
nand ( n8179 , n8178 , n54053 );
and ( n8180 , n8179 , n54022 );
not ( n8181 , n8179 );
and ( n8182 , n8181 , n7851 );
nor ( n8183 , n8180 , n8182 );
and ( n8184 , n7667 , n54060 );
not ( n8185 , n7667 );
and ( n8186 , n8185 , n54057 );
nor ( n8187 , n8184 , n8186 );
nand ( n8188 , n8113 , n7498 );
nand ( n8189 , n7701 , n7696 );
nand ( n8190 , n8188 , n54116 );
nand ( n8191 , C1 , n53656 );
not ( n8192 , n8191 );
and ( n8193 , n8190 , n8192 );
not ( n8194 , n8190 );
and ( n8195 , n8194 , n8191 );
nor ( n8196 , n8193 , n8195 );
nand ( n8197 , n53827 , n53805 );
not ( n8198 , n8197 );
and ( n8199 , n7673 , n8198 );
not ( n8200 , n7673 );
and ( n8201 , n8200 , n8197 );
nor ( n8202 , n8199 , n8201 );
not ( n8203 , n8151 );
or ( n8204 , n8188 , n8203 );
nor ( n8206 , C0 , n8130 );
nand ( n8207 , n8188 , n8206 );
not ( n8208 , n8131 );
and ( n8210 , n8208 , C0 );
nor ( n8211 , n8210 , n8152 );
nand ( n8212 , n8204 , n8207 , n8211 );
nand ( n8213 , n4190 , n8167 );
not ( n8214 , n8213 );
and ( n8215 , n7037 , n8214 );
not ( n8216 , n7037 );
and ( n8217 , n8216 , n8213 );
nor ( n8218 , n8215 , n8217 );
not ( n8219 , n6573 );
not ( n8220 , n401 );
and ( n8221 , n8219 , n8220 );
and ( n8222 , n6573 , n401 );
nor ( n8223 , n8221 , n8222 );
not ( n8224 , n8223 );
not ( n8225 , n52745 );
or ( n8226 , n8224 , n8225 );
or ( n8227 , n52745 , n8223 );
nand ( n8228 , n8226 , n8227 );
not ( n8229 , n54159 );
not ( n8230 , n7548 );
or ( n8231 , n8229 , n8230 );
nand ( n8232 , n8231 , n54075 );
nand ( n8233 , C1 , n7871 );
not ( n8234 , n8233 );
and ( n8235 , n8232 , n8234 );
not ( n8236 , n8232 );
and ( n8237 , n8236 , n8233 );
nor ( n8238 , n8235 , n8237 );
xor ( n8239 , n8153 , n54120 );
buf ( n54299 , n7698 );
buf ( n54300 , n8189 );
xnor ( n8242 , n54299 , n54300 );
buf ( n54302 , n8242 );
not ( C0n , n0 );
and ( C0 , C0n , n0 );
not ( C1n , n0 );
or ( C1 , C1n , n0 );
endmodule
