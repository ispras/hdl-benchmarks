//
// Conformal-LEC Version 15.10-d003 ( 23-Apr-2015) ( 64 bit executable)
//
module top ( 
    n0 , 
    n1 , 
    n2 , 
    n3 , 
    n4 , 
    n5 , 
    n6 , 
    n7 , 
    n8 , 
    n9 , 
    n10 , 
    n11 , 
    n12 , 
    n13 , 
    n14 , 
    n15 , 
    n16 , 
    n17 , 
    n18 , 
    n19 , 
    n20 , 
    n21 , 
    n22 , 
    n23 , 
    n24 , 
    n25 , 
    n26 , 
    n27 , 
    n28 , 
    n29 , 
    n30 , 
    n31 , 
    n32 , 
    n33 , 
    n34 , 
    n35 , 
    n36 , 
    n37 , 
    n38 , 
    n39 , 
    n40 , 
    n41 , 
    n42 , 
    n43 , 
    n44 , 
    n45 , 
    n46 , 
    n47 , 
    n48 , 
    n49 , 
    n50 , 
    n51 , 
    n52 , 
    n53 , 
    n54 , 
    n55 , 
    n56 , 
    n57 , 
    n58 , 
    n59 , 
    n60 , 
    n61 , 
    n62 , 
    n63 , 
    n64 , 
    n65 , 
    n66 , 
    n67 , 
    n68 , 
    n69 , 
    n70 , 
    n71 , 
    n72 , 
    n73 , 
    n74 , 
    n75 , 
    n76 , 
    n77 , 
    n78 , 
    n79 , 
    n80 , 
    n81 , 
    n82 , 
    n83 , 
    n84 , 
    n85 , 
    n86 , 
    n87 , 
    n88 , 
    n89 , 
    n90 , 
    n91 , 
    n92 , 
    n93 , 
    n94 , 
    n95 , 
    n96 , 
    n97 , 
    n98 , 
    n99 , 
    n100 , 
    n101 , 
    n102 , 
    n103 , 
    n104 , 
    n105 , 
    n106 , 
    n107 , 
    n108 , 
    n109 , 
    n110 , 
    n111 , 
    n112 , 
    n113 , 
    n114 , 
    n115 , 
    n116 , 
    n117 , 
    n118 , 
    n119 , 
    n120 , 
    n121 , 
    n122 , 
    n123 , 
    n124 , 
    n125 , 
    n126 , 
    n127 , 
    n128 , 
    n129 , 
    n130 , 
    n131 , 
    n132 , 
    n133 , 
    n134 , 
    n135 , 
    n136 , 
    n137 , 
    n138 , 
    n139 , 
    n140 , 
    n141 , 
    n142 , 
    n143 , 
    n144 , 
    n145 , 
    n146 , 
    n147 , 
    n148 , 
    n149 , 
    n150 , 
    n151 , 
    n152 , 
    n153 , 
    n154 , 
    n155 , 
    n156 , 
    n157 , 
    n158 , 
    n159 , 
    n160 , 
    n161 , 
    n162 , 
    n163 , 
    n164 , 
    n165 , 
    n166 , 
    n167 , 
    n168 , 
    n169 , 
    n170 , 
    n171 , 
    n172 , 
    n173 , 
    n174 , 
    n175 , 
    n176 , 
    n177 , 
    n178 , 
    n179 , 
    n180 , 
    n181 , 
    n182 , 
    n183 , 
    n184 , 
    n185 , 
    n186 , 
    n187 , 
    n188 , 
    n189 , 
    n190 , 
    n191 , 
    n192 , 
    n193 , 
    n194 , 
    n195 , 
    n196 , 
    n197 , 
    n198 , 
    n199 , 
    n200 , 
    n201 , 
    n202 , 
    n203 , 
    n204 , 
    n205 , 
    n206 , 
    n207 , 
    n208 , 
    n209 , 
    n210 , 
    n211 , 
    n212 , 
    n213 , 
    n214 , 
    n215 , 
    n216 , 
    n217 , 
    n218 , 
    n219 , 
    n220 , 
    n221 , 
    n222 , 
    n223 , 
    n224 , 
    n225 , 
    n226 , 
    n227 , 
    n228 , 
    n229 , 
    n230 , 
    n231 , 
    n232 , 
    n233 , 
    n234 , 
    n235 , 
    n236 , 
    n237 , 
    n238 , 
    n239 , 
    n240 , 
    n241 , 
    n242 , 
    n243 , 
    n244 , 
    n245 , 
    n246 , 
    n247 , 
    n248 , 
    n249 , 
    n250 , 
    n251 , 
    n252 , 
    n253 , 
    n254 , 
    n255 , 
    n256 , 
    n257 , 
    n258 , 
    n259 , 
    n260 , 
    n261 , 
    n262 , 
    n263 , 
    n264 , 
    n265 , 
    n266 , 
    n267 , 
    n268 , 
    n269 , 
    n270 , 
    n271 , 
    n272 , 
    n273 , 
    n274 , 
    n275 , 
    n276 , 
    n277 , 
    n278 , 
    n279 , 
    n280 , 
    n281 , 
    n282 , 
    n283 , 
    n284 , 
    n285 , 
    n286 , 
    n287 , 
    n288 , 
    n289 , 
    n290 , 
    n291 , 
    n292 , 
    n293 , 
    n294 , 
    n295 , 
    n296 , 
    n297 , 
    n298 , 
    n299 , 
    n300 , 
    n301 , 
    n302 , 
    n303 , 
    n304 , 
    n305 , 
    n306 , 
    n307 , 
    n308 , 
    n309 , 
    n310 , 
    n311 , 
    n312 , 
    n313 , 
    n314 , 
    n315 , 
    n316 , 
    n317 , 
    n318 , 
    n319 , 
    n320 , 
    n321 , 
    n322 , 
    n323 , 
    n324 , 
    n325 , 
    n326 , 
    n327 , 
    n328 , 
    n329 , 
    n330 , 
    n331 , 
    n332 , 
    n333 , 
    n334 , 
    n335 , 
    n336 , 
    n337 , 
    n338 , 
    n339 , 
    n340 , 
    n341 , 
    n342 , 
    n343 , 
    n344 , 
    n345 , 
    n346 , 
    n347 , 
    n348 , 
    n349 , 
    n350 , 
    n351 , 
    n352 , 
    n353 , 
    n354 , 
    n355 , 
    n356 , 
    n357 , 
    n358 , 
    n359 , 
    n360 , 
    n361 , 
    n362 , 
    n363 , 
    n364 , 
    n365 , 
    n366 , 
    n367 , 
    n368 , 
    n369 , 
    n370 , 
    n371 , 
    n372 , 
    n373 , 
    n374 , 
    n375 , 
    n376 , 
    n377 , 
    n378 , 
    n379 , 
    n380 , 
    n381 , 
    n382 , 
    n383 , 
    n384 , 
    n385 , 
    n386 , 
    n387 , 
    n388 , 
    n389 , 
    n390 , 
    n391 , 
    n392 , 
    n393 , 
    n394 , 
    n395 , 
    n396 , 
    n397 , 
    n398 , 
    n399 , 
    n400 , 
    n401 , 
    n402 , 
    n403 , 
    n404 , 
    n405 , 
    n406 , 
    n407 , 
    n408 , 
    n409 , 
    n410 , 
    n411 , 
    n412 , 
    n413 , 
    n414 , 
    n415 , 
    n416 , 
    n417 , 
    n418 , 
    n419 , 
    n420 , 
    n421 , 
    n422 , 
    n423 , 
    n424 , 
    n425 , 
    n426 , 
    n427 , 
    n428 , 
    n429 , 
    n430 , 
    n431 , 
    n432 , 
    n433 , 
    n434 , 
    n435 , 
    n436 , 
    n437 , 
    n438 , 
    n439 , 
    n440 , 
    n441 , 
    n442 , 
    n443 , 
    n444 , 
    n445 , 
    n446 , 
    n447 , 
    n448 , 
    n449 , 
    n450 , 
    n451 , 
    n452 , 
    n453 , 
    n454 , 
    n455 , 
    n456 , 
    n457 , 
    n458 , 
    n459 , 
    n460 , 
    n461 , 
    n462 , 
    n463 , 
    n464 , 
    n465 , 
    n466 , 
    n467 , 
    n468 , 
    n469 , 
    n470 , 
    n471 , 
    n472 , 
    n473 , 
    n474 , 
    n475 , 
    n476 , 
    n477 , 
    n478 , 
    n479 , 
    n480 , 
    n481 , 
    n482 , 
    n483 , 
    n484 , 
    n485 , 
    n486 , 
    n487 , 
    n488 , 
    n489 , 
    n490 , 
    n491 , 
    n492 , 
    n493 , 
    n494 , 
    n495 , 
    n496 , 
    n497 , 
    n498 , 
    n499 , 
    n500 , 
    n501 , 
    n502 , 
    n503 , 
    n504 , 
    n505 , 
    n506 , 
    n507 , 
    n508 , 
    n509 , 
    n510 , 
    n511 , 
    n512 , 
    n513 , 
    n514 , 
    n515 , 
    n516 , 
    n517 , 
    n518 , 
    n519 , 
    n520 , 
    n521 , 
    n522 , 
    n523 , 
    n524 , 
    n525 , 
    n526 , 
    n527 , 
    n528 , 
    n529 , 
    n530 , 
    n531 , 
    n532 , 
    n533 , 
    n534 , 
    n535 , 
    n536 , 
    n537 , 
    n538 , 
    n539 , 
    n540 , 
    n541 , 
    n542 , 
    n543 , 
    n544 , 
    n545 , 
    n546 , 
    n547 , 
    n548 , 
    n549 , 
    n550 , 
    n551 , 
    n552 , 
    n553 , 
    n554 , 
    n555 , 
    n556 , 
    n557 , 
    n558 , 
    n559 , 
    n560 , 
    n561 , 
    n562 , 
    n563 , 
    n564 , 
    n565 , 
    n566 , 
    n567 , 
    n568 , 
    n569 , 
    n570 , 
    n571 , 
    n572 , 
    n573 , 
    n574 , 
    n575 , 
    n576 , 
    n577 , 
    n578 , 
    n579 , 
    n580 , 
    n581 , 
    n582 , 
    n583 , 
    n584 , 
    n585 , 
    n586 , 
    n587 , 
    n588 , 
    n589 , 
    n590 , 
    n591 , 
    n592 , 
    n593 , 
    n594 , 
    n595 , 
    n596 , 
    n597 , 
    n598 , 
    n599 , 
    n600 , 
    n601 , 
    n602 , 
    n603 , 
    n604 , 
    n605 , 
    n606 , 
    n607 , 
    n608 , 
    n609 , 
    n610 , 
    n611 , 
    n612 , 
    n613 , 
    n614 , 
    n615 , 
    n616 , 
    n617 , 
    n618 , 
    n619 , 
    n620 , 
    n621 , 
    n622 , 
    n623 , 
    n624 , 
    n625 , 
    n626 , 
    n627 , 
    n628 , 
    n629 , 
    n630 , 
    n631 , 
    n632 , 
    n633 , 
    n634 , 
    n635 , 
    n636 , 
    n637 , 
    n638 , 
    n639 , 
    n640 , 
    n641 , 
    n642 , 
    n643 , 
    n644 , 
    n645 , 
    n646 , 
    n647 , 
    n648 , 
    n649 , 
    n650 , 
    n651 , 
    n652 , 
    n653 , 
    n654 , 
    n655 , 
    n656 , 
    n657 , 
    n658 , 
    n659 , 
    n660 , 
    n661 , 
    n662 , 
    n663 , 
    n664 , 
    n665 , 
    n666 , 
    n667 , 
    n668 , 
    n669 , 
    n670 , 
    n671 , 
    n672 , 
    n673 , 
    n674 , 
    n675 , 
    n676 , 
    n677 , 
    n678 , 
    n679 , 
    n680 , 
    n681 , 
    n682 , 
    n683 , 
    n684 , 
    n685 , 
    n686 , 
    n687 , 
    n688 , 
    n689 , 
    n690 , 
    n691 , 
    n692 , 
    n693 , 
    n694 , 
    n695 , 
    n696 , 
    n697 , 
    n698 , 
    n699 , 
    n700 , 
    n701 , 
    n702 , 
    n703 , 
    n704 , 
    n705 , 
    n706 , 
    n707 , 
    n708 , 
    n709 , 
    n710 , 
    n711 , 
    n712 , 
    n713 , 
    n714 , 
    n715 , 
    n716 , 
    n717 , 
    n718 , 
    n719 , 
    n720 , 
    n721 , 
    n722 , 
    n723 , 
    n724 , 
    n725 , 
    n726 , 
    n727 , 
    n728 , 
    n729 , 
    n730 , 
    n731 , 
    n732 , 
    n733 , 
    n734 , 
    n735 , 
    n736 , 
    n737 , 
    n738 , 
    n739 , 
    n740 , 
    n741 , 
    n742 , 
    n743 , 
    n744 , 
    n745 , 
    n746 , 
    n747 , 
    n748 , 
    n749 , 
    n750 , 
    n751 , 
    n752 , 
    n753 , 
    n754 , 
    n755 , 
    n756 , 
    n757 , 
    n758 , 
    n759 , 
    n760 , 
    n761 , 
    n762 , 
    n763 , 
    n764 , 
    n765 , 
    n766 , 
    n767 , 
    n768 , 
    n769 , 
    n770 , 
    n771 , 
    n772 , 
    n773 , 
    n774 , 
    n775 , 
    n776 , 
    n777 , 
    n778 , 
    n779 , 
    n780 , 
    n781 , 
    n782 , 
    n783 , 
    n784 , 
    n785 , 
    n786 , 
    n787 , 
    n788 , 
    n789 , 
    n790 , 
    n791 , 
    n792 , 
    n793 , 
    n794 , 
    n795 , 
    n796 , 
    n797 , 
    n798 , 
    n799 , 
    n800 , 
    n801 , 
    n802 , 
    n803 , 
    n804 , 
    n805 , 
    n806 , 
    n807 , 
    n808 , 
    n809 , 
    n810 , 
    n811 , 
    n812 , 
    n813 , 
    n814 , 
    n815 , 
    n816 , 
    n817 , 
    n818 , 
    n819 , 
    n820 , 
    n821 , 
    n822 , 
    n823 , 
    n824 , 
    n825 , 
    n826 , 
    n827 , 
    n828 , 
    n829 , 
    n830 , 
    n831 , 
    n832 , 
    n833 , 
    n834 , 
    n835 , 
    n836 , 
    n837 , 
    n838 , 
    n839 , 
    n840 , 
    n841 , 
    n842 , 
    n843 , 
    n844 , 
    n845 , 
    n846 , 
    n847 , 
    n848 , 
    n849 , 
    n850 , 
    n851 , 
    n852 , 
    n853 , 
    n854 , 
    n855 , 
    n856 , 
    n857 , 
    n858 , 
    n859 , 
    n860 , 
    n861 , 
    n862 , 
    n863 , 
    n864 , 
    n865 , 
    n866 , 
    n867 , 
    n868 , 
    n869 , 
    n870 , 
    n871 , 
    n872 , 
    n873 , 
    n874 , 
    n875 , 
    n876 , 
    n877 , 
    n878 , 
    n879 , 
    n880 , 
    n881 , 
    n882 , 
    n883 , 
    n884 , 
    n885 , 
    n886 , 
    n887 , 
    n888 , 
    n889 , 
    n890 , 
    n891 , 
    n892 , 
    n893 , 
    n894 , 
    n895 , 
    n896 , 
    n897 , 
    n898 , 
    n899 , 
    n900 , 
    n901 , 
    n902 , 
    n903 , 
    n904 , 
    n905 , 
    n906 , 
    n907 , 
    n908 , 
    n909 , 
    n910 , 
    n911 , 
    n912 , 
    n913 , 
    n914 , 
    n915 , 
    n916 , 
    n917 , 
    n918 , 
    n919 , 
    n920 , 
    n921 , 
    n922 , 
    n923 , 
    n924 , 
    n925 , 
    n926 , 
    n927 , 
    n928 , 
    n929 , 
    n930 , 
    n931 , 
    n932 , 
    n933 , 
    n934 , 
    n935 , 
    n936 , 
    n937 , 
    n938 , 
    n939 , 
    n940 , 
    n941 , 
    n942 , 
    n943 , 
    n944 , 
    n945 , 
    n946 , 
    n947 , 
    n948 , 
    n949 , 
    n950 , 
    n951 , 
    n952 , 
    n953 , 
    n954 , 
    n955 , 
    n956 , 
    n957 , 
    n958 , 
    n959 , 
    n960 , 
    n961 , 
    n962 , 
    n963 , 
    n964 , 
    n965 , 
    n966 , 
    n967 , 
    n968 , 
    n969 , 
    n970 , 
    n971 , 
    n972 , 
    n973 , 
    n974 , 
    n975 , 
    n976 , 
    n977 , 
    n978 , 
    n979 , 
    n980 , 
    n981 , 
    n982 , 
    n983 , 
    n984 , 
    n985 , 
    n986 , 
    n987 , 
    n988 , 
    n989 , 
    n990 , 
    n991 , 
    n992 , 
    n993 , 
    n994 , 
    n995 , 
    n996 , 
    n997 , 
    n998 , 
    n999 , 
    n1000 , 
    n1001 , 
    n1002 , 
    n1003 , 
    n1004 , 
    n1005 , 
    n1006 , 
    n1007 , 
    n1008 , 
    n1009 , 
    n1010 , 
    n1011 , 
    n1012 , 
    n1013 , 
    n1014 , 
    n1015 , 
    n1016 , 
    n1017 , 
    n1018 , 
    n1019 , 
    n1020 , 
    n1021 , 
    n1022 , 
    n1023 , 
    n1024 , 
    n1025 , 
    n1026 , 
    n1027 , 
    n1028 , 
    n1029 , 
    n1030 , 
    n1031 , 
    n1032 , 
    n1033 , 
    n1034 , 
    n1035 , 
    n1036 , 
    n1037 , 
    n1038 , 
    n1039 , 
    n1040 , 
    n1041 , 
    n1042 , 
    n1043 , 
    n1044 , 
    n1045 , 
    n1046 , 
    n1047 , 
    n1048 , 
    n1049 , 
    n1050 , 
    n1051 , 
    n1052 , 
    n1053 , 
    n1054 , 
    n1055 , 
    n1056 , 
    n1057 , 
    n1058 , 
    n1059 , 
    n1060 , 
    n1061 , 
    n1062 , 
    n1063 , 
    n1064 , 
    n1065 , 
    n1066 , 
    n1067 , 
    n1068 , 
    n1069 , 
    n1070 , 
    n1071 , 
    n1072 , 
    n1073 , 
    n1074 , 
    n1075 , 
    n1076 , 
    n1077 , 
    n1078 , 
    n1079 , 
    n1080 , 
    n1081 , 
    n1082 , 
    n1083 , 
    n1084 , 
    n1085 , 
    n1086 , 
    n1087 , 
    n1088 , 
    n1089 , 
    n1090 , 
    n1091 , 
    n1092 , 
    n1093 , 
    n1094 , 
    n1095 , 
    n1096 , 
    n1097 , 
    n1098 , 
    n1099 , 
    n1100 , 
    n1101 , 
    n1102 , 
    n1103 , 
    n1104 , 
    n1105 , 
    n1106 , 
    n1107 , 
    n1108 , 
    n1109 , 
    n1110 , 
    n1111 , 
    n1112 , 
    n1113 , 
    n1114 , 
    n1115 , 
    n1116 , 
    n1117 , 
    n1118 , 
    n1119 , 
    n1120 , 
    n1121 , 
    n1122 , 
    n1123 , 
    n1124 , 
    n1125 , 
    n1126 , 
    n1127 , 
    n1128 , 
    n1129 , 
    n1130 , 
    n1131 , 
    n1132 , 
    n1133 , 
    n1134 , 
    n1135 , 
    n1136 , 
    n1137 , 
    n1138 , 
    n1139 , 
    n1140 , 
    n1141 , 
    n1142 , 
    n1143 , 
    n1144 , 
    n1145 , 
    n1146 , 
    n1147 , 
    n1148 , 
    n1149 , 
    n1150 , 
    n1151 , 
    n1152 , 
    n1153 , 
    n1154 , 
    n1155 , 
    n1156 , 
    n1157 , 
    n1158 , 
    n1159 , 
    n1160 , 
    n1161 , 
    n1162 , 
    n1163 , 
    n1164 , 
    n1165 , 
    n1166 , 
    n1167 , 
    n1168 , 
    n1169 , 
    n1170 , 
    n1171 , 
    n1172 , 
    n1173 , 
    n1174 , 
    n1175 , 
    n1176 , 
    n1177 , 
    n1178 , 
    n1179 , 
    n1180 , 
    n1181 , 
    n1182 , 
    n1183 , 
    n1184 , 
    n1185 , 
    n1186 , 
    n1187 , 
    n1188 , 
    n1189 , 
    n1190 , 
    n1191 , 
    n1192 , 
    n1193 , 
    n1194 , 
    n1195 , 
    n1196 , 
    n1197 , 
    n1198 , 
    n1199 , 
    n1200 , 
    n1201 , 
    n1202 , 
    n1203 , 
    n1204 , 
    n1205 , 
    n1206 , 
    n1207 , 
    n1208 , 
    n1209 , 
    n1210 , 
    n1211 , 
    n1212 , 
    n1213 , 
    n1214 , 
    n1215 , 
    n1216 , 
    n1217 , 
    n1218 , 
    n1219 , 
    n1220 , 
    n1221 , 
    n1222 , 
    n1223 , 
    n1224 , 
    n1225 , 
    n1226 , 
    n1227 , 
    n1228 , 
    n1229 , 
    n1230 , 
    n1231 , 
    n1232 , 
    n1233 , 
    n1234 , 
    n1235 , 
    n1236 , 
    n1237 , 
    n1238 , 
    n1239 , 
    n1240 , 
    n1241 , 
    n1242 , 
    n1243 , 
    n1244 , 
    n1245 , 
    n1246 , 
    n1247 , 
    n1248 , 
    n1249 , 
    n1250 , 
    n1251 , 
    n1252 , 
    n1253 , 
    n1254 , 
    n1255 , 
    n1256 , 
    n1257 , 
    n1258 , 
    n1259 , 
    n1260 , 
    n1261 , 
    n1262 , 
    n1263 , 
    n1264 , 
    n1265 , 
    n1266 , 
    n1267 , 
    n1268 , 
    n1269 , 
    n1270 , 
    n1271 , 
    n1272 , 
    n1273 , 
    n1274 , 
    n1275 , 
    n1276 , 
    n1277 , 
    n1278 , 
    n1279 , 
    n1280 , 
    n1281 , 
    n1282 , 
    n1283 , 
    n1284 , 
    n1285 , 
    n1286 , 
    n1287 , 
    n1288 , 
    n1289 , 
    n1290 , 
    n1291 , 
    n1292 , 
    n1293 , 
    n1294 , 
    n1295 , 
    n1296 , 
    n1297 , 
    n1298 , 
    n1299 , 
    n1300 , 
    n1301 , 
    n1302 , 
    n1303 , 
    n1304 , 
    n1305 , 
    n1306 , 
    n1307 , 
    n1308 , 
    n1309 , 
    n1310 , 
    n1311 , 
    n1312 , 
    n1313 , 
    n1314 , 
    n1315 , 
    n1316 , 
    n1317 , 
    n1318 , 
    n1319 , 
    n1320 , 
    n1321 , 
    n1322 , 
    n1323 , 
    n1324 , 
    n1325 , 
    n1326 , 
    n1327 , 
    n1328 , 
    n1329 , 
    n1330 , 
    n1331 , 
    n1332 , 
    n1333 , 
    n1334 , 
    n1335 , 
    n1336 , 
    n1337 , 
    n1338 , 
    n1339 , 
    n1340 , 
    n1341 , 
    n1342 , 
    n1343 , 
    n1344 , 
    n1345 , 
    n1346 , 
    n1347 , 
    n1348 , 
    n1349 , 
    n1350 , 
    n1351 , 
    n1352 , 
    n1353 , 
    n1354 , 
    n1355 , 
    n1356 , 
    n1357 , 
    n1358 , 
    n1359 , 
    n1360 , 
    n1361 , 
    n1362 , 
    n1363 , 
    n1364 , 
    n1365 , 
    n1366 , 
    n1367 , 
    n1368 , 
    n1369 , 
    n1370 , 
    n1371 , 
    n1372 , 
    n1373 , 
    n1374 , 
    n1375 , 
    n1376 , 
    n1377 , 
    n1378 , 
    n1379 , 
    n1380 , 
    n1381 , 
    n1382 , 
    n1383 , 
    n1384 , 
    n1385 , 
    n1386 , 
    n1387 , 
    n1388 , 
    n1389 , 
    n1390 , 
    n1391 , 
    n1392 , 
    n1393 , 
    n1394 , 
    n1395 , 
    n1396 , 
    n1397 , 
    n1398 , 
    n1399 , 
    n1400 , 
    n1401 , 
    n1402 , 
    n1403 , 
    n1404 , 
    n1405 , 
    n1406 , 
    n1407 , 
    n1408 , 
    n1409 , 
    n1410 , 
    n1411 , 
    n1412 , 
    n1413 , 
    n1414 , 
    n1415 , 
    n1416 , 
    n1417 , 
    n1418 , 
    n1419 , 
    n1420 , 
    n1421 , 
    n1422 , 
    n1423 , 
    n1424 , 
    n1425 , 
    n1426 , 
    n1427 , 
    n1428 , 
    n1429 , 
    n1430 , 
    n1431 , 
    n1432 , 
    n1433 , 
    n1434 , 
    n1435 , 
    n1436 , 
    n1437 , 
    n1438 , 
    n1439 , 
    n1440 , 
    n1441 , 
    n1442 , 
    n1443 , 
    n1444 , 
    n1445 , 
    n1446 , 
    n1447 , 
    n1448 , 
    n1449 , 
    n1450 , 
    n1451 , 
    n1452 , 
    n1453 , 
    n1454 , 
    n1455 , 
    n1456 , 
    n1457 , 
    n1458 , 
    n1459 , 
    n1460 , 
    n1461 , 
    n1462 , 
    n1463 , 
    n1464 , 
    n1465 , 
    n1466 , 
    n1467 , 
    n1468 , 
    n1469 , 
    n1470 , 
    n1471 , 
    n1472 , 
    n1473 , 
    n1474 , 
    n1475 , 
    n1476 , 
    n1477 , 
    n1478 , 
    n1479 , 
    n1480 , 
    n1481 , 
    n1482 , 
    n1483 , 
    n1484 , 
    n1485 , 
    n1486 , 
    n1487 , 
    n1488 , 
    n1489 , 
    n1490 , 
    n1491 , 
    n1492 , 
    n1493 , 
    n1494 , 
    n1495 , 
    n1496 , 
    n1497 , 
    n1498 , 
    n1499 , 
    n1500 , 
    n1501 , 
    n1502 , 
    n1503 , 
    n1504 , 
    n1505 , 
    n1506 , 
    n1507 , 
    n1508 , 
    n1509 , 
    n1510 , 
    n1511 , 
    n1512 , 
    n1513 , 
    n1514 , 
    n1515 , 
    n1516 , 
    n1517 , 
    n1518 , 
    n1519 , 
    n1520 , 
    n1521 , 
    n1522 , 
    n1523 , 
    n1524 , 
    n1525 , 
    n1526 , 
    n1527 , 
    n1528 , 
    n1529 , 
    n1530 , 
    n1531 , 
    n1532 , 
    n1533 , 
    n1534 , 
    n1535 , 
    n1536 , 
    n1537 , 
    n1538 , 
    n1539 , 
    n1540 , 
    n1541 , 
    n1542 , 
    n1543 , 
    n1544 , 
    n1545 , 
    n1546 , 
    n1547 , 
    n1548 , 
    n1549 , 
    n1550 , 
    n1551 , 
    n1552 , 
    n1553 , 
    n1554 , 
    n1555 , 
    n1556 , 
    n1557 , 
    n1558 , 
    n1559 , 
    n1560 , 
    n1561 , 
    n1562 , 
    n1563 , 
    n1564 , 
    n1565 , 
    n1566 , 
    n1567 , 
    n1568 , 
    n1569 , 
    n1570 , 
    n1571 , 
    n1572 , 
    n1573 , 
    n1574 , 
    n1575 , 
    n1576 , 
    n1577 , 
    n1578 , 
    n1579 , 
    n1580 , 
    n1581 , 
    n1582 , 
    n1583 , 
    n1584 , 
    n1585 , 
    n1586 , 
    n1587 , 
    n1588 , 
    n1589 , 
    n1590 , 
    n1591 , 
    n1592 , 
    n1593 , 
    n1594 , 
    n1595 , 
    n1596 , 
    n1597 , 
    n1598 , 
    n1599 , 
    n1600 , 
    n1601 , 
    n1602 , 
    n1603 , 
    n1604 , 
    n1605 , 
    n1606 , 
    n1607 , 
    n1608 , 
    n1609 , 
    n1610 , 
    n1611 , 
    n1612 , 
    n1613 , 
    n1614 , 
    n1615 , 
    n1616 , 
    n1617 , 
    n1618 , 
    n1619 , 
    n1620 , 
    n1621 , 
    n1622 , 
    n1623 , 
    n1624 , 
    n1625 , 
    n1626 , 
    n1627 , 
    n1628 , 
    n1629 , 
    n1630 , 
    n1631 , 
    n1632 , 
    n1633 , 
    n1634 , 
    n1635 , 
    n1636 , 
    n1637 , 
    n1638 , 
    n1639 , 
    n1640 , 
    n1641 , 
    n1642 , 
    n1643 , 
    n1644 , 
    n1645 , 
    n1646 , 
    n1647 , 
    n1648 , 
    n1649 , 
    n1650 , 
    n1651 , 
    n1652 , 
    n1653 , 
    n1654 , 
    n1655 , 
    n1656 , 
    n1657 , 
    n1658 , 
    n1659 , 
    n1660 , 
    n1661 , 
    n1662 , 
    n1663 , 
    n1664 , 
    n1665 , 
    n1666 , 
    n1667 , 
    n1668 , 
    n1669 , 
    n1670 , 
    n1671 , 
    n1672 , 
    n1673 , 
    n1674 , 
    n1675 , 
    n1676 , 
    n1677 , 
    n1678 , 
    n1679 , 
    n1680 , 
    n1681 , 
    n1682 , 
    n1683 , 
    n1684 , 
    n1685 , 
    n1686 , 
    n1687 , 
    n1688 , 
    n1689 , 
    n1690 , 
    n1691 , 
    n1692 , 
    n1693 , 
    n1694 , 
    n1695 , 
    n1696 , 
    n1697 , 
    n1698 , 
    n1699 , 
    n1700 , 
    n1701 , 
    n1702 , 
    n1703 , 
    n1704 , 
    n1705 , 
    n1706 , 
    n1707 , 
    n1708 , 
    n1709 , 
    n1710 , 
    n1711 , 
    n1712 , 
    n1713 , 
    n1714 , 
    n1715 , 
    n1716 , 
    n1717 , 
    n1718 , 
    n1719 , 
    n1720 , 
    n1721 , 
    n1722 , 
    n1723 , 
    n1724 , 
    n1725 , 
    n1726 , 
    n1727 , 
    n1728 , 
    n1729 , 
    n1730 , 
    n1731 , 
    n1732 , 
    n1733 , 
    n1734 , 
    n1735 , 
    n1736 , 
    n1737 , 
    n1738 , 
    n1739 , 
    n1740 , 
    n1741 , 
    n1742 , 
    n1743 , 
    n1744 , 
    n1745 , 
    n1746 , 
    n1747 , 
    n1748 , 
    n1749 , 
    n1750 , 
    n1751 , 
    n1752 , 
    n1753 , 
    n1754 , 
    n1755 , 
    n1756 , 
    n1757 , 
    n1758 , 
    n1759 , 
    n1760 , 
    n1761 , 
    n1762 , 
    n1763 , 
    n1764 , 
    n1765 , 
    n1766 , 
    n1767 , 
    n1768 , 
    n1769 , 
    n1770 , 
    n1771 , 
    n1772 , 
    n1773 , 
    n1774 , 
    n1775 , 
    n1776 , 
    n1777 , 
    n1778 , 
    n1779 , 
    n1780 , 
    n1781 , 
    n1782 , 
    n1783 , 
    n1784 , 
    n1785 , 
    n1786 , 
    n1787 , 
    n1788 , 
    n1789 , 
    n1790 , 
    n1791 , 
    n1792 , 
    n1793 , 
    n1794 , 
    n1795 , 
    n1796 , 
    n1797 , 
    n1798 , 
    n1799 , 
    n1800 , 
    n1801 , 
    n1802 , 
    n1803 , 
    n1804 , 
    n1805 , 
    n1806 , 
    n1807 , 
    n1808 , 
    n1809 , 
    n1810 , 
    n1811 , 
    n1812 , 
    n1813 , 
    n1814 , 
    n1815 , 
    n1816 , 
    n1817 , 
    n1818 , 
    n1819 , 
    n1820 , 
    n1821 , 
    n1822 , 
    n1823 , 
    n1824 , 
    n1825 , 
    n1826 , 
    n1827 , 
    n1828 , 
    n1829 , 
    n1830 , 
    n1831 , 
    n1832 , 
    n1833 , 
    n1834 , 
    n1835 , 
    n1836 , 
    n1837 , 
    n1838 , 
    n1839 , 
    n1840 , 
    n1841 , 
    n1842 , 
    n1843 , 
    n1844 , 
    n1845 , 
    n1846 , 
    n1847 , 
    n1848 , 
    n1849 , 
    n1850 , 
    n1851 , 
    n1852 , 
    n1853 , 
    n1854 , 
    n1855 , 
    n1856 , 
    n1857 , 
    n1858 , 
    n1859 , 
    n1860 , 
    n1861 , 
    n1862 , 
    n1863 , 
    n1864 , 
    n1865 , 
    n1866 , 
    n1867 , 
    n1868 , 
    n1869 , 
    n1870 , 
    n1871 , 
    n1872 , 
    n1873 , 
    n1874 , 
    n1875 , 
    n1876 , 
    n1877 , 
    n1878 , 
    n1879 , 
    n1880 , 
    n1881 , 
    n1882 , 
    n1883 , 
    n1884 , 
    n1885 , 
    n1886 , 
    n1887 , 
    n1888 , 
    n1889 , 
    n1890 , 
    n1891 , 
    n1892 , 
    n1893 , 
    n1894 , 
    n1895 , 
    n1896 , 
    n1897 , 
    n1898 , 
    n1899 , 
    n1900 , 
    n1901 , 
    n1902 , 
    n1903 , 
    n1904 , 
    n1905 , 
    n1906 , 
    n1907 , 
    n1908 , 
    n1909 , 
    n1910 , 
    n1911 , 
    n1912 , 
    n1913 , 
    n1914 , 
    n1915 , 
    n1916 , 
    n1917 , 
    n1918 , 
    n1919 , 
    n1920 , 
    n1921 , 
    n1922 , 
    n1923 , 
    n1924 , 
    n1925 , 
    n1926 , 
    n1927 , 
    n1928 , 
    n1929 , 
    n1930 , 
    n1931 , 
    n1932 , 
    n1933 , 
    n1934 , 
    n1935 , 
    n1936 , 
    n1937 , 
    n1938 , 
    n1939 , 
    n1940 , 
    n1941 , 
    n1942 , 
    n1943 , 
    n1944 , 
    n1945 , 
    n1946 , 
    n1947 , 
    n1948 , 
    n1949 , 
    n1950 , 
    n1951 , 
    n1952 , 
    n1953 , 
    n1954 , 
    n1955 , 
    n1956 , 
    n1957 , 
    n1958 , 
    n1959 , 
    n1960 , 
    n1961 , 
    n1962 , 
    n1963 , 
    n1964 , 
    n1965 , 
    n1966 , 
    n1967 , 
    n1968 , 
    n1969 , 
    n1970 , 
    n1971 , 
    n1972 , 
    n1973 , 
    n1974 , 
    n1975 , 
    n1976 , 
    n1977 , 
    n1978 , 
    n1979 , 
    n1980 , 
    n1981 , 
    n1982 , 
    n1983 , 
    n1984 , 
    n1985 , 
    n1986 , 
    n1987 , 
    n1988 , 
    n1989 , 
    n1990 , 
    n1991 , 
    n1992 , 
    n1993 , 
    n1994 , 
    n1995 , 
    n1996 , 
    n1997 , 
    n1998 , 
    n1999 , 
    n2000 , 
    n2001 , 
    n2002 , 
    n2003 , 
    n2004 , 
    n2005 , 
    n2006 , 
    n2007 , 
    n2008 , 
    n2009 , 
    n2010 , 
    n2011 , 
    n2012 , 
    n2013 , 
    n2014 , 
    n2015 , 
    n2016 , 
    n2017 , 
    n2018 , 
    n2019 , 
    n2020 , 
    n2021 , 
    n2022 , 
    n2023 , 
    n2024 , 
    n2025 , 
    n2026 , 
    n2027 , 
    n2028 , 
    n2029 , 
    n2030 , 
    n2031 , 
    n2032 , 
    n2033 , 
    n2034 , 
    n2035 , 
    n2036 , 
    n2037 , 
    n2038 , 
    n2039 , 
    n2040 , 
    n2041 , 
    n2042 , 
    n2043 , 
    n2044 , 
    n2045 , 
    n2046 , 
    n2047 , 
    n2048 , 
    n2049 , 
    n2050 , 
    n2051 , 
    n2052 , 
    n2053 , 
    n2054 , 
    n2055 , 
    n2056 , 
    n2057 , 
    n2058 , 
    n2059 , 
    n2060 , 
    n2061 , 
    n2062 , 
    n2063 , 
    n2064 , 
    n2065 , 
    n2066 , 
    n2067 , 
    n2068 , 
    n2069 , 
    n2070 , 
    n2071 , 
    n2072 , 
    n2073 , 
    n2074 , 
    n2075 , 
    n2076 , 
    n2077 , 
    n2078 , 
    n2079 , 
    n2080 , 
    n2081 , 
    n2082 , 
    n2083 , 
    n2084 , 
    n2085 , 
    n2086 , 
    n2087 , 
    n2088 , 
    n2089 , 
    n2090 , 
    n2091 , 
    n2092 , 
    n2093 , 
    n2094 , 
    n2095 , 
    n2096 , 
    n2097 , 
    n2098 , 
    n2099 , 
    n2100 , 
    n2101 , 
    n2102 , 
    n2103 , 
    n2104 , 
    n2105 , 
    n2106 , 
    n2107 , 
    n2108 , 
    n2109 , 
    n2110 , 
    n2111 , 
    n2112 , 
    n2113 , 
    n2114 , 
    n2115 , 
    n2116 , 
    n2117 , 
    n2118 , 
    n2119 , 
    n2120 , 
    n2121 , 
    n2122 , 
    n2123 , 
    n2124 , 
    n2125 , 
    n2126 , 
    n2127 , 
    n2128 , 
    n2129 , 
    n2130 , 
    n2131 , 
    n2132 , 
    n2133 , 
    n2134 , 
    n2135 , 
    n2136 , 
    n2137 , 
    n2138 , 
    n2139 , 
    n2140 , 
    n2141 , 
    n2142 , 
    n2143 , 
    n2144 , 
    n2145 , 
    n2146 , 
    n2147 , 
    n2148 , 
    n2149 , 
    n2150 , 
    n2151 , 
    n2152 , 
    n2153 , 
    n2154 , 
    n2155 , 
    n2156 , 
    n2157 , 
    n2158 , 
    n2159 , 
    n2160 , 
    n2161 , 
    n2162 , 
    n2163 , 
    n2164 , 
    n2165 , 
    n2166 , 
    n2167 , 
    n2168 , 
    n2169 , 
    n2170 , 
    n2171 , 
    n2172 , 
    n2173 , 
    n2174 , 
    n2175 , 
    n2176 , 
    n2177 , 
    n2178 , 
    n2179 , 
    n2180 , 
    n2181 , 
    n2182 , 
    n2183 , 
    n2184 , 
    n2185 , 
    n2186 , 
    n2187 , 
    n2188 , 
    n2189 , 
    n2190 , 
    n2191 , 
    n2192 , 
    n2193 , 
    n2194 , 
    n2195 , 
    n2196 , 
    n2197 , 
    n2198 , 
    n2199 , 
    n2200 , 
    n2201 , 
    n2202 , 
    n2203 , 
    n2204 , 
    n2205 , 
    n2206 , 
    n2207 , 
    n2208 , 
    n2209 , 
    n2210 , 
    n2211 , 
    n2212 , 
    n2213 , 
    n2214 , 
    n2215 , 
    n2216 , 
    n2217 , 
    n2218 , 
    n2219 , 
    n2220 , 
    n2221 , 
    n2222 , 
    n2223 , 
    n2224 , 
    n2225 , 
    n2226 , 
    n2227 , 
    n2228 , 
    n2229 , 
    n2230 , 
    n2231 , 
    n2232 , 
    n2233 , 
    n2234 , 
    n2235 , 
    n2236 , 
    n2237 , 
    n2238 , 
    n2239 , 
    n2240 , 
    n2241 , 
    n2242 , 
    n2243 , 
    n2244 , 
    n2245 , 
    n2246 , 
    n2247 , 
    n2248 , 
    n2249 , 
    n2250 , 
    n2251 , 
    n2252 , 
    n2253 , 
    n2254 , 
    n2255 , 
    n2256 , 
    n2257 , 
    n2258 , 
    n2259 , 
    n2260 , 
    n2261 , 
    n2262 , 
    n2263 , 
    n2264 , 
    n2265 , 
    n2266 , 
    n2267 , 
    n2268 , 
    n2269 , 
    n2270 , 
    n2271 , 
    n2272 , 
    n2273 , 
    n2274 , 
    n2275 , 
    n2276 , 
    n2277 , 
    n2278 , 
    n2279 , 
    n2280 , 
    n2281 , 
    n2282 , 
    n2283 , 
    n2284 , 
    n2285 , 
    n2286 , 
    n2287 , 
    n2288 , 
    n2289 , 
    n2290 , 
    n2291 , 
    n2292 , 
    n2293 , 
    n2294 , 
    n2295 , 
    n2296 , 
    n2297 , 
    n2298 , 
    n2299 , 
    n2300 , 
    n2301 , 
    n2302 , 
    n2303 , 
    n2304 , 
    n2305 , 
    n2306 , 
    n2307 , 
    n2308 , 
    n2309 , 
    n2310 , 
    n2311 , 
    n2312 , 
    n2313 , 
    n2314 , 
    n2315 , 
    n2316 , 
    n2317 , 
    n2318 , 
    n2319 , 
    n2320 , 
    n2321 , 
    n2322 , 
    n2323 , 
    n2324 , 
    n2325 , 
    n2326 , 
    n2327 , 
    n2328 , 
    n2329 , 
    n2330 , 
    n2331 , 
    n2332 , 
    n2333 , 
    n2334 , 
    n2335 , 
    n2336 , 
    n2337 , 
    n2338 , 
    n2339 , 
    n2340 , 
    n2341 , 
    n2342 , 
    n2343 , 
    n2344 , 
    n2345 , 
    n2346 , 
    n2347 , 
    n2348 , 
    n2349 , 
    n2350 , 
    n2351 , 
    n2352 , 
    n2353 , 
    n2354 , 
    n2355 , 
    n2356 , 
    n2357 , 
    n2358 , 
    n2359 , 
    n2360 , 
    n2361 , 
    n2362 , 
    n2363 , 
    n2364 , 
    n2365 , 
    n2366 , 
    n2367 , 
    n2368 , 
    n2369 , 
    n2370 , 
    n2371 , 
    n2372 , 
    n2373 , 
    n2374 , 
    n2375 , 
    n2376 , 
    n2377 , 
    n2378 , 
    n2379 , 
    n2380 , 
    n2381 , 
    n2382 , 
    n2383 , 
    n2384 , 
    n2385 , 
    n2386 , 
    n2387 , 
    n2388 , 
    n2389 , 
    n2390 , 
    n2391 , 
    n2392 , 
    n2393 , 
    n2394 , 
    n2395 , 
    n2396 , 
    n2397 , 
    n2398 , 
    n2399 , 
    n2400 , 
    n2401 , 
    n2402 , 
    n2403 , 
    n2404 , 
    n2405 , 
    n2406 , 
    n2407 , 
    n2408 , 
    n2409 , 
    n2410 , 
    n2411 , 
    n2412 , 
    n2413 , 
    n2414 , 
    n2415 , 
    n2416 , 
    n2417 , 
    n2418 , 
    n2419 , 
    n2420 , 
    n2421 , 
    n2422 , 
    n2423 , 
    n2424 , 
    n2425 , 
    n2426 , 
    n2427 , 
    n2428 , 
    n2429 , 
    n2430 , 
    n2431 , 
    n2432 , 
    n2433 , 
    n2434 , 
    n2435 , 
    n2436 , 
    n2437 , 
    n2438 , 
    n2439 , 
    n2440 , 
    n2441 , 
    n2442 , 
    n2443 , 
    n2444 , 
    n2445 , 
    n2446 , 
    n2447 , 
    n2448 , 
    n2449 , 
    n2450 , 
    n2451 , 
    n2452 , 
    n2453 , 
    n2454 , 
    n2455 , 
    n2456 , 
    n2457 , 
    n2458 , 
    n2459 , 
    n2460 , 
    n2461 , 
    n2462 , 
    n2463 , 
    n2464 , 
    n2465 , 
    n2466 , 
    n2467 , 
    n2468 , 
    n2469 , 
    n2470 , 
    n2471 , 
    n2472 , 
    n2473 , 
    n2474 , 
    n2475 , 
    n2476 , 
    n2477 , 
    n2478 , 
    n2479 , 
    n2480 , 
    n2481 , 
    n2482 , 
    n2483 , 
    n2484 , 
    n2485 , 
    n2486 , 
    n2487 , 
    n2488 , 
    n2489 , 
    n2490 , 
    n2491 , 
    n2492 , 
    n2493 , 
    n2494 , 
    n2495 , 
    n2496 , 
    n2497 , 
    n2498 , 
    n2499 , 
    n2500 , 
    n2501 , 
    n2502 , 
    n2503 , 
    n2504 , 
    n2505 , 
    n2506 , 
    n2507 , 
    n2508 , 
    n2509 , 
    n2510 , 
    n2511 , 
    n2512 , 
    n2513 , 
    n2514 , 
    n2515 , 
    n2516 , 
    n2517 , 
    n2518 , 
    n2519 , 
    n2520 , 
    n2521 , 
    n2522 , 
    n2523 , 
    n2524 , 
    n2525 , 
    n2526 , 
    n2527 , 
    n2528 , 
    n2529 , 
    n2530 , 
    n2531 , 
    n2532 , 
    n2533 , 
    n2534 , 
    n2535 , 
    n2536 , 
    n2537 , 
    n2538 , 
    n2539 , 
    n2540 , 
    n2541 , 
    n2542 , 
    n2543 , 
    n2544 , 
    n2545 , 
    n2546 , 
    n2547 , 
    n2548 , 
    n2549 , 
    n2550 , 
    n2551 , 
    n2552 , 
    n2553 , 
    n2554 , 
    n2555 , 
    n2556 , 
    n2557 , 
    n2558 , 
    n2559 , 
    n2560 , 
    n2561 , 
    n2562 , 
    n2563 , 
    n2564 , 
    n2565 , 
    n2566 , 
    n2567 , 
    n2568 , 
    n2569 , 
    n2570 , 
    n2571 , 
    n2572 , 
    n2573 , 
    n2574 , 
    n2575 , 
    n2576 , 
    n2577 , 
    n2578 , 
    n2579 , 
    n2580 , 
    n2581 , 
    n2582 , 
    n2583 , 
    n2584 , 
    n2585 , 
    n2586 , 
    n2587 , 
    n2588 , 
    n2589 , 
    n2590 , 
    n2591 , 
    n2592 , 
    n2593 , 
    n2594 , 
    n2595 , 
    n2596 , 
    n2597 , 
    n2598 , 
    n2599 , 
    n2600 , 
    n2601 , 
    n2602 , 
    n2603 , 
    n2604 , 
    n2605 , 
    n2606 , 
    n2607 , 
    n2608 , 
    n2609 , 
    n2610 , 
    n2611 , 
    n2612 , 
    n2613 , 
    n2614 , 
    n2615 , 
    n2616 , 
    n2617 , 
    n2618 , 
    n2619 , 
    n2620 , 
    n2621 , 
    n2622 , 
    n2623 , 
    n2624 , 
    n2625 , 
    n2626 , 
    n2627 , 
    n2628 , 
    n2629 , 
    n2630 , 
    n2631 , 
    n2632 , 
    n2633 , 
    n2634 , 
    n2635 , 
    n2636 , 
    n2637 , 
    n2638 , 
    n2639 , 
    n2640 , 
    n2641 , 
    n2642 , 
    n2643 , 
    n2644 , 
    n2645 , 
    n2646 , 
    n2647 , 
    n2648 , 
    n2649 , 
    n2650 , 
    n2651 , 
    n2652 , 
    n2653 , 
    n2654 , 
    n2655 , 
    n2656 , 
    n2657 , 
    n2658 , 
    n2659 , 
    n2660 , 
    n2661 , 
    n2662 , 
    n2663 , 
    n2664 , 
    n2665 , 
    n2666 , 
    n2667 , 
    n2668 , 
    n2669 , 
    n2670 , 
    n2671 , 
    n2672 , 
    n2673 , 
    n2674 , 
    n2675 , 
    n2676 , 
    n2677 , 
    n2678 , 
    n2679 , 
    n2680 , 
    n2681 , 
    n2682 , 
    n2683 , 
    n2684 , 
    n2685 , 
    n2686 , 
    n2687 , 
    n2688 , 
    n2689 , 
    n2690 , 
    n2691 , 
    n2692 , 
    n2693 , 
    n2694 , 
    n2695 , 
    n2696 , 
    n2697 , 
    n2698 , 
    n2699 , 
    n2700 , 
    n2701 , 
    n2702 , 
    n2703 , 
    n2704 , 
    n2705 , 
    n2706 , 
    n2707 , 
    n2708 , 
    n2709 , 
    n2710 , 
    n2711 , 
    n2712 , 
    n2713 , 
    n2714 , 
    n2715 , 
    n2716 , 
    n2717 , 
    n2718 , 
    n2719 , 
    n2720 , 
    n2721 , 
    n2722 , 
    n2723 , 
    n2724 , 
    n2725 , 
    n2726 , 
    n2727 , 
    n2728 , 
    n2729 , 
    n2730 , 
    n2731 , 
    n2732 , 
    n2733 , 
    n2734 , 
    n2735 , 
    n2736 , 
    n2737 , 
    n2738 , 
    n2739 , 
    n2740 , 
    n2741 , 
    n2742 , 
    n2743 , 
    n2744 , 
    n2745 , 
    n2746 , 
    n2747 , 
    n2748 , 
    n2749 , 
    n2750 , 
    n2751 , 
    n2752 , 
    n2753 , 
    n2754 , 
    n2755 , 
    n2756 , 
    n2757 , 
    n2758 , 
    n2759 , 
    n2760 , 
    n2761 , 
    n2762 , 
    n2763 , 
    n2764 , 
    n2765 , 
    n2766 , 
    n2767 , 
    n2768 , 
    n2769 , 
    n2770 , 
    n2771 , 
    n2772 , 
    n2773 , 
    n2774 , 
    n2775 , 
    n2776 , 
    n2777 , 
    n2778 , 
    n2779 , 
    n2780 , 
    n2781 , 
    n2782 , 
    n2783 , 
    n2784 , 
    n2785 , 
    n2786 , 
    n2787 , 
    n2788 , 
    n2789 , 
    n2790 , 
    n2791 , 
    n2792 , 
    n2793 , 
    n2794 , 
    n2795 , 
    n2796 , 
    n2797 , 
    n2798 , 
    n2799 , 
    n2800 , 
    n2801 , 
    n2802 , 
    n2803 , 
    n2804 , 
    n2805 , 
    n2806 , 
    n2807 , 
    n2808 , 
    n2809 , 
    n2810 , 
    n2811 , 
    n2812 , 
    n2813 , 
    n2814 , 
    n2815 , 
    n2816 , 
    n2817 , 
    n2818 , 
    n2819 , 
    n2820 , 
    n2821 , 
    n2822 , 
    n2823 , 
    n2824 , 
    n2825 , 
    n2826 , 
    n2827 , 
    n2828 , 
    n2829 , 
    n2830 , 
    n2831 , 
    n2832 , 
    n2833 , 
    n2834 , 
    n2835 , 
    n2836 , 
    n2837 , 
    n2838 , 
    n2839 , 
    n2840 , 
    n2841 , 
    n2842 , 
    n2843 , 
    n2844 , 
    n2845 , 
    n2846 , 
    n2847 , 
    n2848 , 
    n2849 , 
    n2850 , 
    n2851 , 
    n2852 , 
    n2853 , 
    n2854 , 
    n2855 , 
    n2856 , 
    n2857 , 
    n2858 , 
    n2859 , 
    n2860 , 
    n2861 , 
    n2862 , 
    n2863 , 
    n2864 , 
    n2865 , 
    n2866 , 
    n2867 , 
    n2868 , 
    n2869 , 
    n2870 , 
    n2871 , 
    n2872 , 
    n2873 , 
    n2874 , 
    n2875 , 
    n2876 , 
    n2877 , 
    n2878 , 
    n2879 , 
    n2880 , 
    n2881 , 
    n2882 , 
    n2883 , 
    n2884 , 
    n2885 , 
    n2886 , 
    n2887 , 
    n2888 , 
    n2889 , 
    n2890 , 
    n2891 , 
    n2892 , 
    n2893 , 
    n2894 , 
    n2895 , 
    n2896 , 
    n2897 , 
    n2898 , 
    n2899 , 
    n2900 , 
    n2901 , 
    n2902 , 
    n2903 , 
    n2904 , 
    n2905 , 
    n2906 , 
    n2907 , 
    n2908 , 
    n2909 , 
    n2910 , 
    n2911 , 
    n2912 , 
    n2913 , 
    n2914 , 
    n2915 , 
    n2916 , 
    n2917 , 
    n2918 , 
    n2919 , 
    n2920 , 
    n2921 , 
    n2922 , 
    n2923 , 
    n2924 , 
    n2925 , 
    n2926 , 
    n2927 , 
    n2928 , 
    n2929 , 
    n2930 , 
    n2931 , 
    n2932 , 
    n2933 , 
    n2934 , 
    n2935 , 
    n2936 , 
    n2937 , 
    n2938 , 
    n2939 , 
    n2940 , 
    n2941 , 
    n2942 , 
    n2943 , 
    n2944 , 
    n2945 , 
    n2946 , 
    n2947 , 
    n2948 , 
    n2949 , 
    n2950 , 
    n2951 , 
    n2952 , 
    n2953 , 
    n2954 , 
    n2955 , 
    n2956 , 
    n2957 , 
    n2958 , 
    n2959 , 
    n2960 , 
    n2961 , 
    n2962 , 
    n2963 , 
    n2964 , 
    n2965 , 
    n2966 , 
    n2967 , 
    n2968 , 
    n2969 , 
    n2970 , 
    n2971 , 
    n2972 , 
    n2973 , 
    n2974 , 
    n2975 , 
    n2976 , 
    n2977 , 
    n2978 , 
    n2979 , 
    n2980 , 
    n2981 , 
    n2982 , 
    n2983 , 
    n2984 , 
    n2985 , 
    n2986 , 
    n2987 , 
    n2988 , 
    n2989 , 
    n2990 , 
    n2991 , 
    n2992 , 
    n2993 , 
    n2994 , 
    n2995 , 
    n2996 , 
    n2997 , 
    n2998 , 
    n2999 , 
    n3000 , 
    n3001 , 
    n3002 , 
    n3003 , 
    n3004 , 
    n3005 , 
    n3006 , 
    n3007 , 
    n3008 , 
    n3009 , 
    n3010 , 
    n3011 , 
    n3012 , 
    n3013 , 
    n3014 , 
    n3015 , 
    n3016 , 
    n3017 , 
    n3018 , 
    n3019 , 
    n3020 , 
    n3021 , 
    n3022 , 
    n3023 , 
    n3024 , 
    n3025 , 
    n3026 , 
    n3027 , 
    n3028 , 
    n3029 , 
    n3030 , 
    n3031 , 
    n3032 , 
    n3033 , 
    n3034 , 
    n3035 , 
    n3036 , 
    n3037 , 
    n3038 , 
    n3039 , 
    n3040 , 
    n3041 , 
    n3042 , 
    n3043 , 
    n3044 , 
    n3045 , 
    n3046 , 
    n3047 , 
    n3048 , 
    n3049 , 
    n3050 , 
    n3051 , 
    n3052 , 
    n3053 , 
    n3054 , 
    n3055 , 
    n3056 , 
    n3057 , 
    n3058 , 
    n3059 , 
    n3060 , 
    n3061 , 
    n3062 , 
    n3063 , 
    n3064 , 
    n3065 , 
    n3066 , 
    n3067 , 
    n3068 , 
    n3069 , 
    n3070 , 
    n3071 , 
    n3072 , 
    n3073 , 
    n3074 , 
    n3075 , 
    n3076 , 
    n3077 , 
    n3078 , 
    n3079 , 
    n3080 , 
    n3081 , 
    n3082 , 
    n3083 , 
    n3084 , 
    n3085 , 
    n3086 , 
    n3087 , 
    n3088 , 
    n3089 , 
    n3090 , 
    n3091 , 
    n3092 , 
    n3093 , 
    n3094 , 
    n3095 , 
    n3096 , 
    n3097 , 
    n3098 , 
    n3099 , 
    n3100 , 
    n3101 , 
    n3102 , 
    n3103 , 
    n3104 , 
    n3105 , 
    n3106 , 
    n3107 , 
    n3108 , 
    n3109 , 
    n3110 , 
    n3111 , 
    n3112 , 
    n3113 , 
    n3114 , 
    n3115 , 
    n3116 , 
    n3117 , 
    n3118 , 
    n3119 , 
    n3120 , 
    n3121 , 
    n3122 , 
    n3123 , 
    n3124 , 
    n3125 , 
    n3126 , 
    n3127 , 
    n3128 , 
    n3129 , 
    n3130 , 
    n3131 , 
    n3132 , 
    n3133 , 
    n3134 , 
    n3135 , 
    n3136 , 
    n3137 , 
    n3138 , 
    n3139 , 
    n3140 , 
    n3141 , 
    n3142 , 
    n3143 , 
    n3144 , 
    n3145 , 
    n3146 , 
    n3147 , 
    n3148 , 
    n3149 , 
    n3150 , 
    n3151 , 
    n3152 , 
    n3153 , 
    n3154 , 
    n3155 , 
    n3156 , 
    n3157 , 
    n3158 , 
    n3159 , 
    n3160 , 
    n3161 , 
    n3162 , 
    n3163 , 
    n3164 , 
    n3165 , 
    n3166 , 
    n3167 , 
    n3168 , 
    n3169 , 
    n3170 , 
    n3171 , 
    n3172 , 
    n3173 , 
    n3174 , 
    n3175 , 
    n3176 , 
    n3177 , 
    n3178 , 
    n3179 , 
    n3180 , 
    n3181 , 
    n3182 , 
    n3183 , 
    n3184 , 
    n3185 , 
    n3186 , 
    n3187 , 
    n3188 , 
    n3189 , 
    n3190 , 
    n3191 , 
    n3192 , 
    n3193 , 
    n3194 , 
    n3195 , 
    n3196 , 
    n3197 , 
    n3198 , 
    n3199 , 
    n3200 , 
    n3201 , 
    n3202 , 
    n3203 , 
    n3204 , 
    n3205 , 
    n3206 , 
    n3207 , 
    n3208 , 
    n3209 , 
    n3210 , 
    n3211 , 
    n3212 , 
    n3213 , 
    n3214 , 
    n3215 , 
    n3216 , 
    n3217 , 
    n3218 , 
    n3219 , 
    n3220 , 
    n3221 , 
    n3222 , 
    n3223 , 
    n3224 , 
    n3225 , 
    n3226 , 
    n3227 , 
    n3228 , 
    n3229 , 
    n3230 , 
    n3231 , 
    n3232 , 
    n3233 , 
    n3234 , 
    n3235 , 
    n3236 , 
    n3237 , 
    n3238 , 
    n3239 , 
    n3240 , 
    n3241 , 
    n3242 , 
    n3243 , 
    n3244 , 
    n3245 , 
    n3246 , 
    n3247 , 
    n3248 , 
    n3249 , 
    n3250 , 
    n3251 , 
    n3252 , 
    n3253 , 
    n3254 , 
    n3255 , 
    n3256 , 
    n3257 , 
    n3258 , 
    n3259 , 
    n3260 , 
    n3261 , 
    n3262 , 
    n3263 , 
    n3264 , 
    n3265 , 
    n3266 , 
    n3267 , 
    n3268 , 
    n3269 , 
    n3270 , 
    n3271 , 
    n3272 , 
    n3273 , 
    n3274 , 
    n3275 , 
    n3276 , 
    n3277 , 
    n3278 , 
    n3279 , 
    n3280 , 
    n3281 , 
    n3282 , 
    n3283 , 
    n3284 , 
    n3285 , 
    n3286 , 
    n3287 , 
    n3288 , 
    n3289 , 
    n3290 , 
    n3291 , 
    n3292 , 
    n3293 , 
    n3294 , 
    n3295 , 
    n3296 , 
    n3297 , 
    n3298 , 
    n3299 , 
    n3300 , 
    n3301 , 
    n3302 , 
    n3303 , 
    n3304 , 
    n3305 , 
    n3306 , 
    n3307 , 
    n3308 , 
    n3309 , 
    n3310 , 
    n3311 , 
    n3312 , 
    n3313 , 
    n3314 , 
    n3315 , 
    n3316 , 
    n3317 , 
    n3318 , 
    n3319 , 
    n3320 , 
    n3321 , 
    n3322 , 
    n3323 , 
    n3324 , 
    n3325 , 
    n3326 , 
    n3327 , 
    n3328 , 
    n3329 , 
    n3330 , 
    n3331 , 
    n3332 , 
    n3333 , 
    n3334 , 
    n3335 , 
    n3336 , 
    n3337 , 
    n3338 , 
    n3339 , 
    n3340 , 
    n3341 , 
    n3342 , 
    n3343 , 
    n3344 , 
    n3345 , 
    n3346 , 
    n3347 , 
    n3348 , 
    n3349 , 
    n3350 , 
    n3351 , 
    n3352 , 
    n3353 , 
    n3354 , 
    n3355 , 
    n3356 , 
    n3357 , 
    n3358 , 
    n3359 , 
    n3360 , 
    n3361 , 
    n3362 , 
    n3363 , 
    n3364 , 
    n3365 , 
    n3366 , 
    n3367 , 
    n3368 , 
    n3369 , 
    n3370 , 
    n3371 , 
    n3372 , 
    n3373 , 
    n3374 , 
    n3375 , 
    n3376 , 
    n3377 , 
    n3378 , 
    n3379 , 
    n3380 , 
    n3381 , 
    n3382 , 
    n3383 , 
    n3384 , 
    n3385 , 
    n3386 , 
    n3387 , 
    n3388 , 
    n3389 , 
    n3390 , 
    n3391 , 
    n3392 , 
    n3393 , 
    n3394 , 
    n3395 , 
    n3396 , 
    n3397 , 
    n3398 , 
    n3399 , 
    n3400 , 
    n3401 , 
    n3402 , 
    n3403 , 
    n3404 , 
    n3405 , 
    n3406 , 
    n3407 , 
    n3408 , 
    n3409 , 
    n3410 , 
    n3411 , 
    n3412 , 
    n3413 , 
    n3414 , 
    n3415 , 
    n3416 , 
    n3417 , 
    n3418 , 
    n3419 , 
    n3420 , 
    n3421 , 
    n3422 , 
    n3423 , 
    n3424 , 
    n3425 , 
    n3426 , 
    n3427 , 
    n3428 , 
    n3429 , 
    n3430 , 
    n3431 , 
    n3432 , 
    n3433 , 
    n3434 , 
    n3435 , 
    n3436 , 
    n3437 , 
    n3438 , 
    n3439 , 
    n3440 , 
    n3441 , 
    n3442 , 
    n3443 , 
    n3444 , 
    n3445 , 
    n3446 , 
    n3447 , 
    n3448 , 
    n3449 , 
    n3450 , 
    n3451 , 
    n3452 , 
    n3453 , 
    n3454 , 
    n3455 , 
    n3456 , 
    n3457 , 
    n3458 , 
    n3459 , 
    n3460 , 
    n3461 , 
    n3462 , 
    n3463 , 
    n3464 , 
    n3465 , 
    n3466 , 
    n3467 , 
    n3468 , 
    n3469 , 
    n3470 , 
    n3471 , 
    n3472 , 
    n3473 , 
    n3474 , 
    n3475 , 
    n3476 , 
    n3477 , 
    n3478 , 
    n3479 , 
    n3480 , 
    n3481 , 
    n3482 , 
    n3483 , 
    n3484 , 
    n3485 , 
    n3486 , 
    n3487 , 
    n3488 , 
    n3489 , 
    n3490 , 
    n3491 , 
    n3492 , 
    n3493 , 
    n3494 , 
    n3495 , 
    n3496 , 
    n3497 , 
    n3498 , 
    n3499 , 
    n3500 , 
    n3501 , 
    n3502 , 
    n3503 , 
    n3504 , 
    n3505 , 
    n3506 , 
    n3507 , 
    n3508 , 
    n3509 , 
    n3510 , 
    n3511 , 
    n3512 , 
    n3513 , 
    n3514 , 
    n3515 , 
    n3516 , 
    n3517 , 
    n3518 , 
    n3519 , 
    n3520 , 
    n3521 , 
    n3522 , 
    n3523 , 
    n3524 , 
    n3525 , 
    n3526 , 
    n3527 , 
    n3528 , 
    n3529 , 
    n3530 , 
    n3531 , 
    n3532 , 
    n3533 , 
    n3534 , 
    n3535 , 
    n3536 , 
    n3537 , 
    n3538 , 
    n3539 , 
    n3540 , 
    n3541 , 
    n3542 , 
    n3543 , 
    n3544 , 
    n3545 , 
    n3546 , 
    n3547 , 
    n3548 , 
    n3549 , 
    n3550 , 
    n3551 , 
    n3552 , 
    n3553 , 
    n3554 , 
    n3555 , 
    n3556 , 
    n3557 , 
    n3558 , 
    n3559 , 
    n3560 , 
    n3561 , 
    n3562 , 
    n3563 , 
    n3564 , 
    n3565 , 
    n3566 , 
    n3567 , 
    n3568 , 
    n3569 , 
    n3570 , 
    n3571 , 
    n3572 , 
    n3573 , 
    n3574 , 
    n3575 , 
    n3576 , 
    n3577 , 
    n3578 , 
    n3579 , 
    n3580 , 
    n3581 , 
    n3582 , 
    n3583 , 
    n3584 , 
    n3585 , 
    n3586 , 
    n3587 , 
    n3588 , 
    n3589 , 
    n3590 , 
    n3591 , 
    n3592 , 
    n3593 , 
    n3594 , 
    n3595 , 
    n3596 , 
    n3597 , 
    n3598 , 
    n3599 , 
    n3600 , 
    n3601 , 
    n3602 , 
    n3603 , 
    n3604 , 
    n3605 , 
    n3606 , 
    n3607 , 
    n3608 , 
    n3609 , 
    n3610 , 
    n3611 , 
    n3612 , 
    n3613 , 
    n3614 , 
    n3615 , 
    n3616 , 
    n3617 , 
    n3618 , 
    n3619 , 
    n3620 , 
    n3621 , 
    n3622 , 
    n3623 , 
    n3624 , 
    n3625 , 
    n3626 , 
    n3627 , 
    n3628 , 
    n3629 , 
    n3630 , 
    n3631 , 
    n3632 , 
    n3633 , 
    n3634 , 
    n3635 , 
    n3636 , 
    n3637 , 
    n3638 , 
    n3639 , 
    n3640 , 
    n3641 , 
    n3642 , 
    n3643 , 
    n3644 , 
    n3645 , 
    n3646 , 
    n3647 , 
    n3648 , 
    n3649 , 
    n3650 , 
    n3651 , 
    n3652 , 
    n3653 , 
    n3654 , 
    n3655 , 
    n3656 , 
    n3657 , 
    n3658 , 
    n3659 , 
    n3660 , 
    n3661 , 
    n3662 , 
    n3663 , 
    n3664 , 
    n3665 , 
    n3666 , 
    n3667 , 
    n3668 , 
    n3669 , 
    n3670 , 
    n3671 , 
    n3672 , 
    n3673 , 
    n3674 , 
    n3675 , 
    n3676 , 
    n3677 , 
    n3678 , 
    n3679 , 
    n3680 , 
    n3681 , 
    n3682 , 
    n3683 , 
    n3684 , 
    n3685 , 
    n3686 , 
    n3687 , 
    n3688 , 
    n3689 , 
    n3690 , 
    n3691 , 
    n3692 , 
    n3693 , 
    n3694 , 
    n3695 , 
    n3696 , 
    n3697 , 
    n3698 , 
    n3699 , 
    n3700 , 
    n3701 , 
    n3702 , 
    n3703 , 
    n3704 , 
    n3705 , 
    n3706 , 
    n3707 , 
    n3708 , 
    n3709 , 
    n3710 , 
    n3711 , 
    n3712 , 
    n3713 , 
    n3714 , 
    n3715 , 
    n3716 , 
    n3717 , 
    n3718 , 
    n3719 , 
    n3720 , 
    n3721 , 
    n3722 , 
    n3723 , 
    n3724 , 
    n3725 , 
    n3726 , 
    n3727 , 
    n3728 , 
    n3729 , 
    n3730 , 
    n3731 , 
    n3732 , 
    n3733 , 
    n3734 , 
    n3735 , 
    n3736 , 
    n3737 , 
    n3738 , 
    n3739 , 
    n3740 , 
    n3741 , 
    n3742 , 
    n3743 , 
    n3744 , 
    n3745 , 
    n3746 , 
    n3747 , 
    n3748 , 
    n3749 , 
    n3750 , 
    n3751 , 
    n3752 , 
    n3753 , 
    n3754 , 
    n3755 , 
    n3756 , 
    n3757 , 
    n3758 , 
    n3759 , 
    n3760 , 
    n3761 , 
    n3762 , 
    n3763 , 
    n3764 , 
    n3765 , 
    n3766 , 
    n3767 , 
    n3768 , 
    n3769 , 
    n3770 , 
    n3771 , 
    n3772 , 
    n3773 , 
    n3774 , 
    n3775 , 
    n3776 , 
    n3777 , 
    n3778 , 
    n3779 , 
    n3780 , 
    n3781 , 
    n3782 , 
    n3783 , 
    n3784 , 
    n3785 , 
    n3786 , 
    n3787 , 
    n3788 , 
    n3789 , 
    n3790 , 
    n3791 , 
    n3792 , 
    n3793 , 
    n3794 , 
    n3795 , 
    n3796 , 
    n3797 , 
    n3798 , 
    n3799 , 
    n3800 , 
    n3801 , 
    n3802 , 
    n3803 , 
    n3804 , 
    n3805 , 
    n3806 , 
    n3807 , 
    n3808 , 
    n3809 , 
    n3810 , 
    n3811 , 
    n3812 , 
    n3813 , 
    n3814 , 
    n3815 , 
    n3816 , 
    n3817 , 
    n3818 , 
    n3819 , 
    n3820 , 
    n3821 , 
    n3822 , 
    n3823 , 
    n3824 , 
    n3825 , 
    n3826 , 
    n3827 , 
    n3828 , 
    n3829 , 
    n3830 , 
    n3831 , 
    n3832 , 
    n3833 , 
    n3834 , 
    n3835 , 
    n3836 , 
    n3837 , 
    n3838 , 
    n3839 , 
    n3840 , 
    n3841 , 
    n3842 , 
    n3843 , 
    n3844 , 
    n3845 , 
    n3846 , 
    n3847 , 
    n3848 , 
    n3849 , 
    n3850 , 
    n3851 , 
    n3852 , 
    n3853 , 
    n3854 , 
    n3855 , 
    n3856 , 
    n3857 , 
    n3858 , 
    n3859 , 
    n3860 , 
    n3861 , 
    n3862 , 
    n3863 , 
    n3864 , 
    n3865 , 
    n3866 , 
    n3867 , 
    n3868 , 
    n3869 , 
    n3870 , 
    n3871 , 
    n3872 , 
    n3873 , 
    n3874 , 
    n3875 , 
    n3876 , 
    n3877 , 
    n3878 , 
    n3879 , 
    n3880 , 
    n3881 , 
    n3882 , 
    n3883 , 
    n3884 , 
    n3885 , 
    n3886 , 
    n3887 , 
    n3888 , 
    n3889 , 
    n3890 , 
    n3891 , 
    n3892 , 
    n3893 , 
    n3894 , 
    n3895 , 
    n3896 , 
    n3897 , 
    n3898 , 
    n3899 , 
    n3900 , 
    n3901 , 
    n3902 , 
    n3903 , 
    n3904 , 
    n3905 , 
    n3906 , 
    n3907 , 
    n3908 , 
    n3909 , 
    n3910 , 
    n3911 , 
    n3912 , 
    n3913 , 
    n3914 , 
    n3915 , 
    n3916 , 
    n3917 , 
    n3918 , 
    n3919 , 
    n3920 , 
    n3921 , 
    n3922 , 
    n3923 , 
    n3924 , 
    n3925 , 
    n3926 , 
    n3927 , 
    n3928 , 
    n3929 , 
    n3930 , 
    n3931 , 
    n3932 , 
    n3933 , 
    n3934 , 
    n3935 , 
    n3936 , 
    n3937 , 
    n3938 , 
    n3939 , 
    n3940 , 
    n3941 , 
    n3942 , 
    n3943 , 
    n3944 , 
    n3945 , 
    n3946 , 
    n3947 , 
    n3948 , 
    n3949 , 
    n3950 , 
    n3951 , 
    n3952 , 
    n3953 , 
    n3954 , 
    n3955 , 
    n3956 , 
    n3957 , 
    n3958 , 
    n3959 , 
    n3960 , 
    n3961 , 
    n3962 , 
    n3963 , 
    n3964 , 
    n3965 , 
    n3966 , 
    n3967 , 
    n3968 , 
    n3969 , 
    n3970 , 
    n3971 , 
    n3972 , 
    n3973 , 
    n3974 , 
    n3975 , 
    n3976 , 
    n3977 , 
    n3978 , 
    n3979 , 
    n3980 , 
    n3981 , 
    n3982 , 
    n3983 , 
    n3984 , 
    n3985 , 
    n3986 , 
    n3987 , 
    n3988 , 
    n3989 , 
    n3990 , 
    n3991 , 
    n3992 , 
    n3993 , 
    n3994 , 
    n3995 , 
    n3996 , 
    n3997 , 
    n3998 , 
    n3999 , 
    n4000 , 
    n4001 , 
    n4002 , 
    n4003 , 
    n4004 , 
    n4005 , 
    n4006 , 
    n4007 , 
    n4008 , 
    n4009 , 
    n4010 , 
    n4011 , 
    n4012 , 
    n4013 , 
    n4014 , 
    n4015 , 
    n4016 , 
    n4017 , 
    n4018 , 
    n4019 , 
    n4020 , 
    n4021 , 
    n4022 , 
    n4023 , 
    n4024 , 
    n4025 , 
    n4026 , 
    n4027 , 
    n4028 , 
    n4029 , 
    n4030 , 
    n4031 , 
    n4032 , 
    n4033 , 
    n4034 , 
    n4035 , 
    n4036 , 
    n4037 , 
    n4038 , 
    n4039 , 
    n4040 , 
    n4041 , 
    n4042 , 
    n4043 , 
    n4044 , 
    n4045 , 
    n4046 , 
    n4047 , 
    n4048 , 
    n4049 , 
    n4050 , 
    n4051 , 
    n4052 , 
    n4053 , 
    n4054 , 
    n4055 , 
    n4056 , 
    n4057 , 
    n4058 , 
    n4059 , 
    n4060 , 
    n4061 , 
    n4062 , 
    n4063 , 
    n4064 , 
    n4065 , 
    n4066 , 
    n4067 , 
    n4068 , 
    n4069 , 
    n4070 , 
    n4071 , 
    n4072 , 
    n4073 , 
    n4074 , 
    n4075 , 
    n4076 , 
    n4077 , 
    n4078 , 
    n4079 , 
    n4080 , 
    n4081 , 
    n4082 , 
    n4083 , 
    n4084 , 
    n4085 , 
    n4086 , 
    n4087 , 
    n4088 , 
    n4089 , 
    n4090 , 
    n4091 , 
    n4092 , 
    n4093 , 
    n4094 , 
    n4095 , 
    n4096 , 
    n4097 , 
    n4098 , 
    n4099 , 
    n4100 , 
    n4101 , 
    n4102 , 
    n4103 , 
    n4104 , 
    n4105 , 
    n4106 , 
    n4107 , 
    n4108 , 
    n4109 , 
    n4110 , 
    n4111 , 
    n4112 , 
    n4113 , 
    n4114 , 
    n4115 , 
    n4116 , 
    n4117 , 
    n4118 , 
    n4119 , 
    n4120 , 
    n4121 , 
    n4122 , 
    n4123 , 
    n4124 , 
    n4125 , 
    n4126 , 
    n4127 , 
    n4128 , 
    n4129 , 
    n4130 , 
    n4131 , 
    n4132 , 
    n4133 , 
    n4134 , 
    n4135 , 
    n4136 , 
    n4137 , 
    n4138 , 
    n4139 , 
    n4140 , 
    n4141 , 
    n4142 , 
    n4143 , 
    n4144 , 
    n4145 , 
    n4146 , 
    n4147 , 
    n4148 , 
    n4149 , 
    n4150 , 
    n4151 , 
    n4152 , 
    n4153 , 
    n4154 , 
    n4155 , 
    n4156 , 
    n4157 , 
    n4158 , 
    n4159 , 
    n4160 , 
    n4161 , 
    n4162 , 
    n4163 , 
    n4164 , 
    n4165 , 
    n4166 , 
    n4167 , 
    n4168 , 
    n4169 , 
    n4170 , 
    n4171 , 
    n4172 , 
    n4173 , 
    n4174 , 
    n4175 , 
    n4176 , 
    n4177 , 
    n4178 , 
    n4179 , 
    n4180 , 
    n4181 , 
    n4182 , 
    n4183 , 
    n4184 , 
    n4185 , 
    n4186 , 
    n4187 , 
    n4188 , 
    n4189 , 
    n4190 , 
    n4191 , 
    n4192 , 
    n4193 , 
    n4194 , 
    n4195 , 
    n4196 , 
    n4197 , 
    n4198 , 
    n4199 , 
    n4200 , 
    n4201 , 
    n4202 , 
    n4203 , 
    n4204 , 
    n4205 , 
    n4206 , 
    n4207 , 
    n4208 , 
    n4209 , 
    n4210 , 
    n4211 , 
    n4212 , 
    n4213 , 
    n4214 , 
    n4215 , 
    n4216 , 
    n4217 , 
    n4218 , 
    n4219 , 
    n4220 , 
    n4221 , 
    n4222 , 
    n4223 , 
    n4224 , 
    n4225 , 
    n4226 , 
    n4227 , 
    n4228 , 
    n4229 , 
    n4230 , 
    n4231 , 
    n4232 , 
    n4233 , 
    n4234 , 
    n4235 , 
    n4236 , 
    n4237 , 
    n4238 , 
    n4239 , 
    n4240 , 
    n4241 , 
    n4242 , 
    n4243 , 
    n4244 , 
    n4245 , 
    n4246 , 
    n4247 , 
    n4248 , 
    n4249 , 
    n4250 , 
    n4251 , 
    n4252 , 
    n4253 , 
    n4254 , 
    n4255 , 
    n4256 , 
    n4257 , 
    n4258 , 
    n4259 , 
    n4260 , 
    n4261 , 
    n4262 , 
    n4263 , 
    n4264 , 
    n4265 , 
    n4266 , 
    n4267 , 
    n4268 , 
    n4269 , 
    n4270 , 
    n4271 , 
    n4272 , 
    n4273 , 
    n4274 , 
    n4275 , 
    n4276 , 
    n4277 , 
    n4278 , 
    n4279 , 
    n4280 , 
    n4281 , 
    n4282 , 
    n4283 , 
    n4284 , 
    n4285 , 
    n4286 , 
    n4287 , 
    n4288 , 
    n4289 , 
    n4290 , 
    n4291 , 
    n4292 , 
    n4293 , 
    n4294 , 
    n4295 , 
    n4296 , 
    n4297 , 
    n4298 , 
    n4299 , 
    n4300 , 
    n4301 , 
    n4302 , 
    n4303 , 
    n4304 , 
    n4305 , 
    n4306 , 
    n4307 , 
    n4308 , 
    n4309 , 
    n4310 , 
    n4311 , 
    n4312 , 
    n4313 , 
    n4314 , 
    n4315 , 
    n4316 , 
    n4317 , 
    n4318 , 
    n4319 , 
    n4320 , 
    n4321 , 
    n4322 , 
    n4323 , 
    n4324 , 
    n4325 , 
    n4326 , 
    n4327 , 
    n4328 , 
    n4329 , 
    n4330 , 
    n4331 , 
    n4332 , 
    n4333 , 
    n4334 , 
    n4335 , 
    n4336 , 
    n4337 , 
    n4338 , 
    n4339 , 
    n4340 , 
    n4341 , 
    n4342 , 
    n4343 , 
    n4344 , 
    n4345 , 
    n4346 , 
    n4347 , 
    n4348 , 
    n4349 , 
    n4350 , 
    n4351 , 
    n4352 , 
    n4353 , 
    n4354 , 
    n4355 , 
    n4356 , 
    n4357 , 
    n4358 , 
    n4359 , 
    n4360 , 
    n4361 , 
    n4362 , 
    n4363 , 
    n4364 , 
    n4365 , 
    n4366 , 
    n4367 , 
    n4368 , 
    n4369 , 
    n4370 , 
    n4371 , 
    n4372 , 
    n4373 , 
    n4374 , 
    n4375 , 
    n4376 , 
    n4377 , 
    n4378 , 
    n4379 , 
    n4380 , 
    n4381 , 
    n4382 , 
    n4383 , 
    n4384 , 
    n4385 , 
    n4386 , 
    n4387 , 
    n4388 , 
    n4389 , 
    n4390 , 
    n4391 , 
    n4392 , 
    n4393 , 
    n4394 , 
    n4395 , 
    n4396 , 
    n4397 , 
    n4398 , 
    n4399 , 
    n4400 , 
    n4401 , 
    n4402 , 
    n4403 , 
    n4404 , 
    n4405 , 
    n4406 , 
    n4407 , 
    n4408 , 
    n4409 , 
    n4410 , 
    n4411 , 
    n4412 , 
    n4413 , 
    n4414 , 
    n4415 , 
    n4416 , 
    n4417 , 
    n4418 , 
    n4419 , 
    n4420 , 
    n4421 , 
    n4422 , 
    n4423 , 
    n4424 , 
    n4425 , 
    n4426 , 
    n4427 , 
    n4428 , 
    n4429 , 
    n4430 , 
    n4431 , 
    n4432 , 
    n4433 , 
    n4434 , 
    n4435 , 
    n4436 , 
    n4437 , 
    n4438 , 
    n4439 , 
    n4440 , 
    n4441 , 
    n4442 , 
    n4443 , 
    n4444 , 
    n4445 , 
    n4446 , 
    n4447 , 
    n4448 , 
    n4449 , 
    n4450 , 
    n4451 , 
    n4452 , 
    n4453 , 
    n4454 , 
    n4455 , 
    n4456 , 
    n4457 , 
    n4458 , 
    n4459 , 
    n4460 , 
    n4461 , 
    n4462 , 
    n4463 , 
    n4464 , 
    n4465 , 
    n4466 , 
    n4467 , 
    n4468 , 
    n4469 , 
    n4470 , 
    n4471 , 
    n4472 , 
    n4473 , 
    n4474 , 
    n4475 , 
    n4476 , 
    n4477 , 
    n4478 , 
    n4479 , 
    n4480 , 
    n4481 , 
    n4482 , 
    n4483 , 
    n4484 , 
    n4485 , 
    n4486 , 
    n4487 , 
    n4488 , 
    n4489 , 
    n4490 , 
    n4491 , 
    n4492 , 
    n4493 , 
    n4494 , 
    n4495 , 
    n4496 , 
    n4497 , 
    n4498 , 
    n4499 , 
    n4500 , 
    n4501 , 
    n4502 , 
    n4503 , 
    n4504 , 
    n4505 , 
    n4506 , 
    n4507 , 
    n4508 , 
    n4509 , 
    n4510 , 
    n4511 , 
    n4512 , 
    n4513 , 
    n4514 , 
    n4515 , 
    n4516 , 
    n4517 , 
    n4518 , 
    n4519 , 
    n4520 , 
    n4521 , 
    n4522 , 
    n4523 , 
    n4524 , 
    n4525 , 
    n4526 , 
    n4527 , 
    n4528 , 
    n4529 , 
    n4530 , 
    n4531 , 
    n4532 , 
    n4533 , 
    n4534 , 
    n4535 , 
    n4536 , 
    n4537 , 
    n4538 , 
    n4539 , 
    n4540 , 
    n4541 , 
    n4542 , 
    n4543 , 
    n4544 , 
    n4545 , 
    n4546 , 
    n4547 , 
    n4548 , 
    n4549 , 
    n4550 , 
    n4551 , 
    n4552 , 
    n4553 , 
    n4554 , 
    n4555 , 
    n4556 , 
    n4557 , 
    n4558 , 
    n4559 , 
    n4560 , 
    n4561 , 
    n4562 , 
    n4563 , 
    n4564 , 
    n4565 , 
    n4566 , 
    n4567 , 
    n4568 , 
    n4569 , 
    n4570 , 
    n4571 , 
    n4572 , 
    n4573 , 
    n4574 , 
    n4575 , 
    n4576 , 
    n4577 , 
    n4578 , 
    n4579 , 
    n4580 , 
    n4581 , 
    n4582 , 
    n4583 , 
    n4584 , 
    n4585 , 
    n4586 , 
    n4587 , 
    n4588 , 
    n4589 , 
    n4590 , 
    n4591 , 
    n4592 , 
    n4593 , 
    n4594 , 
    n4595 , 
    n4596 , 
    n4597 , 
    n4598 , 
    n4599 , 
    n4600 , 
    n4601 , 
    n4602 , 
    n4603 , 
    n4604 , 
    n4605 , 
    n4606 , 
    n4607 , 
    n4608 , 
    n4609 , 
    n4610 , 
    n4611 , 
    n4612 , 
    n4613 , 
    n4614 , 
    n4615 , 
    n4616 , 
    n4617 , 
    n4618 , 
    n4619 , 
    n4620 , 
    n4621 , 
    n4622 , 
    n4623 , 
    n4624 , 
    n4625 , 
    n4626 , 
    n4627 , 
    n4628 , 
    n4629 , 
    n4630 , 
    n4631 , 
    n4632 , 
    n4633 , 
    n4634 , 
    n4635 , 
    n4636 , 
    n4637 , 
    n4638 , 
    n4639 , 
    n4640 , 
    n4641 , 
    n4642 , 
    n4643 , 
    n4644 , 
    n4645 , 
    n4646 , 
    n4647 , 
    n4648 , 
    n4649 , 
    n4650 , 
    n4651 , 
    n4652 , 
    n4653 , 
    n4654 , 
    n4655 , 
    n4656 , 
    n4657 , 
    n4658 , 
    n4659 , 
    n4660 , 
    n4661 , 
    n4662 , 
    n4663 , 
    n4664 , 
    n4665 , 
    n4666 , 
    n4667 , 
    n4668 , 
    n4669 , 
    n4670 , 
    n4671 , 
    n4672 , 
    n4673 , 
    n4674 , 
    n4675 , 
    n4676 , 
    n4677 , 
    n4678 , 
    n4679 , 
    n4680 , 
    n4681 , 
    n4682 , 
    n4683 , 
    n4684 , 
    n4685 , 
    n4686 , 
    n4687 , 
    n4688 , 
    n4689 , 
    n4690 , 
    n4691 , 
    n4692 , 
    n4693 , 
    n4694 , 
    n4695 , 
    n4696 , 
    n4697 , 
    n4698 , 
    n4699 , 
    n4700 , 
    n4701 , 
    n4702 , 
    n4703 , 
    n4704 , 
    n4705 , 
    n4706 , 
    n4707 , 
    n4708 , 
    n4709 , 
    n4710 , 
    n4711 , 
    n4712 , 
    n4713 , 
    n4714 , 
    n4715 , 
    n4716 , 
    n4717 , 
    n4718 , 
    n4719 , 
    n4720 , 
    n4721 , 
    n4722 , 
    n4723 , 
    n4724 , 
    n4725 , 
    n4726 , 
    n4727 , 
    n4728 , 
    n4729 , 
    n4730 , 
    n4731 , 
    n4732 , 
    n4733 , 
    n4734 , 
    n4735 , 
    n4736 , 
    n4737 , 
    n4738 , 
    n4739 , 
    n4740 , 
    n4741 , 
    n4742 , 
    n4743 , 
    n4744 , 
    n4745 , 
    n4746 , 
    n4747 , 
    n4748 , 
    n4749 , 
    n4750 , 
    n4751 , 
    n4752 , 
    n4753 , 
    n4754 , 
    n4755 , 
    n4756 , 
    n4757 , 
    n4758 , 
    n4759 , 
    n4760 , 
    n4761 , 
    n4762 , 
    n4763 , 
    n4764 , 
    n4765 , 
    n4766 , 
    n4767 , 
    n4768 , 
    n4769 , 
    n4770 , 
    n4771 , 
    n4772 , 
    n4773 , 
    n4774 , 
    n4775 , 
    n4776 , 
    n4777 , 
    n4778 , 
    n4779 , 
    n4780 , 
    n4781 , 
    n4782 , 
    n4783 , 
    n4784 , 
    n4785 , 
    n4786 , 
    n4787 , 
    n4788 , 
    n4789 , 
    n4790 , 
    n4791 , 
    n4792 , 
    n4793 , 
    n4794 , 
    n4795 , 
    n4796 , 
    n4797 , 
    n4798 , 
    n4799 , 
    n4800 , 
    n4801 , 
    n4802 , 
    n4803 , 
    n4804 , 
    n4805 , 
    n4806 , 
    n4807 , 
    n4808 , 
    n4809 , 
    n4810 , 
    n4811 , 
    n4812 , 
    n4813 , 
    n4814 , 
    n4815 , 
    n4816 , 
    n4817 , 
    n4818 , 
    n4819 , 
    n4820 , 
    n4821 , 
    n4822 , 
    n4823 , 
    n4824 , 
    n4825 , 
    n4826 , 
    n4827 , 
    n4828 , 
    n4829 , 
    n4830 , 
    n4831 , 
    n4832 , 
    n4833 , 
    n4834 , 
    n4835 , 
    n4836 , 
    n4837 , 
    n4838 , 
    n4839 , 
    n4840 , 
    n4841 , 
    n4842 , 
    n4843 , 
    n4844 , 
    n4845 , 
    n4846 , 
    n4847 , 
    n4848 , 
    n4849 , 
    n4850 , 
    n4851 , 
    n4852 , 
    n4853 , 
    n4854 , 
    n4855 , 
    n4856 , 
    n4857 , 
    n4858 , 
    n4859 , 
    n4860 , 
    n4861 , 
    n4862 , 
    n4863 , 
    n4864 , 
    n4865 , 
    n4866 , 
    n4867 , 
    n4868 , 
    n4869 , 
    n4870 , 
    n4871 , 
    n4872 , 
    n4873 , 
    n4874 , 
    n4875 , 
    n4876 , 
    n4877 , 
    n4878 , 
    n4879 , 
    n4880 , 
    n4881 , 
    n4882 , 
    n4883 , 
    n4884 , 
    n4885 , 
    n4886 , 
    n4887 , 
    n4888 , 
    n4889 , 
    n4890 , 
    n4891 , 
    n4892 , 
    n4893 , 
    n4894 , 
    n4895 , 
    n4896 , 
    n4897 , 
    n4898 , 
    n4899 , 
    n4900 , 
    n4901 , 
    n4902 , 
    n4903 , 
    n4904 , 
    n4905 , 
    n4906 , 
    n4907 , 
    n4908 , 
    n4909 , 
    n4910 , 
    n4911 , 
    n4912 , 
    n4913 , 
    n4914 , 
    n4915 , 
    n4916 , 
    n4917 , 
    n4918 , 
    n4919 , 
    n4920 , 
    n4921 , 
    n4922 , 
    n4923 , 
    n4924 , 
    n4925 , 
    n4926 , 
    n4927 , 
    n4928 , 
    n4929 , 
    n4930 , 
    n4931 , 
    n4932 , 
    n4933 , 
    n4934 , 
    n4935 , 
    n4936 , 
    n4937 , 
    n4938 , 
    n4939 , 
    n4940 , 
    n4941 , 
    n4942 , 
    n4943 , 
    n4944 , 
    n4945 , 
    n4946 , 
    n4947 , 
    n4948 , 
    n4949 , 
    n4950 , 
    n4951 , 
    n4952 , 
    n4953 , 
    n4954 , 
    n4955 , 
    n4956 , 
    n4957 , 
    n4958 , 
    n4959 , 
    n4960 , 
    n4961 , 
    n4962 , 
    n4963 , 
    n4964 , 
    n4965 , 
    n4966 , 
    n4967 , 
    n4968 , 
    n4969 , 
    n4970 , 
    n4971 , 
    n4972 , 
    n4973 , 
    n4974 , 
    n4975 , 
    n4976 , 
    n4977 , 
    n4978 , 
    n4979 , 
    n4980 , 
    n4981 , 
    n4982 , 
    n4983 , 
    n4984 , 
    n4985 , 
    n4986 , 
    n4987 , 
    n4988 , 
    n4989 , 
    n4990 , 
    n4991 , 
    n4992 , 
    n4993 , 
    n4994 , 
    n4995 , 
    n4996 , 
    n4997 , 
    n4998 , 
    n4999 , 
    n5000 , 
    n5001 , 
    n5002 , 
    n5003 , 
    n5004 , 
    n5005 , 
    n5006 , 
    n5007 , 
    n5008 , 
    n5009 , 
    n5010 , 
    n5011 , 
    n5012 , 
    n5013 , 
    n5014 , 
    n5015 , 
    n5016 , 
    n5017 , 
    n5018 , 
    n5019 , 
    n5020 , 
    n5021 , 
    n5022 , 
    n5023 , 
    n5024 , 
    n5025 , 
    n5026 , 
    n5027 , 
    n5028 , 
    n5029 , 
    n5030 , 
    n5031 , 
    n5032 , 
    n5033 , 
    n5034 , 
    n5035 , 
    n5036 , 
    n5037 , 
    n5038 , 
    n5039 , 
    n5040 , 
    n5041 , 
    n5042 , 
    n5043 , 
    n5044 , 
    n5045 , 
    n5046 , 
    n5047 , 
    n5048 , 
    n5049 , 
    n5050 , 
    n5051 , 
    n5052 , 
    n5053 , 
    n5054 , 
    n5055 , 
    n5056 , 
    n5057 , 
    n5058 , 
    n5059 , 
    n5060 , 
    n5061 , 
    n5062 , 
    n5063 , 
    n5064 , 
    n5065 , 
    n5066 , 
    n5067 , 
    n5068 , 
    n5069 , 
    n5070 , 
    n5071 , 
    n5072 , 
    n5073 , 
    n5074 , 
    n5075 , 
    n5076 , 
    n5077 , 
    n5078 , 
    n5079 , 
    n5080 , 
    n5081 , 
    n5082 , 
    n5083 , 
    n5084 , 
    n5085 , 
    n5086 , 
    n5087 , 
    n5088 , 
    n5089 , 
    n5090 , 
    n5091 , 
    n5092 , 
    n5093 , 
    n5094 , 
    n5095 , 
    n5096 , 
    n5097 , 
    n5098 , 
    n5099 , 
    n5100 , 
    n5101 , 
    n5102 , 
    n5103 , 
    n5104 , 
    n5105 , 
    n5106 , 
    n5107 , 
    n5108 , 
    n5109 , 
    n5110 , 
    n5111 , 
    n5112 , 
    n5113 , 
    n5114 , 
    n5115 , 
    n5116 , 
    n5117 , 
    n5118 , 
    n5119 , 
    n5120 , 
    n5121 , 
    n5122 , 
    n5123 , 
    n5124 , 
    n5125 , 
    n5126 , 
    n5127 , 
    n5128 , 
    n5129 , 
    n5130 , 
    n5131 , 
    n5132 , 
    n5133 , 
    n5134 , 
    n5135 , 
    n5136 , 
    n5137 , 
    n5138 , 
    n5139 , 
    n5140 , 
    n5141 , 
    n5142 , 
    n5143 , 
    n5144 , 
    n5145 , 
    n5146 , 
    n5147 , 
    n5148 , 
    n5149 , 
    n5150 , 
    n5151 , 
    n5152 , 
    n5153 , 
    n5154 , 
    n5155 , 
    n5156 , 
    n5157 , 
    n5158 , 
    n5159 , 
    n5160 , 
    n5161 , 
    n5162 , 
    n5163 , 
    n5164 , 
    n5165 , 
    n5166 , 
    n5167 , 
    n5168 , 
    n5169 , 
    n5170 , 
    n5171 , 
    n5172 , 
    n5173 , 
    n5174 , 
    n5175 , 
    n5176 , 
    n5177 , 
    n5178 , 
    n5179 , 
    n5180 , 
    n5181 , 
    n5182 , 
    n5183 , 
    n5184 , 
    n5185 , 
    n5186 , 
    n5187 , 
    n5188 , 
    n5189 , 
    n5190 , 
    n5191 , 
    n5192 , 
    n5193 , 
    n5194 , 
    n5195 , 
    n5196 , 
    n5197 , 
    n5198 , 
    n5199 , 
    n5200 , 
    n5201 , 
    n5202 , 
    n5203 , 
    n5204 , 
    n5205 , 
    n5206 , 
    n5207 , 
    n5208 , 
    n5209 , 
    n5210 , 
    n5211 , 
    n5212 , 
    n5213 , 
    n5214 , 
    n5215 , 
    n5216 , 
    n5217 , 
    n5218 , 
    n5219 , 
    n5220 , 
    n5221 , 
    n5222 , 
    n5223 , 
    n5224 , 
    n5225 , 
    n5226 , 
    n5227 , 
    n5228 , 
    n5229 , 
    n5230 , 
    n5231 , 
    n5232 , 
    n5233 , 
    n5234 , 
    n5235 , 
    n5236 , 
    n5237 , 
    n5238 , 
    n5239 , 
    n5240 , 
    n5241 , 
    n5242 , 
    n5243 , 
    n5244 , 
    n5245 , 
    n5246 , 
    n5247 , 
    n5248 , 
    n5249 , 
    n5250 , 
    n5251 , 
    n5252 , 
    n5253 , 
    n5254 , 
    n5255 , 
    n5256 , 
    n5257 , 
    n5258 , 
    n5259 , 
    n5260 , 
    n5261 , 
    n5262 , 
    n5263 , 
    n5264 , 
    n5265 , 
    n5266 , 
    n5267 , 
    n5268 , 
    n5269 , 
    n5270 , 
    n5271 , 
    n5272 , 
    n5273 , 
    n5274 , 
    n5275 , 
    n5276 , 
    n5277 , 
    n5278 , 
    n5279 , 
    n5280 , 
    n5281 , 
    n5282 , 
    n5283 , 
    n5284 , 
    n5285 , 
    n5286 , 
    n5287 , 
    n5288 , 
    n5289 , 
    n5290 , 
    n5291 , 
    n5292 , 
    n5293 , 
    n5294 , 
    n5295 , 
    n5296 , 
    n5297 , 
    n5298 , 
    n5299 , 
    n5300 , 
    n5301 , 
    n5302 , 
    n5303 , 
    n5304 , 
    n5305 , 
    n5306 , 
    n5307 , 
    n5308 , 
    n5309 , 
    n5310 , 
    n5311 , 
    n5312 , 
    n5313 , 
    n5314 , 
    n5315 , 
    n5316 , 
    n5317 , 
    n5318 , 
    n5319 , 
    n5320 , 
    n5321 , 
    n5322 , 
    n5323 , 
    n5324 , 
    n5325 , 
    n5326 , 
    n5327 , 
    n5328 , 
    n5329 , 
    n5330 , 
    n5331 , 
    n5332 , 
    n5333 , 
    n5334 , 
    n5335 , 
    n5336 , 
    n5337 , 
    n5338 , 
    n5339 , 
    n5340 , 
    n5341 , 
    n5342 , 
    n5343 , 
    n5344 , 
    n5345 , 
    n5346 , 
    n5347 , 
    n5348 , 
    n5349 , 
    n5350 , 
    n5351 , 
    n5352 , 
    n5353 , 
    n5354 , 
    n5355 , 
    n5356 , 
    n5357 , 
    n5358 , 
    n5359 , 
    n5360 , 
    n5361 , 
    n5362 , 
    n5363 , 
    n5364 , 
    n5365 , 
    n5366 , 
    n5367 , 
    n5368 , 
    n5369 , 
    n5370 , 
    n5371 , 
    n5372 , 
    n5373 , 
    n5374 , 
    n5375 , 
    n5376 , 
    n5377 , 
    n5378 , 
    n5379 , 
    n5380 , 
    n5381 , 
    n5382 , 
    n5383 , 
    n5384 , 
    n5385 , 
    n5386 , 
    n5387 , 
    n5388 , 
    n5389 , 
    n5390 , 
    n5391 , 
    n5392 , 
    n5393 , 
    n5394 , 
    n5395 , 
    n5396 , 
    n5397 , 
    n5398 , 
    n5399 , 
    n5400 , 
    n5401 , 
    n5402 , 
    n5403 , 
    n5404 , 
    n5405 , 
    n5406 , 
    n5407 , 
    n5408 , 
    n5409 , 
    n5410 , 
    n5411 , 
    n5412 , 
    n5413 , 
    n5414 , 
    n5415 , 
    n5416 , 
    n5417 , 
    n5418 , 
    n5419 , 
    n5420 , 
    n5421 , 
    n5422 , 
    n5423 , 
    n5424 , 
    n5425 , 
    n5426 , 
    n5427 , 
    n5428 , 
    n5429 , 
    n5430 , 
    n5431 , 
    n5432 , 
    n5433 , 
    n5434 , 
    n5435 , 
    n5436 , 
    n5437 , 
    n5438 , 
    n5439 , 
    n5440 , 
    n5441 , 
    n5442 , 
    n5443 , 
    n5444 , 
    n5445 , 
    n5446 , 
    n5447 , 
    n5448 , 
    n5449 , 
    n5450 , 
    n5451 , 
    n5452 , 
    n5453 , 
    n5454 , 
    n5455 , 
    n5456 , 
    n5457 , 
    n5458 , 
    n5459 , 
    n5460 , 
    n5461 , 
    n5462 , 
    n5463 , 
    n5464 , 
    n5465 , 
    n5466 , 
    n5467 , 
    n5468 , 
    n5469 , 
    n5470 , 
    n5471 , 
    n5472 , 
    n5473 , 
    n5474 , 
    n5475 , 
    n5476 , 
    n5477 , 
    n5478 , 
    n5479 , 
    n5480 , 
    n5481 , 
    n5482 , 
    n5483 , 
    n5484 , 
    n5485 , 
    n5486 , 
    n5487 , 
    n5488 , 
    n5489 , 
    n5490 , 
    n5491 , 
    n5492 , 
    n5493 , 
    n5494 , 
    n5495 , 
    n5496 , 
    n5497 , 
    n5498 , 
    n5499 , 
    n5500 , 
    n5501 , 
    n5502 , 
    n5503 , 
    n5504 , 
    n5505 , 
    n5506 , 
    n5507 , 
    n5508 , 
    n5509 , 
    n5510 , 
    n5511 , 
    n5512 , 
    n5513 , 
    n5514 , 
    n5515 , 
    n5516 , 
    n5517 , 
    n5518 , 
    n5519 , 
    n5520 , 
    n5521 , 
    n5522 , 
    n5523 , 
    n5524 , 
    n5525 , 
    n5526 , 
    n5527 , 
    n5528 , 
    n5529 , 
    n5530 , 
    n5531 , 
    n5532 , 
    n5533 , 
    n5534 , 
    n5535 , 
    n5536 , 
    n5537 , 
    n5538 , 
    n5539 , 
    n5540 , 
    n5541 , 
    n5542 , 
    n5543 , 
    n5544 , 
    n5545 , 
    n5546 , 
    n5547 , 
    n5548 , 
    n5549 , 
    n5550 , 
    n5551 , 
    n5552 , 
    n5553 , 
    n5554 , 
    n5555 , 
    n5556 , 
    n5557 , 
    n5558 , 
    n5559 , 
    n5560 , 
    n5561 , 
    n5562 , 
    n5563 , 
    n5564 , 
    n5565 , 
    n5566 , 
    n5567 , 
    n5568 , 
    n5569 , 
    n5570 , 
    n5571 , 
    n5572 , 
    n5573 , 
    n5574 , 
    n5575 , 
    n5576 , 
    n5577 , 
    n5578 , 
    n5579 , 
    n5580 , 
    n5581 , 
    n5582 , 
    n5583 , 
    n5584 , 
    n5585 , 
    n5586 , 
    n5587 , 
    n5588 , 
    n5589 , 
    n5590 , 
    n5591 , 
    n5592 , 
    n5593 , 
    n5594 , 
    n5595 , 
    n5596 , 
    n5597 , 
    n5598 , 
    n5599 , 
    n5600 , 
    n5601 , 
    n5602 , 
    n5603 , 
    n5604 , 
    n5605 , 
    n5606 , 
    n5607 , 
    n5608 , 
    n5609 , 
    n5610 , 
    n5611 , 
    n5612 , 
    n5613 , 
    n5614 , 
    n5615 , 
    n5616 , 
    n5617 , 
    n5618 , 
    n5619 , 
    n5620 , 
    n5621 , 
    n5622 , 
    n5623 , 
    n5624 , 
    n5625 , 
    n5626 , 
    n5627 , 
    n5628 , 
    n5629 , 
    n5630 , 
    n5631 , 
    n5632 , 
    n5633 , 
    n5634 , 
    n5635 , 
    n5636 , 
    n5637 , 
    n5638 , 
    n5639 , 
    n5640 , 
    n5641 , 
    n5642 , 
    n5643 , 
    n5644 , 
    n5645 , 
    n5646 , 
    n5647 , 
    n5648 , 
    n5649 , 
    n5650 , 
    n5651 , 
    n5652 , 
    n5653 , 
    n5654 , 
    n5655 , 
    n5656 , 
    n5657 , 
    n5658 , 
    n5659 , 
    n5660 , 
    n5661 , 
    n5662 , 
    n5663 , 
    n5664 , 
    n5665 , 
    n5666 , 
    n5667 , 
    n5668 , 
    n5669 , 
    n5670 , 
    n5671 , 
    n5672 , 
    n5673 , 
    n5674 , 
    n5675 , 
    n5676 , 
    n5677 , 
    n5678 , 
    n5679 , 
    n5680 , 
    n5681 , 
    n5682 , 
    n5683 , 
    n5684 , 
    n5685 , 
    n5686 , 
    n5687 , 
    n5688 , 
    n5689 , 
    n5690 , 
    n5691 , 
    n5692 , 
    n5693 , 
    n5694 , 
    n5695 , 
    n5696 , 
    n5697 , 
    n5698 , 
    n5699 , 
    n5700 , 
    n5701 , 
    n5702 , 
    n5703 , 
    n5704 , 
    n5705 , 
    n5706 , 
    n5707 , 
    n5708 , 
    n5709 , 
    n5710 , 
    n5711 , 
    n5712 , 
    n5713 , 
    n5714 , 
    n5715 , 
    n5716 , 
    n5717 , 
    n5718 , 
    n5719 , 
    n5720 , 
    n5721 , 
    n5722 , 
    n5723 , 
    n5724 , 
    n5725 , 
    n5726 , 
    n5727 , 
    n5728 , 
    n5729 , 
    n5730 , 
    n5731 , 
    n5732 , 
    n5733 , 
    n5734 , 
    n5735 , 
    n5736 , 
    n5737 , 
    n5738 , 
    n5739 , 
    n5740 , 
    n5741 , 
    n5742 , 
    n5743 , 
    n5744 , 
    n5745 , 
    n5746 , 
    n5747 , 
    n5748 , 
    n5749 , 
    n5750 , 
    n5751 , 
    n5752 , 
    n5753 , 
    n5754 , 
    n5755 , 
    n5756 , 
    n5757 , 
    n5758 , 
    n5759 , 
    n5760 , 
    n5761 , 
    n5762 , 
    n5763 , 
    n5764 , 
    n5765 , 
    n5766 , 
    n5767 , 
    n5768 , 
    n5769 , 
    n5770 , 
    n5771 , 
    n5772 , 
    n5773 , 
    n5774 , 
    n5775 , 
    n5776 , 
    n5777 , 
    n5778 , 
    n5779 , 
    n5780 , 
    n5781 , 
    n5782 , 
    n5783 , 
    n5784 , 
    n5785 , 
    n5786 , 
    n5787 , 
    n5788 , 
    n5789 , 
    n5790 , 
    n5791 , 
    n5792 , 
    n5793 , 
    n5794 , 
    n5795 , 
    n5796 , 
    n5797 , 
    n5798 , 
    n5799 , 
    n5800 , 
    n5801 , 
    n5802 , 
    n5803 , 
    n5804 , 
    n5805 , 
    n5806 , 
    n5807 , 
    n5808 , 
    n5809 , 
    n5810 , 
    n5811 , 
    n5812 , 
    n5813 , 
    n5814 , 
    n5815 , 
    n5816 , 
    n5817 , 
    n5818 , 
    n5819 , 
    n5820 , 
    n5821 , 
    n5822 , 
    n5823 , 
    n5824 , 
    n5825 , 
    n5826 , 
    n5827 , 
    n5828 , 
    n5829 , 
    n5830 , 
    n5831 , 
    n5832 , 
    n5833 , 
    n5834 , 
    n5835 , 
    n5836 , 
    n5837 , 
    n5838 , 
    n5839 , 
    n5840 , 
    n5841 , 
    n5842 , 
    n5843 , 
    n5844 , 
    n5845 , 
    n5846 , 
    n5847 , 
    n5848 , 
    n5849 , 
    n5850 , 
    n5851 , 
    n5852 , 
    n5853 , 
    n5854 , 
    n5855 , 
    n5856 , 
    n5857 , 
    n5858 , 
    n5859 , 
    n5860 , 
    n5861 , 
    n5862 , 
    n5863 , 
    n5864 , 
    n5865 , 
    n5866 , 
    n5867 , 
    n5868 , 
    n5869 , 
    n5870 , 
    n5871 , 
    n5872 , 
    n5873 , 
    n5874 , 
    n5875 , 
    n5876 , 
    n5877 , 
    n5878 , 
    n5879 , 
    n5880 , 
    n5881 , 
    n5882 , 
    n5883 , 
    n5884 , 
    n5885 , 
    n5886 , 
    n5887 , 
    n5888 , 
    n5889 , 
    n5890 , 
    n5891 , 
    n5892 , 
    n5893 , 
    n5894 , 
    n5895 , 
    n5896 , 
    n5897 , 
    n5898 , 
    n5899 , 
    n5900 , 
    n5901 , 
    n5902 , 
    n5903 , 
    n5904 , 
    n5905 , 
    n5906 , 
    n5907 , 
    n5908 , 
    n5909 , 
    n5910 , 
    n5911 , 
    n5912 , 
    n5913 , 
    n5914 , 
    n5915 , 
    n5916 , 
    n5917 , 
    n5918 , 
    n5919 , 
    n5920 , 
    n5921 , 
    n5922 , 
    n5923 , 
    n5924 , 
    n5925 , 
    n5926 , 
    n5927 , 
    n5928 , 
    n5929 , 
    n5930 , 
    n5931 , 
    n5932 , 
    n5933 , 
    n5934 , 
    n5935 , 
    n5936 , 
    n5937 , 
    n5938 , 
    n5939 , 
    n5940 , 
    n5941 , 
    n5942 , 
    n5943 , 
    n5944 , 
    n5945 , 
    n5946 , 
    n5947 , 
    n5948 , 
    n5949 , 
    n5950 , 
    n5951 , 
    n5952 , 
    n5953 , 
    n5954 , 
    n5955 , 
    n5956 , 
    n5957 , 
    n5958 , 
    n5959 , 
    n5960 , 
    n5961 , 
    n5962 , 
    n5963 , 
    n5964 , 
    n5965 , 
    n5966 , 
    n5967 , 
    n5968 , 
    n5969 , 
    n5970 , 
    n5971 , 
    n5972 , 
    n5973 , 
    n5974 , 
    n5975 , 
    n5976 , 
    n5977 , 
    n5978 , 
    n5979 , 
    n5980 , 
    n5981 , 
    n5982 , 
    n5983 , 
    n5984 , 
    n5985 , 
    n5986 , 
    n5987 , 
    n5988 , 
    n5989 , 
    n5990 , 
    n5991 , 
    n5992 , 
    n5993 , 
    n5994 , 
    n5995 , 
    n5996 , 
    n5997 , 
    n5998 , 
    n5999 , 
    n6000 , 
    n6001 , 
    n6002 , 
    n6003 , 
    n6004 , 
    n6005 , 
    n6006 , 
    n6007 , 
    n6008 , 
    n6009 , 
    n6010 , 
    n6011 , 
    n6012 , 
    n6013 , 
    n6014 , 
    n6015 , 
    n6016 , 
    n6017 , 
    n6018 , 
    n6019 , 
    n6020 , 
    n6021 , 
    n6022 , 
    n6023 , 
    n6024 , 
    n6025 , 
    n6026 , 
    n6027 , 
    n6028 , 
    n6029 , 
    n6030 , 
    n6031 , 
    n6032 , 
    n6033 , 
    n6034 , 
    n6035 , 
    n6036 , 
    n6037 , 
    n6038 , 
    n6039 , 
    n6040 , 
    n6041 , 
    n6042 , 
    n6043 , 
    n6044 , 
    n6045 , 
    n6046 , 
    n6047 , 
    n6048 , 
    n6049 , 
    n6050 , 
    n6051 , 
    n6052 , 
    n6053 , 
    n6054 , 
    n6055 , 
    n6056 , 
    n6057 , 
    n6058 , 
    n6059 , 
    n6060 , 
    n6061 , 
    n6062 , 
    n6063 , 
    n6064 , 
    n6065 , 
    n6066 , 
    n6067 , 
    n6068 , 
    n6069 , 
    n6070 , 
    n6071 , 
    n6072 , 
    n6073 , 
    n6074 , 
    n6075 , 
    n6076 , 
    n6077 , 
    n6078 , 
    n6079 , 
    n6080 , 
    n6081 , 
    n6082 , 
    n6083 , 
    n6084 , 
    n6085 , 
    n6086 , 
    n6087 , 
    n6088 , 
    n6089 , 
    n6090 , 
    n6091 , 
    n6092 , 
    n6093 , 
    n6094 , 
    n6095 , 
    n6096 , 
    n6097 , 
    n6098 , 
    n6099 , 
    n6100 , 
    n6101 , 
    n6102 , 
    n6103 , 
    n6104 , 
    n6105 , 
    n6106 , 
    n6107 , 
    n6108 , 
    n6109 , 
    n6110 , 
    n6111 , 
    n6112 , 
    n6113 , 
    n6114 , 
    n6115 , 
    n6116 , 
    n6117 , 
    n6118 , 
    n6119 , 
    n6120 , 
    n6121 , 
    n6122 , 
    n6123 , 
    n6124 , 
    n6125 , 
    n6126 , 
    n6127 , 
    n6128 , 
    n6129 , 
    n6130 , 
    n6131 , 
    n6132 , 
    n6133 , 
    n6134 , 
    n6135 , 
    n6136 , 
    n6137 , 
    n6138 , 
    n6139 , 
    n6140 , 
    n6141 , 
    n6142 , 
    n6143 , 
    n6144 , 
    n6145 , 
    n6146 , 
    n6147 , 
    n6148 , 
    n6149 , 
    n6150 , 
    n6151 , 
    n6152 , 
    n6153 , 
    n6154 , 
    n6155 , 
    n6156 , 
    n6157 , 
    n6158 , 
    n6159 , 
    n6160 , 
    n6161 , 
    n6162 , 
    n6163 , 
    n6164 , 
    n6165 , 
    n6166 , 
    n6167 , 
    n6168 , 
    n6169 , 
    n6170 , 
    n6171 , 
    n6172 , 
    n6173 , 
    n6174 , 
    n6175 , 
    n6176 , 
    n6177 , 
    n6178 , 
    n6179 , 
    n6180 , 
    n6181 , 
    n6182 , 
    n6183 , 
    n6184 , 
    n6185 , 
    n6186 , 
    n6187 , 
    n6188 , 
    n6189 , 
    n6190 , 
    n6191 , 
    n6192 , 
    n6193 , 
    n6194 , 
    n6195 , 
    n6196 , 
    n6197 , 
    n6198 , 
    n6199 , 
    n6200 , 
    n6201 , 
    n6202 , 
    n6203 , 
    n6204 , 
    n6205 , 
    n6206 , 
    n6207 , 
    n6208 , 
    n6209 , 
    n6210 , 
    n6211 , 
    n6212 , 
    n6213 , 
    n6214 , 
    n6215 , 
    n6216 , 
    n6217 , 
    n6218 , 
    n6219 , 
    n6220 , 
    n6221 , 
    n6222 , 
    n6223 , 
    n6224 , 
    n6225 , 
    n6226 , 
    n6227 , 
    n6228 , 
    n6229 , 
    n6230 , 
    n6231 , 
    n6232 , 
    n6233 , 
    n6234 , 
    n6235 , 
    n6236 , 
    n6237 , 
    n6238 , 
    n6239 , 
    n6240 , 
    n6241 , 
    n6242 , 
    n6243 , 
    n6244 , 
    n6245 , 
    n6246 , 
    n6247 , 
    n6248 , 
    n6249 , 
    n6250 , 
    n6251 , 
    n6252 , 
    n6253 , 
    n6254 , 
    n6255 , 
    n6256 , 
    n6257 , 
    n6258 , 
    n6259 , 
    n6260 , 
    n6261 , 
    n6262 , 
    n6263 , 
    n6264 , 
    n6265 , 
    n6266 , 
    n6267 , 
    n6268 , 
    n6269 , 
    n6270 , 
    n6271 , 
    n6272 , 
    n6273 , 
    n6274 , 
    n6275 , 
    n6276 , 
    n6277 , 
    n6278 , 
    n6279 , 
    n6280 , 
    n6281 , 
    n6282 , 
    n6283 , 
    n6284 , 
    n6285 , 
    n6286 , 
    n6287 , 
    n6288 , 
    n6289 , 
    n6290 , 
    n6291 , 
    n6292 , 
    n6293 , 
    n6294 , 
    n6295 , 
    n6296 , 
    n6297 , 
    n6298 , 
    n6299 , 
    n6300 , 
    n6301 , 
    n6302 , 
    n6303 , 
    n6304 , 
    n6305 , 
    n6306 , 
    n6307 , 
    n6308 , 
    n6309 , 
    n6310 , 
    n6311 , 
    n6312 , 
    n6313 , 
    n6314 , 
    n6315 , 
    n6316 , 
    n6317 , 
    n6318 , 
    n6319 , 
    n6320 , 
    n6321 , 
    n6322 , 
    n6323 , 
    n6324 , 
    n6325 , 
    n6326 , 
    n6327 , 
    n6328 , 
    n6329 , 
    n6330 , 
    n6331 , 
    n6332 , 
    n6333 , 
    n6334 , 
    n6335 , 
    n6336 , 
    n6337 , 
    n6338 , 
    n6339 , 
    n6340 , 
    n6341 , 
    n6342 , 
    n6343 , 
    n6344 , 
    n6345 , 
    n6346 , 
    n6347 , 
    n6348 , 
    n6349 , 
    n6350 , 
    n6351 , 
    n6352 , 
    n6353 , 
    n6354 , 
    n6355 , 
    n6356 , 
    n6357 , 
    n6358 , 
    n6359 , 
    n6360 , 
    n6361 , 
    n6362 , 
    n6363 , 
    n6364 , 
    n6365 , 
    n6366 , 
    n6367 , 
    n6368 , 
    n6369 , 
    n6370 , 
    n6371 , 
    n6372 , 
    n6373 , 
    n6374 , 
    n6375 , 
    n6376 , 
    n6377 , 
    n6378 , 
    n6379 , 
    n6380 , 
    n6381 , 
    n6382 , 
    n6383 , 
    n6384 , 
    n6385 , 
    n6386 , 
    n6387 , 
    n6388 , 
    n6389 , 
    n6390 , 
    n6391 , 
    n6392 , 
    n6393 , 
    n6394 , 
    n6395 , 
    n6396 , 
    n6397 , 
    n6398 , 
    n6399 , 
    n6400 , 
    n6401 , 
    n6402 , 
    n6403 , 
    n6404 , 
    n6405 , 
    n6406 , 
    n6407 , 
    n6408 , 
    n6409 , 
    n6410 , 
    n6411 , 
    n6412 , 
    n6413 , 
    n6414 , 
    n6415 , 
    n6416 , 
    n6417 , 
    n6418 , 
    n6419 , 
    n6420 , 
    n6421 , 
    n6422 , 
    n6423 , 
    n6424 , 
    n6425 , 
    n6426 , 
    n6427 , 
    n6428 , 
    n6429 , 
    n6430 , 
    n6431 , 
    n6432 , 
    n6433 , 
    n6434 , 
    n6435 , 
    n6436 , 
    n6437 , 
    n6438 , 
    n6439 , 
    n6440 , 
    n6441 , 
    n6442 , 
    n6443 , 
    n6444 , 
    n6445 , 
    n6446 , 
    n6447 , 
    n6448 , 
    n6449 , 
    n6450 , 
    n6451 , 
    n6452 , 
    n6453 , 
    n6454 , 
    n6455 , 
    n6456 , 
    n6457 , 
    n6458 , 
    n6459 , 
    n6460 , 
    n6461 , 
    n6462 , 
    n6463 , 
    n6464 , 
    n6465 , 
    n6466 , 
    n6467 , 
    n6468 , 
    n6469 , 
    n6470 , 
    n6471 , 
    n6472 , 
    n6473 , 
    n6474 , 
    n6475 , 
    n6476 , 
    n6477 , 
    n6478 , 
    n6479 , 
    n6480 , 
    n6481 , 
    n6482 , 
    n6483 , 
    n6484 , 
    n6485 , 
    n6486 , 
    n6487 , 
    n6488 , 
    n6489 , 
    n6490 , 
    n6491 , 
    n6492 , 
    n6493 , 
    n6494 , 
    n6495 , 
    n6496 , 
    n6497 , 
    n6498 , 
    n6499 , 
    n6500 , 
    n6501 , 
    n6502 , 
    n6503 , 
    n6504 , 
    n6505 , 
    n6506 , 
    n6507 , 
    n6508 , 
    n6509 , 
    n6510 , 
    n6511 , 
    n6512 , 
    n6513 , 
    n6514 , 
    n6515 , 
    n6516 , 
    n6517 , 
    n6518 , 
    n6519 , 
    n6520 , 
    n6521 , 
    n6522 , 
    n6523 , 
    n6524 , 
    n6525 , 
    n6526 , 
    n6527 , 
    n6528 , 
    n6529 , 
    n6530 , 
    n6531 , 
    n6532 , 
    n6533 , 
    n6534 , 
    n6535 , 
    n6536 , 
    n6537 , 
    n6538 , 
    n6539 , 
    n6540 , 
    n6541 , 
    n6542 , 
    n6543 , 
    n6544 , 
    n6545 , 
    n6546 , 
    n6547 , 
    n6548 , 
    n6549 , 
    n6550 , 
    n6551 , 
    n6552 , 
    n6553 , 
    n6554 , 
    n6555 , 
    n6556 , 
    n6557 , 
    n6558 , 
    n6559 , 
    n6560 , 
    n6561 , 
    n6562 , 
    n6563 , 
    n6564 , 
    n6565 , 
    n6566 , 
    n6567 , 
    n6568 , 
    n6569 , 
    n6570 , 
    n6571 , 
    n6572 , 
    n6573 , 
    n6574 , 
    n6575 , 
    n6576 , 
    n6577 , 
    n6578 , 
    n6579 , 
    n6580 , 
    n6581 , 
    n6582 , 
    n6583 , 
    n6584 , 
    n6585 , 
    n6586 , 
    n6587 , 
    n6588 , 
    n6589 , 
    n6590 , 
    n6591 , 
    n6592 , 
    n6593 , 
    n6594 , 
    n6595 , 
    n6596 , 
    n6597 , 
    n6598 , 
    n6599 , 
    n6600 , 
    n6601 , 
    n6602 , 
    n6603 , 
    n6604 , 
    n6605 , 
    n6606 , 
    n6607 , 
    n6608 , 
    n6609 , 
    n6610 , 
    n6611 , 
    n6612 , 
    n6613 , 
    n6614 , 
    n6615 , 
    n6616 , 
    n6617 , 
    n6618 , 
    n6619 , 
    n6620 , 
    n6621 , 
    n6622 , 
    n6623 , 
    n6624 , 
    n6625 , 
    n6626 , 
    n6627 , 
    n6628 , 
    n6629 , 
    n6630 , 
    n6631 , 
    n6632 , 
    n6633 , 
    n6634 , 
    n6635 , 
    n6636 , 
    n6637 , 
    n6638 , 
    n6639 , 
    n6640 , 
    n6641 , 
    n6642 , 
    n6643 , 
    n6644 , 
    n6645 , 
    n6646 , 
    n6647 , 
    n6648 , 
    n6649 , 
    n6650 , 
    n6651 , 
    n6652 , 
    n6653 , 
    n6654 , 
    n6655 , 
    n6656 , 
    n6657 , 
    n6658 , 
    n6659 , 
    n6660 , 
    n6661 , 
    n6662 , 
    n6663 , 
    n6664 , 
    n6665 , 
    n6666 , 
    n6667 , 
    n6668 , 
    n6669 , 
    n6670 , 
    n6671 , 
    n6672 , 
    n6673 , 
    n6674 , 
    n6675 , 
    n6676 , 
    n6677 , 
    n6678 , 
    n6679 , 
    n6680 , 
    n6681 , 
    n6682 , 
    n6683 , 
    n6684 , 
    n6685 , 
    n6686 , 
    n6687 , 
    n6688 , 
    n6689 , 
    n6690 , 
    n6691 , 
    n6692 , 
    n6693 , 
    n6694 , 
    n6695 , 
    n6696 , 
    n6697 , 
    n6698 , 
    n6699 , 
    n6700 , 
    n6701 , 
    n6702 , 
    n6703 , 
    n6704 , 
    n6705 , 
    n6706 , 
    n6707 , 
    n6708 , 
    n6709 , 
    n6710 , 
    n6711 , 
    n6712 , 
    n6713 , 
    n6714 , 
    n6715 , 
    n6716 , 
    n6717 , 
    n6718 , 
    n6719 , 
    n6720 , 
    n6721 , 
    n6722 , 
    n6723 , 
    n6724 , 
    n6725 , 
    n6726 , 
    n6727 , 
    n6728 , 
    n6729 , 
    n6730 , 
    n6731 , 
    n6732 , 
    n6733 , 
    n6734 , 
    n6735 , 
    n6736 , 
    n6737 , 
    n6738 , 
    n6739 , 
    n6740 , 
    n6741 , 
    n6742 , 
    n6743 , 
    n6744 , 
    n6745 , 
    n6746 , 
    n6747 , 
    n6748 , 
    n6749 , 
    n6750 , 
    n6751 , 
    n6752 , 
    n6753 , 
    n6754 , 
    n6755 , 
    n6756 , 
    n6757 , 
    n6758 , 
    n6759 , 
    n6760 );
input 
    n0 , 
    n1 , 
    n2 , 
    n3 , 
    n4 , 
    n5 , 
    n6 , 
    n7 , 
    n8 , 
    n9 , 
    n10 , 
    n11 , 
    n12 , 
    n13 , 
    n14 , 
    n15 , 
    n16 , 
    n17 , 
    n18 , 
    n19 , 
    n20 , 
    n21 , 
    n22 , 
    n23 , 
    n24 , 
    n25 , 
    n26 , 
    n27 , 
    n28 , 
    n29 , 
    n30 , 
    n31 , 
    n32 , 
    n33 , 
    n34 , 
    n35 , 
    n36 , 
    n37 , 
    n38 , 
    n39 , 
    n40 , 
    n41 , 
    n42 , 
    n43 , 
    n44 , 
    n45 , 
    n46 , 
    n47 , 
    n48 , 
    n49 , 
    n50 , 
    n51 , 
    n52 , 
    n53 , 
    n54 , 
    n55 , 
    n56 , 
    n57 , 
    n58 , 
    n59 , 
    n60 , 
    n61 , 
    n62 , 
    n63 , 
    n64 , 
    n65 , 
    n66 , 
    n67 , 
    n68 , 
    n69 , 
    n70 , 
    n71 , 
    n72 , 
    n73 , 
    n74 , 
    n75 , 
    n76 , 
    n77 , 
    n78 , 
    n79 , 
    n80 , 
    n81 , 
    n82 , 
    n83 , 
    n84 , 
    n85 , 
    n86 , 
    n87 , 
    n88 , 
    n89 , 
    n90 , 
    n91 , 
    n92 , 
    n93 , 
    n94 , 
    n95 , 
    n96 , 
    n97 , 
    n98 , 
    n99 , 
    n100 , 
    n101 , 
    n102 , 
    n103 , 
    n104 , 
    n105 , 
    n106 , 
    n107 , 
    n108 , 
    n109 , 
    n110 , 
    n111 , 
    n112 , 
    n113 , 
    n114 , 
    n115 , 
    n116 , 
    n117 , 
    n118 , 
    n119 , 
    n120 , 
    n121 , 
    n122 , 
    n123 , 
    n124 , 
    n125 , 
    n126 , 
    n127 , 
    n128 , 
    n129 , 
    n130 , 
    n131 , 
    n132 , 
    n133 , 
    n134 , 
    n135 , 
    n136 , 
    n137 , 
    n138 , 
    n139 , 
    n140 , 
    n141 , 
    n142 , 
    n143 , 
    n144 , 
    n145 , 
    n146 , 
    n147 , 
    n148 , 
    n149 , 
    n150 , 
    n151 , 
    n152 , 
    n153 , 
    n154 , 
    n155 , 
    n156 , 
    n157 , 
    n158 , 
    n159 , 
    n160 , 
    n161 , 
    n162 , 
    n163 , 
    n164 , 
    n165 , 
    n166 , 
    n167 , 
    n168 , 
    n169 , 
    n170 , 
    n171 , 
    n172 , 
    n173 , 
    n174 , 
    n175 , 
    n176 , 
    n177 , 
    n178 , 
    n179 , 
    n180 , 
    n181 , 
    n182 , 
    n183 , 
    n184 , 
    n185 , 
    n186 , 
    n187 , 
    n188 , 
    n189 , 
    n190 , 
    n191 , 
    n192 , 
    n193 , 
    n194 , 
    n195 , 
    n196 , 
    n197 , 
    n198 , 
    n199 , 
    n200 , 
    n201 , 
    n202 , 
    n203 , 
    n204 , 
    n205 , 
    n206 , 
    n207 , 
    n208 , 
    n209 , 
    n210 , 
    n211 , 
    n212 , 
    n213 , 
    n214 , 
    n215 , 
    n216 , 
    n217 , 
    n218 , 
    n219 , 
    n220 , 
    n221 , 
    n222 , 
    n223 , 
    n224 , 
    n225 , 
    n226 , 
    n227 , 
    n228 , 
    n229 , 
    n230 , 
    n231 , 
    n232 , 
    n233 , 
    n234 , 
    n235 , 
    n236 , 
    n237 , 
    n238 , 
    n239 , 
    n240 , 
    n241 , 
    n242 , 
    n243 , 
    n244 , 
    n245 , 
    n246 , 
    n247 , 
    n248 , 
    n249 , 
    n250 , 
    n251 , 
    n252 , 
    n253 , 
    n254 , 
    n255 , 
    n256 , 
    n257 , 
    n258 , 
    n259 , 
    n260 , 
    n261 , 
    n262 , 
    n263 , 
    n264 , 
    n265 , 
    n266 , 
    n267 , 
    n268 , 
    n269 , 
    n270 , 
    n271 , 
    n272 , 
    n273 , 
    n274 , 
    n275 , 
    n276 , 
    n277 , 
    n278 , 
    n279 , 
    n280 , 
    n281 , 
    n282 , 
    n283 , 
    n284 , 
    n285 , 
    n286 , 
    n287 , 
    n288 , 
    n289 , 
    n290 , 
    n291 , 
    n292 , 
    n293 , 
    n294 , 
    n295 , 
    n296 , 
    n297 , 
    n298 , 
    n299 , 
    n300 , 
    n301 , 
    n302 , 
    n303 , 
    n304 , 
    n305 , 
    n306 , 
    n307 , 
    n308 , 
    n309 , 
    n310 , 
    n311 , 
    n312 , 
    n313 , 
    n314 , 
    n315 , 
    n316 , 
    n317 , 
    n318 , 
    n319 , 
    n320 , 
    n321 , 
    n322 , 
    n323 , 
    n324 , 
    n325 , 
    n326 , 
    n327 , 
    n328 , 
    n329 , 
    n330 , 
    n331 , 
    n332 , 
    n333 , 
    n334 , 
    n335 , 
    n336 , 
    n337 , 
    n338 , 
    n339 , 
    n340 , 
    n341 , 
    n342 , 
    n343 , 
    n344 , 
    n345 , 
    n346 , 
    n347 , 
    n348 , 
    n349 , 
    n350 , 
    n351 , 
    n352 , 
    n353 , 
    n354 , 
    n355 , 
    n356 , 
    n357 , 
    n358 , 
    n359 , 
    n360 , 
    n361 , 
    n362 , 
    n363 , 
    n364 , 
    n365 , 
    n366 , 
    n367 , 
    n368 , 
    n369 , 
    n370 , 
    n371 , 
    n372 , 
    n373 , 
    n374 , 
    n375 , 
    n376 , 
    n377 , 
    n378 , 
    n379 , 
    n380 , 
    n381 , 
    n382 , 
    n383 , 
    n384 , 
    n385 , 
    n386 , 
    n387 , 
    n388 , 
    n389 , 
    n390 , 
    n391 , 
    n392 , 
    n393 , 
    n394 , 
    n395 , 
    n396 , 
    n397 , 
    n398 , 
    n399 , 
    n400 , 
    n401 , 
    n402 , 
    n403 , 
    n404 , 
    n405 , 
    n406 , 
    n407 , 
    n408 , 
    n409 , 
    n410 , 
    n411 , 
    n412 , 
    n413 , 
    n414 , 
    n415 , 
    n416 , 
    n417 , 
    n418 , 
    n419 , 
    n420 , 
    n421 , 
    n422 , 
    n423 , 
    n424 , 
    n425 , 
    n426 , 
    n427 , 
    n428 , 
    n429 , 
    n430 , 
    n431 , 
    n432 , 
    n433 , 
    n434 , 
    n435 , 
    n436 , 
    n437 , 
    n438 , 
    n439 , 
    n440 , 
    n441 , 
    n442 , 
    n443 , 
    n444 , 
    n445 , 
    n446 , 
    n447 , 
    n448 , 
    n449 , 
    n450 , 
    n451 , 
    n452 , 
    n453 , 
    n454 , 
    n455 , 
    n456 , 
    n457 , 
    n458 , 
    n459 , 
    n460 , 
    n461 , 
    n462 , 
    n463 , 
    n464 , 
    n465 , 
    n466 , 
    n467 , 
    n468 , 
    n469 , 
    n470 , 
    n471 , 
    n472 , 
    n473 , 
    n474 , 
    n475 , 
    n476 , 
    n477 , 
    n478 , 
    n479 , 
    n480 , 
    n481 , 
    n482 , 
    n483 , 
    n484 , 
    n485 , 
    n486 , 
    n487 , 
    n488 , 
    n489 , 
    n490 , 
    n491 , 
    n492 , 
    n493 , 
    n494 , 
    n495 , 
    n496 , 
    n497 , 
    n498 , 
    n499 , 
    n500 , 
    n501 , 
    n502 , 
    n503 , 
    n504 , 
    n505 , 
    n506 , 
    n507 , 
    n508 , 
    n509 , 
    n510 , 
    n511 , 
    n512 , 
    n513 , 
    n514 , 
    n515 , 
    n516 , 
    n517 , 
    n518 , 
    n519 , 
    n520 , 
    n521 , 
    n522 , 
    n523 , 
    n524 , 
    n525 , 
    n526 , 
    n527 , 
    n528 , 
    n529 , 
    n530 , 
    n531 , 
    n532 , 
    n533 , 
    n534 , 
    n535 , 
    n536 , 
    n537 , 
    n538 , 
    n539 , 
    n540 , 
    n541 , 
    n542 , 
    n543 , 
    n544 , 
    n545 , 
    n546 , 
    n547 , 
    n548 , 
    n549 , 
    n550 , 
    n551 , 
    n552 , 
    n553 , 
    n554 , 
    n555 , 
    n556 , 
    n557 , 
    n558 , 
    n559 , 
    n560 , 
    n561 , 
    n562 , 
    n563 , 
    n564 , 
    n565 , 
    n566 , 
    n567 , 
    n568 , 
    n569 , 
    n570 , 
    n571 , 
    n572 , 
    n573 , 
    n574 , 
    n575 , 
    n576 , 
    n577 , 
    n578 , 
    n579 , 
    n580 , 
    n581 , 
    n582 , 
    n583 , 
    n584 , 
    n585 , 
    n586 , 
    n587 , 
    n588 , 
    n589 , 
    n590 , 
    n591 , 
    n592 , 
    n593 , 
    n594 , 
    n595 , 
    n596 , 
    n597 , 
    n598 , 
    n599 , 
    n600 , 
    n601 , 
    n602 , 
    n603 , 
    n604 , 
    n605 , 
    n606 , 
    n607 , 
    n608 , 
    n609 , 
    n610 , 
    n611 , 
    n612 , 
    n613 , 
    n614 , 
    n615 , 
    n616 , 
    n617 , 
    n618 , 
    n619 , 
    n620 , 
    n621 , 
    n622 , 
    n623 , 
    n624 , 
    n625 , 
    n626 , 
    n627 , 
    n628 , 
    n629 , 
    n630 , 
    n631 , 
    n632 , 
    n633 , 
    n634 , 
    n635 , 
    n636 , 
    n637 , 
    n638 , 
    n639 , 
    n640 , 
    n641 , 
    n642 , 
    n643 , 
    n644 , 
    n645 , 
    n646 , 
    n647 , 
    n648 , 
    n649 , 
    n650 , 
    n651 , 
    n652 , 
    n653 , 
    n654 , 
    n655 , 
    n656 , 
    n657 , 
    n658 , 
    n659 , 
    n660 , 
    n661 , 
    n662 , 
    n663 , 
    n664 , 
    n665 , 
    n666 , 
    n667 , 
    n668 , 
    n669 , 
    n670 , 
    n671 , 
    n672 , 
    n673 , 
    n674 , 
    n675 , 
    n676 , 
    n677 , 
    n678 , 
    n679 , 
    n680 , 
    n681 , 
    n682 , 
    n683 , 
    n684 , 
    n685 , 
    n686 , 
    n687 , 
    n688 , 
    n689 , 
    n690 , 
    n691 , 
    n692 , 
    n693 , 
    n694 , 
    n695 , 
    n696 , 
    n697 , 
    n698 , 
    n699 , 
    n700 , 
    n701 , 
    n702 , 
    n703 , 
    n704 , 
    n705 , 
    n706 , 
    n707 , 
    n708 , 
    n709 , 
    n710 , 
    n711 , 
    n712 , 
    n713 , 
    n714 , 
    n715 , 
    n716 , 
    n717 , 
    n718 , 
    n719 , 
    n720 , 
    n721 , 
    n722 , 
    n723 , 
    n724 , 
    n725 , 
    n726 , 
    n727 , 
    n728 , 
    n729 , 
    n730 , 
    n731 , 
    n732 , 
    n733 , 
    n734 , 
    n735 , 
    n736 , 
    n737 , 
    n738 , 
    n739 , 
    n740 , 
    n741 , 
    n742 , 
    n743 , 
    n744 , 
    n745 , 
    n746 , 
    n747 , 
    n748 , 
    n749 , 
    n750 , 
    n751 , 
    n752 , 
    n753 , 
    n754 , 
    n755 , 
    n756 , 
    n757 , 
    n758 , 
    n759 , 
    n760 , 
    n761 , 
    n762 , 
    n763 , 
    n764 , 
    n765 , 
    n766 , 
    n767 , 
    n768 , 
    n769 , 
    n770 , 
    n771 , 
    n772 , 
    n773 , 
    n774 , 
    n775 , 
    n776 , 
    n777 , 
    n778 , 
    n779 , 
    n780 , 
    n781 , 
    n782 , 
    n783 , 
    n784 , 
    n785 , 
    n786 , 
    n787 , 
    n788 , 
    n789 , 
    n790 , 
    n791 , 
    n792 , 
    n793 , 
    n794 , 
    n795 , 
    n796 , 
    n797 , 
    n798 , 
    n799 , 
    n800 , 
    n801 , 
    n802 , 
    n803 , 
    n804 , 
    n805 , 
    n806 , 
    n807 , 
    n808 , 
    n809 , 
    n810 , 
    n811 , 
    n812 , 
    n813 , 
    n814 , 
    n815 , 
    n816 , 
    n817 , 
    n818 , 
    n819 , 
    n820 , 
    n821 , 
    n822 , 
    n823 , 
    n824 , 
    n825 , 
    n826 , 
    n827 , 
    n828 , 
    n829 , 
    n830 , 
    n831 , 
    n832 , 
    n833 , 
    n834 , 
    n835 , 
    n836 , 
    n837 , 
    n838 , 
    n839 , 
    n840 , 
    n841 , 
    n842 , 
    n843 , 
    n844 , 
    n845 , 
    n846 , 
    n847 , 
    n848 , 
    n849 , 
    n850 , 
    n851 , 
    n852 , 
    n853 , 
    n854 , 
    n855 , 
    n856 , 
    n857 , 
    n858 , 
    n859 , 
    n860 , 
    n861 , 
    n862 , 
    n863 , 
    n864 , 
    n865 , 
    n866 , 
    n867 , 
    n868 , 
    n869 , 
    n870 , 
    n871 , 
    n872 , 
    n873 , 
    n874 , 
    n875 , 
    n876 , 
    n877 , 
    n878 , 
    n879 , 
    n880 , 
    n881 , 
    n882 , 
    n883 , 
    n884 , 
    n885 , 
    n886 , 
    n887 , 
    n888 , 
    n889 , 
    n890 , 
    n891 , 
    n892 , 
    n893 , 
    n894 , 
    n895 , 
    n896 , 
    n897 , 
    n898 , 
    n899 , 
    n900 , 
    n901 , 
    n902 , 
    n903 , 
    n904 , 
    n905 , 
    n906 , 
    n907 , 
    n908 , 
    n909 , 
    n910 , 
    n911 , 
    n912 , 
    n913 , 
    n914 , 
    n915 , 
    n916 , 
    n917 , 
    n918 , 
    n919 , 
    n920 , 
    n921 , 
    n922 , 
    n923 , 
    n924 , 
    n925 , 
    n926 , 
    n927 , 
    n928 , 
    n929 , 
    n930 , 
    n931 , 
    n932 , 
    n933 , 
    n934 , 
    n935 , 
    n936 , 
    n937 , 
    n938 , 
    n939 , 
    n940 , 
    n941 , 
    n942 , 
    n943 , 
    n944 , 
    n945 , 
    n946 , 
    n947 , 
    n948 , 
    n949 , 
    n950 , 
    n951 , 
    n952 , 
    n953 , 
    n954 , 
    n955 , 
    n956 , 
    n957 , 
    n958 , 
    n959 , 
    n960 , 
    n961 , 
    n962 , 
    n963 , 
    n964 , 
    n965 , 
    n966 , 
    n967 , 
    n968 , 
    n969 , 
    n970 , 
    n971 , 
    n972 , 
    n973 , 
    n974 , 
    n975 , 
    n976 , 
    n977 , 
    n978 , 
    n979 , 
    n980 , 
    n981 , 
    n982 , 
    n983 , 
    n984 , 
    n985 , 
    n986 , 
    n987 , 
    n988 , 
    n989 , 
    n990 , 
    n991 , 
    n992 , 
    n993 , 
    n994 , 
    n995 , 
    n996 , 
    n997 , 
    n998 , 
    n999 , 
    n1000 , 
    n1001 , 
    n1002 , 
    n1003 , 
    n1004 , 
    n1005 , 
    n1006 , 
    n1007 , 
    n1008 , 
    n1009 , 
    n1010 , 
    n1011 , 
    n1012 , 
    n1013 , 
    n1014 , 
    n1015 , 
    n1016 , 
    n1017 , 
    n1018 , 
    n1019 , 
    n1020 , 
    n1021 , 
    n1022 , 
    n1023 , 
    n1024 , 
    n1025 , 
    n1026 , 
    n1027 , 
    n1028 , 
    n1029 , 
    n1030 , 
    n1031 , 
    n1032 , 
    n1033 , 
    n1034 , 
    n1035 , 
    n1036 , 
    n1037 , 
    n1038 , 
    n1039 , 
    n1040 , 
    n1041 , 
    n1042 , 
    n1043 , 
    n1044 , 
    n1045 , 
    n1046 , 
    n1047 , 
    n1048 , 
    n1049 , 
    n1050 , 
    n1051 , 
    n1052 , 
    n1053 , 
    n1054 , 
    n1055 , 
    n1056 , 
    n1057 , 
    n1058 , 
    n1059 , 
    n1060 , 
    n1061 , 
    n1062 , 
    n1063 , 
    n1064 , 
    n1065 , 
    n1066 , 
    n1067 , 
    n1068 , 
    n1069 , 
    n1070 , 
    n1071 , 
    n1072 , 
    n1073 , 
    n1074 , 
    n1075 , 
    n1076 , 
    n1077 , 
    n1078 , 
    n1079 , 
    n1080 , 
    n1081 , 
    n1082 , 
    n1083 , 
    n1084 , 
    n1085 , 
    n1086 , 
    n1087 , 
    n1088 , 
    n1089 , 
    n1090 , 
    n1091 , 
    n1092 , 
    n1093 , 
    n1094 , 
    n1095 , 
    n1096 , 
    n1097 , 
    n1098 , 
    n1099 , 
    n1100 , 
    n1101 , 
    n1102 , 
    n1103 , 
    n1104 , 
    n1105 , 
    n1106 , 
    n1107 , 
    n1108 , 
    n1109 , 
    n1110 , 
    n1111 , 
    n1112 , 
    n1113 , 
    n1114 , 
    n1115 , 
    n1116 , 
    n1117 , 
    n1118 , 
    n1119 , 
    n1120 , 
    n1121 , 
    n1122 , 
    n1123 , 
    n1124 , 
    n1125 , 
    n1126 , 
    n1127 , 
    n1128 , 
    n1129 , 
    n1130 , 
    n1131 , 
    n1132 , 
    n1133 , 
    n1134 , 
    n1135 , 
    n1136 , 
    n1137 , 
    n1138 , 
    n1139 , 
    n1140 , 
    n1141 , 
    n1142 , 
    n1143 , 
    n1144 , 
    n1145 , 
    n1146 , 
    n1147 , 
    n1148 , 
    n1149 , 
    n1150 , 
    n1151 , 
    n1152 , 
    n1153 , 
    n1154 , 
    n1155 , 
    n1156 , 
    n1157 , 
    n1158 , 
    n1159 , 
    n1160 , 
    n1161 , 
    n1162 , 
    n1163 , 
    n1164 , 
    n1165 , 
    n1166 , 
    n1167 , 
    n1168 , 
    n1169 , 
    n1170 , 
    n1171 , 
    n1172 , 
    n1173 , 
    n1174 , 
    n1175 , 
    n1176 , 
    n1177 , 
    n1178 , 
    n1179 , 
    n1180 , 
    n1181 , 
    n1182 , 
    n1183 , 
    n1184 , 
    n1185 , 
    n1186 , 
    n1187 , 
    n1188 , 
    n1189 , 
    n1190 , 
    n1191 , 
    n1192 , 
    n1193 , 
    n1194 , 
    n1195 , 
    n1196 , 
    n1197 , 
    n1198 , 
    n1199 , 
    n1200 , 
    n1201 , 
    n1202 , 
    n1203 , 
    n1204 , 
    n1205 , 
    n1206 , 
    n1207 , 
    n1208 , 
    n1209 , 
    n1210 , 
    n1211 , 
    n1212 , 
    n1213 , 
    n1214 , 
    n1215 , 
    n1216 , 
    n1217 , 
    n1218 , 
    n1219 , 
    n1220 , 
    n1221 , 
    n1222 , 
    n1223 , 
    n1224 , 
    n1225 , 
    n1226 , 
    n1227 , 
    n1228 , 
    n1229 , 
    n1230 , 
    n1231 , 
    n1232 , 
    n1233 , 
    n1234 , 
    n1235 , 
    n1236 , 
    n1237 , 
    n1238 , 
    n1239 , 
    n1240 , 
    n1241 , 
    n1242 , 
    n1243 , 
    n1244 , 
    n1245 , 
    n1246 , 
    n1247 , 
    n1248 , 
    n1249 , 
    n1250 , 
    n1251 , 
    n1252 , 
    n1253 , 
    n1254 , 
    n1255 , 
    n1256 , 
    n1257 , 
    n1258 , 
    n1259 , 
    n1260 , 
    n1261 , 
    n1262 , 
    n1263 , 
    n1264 , 
    n1265 , 
    n1266 , 
    n1267 , 
    n1268 , 
    n1269 , 
    n1270 , 
    n1271 , 
    n1272 , 
    n1273 , 
    n1274 , 
    n1275 , 
    n1276 , 
    n1277 , 
    n1278 , 
    n1279 , 
    n1280 , 
    n1281 , 
    n1282 , 
    n1283 , 
    n1284 , 
    n1285 , 
    n1286 , 
    n1287 , 
    n1288 , 
    n1289 , 
    n1290 , 
    n1291 , 
    n1292 , 
    n1293 , 
    n1294 , 
    n1295 , 
    n1296 , 
    n1297 , 
    n1298 , 
    n1299 , 
    n1300 , 
    n1301 , 
    n1302 , 
    n1303 , 
    n1304 , 
    n1305 , 
    n1306 , 
    n1307 , 
    n1308 , 
    n1309 , 
    n1310 , 
    n1311 , 
    n1312 , 
    n1313 , 
    n1314 , 
    n1315 , 
    n1316 , 
    n1317 , 
    n1318 , 
    n1319 , 
    n1320 , 
    n1321 , 
    n1322 , 
    n1323 , 
    n1324 , 
    n1325 , 
    n1326 , 
    n1327 , 
    n1328 , 
    n1329 , 
    n1330 , 
    n1331 , 
    n1332 , 
    n1333 , 
    n1334 , 
    n1335 , 
    n1336 , 
    n1337 , 
    n1338 , 
    n1339 , 
    n1340 , 
    n1341 , 
    n1342 , 
    n1343 , 
    n1344 , 
    n1345 , 
    n1346 , 
    n1347 , 
    n1348 , 
    n1349 , 
    n1350 , 
    n1351 , 
    n1352 , 
    n1353 , 
    n1354 , 
    n1355 , 
    n1356 , 
    n1357 , 
    n1358 , 
    n1359 , 
    n1360 , 
    n1361 , 
    n1362 , 
    n1363 ;
output 
    n1364 , 
    n1365 , 
    n1366 , 
    n1367 , 
    n1368 , 
    n1369 , 
    n1370 , 
    n1371 , 
    n1372 , 
    n1373 , 
    n1374 , 
    n1375 , 
    n1376 , 
    n1377 , 
    n1378 , 
    n1379 , 
    n1380 , 
    n1381 , 
    n1382 , 
    n1383 , 
    n1384 , 
    n1385 , 
    n1386 , 
    n1387 , 
    n1388 , 
    n1389 , 
    n1390 , 
    n1391 , 
    n1392 , 
    n1393 , 
    n1394 , 
    n1395 , 
    n1396 , 
    n1397 , 
    n1398 , 
    n1399 , 
    n1400 , 
    n1401 , 
    n1402 , 
    n1403 , 
    n1404 , 
    n1405 , 
    n1406 , 
    n1407 , 
    n1408 , 
    n1409 , 
    n1410 , 
    n1411 , 
    n1412 , 
    n1413 , 
    n1414 , 
    n1415 , 
    n1416 , 
    n1417 , 
    n1418 , 
    n1419 , 
    n1420 , 
    n1421 , 
    n1422 , 
    n1423 , 
    n1424 , 
    n1425 , 
    n1426 , 
    n1427 , 
    n1428 , 
    n1429 , 
    n1430 , 
    n1431 , 
    n1432 , 
    n1433 , 
    n1434 , 
    n1435 , 
    n1436 , 
    n1437 , 
    n1438 , 
    n1439 , 
    n1440 , 
    n1441 , 
    n1442 , 
    n1443 , 
    n1444 , 
    n1445 , 
    n1446 , 
    n1447 , 
    n1448 , 
    n1449 , 
    n1450 , 
    n1451 , 
    n1452 , 
    n1453 , 
    n1454 , 
    n1455 , 
    n1456 , 
    n1457 , 
    n1458 , 
    n1459 , 
    n1460 , 
    n1461 , 
    n1462 , 
    n1463 , 
    n1464 , 
    n1465 , 
    n1466 , 
    n1467 , 
    n1468 , 
    n1469 , 
    n1470 , 
    n1471 , 
    n1472 , 
    n1473 , 
    n1474 , 
    n1475 , 
    n1476 , 
    n1477 , 
    n1478 , 
    n1479 , 
    n1480 , 
    n1481 , 
    n1482 , 
    n1483 , 
    n1484 , 
    n1485 , 
    n1486 , 
    n1487 , 
    n1488 , 
    n1489 , 
    n1490 , 
    n1491 , 
    n1492 , 
    n1493 , 
    n1494 , 
    n1495 , 
    n1496 , 
    n1497 , 
    n1498 , 
    n1499 , 
    n1500 , 
    n1501 , 
    n1502 , 
    n1503 , 
    n1504 , 
    n1505 , 
    n1506 , 
    n1507 , 
    n1508 , 
    n1509 , 
    n1510 , 
    n1511 , 
    n1512 , 
    n1513 , 
    n1514 , 
    n1515 , 
    n1516 , 
    n1517 , 
    n1518 , 
    n1519 , 
    n1520 , 
    n1521 , 
    n1522 , 
    n1523 , 
    n1524 , 
    n1525 , 
    n1526 , 
    n1527 , 
    n1528 , 
    n1529 , 
    n1530 , 
    n1531 , 
    n1532 , 
    n1533 , 
    n1534 , 
    n1535 , 
    n1536 , 
    n1537 , 
    n1538 , 
    n1539 , 
    n1540 , 
    n1541 , 
    n1542 , 
    n1543 , 
    n1544 , 
    n1545 , 
    n1546 , 
    n1547 , 
    n1548 , 
    n1549 , 
    n1550 , 
    n1551 , 
    n1552 , 
    n1553 , 
    n1554 , 
    n1555 , 
    n1556 , 
    n1557 , 
    n1558 , 
    n1559 , 
    n1560 , 
    n1561 , 
    n1562 , 
    n1563 , 
    n1564 , 
    n1565 , 
    n1566 , 
    n1567 , 
    n1568 , 
    n1569 , 
    n1570 , 
    n1571 , 
    n1572 , 
    n1573 , 
    n1574 , 
    n1575 , 
    n1576 , 
    n1577 , 
    n1578 , 
    n1579 , 
    n1580 , 
    n1581 , 
    n1582 , 
    n1583 , 
    n1584 , 
    n1585 , 
    n1586 , 
    n1587 , 
    n1588 , 
    n1589 , 
    n1590 , 
    n1591 , 
    n1592 , 
    n1593 , 
    n1594 , 
    n1595 , 
    n1596 , 
    n1597 , 
    n1598 , 
    n1599 , 
    n1600 , 
    n1601 , 
    n1602 , 
    n1603 , 
    n1604 , 
    n1605 , 
    n1606 , 
    n1607 , 
    n1608 , 
    n1609 , 
    n1610 , 
    n1611 , 
    n1612 , 
    n1613 , 
    n1614 , 
    n1615 , 
    n1616 , 
    n1617 , 
    n1618 , 
    n1619 , 
    n1620 , 
    n1621 , 
    n1622 , 
    n1623 , 
    n1624 , 
    n1625 , 
    n1626 , 
    n1627 , 
    n1628 , 
    n1629 , 
    n1630 , 
    n1631 , 
    n1632 , 
    n1633 , 
    n1634 , 
    n1635 , 
    n1636 , 
    n1637 , 
    n1638 , 
    n1639 , 
    n1640 , 
    n1641 , 
    n1642 , 
    n1643 , 
    n1644 , 
    n1645 , 
    n1646 , 
    n1647 , 
    n1648 , 
    n1649 , 
    n1650 , 
    n1651 , 
    n1652 , 
    n1653 , 
    n1654 , 
    n1655 , 
    n1656 , 
    n1657 , 
    n1658 , 
    n1659 , 
    n1660 , 
    n1661 , 
    n1662 , 
    n1663 , 
    n1664 , 
    n1665 , 
    n1666 , 
    n1667 , 
    n1668 , 
    n1669 , 
    n1670 , 
    n1671 , 
    n1672 , 
    n1673 , 
    n1674 , 
    n1675 , 
    n1676 , 
    n1677 , 
    n1678 , 
    n1679 , 
    n1680 , 
    n1681 , 
    n1682 , 
    n1683 , 
    n1684 , 
    n1685 , 
    n1686 , 
    n1687 , 
    n1688 , 
    n1689 , 
    n1690 , 
    n1691 , 
    n1692 , 
    n1693 , 
    n1694 , 
    n1695 , 
    n1696 , 
    n1697 , 
    n1698 , 
    n1699 , 
    n1700 , 
    n1701 , 
    n1702 , 
    n1703 , 
    n1704 , 
    n1705 , 
    n1706 , 
    n1707 , 
    n1708 , 
    n1709 , 
    n1710 , 
    n1711 , 
    n1712 , 
    n1713 , 
    n1714 , 
    n1715 , 
    n1716 , 
    n1717 , 
    n1718 , 
    n1719 , 
    n1720 , 
    n1721 , 
    n1722 , 
    n1723 , 
    n1724 , 
    n1725 , 
    n1726 , 
    n1727 , 
    n1728 , 
    n1729 , 
    n1730 , 
    n1731 , 
    n1732 , 
    n1733 , 
    n1734 , 
    n1735 , 
    n1736 , 
    n1737 , 
    n1738 , 
    n1739 , 
    n1740 , 
    n1741 , 
    n1742 , 
    n1743 , 
    n1744 , 
    n1745 , 
    n1746 , 
    n1747 , 
    n1748 , 
    n1749 , 
    n1750 , 
    n1751 , 
    n1752 , 
    n1753 , 
    n1754 , 
    n1755 , 
    n1756 , 
    n1757 , 
    n1758 , 
    n1759 , 
    n1760 , 
    n1761 , 
    n1762 , 
    n1763 , 
    n1764 , 
    n1765 , 
    n1766 , 
    n1767 , 
    n1768 , 
    n1769 , 
    n1770 , 
    n1771 , 
    n1772 , 
    n1773 , 
    n1774 , 
    n1775 , 
    n1776 , 
    n1777 , 
    n1778 , 
    n1779 , 
    n1780 , 
    n1781 , 
    n1782 , 
    n1783 , 
    n1784 , 
    n1785 , 
    n1786 , 
    n1787 , 
    n1788 , 
    n1789 , 
    n1790 , 
    n1791 , 
    n1792 , 
    n1793 , 
    n1794 , 
    n1795 , 
    n1796 , 
    n1797 , 
    n1798 , 
    n1799 , 
    n1800 , 
    n1801 , 
    n1802 , 
    n1803 , 
    n1804 , 
    n1805 , 
    n1806 , 
    n1807 , 
    n1808 , 
    n1809 , 
    n1810 , 
    n1811 , 
    n1812 , 
    n1813 , 
    n1814 , 
    n1815 , 
    n1816 , 
    n1817 , 
    n1818 , 
    n1819 , 
    n1820 , 
    n1821 , 
    n1822 , 
    n1823 , 
    n1824 , 
    n1825 , 
    n1826 , 
    n1827 , 
    n1828 , 
    n1829 , 
    n1830 , 
    n1831 , 
    n1832 , 
    n1833 , 
    n1834 , 
    n1835 , 
    n1836 , 
    n1837 , 
    n1838 , 
    n1839 , 
    n1840 , 
    n1841 , 
    n1842 , 
    n1843 , 
    n1844 , 
    n1845 , 
    n1846 , 
    n1847 , 
    n1848 , 
    n1849 , 
    n1850 , 
    n1851 , 
    n1852 , 
    n1853 , 
    n1854 , 
    n1855 , 
    n1856 , 
    n1857 , 
    n1858 , 
    n1859 , 
    n1860 , 
    n1861 , 
    n1862 , 
    n1863 , 
    n1864 , 
    n1865 , 
    n1866 , 
    n1867 , 
    n1868 , 
    n1869 , 
    n1870 , 
    n1871 , 
    n1872 , 
    n1873 , 
    n1874 , 
    n1875 , 
    n1876 , 
    n1877 , 
    n1878 , 
    n1879 , 
    n1880 , 
    n1881 , 
    n1882 , 
    n1883 , 
    n1884 , 
    n1885 , 
    n1886 , 
    n1887 , 
    n1888 , 
    n1889 , 
    n1890 , 
    n1891 , 
    n1892 , 
    n1893 , 
    n1894 , 
    n1895 , 
    n1896 , 
    n1897 , 
    n1898 , 
    n1899 , 
    n1900 , 
    n1901 , 
    n1902 , 
    n1903 , 
    n1904 , 
    n1905 , 
    n1906 , 
    n1907 , 
    n1908 , 
    n1909 , 
    n1910 , 
    n1911 , 
    n1912 , 
    n1913 , 
    n1914 , 
    n1915 , 
    n1916 , 
    n1917 , 
    n1918 , 
    n1919 , 
    n1920 , 
    n1921 , 
    n1922 , 
    n1923 , 
    n1924 , 
    n1925 , 
    n1926 , 
    n1927 , 
    n1928 , 
    n1929 , 
    n1930 , 
    n1931 , 
    n1932 , 
    n1933 , 
    n1934 , 
    n1935 , 
    n1936 , 
    n1937 , 
    n1938 , 
    n1939 , 
    n1940 , 
    n1941 , 
    n1942 , 
    n1943 , 
    n1944 , 
    n1945 , 
    n1946 , 
    n1947 , 
    n1948 , 
    n1949 , 
    n1950 , 
    n1951 , 
    n1952 , 
    n1953 , 
    n1954 , 
    n1955 , 
    n1956 , 
    n1957 , 
    n1958 , 
    n1959 , 
    n1960 , 
    n1961 , 
    n1962 , 
    n1963 , 
    n1964 , 
    n1965 , 
    n1966 , 
    n1967 , 
    n1968 , 
    n1969 , 
    n1970 , 
    n1971 , 
    n1972 , 
    n1973 , 
    n1974 , 
    n1975 , 
    n1976 , 
    n1977 , 
    n1978 , 
    n1979 , 
    n1980 , 
    n1981 , 
    n1982 , 
    n1983 , 
    n1984 , 
    n1985 , 
    n1986 , 
    n1987 , 
    n1988 , 
    n1989 , 
    n1990 , 
    n1991 , 
    n1992 , 
    n1993 , 
    n1994 , 
    n1995 , 
    n1996 , 
    n1997 , 
    n1998 , 
    n1999 , 
    n2000 , 
    n2001 , 
    n2002 , 
    n2003 , 
    n2004 , 
    n2005 , 
    n2006 , 
    n2007 , 
    n2008 , 
    n2009 , 
    n2010 , 
    n2011 , 
    n2012 , 
    n2013 , 
    n2014 , 
    n2015 , 
    n2016 , 
    n2017 , 
    n2018 , 
    n2019 , 
    n2020 , 
    n2021 , 
    n2022 , 
    n2023 , 
    n2024 , 
    n2025 , 
    n2026 , 
    n2027 , 
    n2028 , 
    n2029 , 
    n2030 , 
    n2031 , 
    n2032 , 
    n2033 , 
    n2034 , 
    n2035 , 
    n2036 , 
    n2037 , 
    n2038 , 
    n2039 , 
    n2040 , 
    n2041 , 
    n2042 , 
    n2043 , 
    n2044 , 
    n2045 , 
    n2046 , 
    n2047 , 
    n2048 , 
    n2049 , 
    n2050 , 
    n2051 , 
    n2052 , 
    n2053 , 
    n2054 , 
    n2055 , 
    n2056 , 
    n2057 , 
    n2058 , 
    n2059 , 
    n2060 , 
    n2061 , 
    n2062 , 
    n2063 , 
    n2064 , 
    n2065 , 
    n2066 , 
    n2067 , 
    n2068 , 
    n2069 , 
    n2070 , 
    n2071 , 
    n2072 , 
    n2073 , 
    n2074 , 
    n2075 , 
    n2076 , 
    n2077 , 
    n2078 , 
    n2079 , 
    n2080 , 
    n2081 , 
    n2082 , 
    n2083 , 
    n2084 , 
    n2085 , 
    n2086 , 
    n2087 , 
    n2088 , 
    n2089 , 
    n2090 , 
    n2091 , 
    n2092 , 
    n2093 , 
    n2094 , 
    n2095 , 
    n2096 , 
    n2097 , 
    n2098 , 
    n2099 , 
    n2100 , 
    n2101 , 
    n2102 , 
    n2103 , 
    n2104 , 
    n2105 , 
    n2106 , 
    n2107 , 
    n2108 , 
    n2109 , 
    n2110 , 
    n2111 , 
    n2112 , 
    n2113 , 
    n2114 , 
    n2115 , 
    n2116 , 
    n2117 , 
    n2118 , 
    n2119 , 
    n2120 , 
    n2121 , 
    n2122 , 
    n2123 , 
    n2124 , 
    n2125 , 
    n2126 , 
    n2127 , 
    n2128 , 
    n2129 , 
    n2130 , 
    n2131 , 
    n2132 , 
    n2133 , 
    n2134 , 
    n2135 , 
    n2136 , 
    n2137 , 
    n2138 , 
    n2139 , 
    n2140 , 
    n2141 , 
    n2142 , 
    n2143 , 
    n2144 , 
    n2145 , 
    n2146 , 
    n2147 , 
    n2148 , 
    n2149 , 
    n2150 , 
    n2151 , 
    n2152 , 
    n2153 , 
    n2154 , 
    n2155 , 
    n2156 , 
    n2157 , 
    n2158 , 
    n2159 , 
    n2160 , 
    n2161 , 
    n2162 , 
    n2163 , 
    n2164 , 
    n2165 , 
    n2166 , 
    n2167 , 
    n2168 , 
    n2169 , 
    n2170 , 
    n2171 , 
    n2172 , 
    n2173 , 
    n2174 , 
    n2175 , 
    n2176 , 
    n2177 , 
    n2178 , 
    n2179 , 
    n2180 , 
    n2181 , 
    n2182 , 
    n2183 , 
    n2184 , 
    n2185 , 
    n2186 , 
    n2187 , 
    n2188 , 
    n2189 , 
    n2190 , 
    n2191 , 
    n2192 , 
    n2193 , 
    n2194 , 
    n2195 , 
    n2196 , 
    n2197 , 
    n2198 , 
    n2199 , 
    n2200 , 
    n2201 , 
    n2202 , 
    n2203 , 
    n2204 , 
    n2205 , 
    n2206 , 
    n2207 , 
    n2208 , 
    n2209 , 
    n2210 , 
    n2211 , 
    n2212 , 
    n2213 , 
    n2214 , 
    n2215 , 
    n2216 , 
    n2217 , 
    n2218 , 
    n2219 , 
    n2220 , 
    n2221 , 
    n2222 , 
    n2223 , 
    n2224 , 
    n2225 , 
    n2226 , 
    n2227 , 
    n2228 , 
    n2229 , 
    n2230 , 
    n2231 , 
    n2232 , 
    n2233 , 
    n2234 , 
    n2235 , 
    n2236 , 
    n2237 , 
    n2238 , 
    n2239 , 
    n2240 , 
    n2241 , 
    n2242 , 
    n2243 , 
    n2244 , 
    n2245 , 
    n2246 , 
    n2247 , 
    n2248 , 
    n2249 , 
    n2250 , 
    n2251 , 
    n2252 , 
    n2253 , 
    n2254 , 
    n2255 , 
    n2256 , 
    n2257 , 
    n2258 , 
    n2259 , 
    n2260 , 
    n2261 , 
    n2262 , 
    n2263 , 
    n2264 , 
    n2265 , 
    n2266 , 
    n2267 , 
    n2268 , 
    n2269 , 
    n2270 , 
    n2271 , 
    n2272 , 
    n2273 , 
    n2274 , 
    n2275 , 
    n2276 , 
    n2277 , 
    n2278 , 
    n2279 , 
    n2280 , 
    n2281 , 
    n2282 , 
    n2283 , 
    n2284 , 
    n2285 , 
    n2286 , 
    n2287 , 
    n2288 , 
    n2289 , 
    n2290 , 
    n2291 , 
    n2292 , 
    n2293 , 
    n2294 , 
    n2295 , 
    n2296 , 
    n2297 , 
    n2298 , 
    n2299 , 
    n2300 , 
    n2301 , 
    n2302 , 
    n2303 , 
    n2304 , 
    n2305 , 
    n2306 , 
    n2307 , 
    n2308 , 
    n2309 , 
    n2310 , 
    n2311 , 
    n2312 , 
    n2313 , 
    n2314 , 
    n2315 , 
    n2316 , 
    n2317 , 
    n2318 , 
    n2319 , 
    n2320 , 
    n2321 , 
    n2322 , 
    n2323 , 
    n2324 , 
    n2325 , 
    n2326 , 
    n2327 , 
    n2328 , 
    n2329 , 
    n2330 , 
    n2331 , 
    n2332 , 
    n2333 , 
    n2334 , 
    n2335 , 
    n2336 , 
    n2337 , 
    n2338 , 
    n2339 , 
    n2340 , 
    n2341 , 
    n2342 , 
    n2343 , 
    n2344 , 
    n2345 , 
    n2346 , 
    n2347 , 
    n2348 , 
    n2349 , 
    n2350 , 
    n2351 , 
    n2352 , 
    n2353 , 
    n2354 , 
    n2355 , 
    n2356 , 
    n2357 , 
    n2358 , 
    n2359 , 
    n2360 , 
    n2361 , 
    n2362 , 
    n2363 , 
    n2364 , 
    n2365 , 
    n2366 , 
    n2367 , 
    n2368 , 
    n2369 , 
    n2370 , 
    n2371 , 
    n2372 , 
    n2373 , 
    n2374 , 
    n2375 , 
    n2376 , 
    n2377 , 
    n2378 , 
    n2379 , 
    n2380 , 
    n2381 , 
    n2382 , 
    n2383 , 
    n2384 , 
    n2385 , 
    n2386 , 
    n2387 , 
    n2388 , 
    n2389 , 
    n2390 , 
    n2391 , 
    n2392 , 
    n2393 , 
    n2394 , 
    n2395 , 
    n2396 , 
    n2397 , 
    n2398 , 
    n2399 , 
    n2400 , 
    n2401 , 
    n2402 , 
    n2403 , 
    n2404 , 
    n2405 , 
    n2406 , 
    n2407 , 
    n2408 , 
    n2409 , 
    n2410 , 
    n2411 , 
    n2412 , 
    n2413 , 
    n2414 , 
    n2415 , 
    n2416 , 
    n2417 , 
    n2418 , 
    n2419 , 
    n2420 , 
    n2421 , 
    n2422 , 
    n2423 , 
    n2424 , 
    n2425 , 
    n2426 , 
    n2427 , 
    n2428 , 
    n2429 , 
    n2430 , 
    n2431 , 
    n2432 , 
    n2433 , 
    n2434 , 
    n2435 , 
    n2436 , 
    n2437 , 
    n2438 , 
    n2439 , 
    n2440 , 
    n2441 , 
    n2442 , 
    n2443 , 
    n2444 , 
    n2445 , 
    n2446 , 
    n2447 , 
    n2448 , 
    n2449 , 
    n2450 , 
    n2451 , 
    n2452 , 
    n2453 , 
    n2454 , 
    n2455 , 
    n2456 , 
    n2457 , 
    n2458 , 
    n2459 , 
    n2460 , 
    n2461 , 
    n2462 , 
    n2463 , 
    n2464 , 
    n2465 , 
    n2466 , 
    n2467 , 
    n2468 , 
    n2469 , 
    n2470 , 
    n2471 , 
    n2472 , 
    n2473 , 
    n2474 , 
    n2475 , 
    n2476 , 
    n2477 , 
    n2478 , 
    n2479 , 
    n2480 , 
    n2481 , 
    n2482 , 
    n2483 , 
    n2484 , 
    n2485 , 
    n2486 , 
    n2487 , 
    n2488 , 
    n2489 , 
    n2490 , 
    n2491 , 
    n2492 , 
    n2493 , 
    n2494 , 
    n2495 , 
    n2496 , 
    n2497 , 
    n2498 , 
    n2499 , 
    n2500 , 
    n2501 , 
    n2502 , 
    n2503 , 
    n2504 , 
    n2505 , 
    n2506 , 
    n2507 , 
    n2508 , 
    n2509 , 
    n2510 , 
    n2511 , 
    n2512 , 
    n2513 , 
    n2514 , 
    n2515 , 
    n2516 , 
    n2517 , 
    n2518 , 
    n2519 , 
    n2520 , 
    n2521 , 
    n2522 , 
    n2523 , 
    n2524 , 
    n2525 , 
    n2526 , 
    n2527 , 
    n2528 , 
    n2529 , 
    n2530 , 
    n2531 , 
    n2532 , 
    n2533 , 
    n2534 , 
    n2535 , 
    n2536 , 
    n2537 , 
    n2538 , 
    n2539 , 
    n2540 , 
    n2541 , 
    n2542 , 
    n2543 , 
    n2544 , 
    n2545 , 
    n2546 , 
    n2547 , 
    n2548 , 
    n2549 , 
    n2550 , 
    n2551 , 
    n2552 , 
    n2553 , 
    n2554 , 
    n2555 , 
    n2556 , 
    n2557 , 
    n2558 , 
    n2559 , 
    n2560 , 
    n2561 , 
    n2562 , 
    n2563 , 
    n2564 , 
    n2565 , 
    n2566 , 
    n2567 , 
    n2568 , 
    n2569 , 
    n2570 , 
    n2571 , 
    n2572 , 
    n2573 , 
    n2574 , 
    n2575 , 
    n2576 , 
    n2577 , 
    n2578 , 
    n2579 , 
    n2580 , 
    n2581 , 
    n2582 , 
    n2583 , 
    n2584 , 
    n2585 , 
    n2586 , 
    n2587 , 
    n2588 , 
    n2589 , 
    n2590 , 
    n2591 , 
    n2592 , 
    n2593 , 
    n2594 , 
    n2595 , 
    n2596 , 
    n2597 , 
    n2598 , 
    n2599 , 
    n2600 , 
    n2601 , 
    n2602 , 
    n2603 , 
    n2604 , 
    n2605 , 
    n2606 , 
    n2607 , 
    n2608 , 
    n2609 , 
    n2610 , 
    n2611 , 
    n2612 , 
    n2613 , 
    n2614 , 
    n2615 , 
    n2616 , 
    n2617 , 
    n2618 , 
    n2619 , 
    n2620 , 
    n2621 , 
    n2622 , 
    n2623 , 
    n2624 , 
    n2625 , 
    n2626 , 
    n2627 , 
    n2628 , 
    n2629 , 
    n2630 , 
    n2631 , 
    n2632 , 
    n2633 , 
    n2634 , 
    n2635 , 
    n2636 , 
    n2637 , 
    n2638 , 
    n2639 , 
    n2640 , 
    n2641 , 
    n2642 , 
    n2643 , 
    n2644 , 
    n2645 , 
    n2646 , 
    n2647 , 
    n2648 , 
    n2649 , 
    n2650 , 
    n2651 , 
    n2652 , 
    n2653 , 
    n2654 , 
    n2655 , 
    n2656 , 
    n2657 , 
    n2658 , 
    n2659 , 
    n2660 , 
    n2661 , 
    n2662 , 
    n2663 , 
    n2664 , 
    n2665 , 
    n2666 , 
    n2667 , 
    n2668 , 
    n2669 , 
    n2670 , 
    n2671 , 
    n2672 , 
    n2673 , 
    n2674 , 
    n2675 , 
    n2676 , 
    n2677 , 
    n2678 , 
    n2679 , 
    n2680 , 
    n2681 , 
    n2682 , 
    n2683 , 
    n2684 , 
    n2685 , 
    n2686 , 
    n2687 , 
    n2688 , 
    n2689 , 
    n2690 , 
    n2691 , 
    n2692 , 
    n2693 , 
    n2694 , 
    n2695 , 
    n2696 , 
    n2697 , 
    n2698 , 
    n2699 , 
    n2700 , 
    n2701 , 
    n2702 , 
    n2703 , 
    n2704 , 
    n2705 , 
    n2706 , 
    n2707 , 
    n2708 , 
    n2709 , 
    n2710 , 
    n2711 , 
    n2712 , 
    n2713 , 
    n2714 , 
    n2715 , 
    n2716 , 
    n2717 , 
    n2718 , 
    n2719 , 
    n2720 , 
    n2721 , 
    n2722 , 
    n2723 , 
    n2724 , 
    n2725 , 
    n2726 , 
    n2727 , 
    n2728 , 
    n2729 , 
    n2730 , 
    n2731 , 
    n2732 , 
    n2733 , 
    n2734 , 
    n2735 , 
    n2736 , 
    n2737 , 
    n2738 , 
    n2739 , 
    n2740 , 
    n2741 , 
    n2742 , 
    n2743 , 
    n2744 , 
    n2745 , 
    n2746 , 
    n2747 , 
    n2748 , 
    n2749 , 
    n2750 , 
    n2751 , 
    n2752 , 
    n2753 , 
    n2754 , 
    n2755 , 
    n2756 , 
    n2757 , 
    n2758 , 
    n2759 , 
    n2760 , 
    n2761 , 
    n2762 , 
    n2763 , 
    n2764 , 
    n2765 , 
    n2766 , 
    n2767 , 
    n2768 , 
    n2769 , 
    n2770 , 
    n2771 , 
    n2772 , 
    n2773 , 
    n2774 , 
    n2775 , 
    n2776 , 
    n2777 , 
    n2778 , 
    n2779 , 
    n2780 , 
    n2781 , 
    n2782 , 
    n2783 , 
    n2784 , 
    n2785 , 
    n2786 , 
    n2787 , 
    n2788 , 
    n2789 , 
    n2790 , 
    n2791 , 
    n2792 , 
    n2793 , 
    n2794 , 
    n2795 , 
    n2796 , 
    n2797 , 
    n2798 , 
    n2799 , 
    n2800 , 
    n2801 , 
    n2802 , 
    n2803 , 
    n2804 , 
    n2805 , 
    n2806 , 
    n2807 , 
    n2808 , 
    n2809 , 
    n2810 , 
    n2811 , 
    n2812 , 
    n2813 , 
    n2814 , 
    n2815 , 
    n2816 , 
    n2817 , 
    n2818 , 
    n2819 , 
    n2820 , 
    n2821 , 
    n2822 , 
    n2823 , 
    n2824 , 
    n2825 , 
    n2826 , 
    n2827 , 
    n2828 , 
    n2829 , 
    n2830 , 
    n2831 , 
    n2832 , 
    n2833 , 
    n2834 , 
    n2835 , 
    n2836 , 
    n2837 , 
    n2838 , 
    n2839 , 
    n2840 , 
    n2841 , 
    n2842 , 
    n2843 , 
    n2844 , 
    n2845 , 
    n2846 , 
    n2847 , 
    n2848 , 
    n2849 , 
    n2850 , 
    n2851 , 
    n2852 , 
    n2853 , 
    n2854 , 
    n2855 , 
    n2856 , 
    n2857 , 
    n2858 , 
    n2859 , 
    n2860 , 
    n2861 , 
    n2862 , 
    n2863 , 
    n2864 , 
    n2865 , 
    n2866 , 
    n2867 , 
    n2868 , 
    n2869 , 
    n2870 , 
    n2871 , 
    n2872 , 
    n2873 , 
    n2874 , 
    n2875 , 
    n2876 , 
    n2877 , 
    n2878 , 
    n2879 , 
    n2880 , 
    n2881 , 
    n2882 , 
    n2883 , 
    n2884 , 
    n2885 , 
    n2886 , 
    n2887 , 
    n2888 , 
    n2889 , 
    n2890 , 
    n2891 , 
    n2892 , 
    n2893 , 
    n2894 , 
    n2895 , 
    n2896 , 
    n2897 , 
    n2898 , 
    n2899 , 
    n2900 , 
    n2901 , 
    n2902 , 
    n2903 , 
    n2904 , 
    n2905 , 
    n2906 , 
    n2907 , 
    n2908 , 
    n2909 , 
    n2910 , 
    n2911 , 
    n2912 , 
    n2913 , 
    n2914 , 
    n2915 , 
    n2916 , 
    n2917 , 
    n2918 , 
    n2919 , 
    n2920 , 
    n2921 , 
    n2922 , 
    n2923 , 
    n2924 , 
    n2925 , 
    n2926 , 
    n2927 , 
    n2928 , 
    n2929 , 
    n2930 , 
    n2931 , 
    n2932 , 
    n2933 , 
    n2934 , 
    n2935 , 
    n2936 , 
    n2937 , 
    n2938 , 
    n2939 , 
    n2940 , 
    n2941 , 
    n2942 , 
    n2943 , 
    n2944 , 
    n2945 , 
    n2946 , 
    n2947 , 
    n2948 , 
    n2949 , 
    n2950 , 
    n2951 , 
    n2952 , 
    n2953 , 
    n2954 , 
    n2955 , 
    n2956 , 
    n2957 , 
    n2958 , 
    n2959 , 
    n2960 , 
    n2961 , 
    n2962 , 
    n2963 , 
    n2964 , 
    n2965 , 
    n2966 , 
    n2967 , 
    n2968 , 
    n2969 , 
    n2970 , 
    n2971 , 
    n2972 , 
    n2973 , 
    n2974 , 
    n2975 , 
    n2976 , 
    n2977 , 
    n2978 , 
    n2979 , 
    n2980 , 
    n2981 , 
    n2982 , 
    n2983 , 
    n2984 , 
    n2985 , 
    n2986 , 
    n2987 , 
    n2988 , 
    n2989 , 
    n2990 , 
    n2991 , 
    n2992 , 
    n2993 , 
    n2994 , 
    n2995 , 
    n2996 , 
    n2997 , 
    n2998 , 
    n2999 , 
    n3000 , 
    n3001 , 
    n3002 , 
    n3003 , 
    n3004 , 
    n3005 , 
    n3006 , 
    n3007 , 
    n3008 , 
    n3009 , 
    n3010 , 
    n3011 , 
    n3012 , 
    n3013 , 
    n3014 , 
    n3015 , 
    n3016 , 
    n3017 , 
    n3018 , 
    n3019 , 
    n3020 , 
    n3021 , 
    n3022 , 
    n3023 , 
    n3024 , 
    n3025 , 
    n3026 , 
    n3027 , 
    n3028 , 
    n3029 , 
    n3030 , 
    n3031 , 
    n3032 , 
    n3033 , 
    n3034 , 
    n3035 , 
    n3036 , 
    n3037 , 
    n3038 , 
    n3039 , 
    n3040 , 
    n3041 , 
    n3042 , 
    n3043 , 
    n3044 , 
    n3045 , 
    n3046 , 
    n3047 , 
    n3048 , 
    n3049 , 
    n3050 , 
    n3051 , 
    n3052 , 
    n3053 , 
    n3054 , 
    n3055 , 
    n3056 , 
    n3057 , 
    n3058 , 
    n3059 , 
    n3060 , 
    n3061 , 
    n3062 , 
    n3063 , 
    n3064 , 
    n3065 , 
    n3066 , 
    n3067 , 
    n3068 , 
    n3069 , 
    n3070 , 
    n3071 , 
    n3072 , 
    n3073 , 
    n3074 , 
    n3075 , 
    n3076 , 
    n3077 , 
    n3078 , 
    n3079 , 
    n3080 , 
    n3081 , 
    n3082 , 
    n3083 , 
    n3084 , 
    n3085 , 
    n3086 , 
    n3087 , 
    n3088 , 
    n3089 , 
    n3090 , 
    n3091 , 
    n3092 , 
    n3093 , 
    n3094 , 
    n3095 , 
    n3096 , 
    n3097 , 
    n3098 , 
    n3099 , 
    n3100 , 
    n3101 , 
    n3102 , 
    n3103 , 
    n3104 , 
    n3105 , 
    n3106 , 
    n3107 , 
    n3108 , 
    n3109 , 
    n3110 , 
    n3111 , 
    n3112 , 
    n3113 , 
    n3114 , 
    n3115 , 
    n3116 , 
    n3117 , 
    n3118 , 
    n3119 , 
    n3120 , 
    n3121 , 
    n3122 , 
    n3123 , 
    n3124 , 
    n3125 , 
    n3126 , 
    n3127 , 
    n3128 , 
    n3129 , 
    n3130 , 
    n3131 , 
    n3132 , 
    n3133 , 
    n3134 , 
    n3135 , 
    n3136 , 
    n3137 , 
    n3138 , 
    n3139 , 
    n3140 , 
    n3141 , 
    n3142 , 
    n3143 , 
    n3144 , 
    n3145 , 
    n3146 , 
    n3147 , 
    n3148 , 
    n3149 , 
    n3150 , 
    n3151 , 
    n3152 , 
    n3153 , 
    n3154 , 
    n3155 , 
    n3156 , 
    n3157 , 
    n3158 , 
    n3159 , 
    n3160 , 
    n3161 , 
    n3162 , 
    n3163 , 
    n3164 , 
    n3165 , 
    n3166 , 
    n3167 , 
    n3168 , 
    n3169 , 
    n3170 , 
    n3171 , 
    n3172 , 
    n3173 , 
    n3174 , 
    n3175 , 
    n3176 , 
    n3177 , 
    n3178 , 
    n3179 , 
    n3180 , 
    n3181 , 
    n3182 , 
    n3183 , 
    n3184 , 
    n3185 , 
    n3186 , 
    n3187 , 
    n3188 , 
    n3189 , 
    n3190 , 
    n3191 , 
    n3192 , 
    n3193 , 
    n3194 , 
    n3195 , 
    n3196 , 
    n3197 , 
    n3198 , 
    n3199 , 
    n3200 , 
    n3201 , 
    n3202 , 
    n3203 , 
    n3204 , 
    n3205 , 
    n3206 , 
    n3207 , 
    n3208 , 
    n3209 , 
    n3210 , 
    n3211 , 
    n3212 , 
    n3213 , 
    n3214 , 
    n3215 , 
    n3216 , 
    n3217 , 
    n3218 , 
    n3219 , 
    n3220 , 
    n3221 , 
    n3222 , 
    n3223 , 
    n3224 , 
    n3225 , 
    n3226 , 
    n3227 , 
    n3228 , 
    n3229 , 
    n3230 , 
    n3231 , 
    n3232 , 
    n3233 , 
    n3234 , 
    n3235 , 
    n3236 , 
    n3237 , 
    n3238 , 
    n3239 , 
    n3240 , 
    n3241 , 
    n3242 , 
    n3243 , 
    n3244 , 
    n3245 , 
    n3246 , 
    n3247 , 
    n3248 , 
    n3249 , 
    n3250 , 
    n3251 , 
    n3252 , 
    n3253 , 
    n3254 , 
    n3255 , 
    n3256 , 
    n3257 , 
    n3258 , 
    n3259 , 
    n3260 , 
    n3261 , 
    n3262 , 
    n3263 , 
    n3264 , 
    n3265 , 
    n3266 , 
    n3267 , 
    n3268 , 
    n3269 , 
    n3270 , 
    n3271 , 
    n3272 , 
    n3273 , 
    n3274 , 
    n3275 , 
    n3276 , 
    n3277 , 
    n3278 , 
    n3279 , 
    n3280 , 
    n3281 , 
    n3282 , 
    n3283 , 
    n3284 , 
    n3285 , 
    n3286 , 
    n3287 , 
    n3288 , 
    n3289 , 
    n3290 , 
    n3291 , 
    n3292 , 
    n3293 , 
    n3294 , 
    n3295 , 
    n3296 , 
    n3297 , 
    n3298 , 
    n3299 , 
    n3300 , 
    n3301 , 
    n3302 , 
    n3303 , 
    n3304 , 
    n3305 , 
    n3306 , 
    n3307 , 
    n3308 , 
    n3309 , 
    n3310 , 
    n3311 , 
    n3312 , 
    n3313 , 
    n3314 , 
    n3315 , 
    n3316 , 
    n3317 , 
    n3318 , 
    n3319 , 
    n3320 , 
    n3321 , 
    n3322 , 
    n3323 , 
    n3324 , 
    n3325 , 
    n3326 , 
    n3327 , 
    n3328 , 
    n3329 , 
    n3330 , 
    n3331 , 
    n3332 , 
    n3333 , 
    n3334 , 
    n3335 , 
    n3336 , 
    n3337 , 
    n3338 , 
    n3339 , 
    n3340 , 
    n3341 , 
    n3342 , 
    n3343 , 
    n3344 , 
    n3345 , 
    n3346 , 
    n3347 , 
    n3348 , 
    n3349 , 
    n3350 , 
    n3351 , 
    n3352 , 
    n3353 , 
    n3354 , 
    n3355 , 
    n3356 , 
    n3357 , 
    n3358 , 
    n3359 , 
    n3360 , 
    n3361 , 
    n3362 , 
    n3363 , 
    n3364 , 
    n3365 , 
    n3366 , 
    n3367 , 
    n3368 , 
    n3369 , 
    n3370 , 
    n3371 , 
    n3372 , 
    n3373 , 
    n3374 , 
    n3375 , 
    n3376 , 
    n3377 , 
    n3378 , 
    n3379 , 
    n3380 , 
    n3381 , 
    n3382 , 
    n3383 , 
    n3384 , 
    n3385 , 
    n3386 , 
    n3387 , 
    n3388 , 
    n3389 , 
    n3390 , 
    n3391 , 
    n3392 , 
    n3393 , 
    n3394 , 
    n3395 , 
    n3396 , 
    n3397 , 
    n3398 , 
    n3399 , 
    n3400 , 
    n3401 , 
    n3402 , 
    n3403 , 
    n3404 , 
    n3405 , 
    n3406 , 
    n3407 , 
    n3408 , 
    n3409 , 
    n3410 , 
    n3411 , 
    n3412 , 
    n3413 , 
    n3414 , 
    n3415 , 
    n3416 , 
    n3417 , 
    n3418 , 
    n3419 , 
    n3420 , 
    n3421 , 
    n3422 , 
    n3423 , 
    n3424 , 
    n3425 , 
    n3426 , 
    n3427 , 
    n3428 , 
    n3429 , 
    n3430 , 
    n3431 , 
    n3432 , 
    n3433 , 
    n3434 , 
    n3435 , 
    n3436 , 
    n3437 , 
    n3438 , 
    n3439 , 
    n3440 , 
    n3441 , 
    n3442 , 
    n3443 , 
    n3444 , 
    n3445 , 
    n3446 , 
    n3447 , 
    n3448 , 
    n3449 , 
    n3450 , 
    n3451 , 
    n3452 , 
    n3453 , 
    n3454 , 
    n3455 , 
    n3456 , 
    n3457 , 
    n3458 , 
    n3459 , 
    n3460 , 
    n3461 , 
    n3462 , 
    n3463 , 
    n3464 , 
    n3465 , 
    n3466 , 
    n3467 , 
    n3468 , 
    n3469 , 
    n3470 , 
    n3471 , 
    n3472 , 
    n3473 , 
    n3474 , 
    n3475 , 
    n3476 , 
    n3477 , 
    n3478 , 
    n3479 , 
    n3480 , 
    n3481 , 
    n3482 , 
    n3483 , 
    n3484 , 
    n3485 , 
    n3486 , 
    n3487 , 
    n3488 , 
    n3489 , 
    n3490 , 
    n3491 , 
    n3492 , 
    n3493 , 
    n3494 , 
    n3495 , 
    n3496 , 
    n3497 , 
    n3498 , 
    n3499 , 
    n3500 , 
    n3501 , 
    n3502 , 
    n3503 , 
    n3504 , 
    n3505 , 
    n3506 , 
    n3507 , 
    n3508 , 
    n3509 , 
    n3510 , 
    n3511 , 
    n3512 , 
    n3513 , 
    n3514 , 
    n3515 , 
    n3516 , 
    n3517 , 
    n3518 , 
    n3519 , 
    n3520 , 
    n3521 , 
    n3522 , 
    n3523 , 
    n3524 , 
    n3525 , 
    n3526 , 
    n3527 , 
    n3528 , 
    n3529 , 
    n3530 , 
    n3531 , 
    n3532 , 
    n3533 , 
    n3534 , 
    n3535 , 
    n3536 , 
    n3537 , 
    n3538 , 
    n3539 , 
    n3540 , 
    n3541 , 
    n3542 , 
    n3543 , 
    n3544 , 
    n3545 , 
    n3546 , 
    n3547 , 
    n3548 , 
    n3549 , 
    n3550 , 
    n3551 , 
    n3552 , 
    n3553 , 
    n3554 , 
    n3555 , 
    n3556 , 
    n3557 , 
    n3558 , 
    n3559 , 
    n3560 , 
    n3561 , 
    n3562 , 
    n3563 , 
    n3564 , 
    n3565 , 
    n3566 , 
    n3567 , 
    n3568 , 
    n3569 , 
    n3570 , 
    n3571 , 
    n3572 , 
    n3573 , 
    n3574 , 
    n3575 , 
    n3576 , 
    n3577 , 
    n3578 , 
    n3579 , 
    n3580 , 
    n3581 , 
    n3582 , 
    n3583 , 
    n3584 , 
    n3585 , 
    n3586 , 
    n3587 , 
    n3588 , 
    n3589 , 
    n3590 , 
    n3591 , 
    n3592 , 
    n3593 , 
    n3594 , 
    n3595 , 
    n3596 , 
    n3597 , 
    n3598 , 
    n3599 , 
    n3600 , 
    n3601 , 
    n3602 , 
    n3603 , 
    n3604 , 
    n3605 , 
    n3606 , 
    n3607 , 
    n3608 , 
    n3609 , 
    n3610 , 
    n3611 , 
    n3612 , 
    n3613 , 
    n3614 , 
    n3615 , 
    n3616 , 
    n3617 , 
    n3618 , 
    n3619 , 
    n3620 , 
    n3621 , 
    n3622 , 
    n3623 , 
    n3624 , 
    n3625 , 
    n3626 , 
    n3627 , 
    n3628 , 
    n3629 , 
    n3630 , 
    n3631 , 
    n3632 , 
    n3633 , 
    n3634 , 
    n3635 , 
    n3636 , 
    n3637 , 
    n3638 , 
    n3639 , 
    n3640 , 
    n3641 , 
    n3642 , 
    n3643 , 
    n3644 , 
    n3645 , 
    n3646 , 
    n3647 , 
    n3648 , 
    n3649 , 
    n3650 , 
    n3651 , 
    n3652 , 
    n3653 , 
    n3654 , 
    n3655 , 
    n3656 , 
    n3657 , 
    n3658 , 
    n3659 , 
    n3660 , 
    n3661 , 
    n3662 , 
    n3663 , 
    n3664 , 
    n3665 , 
    n3666 , 
    n3667 , 
    n3668 , 
    n3669 , 
    n3670 , 
    n3671 , 
    n3672 , 
    n3673 , 
    n3674 , 
    n3675 , 
    n3676 , 
    n3677 , 
    n3678 , 
    n3679 , 
    n3680 , 
    n3681 , 
    n3682 , 
    n3683 , 
    n3684 , 
    n3685 , 
    n3686 , 
    n3687 , 
    n3688 , 
    n3689 , 
    n3690 , 
    n3691 , 
    n3692 , 
    n3693 , 
    n3694 , 
    n3695 , 
    n3696 , 
    n3697 , 
    n3698 , 
    n3699 , 
    n3700 , 
    n3701 , 
    n3702 , 
    n3703 , 
    n3704 , 
    n3705 , 
    n3706 , 
    n3707 , 
    n3708 , 
    n3709 , 
    n3710 , 
    n3711 , 
    n3712 , 
    n3713 , 
    n3714 , 
    n3715 , 
    n3716 , 
    n3717 , 
    n3718 , 
    n3719 , 
    n3720 , 
    n3721 , 
    n3722 , 
    n3723 , 
    n3724 , 
    n3725 , 
    n3726 , 
    n3727 , 
    n3728 , 
    n3729 , 
    n3730 , 
    n3731 , 
    n3732 , 
    n3733 , 
    n3734 , 
    n3735 , 
    n3736 , 
    n3737 , 
    n3738 , 
    n3739 , 
    n3740 , 
    n3741 , 
    n3742 , 
    n3743 , 
    n3744 , 
    n3745 , 
    n3746 , 
    n3747 , 
    n3748 , 
    n3749 , 
    n3750 , 
    n3751 , 
    n3752 , 
    n3753 , 
    n3754 , 
    n3755 , 
    n3756 , 
    n3757 , 
    n3758 , 
    n3759 , 
    n3760 , 
    n3761 , 
    n3762 , 
    n3763 , 
    n3764 , 
    n3765 , 
    n3766 , 
    n3767 , 
    n3768 , 
    n3769 , 
    n3770 , 
    n3771 , 
    n3772 , 
    n3773 , 
    n3774 , 
    n3775 , 
    n3776 , 
    n3777 , 
    n3778 , 
    n3779 , 
    n3780 , 
    n3781 , 
    n3782 , 
    n3783 , 
    n3784 , 
    n3785 , 
    n3786 , 
    n3787 , 
    n3788 , 
    n3789 , 
    n3790 , 
    n3791 , 
    n3792 , 
    n3793 , 
    n3794 , 
    n3795 , 
    n3796 , 
    n3797 , 
    n3798 , 
    n3799 , 
    n3800 , 
    n3801 , 
    n3802 , 
    n3803 , 
    n3804 , 
    n3805 , 
    n3806 , 
    n3807 , 
    n3808 , 
    n3809 , 
    n3810 , 
    n3811 , 
    n3812 , 
    n3813 , 
    n3814 , 
    n3815 , 
    n3816 , 
    n3817 , 
    n3818 , 
    n3819 , 
    n3820 , 
    n3821 , 
    n3822 , 
    n3823 , 
    n3824 , 
    n3825 , 
    n3826 , 
    n3827 , 
    n3828 , 
    n3829 , 
    n3830 , 
    n3831 , 
    n3832 , 
    n3833 , 
    n3834 , 
    n3835 , 
    n3836 , 
    n3837 , 
    n3838 , 
    n3839 , 
    n3840 , 
    n3841 , 
    n3842 , 
    n3843 , 
    n3844 , 
    n3845 , 
    n3846 , 
    n3847 , 
    n3848 , 
    n3849 , 
    n3850 , 
    n3851 , 
    n3852 , 
    n3853 , 
    n3854 , 
    n3855 , 
    n3856 , 
    n3857 , 
    n3858 , 
    n3859 , 
    n3860 , 
    n3861 , 
    n3862 , 
    n3863 , 
    n3864 , 
    n3865 , 
    n3866 , 
    n3867 , 
    n3868 , 
    n3869 , 
    n3870 , 
    n3871 , 
    n3872 , 
    n3873 , 
    n3874 , 
    n3875 , 
    n3876 , 
    n3877 , 
    n3878 , 
    n3879 , 
    n3880 , 
    n3881 , 
    n3882 , 
    n3883 , 
    n3884 , 
    n3885 , 
    n3886 , 
    n3887 , 
    n3888 , 
    n3889 , 
    n3890 , 
    n3891 , 
    n3892 , 
    n3893 , 
    n3894 , 
    n3895 , 
    n3896 , 
    n3897 , 
    n3898 , 
    n3899 , 
    n3900 , 
    n3901 , 
    n3902 , 
    n3903 , 
    n3904 , 
    n3905 , 
    n3906 , 
    n3907 , 
    n3908 , 
    n3909 , 
    n3910 , 
    n3911 , 
    n3912 , 
    n3913 , 
    n3914 , 
    n3915 , 
    n3916 , 
    n3917 , 
    n3918 , 
    n3919 , 
    n3920 , 
    n3921 , 
    n3922 , 
    n3923 , 
    n3924 , 
    n3925 , 
    n3926 , 
    n3927 , 
    n3928 , 
    n3929 , 
    n3930 , 
    n3931 , 
    n3932 , 
    n3933 , 
    n3934 , 
    n3935 , 
    n3936 , 
    n3937 , 
    n3938 , 
    n3939 , 
    n3940 , 
    n3941 , 
    n3942 , 
    n3943 , 
    n3944 , 
    n3945 , 
    n3946 , 
    n3947 , 
    n3948 , 
    n3949 , 
    n3950 , 
    n3951 , 
    n3952 , 
    n3953 , 
    n3954 , 
    n3955 , 
    n3956 , 
    n3957 , 
    n3958 , 
    n3959 , 
    n3960 , 
    n3961 , 
    n3962 , 
    n3963 , 
    n3964 , 
    n3965 , 
    n3966 , 
    n3967 , 
    n3968 , 
    n3969 , 
    n3970 , 
    n3971 , 
    n3972 , 
    n3973 , 
    n3974 , 
    n3975 , 
    n3976 , 
    n3977 , 
    n3978 , 
    n3979 , 
    n3980 , 
    n3981 , 
    n3982 , 
    n3983 , 
    n3984 , 
    n3985 , 
    n3986 , 
    n3987 , 
    n3988 , 
    n3989 , 
    n3990 , 
    n3991 , 
    n3992 , 
    n3993 , 
    n3994 , 
    n3995 , 
    n3996 , 
    n3997 , 
    n3998 , 
    n3999 , 
    n4000 , 
    n4001 , 
    n4002 , 
    n4003 , 
    n4004 , 
    n4005 , 
    n4006 , 
    n4007 , 
    n4008 , 
    n4009 , 
    n4010 , 
    n4011 , 
    n4012 , 
    n4013 , 
    n4014 , 
    n4015 , 
    n4016 , 
    n4017 , 
    n4018 , 
    n4019 , 
    n4020 , 
    n4021 , 
    n4022 , 
    n4023 , 
    n4024 , 
    n4025 , 
    n4026 , 
    n4027 , 
    n4028 , 
    n4029 , 
    n4030 , 
    n4031 , 
    n4032 , 
    n4033 , 
    n4034 , 
    n4035 , 
    n4036 , 
    n4037 , 
    n4038 , 
    n4039 , 
    n4040 , 
    n4041 , 
    n4042 , 
    n4043 , 
    n4044 , 
    n4045 , 
    n4046 , 
    n4047 , 
    n4048 , 
    n4049 , 
    n4050 , 
    n4051 , 
    n4052 , 
    n4053 , 
    n4054 , 
    n4055 , 
    n4056 , 
    n4057 , 
    n4058 , 
    n4059 , 
    n4060 , 
    n4061 , 
    n4062 , 
    n4063 , 
    n4064 , 
    n4065 , 
    n4066 , 
    n4067 , 
    n4068 , 
    n4069 , 
    n4070 , 
    n4071 , 
    n4072 , 
    n4073 , 
    n4074 , 
    n4075 , 
    n4076 , 
    n4077 , 
    n4078 , 
    n4079 , 
    n4080 , 
    n4081 , 
    n4082 , 
    n4083 , 
    n4084 , 
    n4085 , 
    n4086 , 
    n4087 , 
    n4088 , 
    n4089 , 
    n4090 , 
    n4091 , 
    n4092 , 
    n4093 , 
    n4094 , 
    n4095 , 
    n4096 , 
    n4097 , 
    n4098 , 
    n4099 , 
    n4100 , 
    n4101 , 
    n4102 , 
    n4103 , 
    n4104 , 
    n4105 , 
    n4106 , 
    n4107 , 
    n4108 , 
    n4109 , 
    n4110 , 
    n4111 , 
    n4112 , 
    n4113 , 
    n4114 , 
    n4115 , 
    n4116 , 
    n4117 , 
    n4118 , 
    n4119 , 
    n4120 , 
    n4121 , 
    n4122 , 
    n4123 , 
    n4124 , 
    n4125 , 
    n4126 , 
    n4127 , 
    n4128 , 
    n4129 , 
    n4130 , 
    n4131 , 
    n4132 , 
    n4133 , 
    n4134 , 
    n4135 , 
    n4136 , 
    n4137 , 
    n4138 , 
    n4139 , 
    n4140 , 
    n4141 , 
    n4142 , 
    n4143 , 
    n4144 , 
    n4145 , 
    n4146 , 
    n4147 , 
    n4148 , 
    n4149 , 
    n4150 , 
    n4151 , 
    n4152 , 
    n4153 , 
    n4154 , 
    n4155 , 
    n4156 , 
    n4157 , 
    n4158 , 
    n4159 , 
    n4160 , 
    n4161 , 
    n4162 , 
    n4163 , 
    n4164 , 
    n4165 , 
    n4166 , 
    n4167 , 
    n4168 , 
    n4169 , 
    n4170 , 
    n4171 , 
    n4172 , 
    n4173 , 
    n4174 , 
    n4175 , 
    n4176 , 
    n4177 , 
    n4178 , 
    n4179 , 
    n4180 , 
    n4181 , 
    n4182 , 
    n4183 , 
    n4184 , 
    n4185 , 
    n4186 , 
    n4187 , 
    n4188 , 
    n4189 , 
    n4190 , 
    n4191 , 
    n4192 , 
    n4193 , 
    n4194 , 
    n4195 , 
    n4196 , 
    n4197 , 
    n4198 , 
    n4199 , 
    n4200 , 
    n4201 , 
    n4202 , 
    n4203 , 
    n4204 , 
    n4205 , 
    n4206 , 
    n4207 , 
    n4208 , 
    n4209 , 
    n4210 , 
    n4211 , 
    n4212 , 
    n4213 , 
    n4214 , 
    n4215 , 
    n4216 , 
    n4217 , 
    n4218 , 
    n4219 , 
    n4220 , 
    n4221 , 
    n4222 , 
    n4223 , 
    n4224 , 
    n4225 , 
    n4226 , 
    n4227 , 
    n4228 , 
    n4229 , 
    n4230 , 
    n4231 , 
    n4232 , 
    n4233 , 
    n4234 , 
    n4235 , 
    n4236 , 
    n4237 , 
    n4238 , 
    n4239 , 
    n4240 , 
    n4241 , 
    n4242 , 
    n4243 , 
    n4244 , 
    n4245 , 
    n4246 , 
    n4247 , 
    n4248 , 
    n4249 , 
    n4250 , 
    n4251 , 
    n4252 , 
    n4253 , 
    n4254 , 
    n4255 , 
    n4256 , 
    n4257 , 
    n4258 , 
    n4259 , 
    n4260 , 
    n4261 , 
    n4262 , 
    n4263 , 
    n4264 , 
    n4265 , 
    n4266 , 
    n4267 , 
    n4268 , 
    n4269 , 
    n4270 , 
    n4271 , 
    n4272 , 
    n4273 , 
    n4274 , 
    n4275 , 
    n4276 , 
    n4277 , 
    n4278 , 
    n4279 , 
    n4280 , 
    n4281 , 
    n4282 , 
    n4283 , 
    n4284 , 
    n4285 , 
    n4286 , 
    n4287 , 
    n4288 , 
    n4289 , 
    n4290 , 
    n4291 , 
    n4292 , 
    n4293 , 
    n4294 , 
    n4295 , 
    n4296 , 
    n4297 , 
    n4298 , 
    n4299 , 
    n4300 , 
    n4301 , 
    n4302 , 
    n4303 , 
    n4304 , 
    n4305 , 
    n4306 , 
    n4307 , 
    n4308 , 
    n4309 , 
    n4310 , 
    n4311 , 
    n4312 , 
    n4313 , 
    n4314 , 
    n4315 , 
    n4316 , 
    n4317 , 
    n4318 , 
    n4319 , 
    n4320 , 
    n4321 , 
    n4322 , 
    n4323 , 
    n4324 , 
    n4325 , 
    n4326 , 
    n4327 , 
    n4328 , 
    n4329 , 
    n4330 , 
    n4331 , 
    n4332 , 
    n4333 , 
    n4334 , 
    n4335 , 
    n4336 , 
    n4337 , 
    n4338 , 
    n4339 , 
    n4340 , 
    n4341 , 
    n4342 , 
    n4343 , 
    n4344 , 
    n4345 , 
    n4346 , 
    n4347 , 
    n4348 , 
    n4349 , 
    n4350 , 
    n4351 , 
    n4352 , 
    n4353 , 
    n4354 , 
    n4355 , 
    n4356 , 
    n4357 , 
    n4358 , 
    n4359 , 
    n4360 , 
    n4361 , 
    n4362 , 
    n4363 , 
    n4364 , 
    n4365 , 
    n4366 , 
    n4367 , 
    n4368 , 
    n4369 , 
    n4370 , 
    n4371 , 
    n4372 , 
    n4373 , 
    n4374 , 
    n4375 , 
    n4376 , 
    n4377 , 
    n4378 , 
    n4379 , 
    n4380 , 
    n4381 , 
    n4382 , 
    n4383 , 
    n4384 , 
    n4385 , 
    n4386 , 
    n4387 , 
    n4388 , 
    n4389 , 
    n4390 , 
    n4391 , 
    n4392 , 
    n4393 , 
    n4394 , 
    n4395 , 
    n4396 , 
    n4397 , 
    n4398 , 
    n4399 , 
    n4400 , 
    n4401 , 
    n4402 , 
    n4403 , 
    n4404 , 
    n4405 , 
    n4406 , 
    n4407 , 
    n4408 , 
    n4409 , 
    n4410 , 
    n4411 , 
    n4412 , 
    n4413 , 
    n4414 , 
    n4415 , 
    n4416 , 
    n4417 , 
    n4418 , 
    n4419 , 
    n4420 , 
    n4421 , 
    n4422 , 
    n4423 , 
    n4424 , 
    n4425 , 
    n4426 , 
    n4427 , 
    n4428 , 
    n4429 , 
    n4430 , 
    n4431 , 
    n4432 , 
    n4433 , 
    n4434 , 
    n4435 , 
    n4436 , 
    n4437 , 
    n4438 , 
    n4439 , 
    n4440 , 
    n4441 , 
    n4442 , 
    n4443 , 
    n4444 , 
    n4445 , 
    n4446 , 
    n4447 , 
    n4448 , 
    n4449 , 
    n4450 , 
    n4451 , 
    n4452 , 
    n4453 , 
    n4454 , 
    n4455 , 
    n4456 , 
    n4457 , 
    n4458 , 
    n4459 , 
    n4460 , 
    n4461 , 
    n4462 , 
    n4463 , 
    n4464 , 
    n4465 , 
    n4466 , 
    n4467 , 
    n4468 , 
    n4469 , 
    n4470 , 
    n4471 , 
    n4472 , 
    n4473 , 
    n4474 , 
    n4475 , 
    n4476 , 
    n4477 , 
    n4478 , 
    n4479 , 
    n4480 , 
    n4481 , 
    n4482 , 
    n4483 , 
    n4484 , 
    n4485 , 
    n4486 , 
    n4487 , 
    n4488 , 
    n4489 , 
    n4490 , 
    n4491 , 
    n4492 , 
    n4493 , 
    n4494 , 
    n4495 , 
    n4496 , 
    n4497 , 
    n4498 , 
    n4499 , 
    n4500 , 
    n4501 , 
    n4502 , 
    n4503 , 
    n4504 , 
    n4505 , 
    n4506 , 
    n4507 , 
    n4508 , 
    n4509 , 
    n4510 , 
    n4511 , 
    n4512 , 
    n4513 , 
    n4514 , 
    n4515 , 
    n4516 , 
    n4517 , 
    n4518 , 
    n4519 , 
    n4520 , 
    n4521 , 
    n4522 , 
    n4523 , 
    n4524 , 
    n4525 , 
    n4526 , 
    n4527 , 
    n4528 , 
    n4529 , 
    n4530 , 
    n4531 , 
    n4532 , 
    n4533 , 
    n4534 , 
    n4535 , 
    n4536 , 
    n4537 , 
    n4538 , 
    n4539 , 
    n4540 , 
    n4541 , 
    n4542 , 
    n4543 , 
    n4544 , 
    n4545 , 
    n4546 , 
    n4547 , 
    n4548 , 
    n4549 , 
    n4550 , 
    n4551 , 
    n4552 , 
    n4553 , 
    n4554 , 
    n4555 , 
    n4556 , 
    n4557 , 
    n4558 , 
    n4559 , 
    n4560 , 
    n4561 , 
    n4562 , 
    n4563 , 
    n4564 , 
    n4565 , 
    n4566 , 
    n4567 , 
    n4568 , 
    n4569 , 
    n4570 , 
    n4571 , 
    n4572 , 
    n4573 , 
    n4574 , 
    n4575 , 
    n4576 , 
    n4577 , 
    n4578 , 
    n4579 , 
    n4580 , 
    n4581 , 
    n4582 , 
    n4583 , 
    n4584 , 
    n4585 , 
    n4586 , 
    n4587 , 
    n4588 , 
    n4589 , 
    n4590 , 
    n4591 , 
    n4592 , 
    n4593 , 
    n4594 , 
    n4595 , 
    n4596 , 
    n4597 , 
    n4598 , 
    n4599 , 
    n4600 , 
    n4601 , 
    n4602 , 
    n4603 , 
    n4604 , 
    n4605 , 
    n4606 , 
    n4607 , 
    n4608 , 
    n4609 , 
    n4610 , 
    n4611 , 
    n4612 , 
    n4613 , 
    n4614 , 
    n4615 , 
    n4616 , 
    n4617 , 
    n4618 , 
    n4619 , 
    n4620 , 
    n4621 , 
    n4622 , 
    n4623 , 
    n4624 , 
    n4625 , 
    n4626 , 
    n4627 , 
    n4628 , 
    n4629 , 
    n4630 , 
    n4631 , 
    n4632 , 
    n4633 , 
    n4634 , 
    n4635 , 
    n4636 , 
    n4637 , 
    n4638 , 
    n4639 , 
    n4640 , 
    n4641 , 
    n4642 , 
    n4643 , 
    n4644 , 
    n4645 , 
    n4646 , 
    n4647 , 
    n4648 , 
    n4649 , 
    n4650 , 
    n4651 , 
    n4652 , 
    n4653 , 
    n4654 , 
    n4655 , 
    n4656 , 
    n4657 , 
    n4658 , 
    n4659 , 
    n4660 , 
    n4661 , 
    n4662 , 
    n4663 , 
    n4664 , 
    n4665 , 
    n4666 , 
    n4667 , 
    n4668 , 
    n4669 , 
    n4670 , 
    n4671 , 
    n4672 , 
    n4673 , 
    n4674 , 
    n4675 , 
    n4676 , 
    n4677 , 
    n4678 , 
    n4679 , 
    n4680 , 
    n4681 , 
    n4682 , 
    n4683 , 
    n4684 , 
    n4685 , 
    n4686 , 
    n4687 , 
    n4688 , 
    n4689 , 
    n4690 , 
    n4691 , 
    n4692 , 
    n4693 , 
    n4694 , 
    n4695 , 
    n4696 , 
    n4697 , 
    n4698 , 
    n4699 , 
    n4700 , 
    n4701 , 
    n4702 , 
    n4703 , 
    n4704 , 
    n4705 , 
    n4706 , 
    n4707 , 
    n4708 , 
    n4709 , 
    n4710 , 
    n4711 , 
    n4712 , 
    n4713 , 
    n4714 , 
    n4715 , 
    n4716 , 
    n4717 , 
    n4718 , 
    n4719 , 
    n4720 , 
    n4721 , 
    n4722 , 
    n4723 , 
    n4724 , 
    n4725 , 
    n4726 , 
    n4727 , 
    n4728 , 
    n4729 , 
    n4730 , 
    n4731 , 
    n4732 , 
    n4733 , 
    n4734 , 
    n4735 , 
    n4736 , 
    n4737 , 
    n4738 , 
    n4739 , 
    n4740 , 
    n4741 , 
    n4742 , 
    n4743 , 
    n4744 , 
    n4745 , 
    n4746 , 
    n4747 , 
    n4748 , 
    n4749 , 
    n4750 , 
    n4751 , 
    n4752 , 
    n4753 , 
    n4754 , 
    n4755 , 
    n4756 , 
    n4757 , 
    n4758 , 
    n4759 , 
    n4760 , 
    n4761 , 
    n4762 , 
    n4763 , 
    n4764 , 
    n4765 , 
    n4766 , 
    n4767 , 
    n4768 , 
    n4769 , 
    n4770 , 
    n4771 , 
    n4772 , 
    n4773 , 
    n4774 , 
    n4775 , 
    n4776 , 
    n4777 , 
    n4778 , 
    n4779 , 
    n4780 , 
    n4781 , 
    n4782 , 
    n4783 , 
    n4784 , 
    n4785 , 
    n4786 , 
    n4787 , 
    n4788 , 
    n4789 , 
    n4790 , 
    n4791 , 
    n4792 , 
    n4793 , 
    n4794 , 
    n4795 , 
    n4796 , 
    n4797 , 
    n4798 , 
    n4799 , 
    n4800 , 
    n4801 , 
    n4802 , 
    n4803 , 
    n4804 , 
    n4805 , 
    n4806 , 
    n4807 , 
    n4808 , 
    n4809 , 
    n4810 , 
    n4811 , 
    n4812 , 
    n4813 , 
    n4814 , 
    n4815 , 
    n4816 , 
    n4817 , 
    n4818 , 
    n4819 , 
    n4820 , 
    n4821 , 
    n4822 , 
    n4823 , 
    n4824 , 
    n4825 , 
    n4826 , 
    n4827 , 
    n4828 , 
    n4829 , 
    n4830 , 
    n4831 , 
    n4832 , 
    n4833 , 
    n4834 , 
    n4835 , 
    n4836 , 
    n4837 , 
    n4838 , 
    n4839 , 
    n4840 , 
    n4841 , 
    n4842 , 
    n4843 , 
    n4844 , 
    n4845 , 
    n4846 , 
    n4847 , 
    n4848 , 
    n4849 , 
    n4850 , 
    n4851 , 
    n4852 , 
    n4853 , 
    n4854 , 
    n4855 , 
    n4856 , 
    n4857 , 
    n4858 , 
    n4859 , 
    n4860 , 
    n4861 , 
    n4862 , 
    n4863 , 
    n4864 , 
    n4865 , 
    n4866 , 
    n4867 , 
    n4868 , 
    n4869 , 
    n4870 , 
    n4871 , 
    n4872 , 
    n4873 , 
    n4874 , 
    n4875 , 
    n4876 , 
    n4877 , 
    n4878 , 
    n4879 , 
    n4880 , 
    n4881 , 
    n4882 , 
    n4883 , 
    n4884 , 
    n4885 , 
    n4886 , 
    n4887 , 
    n4888 , 
    n4889 , 
    n4890 , 
    n4891 , 
    n4892 , 
    n4893 , 
    n4894 , 
    n4895 , 
    n4896 , 
    n4897 , 
    n4898 , 
    n4899 , 
    n4900 , 
    n4901 , 
    n4902 , 
    n4903 , 
    n4904 , 
    n4905 , 
    n4906 , 
    n4907 , 
    n4908 , 
    n4909 , 
    n4910 , 
    n4911 , 
    n4912 , 
    n4913 , 
    n4914 , 
    n4915 , 
    n4916 , 
    n4917 , 
    n4918 , 
    n4919 , 
    n4920 , 
    n4921 , 
    n4922 , 
    n4923 , 
    n4924 , 
    n4925 , 
    n4926 , 
    n4927 , 
    n4928 , 
    n4929 , 
    n4930 , 
    n4931 , 
    n4932 , 
    n4933 , 
    n4934 , 
    n4935 , 
    n4936 , 
    n4937 , 
    n4938 , 
    n4939 , 
    n4940 , 
    n4941 , 
    n4942 , 
    n4943 , 
    n4944 , 
    n4945 , 
    n4946 , 
    n4947 , 
    n4948 , 
    n4949 , 
    n4950 , 
    n4951 , 
    n4952 , 
    n4953 , 
    n4954 , 
    n4955 , 
    n4956 , 
    n4957 , 
    n4958 , 
    n4959 , 
    n4960 , 
    n4961 , 
    n4962 , 
    n4963 , 
    n4964 , 
    n4965 , 
    n4966 , 
    n4967 , 
    n4968 , 
    n4969 , 
    n4970 , 
    n4971 , 
    n4972 , 
    n4973 , 
    n4974 , 
    n4975 , 
    n4976 , 
    n4977 , 
    n4978 , 
    n4979 , 
    n4980 , 
    n4981 , 
    n4982 , 
    n4983 , 
    n4984 , 
    n4985 , 
    n4986 , 
    n4987 , 
    n4988 , 
    n4989 , 
    n4990 , 
    n4991 , 
    n4992 , 
    n4993 , 
    n4994 , 
    n4995 , 
    n4996 , 
    n4997 , 
    n4998 , 
    n4999 , 
    n5000 , 
    n5001 , 
    n5002 , 
    n5003 , 
    n5004 , 
    n5005 , 
    n5006 , 
    n5007 , 
    n5008 , 
    n5009 , 
    n5010 , 
    n5011 , 
    n5012 , 
    n5013 , 
    n5014 , 
    n5015 , 
    n5016 , 
    n5017 , 
    n5018 , 
    n5019 , 
    n5020 , 
    n5021 , 
    n5022 , 
    n5023 , 
    n5024 , 
    n5025 , 
    n5026 , 
    n5027 , 
    n5028 , 
    n5029 , 
    n5030 , 
    n5031 , 
    n5032 , 
    n5033 , 
    n5034 , 
    n5035 , 
    n5036 , 
    n5037 , 
    n5038 , 
    n5039 , 
    n5040 , 
    n5041 , 
    n5042 , 
    n5043 , 
    n5044 , 
    n5045 , 
    n5046 , 
    n5047 , 
    n5048 , 
    n5049 , 
    n5050 , 
    n5051 , 
    n5052 , 
    n5053 , 
    n5054 , 
    n5055 , 
    n5056 , 
    n5057 , 
    n5058 , 
    n5059 , 
    n5060 , 
    n5061 , 
    n5062 , 
    n5063 , 
    n5064 , 
    n5065 , 
    n5066 , 
    n5067 , 
    n5068 , 
    n5069 , 
    n5070 , 
    n5071 , 
    n5072 , 
    n5073 , 
    n5074 , 
    n5075 , 
    n5076 , 
    n5077 , 
    n5078 , 
    n5079 , 
    n5080 , 
    n5081 , 
    n5082 , 
    n5083 , 
    n5084 , 
    n5085 , 
    n5086 , 
    n5087 , 
    n5088 , 
    n5089 , 
    n5090 , 
    n5091 , 
    n5092 , 
    n5093 , 
    n5094 , 
    n5095 , 
    n5096 , 
    n5097 , 
    n5098 , 
    n5099 , 
    n5100 , 
    n5101 , 
    n5102 , 
    n5103 , 
    n5104 , 
    n5105 , 
    n5106 , 
    n5107 , 
    n5108 , 
    n5109 , 
    n5110 , 
    n5111 , 
    n5112 , 
    n5113 , 
    n5114 , 
    n5115 , 
    n5116 , 
    n5117 , 
    n5118 , 
    n5119 , 
    n5120 , 
    n5121 , 
    n5122 , 
    n5123 , 
    n5124 , 
    n5125 , 
    n5126 , 
    n5127 , 
    n5128 , 
    n5129 , 
    n5130 , 
    n5131 , 
    n5132 , 
    n5133 , 
    n5134 , 
    n5135 , 
    n5136 , 
    n5137 , 
    n5138 , 
    n5139 , 
    n5140 , 
    n5141 , 
    n5142 , 
    n5143 , 
    n5144 , 
    n5145 , 
    n5146 , 
    n5147 , 
    n5148 , 
    n5149 , 
    n5150 , 
    n5151 , 
    n5152 , 
    n5153 , 
    n5154 , 
    n5155 , 
    n5156 , 
    n5157 , 
    n5158 , 
    n5159 , 
    n5160 , 
    n5161 , 
    n5162 , 
    n5163 , 
    n5164 , 
    n5165 , 
    n5166 , 
    n5167 , 
    n5168 , 
    n5169 , 
    n5170 , 
    n5171 , 
    n5172 , 
    n5173 , 
    n5174 , 
    n5175 , 
    n5176 , 
    n5177 , 
    n5178 , 
    n5179 , 
    n5180 , 
    n5181 , 
    n5182 , 
    n5183 , 
    n5184 , 
    n5185 , 
    n5186 , 
    n5187 , 
    n5188 , 
    n5189 , 
    n5190 , 
    n5191 , 
    n5192 , 
    n5193 , 
    n5194 , 
    n5195 , 
    n5196 , 
    n5197 , 
    n5198 , 
    n5199 , 
    n5200 , 
    n5201 , 
    n5202 , 
    n5203 , 
    n5204 , 
    n5205 , 
    n5206 , 
    n5207 , 
    n5208 , 
    n5209 , 
    n5210 , 
    n5211 , 
    n5212 , 
    n5213 , 
    n5214 , 
    n5215 , 
    n5216 , 
    n5217 , 
    n5218 , 
    n5219 , 
    n5220 , 
    n5221 , 
    n5222 , 
    n5223 , 
    n5224 , 
    n5225 , 
    n5226 , 
    n5227 , 
    n5228 , 
    n5229 , 
    n5230 , 
    n5231 , 
    n5232 , 
    n5233 , 
    n5234 , 
    n5235 , 
    n5236 , 
    n5237 , 
    n5238 , 
    n5239 , 
    n5240 , 
    n5241 , 
    n5242 , 
    n5243 , 
    n5244 , 
    n5245 , 
    n5246 , 
    n5247 , 
    n5248 , 
    n5249 , 
    n5250 , 
    n5251 , 
    n5252 , 
    n5253 , 
    n5254 , 
    n5255 , 
    n5256 , 
    n5257 , 
    n5258 , 
    n5259 , 
    n5260 , 
    n5261 , 
    n5262 , 
    n5263 , 
    n5264 , 
    n5265 , 
    n5266 , 
    n5267 , 
    n5268 , 
    n5269 , 
    n5270 , 
    n5271 , 
    n5272 , 
    n5273 , 
    n5274 , 
    n5275 , 
    n5276 , 
    n5277 , 
    n5278 , 
    n5279 , 
    n5280 , 
    n5281 , 
    n5282 , 
    n5283 , 
    n5284 , 
    n5285 , 
    n5286 , 
    n5287 , 
    n5288 , 
    n5289 , 
    n5290 , 
    n5291 , 
    n5292 , 
    n5293 , 
    n5294 , 
    n5295 , 
    n5296 , 
    n5297 , 
    n5298 , 
    n5299 , 
    n5300 , 
    n5301 , 
    n5302 , 
    n5303 , 
    n5304 , 
    n5305 , 
    n5306 , 
    n5307 , 
    n5308 , 
    n5309 , 
    n5310 , 
    n5311 , 
    n5312 , 
    n5313 , 
    n5314 , 
    n5315 , 
    n5316 , 
    n5317 , 
    n5318 , 
    n5319 , 
    n5320 , 
    n5321 , 
    n5322 , 
    n5323 , 
    n5324 , 
    n5325 , 
    n5326 , 
    n5327 , 
    n5328 , 
    n5329 , 
    n5330 , 
    n5331 , 
    n5332 , 
    n5333 , 
    n5334 , 
    n5335 , 
    n5336 , 
    n5337 , 
    n5338 , 
    n5339 , 
    n5340 , 
    n5341 , 
    n5342 , 
    n5343 , 
    n5344 , 
    n5345 , 
    n5346 , 
    n5347 , 
    n5348 , 
    n5349 , 
    n5350 , 
    n5351 , 
    n5352 , 
    n5353 , 
    n5354 , 
    n5355 , 
    n5356 , 
    n5357 , 
    n5358 , 
    n5359 , 
    n5360 , 
    n5361 , 
    n5362 , 
    n5363 , 
    n5364 , 
    n5365 , 
    n5366 , 
    n5367 , 
    n5368 , 
    n5369 , 
    n5370 , 
    n5371 , 
    n5372 , 
    n5373 , 
    n5374 , 
    n5375 , 
    n5376 , 
    n5377 , 
    n5378 , 
    n5379 , 
    n5380 , 
    n5381 , 
    n5382 , 
    n5383 , 
    n5384 , 
    n5385 , 
    n5386 , 
    n5387 , 
    n5388 , 
    n5389 , 
    n5390 , 
    n5391 , 
    n5392 , 
    n5393 , 
    n5394 , 
    n5395 , 
    n5396 , 
    n5397 , 
    n5398 , 
    n5399 , 
    n5400 , 
    n5401 , 
    n5402 , 
    n5403 , 
    n5404 , 
    n5405 , 
    n5406 , 
    n5407 , 
    n5408 , 
    n5409 , 
    n5410 , 
    n5411 , 
    n5412 , 
    n5413 , 
    n5414 , 
    n5415 , 
    n5416 , 
    n5417 , 
    n5418 , 
    n5419 , 
    n5420 , 
    n5421 , 
    n5422 , 
    n5423 , 
    n5424 , 
    n5425 , 
    n5426 , 
    n5427 , 
    n5428 , 
    n5429 , 
    n5430 , 
    n5431 , 
    n5432 , 
    n5433 , 
    n5434 , 
    n5435 , 
    n5436 , 
    n5437 , 
    n5438 , 
    n5439 , 
    n5440 , 
    n5441 , 
    n5442 , 
    n5443 , 
    n5444 , 
    n5445 , 
    n5446 , 
    n5447 , 
    n5448 , 
    n5449 , 
    n5450 , 
    n5451 , 
    n5452 , 
    n5453 , 
    n5454 , 
    n5455 , 
    n5456 , 
    n5457 , 
    n5458 , 
    n5459 , 
    n5460 , 
    n5461 , 
    n5462 , 
    n5463 , 
    n5464 , 
    n5465 , 
    n5466 , 
    n5467 , 
    n5468 , 
    n5469 , 
    n5470 , 
    n5471 , 
    n5472 , 
    n5473 , 
    n5474 , 
    n5475 , 
    n5476 , 
    n5477 , 
    n5478 , 
    n5479 , 
    n5480 , 
    n5481 , 
    n5482 , 
    n5483 , 
    n5484 , 
    n5485 , 
    n5486 , 
    n5487 , 
    n5488 , 
    n5489 , 
    n5490 , 
    n5491 , 
    n5492 , 
    n5493 , 
    n5494 , 
    n5495 , 
    n5496 , 
    n5497 , 
    n5498 , 
    n5499 , 
    n5500 , 
    n5501 , 
    n5502 , 
    n5503 , 
    n5504 , 
    n5505 , 
    n5506 , 
    n5507 , 
    n5508 , 
    n5509 , 
    n5510 , 
    n5511 , 
    n5512 , 
    n5513 , 
    n5514 , 
    n5515 , 
    n5516 , 
    n5517 , 
    n5518 , 
    n5519 , 
    n5520 , 
    n5521 , 
    n5522 , 
    n5523 , 
    n5524 , 
    n5525 , 
    n5526 , 
    n5527 , 
    n5528 , 
    n5529 , 
    n5530 , 
    n5531 , 
    n5532 , 
    n5533 , 
    n5534 , 
    n5535 , 
    n5536 , 
    n5537 , 
    n5538 , 
    n5539 , 
    n5540 , 
    n5541 , 
    n5542 , 
    n5543 , 
    n5544 , 
    n5545 , 
    n5546 , 
    n5547 , 
    n5548 , 
    n5549 , 
    n5550 , 
    n5551 , 
    n5552 , 
    n5553 , 
    n5554 , 
    n5555 , 
    n5556 , 
    n5557 , 
    n5558 , 
    n5559 , 
    n5560 , 
    n5561 , 
    n5562 , 
    n5563 , 
    n5564 , 
    n5565 , 
    n5566 , 
    n5567 , 
    n5568 , 
    n5569 , 
    n5570 , 
    n5571 , 
    n5572 , 
    n5573 , 
    n5574 , 
    n5575 , 
    n5576 , 
    n5577 , 
    n5578 , 
    n5579 , 
    n5580 , 
    n5581 , 
    n5582 , 
    n5583 , 
    n5584 , 
    n5585 , 
    n5586 , 
    n5587 , 
    n5588 , 
    n5589 , 
    n5590 , 
    n5591 , 
    n5592 , 
    n5593 , 
    n5594 , 
    n5595 , 
    n5596 , 
    n5597 , 
    n5598 , 
    n5599 , 
    n5600 , 
    n5601 , 
    n5602 , 
    n5603 , 
    n5604 , 
    n5605 , 
    n5606 , 
    n5607 , 
    n5608 , 
    n5609 , 
    n5610 , 
    n5611 , 
    n5612 , 
    n5613 , 
    n5614 , 
    n5615 , 
    n5616 , 
    n5617 , 
    n5618 , 
    n5619 , 
    n5620 , 
    n5621 , 
    n5622 , 
    n5623 , 
    n5624 , 
    n5625 , 
    n5626 , 
    n5627 , 
    n5628 , 
    n5629 , 
    n5630 , 
    n5631 , 
    n5632 , 
    n5633 , 
    n5634 , 
    n5635 , 
    n5636 , 
    n5637 , 
    n5638 , 
    n5639 , 
    n5640 , 
    n5641 , 
    n5642 , 
    n5643 , 
    n5644 , 
    n5645 , 
    n5646 , 
    n5647 , 
    n5648 , 
    n5649 , 
    n5650 , 
    n5651 , 
    n5652 , 
    n5653 , 
    n5654 , 
    n5655 , 
    n5656 , 
    n5657 , 
    n5658 , 
    n5659 , 
    n5660 , 
    n5661 , 
    n5662 , 
    n5663 , 
    n5664 , 
    n5665 , 
    n5666 , 
    n5667 , 
    n5668 , 
    n5669 , 
    n5670 , 
    n5671 , 
    n5672 , 
    n5673 , 
    n5674 , 
    n5675 , 
    n5676 , 
    n5677 , 
    n5678 , 
    n5679 , 
    n5680 , 
    n5681 , 
    n5682 , 
    n5683 , 
    n5684 , 
    n5685 , 
    n5686 , 
    n5687 , 
    n5688 , 
    n5689 , 
    n5690 , 
    n5691 , 
    n5692 , 
    n5693 , 
    n5694 , 
    n5695 , 
    n5696 , 
    n5697 , 
    n5698 , 
    n5699 , 
    n5700 , 
    n5701 , 
    n5702 , 
    n5703 , 
    n5704 , 
    n5705 , 
    n5706 , 
    n5707 , 
    n5708 , 
    n5709 , 
    n5710 , 
    n5711 , 
    n5712 , 
    n5713 , 
    n5714 , 
    n5715 , 
    n5716 , 
    n5717 , 
    n5718 , 
    n5719 , 
    n5720 , 
    n5721 , 
    n5722 , 
    n5723 , 
    n5724 , 
    n5725 , 
    n5726 , 
    n5727 , 
    n5728 , 
    n5729 , 
    n5730 , 
    n5731 , 
    n5732 , 
    n5733 , 
    n5734 , 
    n5735 , 
    n5736 , 
    n5737 , 
    n5738 , 
    n5739 , 
    n5740 , 
    n5741 , 
    n5742 , 
    n5743 , 
    n5744 , 
    n5745 , 
    n5746 , 
    n5747 , 
    n5748 , 
    n5749 , 
    n5750 , 
    n5751 , 
    n5752 , 
    n5753 , 
    n5754 , 
    n5755 , 
    n5756 , 
    n5757 , 
    n5758 , 
    n5759 , 
    n5760 , 
    n5761 , 
    n5762 , 
    n5763 , 
    n5764 , 
    n5765 , 
    n5766 , 
    n5767 , 
    n5768 , 
    n5769 , 
    n5770 , 
    n5771 , 
    n5772 , 
    n5773 , 
    n5774 , 
    n5775 , 
    n5776 , 
    n5777 , 
    n5778 , 
    n5779 , 
    n5780 , 
    n5781 , 
    n5782 , 
    n5783 , 
    n5784 , 
    n5785 , 
    n5786 , 
    n5787 , 
    n5788 , 
    n5789 , 
    n5790 , 
    n5791 , 
    n5792 , 
    n5793 , 
    n5794 , 
    n5795 , 
    n5796 , 
    n5797 , 
    n5798 , 
    n5799 , 
    n5800 , 
    n5801 , 
    n5802 , 
    n5803 , 
    n5804 , 
    n5805 , 
    n5806 , 
    n5807 , 
    n5808 , 
    n5809 , 
    n5810 , 
    n5811 , 
    n5812 , 
    n5813 , 
    n5814 , 
    n5815 , 
    n5816 , 
    n5817 , 
    n5818 , 
    n5819 , 
    n5820 , 
    n5821 , 
    n5822 , 
    n5823 , 
    n5824 , 
    n5825 , 
    n5826 , 
    n5827 , 
    n5828 , 
    n5829 , 
    n5830 , 
    n5831 , 
    n5832 , 
    n5833 , 
    n5834 , 
    n5835 , 
    n5836 , 
    n5837 , 
    n5838 , 
    n5839 , 
    n5840 , 
    n5841 , 
    n5842 , 
    n5843 , 
    n5844 , 
    n5845 , 
    n5846 , 
    n5847 , 
    n5848 , 
    n5849 , 
    n5850 , 
    n5851 , 
    n5852 , 
    n5853 , 
    n5854 , 
    n5855 , 
    n5856 , 
    n5857 , 
    n5858 , 
    n5859 , 
    n5860 , 
    n5861 , 
    n5862 , 
    n5863 , 
    n5864 , 
    n5865 , 
    n5866 , 
    n5867 , 
    n5868 , 
    n5869 , 
    n5870 , 
    n5871 , 
    n5872 , 
    n5873 , 
    n5874 , 
    n5875 , 
    n5876 , 
    n5877 , 
    n5878 , 
    n5879 , 
    n5880 , 
    n5881 , 
    n5882 , 
    n5883 , 
    n5884 , 
    n5885 , 
    n5886 , 
    n5887 , 
    n5888 , 
    n5889 , 
    n5890 , 
    n5891 , 
    n5892 , 
    n5893 , 
    n5894 , 
    n5895 , 
    n5896 , 
    n5897 , 
    n5898 , 
    n5899 , 
    n5900 , 
    n5901 , 
    n5902 , 
    n5903 , 
    n5904 , 
    n5905 , 
    n5906 , 
    n5907 , 
    n5908 , 
    n5909 , 
    n5910 , 
    n5911 , 
    n5912 , 
    n5913 , 
    n5914 , 
    n5915 , 
    n5916 , 
    n5917 , 
    n5918 , 
    n5919 , 
    n5920 , 
    n5921 , 
    n5922 , 
    n5923 , 
    n5924 , 
    n5925 , 
    n5926 , 
    n5927 , 
    n5928 , 
    n5929 , 
    n5930 , 
    n5931 , 
    n5932 , 
    n5933 , 
    n5934 , 
    n5935 , 
    n5936 , 
    n5937 , 
    n5938 , 
    n5939 , 
    n5940 , 
    n5941 , 
    n5942 , 
    n5943 , 
    n5944 , 
    n5945 , 
    n5946 , 
    n5947 , 
    n5948 , 
    n5949 , 
    n5950 , 
    n5951 , 
    n5952 , 
    n5953 , 
    n5954 , 
    n5955 , 
    n5956 , 
    n5957 , 
    n5958 , 
    n5959 , 
    n5960 , 
    n5961 , 
    n5962 , 
    n5963 , 
    n5964 , 
    n5965 , 
    n5966 , 
    n5967 , 
    n5968 , 
    n5969 , 
    n5970 , 
    n5971 , 
    n5972 , 
    n5973 , 
    n5974 , 
    n5975 , 
    n5976 , 
    n5977 , 
    n5978 , 
    n5979 , 
    n5980 , 
    n5981 , 
    n5982 , 
    n5983 , 
    n5984 , 
    n5985 , 
    n5986 , 
    n5987 , 
    n5988 , 
    n5989 , 
    n5990 , 
    n5991 , 
    n5992 , 
    n5993 , 
    n5994 , 
    n5995 , 
    n5996 , 
    n5997 , 
    n5998 , 
    n5999 , 
    n6000 , 
    n6001 , 
    n6002 , 
    n6003 , 
    n6004 , 
    n6005 , 
    n6006 , 
    n6007 , 
    n6008 , 
    n6009 , 
    n6010 , 
    n6011 , 
    n6012 , 
    n6013 , 
    n6014 , 
    n6015 , 
    n6016 , 
    n6017 , 
    n6018 , 
    n6019 , 
    n6020 , 
    n6021 , 
    n6022 , 
    n6023 , 
    n6024 , 
    n6025 , 
    n6026 , 
    n6027 , 
    n6028 , 
    n6029 , 
    n6030 , 
    n6031 , 
    n6032 , 
    n6033 , 
    n6034 , 
    n6035 , 
    n6036 , 
    n6037 , 
    n6038 , 
    n6039 , 
    n6040 , 
    n6041 , 
    n6042 , 
    n6043 , 
    n6044 , 
    n6045 , 
    n6046 , 
    n6047 , 
    n6048 , 
    n6049 , 
    n6050 , 
    n6051 , 
    n6052 , 
    n6053 , 
    n6054 , 
    n6055 , 
    n6056 , 
    n6057 , 
    n6058 , 
    n6059 , 
    n6060 , 
    n6061 , 
    n6062 , 
    n6063 , 
    n6064 , 
    n6065 , 
    n6066 , 
    n6067 , 
    n6068 , 
    n6069 , 
    n6070 , 
    n6071 , 
    n6072 , 
    n6073 , 
    n6074 , 
    n6075 , 
    n6076 , 
    n6077 , 
    n6078 , 
    n6079 , 
    n6080 , 
    n6081 , 
    n6082 , 
    n6083 , 
    n6084 , 
    n6085 , 
    n6086 , 
    n6087 , 
    n6088 , 
    n6089 , 
    n6090 , 
    n6091 , 
    n6092 , 
    n6093 , 
    n6094 , 
    n6095 , 
    n6096 , 
    n6097 , 
    n6098 , 
    n6099 , 
    n6100 , 
    n6101 , 
    n6102 , 
    n6103 , 
    n6104 , 
    n6105 , 
    n6106 , 
    n6107 , 
    n6108 , 
    n6109 , 
    n6110 , 
    n6111 , 
    n6112 , 
    n6113 , 
    n6114 , 
    n6115 , 
    n6116 , 
    n6117 , 
    n6118 , 
    n6119 , 
    n6120 , 
    n6121 , 
    n6122 , 
    n6123 , 
    n6124 , 
    n6125 , 
    n6126 , 
    n6127 , 
    n6128 , 
    n6129 , 
    n6130 , 
    n6131 , 
    n6132 , 
    n6133 , 
    n6134 , 
    n6135 , 
    n6136 , 
    n6137 , 
    n6138 , 
    n6139 , 
    n6140 , 
    n6141 , 
    n6142 , 
    n6143 , 
    n6144 , 
    n6145 , 
    n6146 , 
    n6147 , 
    n6148 , 
    n6149 , 
    n6150 , 
    n6151 , 
    n6152 , 
    n6153 , 
    n6154 , 
    n6155 , 
    n6156 , 
    n6157 , 
    n6158 , 
    n6159 , 
    n6160 , 
    n6161 , 
    n6162 , 
    n6163 , 
    n6164 , 
    n6165 , 
    n6166 , 
    n6167 , 
    n6168 , 
    n6169 , 
    n6170 , 
    n6171 , 
    n6172 , 
    n6173 , 
    n6174 , 
    n6175 , 
    n6176 , 
    n6177 , 
    n6178 , 
    n6179 , 
    n6180 , 
    n6181 , 
    n6182 , 
    n6183 , 
    n6184 , 
    n6185 , 
    n6186 , 
    n6187 , 
    n6188 , 
    n6189 , 
    n6190 , 
    n6191 , 
    n6192 , 
    n6193 , 
    n6194 , 
    n6195 , 
    n6196 , 
    n6197 , 
    n6198 , 
    n6199 , 
    n6200 , 
    n6201 , 
    n6202 , 
    n6203 , 
    n6204 , 
    n6205 , 
    n6206 , 
    n6207 , 
    n6208 , 
    n6209 , 
    n6210 , 
    n6211 , 
    n6212 , 
    n6213 , 
    n6214 , 
    n6215 , 
    n6216 , 
    n6217 , 
    n6218 , 
    n6219 , 
    n6220 , 
    n6221 , 
    n6222 , 
    n6223 , 
    n6224 , 
    n6225 , 
    n6226 , 
    n6227 , 
    n6228 , 
    n6229 , 
    n6230 , 
    n6231 , 
    n6232 , 
    n6233 , 
    n6234 , 
    n6235 , 
    n6236 , 
    n6237 , 
    n6238 , 
    n6239 , 
    n6240 , 
    n6241 , 
    n6242 , 
    n6243 , 
    n6244 , 
    n6245 , 
    n6246 , 
    n6247 , 
    n6248 , 
    n6249 , 
    n6250 , 
    n6251 , 
    n6252 , 
    n6253 , 
    n6254 , 
    n6255 , 
    n6256 , 
    n6257 , 
    n6258 , 
    n6259 , 
    n6260 , 
    n6261 , 
    n6262 , 
    n6263 , 
    n6264 , 
    n6265 , 
    n6266 , 
    n6267 , 
    n6268 , 
    n6269 , 
    n6270 , 
    n6271 , 
    n6272 , 
    n6273 , 
    n6274 , 
    n6275 , 
    n6276 , 
    n6277 , 
    n6278 , 
    n6279 , 
    n6280 , 
    n6281 , 
    n6282 , 
    n6283 , 
    n6284 , 
    n6285 , 
    n6286 , 
    n6287 , 
    n6288 , 
    n6289 , 
    n6290 , 
    n6291 , 
    n6292 , 
    n6293 , 
    n6294 , 
    n6295 , 
    n6296 , 
    n6297 , 
    n6298 , 
    n6299 , 
    n6300 , 
    n6301 , 
    n6302 , 
    n6303 , 
    n6304 , 
    n6305 , 
    n6306 , 
    n6307 , 
    n6308 , 
    n6309 , 
    n6310 , 
    n6311 , 
    n6312 , 
    n6313 , 
    n6314 , 
    n6315 , 
    n6316 , 
    n6317 , 
    n6318 , 
    n6319 , 
    n6320 , 
    n6321 , 
    n6322 , 
    n6323 , 
    n6324 , 
    n6325 , 
    n6326 , 
    n6327 , 
    n6328 , 
    n6329 , 
    n6330 , 
    n6331 , 
    n6332 , 
    n6333 , 
    n6334 , 
    n6335 , 
    n6336 , 
    n6337 , 
    n6338 , 
    n6339 , 
    n6340 , 
    n6341 , 
    n6342 , 
    n6343 , 
    n6344 , 
    n6345 , 
    n6346 , 
    n6347 , 
    n6348 , 
    n6349 , 
    n6350 , 
    n6351 , 
    n6352 , 
    n6353 , 
    n6354 , 
    n6355 , 
    n6356 , 
    n6357 , 
    n6358 , 
    n6359 , 
    n6360 , 
    n6361 , 
    n6362 , 
    n6363 , 
    n6364 , 
    n6365 , 
    n6366 , 
    n6367 , 
    n6368 , 
    n6369 , 
    n6370 , 
    n6371 , 
    n6372 , 
    n6373 , 
    n6374 , 
    n6375 , 
    n6376 , 
    n6377 , 
    n6378 , 
    n6379 , 
    n6380 , 
    n6381 , 
    n6382 , 
    n6383 , 
    n6384 , 
    n6385 , 
    n6386 , 
    n6387 , 
    n6388 , 
    n6389 , 
    n6390 , 
    n6391 , 
    n6392 , 
    n6393 , 
    n6394 , 
    n6395 , 
    n6396 , 
    n6397 , 
    n6398 , 
    n6399 , 
    n6400 , 
    n6401 , 
    n6402 , 
    n6403 , 
    n6404 , 
    n6405 , 
    n6406 , 
    n6407 , 
    n6408 , 
    n6409 , 
    n6410 , 
    n6411 , 
    n6412 , 
    n6413 , 
    n6414 , 
    n6415 , 
    n6416 , 
    n6417 , 
    n6418 , 
    n6419 , 
    n6420 , 
    n6421 , 
    n6422 , 
    n6423 , 
    n6424 , 
    n6425 , 
    n6426 , 
    n6427 , 
    n6428 , 
    n6429 , 
    n6430 , 
    n6431 , 
    n6432 , 
    n6433 , 
    n6434 , 
    n6435 , 
    n6436 , 
    n6437 , 
    n6438 , 
    n6439 , 
    n6440 , 
    n6441 , 
    n6442 , 
    n6443 , 
    n6444 , 
    n6445 , 
    n6446 , 
    n6447 , 
    n6448 , 
    n6449 , 
    n6450 , 
    n6451 , 
    n6452 , 
    n6453 , 
    n6454 , 
    n6455 , 
    n6456 , 
    n6457 , 
    n6458 , 
    n6459 , 
    n6460 , 
    n6461 , 
    n6462 , 
    n6463 , 
    n6464 , 
    n6465 , 
    n6466 , 
    n6467 , 
    n6468 , 
    n6469 , 
    n6470 , 
    n6471 , 
    n6472 , 
    n6473 , 
    n6474 , 
    n6475 , 
    n6476 , 
    n6477 , 
    n6478 , 
    n6479 , 
    n6480 , 
    n6481 , 
    n6482 , 
    n6483 , 
    n6484 , 
    n6485 , 
    n6486 , 
    n6487 , 
    n6488 , 
    n6489 , 
    n6490 , 
    n6491 , 
    n6492 , 
    n6493 , 
    n6494 , 
    n6495 , 
    n6496 , 
    n6497 , 
    n6498 , 
    n6499 , 
    n6500 , 
    n6501 , 
    n6502 , 
    n6503 , 
    n6504 , 
    n6505 , 
    n6506 , 
    n6507 , 
    n6508 , 
    n6509 , 
    n6510 , 
    n6511 , 
    n6512 , 
    n6513 , 
    n6514 , 
    n6515 , 
    n6516 , 
    n6517 , 
    n6518 , 
    n6519 , 
    n6520 , 
    n6521 , 
    n6522 , 
    n6523 , 
    n6524 , 
    n6525 , 
    n6526 , 
    n6527 , 
    n6528 , 
    n6529 , 
    n6530 , 
    n6531 , 
    n6532 , 
    n6533 , 
    n6534 , 
    n6535 , 
    n6536 , 
    n6537 , 
    n6538 , 
    n6539 , 
    n6540 , 
    n6541 , 
    n6542 , 
    n6543 , 
    n6544 , 
    n6545 , 
    n6546 , 
    n6547 , 
    n6548 , 
    n6549 , 
    n6550 , 
    n6551 , 
    n6552 , 
    n6553 , 
    n6554 , 
    n6555 , 
    n6556 , 
    n6557 , 
    n6558 , 
    n6559 , 
    n6560 , 
    n6561 , 
    n6562 , 
    n6563 , 
    n6564 , 
    n6565 , 
    n6566 , 
    n6567 , 
    n6568 , 
    n6569 , 
    n6570 , 
    n6571 , 
    n6572 , 
    n6573 , 
    n6574 , 
    n6575 , 
    n6576 , 
    n6577 , 
    n6578 , 
    n6579 , 
    n6580 , 
    n6581 , 
    n6582 , 
    n6583 , 
    n6584 , 
    n6585 , 
    n6586 , 
    n6587 , 
    n6588 , 
    n6589 , 
    n6590 , 
    n6591 , 
    n6592 , 
    n6593 , 
    n6594 , 
    n6595 , 
    n6596 , 
    n6597 , 
    n6598 , 
    n6599 , 
    n6600 , 
    n6601 , 
    n6602 , 
    n6603 , 
    n6604 , 
    n6605 , 
    n6606 , 
    n6607 , 
    n6608 , 
    n6609 , 
    n6610 , 
    n6611 , 
    n6612 , 
    n6613 , 
    n6614 , 
    n6615 , 
    n6616 , 
    n6617 , 
    n6618 , 
    n6619 , 
    n6620 , 
    n6621 , 
    n6622 , 
    n6623 , 
    n6624 , 
    n6625 , 
    n6626 , 
    n6627 , 
    n6628 , 
    n6629 , 
    n6630 , 
    n6631 , 
    n6632 , 
    n6633 , 
    n6634 , 
    n6635 , 
    n6636 , 
    n6637 , 
    n6638 , 
    n6639 , 
    n6640 , 
    n6641 , 
    n6642 , 
    n6643 , 
    n6644 , 
    n6645 , 
    n6646 , 
    n6647 , 
    n6648 , 
    n6649 , 
    n6650 , 
    n6651 , 
    n6652 , 
    n6653 , 
    n6654 , 
    n6655 , 
    n6656 , 
    n6657 , 
    n6658 , 
    n6659 , 
    n6660 , 
    n6661 , 
    n6662 , 
    n6663 , 
    n6664 , 
    n6665 , 
    n6666 , 
    n6667 , 
    n6668 , 
    n6669 , 
    n6670 , 
    n6671 , 
    n6672 , 
    n6673 , 
    n6674 , 
    n6675 , 
    n6676 , 
    n6677 , 
    n6678 , 
    n6679 , 
    n6680 , 
    n6681 , 
    n6682 , 
    n6683 , 
    n6684 , 
    n6685 , 
    n6686 , 
    n6687 , 
    n6688 , 
    n6689 , 
    n6690 , 
    n6691 , 
    n6692 , 
    n6693 , 
    n6694 , 
    n6695 , 
    n6696 , 
    n6697 , 
    n6698 , 
    n6699 , 
    n6700 , 
    n6701 , 
    n6702 , 
    n6703 , 
    n6704 , 
    n6705 , 
    n6706 , 
    n6707 , 
    n6708 , 
    n6709 , 
    n6710 , 
    n6711 , 
    n6712 , 
    n6713 , 
    n6714 , 
    n6715 , 
    n6716 , 
    n6717 , 
    n6718 , 
    n6719 , 
    n6720 , 
    n6721 , 
    n6722 , 
    n6723 , 
    n6724 , 
    n6725 , 
    n6726 , 
    n6727 , 
    n6728 , 
    n6729 , 
    n6730 , 
    n6731 , 
    n6732 , 
    n6733 , 
    n6734 , 
    n6735 , 
    n6736 , 
    n6737 , 
    n6738 , 
    n6739 , 
    n6740 , 
    n6741 , 
    n6742 , 
    n6743 , 
    n6744 , 
    n6745 , 
    n6746 , 
    n6747 , 
    n6748 , 
    n6749 , 
    n6750 , 
    n6751 , 
    n6752 , 
    n6753 , 
    n6754 , 
    n6755 , 
    n6756 , 
    n6757 , 
    n6758 , 
    n6759 , 
    n6760 ;

wire  C0 , 
    RI15b3e9d0_1 , 
    RI15b51198_632 , 
    RI15b51210_633 , 
    RI15b51120_631 , 
    RI15b51288_634 , 
    RI15b54690_745 , 
    RI15b56760_815 , 
    RI15b567d8_816 , 
    RI15b566e8_814 , 
    RI15b570c0_835 , 
    RI15b57138_836 , 
    RI15b571b0_837 , 
    RI15b57228_838 , 
    RI15b572a0_839 , 
    RI15b57318_840 , 
    RI15b57390_841 , 
    RI15b57408_842 , 
    RI15b56850_817 , 
    RI15b568c8_818 , 
    RI15b56940_819 , 
    RI15b569b8_820 , 
    RI15b56a30_821 , 
    RI15b56aa8_822 , 
    RI15b56b20_823 , 
    RI15b56b98_824 , 
    RI15b56c10_825 , 
    RI15b56c88_826 , 
    RI15b56d00_827 , 
    RI15b56d78_828 , 
    RI15b56df0_829 , 
    RI15b56e68_830 , 
    RI15b56ee0_831 , 
    RI15b56f58_832 , 
    RI15b56fd0_833 , 
    RI15b57048_834 , 
    RI15b57480_843 , 
    RI15b574f8_844 , 
    RI15b57570_845 , 
    RI15b4d340_499 , 
    RI15b50e50_625 , 
    RI15b50ec8_626 , 
    RI15b50f40_627 , 
    RI15b50fb8_628 , 
    RI15b51030_629 , 
    RI15b4dac0_515 , 
    RI15b4e9c0_547 , 
    RI15b4ed80_555 , 
    RI15b4fc80_587 , 
    RI15b4e600_539 , 
    RI15b4c800_475 , 
    RI15b4d700_507 , 
    RI15b4c440_467 , 
    RI15b4cbc0_483 , 
    RI15b4cf80_491 , 
    RI15b4f140_563 , 
    RI15b4f8c0_579 , 
    RI15b4e240_531 , 
    RI15b4f500_571 , 
    RI15b4de80_523 , 
    RI15b4d3b8_500 , 
    RI15b4db38_516 , 
    RI15b4ea38_548 , 
    RI15b4edf8_556 , 
    RI15b4fcf8_588 , 
    RI15b4e678_540 , 
    RI15b4c878_476 , 
    RI15b4d778_508 , 
    RI15b4cc38_484 , 
    RI15b4c4b8_468 , 
    RI15b4cff8_492 , 
    RI15b4f1b8_564 , 
    RI15b4f938_580 , 
    RI15b4e2b8_532 , 
    RI15b4f578_572 , 
    RI15b4def8_524 , 
    RI15b4d598_504 , 
    RI15b4dd18_520 , 
    RI15b4ec18_552 , 
    RI15b4efd8_560 , 
    RI15b4fed8_592 , 
    RI15b4e858_544 , 
    RI15b4ca58_480 , 
    RI15b4d958_512 , 
    RI15b4ce18_488 , 
    RI15b4c698_472 , 
    RI15b4d1d8_496 , 
    RI15b4f398_568 , 
    RI15b4fb18_584 , 
    RI15b4e498_536 , 
    RI15b4f758_576 , 
    RI15b4e0d8_528 , 
    RI15b4d4a8_502 , 
    RI15b4dc28_518 , 
    RI15b4eb28_550 , 
    RI15b4eee8_558 , 
    RI15b4fde8_590 , 
    RI15b4c968_478 , 
    RI15b4d868_510 , 
    RI15b4cd28_486 , 
    RI15b4c5a8_470 , 
    RI15b4d0e8_494 , 
    RI15b4e768_542 , 
    RI15b4f2a8_566 , 
    RI15b4fa28_582 , 
    RI15b4e3a8_534 , 
    RI15b4f668_574 , 
    RI15b4dfe8_526 , 
    RI15b4d430_501 , 
    RI15b4dbb0_517 , 
    RI15b4eab0_549 , 
    RI15b4ee70_557 , 
    RI15b4fd70_589 , 
    RI15b4c8f0_477 , 
    RI15b4d7f0_509 , 
    RI15b4d070_493 , 
    RI15b4e6f0_541 , 
    RI15b4c530_469 , 
    RI15b4ccb0_485 , 
    RI15b4f230_565 , 
    RI15b4f9b0_581 , 
    RI15b4e330_533 , 
    RI15b4f5f0_573 , 
    RI15b4df70_525 , 
    RI15b4d520_503 , 
    RI15b4dca0_519 , 
    RI15b4eba0_551 , 
    RI15b4ef60_559 , 
    RI15b4fe60_591 , 
    RI15b4e7e0_543 , 
    RI15b4c9e0_479 , 
    RI15b4d8e0_511 , 
    RI15b4cda0_487 , 
    RI15b4c620_471 , 
    RI15b4d160_495 , 
    RI15b4f320_567 , 
    RI15b4faa0_583 , 
    RI15b4e420_535 , 
    RI15b4f6e0_575 , 
    RI15b4e060_527 , 
    RI15b4c788_474 , 
    RI15b4cf08_490 , 
    RI15b4d688_506 , 
    RI15b4c3c8_466 , 
    RI15b4cb48_482 , 
    RI15b4f0c8_562 , 
    RI15b4e588_538 , 
    RI15b4f848_578 , 
    RI15b4f488_570 , 
    RI15b4de08_522 , 
    RI15b4e1c8_530 , 
    RI15b4d2c8_498 , 
    RI15b4ed08_554 , 
    RI15b4fc08_586 , 
    RI15b4e948_546 , 
    RI15b4da48_514 , 
    RI15b4d250_497 , 
    RI15b4d9d0_513 , 
    RI15b4e8d0_545 , 
    RI15b4ec90_553 , 
    RI15b4fb90_585 , 
    RI15b4e510_537 , 
    RI15b4c710_473 , 
    RI15b4d610_505 , 
    RI15b4cad0_481 , 
    RI15b4c350_465 , 
    RI15b4ce90_489 , 
    RI15b4f050_561 , 
    RI15b4f7d0_577 , 
    RI15b4e150_529 , 
    RI15b4f410_569 , 
    RI15b4dd90_521 , 
    RI15b4c1e8_462 , 
    RI15b4c0f8_460 , 
    RI15b4c170_461 , 
    RI15b4c260_463 , 
    RI15b4c2d8_464 , 
    RI15b667c8_1362 , 
    RI15b66840_1363 , 
    RI15b557e8_782 , 
    RI15b55860_783 , 
    RI15b558d8_784 , 
    RI15b56670_813 , 
    RI15b547f8_748 , 
    RI15b54870_749 , 
    RI15b54780_747 , 
    RI15b55950_785 , 
    RI15b57750_849 , 
    RI15b57660_847 , 
    RI15b576d8_848 , 
    RI15b3ea48_2 , 
    RI15b5c4a8_1014 , 
    RI15b5c520_1015 , 
    RI15b5c598_1016 , 
    RI15b5c430_1013 , 
    RI15b5c610_1017 , 
    RI15b5c688_1018 , 
    RI15b5c700_1019 , 
    RI15b5c778_1020 , 
    RI15b5d2b8_1044 , 
    RI15b5d330_1045 , 
    RI15b5d420_1047 , 
    RI15b5d3a8_1046 , 
    RI15b5b440_979 , 
    RI15b5b080_971 , 
    RI15b5a900_955 , 
    RI15b5acc0_963 , 
    RI15b5b800_987 , 
    RI15b5bbc0_995 , 
    RI15b5bf80_1003 , 
    RI15b5c340_1011 , 
    RI15b59a00_923 , 
    RI15b59dc0_931 , 
    RI15b5a180_939 , 
    RI15b5a540_947 , 
    RI15b59640_915 , 
    RI15b59280_907 , 
    RI15b58b00_891 , 
    RI15b58ec0_899 , 
    RI15b5b008_970 , 
    RI15b5b3c8_978 , 
    RI15b5a4c8_946 , 
    RI15b5a108_938 , 
    RI15b5a888_954 , 
    RI15b5ac48_962 , 
    RI15b59988_922 , 
    RI15b59d48_930 , 
    RI15b5bf08_1002 , 
    RI15b5c2c8_1010 , 
    RI15b595c8_914 , 
    RI15b59208_906 , 
    RI15b58a88_890 , 
    RI15b58e48_898 , 
    RI15b5b788_986 , 
    RI15b5bb48_994 , 
    RI15b5be18_1000 , 
    RI15b5c1d8_1008 , 
    RI15b59118_904 , 
    RI15b594d8_912 , 
    RI15b5a798_952 , 
    RI15b5ab58_960 , 
    RI15b59898_920 , 
    RI15b59c58_928 , 
    RI15b5b2d8_976 , 
    RI15b5af18_968 , 
    RI15b5a3d8_944 , 
    RI15b5a018_936 , 
    RI15b58998_888 , 
    RI15b58d58_896 , 
    RI15b5b698_984 , 
    RI15b5ba58_992 , 
    RI15b59820_919 , 
    RI15b59be0_927 , 
    RI15b5b260_975 , 
    RI15b5aea0_967 , 
    RI15b5a360_943 , 
    RI15b59fa0_935 , 
    RI15b5a720_951 , 
    RI15b5aae0_959 , 
    RI15b58920_887 , 
    RI15b58ce0_895 , 
    RI15b5c160_1007 , 
    RI15b5bda0_999 , 
    RI15b5b620_983 , 
    RI15b5b9e0_991 , 
    RI15b59460_911 , 
    RI15b590a0_903 , 
    RI15b5ae28_966 , 
    RI15b5b1e8_974 , 
    RI15b5c0e8_1006 , 
    RI15b5bd28_998 , 
    RI15b5b5a8_982 , 
    RI15b5b968_990 , 
    RI15b593e8_910 , 
    RI15b59028_902 , 
    RI15b5a6a8_950 , 
    RI15b5a2e8_942 , 
    RI15b59f28_934 , 
    RI15b5aa68_958 , 
    RI15b588a8_886 , 
    RI15b58c68_894 , 
    RI15b597a8_918 , 
    RI15b59b68_926 , 
    RI15b5b170_973 , 
    RI15b5adb0_965 , 
    RI15b59370_909 , 
    RI15b58fb0_901 , 
    RI15b5c070_1005 , 
    RI15b5bcb0_997 , 
    RI15b5a270_941 , 
    RI15b59eb0_933 , 
    RI15b5a630_949 , 
    RI15b58830_885 , 
    RI15b58bf0_893 , 
    RI15b5a9f0_957 , 
    RI15b5b530_981 , 
    RI15b59730_917 , 
    RI15b59af0_925 , 
    RI15b5b8f0_989 , 
    RI15b5bff8_1004 , 
    RI15b5bc38_996 , 
    RI15b592f8_908 , 
    RI15b58f38_900 , 
    RI15b5b0f8_972 , 
    RI15b5ad38_964 , 
    RI15b5a1f8_940 , 
    RI15b59e38_932 , 
    RI15b5a5b8_948 , 
    RI15b596b8_916 , 
    RI15b5b4b8_980 , 
    RI15b5a978_956 , 
    RI15b587b8_884 , 
    RI15b59a78_924 , 
    RI15b5b878_988 , 
    RI15b58b78_892 , 
    RI15b5c3b8_1012 , 
    RI15b5c250_1009 , 
    RI15b5be90_1001 , 
    RI15b5b350_977 , 
    RI15b5af90_969 , 
    RI15b5a810_953 , 
    RI15b5abd0_961 , 
    RI15b5b710_985 , 
    RI15b5bad0_993 , 
    RI15b5a450_945 , 
    RI15b5a090_937 , 
    RI15b59550_913 , 
    RI15b59190_905 , 
    RI15b58a10_889 , 
    RI15b58dd0_897 , 
    RI15b59910_921 , 
    RI15b59cd0_929 , 
    RI15b5d498_1048 , 
    RI15b5d588_1050 , 
    RI15b5d6f0_1053 , 
    RI15b5d600_1051 , 
    RI15b5d678_1052 , 
    RI15b58740_883 , 
    RI15b586c8_882 , 
    RI15b58650_881 , 
    RI15b58560_879 , 
    RI15b585d8_880 , 
    RI15b63e10_1273 , 
    RI15b62f10_1241 , 
    RI15b62c40_1235 , 
    RI15b62cb8_1236 , 
    RI15b62d30_1237 , 
    RI15b62da8_1238 , 
    RI15b62e20_1239 , 
    RI15b62e98_1240 , 
    RI15b62bc8_1234 , 
    RI15b606c0_1155 , 
    RI15b4a370_397 , 
    RI15b4a3e8_398 , 
    RI15b4a460_399 , 
    RI15b4a4d8_400 , 
    RI15b4a550_401 , 
    RI15b4a5c8_402 , 
    RI15b4a640_403 , 
    RI15b4a6b8_404 , 
    RI15b4a730_405 , 
    RI15b4a7a8_406 , 
    RI15b4a820_407 , 
    RI15b4a898_408 , 
    RI15b4a910_409 , 
    RI15b4a988_410 , 
    RI15b4a2f8_396 , 
    RI15b4aa00_411 , 
    RI15b4aa78_412 , 
    RI15b4aaf0_413 , 
    RI15b4ab68_414 , 
    RI15b4abe0_415 , 
    RI15b4ac58_416 , 
    RI15b4acd0_417 , 
    RI15b4ad48_418 , 
    RI15b4adc0_419 , 
    RI15b4ae38_420 , 
    RI15b4aeb0_421 , 
    RI15b4af28_422 , 
    RI15b4afa0_423 , 
    RI15b4b018_424 , 
    RI15b4a280_395 , 
    RI15b44d30_213 , 
    RI15b44cb8_212 , 
    RI15b44da8_214 , 
    RI15b44e20_215 , 
    RI15b47df0_317 , 
    RI15b4b090_425 , 
    RI15b4b108_426 , 
    RI15b4a0a0_391 , 
    RI15b49380_363 , 
    RI15b493f8_364 , 
    RI15b49470_365 , 
    RI15b494e8_366 , 
    RI15b49560_367 , 
    RI15b495d8_368 , 
    RI15b49650_369 , 
    RI15b496c8_370 , 
    RI15b49740_371 , 
    RI15b497b8_372 , 
    RI15b49830_373 , 
    RI15b498a8_374 , 
    RI15b49920_375 , 
    RI15b49998_376 , 
    RI15b49a10_377 , 
    RI15b49a88_378 , 
    RI15b49b00_379 , 
    RI15b49b78_380 , 
    RI15b49bf0_381 , 
    RI15b49c68_382 , 
    RI15b49ce0_383 , 
    RI15b49d58_384 , 
    RI15b49dd0_385 , 
    RI15b49e48_386 , 
    RI15b49ec0_387 , 
    RI15b49f38_388 , 
    RI15b49fb0_389 , 
    RI15b4a028_390 , 
    RI15b4a118_392 , 
    RI15b42918_136 , 
    RI15b449e8_206 , 
    RI15b44a60_207 , 
    RI15b44b50_209 , 
    RI15b44ad8_208 , 
    RI15b44bc8_210 , 
    RI15b41298_88 , 
    RI15b40ed8_80 , 
    RI15b41658_96 , 
    RI15b40758_64 , 
    RI15b41a18_104 , 
    RI15b42198_120 , 
    RI15b42558_128 , 
    RI15b42cd8_144 , 
    RI15b43098_152 , 
    RI15b43458_160 , 
    RI15b43818_168 , 
    RI15b41dd8_112 , 
    RI15b40b18_72 , 
    RI15b40398_56 , 
    RI15b3ffd8_48 , 
    RI15b432f0_157 , 
    RI15b42f30_149 , 
    RI15b43a70_173 , 
    RI15b436b0_165 , 
    RI15b42030_117 , 
    RI15b40d70_77 , 
    RI15b405f0_61 , 
    RI15b40230_53 , 
    RI15b42b70_141 , 
    RI15b414f0_93 , 
    RI15b41130_85 , 
    RI15b418b0_101 , 
    RI15b409b0_69 , 
    RI15b41c70_109 , 
    RI15b423f0_125 , 
    RI15b427b0_133 , 
    RI15b43110_153 , 
    RI15b42d50_145 , 
    RI15b43890_169 , 
    RI15b434d0_161 , 
    RI15b41e50_113 , 
    RI15b40b90_73 , 
    RI15b40410_57 , 
    RI15b40050_49 , 
    RI15b42990_137 , 
    RI15b41310_89 , 
    RI15b40f50_81 , 
    RI15b416d0_97 , 
    RI15b407d0_65 , 
    RI15b41a90_105 , 
    RI15b42210_121 , 
    RI15b425d0_129 , 
    RI15b42828_134 , 
    RI15b411a8_86 , 
    RI15b40de8_78 , 
    RI15b41568_94 , 
    RI15b40668_62 , 
    RI15b41928_102 , 
    RI15b420a8_118 , 
    RI15b42468_126 , 
    RI15b42be8_142 , 
    RI15b42fa8_150 , 
    RI15b43368_158 , 
    RI15b43728_166 , 
    RI15b41ce8_110 , 
    RI15b40a28_70 , 
    RI15b402a8_54 , 
    RI15b3fee8_46 , 
    RI15b42a08_138 , 
    RI15b41388_90 , 
    RI15b40fc8_82 , 
    RI15b41748_98 , 
    RI15b40848_66 , 
    RI15b41b08_106 , 
    RI15b42288_122 , 
    RI15b42648_130 , 
    RI15b42dc8_146 , 
    RI15b43188_154 , 
    RI15b43548_162 , 
    RI15b43908_170 , 
    RI15b41ec8_114 , 
    RI15b40c08_74 , 
    RI15b400c8_50 , 
    RI15b40488_58 , 
    RI15b428a0_135 , 
    RI15b41220_87 , 
    RI15b40e60_79 , 
    RI15b415e0_95 , 
    RI15b406e0_63 , 
    RI15b419a0_103 , 
    RI15b42120_119 , 
    RI15b424e0_127 , 
    RI15b42c60_143 , 
    RI15b43020_151 , 
    RI15b433e0_159 , 
    RI15b437a0_167 , 
    RI15b41d60_111 , 
    RI15b40aa0_71 , 
    RI15b3ff60_47 , 
    RI15b40320_55 , 
    RI15b42e40_147 , 
    RI15b43200_155 , 
    RI15b43980_171 , 
    RI15b435c0_163 , 
    RI15b41f40_115 , 
    RI15b40c80_75 , 
    RI15b40500_59 , 
    RI15b40140_51 , 
    RI15b41b80_107 , 
    RI15b42300_123 , 
    RI15b426c0_131 , 
    RI15b41400_91 , 
    RI15b42a80_139 , 
    RI15b417c0_99 , 
    RI15b408c0_67 , 
    RI15b41040_83 , 
    RI15b42af8_140 , 
    RI15b41478_92 , 
    RI15b410b8_84 , 
    RI15b41838_100 , 
    RI15b40938_68 , 
    RI15b41bf8_108 , 
    RI15b42378_124 , 
    RI15b42738_132 , 
    RI15b42eb8_148 , 
    RI15b43278_156 , 
    RI15b43638_164 , 
    RI15b439f8_172 , 
    RI15b41fb8_116 , 
    RI15b40cf8_76 , 
    RI15b40578_60 , 
    RI15b401b8_52 , 
    RI15b3fd80_43 , 
    RI15b3fc90_41 , 
    RI15b3fd08_42 , 
    RI15b3fe70_45 , 
    RI15b3fdf8_44 , 
    RI15b3fba0_39 , 
    RI15b668b8_1364 , 
    RI15b4a208_394 , 
    RI15b48390_329 , 
    RI15b48408_330 , 
    RI15b48318_328 , 
    RI15b4a190_393 , 
    RI15b4b2e8_430 , 
    RI15b4b1f8_428 , 
    RI15b4b270_429 , 
    RI15b4b360_431 , 
    RI15b4b3d8_432 , 
    RI15b4b450_433 , 
    RI15b4b4c8_434 , 
    RI15b4b540_435 , 
    RI15b4b5b8_436 , 
    RI15b4b630_437 , 
    RI15b4b6a8_438 , 
    RI15b4b720_439 , 
    RI15b4b798_440 , 
    RI15b4b888_442 , 
    RI15b4b810_441 , 
    RI15b4b900_443 , 
    RI15b4b978_444 , 
    RI15b4b9f0_445 , 
    RI15b4ba68_446 , 
    RI15b4bae0_447 , 
    RI15b4bb58_448 , 
    RI15b4bbd0_449 , 
    RI15b4bc48_450 , 
    RI15b4bcc0_451 , 
    RI15b4bd38_452 , 
    RI15b4bdb0_453 , 
    RI15b4be28_454 , 
    RI15b4bea0_455 , 
    RI15b4bf18_456 , 
    RI15b4bf90_457 , 
    RI15b508b0_613 , 
    RI15b4ffc8_594 , 
    RI15b50040_595 , 
    RI15b500b8_596 , 
    RI15b50130_597 , 
    RI15b501a8_598 , 
    RI15b50220_599 , 
    RI15b50298_600 , 
    RI15b50310_601 , 
    RI15b50388_602 , 
    RI15b50400_603 , 
    RI15b50478_604 , 
    RI15b504f0_605 , 
    RI15b50568_606 , 
    RI15b505e0_607 , 
    RI15b50658_608 , 
    RI15b506d0_609 , 
    RI15b50748_610 , 
    RI15b507c0_611 , 
    RI15b50838_612 , 
    RI15b4ff50_593 , 
    RI15b50928_614 , 
    RI15b57fc0_867 , 
    RI15b577c8_850 , 
    RI15b57840_851 , 
    RI15b578b8_852 , 
    RI15b57930_853 , 
    RI15b579a8_854 , 
    RI15b57a20_855 , 
    RI15b57a98_856 , 
    RI15b57b10_857 , 
    RI15b57b88_858 , 
    RI15b57c00_859 , 
    RI15b57c78_860 , 
    RI15b57cf0_861 , 
    RI15b57de0_863 , 
    RI15b559c8_786 , 
    RI15b55a40_787 , 
    RI15b55ab8_788 , 
    RI15b55b30_789 , 
    RI15b55ba8_790 , 
    RI15b55c20_791 , 
    RI15b55c98_792 , 
    RI15b55d10_793 , 
    RI15b55d88_794 , 
    RI15b55e00_795 , 
    RI15b55e78_796 , 
    RI15b55ef0_797 , 
    RI15b55f68_798 , 
    RI15b55fe0_799 , 
    RI15b57d68_862 , 
    RI15b66408_1354 , 
    RI15b65850_1329 , 
    RI15b658c8_1330 , 
    RI15b65940_1331 , 
    RI15b659b8_1332 , 
    RI15b65a30_1333 , 
    RI15b65aa8_1334 , 
    RI15b65b20_1335 , 
    RI15b65b98_1336 , 
    RI15b65c10_1337 , 
    RI15b65c88_1338 , 
    RI15b65d00_1339 , 
    RI15b65d78_1340 , 
    RI15b65df0_1341 , 
    RI15b65e68_1342 , 
    RI15b65ee0_1343 , 
    RI15b65f58_1344 , 
    RI15b65fd0_1345 , 
    RI15b66048_1346 , 
    RI15b660c0_1347 , 
    RI15b66138_1348 , 
    RI15b661b0_1349 , 
    RI15b66228_1350 , 
    RI15b662a0_1351 , 
    RI15b66318_1352 , 
    RI15b66390_1353 , 
    RI15b66480_1355 , 
    RI15b666d8_1360 , 
    RI15b664f8_1356 , 
    RI15b66570_1357 , 
    RI15b3fb28_38 , 
    RI15b66750_1361 , 
    RI15b60be8_1166 , 
    RI15b60c60_1167 , 
    RI15b60cd8_1168 , 
    RI15b63a50_1265 , 
    RI15b61c50_1201 , 
    RI15b62b50_1233 , 
    RI15b56058_800 , 
    RI15b560d0_801 , 
    RI15b56148_802 , 
    RI15b561c0_803 , 
    RI15b56238_804 , 
    RI15b562b0_805 , 
    RI15b56328_806 , 
    RI15b563a0_807 , 
    RI15b56418_808 , 
    RI15b56490_809 , 
    RI15b56508_810 , 
    RI15b56580_811 , 
    RI15b565f8_812 , 
    RI15b58470_877 , 
    RI15b583f8_876 , 
    RI15b57e58_864 , 
    RI15b57ed0_865 , 
    RI15b57f48_866 , 
    RI15b58038_868 , 
    RI15b580b0_869 , 
    RI15b58128_870 , 
    RI15b581a0_871 , 
    RI15b58218_872 , 
    RI15b58290_873 , 
    RI15b58308_874 , 
    RI15b58380_875 , 
    RI15b60648_1154 , 
    RI15b605d0_1153 , 
    RI15b47d78_316 , 
    RI15b47d00_315 , 
    RI15b541e0_735 , 
    RI15b54168_734 , 
    RI15b450f0_221 , 
    RI15b51558_640 , 
    RI15b4c008_458 , 
    RI15b63d98_1272 , 
    RI15b575e8_846 , 
    RI15b63ac8_1266 , 
    RI15b648d8_1296 , 
    RI15b63b40_1267 , 
    RI15b64860_1295 , 
    RI15b63c30_1269 , 
    RI15b63ca8_1270 , 
    RI15b63bb8_1268 , 
    RI15b63e88_1274 , 
    RI15b63f00_1275 , 
    RI15b63d20_1271 , 
    RI15b63f78_1276 , 
    RI15b63ff0_1277 , 
    RI15b64068_1278 , 
    RI15b640e0_1279 , 
    RI15b64158_1280 , 
    RI15b641d0_1281 , 
    RI15b64248_1282 , 
    RI15b642c0_1283 , 
    RI15b64338_1284 , 
    RI15b643b0_1285 , 
    RI15b64428_1286 , 
    RI15b644a0_1287 , 
    RI15b64518_1288 , 
    RI15b64590_1289 , 
    RI15b64608_1290 , 
    RI15b64680_1291 , 
    RI15b646f8_1292 , 
    RI15b64770_1293 , 
    RI15b647e8_1294 , 
    RI15b5d948_1058 , 
    RI15b484f8_332 , 
    RI15b467e8_270 , 
    RI15b5e5f0_1085 , 
    RI15b5ddf8_1068 , 
    RI15b5de70_1069 , 
    RI15b5dee8_1070 , 
    RI15b5df60_1071 , 
    RI15b5dfd8_1072 , 
    RI15b5e050_1073 , 
    RI15b5e0c8_1074 , 
    RI15b5e140_1075 , 
    RI15b5da38_1060 , 
    RI15b5dab0_1061 , 
    RI15b5db28_1062 , 
    RI15b5dba0_1063 , 
    RI15b5e398_1080 , 
    RI15b5e410_1081 , 
    RI15b5e488_1082 , 
    RI15b5e500_1083 , 
    RI15b5dc18_1064 , 
    RI15b5dc90_1065 , 
    RI15b5dd08_1066 , 
    RI15b5dd80_1067 , 
    RI15b5e1b8_1076 , 
    RI15b5e230_1077 , 
    RI15b5e2a8_1078 , 
    RI15b5e320_1079 , 
    RI15b5e578_1084 , 
    RI15b5d9c0_1059 , 
    RI15b5e668_1086 , 
    RI15b5e6e0_1087 , 
    RI15b657d8_1328 , 
    RI15b3eac0_3 , 
    RI15b64ab8_1300 , 
    RI15b3f7e0_31 , 
    RI15b64b30_1301 , 
    RI15b3f768_30 , 
    RI15b64ba8_1302 , 
    RI15b3f6f0_29 , 
    RI15b649c8_1298 , 
    RI15b3f8d0_33 , 
    RI15b64950_1297 , 
    RI15b3f948_34 , 
    RI15b64a40_1299 , 
    RI15b3f858_32 , 
    RI15b64c20_1303 , 
    RI15b3f678_28 , 
    RI15b64c98_1304 , 
    RI15b3f600_27 , 
    RI15b64d10_1305 , 
    RI15b3f588_26 , 
    RI15b64d88_1306 , 
    RI15b3f510_25 , 
    RI15b64e00_1307 , 
    RI15b3f498_24 , 
    RI15b64e78_1308 , 
    RI15b3f420_23 , 
    RI15b64ef0_1309 , 
    RI15b3f3a8_22 , 
    RI15b64f68_1310 , 
    RI15b3f330_21 , 
    RI15b64fe0_1311 , 
    RI15b3f2b8_20 , 
    RI15b65058_1312 , 
    RI15b3f240_19 , 
    RI15b650d0_1313 , 
    RI15b3f1c8_18 , 
    RI15b65148_1314 , 
    RI15b3f150_17 , 
    RI15b65328_1318 , 
    RI15b3ef70_13 , 
    RI15b65238_1316 , 
    RI15b3f060_15 , 
    RI15b652b0_1317 , 
    RI15b3efe8_14 , 
    RI15b651c0_1315 , 
    RI15b3f0d8_16 , 
    RI15b65490_1321 , 
    RI15b3ee08_10 , 
    RI15b65508_1322 , 
    RI15b3ed90_9 , 
    RI15b3eef8_12 , 
    RI15b653a0_1319 , 
    RI15b65418_1320 , 
    RI15b3ee80_11 , 
    RI15b65580_1323 , 
    RI15b655f8_1324 , 
    RI15b3eca0_7 , 
    RI15b3ed18_8 , 
    RI15b3ec28_6 , 
    RI15b65670_1325 , 
    RI15b656e8_1326 , 
    RI15b3ebb0_5 , 
    RI15b65760_1327 , 
    RI15b3eb38_4 , 
    RI15b5c7f0_1021 , 
    RI15b62f88_1242 , 
    RI15b479b8_308 , 
    RI15b665e8_1358 , 
    RI15b47b98_312 , 
    RI15b523e0_671 , 
    RI15b51300_635 , 
    RI15b51378_636 , 
    RI15b513f0_637 , 
    RI15b51468_638 , 
    RI15b52368_670 , 
    RI15b522f0_669 , 
    RI15b52458_672 , 
    RI15b52278_668 , 
    RI15b534c0_707 , 
    RI15b515d0_641 , 
    RI15b51648_642 , 
    RI15b516c0_643 , 
    RI15b51738_644 , 
    RI15b517b0_645 , 
    RI15b51828_646 , 
    RI15b518a0_647 , 
    RI15b51918_648 , 
    RI15b52110_665 , 
    RI15b52188_666 , 
    RI15b514e0_639 , 
    RI15b52200_667 , 
    RI15b51990_649 , 
    RI15b51a08_650 , 
    RI15b51a80_651 , 
    RI15b51af8_652 , 
    RI15b51b70_653 , 
    RI15b51be8_654 , 
    RI15b51c60_655 , 
    RI15b51cd8_656 , 
    RI15b51d50_657 , 
    RI15b51dc8_658 , 
    RI15b51e40_659 , 
    RI15b51eb8_660 , 
    RI15b51f30_661 , 
    RI15b51fa8_662 , 
    RI15b52020_663 , 
    RI15b52098_664 , 
    RI15b548e8_750 , 
    RI15b54b40_755 , 
    RI15b54bb8_756 , 
    RI15b54960_751 , 
    RI15b549d8_752 , 
    RI15b54a50_753 , 
    RI15b54ac8_754 , 
    RI15b55770_781 , 
    RI15b54c30_757 , 
    RI15b54ca8_758 , 
    RI15b52f98_696 , 
    RI15b509a0_615 , 
    RI15b50a18_616 , 
    RI15b50a90_617 , 
    RI15b50b08_618 , 
    RI15b46e00_283 , 
    RI15b48480_331 , 
    RI15b486d8_336 , 
    RI15b48570_333 , 
    RI15b48750_337 , 
    RI15b488b8_340 , 
    RI15b48a20_343 , 
    RI15b48930_341 , 
    RI15b48a98_344 , 
    RI15b48660_335 , 
    RI15b485e8_334 , 
    RI15b48840_339 , 
    RI15b487c8_338 , 
    RI15b489a8_342 , 
    RI15b48b10_345 , 
    RI15b49308_362 , 
    RI15b48228_326 , 
    RI15b482a0_327 , 
    RI15b4b180_427 , 
    RI15b45348_226 , 
    RI15b4c080_459 , 
    RI15b54d20_759 , 
    RI15b54d98_760 , 
    RI15b54e10_761 , 
    RI15b54e88_762 , 
    RI15b54f00_763 , 
    RI15b54f78_764 , 
    RI15b54ff0_765 , 
    RI15b55068_766 , 
    RI15b550e0_767 , 
    RI15b55158_768 , 
    RI15b551d0_769 , 
    RI15b55248_770 , 
    RI15b552c0_771 , 
    RI15b55338_772 , 
    RI15b553b0_773 , 
    RI15b554a0_775 , 
    RI15b55428_774 , 
    RI15b55518_776 , 
    RI15b55590_777 , 
    RI15b55608_778 , 
    RI15b55680_779 , 
    RI15b52908_682 , 
    RI15b53f10_729 , 
    RI15b556f8_780 , 
    RI15b52b60_687 , 
    RI15b61cc8_1202 , 
    RI15b62ad8_1232 , 
    RI15b61d40_1203 , 
    RI15b63528_1254 , 
    RI15b635a0_1255 , 
    RI15b63618_1256 , 
    RI15b63690_1257 , 
    RI15b63708_1258 , 
    RI15b63780_1259 , 
    RI15b637f8_1260 , 
    RI15b63870_1261 , 
    RI15b638e8_1262 , 
    RI15b63960_1263 , 
    RI15b63168_1246 , 
    RI15b631e0_1247 , 
    RI15b63258_1248 , 
    RI15b632d0_1249 , 
    RI15b63348_1250 , 
    RI15b633c0_1251 , 
    RI15b63438_1252 , 
    RI15b63000_1243 , 
    RI15b63078_1244 , 
    RI15b630f0_1245 , 
    RI15b634b0_1253 , 
    RI15b639d8_1264 , 
    RI15b60d50_1169 , 
    RI15b60fa8_1174 , 
    RI15b61020_1175 , 
    RI15b60dc8_1170 , 
    RI15b60e40_1171 , 
    RI15b60eb8_1172 , 
    RI15b60f30_1173 , 
    RI15b61bd8_1200 , 
    RI15b61098_1176 , 
    RI15b61110_1177 , 
    RI15b61188_1178 , 
    RI15b61200_1179 , 
    RI15b61278_1180 , 
    RI15b612f0_1181 , 
    RI15b61368_1182 , 
    RI15b5fdd8_1136 , 
    RI15b5f658_1120 , 
    RI15b66660_1359 , 
    RI15b62100_1211 , 
    RI15b61db8_1204 , 
    RI15b61e30_1205 , 
    RI15b61ea8_1206 , 
    RI15b61f20_1207 , 
    RI15b61f98_1208 , 
    RI15b62010_1209 , 
    RI15b62088_1210 , 
    RI15b45438_228 , 
    RI15b477d8_304 , 
    RI15b5c868_1022 , 
    RI15b5c8e0_1023 , 
    RI15b5c958_1024 , 
    RI15b5c9d0_1025 , 
    RI15b5ca48_1026 , 
    RI15b5cac0_1027 , 
    RI15b5cb38_1028 , 
    RI15b5cbb0_1029 , 
    RI15b5cc28_1030 , 
    RI15b5cca0_1031 , 
    RI15b5cd18_1032 , 
    RI15b5cd90_1033 , 
    RI15b5ce08_1034 , 
    RI15b5ce80_1035 , 
    RI15b5cef8_1036 , 
    RI15b5cf70_1037 , 
    RI15b5f388_1114 , 
    RI15b3f9c0_35 , 
    RI15b60738_1156 , 
    RI15b3fa38_36 , 
    RI15b5e848_1090 , 
    RI15b60828_1158 , 
    RI15b470d0_289 , 
    RI15b46950_273 , 
    RI15b43bd8_176 , 
    RI15b43c50_177 , 
    RI15b43cc8_178 , 
    RI15b43b60_175 , 
    RI15b43d40_179 , 
    RI15b43db8_180 , 
    RI15b43e30_181 , 
    RI15b43ea8_182 , 
    RI15b43f20_183 , 
    RI15b43f98_184 , 
    RI15b44010_185 , 
    RI15b44268_190 , 
    RI15b44088_186 , 
    RI15b44100_187 , 
    RI15b44178_188 , 
    RI15b441f0_189 , 
    RI15b43ae8_174 , 
    RI15b442e0_191 , 
    RI15b44358_192 , 
    RI15b443d0_193 , 
    RI15b445b0_197 , 
    RI15b44448_194 , 
    RI15b444c0_195 , 
    RI15b44538_196 , 
    RI15b44628_198 , 
    RI15b446a0_199 , 
    RI15b44718_200 , 
    RI15b44790_201 , 
    RI15b44808_202 , 
    RI15b44880_203 , 
    RI15b62178_1212 , 
    RI15b621f0_1213 , 
    RI15b62268_1214 , 
    RI15b622e0_1215 , 
    RI15b62358_1216 , 
    RI15b623d0_1217 , 
    RI15b62448_1218 , 
    RI15b624c0_1219 , 
    RI15b62538_1220 , 
    RI15b625b0_1221 , 
    RI15b62628_1222 , 
    RI15b626a0_1223 , 
    RI15b62718_1224 , 
    RI15b62790_1225 , 
    RI15b62808_1226 , 
    RI15b62880_1227 , 
    RI15b628f8_1228 , 
    RI15b62970_1229 , 
    RI15b629e8_1230 , 
    RI15b62a60_1231 , 
    RI15b613e0_1183 , 
    RI15b5cfe8_1038 , 
    RI15b5d060_1039 , 
    RI15b5d0d8_1040 , 
    RI15b5d150_1041 , 
    RI15b5d1c8_1042 , 
    RI15b45618_232 , 
    RI15b53538_708 , 
    RI15b5d768_1054 , 
    RI15b5d7e0_1055 , 
    RI15b5d858_1056 , 
    RI15b5d8d0_1057 , 
    RI15b5e758_1088 , 
    RI15b5e7d0_1089 , 
    RI15b5e8c0_1091 , 
    RI15b5f9a0_1127 , 
    RI15b615c0_1187 , 
    RI15b61458_1184 , 
    RI15b614d0_1185 , 
    RI15b61548_1186 , 
    RI15b61638_1188 , 
    RI15b616b0_1189 , 
    RI15b61728_1190 , 
    RI15b617a0_1191 , 
    RI15b5ec08_1098 , 
    RI15b526b0_677 , 
    RI15b46ba8_278 , 
    RI15b53f88_730 , 
    RI15b603f0_1149 , 
    RI15b45d98_248 , 
    RI15b475f8_300 , 
    RI15b3fab0_37 , 
    RI15b45168_222 , 
    RI15b542d0_737 , 
    RI15b45ac8_242 , 
    RI15b527a0_679 , 
    RI15b53808_714 , 
    RI15b53088_698 , 
    RI15b61818_1192 , 
    RI15b61890_1193 , 
    RI15b61908_1194 , 
    RI15b61980_1195 , 
    RI15b619f8_1196 , 
    RI15b60468_1150 , 
    RI15b5ee60_1103 , 
    RI15b54618_744 , 
    RI15b54708_746 , 
    RI15b46fe0_287 , 
    RI15b60918_1160 , 
    RI15b48b88_346 , 
    RI15b48c00_347 , 
    RI15b48c78_348 , 
    RI15b48cf0_349 , 
    RI15b48d68_350 , 
    RI15b48de0_351 , 
    RI15b48e58_352 , 
    RI15b48ed0_353 , 
    RI15b48f48_354 , 
    RI15b48fc0_355 , 
    RI15b490b0_357 , 
    RI15b49128_358 , 
    RI15b49038_356 , 
    RI15b49290_361 , 
    RI15b491a0_359 , 
    RI15b49218_360 , 
    RI15b460e0_255 , 
    RI15b476e8_302 , 
    RI15b53c40_723 , 
    RI15b52638_676 , 
    RI15b45f78_252 , 
    RI15b45e88_250 , 
    RI15b45f00_251 , 
    RI15b45ff0_253 , 
    RI15b44e98_216 , 
    RI15b44f10_217 , 
    RI15b44f88_218 , 
    RI15b45000_219 , 
    RI15b54258_736 , 
    RI15b53b50_721 , 
    RI15b53da8_726 , 
    RI15b5f220_1111 , 
    RI15b47328_294 , 
    RI15b45a50_241 , 
    RI15b584e8_878 , 
    RI15b535b0_709 , 
    RI15b52e30_693 , 
    RI15b53e20_727 , 
    RI15b60288_1146 , 
    RI15b3fc18_40 , 
    RI15b608a0_1159 , 
    RI15b45780_235 , 
    RI15b52cc8_690 , 
    RI15b525c0_675 , 
    RI15b47418_296 , 
    RI15b50b80_619 , 
    RI15b50bf8_620 , 
    RI15b50c70_621 , 
    RI15b50ce8_622 , 
    RI15b44c40_211 , 
    RI15b46a40_275 , 
    RI15b60af8_1164 , 
    RI15b47f58_320 , 
    RI15b53718_712 , 
    RI15b5fb80_1131 , 
    RI15b45d20_247 , 
    RI15b52f20_695 , 
    RI15b47ee0_319 , 
    RI15b543c0_739 , 
    RI15b61a70_1197 , 
    RI15b61ae8_1198 , 
    RI15b5ef50_1105 , 
    RI15b5ec80_1099 , 
    RI15b50d60_623 , 
    RI15b50dd8_624 , 
    RI15b53448_706 , 
    RI15b54000_731 , 
    RI15b529f8_684 , 
    RI15b5f838_1124 , 
    RI15b5f0b8_1108 , 
    RI15b53880_715 , 
    RI15b5fce8_1134 , 
    RI15b46d10_281 , 
    RI15b52890_681 , 
    RI15b5fd60_1135 , 
    RI15b5f5e0_1119 , 
    RI15b454b0_229 , 
    RI15b46860_271 , 
    RI15b540f0_733 , 
    RI15b60558_1152 , 
    RI15b47490_297 , 
    RI15b471c0_291 , 
    RI15b47238_292 , 
    RI15b539e8_718 , 
    RI15b53268_702 , 
    RI15b5f130_1109 , 
    RI15b5fb08_1130 , 
    RI15b607b0_1157 , 
    RI15b544b0_741 , 
    RI15b604e0_1151 , 
    RI15b5eed8_1104 , 
    RI15b510a8_630 , 
    RI15b5d240_1043 , 
    RI15b463b0_261 , 
    RI15b46428_262 , 
    RI15b5f298_1112 , 
    RI15b47a30_309 , 
    RI15b53bc8_722 , 
    RI15b46338_260 , 
    RI15b47c10_313 , 
    RI15b48048_322 , 
    RI15b464a0_263 , 
    RI15b5ecf8_1100 , 
    RI15b53628_710 , 
    RI15b52ea8_694 , 
    RI15b47850_305 , 
    RI15b47670_301 , 
    RI15b46068_254 , 
    RI15b524d0_673 , 
    RI15b52ae8_686 , 
    RI15b451e0_223 , 
    RI15b52548_674 , 
    RI15b60030_1141 , 
    RI15b457f8_236 , 
    RI15b60990_1161 , 
    RI15b53ad8_720 , 
    RI15b5ff40_1139 , 
    RI15b45528_230 , 
    RI15b5fa18_1128 , 
    RI15b53358_704 , 
    RI15b5f7c0_1123 , 
    RI15b462c0_259 , 
    RI15b453c0_227 , 
    RI15b45870_237 , 
    RI15b46518_264 , 
    RI15b47058_288 , 
    RI15b60b70_1165 , 
    RI15b45bb8_244 , 
    RI15b533d0_705 , 
    RI15b47e68_318 , 
    RI15b44970_205 , 
    RI15b53100_699 , 
    RI15b47fd0_321 , 
    RI15b5f568_1118 , 
    RI15b480c0_323 , 
    RI15b45960_239 , 
    RI15b52980_683 , 
    RI15b53cb8_724 , 
    RI15b60120_1143 , 
    RI15b5f4f0_1117 , 
    RI15b46248_258 , 
    RI15b46590_265 , 
    RI15b5fe50_1137 , 
    RI15b52c50_689 , 
    RI15b47aa8_310 , 
    RI15b47b20_311 , 
    RI15b61b60_1199 , 
    RI15b5efc8_1106 , 
    RI15b468d8_272 , 
    RI15b60378_1148 , 
    RI15b5ed70_1101 , 
    RI15b5f6d0_1121 , 
    RI15b46c20_279 , 
    RI15b5d510_1049 , 
    RI15b46ab8_276 , 
    RI15b45258_224 , 
    RI15b46f68_286 , 
    RI15b461d0_257 , 
    RI15b472b0_293 , 
    RI15b5f928_1126 , 
    RI15b5f1a8_1110 , 
    RI15b536a0_711 , 
    RI15b45b40_243 , 
    RI15b48138_324 , 
    RI15b5f400_1115 , 
    RI15b46b30_277 , 
    RI15b46608_266 , 
    RI15b45690_233 , 
    RI15b53790_713 , 
    RI15b5fbf8_1132 , 
    RI15b54078_732 , 
    RI15b46e78_284 , 
    RI15b46c98_280 , 
    RI15b53e98_728 , 
    RI15b455a0_231 , 
    RI15b47940_307 , 
    RI15b45e10_249 , 
    RI15b5fa90_1129 , 
    RI15b5f310_1113 , 
    RI15b54348_738 , 
    RI15b60a08_1162 , 
    RI15b60210_1145 , 
    RI15b478c8_306 , 
    RI15b47c88_314 , 
    RI15b46680_267 , 
    RI15b46158_256 , 
    RI15b5fc70_1133 , 
    RI15b53a60_719 , 
    RI15b532e0_703 , 
    RI15b538f8_716 , 
    RI15b5eb18_1096 , 
    RI15b52728_678 , 
    RI15b600a8_1142 , 
    RI15b5eaa0_1095 , 
    RI15b5ede8_1102 , 
    RI15b5f040_1107 , 
    RI15b5eb90_1097 , 
    RI15b60198_1144 , 
    RI15b481b0_325 , 
    RI15b545a0_743 , 
    RI15b452d0_225 , 
    RI15b46d88_282 , 
    RI15b5ea28_1094 , 
    RI15b54438_740 , 
    RI15b47508_298 , 
    RI15b466f8_268 , 
    RI15b53178_700 , 
    RI15b47148_290 , 
    RI15b469c8_274 , 
    RI15b458e8_238 , 
    RI15b448f8_204 , 
    RI15b52a70_685 , 
    RI15b52818_680 , 
    RI15b5ffb8_1140 , 
    RI15b5e9b0_1093 , 
    RI15b5f8b0_1125 , 
    RI15b531f0_701 , 
    RI15b46ef0_285 , 
    RI15b45ca8_246 , 
    RI15b52bd8_688 , 
    RI15b53970_717 , 
    RI15b52db8_692 , 
    RI15b47580_299 , 
    RI15b5e938_1092 , 
    RI15b45078_220 , 
    RI15b60300_1147 , 
    RI15b60a80_1163 , 
    RI15b5f478_1116 , 
    RI15b473a0_295 , 
    RI15b47760_303 , 
    RI15b5fec8_1138 , 
    RI15b5f748_1122 , 
    RI15b45c30_245 , 
    RI15b46770_269 , 
    RI15b53010_697 , 
    RI15b53d30_725 , 
    RI15b52d40_691 , 
    RI15b45708_234 , 
    RI15b54528_742 , 
    RI15b459d8_240 , 
    R_187c_13cca558 , 
    R_125d_156aaaf8 , 
    R_c3e_13d2c178 , 
    R_61f_117eb278 , 
    R_187d_117f5b38 , 
    R_125e_13b8fe18 , 
    R_c3f_123b4358 , 
    R_187b_13ccb278 , 
    R_620_13dfb518 , 
    R_125c_15816b78 , 
    R_c3d_13c22918 , 
    R_61e_14a0c538 , 
    R_5e7_10080958 , 
    R_c06_170189e8 , 
    R_18b4_1162f978 , 
    R_1225_13c08298 , 
    R_1844_117ef378 , 
    R_1295_123bcf58 , 
    R_c76_15ff42e8 , 
    R_657_13bf5c78 , 
    R_187e_140ac0d8 , 
    R_125f_13c0f638 , 
    R_c40_1580a9b8 , 
    R_621_11c70318 , 
    R_187a_13ddd2d8 , 
    R_61d_123b84f8 , 
    R_125b_1162bf58 , 
    R_c3c_15ff9928 , 
    R_12be_13ccf378 , 
    R_5be_11c6a738 , 
    R_bdd_17016508 , 
    R_c9f_11636598 , 
    R_11fc_13ddf7b8 , 
    R_680_10085638 , 
    R_181b_13d430d8 , 
    R_18dd_13c062b8 , 
    R_180c_156b4eb8 , 
    R_12cd_13d535d8 , 
    R_5af_1700c3c8 , 
    R_cae_14a14ff8 , 
    R_bce_15ff4608 , 
    R_68f_13befcd8 , 
    R_18ec_13d204b8 , 
    R_11ed_116361d8 , 
    R_187f_15811038 , 
    R_1260_13d3b6f8 , 
    R_c41_14a0bef8 , 
    R_622_123b3bd8 , 
    R_61c_13d56378 , 
    R_c3b_150e7c58 , 
    R_1879_15ff5c88 , 
    R_125a_13bf58b8 , 
    R_f82_13c1cd38 , 
    R_963_13c209d8 , 
    R_8fa_117ec678 , 
    R_f19_15ff0648 , 
    R_1538_13d29bf8 , 
    R_15a1_150e22f8 , 
    R_158f_13cd9058 , 
    R_f70_17015608 , 
    R_951_156b2578 , 
    R_90c_13c0e0f8 , 
    R_f2b_140b8838 , 
    R_154a_1587f278 , 
    R_1880_13c22738 , 
    R_1261_13ccc0d8 , 
    R_c42_117eb818 , 
    R_623_140b3158 , 
    R_61b_11c70458 , 
    R_c3a_13b96218 , 
    R_1259_13d23578 , 
    R_1878_1162da38 , 
    R_ce6_14875d78 , 
    R_1924_13d1df38 , 
    R_11b5_13d56f58 , 
    R_577_1162c818 , 
    R_6c7_10082438 , 
    R_17d4_13cda278 , 
    R_1305_10081fd8 , 
    R_b96_15812b18 , 
    R_1881_156b0638 , 
    R_1262_12fc1698 , 
    R_c43_140b0138 , 
    R_624_13d421d8 , 
    R_61a_14b2a318 , 
    R_c39_117eaeb8 , 
    R_1258_117e8618 , 
    R_1877_1162cdb8 , 
    R_119b_15ffa3c8 , 
    R_55d_13b8e5b8 , 
    R_131f_158106d8 , 
    R_6e1_13c0fb38 , 
    R_17ba_15fed6c8 , 
    R_b7c_13b96e98 , 
    R_193e_123b6018 , 
    R_d00_117ec358 , 
    R_1323_13d5b878 , 
    R_6e5_15ff5328 , 
    R_559_13c024d8 , 
    R_1197_13bf4918 , 
    R_1942_11c6dd98 , 
    R_d04_14a16df8 , 
    R_17b6_13dec158 , 
    R_b78_13c10c18 , 
    R_13ca_13d2c718 , 
    R_19e9_13bf62b8 , 
    R_170f_150defb8 , 
    R_10f0_140b1ad8 , 
    R_ad1_11c6ac38 , 
    R_78c_13d5d3f8 , 
    R_dab_140b3dd8 , 
    R_883_13b936f8 , 
    R_ff9_11631958 , 
    R_ea2_150dd758 , 
    R_9da_13cd8018 , 
    R_1618_117f3658 , 
    R_14c1_123ba4d8 , 
    R_b5e_14a0f918 , 
    R_179c_123bb018 , 
    R_133d_13cd4e18 , 
    R_6ff_14a0a918 , 
    R_195c_150ddf78 , 
    R_117d_123b8c78 , 
    R_d1e_124c2cd8 , 
    R_5f7_12fbf758 , 
    R_c16_13df9858 , 
    R_1235_15880cb8 , 
    R_1854_1580fd78 , 
    R_18a4_13bf2d98 , 
    R_1285_100890f8 , 
    R_c66_13bed2f8 , 
    R_647_13d51af8 , 
    R_1882_13d1fbf8 , 
    R_1263_123be498 , 
    R_c44_13c229b8 , 
    R_625_13c1e638 , 
    R_619_156b6718 , 
    R_c38_117efd78 , 
    R_1257_14a0f0f8 , 
    R_1876_15ffcb28 , 
    R_985_1587c4d8 , 
    R_1516_12fc1eb8 , 
    R_15c3_13c02078 , 
    R_8d8_13d22fd8 , 
    R_fa4_13d1e898 , 
    R_ef7_1162bd78 , 
    R_1663_124c2698 , 
    R_838_1580b8b8 , 
    R_a25_13bf4ff8 , 
    R_1476_1486bd78 , 
    R_1044_13d57818 , 
    R_e57_13b8f738 , 
    R_15fa_13c0bb78 , 
    R_ec0_13c1bf78 , 
    R_fdb_15ff7308 , 
    R_14df_14a0cdf8 , 
    R_9bc_15812758 , 
    R_8a1_13d21818 , 
    R_1883_13d41058 , 
    R_1264_13c02758 , 
    R_c45_13d24c98 , 
    R_626_123b86d8 , 
    R_618_1587ea58 , 
    R_c37_13c0bfd8 , 
    R_1256_13d54258 , 
    R_1875_158179d8 , 
    R_1145_13b98658 , 
    R_737_116313b8 , 
    R_b26_1486a518 , 
    R_d56_117e9d38 , 
    R_1764_13ccf7d8 , 
    R_1375_13c275f8 , 
    R_1994_123bac58 , 
    R_143d_13bf2258 , 
    R_a5e_1587ed78 , 
    R_e1e_13c1bbb8 , 
    R_107d_15888418 , 
    R_7ff_13cd45f8 , 
    R_169c_15885fd8 , 
    R_1a5c_13de04d8 , 
    R_1a48_13c1ff38 , 
    R_a72_1486d358 , 
    R_1429_13d23438 , 
    R_1091_14a11d58 , 
    R_e0a_13bfa3b8 , 
    R_16b0_140aae18 , 
    R_7eb_123b8278 , 
    R_12c6_13cd49b8 , 
    R_5b6_117f1f38 , 
    R_ca7_140b4418 , 
    R_bd5_13d51698 , 
    R_688_13b99af8 , 
    R_11f4_13d1e6b8 , 
    R_18e5_13d45658 , 
    R_1813_13d29c98 , 
    R_16d9_14a17cf8 , 
    R_1a1f_11c70958 , 
    R_1400_14b29b98 , 
    R_de1_13cd0638 , 
    R_7c2_15ffa508 , 
    R_a9b_100865d8 , 
    R_10ba_15881938 , 
    R_1805_14b271b8 , 
    R_5a8_123b8318 , 
    R_cb5_170107e8 , 
    R_bc7_13c2a758 , 
    R_696_10082ed8 , 
    R_18f3_15ffc628 , 
    R_11e6_14b222f8 , 
    R_12d4_11634d38 , 
    R_119f_156b4738 , 
    R_561_1162a658 , 
    R_6dd_117f36f8 , 
    R_131b_15ff76c8 , 
    R_17be_15816538 , 
    R_b80_13cd8338 , 
    R_cfc_1700d2c8 , 
    R_193a_15885718 , 
    R_5da_13df70f8 , 
    R_18c1_11c6f738 , 
    R_bf9_13d28ed8 , 
    R_12a2_13bf2578 , 
    R_1218_13d28078 , 
    R_c83_13d59f78 , 
    R_1837_13deb9d8 , 
    R_664_123b47b8 , 
    R_e39_156b3518 , 
    R_a43_14b1feb8 , 
    R_81a_13cceb58 , 
    R_1062_117eedd8 , 
    R_1458_13df07f8 , 
    R_1681_140b99b8 , 
    R_1327_124c2b98 , 
    R_6e9_156b3158 , 
    R_555_13d59b18 , 
    R_1193_13b97438 , 
    R_1946_14a16858 , 
    R_d08_13d59938 , 
    R_b74_123c0478 , 
    R_17b2_13cd6498 , 
    R_113a_117eb458 , 
    R_742_14a129d8 , 
    R_b1b_11629758 , 
    R_d61_11633618 , 
    R_1380_15887338 , 
    R_1759_14874518 , 
    R_199f_13d3c9b8 , 
    R_1884_13cd1c18 , 
    R_1265_156b0818 , 
    R_c46_1580b598 , 
    R_627_117efb98 , 
    R_617_158807b8 , 
    R_c36_156b63f8 , 
    R_1255_1580dbb8 , 
    R_1874_13df9c18 , 
    R_87a_13c286d8 , 
    R_1002_14a17938 , 
    R_e99_123ba258 , 
    R_9e3_170110a8 , 
    R_1621_117eacd8 , 
    R_14b8_123b31d8 , 
    R_edf_117f5bd8 , 
    R_14fe_13d55518 , 
    R_15db_117f7258 , 
    R_fbc_13beb9f8 , 
    R_8c0_11631ef8 , 
    R_99d_13cd4d78 , 
    R_845_15888918 , 
    R_1656_117f4af8 , 
    R_1483_13d53d58 , 
    R_a18_12fbdef8 , 
    R_e64_14875058 , 
    R_1037_15815098 , 
    R_d8e_11630878 , 
    R_172c_13d39d58 , 
    R_13ad_14a12618 , 
    R_19cc_13cda1d8 , 
    R_110d_13dd5cb8 , 
    R_aee_117e9478 , 
    R_76f_117f4378 , 
    R_ccd_13b8c8f8 , 
    R_590_13dd64d8 , 
    R_17ed_156b36f8 , 
    R_190b_14872038 , 
    R_6ae_156ab958 , 
    R_baf_1700cd28 , 
    R_12ec_124c3778 , 
    R_11ce_11c6cad8 , 
    R_17a3_150e7398 , 
    R_1336_148754b8 , 
    R_6f8_13c1c018 , 
    R_1184_150e6498 , 
    R_1955_14b235b8 , 
    R_d17_14b27398 , 
    R_b65_13dde318 , 
    R_1885_1486cdb8 , 
    R_1266_14a12438 , 
    R_c47_100803b8 , 
    R_628_117eb098 , 
    R_616_170152e8 , 
    R_c35_123b88b8 , 
    R_1254_150e59f8 , 
    R_1873_12fc2278 , 
    R_74a_1008cb18 , 
    R_1132_15880e98 , 
    R_d69_14b23158 , 
    R_b13_140b3d38 , 
    R_1388_140aaf58 , 
    R_19a7_140b9b98 , 
    R_1751_1007feb8 , 
    R_b57_13ccd6b8 , 
    R_1344_117f3018 , 
    R_1795_1008b678 , 
    R_706_1580bd18 , 
    R_1963_13d1f478 , 
    R_1176_17015b08 , 
    R_d25_15882298 , 
    R_1590_150e4b98 , 
    R_f71_124c4998 , 
    R_952_14b26e98 , 
    R_90b_13d41af8 , 
    R_f2a_1162a158 , 
    R_1549_1587ff98 , 
    R_5c6_15816218 , 
    R_12b6_1587db58 , 
    R_be5_140b5818 , 
    R_c97_156b09f8 , 
    R_1204_13c23b38 , 
    R_678_15884ef8 , 
    R_1823_13d53df8 , 
    R_18d5_11636098 , 
    R_ed8_117e9c98 , 
    R_15e2_14a140f8 , 
    R_14f7_13b965d8 , 
    R_fc3_14b27e38 , 
    R_8b9_14875e18 , 
    R_9a4_117ee018 , 
    R_1a04_13c22b98 , 
    R_13e5_13de07f8 , 
    R_16f4_123b9fd8 , 
    R_dc6_14873f78 , 
    R_10d5_13b94a58 , 
    R_7a7_116355f8 , 
    R_ab6_15814e18 , 
    R_1886_11638c58 , 
    R_1267_14b23f18 , 
    R_c48_13bf5e58 , 
    R_629_150e7e38 , 
    R_615_13c1d7d8 , 
    R_c34_15ff1228 , 
    R_1253_13d222b8 , 
    R_1872_13ccb4f8 , 
    R_16f6_116389d8 , 
    R_10d7_156b5778 , 
    R_ab8_156ac8f8 , 
    R_1a02_13cd8298 , 
    R_13e3_14a0a7d8 , 
    R_7a5_13d456f8 , 
    R_dc4_11634b58 , 
    R_b4d_1700f208 , 
    R_710_156ac718 , 
    R_178b_1580ca38 , 
    R_196d_117eb8b8 , 
    R_d2f_13dedf58 , 
    R_116c_140b8338 , 
    R_134e_13d282f8 , 
    R_1a06_1486e1b8 , 
    R_13e7_116377b8 , 
    R_dc8_1162b058 , 
    R_7a9_123bd458 , 
    R_16f2_158857b8 , 
    R_ab4_12fbed58 , 
    R_10d3_158899f8 , 
    R_85a_156b1a38 , 
    R_1498_15811c18 , 
    R_1641_150db8b8 , 
    R_a03_123bd818 , 
    R_e79_13cd8658 , 
    R_1022_11c6cf38 , 
    R_150d_14b21678 , 
    R_15cc_14a0ba98 , 
    R_8cf_13ded9b8 , 
    R_fad_140ac038 , 
    R_eee_11632e98 , 
    R_98e_12fbecb8 , 
    R_13bd_13df6c98 , 
    R_19dc_156b6858 , 
    R_171c_117ecb78 , 
    R_10fd_117eef18 , 
    R_ade_13dd7658 , 
    R_77f_117f4558 , 
    R_d9e_13ddc3d8 , 
    R_16f8_14a0e018 , 
    R_10d9_123b9538 , 
    R_aba_13c29678 , 
    R_7a3_13ccb138 , 
    R_dc2_158108b8 , 
    R_13e1_156b8478 , 
    R_1a00_123b7f58 , 
    R_971_13df5618 , 
    R_8ec_123bbd38 , 
    R_15af_14866eb8 , 
    R_f0b_13cd72f8 , 
    R_f90_15812438 , 
    R_152a_13df8818 , 
    R_c15_15fee528 , 
    R_1234_15ff9e28 , 
    R_1853_13dd8738 , 
    R_18a5_170177c8 , 
    R_1286_124c4858 , 
    R_c67_13ccba98 , 
    R_648_15814058 , 
    R_5f6_13cce018 , 
    R_c05_14866d78 , 
    R_18b5_10087cf8 , 
    R_1224_13ccff58 , 
    R_1296_13dda7b8 , 
    R_1843_1580a878 , 
    R_c77_13d523b8 , 
    R_658_140ae1f8 , 
    R_5e6_13d46698 , 
    R_1a08_14b1b958 , 
    R_13e9_13d22358 , 
    R_dca_14b297d8 , 
    R_7ab_15887ab8 , 
    R_ab2_13df75f8 , 
    R_10d1_13d55d38 , 
    R_16f0_14b1e978 , 
    R_d87_123bae38 , 
    R_1733_15ff79e8 , 
    R_13a6_156b1718 , 
    R_1114_13d46ff8 , 
    R_19c5_13bf6ad8 , 
    R_af5_13c1b6b8 , 
    R_768_158896d8 , 
    R_964_123c1f58 , 
    R_8f9_117ee658 , 
    R_f18_14a19d78 , 
    R_1537_117e9b58 , 
    R_15a2_13ccce98 , 
    R_f83_14a0e978 , 
    R_1887_17018da8 , 
    R_1268_13d38278 , 
    R_c49_123b36d8 , 
    R_62a_13d42278 , 
    R_614_13c2a258 , 
    R_c33_150e7bb8 , 
    R_1252_116378f8 , 
    R_1871_13defad8 , 
    R_11a3_13c1be38 , 
    R_565_13ddbb18 , 
    R_6d9_11636818 , 
    R_1317_1580c5d8 , 
    R_17c2_13c03518 , 
    R_b84_156b5278 , 
    R_cf8_15881a78 , 
    R_1936_13d2a558 , 
    R_13b4_156abb38 , 
    R_19d3_13bf92d8 , 
    R_1725_13cd9a58 , 
    R_1106_14b1c718 , 
    R_ae7_13cd22f8 , 
    R_776_14873bb8 , 
    R_d95_15815778 , 
    R_feb_1486c818 , 
    R_eb0_13d53498 , 
    R_14cf_14b1bd18 , 
    R_9cc_158172f8 , 
    R_160a_17010ce8 , 
    R_891_13b8ab98 , 
    R_132b_1007f7d8 , 
    R_6ed_140b6538 , 
    R_118f_14b1ee78 , 
    R_194a_13d2ae18 , 
    R_d0c_13dee8b8 , 
    R_b70_13d20f58 , 
    R_17ae_13d29a18 , 
    R_1a3c_13b95278 , 
    R_109d_10084878 , 
    R_141d_13d441b8 , 
    R_16bc_14a0bdb8 , 
    R_dfe_15ff38e8 , 
    R_7df_1587d338 , 
    R_a7e_14a0bb38 , 
    R_151f_12fbe998 , 
    R_97c_13d528b8 , 
    R_15ba_1008b0d8 , 
    R_8e1_15889818 , 
    R_f00_17017ae8 , 
    R_f9b_13b974d8 , 
    R_16fa_14b299b8 , 
    R_10db_13cd6cb8 , 
    R_abc_15882b58 , 
    R_7a1_15ffcd08 , 
    R_dc0_117f53b8 , 
    R_13df_156b9238 , 
    R_19fe_13c01fd8 , 
    R_5cf_124c4678 , 
    R_12ad_13cca878 , 
    R_bee_156ac498 , 
    R_c8e_156b6cb8 , 
    R_120d_123be218 , 
    R_66f_13df8d18 , 
    R_182c_13b90598 , 
    R_18cc_170190c8 , 
    R_1505_13d27858 , 
    R_15d4_13d3a078 , 
    R_fb5_13c265b8 , 
    R_8c7_13ccf738 , 
    R_996_13cd1498 , 
    R_ee6_156ae158 , 
    R_1a0a_140b9238 , 
    R_13eb_150e7438 , 
    R_dcc_15815c78 , 
    R_7ad_1008c078 , 
    R_ab0_11629618 , 
    R_10cf_1580df78 , 
    R_16ee_123bf758 , 
    R_1660_13dd6258 , 
    R_83b_117f03b8 , 
    R_a22_156b92d8 , 
    R_1479_13ddc518 , 
    R_1041_14a0db18 , 
    R_e5a_11633118 , 
    R_1711_11c69d38 , 
    R_10f2_1486ad38 , 
    R_ad3_13d5a5b8 , 
    R_78a_13dfa2f8 , 
    R_da9_123bc9b8 , 
    R_13c8_11628e98 , 
    R_19e7_14a10098 , 
    R_eb5_13cd9cd8 , 
    R_fe6_13df1d38 , 
    R_14d4_13c27a58 , 
    R_9c7_140af5f8 , 
    R_896_123b6658 , 
    R_1605_156b1b78 , 
    R_1888_1580c858 , 
    R_1269_13b99c38 , 
    R_c4a_14a0cb78 , 
    R_62b_1162a1f8 , 
    R_613_124c47b8 , 
    R_c32_14b23518 , 
    R_1251_13d3fed8 , 
    R_1870_13b92bb8 , 
    R_16cc_156ba318 , 
    R_1a2c_156b08b8 , 
    R_140d_11638258 , 
    R_dee_13c0e058 , 
    R_7cf_123bbe78 , 
    R_a8e_170160a8 , 
    R_10ad_10082618 , 
    R_11b0_13b99f58 , 
    R_572_140ab458 , 
    R_6cc_117e8a78 , 
    R_130a_13dda498 , 
    R_17cf_13d389f8 , 
    R_b91_14b1f418 , 
    R_ceb_13d56d78 , 
    R_1929_13cd4af8 , 
    R_f72_13c2a1b8 , 
    R_953_14b20a98 , 
    R_90a_156ae658 , 
    R_f29_11630698 , 
    R_1548_140ac538 , 
    R_1591_13c25618 , 
    R_16fc_156b9a58 , 
    R_10dd_13d551f8 , 
    R_abe_14a15958 , 
    R_79f_140af7d8 , 
    R_dbe_13cd4c38 , 
    R_13dd_15884b38 , 
    R_19fc_13b96fd8 , 
    R_ff0_123b3b38 , 
    R_eab_11634518 , 
    R_9d1_13d4ed58 , 
    R_14ca_11631e58 , 
    R_160f_170102e8 , 
    R_88c_116319f8 , 
    R_e36_13c05b38 , 
    R_a46_11637e98 , 
    R_817_116294d8 , 
    R_1065_13c0b218 , 
    R_1455_117ef238 , 
    R_1684_13dd5ad8 , 
    R_e2b_13d28578 , 
    R_a51_11630ff8 , 
    R_80c_13d2acd8 , 
    R_1070_150e2d98 , 
    R_1a69_11c6fe18 , 
    R_168f_13d295b8 , 
    R_144a_1580c678 , 
    R_1a0c_13ccacd8 , 
    R_13ed_13cd4ff8 , 
    R_dce_14871f98 , 
    R_7af_11633578 , 
    R_aae_15814238 , 
    R_10cd_13d20878 , 
    R_16ec_13df6a18 , 
    R_1889_13bf9c38 , 
    R_126a_15886a78 , 
    R_c4b_13cd76b8 , 
    R_62c_10086038 , 
    R_612_10088dd8 , 
    R_c31_13b90778 , 
    R_1250_13d58c18 , 
    R_186f_1162dcb8 , 
    R_1a21_150e5598 , 
    R_1402_140b1cb8 , 
    R_de3_140b0778 , 
    R_7c4_13cd5138 , 
    R_a99_13cd0a98 , 
    R_10b8_13bea7d8 , 
    R_16d7_15888a58 , 
    R_b23_1587bc18 , 
    R_d59_14868cb8 , 
    R_1378_14b28158 , 
    R_1761_11631f98 , 
    R_1997_13d45158 , 
    R_1142_117f06d8 , 
    R_73a_13de1158 , 
    R_1a35_1486d7b8 , 
    R_16c3_13c01498 , 
    R_1416_1162ee38 , 
    R_df7_117f35b8 , 
    R_7d8_156abc78 , 
    R_a85_17014168 , 
    R_10a4_1486b0f8 , 
    R_a59_14a1a1d8 , 
    R_e23_13df5f78 , 
    R_1078_1580f558 , 
    R_804_156b6f38 , 
    R_1697_13d59d98 , 
    R_1a61_14a195f8 , 
    R_1442_14a18c98 , 
    R_1096_13dd6f78 , 
    R_1424_13b906d8 , 
    R_16b5_13c045f8 , 
    R_e05_140ad938 , 
    R_7e6_1486dd58 , 
    R_a77_100895f8 , 
    R_1a43_170104c8 , 
    R_15ef_15889318 , 
    R_ecb_13df7198 , 
    R_14ea_13cd2078 , 
    R_fd0_13cd59f8 , 
    R_8ac_15889278 , 
    R_9b1_1008a3b8 , 
    R_cc2_14a11218 , 
    R_17f8_13c28d18 , 
    R_59b_15812bb8 , 
    R_1900_1486c318 , 
    R_6a3_11c69658 , 
    R_bba_13deb7f8 , 
    R_12e1_123bbf18 , 
    R_11d9_14a18518 , 
    R_1125_124c3e58 , 
    R_d76_156b6218 , 
    R_b06_14b24af8 , 
    R_1395_13c0d978 , 
    R_19b4_14a10598 , 
    R_1744_11c6e3d8 , 
    R_757_13d3ceb8 , 
    R_16fe_123b51b8 , 
    R_10df_156b31f8 , 
    R_ac0_123c19b8 , 
    R_79d_13ddd698 , 
    R_dbc_13d207d8 , 
    R_13db_13d412d8 , 
    R_19fa_140afeb8 , 
    R_188a_14a0dd98 , 
    R_126b_170193e8 , 
    R_c4c_14874a18 , 
    R_62d_123c23b8 , 
    R_611_156aa558 , 
    R_c30_13cd8158 , 
    R_124f_13cd9418 , 
    R_186e_1162cb38 , 
    R_1233_13d5c318 , 
    R_1852_11635698 , 
    R_18a6_15885218 , 
    R_1287_13c29e98 , 
    R_c68_12fc1cd8 , 
    R_649_150e1f38 , 
    R_5f5_13bf7398 , 
    R_c14_13defe98 , 
    R_18c2_13d5d998 , 
    R_bf8_13bf77f8 , 
    R_12a3_14b20278 , 
    R_1217_123bdd18 , 
    R_c84_123bee98 , 
    R_1836_14a16038 , 
    R_665_117eefb8 , 
    R_5d9_15fed588 , 
    R_84f_1587bdf8 , 
    R_148d_156b2d98 , 
    R_164c_156b65d8 , 
    R_a0e_13cd5098 , 
    R_e6e_13c1e818 , 
    R_102d_14a14878 , 
    R_d7b_1007dbb8 , 
    R_1120_13cd3158 , 
    R_139a_12fbf398 , 
    R_b01_1587af98 , 
    R_19b9_116327b8 , 
    R_75c_13d54b18 , 
    R_173f_14a0d1b8 , 
    R_ca0_117f3978 , 
    R_bdc_14867a98 , 
    R_11fb_13d26638 , 
    R_681_13c02c58 , 
    R_18de_1162c638 , 
    R_181a_15887fb8 , 
    R_12bf_12fbe3f8 , 
    R_5bd_123b9678 , 
    R_1a0e_1486b698 , 
    R_13ef_156ba1d8 , 
    R_dd0_12fc0798 , 
    R_7b1_14a13478 , 
    R_aac_116311d8 , 
    R_10cb_150dccb8 , 
    R_16ea_140b6cb8 , 
    R_ffe_13ccf198 , 
    R_e9d_13d27038 , 
    R_9df_14a17398 , 
    R_161d_13b962b8 , 
    R_14bc_117f0598 , 
    R_87e_140b08b8 , 
    R_5a1_13d446b8 , 
    R_cbc_12fc1b98 , 
    R_bc0_13dfb338 , 
    R_69d_11c69798 , 
    R_18fa_140b5098 , 
    R_11df_15880998 , 
    R_12db_156b4af8 , 
    R_17fe_1580f5f8 , 
    R_191b_13c25f78 , 
    R_580_1162b4b8 , 
    R_6be_158101d8 , 
    R_17dd_14872358 , 
    R_12fc_15813dd8 , 
    R_b9f_140b49b8 , 
    R_cdd_13bf42d8 , 
    R_11be_150e4378 , 
    R_eba_13d29158 , 
    R_fe1_13d2bef8 , 
    R_14d9_13c21338 , 
    R_9c2_116297f8 , 
    R_89b_117ed118 , 
    R_1600_117e96f8 , 
    R_585_14a19b98 , 
    R_1916_150e99b8 , 
    R_17e2_123c1d78 , 
    R_6b9_150dc998 , 
    R_ba4_13c04d78 , 
    R_12f7_117f4ff8 , 
    R_11c3_117ee158 , 
    R_cd8_150deab8 , 
    R_15c4_13d46e18 , 
    R_8d7_13de10b8 , 
    R_fa5_13df4858 , 
    R_ef6_13c1f358 , 
    R_986_11631278 , 
    R_1515_13ccb8b8 , 
    R_11a7_123b9b78 , 
    R_569_12fbfd98 , 
    R_6d5_14b25958 , 
    R_1313_1587dab8 , 
    R_17c6_13d290b8 , 
    R_b88_14a0d9d8 , 
    R_cf4_13bea558 , 
    R_1932_13cd1538 , 
    R_1778_11631598 , 
    R_d42_1580f918 , 
    R_1159_148722b8 , 
    R_1361_14a18658 , 
    R_b3a_11637678 , 
    R_1980_15883a58 , 
    R_723_14a0aeb8 , 
    R_ec5_123c1eb8 , 
    R_fd6_15ff7448 , 
    R_14e4_14a121b8 , 
    R_9b7_117eaaf8 , 
    R_8a6_156b3018 , 
    R_15f5_140ade38 , 
    R_d45_117f4418 , 
    R_1775_140b5d18 , 
    R_1364_13c1d918 , 
    R_1156_15ff6fe8 , 
    R_1983_100863f8 , 
    R_726_13d39498 , 
    R_b37_10089b98 , 
    R_15e9_11636db8 , 
    R_14f0_13b92398 , 
    R_fca_156b44b8 , 
    R_8b2_11629078 , 
    R_9ab_14866698 , 
    R_ed1_158870b8 , 
    R_1632_117f1178 , 
    R_9f4_1486d2b8 , 
    R_e88_124c4498 , 
    R_1013_14a135b8 , 
    R_14a7_15814af8 , 
    R_869_14a19e18 , 
    R_132f_13c0b8f8 , 
    R_6f1_150df878 , 
    R_118b_14b27618 , 
    R_194e_14b236f8 , 
    R_d10_123b2d78 , 
    R_b6c_123b8138 , 
    R_17aa_13dfac58 , 
    R_188b_117e9978 , 
    R_126c_1580edd8 , 
    R_c4d_13d24b58 , 
    R_62e_13bf7438 , 
    R_610_14a186f8 , 
    R_c2f_14a0c038 , 
    R_124e_117ee338 , 
    R_186d_15fee348 , 
    R_e8c_1587e738 , 
    R_162e_123b25f8 , 
    R_9f0_140abe58 , 
    R_14ab_13dd50d8 , 
    R_86d_14a18dd8 , 
    R_100f_13d5dad8 , 
    R_8f8_15ff8668 , 
    R_f17_14a18e78 , 
    R_1536_14a0dc58 , 
    R_15a3_12fc08d8 , 
    R_f84_117e8d98 , 
    R_965_140b2578 , 
    R_d71_14b23018 , 
    R_b0b_13c21e78 , 
    R_1390_17016a08 , 
    R_19af_11636458 , 
    R_1749_117ec178 , 
    R_752_15ff64a8 , 
    R_112a_1587e0f8 , 
    R_18b6_13bf3018 , 
    R_1223_13dd8418 , 
    R_1297_13b99738 , 
    R_1842_123b43f8 , 
    R_c78_15887018 , 
    R_659_123b34f8 , 
    R_5e5_13df0578 , 
    R_c04_13cd6f38 , 
    R_954_17014988 , 
    R_909_13d3efd8 , 
    R_f28_13bf6fd8 , 
    R_1547_13df7b98 , 
    R_1592_156b9918 , 
    R_f73_13d22a38 , 
    R_70d_13beb098 , 
    R_178e_13c1cb58 , 
    R_196a_156b6d58 , 
    R_d2c_14a0ec98 , 
    R_116f_13d3e7b8 , 
    R_134b_15ff6cc8 , 
    R_b50_15815598 , 
    R_caf_156adc58 , 
    R_bcd_1162baf8 , 
    R_690_13c1e098 , 
    R_18ed_124c3278 , 
    R_11ec_1008d0b8 , 
    R_12ce_13c071b8 , 
    R_180b_1008abd8 , 
    R_5ae_13cd7ed8 , 
    R_177b_1007d6b8 , 
    R_d3f_13cd10d8 , 
    R_115c_150e8f18 , 
    R_135e_11c696f8 , 
    R_b3d_13dddeb8 , 
    R_720_13d395d8 , 
    R_197d_14a15458 , 
    R_1700_140ae8d8 , 
    R_10e1_13c07758 , 
    R_ac2_156ad2f8 , 
    R_79b_15886398 , 
    R_dba_116373f8 , 
    R_13d9_14a14378 , 
    R_19f8_117ef558 , 
    R_595_13def178 , 
    R_17f2_1580c998 , 
    R_1906_13ccad78 , 
    R_6a9_15ff4ba8 , 
    R_bb4_117f4d78 , 
    R_12e7_13cd42d8 , 
    R_11d3_1162b0f8 , 
    R_cc8_123b7738 , 
    R_d48_13c21c98 , 
    R_1772_14a16998 , 
    R_1367_15880858 , 
    R_1153_117f1678 , 
    R_1986_11c6c038 , 
    R_729_117f72f8 , 
    R_b34_158825b8 , 
    R_ff5_13c2a618 , 
    R_ea6_150dd7f8 , 
    R_9d6_13c01f38 , 
    R_14c5_14a0e518 , 
    R_1614_156b2b18 , 
    R_887_14a18298 , 
    R_848_13ddf218 , 
    R_1653_14869438 , 
    R_1486_156afe18 , 
    R_a15_1700ed08 , 
    R_e67_117f4e18 , 
    R_1034_156ac5d8 , 
    R_8eb_150db1d8 , 
    R_15b0_1580bdb8 , 
    R_f0a_14a0ce98 , 
    R_f91_117f6f38 , 
    R_1529_123bca58 , 
    R_972_13ccc038 , 
    R_1a10_123b4718 , 
    R_13f1_13d24298 , 
    R_dd2_14a19198 , 
    R_7b3_13c07938 , 
    R_aaa_13b8cfd8 , 
    R_10c9_15812a78 , 
    R_16e8_13cd8d38 , 
    R_d64_15ff5968 , 
    R_b18_117f40f8 , 
    R_1383_13c2a438 , 
    R_19a2_117f01d8 , 
    R_1756_123c0f18 , 
    R_1137_13d20ff8 , 
    R_745_13c1d5f8 , 
    R_1636_14b22618 , 
    R_9f8_13decdd8 , 
    R_e84_14875b98 , 
    R_1017_13d3bbf8 , 
    R_865_13d4e7b8 , 
    R_14a3_11c6d078 , 
    R_83e_13d43ad8 , 
    R_a1f_13d22d58 , 
    R_147c_1580d398 , 
    R_103e_13d57958 , 
    R_e5d_1486ddf8 , 
    R_165d_13bec038 , 
    R_1494_117f6718 , 
    R_1645_11c6c178 , 
    R_a07_14b251d8 , 
    R_e75_1580a5f8 , 
    R_1026_158103b8 , 
    R_856_13cd2a78 , 
    R_188c_13d39ad8 , 
    R_126d_11636638 , 
    R_c4e_13c0fe58 , 
    R_62f_116305f8 , 
    R_60f_13bf44b8 , 
    R_c2e_156b6c18 , 
    R_124d_123b5438 , 
    R_186c_15817758 , 
    R_57b_12fc1f58 , 
    R_6c3_14a11718 , 
    R_17d8_13bf24d8 , 
    R_1301_13ccee78 , 
    R_b9a_140b40f8 , 
    R_ce2_156b49b8 , 
    R_11b9_13d5d5d8 , 
    R_1920_117ea198 , 
    R_1713_14a0f878 , 
    R_10f4_13de4c18 , 
    R_ad5_117ed1b8 , 
    R_788_117e8ed8 , 
    R_da7_11635ff8 , 
    R_13c6_123c10f8 , 
    R_19e5_1580eb58 , 
    R_e90_11637038 , 
    R_9ec_117eb958 , 
    R_162a_117ec0d8 , 
    R_14af_156abdb8 , 
    R_871_1587f138 , 
    R_100b_11631d18 , 
    R_111b_1580faf8 , 
    R_139f_150df058 , 
    R_afc_117f8158 , 
    R_19be_13ccfff8 , 
    R_761_12fbf078 , 
    R_173a_156b5a98 , 
    R_d80_13c1d418 , 
    R_58a_13ddaf38 , 
    R_1911_124c4038 , 
    R_17e7_15883198 , 
    R_6b4_15881bb8 , 
    R_ba9_13d5c958 , 
    R_12f2_17013c68 , 
    R_11c8_11634fb8 , 
    R_cd3_13c06178 , 
    R_6fc_13de34f8 , 
    R_1180_13ddc298 , 
    R_1959_14a14698 , 
    R_d1b_13cd9558 , 
    R_b61_13d22538 , 
    R_179f_150e5818 , 
    R_133a_13d57138 , 
    R_be4_15817bb8 , 
    R_c98_13dec298 , 
    R_1203_1587d978 , 
    R_679_123b7918 , 
    R_1822_117e9018 , 
    R_18d6_13c2ad98 , 
    R_5c5_1162b5f8 , 
    R_12b7_117f83d8 , 
    R_ca8_14a11038 , 
    R_bd4_11637ad8 , 
    R_689_158869d8 , 
    R_11f3_116300f8 , 
    R_18e6_156b1678 , 
    R_1812_11c6f558 , 
    R_12c7_13b97c58 , 
    R_5b5_11637fd8 , 
    R_177e_14b1a738 , 
    R_d3c_13b8b278 , 
    R_115f_156ac7b8 , 
    R_135b_13d38b38 , 
    R_b40_158142d8 , 
    R_71d_13c1ea98 , 
    R_197a_13c0a318 , 
    R_e16_17018088 , 
    R_1085_13c03e78 , 
    R_7f7_15888b98 , 
    R_16a4_158821f8 , 
    R_1a54_13de0438 , 
    R_1435_10082258 , 
    R_a66_15882838 , 
    R_703_14867bd8 , 
    R_1960_1162c958 , 
    R_1179_13d3c7d8 , 
    R_d22_13d599d8 , 
    R_b5a_13bf68f8 , 
    R_1341_13d458d8 , 
    R_1798_1700e9e8 , 
    R_171e_13df60b8 , 
    R_10ff_13ddcab8 , 
    R_ae0_14a11f38 , 
    R_77d_13d27df8 , 
    R_d9c_13ccd4d8 , 
    R_13bb_1587d478 , 
    R_19da_13dd5a38 , 
    R_108a_1486e938 , 
    R_e11_13cd8c98 , 
    R_16a9_14a130b8 , 
    R_7f2_156b2938 , 
    R_1a4f_13d3a618 , 
    R_a6b_13b8e1f8 , 
    R_1430_13dd84b8 , 
    R_d4b_117f6178 , 
    R_176f_13d447f8 , 
    R_136a_13c26838 , 
    R_1150_15ff71c8 , 
    R_1989_13ccbc78 , 
    R_72c_10083c98 , 
    R_b31_13d44c58 , 
    R_814_13d51eb8 , 
    R_1068_1580ea18 , 
    R_1687_123b81d8 , 
    R_1452_13df0938 , 
    R_e33_14a0c3f8 , 
    R_a49_14a0eb58 , 
    R_1851_13d5b058 , 
    R_18a7_13b96858 , 
    R_1288_13c1daf8 , 
    R_c69_156af738 , 
    R_64a_11629438 , 
    R_5f4_140b13f8 , 
    R_c13_1162db78 , 
    R_1232_156aaa58 , 
    R_15bb_117f3338 , 
    R_8e0_14a0f698 , 
    R_f9c_14a104f8 , 
    R_eff_13d381d8 , 
    R_151e_15883af8 , 
    R_97d_14a16178 , 
    R_1702_13cd9198 , 
    R_10e3_117f2f78 , 
    R_ac4_1700f028 , 
    R_799_13d5a018 , 
    R_db8_150e6998 , 
    R_13d7_14b1d1b8 , 
    R_19f6_1580aa58 , 
    R_14fd_156b56d8 , 
    R_15dc_123bfd98 , 
    R_fbd_14a0b098 , 
    R_8bf_14875f58 , 
    R_99e_15ff9388 , 
    R_ede_11634338 , 
    R_188d_17018e48 , 
    R_126e_150e04f8 , 
    R_c4f_15814918 , 
    R_630_13d25558 , 
    R_60e_13cd3d38 , 
    R_c2d_1580aaf8 , 
    R_124c_13d40018 , 
    R_186b_13d42bd8 , 
    R_1a23_13d52458 , 
    R_1404_1486a8d8 , 
    R_de5_11633a78 , 
    R_7c6_156b9738 , 
    R_a97_13c05e58 , 
    R_10b6_124c3638 , 
    R_16d5_123bc4b8 , 
    R_bed_13b90db8 , 
    R_c8f_117ef4b8 , 
    R_120c_13ddcd38 , 
    R_670_13ccfaf8 , 
    R_182b_13cd80b8 , 
    R_18cd_13c1ca18 , 
    R_5ce_14b1ded8 , 
    R_12ae_13c1f178 , 
    R_bc6_13cd7bb8 , 
    R_697_13bf83d8 , 
    R_18f4_15881cf8 , 
    R_11e5_1162add8 , 
    R_12d5_17015928 , 
    R_1804_150e44b8 , 
    R_5a7_12fbe178 , 
    R_cb6_1162e398 , 
    R_110f_15887518 , 
    R_19ca_156b8a18 , 
    R_af0_17012a48 , 
    R_76d_156b1df8 , 
    R_d8c_15814b98 , 
    R_172e_117ed438 , 
    R_13ab_13b99878 , 
    R_1a12_13d52ef8 , 
    R_13f3_156b74d8 , 
    R_dd4_140ac5d8 , 
    R_7b5_13c1f718 , 
    R_aa8_14a0ea18 , 
    R_10c7_13df2c38 , 
    R_16e6_156b9eb8 , 
    R_15cd_13cd86f8 , 
    R_8ce_13d1e2f8 , 
    R_fae_13bf6df8 , 
    R_eed_15812578 , 
    R_98f_117f62b8 , 
    R_150c_15ff3848 , 
    R_908_123c0658 , 
    R_f27_13cd08b8 , 
    R_1546_14a18f18 , 
    R_1593_13d58e98 , 
    R_f74_158805d8 , 
    R_955_1580f0f8 , 
    R_d5c_1580ed38 , 
    R_137b_13d5cc78 , 
    R_175e_15813478 , 
    R_199a_117e8b18 , 
    R_113f_123b3098 , 
    R_73d_13c220f8 , 
    R_b20_13c06c18 , 
    R_163a_13d3ddb8 , 
    R_9fc_14a0b818 , 
    R_e80_11633ed8 , 
    R_101b_123b6518 , 
    R_861_124c3bd8 , 
    R_149f_123b5e38 , 
    R_1080_14a149b8 , 
    R_7fc_13d3f258 , 
    R_169f_124c2d78 , 
    R_1a59_117eded8 , 
    R_143a_14a0edd8 , 
    R_a61_1700dd68 , 
    R_e1b_13cd1178 , 
    R_140f_117f1cb8 , 
    R_df0_13c09cd8 , 
    R_7d1_14b28978 , 
    R_a8c_123c0338 , 
    R_10ab_13df0398 , 
    R_16ca_13d52f98 , 
    R_1a2e_13c22698 , 
    R_b10_14b21fd8 , 
    R_138b_156b0318 , 
    R_19aa_14a194b8 , 
    R_174e_15811a38 , 
    R_74d_117f0e58 , 
    R_112f_156aac38 , 
    R_d6c_156b62b8 , 
    R_1781_1162d5d8 , 
    R_d39_15811b78 , 
    R_1162_124c2558 , 
    R_1358_156b8e78 , 
    R_b43_13c06858 , 
    R_71a_117ee798 , 
    R_1977_15880b78 , 
    R_1108_13ccfb98 , 
    R_ae9_1580cd58 , 
    R_774_1700a7a8 , 
    R_d93_13cce0b8 , 
    R_13b2_15886898 , 
    R_1727_14870e18 , 
    R_19d1_123b5b18 , 
    R_188e_11c6a698 , 
    R_126f_14b23c98 , 
    R_c50_13d471d8 , 
    R_631_13ddd7d8 , 
    R_60d_117f3a18 , 
    R_c2c_13d2c498 , 
    R_124b_156b97d8 , 
    R_186a_13ddb118 , 
    R_fdc_1162ca98 , 
    R_14de_13c202f8 , 
    R_9bd_11632cb8 , 
    R_8a0_13bf81f8 , 
    R_15fb_123ba078 , 
    R_ebf_13b91678 , 
    R_e94_148719f8 , 
    R_9e8_15ff97e8 , 
    R_1626_13de2918 , 
    R_14b3_13dde9f8 , 
    R_875_156aea18 , 
    R_1007_15881578 , 
    R_14f6_11638938 , 
    R_fc4_1580d578 , 
    R_8b8_123ba2f8 , 
    R_9a5_117ecc18 , 
    R_ed7_14a0da78 , 
    R_15e3_123c0158 , 
    R_e0c_1700d0e8 , 
    R_16ae_123b38b8 , 
    R_7ed_117ef738 , 
    R_1a4a_12fc1c38 , 
    R_a70_150dbc78 , 
    R_142b_15889bd8 , 
    R_108f_13de36d8 , 
    R_d4e_11c6b6d8 , 
    R_176c_13ddfcb8 , 
    R_136d_11634dd8 , 
    R_114d_158861b8 , 
    R_198c_13d53a38 , 
    R_72f_11637498 , 
    R_b2e_170098a8 , 
    R_8f7_13b8e298 , 
    R_f16_1587d838 , 
    R_1535_13ded2d8 , 
    R_15a4_1162bcd8 , 
    R_f85_170174a8 , 
    R_966_156acd58 , 
    R_12a4_13cd0db8 , 
    R_1216_13c26518 , 
    R_c85_13d505b8 , 
    R_1835_13b8eb58 , 
    R_666_13cd8798 , 
    R_5d8_14a11fd8 , 
    R_18c3_156b8c98 , 
    R_bf7_156b4418 , 
    R_15d5_117ed898 , 
    R_fb6_14b24558 , 
    R_8c6_13d442f8 , 
    R_997_123bb478 , 
    R_ee5_14a14af8 , 
    R_1504_13d553d8 , 
    R_6d1_158167b8 , 
    R_130f_156ab4f8 , 
    R_17ca_150df9b8 , 
    R_b8c_124c3ef8 , 
    R_cf0_11c6a878 , 
    R_192e_150e8a18 , 
    R_11ab_13d29d38 , 
    R_56d_156b76b8 , 
    R_1704_13bf4238 , 
    R_10e5_14871778 , 
    R_ac6_1587bcb8 , 
    R_797_14b1c178 , 
    R_db6_13ddd058 , 
    R_13d5_1587c618 , 
    R_19f4_150e3ab8 , 
    R_1298_156b1d58 , 
    R_1841_13d2c538 , 
    R_c79_156b5598 , 
    R_65a_14874ab8 , 
    R_5e4_13bf0278 , 
    R_c03_14a0d2f8 , 
    R_18b7_13ccd1b8 , 
    R_1222_14b1acd8 , 
    R_1073_14b20f98 , 
    R_809_13d3e678 , 
    R_1a66_123b6158 , 
    R_1692_117f31f8 , 
    R_1447_13b93338 , 
    R_e28_156abbd8 , 
    R_a54_13cce838 , 
    R_1054_13bf8ab8 , 
    R_1466_13d5abf8 , 
    R_1673_1580e798 , 
    R_e47_1587b178 , 
    R_a35_117f5db8 , 
    R_828_10081f38 , 
    R_1469_1587ee18 , 
    R_1051_11635c38 , 
    R_e4a_11629118 , 
    R_1670_1007f238 , 
    R_82b_13cd7258 , 
    R_a32_1486afb8 , 
    R_1187_117f4198 , 
    R_1952_14a0c0d8 , 
    R_d14_13dee778 , 
    R_b68_10089d78 , 
    R_17a6_15811f38 , 
    R_1333_117f21b8 , 
    R_6f5_13d43678 , 
    R_6c8_1580d758 , 
    R_1306_1580d938 , 
    R_17d3_13d3a578 , 
    R_b95_117f7618 , 
    R_ce7_13d27218 , 
    R_1925_15ff0328 , 
    R_11b4_13b8ec98 , 
    R_576_13d2bf98 , 
    R_e00_13cd8bf8 , 
    R_7e1_150e4058 , 
    R_a7c_156b7118 , 
    R_1a3e_14a0b278 , 
    R_109b_123bd4f8 , 
    R_141f_1008c578 , 
    R_16ba_156b6e98 , 
    R_188f_156b5458 , 
    R_1270_14a103b8 , 
    R_c51_11630af8 , 
    R_632_13ccde38 , 
    R_60c_13dd9c78 , 
    R_c2b_14b23478 , 
    R_124a_140b7898 , 
    R_1869_14b29cd8 , 
    R_1a14_117ebbd8 , 
    R_13f5_13cd8a18 , 
    R_dd6_13de0d98 , 
    R_7b7_15816a38 , 
    R_aa6_13d28c58 , 
    R_10c5_11632998 , 
    R_16e4_10087078 , 
    R_190c_13d1d998 , 
    R_6af_124c33b8 , 
    R_bae_1587b5d8 , 
    R_12ed_14a176b8 , 
    R_11cd_13cd27f8 , 
    R_cce_116331b8 , 
    R_58f_156b9558 , 
    R_17ec_13dd7fb8 , 
    R_1057_123bd278 , 
    R_1463_124c4b78 , 
    R_1676_140ae6f8 , 
    R_e44_148741f8 , 
    R_a38_150dc3f8 , 
    R_825_123b3278 , 
    R_18a8_1580c8f8 , 
    R_1289_13c09738 , 
    R_c6a_15811fd8 , 
    R_64b_1007d938 , 
    R_5f3_116307d8 , 
    R_c12_1162cc78 , 
    R_1231_13dee9f8 , 
    R_1850_1587f778 , 
    R_146c_14872f38 , 
    R_104e_1580f7d8 , 
    R_e4d_14b20d18 , 
    R_166d_13d20058 , 
    R_82e_1580f2d8 , 
    R_a2f_123b3db8 , 
    R_19c3_116340b8 , 
    R_af7_13cd2d98 , 
    R_766_13c07618 , 
    R_1735_13bf9f58 , 
    R_d85_13dd7518 , 
    R_13a4_150ea138 , 
    R_1116_13c02438 , 
    R_df9_13dd9458 , 
    R_7da_14a16fd8 , 
    R_a83_13b9a278 , 
    R_10a2_123b3d18 , 
    R_1a37_1587f958 , 
    R_16c1_13d3d458 , 
    R_1418_13d2b1d8 , 
    R_ea1_156b5c78 , 
    R_9db_13c05bd8 , 
    R_1619_15888d78 , 
    R_14c0_17012fe8 , 
    R_882_13dee458 , 
    R_ffa_11c68f78 , 
    R_1967_15ff9608 , 
    R_1172_170122c8 , 
    R_d29_13bed898 , 
    R_1348_156b1178 , 
    R_b53_1162fe78 , 
    R_1791_15ff73a8 , 
    R_70a_13dee818 , 
    R_8ea_13b91c18 , 
    R_15b1_140b0d18 , 
    R_f09_13d4f9d8 , 
    R_f92_13b99238 , 
    R_1528_13cca918 , 
    R_973_12fc1738 , 
    R_907_13d1cef8 , 
    R_f26_13d51378 , 
    R_1545_13ddab78 , 
    R_1594_123b52f8 , 
    R_f75_1587ec38 , 
    R_956_117f3bf8 , 
    R_a1c_13d42098 , 
    R_147f_15ffd208 , 
    R_103b_12fbfbb8 , 
    R_e60_13b98dd8 , 
    R_165a_156b9418 , 
    R_841_13de1e78 , 
    R_1715_13c03ab8 , 
    R_10f6_1587fc78 , 
    R_ad7_11c6aaf8 , 
    R_786_13bf7938 , 
    R_da5_13c24c18 , 
    R_13c4_156adbb8 , 
    R_19e3_13b8b4f8 , 
    R_15c5_13cce478 , 
    R_8d6_14a156d8 , 
    R_fa6_13ccd7f8 , 
    R_ef5_13c0f8b8 , 
    R_987_148737f8 , 
    R_1514_13d4ea38 , 
    R_d36_13cd2938 , 
    R_1165_1700dae8 , 
    R_1355_13c0e2d8 , 
    R_b46_12fbedf8 , 
    R_717_13c1ebd8 , 
    R_1974_13b938d8 , 
    R_1784_14b1b3b8 , 
    R_156d_13b91d58 , 
    R_f4e_13d2bb38 , 
    R_156c_1486f8d8 , 
    R_92f_1587e418 , 
    R_f4d_158174d8 , 
    R_92e_15880df8 , 
    R_156e_13bee0b8 , 
    R_f4f_13d1f298 , 
    R_930_117f5818 , 
    R_156b_13cd6a38 , 
    R_f4c_13d4edf8 , 
    R_92d_13b93838 , 
    R_156f_1700c828 , 
    R_f50_13d5d038 , 
    R_931_1007f198 , 
    R_92c_13bef238 , 
    R_156a_14a0d7f8 , 
    R_f4b_1162df38 , 
    R_682_13dd6a78 , 
    R_11fa_12fbfe38 , 
    R_18df_1162e1b8 , 
    R_1819_117f44b8 , 
    R_12c0_156b3478 , 
    R_5bc_150db098 , 
    R_ca1_15888af8 , 
    R_bdb_123b9178 , 
    R_1890_13c0a4f8 , 
    R_1271_13cd3e78 , 
    R_c52_11629cf8 , 
    R_633_1587c6b8 , 
    R_60b_17014c08 , 
    R_c2a_13c01d58 , 
    R_1249_150de798 , 
    R_1868_13cd62b8 , 
    R_105a_14a112b8 , 
    R_1460_158862f8 , 
    R_1679_13cd44b8 , 
    R_e41_14a14e18 , 
    R_a3b_13cd1998 , 
    R_822_117e9158 , 
    R_1570_13d44118 , 
    R_f51_13ccb778 , 
    R_932_15810d18 , 
    R_92b_14a180b8 , 
    R_f4a_1162c8b8 , 
    R_1569_13bede38 , 
    R_163e_12fc0338 , 
    R_a00_13df4df8 , 
    R_e7c_13c08798 , 
    R_101f_117ed9d8 , 
    R_85d_117f4738 , 
    R_149b_13cd1038 , 
    R_146f_117f47d8 , 
    R_104b_158885f8 , 
    R_e50_12fbe858 , 
    R_166a_1587c938 , 
    R_831_156b2398 , 
    R_a2c_11c701d8 , 
    R_801_150e6e98 , 
    R_169a_13b94878 , 
    R_1a5e_1162d3f8 , 
    R_143f_13b8c218 , 
    R_a5c_13b8c178 , 
    R_e20_13ddd0f8 , 
    R_107b_156b2118 , 
    R_d51_13df3b38 , 
    R_1769_14b21038 , 
    R_1370_13cd2618 , 
    R_114a_13c218d8 , 
    R_198f_13d28bb8 , 
    R_732_13d55fb8 , 
    R_b2b_13ccd2f8 , 
    R_1571_1580af58 , 
    R_f52_12fc1ff8 , 
    R_933_14868718 , 
    R_92a_13c01a38 , 
    R_f49_13d4f4d8 , 
    R_1568_1580c218 , 
    R_1706_15814eb8 , 
    R_10e7_14a160d8 , 
    R_ac8_156afa58 , 
    R_795_14a12b18 , 
    R_db4_117edd98 , 
    R_13d3_13b90f98 , 
    R_19f2_12fbf258 , 
    R_17b9_156b0b38 , 
    R_193f_13d3aa78 , 
    R_b7b_13befeb8 , 
    R_d01_140ab318 , 
    R_119a_13b8a5f8 , 
    R_1320_14b27f78 , 
    R_55c_11630e18 , 
    R_6e2_158149b8 , 
    R_106b_117f3518 , 
    R_168a_117eb598 , 
    R_144f_14b26718 , 
    R_e30_123b3e58 , 
    R_a4c_170172c8 , 
    R_811_15882478 , 
    R_1406_148665f8 , 
    R_de7_1007fcd8 , 
    R_7c8_156b7f78 , 
    R_a95_117f6cb8 , 
    R_10b4_13d3d598 , 
    R_16d3_1700be28 , 
    R_1a25_13b9a318 , 
    R_1572_156b67b8 , 
    R_f53_123c01f8 , 
    R_934_156b0958 , 
    R_929_13d5bf58 , 
    R_f48_13c256b8 , 
    R_1567_13b91e98 , 
    R_1943_11c70598 , 
    R_d05_13c0cd98 , 
    R_b77_13d415f8 , 
    R_17b5_14a12118 , 
    R_1324_15887298 , 
    R_6e6_13becb78 , 
    R_558_116299d8 , 
    R_1196_13d4f398 , 
    R_e98_13d433f8 , 
    R_9e4_13cccdf8 , 
    R_1622_13c044b8 , 
    R_14b7_13d21318 , 
    R_879_15884c78 , 
    R_1003_124c39f8 , 
    R_1a16_1486b418 , 
    R_13f7_13d24338 , 
    R_dd8_1587fd18 , 
    R_7b9_13c0f458 , 
    R_aa4_13c1d0f8 , 
    R_10c3_13ccbef8 , 
    R_16e2_140b6df8 , 
    R_1573_14a0c498 , 
    R_f54_11632858 , 
    R_935_150e5318 , 
    R_928_156aab98 , 
    R_f47_13cd9238 , 
    R_1566_123b2a58 , 
    R_a0b_11637858 , 
    R_e71_14b21a38 , 
    R_102a_11c6ccb8 , 
    R_852_14b1d938 , 
    R_1490_13bf8158 , 
    R_1649_13dd4f98 , 
    R_a12_1008b358 , 
    R_e6a_156b7a78 , 
    R_1031_14b25778 , 
    R_84b_156ad1b8 , 
    R_1650_13dd4e58 , 
    R_1489_13c21978 , 
    R_7e8_1486a0b8 , 
    R_1a45_1162e2f8 , 
    R_a75_156b0778 , 
    R_1426_11637718 , 
    R_1094_13d28398 , 
    R_16b3_117efeb8 , 
    R_e07_13d453d8 , 
    R_17bd_1162b918 , 
    R_b7f_14a0be58 , 
    R_cfd_13d1d038 , 
    R_193b_13d39f38 , 
    R_119e_13c1bcf8 , 
    R_560_12fbf118 , 
    R_6de_13cd4058 , 
    R_131c_13c245d8 , 
    R_1891_123b9858 , 
    R_1272_13dd9ef8 , 
    R_c53_15ff5148 , 
    R_634_11631818 , 
    R_60a_156b2758 , 
    R_c29_13cd0598 , 
    R_1248_12fbfcf8 , 
    R_1867_14a0ded8 , 
    R_9cd_13d1f518 , 
    R_14ce_1008b5d8 , 
    R_160b_14b24cd8 , 
    R_890_11628df8 , 
    R_fec_13ccc5d8 , 
    R_eaf_13d5baf8 , 
    R_15bc_15889138 , 
    R_8df_11637358 , 
    R_f9d_158889b8 , 
    R_efe_11632b78 , 
    R_97e_13c29718 , 
    R_151d_1700bc48 , 
    R_ae2_123bdef8 , 
    R_77b_17011828 , 
    R_d9a_13c047d8 , 
    R_13b9_15ffc948 , 
    R_19d8_14870b98 , 
    R_1720_156b9198 , 
    R_1101_140b7398 , 
    R_1202_15881898 , 
    R_67a_13de2878 , 
    R_1821_117f1c18 , 
    R_18d7_1580f378 , 
    R_5c4_14868fd8 , 
    R_12b8_11631b38 , 
    R_be3_13de2198 , 
    R_c99_13c029d8 , 
    R_fd1_13c1d058 , 
    R_14e9_14868538 , 
    R_9b2_1580b6d8 , 
    R_8ab_14a0fc38 , 
    R_15f0_140ae3d8 , 
    R_eca_14a11df8 , 
    R_1574_13cd7cf8 , 
    R_f55_14b1ac38 , 
    R_936_140acf38 , 
    R_927_124c4178 , 
    R_f46_14a0af58 , 
    R_1565_1700e808 , 
    R_14d3_1580e5b8 , 
    R_9c8_15fef248 , 
    R_895_13d532b8 , 
    R_1606_1007ef18 , 
    R_eb4_117eda78 , 
    R_fe7_1162ba58 , 
    R_8f6_156b7b18 , 
    R_f15_158819d8 , 
    R_15a5_158168f8 , 
    R_1534_123b9c18 , 
    R_f86_13c1ce78 , 
    R_967_11c68938 , 
    R_1901_15817ed8 , 
    R_6a4_1162c1d8 , 
    R_bb9_156ab1d8 , 
    R_12e2_11636a98 , 
    R_11d8_156aa738 , 
    R_cc3_15887c98 , 
    R_59a_117f76b8 , 
    R_17f7_117e9838 , 
    R_105d_123b4998 , 
    R_145d_123bec18 , 
    R_167c_140b6178 , 
    R_e3e_150da7d8 , 
    R_a3e_11635cd8 , 
    R_81f_156b45f8 , 
    R_120b_13def358 , 
    R_671_140b4058 , 
    R_182a_117ef698 , 
    R_18ce_156b4e18 , 
    R_5cd_14a185b8 , 
    R_12af_15ff69a8 , 
    R_bec_124c2878 , 
    R_c90_117eb778 , 
    R_1386_14a0c7b8 , 
    R_19a5_1008a598 , 
    R_1753_13cd1218 , 
    R_748_13d3b518 , 
    R_1134_1580ad78 , 
    R_d67_13d3caf8 , 
    R_b15_156b2078 , 
    R_128a_15880718 , 
    R_c6b_14a13518 , 
    R_64c_148739d8 , 
    R_5f2_13dd5538 , 
    R_c11_15ff5aa8 , 
    R_1230_124c42b8 , 
    R_184f_1587fa98 , 
    R_18a9_11c6f918 , 
    R_bbf_1587ddd8 , 
    R_69e_123b5bb8 , 
    R_18fb_13df16f8 , 
    R_11de_10089058 , 
    R_12dc_13c0bc18 , 
    R_17fd_13d408d8 , 
    R_5a0_11631db8 , 
    R_cbd_14872df8 , 
    R_691_15883378 , 
    R_18ee_14a171b8 , 
    R_11eb_13d4f078 , 
    R_12cf_158850d8 , 
    R_180a_13d3fc58 , 
    R_5ad_14a0c2b8 , 
    R_cb0_13de1658 , 
    R_bcc_13df1f18 , 
    R_1472_13d3c698 , 
    R_1048_13df8bd8 , 
    R_e53_10087b18 , 
    R_1667_13beaf58 , 
    R_834_15888698 , 
    R_a29_13de0618 , 
    R_1575_13d42598 , 
    R_f56_13c0c578 , 
    R_937_15886c58 , 
    R_926_158846d8 , 
    R_f45_13d4f438 , 
    R_1564_1587b038 , 
    R_906_14a145f8 , 
    R_f25_13d24e78 , 
    R_1544_124c4fd8 , 
    R_1595_14b1f698 , 
    R_f76_117f6fd8 , 
    R_957_15888878 , 
    R_c7a_140ac998 , 
    R_65b_1580b778 , 
    R_5e3_117eba98 , 
    R_c02_123b2f58 , 
    R_18b8_12fc05b8 , 
    R_1221_15812cf8 , 
    R_1299_14b1fc38 , 
    R_1840_13d549d8 , 
    R_1947_156ac3f8 , 
    R_d09_150dd438 , 
    R_b73_117f7938 , 
    R_17b1_14a0dcf8 , 
    R_1328_13d2aeb8 , 
    R_6ea_123bbb58 , 
    R_1192_1587dbf8 , 
    R_137e_13c27738 , 
    R_175b_15883ff8 , 
    R_199d_1008a6d8 , 
    R_113c_13d20eb8 , 
    R_740_13bf6b78 , 
    R_b1d_123c1918 , 
    R_d5f_15888c38 , 
    R_fcb_13def8f8 , 
    R_8b1_170124a8 , 
    R_9ac_14a190f8 , 
    R_ed0_13d23d98 , 
    R_15ea_1580e658 , 
    R_14ef_123bead8 , 
    R_d33_123bd8b8 , 
    R_1168_156b6fd8 , 
    R_1352_13c10b78 , 
    R_b49_14a158b8 , 
    R_714_1587c898 , 
    R_1971_13ddfe98 , 
    R_1787_1486e2f8 , 
    R_68a_14a15b38 , 
    R_11f2_1162a6f8 , 
    R_18e7_13c08c98 , 
    R_1811_117e9a18 , 
    R_12c8_140aa878 , 
    R_5b4_140b2a78 , 
    R_ca9_15887e78 , 
    R_bd3_13c0e9b8 , 
    R_195d_15884818 , 
    R_117c_14874838 , 
    R_d1f_1007f698 , 
    R_b5d_123bb8d8 , 
    R_133e_13d55dd8 , 
    R_179b_12fbde58 , 
    R_700_13cd9878 , 
    R_1576_1700c6e8 , 
    R_f57_14a14198 , 
    R_938_13bedc58 , 
    R_925_13df1338 , 
    R_f44_156b99b8 , 
    R_1563_158841d8 , 
    R_c86_14a12e38 , 
    R_1834_13cd3f18 , 
    R_667_1486b558 , 
    R_5d7_156b0c78 , 
    R_18c4_11c709f8 , 
    R_bf6_11c6f378 , 
    R_12a5_1162d718 , 
    R_1215_117f51d8 , 
    R_1892_13d3b1f8 , 
    R_1273_13dd5c18 , 
    R_c54_13becd58 , 
    R_635_13d2c678 , 
    R_609_1580ef18 , 
    R_c28_140ba098 , 
    R_1247_13ccda78 , 
    R_1866_13bf9eb8 , 
    R_9d2_13ccb958 , 
    R_14c9_117f80b8 , 
    R_1610_1700a988 , 
    R_88b_1587e5f8 , 
    R_ff1_13b8bd18 , 
    R_eaa_13dd6618 , 
    R_1708_11630558 , 
    R_10e9_123c2138 , 
    R_aca_14a131f8 , 
    R_793_12fc2138 , 
    R_db2_123b68d8 , 
    R_13d1_156ac998 , 
    R_19f0_13d47138 , 
    R_7d3_13dd99f8 , 
    R_a8a_150e0ef8 , 
    R_10a9_1486ae78 , 
    R_16c8_13dfaed8 , 
    R_1a30_14a19698 , 
    R_1411_13dfa438 , 
    R_df2_150e09f8 , 
    R_14e3_11634838 , 
    R_9b8_13d43b78 , 
    R_8a5_13bee798 , 
    R_15f6_117f0458 , 
    R_ec4_11c68a78 , 
    R_fd7_116387f8 , 
    R_17c1_13d57d18 , 
    R_b83_13bedd98 , 
    R_cf9_1587d798 , 
    R_1937_150e3c98 , 
    R_11a2_13c05138 , 
    R_564_15815278 , 
    R_6da_13c00f98 , 
    R_1318_1008a9f8 , 
    R_faf_158866b8 , 
    R_8cd_15ff2ee8 , 
    R_eec_117f7078 , 
    R_990_11633c58 , 
    R_150b_13cd8dd8 , 
    R_15ce_13df0898 , 
    R_1766_116318b8 , 
    R_1373_15810598 , 
    R_1147_13b8d438 , 
    R_1992_13b8d1b8 , 
    R_735_13cd4cd8 , 
    R_b28_1162fab8 , 
    R_d54_150e15d8 , 
    R_1577_13d44ed8 , 
    R_f58_13d3e178 , 
    R_939_123b2878 , 
    R_924_140b7118 , 
    R_f43_140aeab8 , 
    R_1562_100874d8 , 
    R_17ce_13d50b58 , 
    R_b90_14a17e38 , 
    R_cec_156b8fb8 , 
    R_192a_13df93f8 , 
    R_11af_156b2a78 , 
    R_571_13b96ad8 , 
    R_6cd_150dc5d8 , 
    R_130b_14b1eab8 , 
    R_19b7_117f7758 , 
    R_75a_150de5b8 , 
    R_1741_100824d8 , 
    R_d79_1008a638 , 
    R_1122_150e9a58 , 
    R_1398_10083978 , 
    R_b03_158129d8 , 
    R_14d8_13cd4698 , 
    R_9c3_13befa58 , 
    R_89a_117edb18 , 
    R_1601_13d272b8 , 
    R_eb9_11638438 , 
    R_fe2_13defdf8 , 
    R_13f9_1580cb78 , 
    R_dda_117f7118 , 
    R_7bb_13bf54f8 , 
    R_aa2_12fc1a58 , 
    R_10c1_13b901d8 , 
    R_16e0_158811b8 , 
    R_1a18_156b8bf8 , 
    R_fbe_13cd90f8 , 
    R_8be_13df3278 , 
    R_99f_123b6b58 , 
    R_edd_13b99cd8 , 
    R_15dd_156aef18 , 
    R_14fc_140b09f8 , 
    R_19b2_150e0318 , 
    R_1746_123b75f8 , 
    R_755_14a13338 , 
    R_1127_13de3318 , 
    R_d74_17011d28 , 
    R_b08_150dce98 , 
    R_1393_11c68c58 , 
    R_1956_15813158 , 
    R_d18_156b9698 , 
    R_b64_156b3a18 , 
    R_17a2_117e8758 , 
    R_1337_13d20af8 , 
    R_6f9_17012b88 , 
    R_1183_1580f698 , 
    R_bb3_17013d08 , 
    R_12e8_14b1e158 , 
    R_11d2_124c3318 , 
    R_cc9_11c6e018 , 
    R_594_13cd9698 , 
    R_17f1_13c0bdf8 , 
    R_1907_13ccaa58 , 
    R_6aa_13de4038 , 
    R_ba3_13cd5bd8 , 
    R_12f8_13cd2758 , 
    R_11c2_13c1fc18 , 
    R_cd9_14b1f878 , 
    R_584_12fc0bf8 , 
    R_1917_13d21f98 , 
    R_17e1_13d37878 , 
    R_6ba_11637b78 , 
    R_8e9_13cd6b78 , 
    R_15b2_117f08b8 , 
    R_f08_156b5db8 , 
    R_f93_13b92758 , 
    R_1527_13ccaeb8 , 
    R_974_13c0c2f8 , 
    R_ad9_150e2a78 , 
    R_784_13dfa4d8 , 
    R_da3_14a0cd58 , 
    R_13c2_13d2a4b8 , 
    R_19e1_1700c5a8 , 
    R_1717_13df61f8 , 
    R_10f8_156b7258 , 
    R_1578_123bab18 , 
    R_f59_13c10358 , 
    R_93a_1486f978 , 
    R_923_11632178 , 
    R_f42_14b1f9b8 , 
    R_1561_13bf4a58 , 
    R_1060_13c0b358 , 
    R_145a_14a12bb8 , 
    R_167f_14a19378 , 
    R_e3b_13dd7f18 , 
    R_a41_14a10d18 , 
    R_81c_13bf79d8 , 
    R_12fd_1007d9d8 , 
    R_b9e_123ba618 , 
    R_cde_13d39218 , 
    R_11bd_11c6dcf8 , 
    R_191c_1580c038 , 
    R_57f_158160d8 , 
    R_6bf_13df4e98 , 
    R_17dc_15ff5508 , 
    R_1893_117f0d18 , 
    R_1274_156b1218 , 
    R_c55_13cce338 , 
    R_636_123c1238 , 
    R_608_13d58678 , 
    R_c27_13bf2a78 , 
    R_1246_14b229d8 , 
    R_1865_156b4d78 , 
    R_772_11634a18 , 
    R_d91_13c0fdb8 , 
    R_13b0_1486d0d8 , 
    R_1729_123b6338 , 
    R_19cf_11c70c78 , 
    R_110a_156b12b8 , 
    R_aeb_11638758 , 
    R_e78_117ef0f8 , 
    R_1023_15ff3ac8 , 
    R_859_13c0f098 , 
    R_1497_116337f8 , 
    R_1642_1162e578 , 
    R_a04_13c22e18 , 
    R_76b_13ddaad8 , 
    R_d8a_10085458 , 
    R_1730_11c6fd78 , 
    R_13a9_15887978 , 
    R_1111_11629c58 , 
    R_19c8_123b61f8 , 
    R_af2_11635558 , 
    R_1045_13c2abb8 , 
    R_e56_13c1f0d8 , 
    R_1664_1700d9a8 , 
    R_837_13d43c18 , 
    R_a26_13c28c78 , 
    R_1475_123b8bd8 , 
    R_e63_156b1358 , 
    R_1038_10085f98 , 
    R_1657_13cd2c58 , 
    R_844_117f3ab8 , 
    R_1482_140b29d8 , 
    R_a19_156ad4d8 , 
    R_18f5_1587d518 , 
    R_11e4_158159f8 , 
    R_12d6_11c6c5d8 , 
    R_1803_123b54d8 , 
    R_5a6_13ccf5f8 , 
    R_cb7_1162c458 , 
    R_bc5_14a0c5d8 , 
    R_698_14a0feb8 , 
    R_194b_15882658 , 
    R_d0d_1580bef8 , 
    R_b6f_117eb638 , 
    R_17ad_156b4f58 , 
    R_132c_158823d8 , 
    R_6ee_14a0faf8 , 
    R_118e_156ab3b8 , 
    R_75f_14870918 , 
    R_173c_123b9218 , 
    R_d7e_11634018 , 
    R_111d_13beeb58 , 
    R_139d_100868f8 , 
    R_afe_15ff7ee8 , 
    R_19bc_17010248 , 
    R_1175_11634c98 , 
    R_d26_1587cf78 , 
    R_b56_13c236d8 , 
    R_1345_13cd4738 , 
    R_1794_15813338 , 
    R_707_13d580d8 , 
    R_1964_13d42b38 , 
    R_f24_13b92938 , 
    R_1543_15ff0828 , 
    R_1596_15ff8a28 , 
    R_f77_158124d8 , 
    R_958_13df5bb8 , 
    R_905_13d4f758 , 
    R_1579_13b8d078 , 
    R_f5a_15884d18 , 
    R_93b_1580c3f8 , 
    R_922_140af198 , 
    R_f41_156b7cf8 , 
    R_1560_14a14cd8 , 
    R_c6c_14b20318 , 
    R_64d_13ccebf8 , 
    R_5f1_15814c38 , 
    R_c10_15817898 , 
    R_122f_13d22038 , 
    R_184e_14b1b8b8 , 
    R_18aa_11638b18 , 
    R_128b_1587eaf8 , 
    R_1695_14a12ed8 , 
    R_1a63_1486ec58 , 
    R_1444_15ff0788 , 
    R_a57_13d5aa18 , 
    R_e25_14a17078 , 
    R_1076_1587b678 , 
    R_806_14a0bd18 , 
    R_fb7_15887158 , 
    R_8c5_1008b2b8 , 
    R_998_13d573b8 , 
    R_ee4_15ff7da8 , 
    R_1503_150daf58 , 
    R_15d6_117ed398 , 
    R_7ca_150de978 , 
    R_a93_156af4b8 , 
    R_10b2_100826b8 , 
    R_16d1_156b27f8 , 
    R_1a27_13cd2118 , 
    R_1408_1587fbd8 , 
    R_de9_13cd12b8 , 
    R_9e0_15ffc9e8 , 
    R_161e_123b8a98 , 
    R_14bb_10081cb8 , 
    R_87d_123b9498 , 
    R_fff_12fbe5d8 , 
    R_e9c_13df34f8 , 
    R_ba8_123c12d8 , 
    R_12f3_11634f18 , 
    R_11c7_17013b28 , 
    R_cd4_13c2b018 , 
    R_589_14a19058 , 
    R_1912_156aacd8 , 
    R_17e6_140b2758 , 
    R_6b5_1587d658 , 
    R_f14_13d26458 , 
    R_15a6_1162eb18 , 
    R_1533_14b268f8 , 
    R_f87_11637998 , 
    R_968_13d2b958 , 
    R_8f5_13bebe58 , 
    R_8d5_150e1c18 , 
    R_fa7_12fbff78 , 
    R_ef4_1162ea78 , 
    R_988_15814198 , 
    R_1513_13c06498 , 
    R_15c6_12fbf2f8 , 
    R_8b7_15ffa468 , 
    R_9a6_13d46058 , 
    R_ed6_13d57598 , 
    R_15e4_156aeb58 , 
    R_14f5_13c29178 , 
    R_fc5_13b8d258 , 
    R_acc_13df8638 , 
    R_791_13d42818 , 
    R_db0_13bf9418 , 
    R_13cf_123c2318 , 
    R_19ee_11630cd8 , 
    R_170a_13d25698 , 
    R_10eb_13debbb8 , 
    R_19ad_1587f9f8 , 
    R_174b_15ff3528 , 
    R_750_1008c9d8 , 
    R_112c_13c015d8 , 
    R_d6f_117eae18 , 
    R_b0d_13d41c38 , 
    R_138e_158113f8 , 
    R_168d_156b2f78 , 
    R_144c_14a0dbb8 , 
    R_e2d_1587d3d8 , 
    R_a4f_15814418 , 
    R_80e_156ac218 , 
    R_106e_14a15318 , 
    R_157a_156b4198 , 
    R_f5b_1162d7b8 , 
    R_93c_13b933d8 , 
    R_921_15813298 , 
    R_f40_13cd1fd8 , 
    R_155f_148745b8 , 
    R_1275_13d26bd8 , 
    R_c56_12fbf438 , 
    R_637_14b20db8 , 
    R_607_15886258 , 
    R_c26_13d3ac58 , 
    R_1245_13d261d8 , 
    R_1864_13ddb2f8 , 
    R_1894_13cd6998 , 
    R_9d7_1580ac38 , 
    R_1615_150e0598 , 
    R_14c4_15ffa148 , 
    R_886_156aa9b8 , 
    R_ff6_13d424f8 , 
    R_ea5_13d23b18 , 
    R_1a51_13cda098 , 
    R_a69_123b4f38 , 
    R_1432_14b1d258 , 
    R_1088_13bec3f8 , 
    R_e13_140ab1d8 , 
    R_16a7_156afb98 , 
    R_7f4_14b238d8 , 
    R_17c5_12fc1058 , 
    R_b87_140b0db8 , 
    R_cf5_156ab818 , 
    R_1933_11633258 , 
    R_11a6_13c243f8 , 
    R_568_13ccd9d8 , 
    R_6d6_13ccc498 , 
    R_1314_13b93158 , 
    R_a81_11c6b098 , 
    R_10a0_148694d8 , 
    R_1a39_150e4cd8 , 
    R_16bf_13d3e8f8 , 
    R_141a_13ccc678 , 
    R_dfb_123b4c18 , 
    R_7dc_14b22578 , 
    R_116b_13ddcb58 , 
    R_134f_14b1c7b8 , 
    R_b4c_13d41eb8 , 
    R_711_140b8798 , 
    R_178a_13b96538 , 
    R_196e_150e3658 , 
    R_d30_13df5118 , 
    R_b99_13df2ff8 , 
    R_ce3_10088b58 , 
    R_11b8_156b8798 , 
    R_1921_13b91df8 , 
    R_57a_13ccb818 , 
    R_6c4_15887798 , 
    R_17d7_11c6faf8 , 
    R_1302_12fbe8f8 , 
    R_65c_117f0278 , 
    R_5e2_117ef198 , 
    R_c01_13df0118 , 
    R_18b9_13ded058 , 
    R_1220_117f77f8 , 
    R_129a_14a10ef8 , 
    R_183f_140b7f78 , 
    R_c7b_1580c178 , 
    R_7bd_12fc1558 , 
    R_aa0_11c6be58 , 
    R_10bf_13df54d8 , 
    R_16de_13de3138 , 
    R_1a1a_156b8ab8 , 
    R_13fb_156b4b98 , 
    R_ddc_11632df8 , 
    R_a7a_11c6b1d8 , 
    R_1a40_140b6d58 , 
    R_1099_116354b8 , 
    R_1421_117ef7d8 , 
    R_16b8_13d3ea38 , 
    R_e02_15ff37a8 , 
    R_7e3_15812118 , 
    R_1a56_13bf0818 , 
    R_1437_123bad98 , 
    R_a64_13beb318 , 
    R_e18_156afc38 , 
    R_1083_123c0a18 , 
    R_7f9_156b30b8 , 
    R_16a2_150e9418 , 
    R_18e0_13c201b8 , 
    R_1818_140b47d8 , 
    R_12c1_123bb838 , 
    R_5bb_156b5638 , 
    R_ca2_13dd9d18 , 
    R_bda_13b985b8 , 
    R_683_11634478 , 
    R_11f9_13ccd938 , 
    R_157b_1486f0b8 , 
    R_f5c_13de2378 , 
    R_93d_117f0ef8 , 
    R_920_13df90d8 , 
    R_f3f_13bf1a38 , 
    R_155e_123c0d38 , 
    R_8de_13d4e0d8 , 
    R_f9e_13b8a738 , 
    R_efd_123bfed8 , 
    R_97f_123c21d8 , 
    R_151c_13d5c4f8 , 
    R_15bd_13df43f8 , 
    R_1763_13d44618 , 
    R_1995_17017548 , 
    R_1144_17018948 , 
    R_738_1700bce8 , 
    R_b25_1162ad38 , 
    R_d57_13c242b8 , 
    R_1376_117f5098 , 
    R_9be_140aaaf8 , 
    R_89f_156b2ed8 , 
    R_15fc_13c28db8 , 
    R_ebe_13cd5c78 , 
    R_fdd_1162dd58 , 
    R_14dd_123b8db8 , 
    R_14aa_13c0f9f8 , 
    R_86c_13df77d8 , 
    R_1010_15884278 , 
    R_e8b_15880ad8 , 
    R_162f_15ff7808 , 
    R_9f1_123be718 , 
    R_1457_13d54758 , 
    R_1682_1587fb38 , 
    R_e38_150debf8 , 
    R_a44_1580d618 , 
    R_819_14873898 , 
    R_1063_13cd8978 , 
    R_1a4c_156b8b58 , 
    R_a6e_117ec3f8 , 
    R_142d_14b1c998 , 
    R_108d_14a0a878 , 
    R_e0e_156b9f58 , 
    R_16ac_13bf1218 , 
    R_7ef_1700c788 , 
    R_1014_13c079d8 , 
    R_868_1587de78 , 
    R_14a6_10081998 , 
    R_1633_117e9ab8 , 
    R_9f5_13d25c38 , 
    R_e87_15ff9ce8 , 
    R_1829_123b40d8 , 
    R_18cf_13ded238 , 
    R_5cc_156aa698 , 
    R_12b0_14a177f8 , 
    R_beb_13cca738 , 
    R_c91_15ff1cc8 , 
    R_120a_13cd9738 , 
    R_672_13c06fd8 , 
    R_779_13cd2258 , 
    R_d98_13b958b8 , 
    R_13b7_1700e308 , 
    R_19d6_117ecfd8 , 
    R_1722_123b5a78 , 
    R_1103_117f7bb8 , 
    R_ae4_11634ab8 , 
    R_c57_15814f58 , 
    R_638_14a151d8 , 
    R_606_13d50838 , 
    R_c25_10083bf8 , 
    R_1244_13ddb898 , 
    R_1863_123b9f38 , 
    R_1895_13df3a98 , 
    R_1276_123bda98 , 
    R_1042_13cd6718 , 
    R_e59_1587dd38 , 
    R_1661_13de0758 , 
    R_83a_13d21598 , 
    R_a23_14869cf8 , 
    R_1478_13cd7618 , 
    R_668_11c6aff8 , 
    R_5d6_13d24158 , 
    R_18c5_123b5f78 , 
    R_bf5_123ba7f8 , 
    R_12a6_148674f8 , 
    R_1214_15886cf8 , 
    R_c87_13c21bf8 , 
    R_1833_117f3838 , 
    R_1820_14872a38 , 
    R_18d8_13b8ef18 , 
    R_5c3_10080778 , 
    R_12b9_140abb38 , 
    R_be2_13b98338 , 
    R_c9a_13cd1f38 , 
    R_1201_15ff65e8 , 
    R_67b_13c02bb8 , 
    R_1542_14a19cd8 , 
    R_1597_117ee478 , 
    R_f78_156af198 , 
    R_959_11631bd8 , 
    R_904_13bebbd8 , 
    R_f23_13c2b338 , 
    R_157c_14a0eab8 , 
    R_f5d_15817c58 , 
    R_93e_13cd6858 , 
    R_91f_117f7d98 , 
    R_f3e_1700a708 , 
    R_155d_1700fa28 , 
    R_764_150dee78 , 
    R_1737_13cd6538 , 
    R_d83_150dc678 , 
    R_1118_13cce3d8 , 
    R_13a2_13df95d8 , 
    R_af9_14b1bc78 , 
    R_19c1_15811358 , 
    R_14ae_14b22438 , 
    R_870_158800d8 , 
    R_100c_14b1bef8 , 
    R_e8f_13c27cd8 , 
    R_9ed_150e3a18 , 
    R_162b_13d24478 , 
    R_64e_12fbeb78 , 
    R_5f0_13d25738 , 
    R_c0f_1587ef58 , 
    R_122e_14a181f8 , 
    R_184d_1486ac98 , 
    R_18ab_13bf9d78 , 
    R_128c_11c6a378 , 
    R_c6d_13d3be78 , 
    R_d11_117f09f8 , 
    R_b6b_13c0e878 , 
    R_17a9_15ff62c8 , 
    R_1330_1580d6b8 , 
    R_6f2_123ba398 , 
    R_118a_13c1eef8 , 
    R_194f_13c0e738 , 
    R_1758_14a14eb8 , 
    R_19a0_13c204d8 , 
    R_1139_117ef878 , 
    R_743_13d5a478 , 
    R_b1a_13c01038 , 
    R_d62_15811df8 , 
    R_1381_123b3a98 , 
    R_e6d_123b7238 , 
    R_102e_150ddd98 , 
    R_84e_15883418 , 
    R_164d_14a0c678 , 
    R_148c_1580e8d8 , 
    R_a0f_15ffbae8 , 
    R_12ee_13d3d958 , 
    R_11cc_14a11a38 , 
    R_ccf_15812258 , 
    R_58e_150e4558 , 
    R_17eb_150e6538 , 
    R_190d_14b294b8 , 
    R_6b0_14a172f8 , 
    R_bad_15883c38 , 
    R_1018_13d2a878 , 
    R_864_13c09238 , 
    R_14a2_13cd9e18 , 
    R_1637_1162fbf8 , 
    R_9f9_156b7438 , 
    R_e83_15886438 , 
    R_1a5b_13df6158 , 
    R_143c_15ff2a88 , 
    R_a5f_13df1518 , 
    R_e1d_13c288b8 , 
    R_107e_13c1c298 , 
    R_7fe_117f30b8 , 
    R_169d_156abf98 , 
    R_15b3_13cd6e98 , 
    R_f07_13b953b8 , 
    R_f94_13d25198 , 
    R_1526_1486bf58 , 
    R_975_13d529f8 , 
    R_8e8_117f0bd8 , 
    R_78f_1162c9f8 , 
    R_dae_11c6d578 , 
    R_13cd_14a162b8 , 
    R_19ec_15814738 , 
    R_170c_13ccdd98 , 
    R_10ed_15882dd8 , 
    R_ace_15885cb8 , 
    R_157d_13cd56d8 , 
    R_f5e_140b53b8 , 
    R_93f_13d57778 , 
    R_91e_15886f78 , 
    R_f3d_11634798 , 
    R_155c_156adf78 , 
    R_782_15ffd168 , 
    R_da1_14b290f8 , 
    R_13c0_117f6b78 , 
    R_19df_117eb318 , 
    R_1719_13c1f8f8 , 
    R_10fa_13decd38 , 
    R_adb_17014708 , 
    R_a88_13cd40f8 , 
    R_10a7_117eb1d8 , 
    R_16c6_158880f8 , 
    R_1a32_15818018 , 
    R_1413_13d57ef8 , 
    R_df4_17013f88 , 
    R_7d5_15889098 , 
    R_639_13df0cf8 , 
    R_605_14b1c3f8 , 
    R_c24_11632d58 , 
    R_1243_158151d8 , 
    R_1862_140b94b8 , 
    R_1896_13c0a598 , 
    R_1277_13c27378 , 
    R_c58_13dddc38 , 
    R_15a7_17013448 , 
    R_1532_156b4ff8 , 
    R_f88_13d225d8 , 
    R_969_13cce298 , 
    R_8f4_156b9af8 , 
    R_f13_13c2b478 , 
    R_1750_14a13018 , 
    R_74b_123b9998 , 
    R_1131_13d21c78 , 
    R_d6a_13c0c118 , 
    R_b12_1587bb78 , 
    R_1389_13c2a4d8 , 
    R_19a8_124c5578 , 
    R_a9e_13de43f8 , 
    R_10bd_1162e6b8 , 
    R_16dc_14b1f058 , 
    R_1a1c_13cda138 , 
    R_13fd_14a0e0b8 , 
    R_dde_15ffc448 , 
    R_7bf_123bb0b8 , 
    R_1027_13c277d8 , 
    R_855_14a117b8 , 
    R_1493_13bee3d8 , 
    R_1646_13ccbdb8 , 
    R_a08_15ffa5a8 , 
    R_e74_123b4678 , 
    R_12d0_14a11cb8 , 
    R_1809_13d4f7f8 , 
    R_5ac_11c6e838 , 
    R_cb1_13d2c998 , 
    R_bcb_1007e3d8 , 
    R_692_1587be98 , 
    R_18ef_13d28758 , 
    R_11ea_1580f238 , 
    R_991_1007ff58 , 
    R_eeb_12fbe0d8 , 
    R_150a_14a0b3b8 , 
    R_15cf_10085958 , 
    R_fb0_117f5318 , 
    R_8cc_13bf3338 , 
    R_ce8_11c6a7d8 , 
    R_1926_116372b8 , 
    R_11b3_13cd3fb8 , 
    R_575_15817438 , 
    R_6c9_13dee318 , 
    R_1307_15ff2da8 , 
    R_17d2_156b8978 , 
    R_b94_1587e198 , 
    R_1810_117f12b8 , 
    R_12c9_17017868 , 
    R_5b3_123baa78 , 
    R_caa_15fedbc8 , 
    R_bd2_1580d9d8 , 
    R_68b_13ddf038 , 
    R_11f1_13c2a938 , 
    R_18e8_123bd638 , 
    R_157e_13dee278 , 
    R_f5f_1162d038 , 
    R_940_1486f838 , 
    R_91d_14b1cdf8 , 
    R_f3c_148682b8 , 
    R_155b_12fc0158 , 
    R_14b2_15ff2628 , 
    R_874_123c0298 , 
    R_1008_1587dc98 , 
    R_e93_13cd4878 , 
    R_9e9_123b4498 , 
    R_1627_156b7578 , 
    R_cf1_124c34f8 , 
    R_192f_14a12cf8 , 
    R_11aa_117e9bf8 , 
    R_56c_140ab598 , 
    R_6d2_1162ec58 , 
    R_1310_13ddf538 , 
    R_17c9_11638578 , 
    R_b8b_13df36d8 , 
    R_a91_13ccfeb8 , 
    R_10b0_117ea418 , 
    R_16cf_11c6b138 , 
    R_1a29_13d384f8 , 
    R_140a_140aa5f8 , 
    R_deb_140b71b8 , 
    R_7cc_13cd94b8 , 
    R_1a47_100862b8 , 
    R_a73_123be538 , 
    R_1428_13dde3b8 , 
    R_1092_15ff41a8 , 
    R_e09_15887a18 , 
    R_16b1_13c0c258 , 
    R_7ea_11c6e518 , 
    R_e66_170138a8 , 
    R_1035_1162a478 , 
    R_847_14a15a98 , 
    R_1654_1580fff8 , 
    R_1485_117f6358 , 
    R_a16_14b25638 , 
    R_b60_13b97b18 , 
    R_179e_156b3c98 , 
    R_133b_13ddde18 , 
    R_6fd_156b8338 , 
    R_117f_13cd7578 , 
    R_195a_150e1218 , 
    R_d1c_13d3fd98 , 
    R_134c_14a11ad8 , 
    R_b4f_12fbee98 , 
    R_70e_124c25f8 , 
    R_178d_11638a78 , 
    R_196b_1580a918 , 
    R_d2d_13cd54f8 , 
    R_116e_117ebb38 , 
    R_5e1_14b286f8 , 
    R_c00_150df558 , 
    R_18ba_11638bb8 , 
    R_121f_13dfa1b8 , 
    R_129b_13cd3298 , 
    R_183e_1587c398 , 
    R_c7c_11c6a558 , 
    R_65d_13cd74d8 , 
    R_9b3_13df8138 , 
    R_8aa_13dd9a98 , 
    R_15f1_156b5d18 , 
    R_ec9_1587c1b8 , 
    R_fd2_13c05098 , 
    R_14e8_1700a528 , 
    R_11dd_14875918 , 
    R_12dd_14a0e158 , 
    R_17fc_11635eb8 , 
    R_59f_14a14c38 , 
    R_cbe_116357d8 , 
    R_bbe_15881438 , 
    R_18fc_17009bc8 , 
    R_69f_13d56b98 , 
    R_1598_13cd92d8 , 
    R_f79_13bf2e38 , 
    R_95a_13d37698 , 
    R_903_117ec7b8 , 
    R_f22_14a13978 , 
    R_1541_15886758 , 
    R_12e3_17014028 , 
    R_11d7_1587d5b8 , 
    R_cc4_13bead78 , 
    R_599_150dcf38 , 
    R_17f6_117f1498 , 
    R_1902_14b1af58 , 
    R_6a5_13df56b8 , 
    R_bb8_124c3b38 , 
    R_14bf_150dd938 , 
    R_881_150db278 , 
    R_ffb_15813ab8 , 
    R_ea0_13b95778 , 
    R_9dc_15ff19a8 , 
    R_161a_14b23bf8 , 
    R_1454_123b4538 , 
    R_e35_11c70098 , 
    R_a47_1486f3d8 , 
    R_816_13c06cb8 , 
    R_1066_13bee838 , 
    R_1685_15ff1d68 , 
    R_8b0_15813c98 , 
    R_9ad_13de0bb8 , 
    R_ecf_13c26798 , 
    R_15eb_140b6498 , 
    R_14ee_13d5a298 , 
    R_fcc_150e33d8 , 
    R_101c_11c6ce98 , 
    R_860_14a17b18 , 
    R_149e_11c6edd8 , 
    R_163b_13c04b98 , 
    R_9fd_117ebf98 , 
    R_e7f_117f6038 , 
    R_604_15811718 , 
    R_c23_123bfc58 , 
    R_1242_10080c78 , 
    R_1861_12fbf7f8 , 
    R_1897_13d3d1d8 , 
    R_1278_117f4f58 , 
    R_c59_116304b8 , 
    R_63a_13c0a278 , 
    R_b59_15feff68 , 
    R_1342_148716d8 , 
    R_1797_117f7e38 , 
    R_704_123b2ff8 , 
    R_1961_1162de98 , 
    R_1178_13cd24d8 , 
    R_d23_11c68618 , 
    R_157f_13b8ce98 , 
    R_f60_140af9b8 , 
    R_941_13df8b38 , 
    R_91c_13df6d38 , 
    R_f3b_15810c78 , 
    R_155a_15882338 , 
    R_e5c_117f6df8 , 
    R_165e_117edf78 , 
    R_83d_13c24ad8 , 
    R_a20_15883738 , 
    R_147b_1700f5c8 , 
    R_103f_123b9ad8 , 
    R_5ef_1162a018 , 
    R_c0e_158802b8 , 
    R_122d_150e4eb8 , 
    R_184c_14a19418 , 
    R_18ac_117f13f8 , 
    R_128d_123b2af8 , 
    R_c6e_15ff6408 , 
    R_64f_13bf1ad8 , 
    R_9a0_13dd6078 , 
    R_edc_123be678 , 
    R_15de_15ff2268 , 
    R_14fb_13c29038 , 
    R_fbf_150e4f58 , 
    R_8bd_13cd5ef8 , 
    R_1998_14b279d8 , 
    R_1141_1580bbd8 , 
    R_73b_14a15638 , 
    R_b22_13cce8d8 , 
    R_d5a_13bf6178 , 
    R_1379_123bdbd8 , 
    R_1760_117f7f78 , 
    R_1981_1587b7b8 , 
    R_b39_15ffae68 , 
    R_724_117ec8f8 , 
    R_1777_1587ccf8 , 
    R_d43_13beedd8 , 
    R_1362_150dfcd8 , 
    R_1158_13bf0f98 , 
    R_770_15888058 , 
    R_d8f_11629f78 , 
    R_13ae_13bf3478 , 
    R_172b_156b88d8 , 
    R_19cd_117ed578 , 
    R_110c_15810458 , 
    R_aed_14a0e298 , 
    R_1449_14b26678 , 
    R_e2a_13c29858 , 
    R_a52_140af378 , 
    R_80b_158154f8 , 
    R_1071_123c1378 , 
    R_1a68_117ed618 , 
    R_1690_13c216f8 , 
    R_ef3_13cd06d8 , 
    R_989_13c068f8 , 
    R_1512_1162e078 , 
    R_15c7_13d3c4b8 , 
    R_8d4_123c1738 , 
    R_fa8_123be858 , 
    R_1984_1162e438 , 
    R_727_1700aca8 , 
    R_b36_123bb338 , 
    R_d46_13cd3338 , 
    R_1774_13c26c98 , 
    R_1365_150db818 , 
    R_1155_17012868 , 
    R_b3c_13cd4eb8 , 
    R_721_156b7d98 , 
    R_197e_13d5c8b8 , 
    R_177a_123c1418 , 
    R_d40_11635af8 , 
    R_115b_123bf2f8 , 
    R_135f_11c6da78 , 
    R_894_1587b2b8 , 
    R_1607_123bd138 , 
    R_eb3_123b5cf8 , 
    R_fe8_15816678 , 
    R_14d2_11636e58 , 
    R_9c9_13cce798 , 
    R_160c_117f74d8 , 
    R_88f_13c0d338 , 
    R_fed_12fc1198 , 
    R_eae_13cd1d58 , 
    R_9ce_1162c6d8 , 
    R_14cd_10081178 , 
    R_dac_14a109f8 , 
    R_13cb_13ccf0f8 , 
    R_19ea_11629b18 , 
    R_170e_1580e338 , 
    R_10ef_14a199b8 , 
    R_ad0_123b65b8 , 
    R_78d_15817618 , 
    R_999_1008a138 , 
    R_ee3_158135b8 , 
    R_1502_117ea238 , 
    R_15d7_11c6ab98 , 
    R_fb8_156b7bb8 , 
    R_8c4_117f8018 , 
    R_efc_12fc14b8 , 
    R_980_13d2b9f8 , 
    R_151b_14a153b8 , 
    R_15be_11629bb8 , 
    R_8dd_13d1dcb8 , 
    R_f9f_13bf1858 , 
    R_8a4_13cd4418 , 
    R_15f7_117ea878 , 
    R_ec3_14a15e58 , 
    R_fd8_117f1718 , 
    R_14e2_13ddc478 , 
    R_9b9_1008a458 , 
    R_1580_123b3958 , 
    R_f61_14867318 , 
    R_942_140b3a18 , 
    R_91b_156b0d18 , 
    R_f3a_1007f4b8 , 
    R_1559_13c234f8 , 
    R_1441_13ded378 , 
    R_a5a_13c097d8 , 
    R_e22_117eccb8 , 
    R_1079_13beb6d8 , 
    R_803_140b8158 , 
    R_1698_15811998 , 
    R_1a60_14b1b778 , 
    R_1987_140b7cf8 , 
    R_72a_158127f8 , 
    R_b33_13d2aaf8 , 
    R_d49_15811678 , 
    R_1771_17009c68 , 
    R_1368_1587e9b8 , 
    R_1152_13c0bd58 , 
    R_5d5_123be038 , 
    R_18c6_13d3a1b8 , 
    R_bf4_1587cb18 , 
    R_12a7_15817cf8 , 
    R_1213_140ad078 , 
    R_c88_17017cc8 , 
    R_1832_123bc2d8 , 
    R_669_116322b8 , 
    R_769_150da558 , 
    R_d88_117f22f8 , 
    R_1732_123b2558 , 
    R_13a7_13c08ab8 , 
    R_1113_123c1e18 , 
    R_19c6_13cd18f8 , 
    R_af4_1580feb8 , 
    R_b3f_13c22198 , 
    R_71e_140aec98 , 
    R_197b_123c14b8 , 
    R_177d_17012728 , 
    R_d3d_13c053b8 , 
    R_115e_15885c18 , 
    R_135c_13cda3b8 , 
    R_12d7_13cd2578 , 
    R_1802_13d3fbb8 , 
    R_5a5_13d375f8 , 
    R_cb8_11c6c218 , 
    R_bc4_14b2a138 , 
    R_699_15888ff8 , 
    R_18f6_124c27d8 , 
    R_11e3_1162fa18 , 
    R_b67_13cd4f58 , 
    R_17a5_116334d8 , 
    R_1334_13cd5598 , 
    R_6f6_117f1858 , 
    R_1186_11635d78 , 
    R_1953_117eb6d8 , 
    R_d15_123b5578 , 
    R_603_13ddbe38 , 
    R_c22_117f71b8 , 
    R_1241_1162a5b8 , 
    R_1860_13ccdf78 , 
    R_1898_11c6bb38 , 
    R_1279_15887478 , 
    R_c5a_14a16538 , 
    R_63b_15883cd8 , 
    R_10bb_1587d8d8 , 
    R_16da_124c3db8 , 
    R_1a1e_11c6ed38 , 
    R_13ff_17012c28 , 
    R_de0_13d3abb8 , 
    R_7c1_156b3bf8 , 
    R_a9c_1162e4d8 , 
    R_18d0_117f1358 , 
    R_5cb_12fc0d38 , 
    R_12b1_124c38b8 , 
    R_bea_13ccb098 , 
    R_c92_150e3838 , 
    R_1209_14a0aa58 , 
    R_673_14a13fb8 , 
    R_1828_1580ab98 , 
    R_14b6_1587d1f8 , 
    R_878_13c100d8 , 
    R_1004_156ab318 , 
    R_e97_14866918 , 
    R_9e5_1587d6f8 , 
    R_1623_13b96178 , 
    R_11d1_1162f6f8 , 
    R_cca_117eebf8 , 
    R_593_117ee0b8 , 
    R_17f0_100833d8 , 
    R_1908_1162f5b8 , 
    R_6ab_13ccbe58 , 
    R_bb2_15810278 , 
    R_12e9_13d26818 , 
    R_f89_13d51738 , 
    R_96a_1587c258 , 
    R_8f3_10082b18 , 
    R_f12_1162b2d8 , 
    R_15a8_14b25db8 , 
    R_1531_13c0ac78 , 
    R_12c2_13d4e2b8 , 
    R_5ba_13b94d78 , 
    R_ca3_13ddaa38 , 
    R_bd9_13d54398 , 
    R_684_117f5a98 , 
    R_11f8_13bf1538 , 
    R_18e1_17010388 , 
    R_1817_1580f9b8 , 
    R_a7f_117ebc78 , 
    R_1a3b_13d275d8 , 
    R_109e_14a11538 , 
    R_16bd_117eb9f8 , 
    R_141c_123b3f98 , 
    R_dfd_1700cf08 , 
    R_7de_15881ed8 , 
    R_f95_13d51058 , 
    R_1525_140b5598 , 
    R_976_140b2f78 , 
    R_8e7_13dd8ff8 , 
    R_15b4_13dee598 , 
    R_f06_14b29238 , 
    R_899_13d5a8d8 , 
    R_1602_13c28ef8 , 
    R_eb8_13c1c0b8 , 
    R_fe3_13ccb598 , 
    R_14d7_14a0fb98 , 
    R_9c4_123c1a58 , 
    R_1599_13bf40f8 , 
    R_f7a_13d510f8 , 
    R_95b_15813838 , 
    R_902_14a0aff8 , 
    R_f21_15812398 , 
    R_1540_14871458 , 
    R_1321_156b1038 , 
    R_1199_13cd3bf8 , 
    R_6e3_140b27f8 , 
    R_55b_13d54f78 , 
    R_1940_117ed758 , 
    R_17b8_14b1ca38 , 
    R_d02_14b21998 , 
    R_b7a_140b8298 , 
    R_ed5_123b27d8 , 
    R_15e5_13d3e0d8 , 
    R_14f4_1580cad8 , 
    R_fc6_117f2078 , 
    R_8b6_12fbe7b8 , 
    R_9a7_13dd6118 , 
    R_d96_13c23778 , 
    R_13b5_124c31d8 , 
    R_19d4_123b6798 , 
    R_1724_117edcf8 , 
    R_1105_158130b8 , 
    R_ae6_14873e38 , 
    R_777_17012228 , 
    R_1581_10080458 , 
    R_f62_13ccaff8 , 
    R_943_156b21b8 , 
    R_91a_13d23e38 , 
    R_f39_117f5778 , 
    R_1558_15ffb2c8 , 
    R_88a_15880c18 , 
    R_ff2_13d42638 , 
    R_ea9_15810ef8 , 
    R_9d3_12fc1e18 , 
    R_14c8_13d50d38 , 
    R_1611_13df2b98 , 
    R_5c2_150db138 , 
    R_12ba_158138d8 , 
    R_be1_10082898 , 
    R_c9b_13b977f8 , 
    R_1200_13d3d778 , 
    R_67c_13dec978 , 
    R_181f_156b4558 , 
    R_18d9_117f3e78 , 
    R_1743_15ff3488 , 
    R_758_13cd0ef8 , 
    R_1124_14a17d98 , 
    R_d77_14a0ca38 , 
    R_1396_156ace98 , 
    R_b05_13d37d78 , 
    R_19b5_13cd3c98 , 
    R_d9f_1580b818 , 
    R_13be_156af5f8 , 
    R_19dd_13d56238 , 
    R_171b_14a0ac38 , 
    R_10fc_13d52c78 , 
    R_add_17015ce8 , 
    R_780_13cd31f8 , 
    R_198a_12fc1af8 , 
    R_72d_13d467d8 , 
    R_b30_156ac358 , 
    R_d4c_11633d98 , 
    R_176e_12fbe678 , 
    R_136b_15810638 , 
    R_114f_123ba1b8 , 
    R_119d_123ba578 , 
    R_55f_13cce658 , 
    R_6df_13bf5ef8 , 
    R_131d_14a11c18 , 
    R_17bc_15886d98 , 
    R_b7e_123b7eb8 , 
    R_cfe_123b7418 , 
    R_193c_123b6298 , 
    R_b42_116296b8 , 
    R_71b_13cd8fb8 , 
    R_1978_1587e698 , 
    R_1780_1587b718 , 
    R_d3a_117f6678 , 
    R_1161_13beb3b8 , 
    R_1359_11c6d9d8 , 
    R_1325_156ac178 , 
    R_6e7_15882fb8 , 
    R_557_15885f38 , 
    R_1195_116363b8 , 
    R_1944_124c2918 , 
    R_d06_13dde818 , 
    R_b76_13d41b98 , 
    R_17b4_13d29ab8 , 
    R_1020_117ed258 , 
    R_85c_1580fc38 , 
    R_149a_13bf0ef8 , 
    R_163f_13de4218 , 
    R_a01_156b1498 , 
    R_e7b_1486b738 , 
    R_11c1_123b5618 , 
    R_cda_156b9878 , 
    R_1918_15880f38 , 
    R_583_13cccb78 , 
    R_17e0_14a15d18 , 
    R_6bb_117f2398 , 
    R_ba2_14a0e5b8 , 
    R_12f9_13d5c9f8 , 
    R_5ee_12fc0c98 , 
    R_c0d_13b93fb8 , 
    R_122c_14b217b8 , 
    R_18ad_13cd6358 , 
    R_184b_1486d3f8 , 
    R_128e_13b91a38 , 
    R_c6f_150e83d8 , 
    R_650_116346f8 , 
    R_5e0_13df04d8 , 
    R_bff_123b92b8 , 
    R_18bb_11c6f698 , 
    R_121e_14b1d438 , 
    R_129c_1007ebf8 , 
    R_183d_15882e78 , 
    R_c7d_13c108f8 , 
    R_65e_13d43998 , 
    R_75d_156ad118 , 
    R_173e_148678b8 , 
    R_d7c_123be998 , 
    R_111f_14a110d8 , 
    R_139b_156b35b8 , 
    R_b00_13ccf558 , 
    R_19ba_17014d48 , 
    R_a78_13cd1cb8 , 
    R_1a42_15817118 , 
    R_1097_13d240b8 , 
    R_1423_13c05a98 , 
    R_16b6_140aab98 , 
    R_e04_156b17b8 , 
    R_7e5_14b1e798 , 
    R_746_170166e8 , 
    R_1136_13d56558 , 
    R_d65_1008bb78 , 
    R_b17_123bcc38 , 
    R_1384_140b3298 , 
    R_19a3_117eaa58 , 
    R_1755_10087258 , 
    R_c21_1700d4a8 , 
    R_1240_11630238 , 
    R_185f_13bf7118 , 
    R_1899_156b1fd8 , 
    R_127a_14b28298 , 
    R_c5b_13d26278 , 
    R_63c_1587b538 , 
    R_602_156afff8 , 
    R_753_116336b8 , 
    R_1129_13ccc3f8 , 
    R_d72_13b95e58 , 
    R_b0a_156ad438 , 
    R_1391_15886578 , 
    R_19b0_17014a28 , 
    R_1748_117eeab8 , 
    R_e32_13c05c78 , 
    R_a4a_117e8bb8 , 
    R_813_11631318 , 
    R_1069_116369f8 , 
    R_1688_156b6a38 , 
    R_1451_150e6b78 , 
    R_cdf_150dfa58 , 
    R_11bc_11c6a9b8 , 
    R_191d_13c10678 , 
    R_57e_1162f338 , 
    R_6c0_13b98c98 , 
    R_17db_117f6858 , 
    R_12fe_116291b8 , 
    R_b9d_14872678 , 
    R_1349_13d26db8 , 
    R_b52_1162a978 , 
    R_1790_117e9798 , 
    R_70b_17018808 , 
    R_1968_13bf0318 , 
    R_d2a_15fef568 , 
    R_1171_117f5278 , 
    R_192b_11633cf8 , 
    R_11ae_123bc238 , 
    R_570_117ec218 , 
    R_6ce_13dee1d8 , 
    R_130c_15ff67c8 , 
    R_17cd_13b91858 , 
    R_b8f_14b25b38 , 
    R_ced_14a0a558 , 
    R_1582_150e7ed8 , 
    R_f63_13cca7d8 , 
    R_944_13d1fab8 , 
    R_919_123bdf98 , 
    R_f38_13d26958 , 
    R_1557_14a16c18 , 
    R_10ae_123b9358 , 
    R_16cd_117eee78 , 
    R_1a2b_140accb8 , 
    R_140c_11c6f058 , 
    R_ded_14a14738 , 
    R_7ce_13d45d38 , 
    R_a8f_17014de8 , 
    R_10a5_13d564b8 , 
    R_16c4_1580f878 , 
    R_1a34_14a19558 , 
    R_1415_158165d8 , 
    R_df6_156b2bb8 , 
    R_7d7_13c29998 , 
    R_a86_123bc0f8 , 
    R_165b_13de0898 , 
    R_840_156b26b8 , 
    R_a1d_14a15778 , 
    R_147e_11638078 , 
    R_103c_140b0ef8 , 
    R_e5f_150e3d38 , 
    R_11c6_13def038 , 
    R_cd5_13cd09f8 , 
    R_588_13de09d8 , 
    R_1913_13beef18 , 
    R_17e5_150de518 , 
    R_6b6_13d519b8 , 
    R_ba7_13d2ca38 , 
    R_12f4_11c6ca38 , 
    R_19e8_15888e18 , 
    R_1710_13bf6718 , 
    R_10f1_124c52f8 , 
    R_ad2_156b8658 , 
    R_78b_1162ddf8 , 
    R_daa_1008ced8 , 
    R_13c9_13de18d8 , 
    R_11a1_117e91f8 , 
    R_563_13d1ea78 , 
    R_6db_13dd91d8 , 
    R_1319_117f10d8 , 
    R_17c0_15ff4888 , 
    R_b82_13beff58 , 
    R_cfa_14b21ad8 , 
    R_1938_13df6ab8 , 
    R_82a_14a0cfd8 , 
    R_a33_11c70278 , 
    R_1468_158803f8 , 
    R_1052_117f42d8 , 
    R_1671_13dd6898 , 
    R_e49_15ff8f28 , 
    R_1329_14a16ad8 , 
    R_6eb_13d45b58 , 
    R_1191_15881618 , 
    R_1948_13c26a18 , 
    R_d0a_158820b8 , 
    R_b72_13c103f8 , 
    R_17b0_13decf18 , 
    R_a36_13b92438 , 
    R_827_123b8f98 , 
    R_1055_11635738 , 
    R_1465_14a18ab8 , 
    R_1674_11636c78 , 
    R_e46_15884098 , 
    R_851_11635238 , 
    R_148f_13df4358 , 
    R_164a_13c1e318 , 
    R_a0c_100899b8 , 
    R_e70_117ec538 , 
    R_102b_13d38d18 , 
    R_198d_156b4378 , 
    R_730_123bb518 , 
    R_b2d_124c29b8 , 
    R_d4f_13cd15d8 , 
    R_176b_150e5bd8 , 
    R_136e_15ff6b88 , 
    R_114c_140b06d8 , 
    R_16f5_13d39b78 , 
    R_1a03_14b23338 , 
    R_10d6_150df4b8 , 
    R_13e4_13cd99b8 , 
    R_ab7_1700b748 , 
    R_dc5_15ff3f28 , 
    R_7a6_150dad78 , 
    R_1a05_1162d498 , 
    R_13e6_1486e578 , 
    R_dc7_13cd2398 , 
    R_16f3_10088bf8 , 
    R_7a8_13beac38 , 
    R_10d4_13d1de98 , 
    R_ab5_13df25f8 , 
    R_82d_13c24b78 , 
    R_a30_117ef9b8 , 
    R_146b_150da9b8 , 
    R_104f_170118c8 , 
    R_e4c_13ddfd58 , 
    R_166e_123be3f8 , 
    R_73e_15883878 , 
    R_b1f_11631098 , 
    R_d5d_11636778 , 
    R_137c_11634e78 , 
    R_175d_13df13d8 , 
    R_199b_150dc8f8 , 
    R_113e_10081ad8 , 
    R_b45_13cce978 , 
    R_718_123b4fd8 , 
    R_1975_13deedb8 , 
    R_1783_15817e38 , 
    R_d37_13d26d18 , 
    R_1164_13df29b8 , 
    R_1356_15884958 , 
    R_16f7_140b9558 , 
    R_10d8_13d55158 , 
    R_ab9_14a16358 , 
    R_1a01_14a0bf98 , 
    R_7a4_13cca698 , 
    R_13e2_13d50338 , 
    R_dc3_13d5b918 , 
    R_1509_13c080b8 , 
    R_15d0_13d5d7b8 , 
    R_fb1_17011fa8 , 
    R_8cb_1162afb8 , 
    R_992_158117b8 , 
    R_eea_158843b8 , 
    R_1a07_15817f78 , 
    R_13e8_13d57458 , 
    R_dc9_13dedb98 , 
    R_7aa_14a113f8 , 
    R_ab3_13ccea18 , 
    R_16f1_13c2b298 , 
    R_10d2_14a0f4b8 , 
    R_84a_1700eee8 , 
    R_1651_100849b8 , 
    R_1488_15811858 , 
    R_a13_117f7ed8 , 
    R_e69_14b24ff8 , 
    R_1032_15884638 , 
    R_1434_15884a98 , 
    R_a67_1587c9d8 , 
    R_e15_117f6538 , 
    R_1086_158844f8 , 
    R_16a5_1587d018 , 
    R_7f6_14a10318 , 
    R_1a53_11c70b38 , 
    R_f7b_13c24f38 , 
    R_95c_13b8ad78 , 
    R_901_15ff0dc8 , 
    R_f20_11633078 , 
    R_153f_140abef8 , 
    R_159a_13d58d58 , 
    R_1a20_117f5638 , 
    R_1401_14a19918 , 
    R_de2_123bef38 , 
    R_7c3_14a0f058 , 
    R_a9a_15816f38 , 
    R_10b9_15ff6908 , 
    R_16d8_14b209f8 , 
    R_1583_13b8ba98 , 
    R_f64_123b9718 , 
    R_945_123bcaf8 , 
    R_918_13c20ed8 , 
    R_f37_158875b8 , 
    R_1556_140b5db8 , 
    R_a39_17016d28 , 
    R_824_140b4b98 , 
    R_1058_13b8c7b8 , 
    R_1462_13d228f8 , 
    R_1677_1008aef8 , 
    R_e43_140ab8b8 , 
    R_123f_12fc2458 , 
    R_185e_100815d8 , 
    R_189a_15ff14a8 , 
    R_127b_13de1a18 , 
    R_c5c_140b8518 , 
    R_63d_13df0438 , 
    R_601_14a12c58 , 
    R_c20_1486b7d8 , 
    R_15fd_156b4c38 , 
    R_ebd_117f1ad8 , 
    R_fde_13d429f8 , 
    R_14dc_13ddc5b8 , 
    R_9bf_15ff2128 , 
    R_89e_123bbdd8 , 
    R_16f9_13cd6218 , 
    R_10da_14a0d4d8 , 
    R_abb_14b262b8 , 
    R_7a2_13de1fb8 , 
    R_dc1_13c211f8 , 
    R_13e0_1486e4d8 , 
    R_19ff_123b42b8 , 
    R_1739_15ff78a8 , 
    R_d81_140ad4d8 , 
    R_111a_13d42ef8 , 
    R_13a0_117f2bb8 , 
    R_afb_13bf4af8 , 
    R_19bf_117f5e58 , 
    R_762_156b33d8 , 
    R_1a09_1162d358 , 
    R_13ea_1580dc58 , 
    R_dcb_1162f798 , 
    R_7ac_13c08838 , 
    R_ab1_150e1b78 , 
    R_10d0_150e7938 , 
    R_16ef_14a136f8 , 
    R_a6c_123b7378 , 
    R_142f_117f79d8 , 
    R_108b_156b83d8 , 
    R_e10_14a0b4f8 , 
    R_16aa_150e47d8 , 
    R_7f1_123bc378 , 
    R_1a4e_123b60b8 , 
    R_5b2_1486f018 , 
    R_cab_15fee028 , 
    R_bd1_1587dfb8 , 
    R_68c_123c1b98 , 
    R_11f0_13cd3a18 , 
    R_18e9_13b98a18 , 
    R_180f_13c1cbf8 , 
    R_12ca_14a13dd8 , 
    R_1000_13d4e858 , 
    R_e9b_13cd5f98 , 
    R_9e1_13bea878 , 
    R_161f_10080098 , 
    R_14ba_1580ba98 , 
    R_87c_13dee6d8 , 
    R_830_1008cc58 , 
    R_a2d_13d43f38 , 
    R_146e_17010ba8 , 
    R_104c_13d1f658 , 
    R_e4f_13ccef18 , 
    R_166b_116345b8 , 
    R_ff7_13c0cf78 , 
    R_ea4_117ea738 , 
    R_9d8_156b6ad8 , 
    R_1616_17009da8 , 
    R_14c3_116384d8 , 
    R_885_13de02f8 , 
    R_11b7_11c6de38 , 
    R_1922_13c26018 , 
    R_579_13d5d358 , 
    R_6c5_13d59398 , 
    R_17d6_11c6d258 , 
    R_1303_156b3d38 , 
    R_b98_14b1aeb8 , 
    R_ce4_117f17b8 , 
    R_96b_15816c18 , 
    R_8f2_158891d8 , 
    R_f11_124c3598 , 
    R_15a9_1007e0b8 , 
    R_1530_13c1c5b8 , 
    R_f8a_1580da78 , 
    R_5ab_13d20b98 , 
    R_cb2_15883eb8 , 
    R_bca_1162ecf8 , 
    R_693_1580e978 , 
    R_18f0_14868178 , 
    R_11e9_12fc0518 , 
    R_12d1_15ff4388 , 
    R_1808_117ec998 , 
    R_112e_124c40d8 , 
    R_d6d_10080278 , 
    R_b0f_150e1e98 , 
    R_138c_14a12938 , 
    R_19ab_1486d5d8 , 
    R_174d_13c05318 , 
    R_74e_117e9dd8 , 
    R_5d4_1587e918 , 
    R_18c7_117ed7f8 , 
    R_bf3_158826f8 , 
    R_12a8_140b92d8 , 
    R_1212_13debed8 , 
    R_c89_15886078 , 
    R_1831_13b99eb8 , 
    R_66a_117f7c58 , 
    R_16fb_13d39a38 , 
    R_10dc_140acad8 , 
    R_abd_12fbf938 , 
    R_7a0_1162cef8 , 
    R_dbf_13d1dd58 , 
    R_13de_13bf51d8 , 
    R_19fd_13c22cd8 , 
    R_a62_11630378 , 
    R_e1a_13d29f18 , 
    R_1081_156ae298 , 
    R_7fb_13c27c38 , 
    R_16a0_1007f9b8 , 
    R_1a58_123b6a18 , 
    R_1439_11637c18 , 
    R_1511_1162c778 , 
    R_15c8_10085a98 , 
    R_8d3_15fefba8 , 
    R_fa9_150dc218 , 
    R_ef2_13d3af78 , 
    R_98a_11629578 , 
    R_151a_15ff8d48 , 
    R_15bf_15ff4f68 , 
    R_8dc_13dd7b58 , 
    R_fa0_1162a838 , 
    R_efb_13ccc2b8 , 
    R_981_156acad8 , 
    R_133f_11636ef8 , 
    R_179a_13ccf918 , 
    R_701_13dd6438 , 
    R_195e_15817578 , 
    R_117b_156b5f98 , 
    R_d20_1162aa18 , 
    R_b5c_116370d8 , 
    R_c0c_13d3f7f8 , 
    R_122b_117ec498 , 
    R_18ae_13d39998 , 
    R_184a_124c54d8 , 
    R_128f_123b97b8 , 
    R_c70_15885998 , 
    R_651_14a122f8 , 
    R_5ed_13cccad8 , 
    R_1a0b_1486ee38 , 
    R_13ec_117f2758 , 
    R_dcd_13d1e438 , 
    R_7ae_13d3c058 , 
    R_aaf_140af698 , 
    R_10ce_11637538 , 
    R_16ed_156af558 , 
    R_a55_12fbef38 , 
    R_e27_13d405b8 , 
    R_1074_14b1a878 , 
    R_808_13c22c38 , 
    R_1693_13cd4558 , 
    R_1a65_1587f8b8 , 
    R_1446_1587eff8 , 
    R_a3c_150e6038 , 
    R_821_117f1b78 , 
    R_105b_13cd2f78 , 
    R_145f_13b8d398 , 
    R_167a_13df45d8 , 
    R_e40_13c26f18 , 
    R_1584_1580b318 , 
    R_f65_13d3b5b8 , 
    R_946_14a10a98 , 
    R_917_117f5458 , 
    R_f36_14a118f8 , 
    R_1555_15815638 , 
    R_cd0_117f6d58 , 
    R_58d_1587f3b8 , 
    R_17ea_15ffadc8 , 
    R_190e_13bf3d38 , 
    R_6b1_15ffc808 , 
    R_bac_13c0a098 , 
    R_12ef_14b277f8 , 
    R_11cb_15ff6f48 , 
    R_977_1580b1d8 , 
    R_8e6_1580c0d8 , 
    R_15b5_14866f58 , 
    R_f05_123b8ef8 , 
    R_f96_15885538 , 
    R_1524_1162d178 , 
    R_11a5_156b5138 , 
    R_567_13bf17b8 , 
    R_6d7_12fc12d8 , 
    R_1315_123b2698 , 
    R_17c4_13ccc718 , 
    R_b86_123b9a38 , 
    R_cf6_14b29738 , 
    R_1934_123bf7f8 , 
    R_1338_116375d8 , 
    R_6fa_13bec218 , 
    R_1182_13c1c658 , 
    R_1957_13d3ec18 , 
    R_d19_13def3f8 , 
    R_b63_15ffbb88 , 
    R_17a1_117f24d8 , 
    R_132d_1587ce38 , 
    R_6ef_158893b8 , 
    R_118d_124c3958 , 
    R_194c_1587cbb8 , 
    R_d0e_13c10998 , 
    R_b6e_117ef5f8 , 
    R_17ac_1486cb38 , 
    R_12b2_156ab458 , 
    R_be9_14867638 , 
    R_c93_14a12258 , 
    R_1208_13bec358 , 
    R_674_123c0018 , 
    R_1827_13c01b78 , 
    R_18d1_117e98d8 , 
    R_5ca_13ccca38 , 
    R_16fd_13bf4378 , 
    R_10de_140b68f8 , 
    R_abf_13befd78 , 
    R_79e_15817b18 , 
    R_dbd_117f2b18 , 
    R_13dc_13d1ce58 , 
    R_19fb_150e3978 , 
    R_858_150dae18 , 
    R_1496_13b8b098 , 
    R_1643_1162c278 , 
    R_a05_117f4cd8 , 
    R_e77_1486b878 , 
    R_1024_11635058 , 
    R_733_10086998 , 
    R_b2a_150dd2f8 , 
    R_d52_1580c498 , 
    R_1768_15813b58 , 
    R_1371_156b10d8 , 
    R_1149_156aff58 , 
    R_1990_117f1df8 , 
    R_185d_1162a0b8 , 
    R_189b_123bccd8 , 
    R_127c_1580f198 , 
    R_c5d_13bf88d8 , 
    R_63e_170163c8 , 
    R_600_150e8798 , 
    R_c1f_117ebdb8 , 
    R_123e_13ccb318 , 
    R_bfe_17018b28 , 
    R_18bc_123b9df8 , 
    R_121d_11632718 , 
    R_129d_117f6998 , 
    R_183c_14b21498 , 
    R_c7e_14a0d6b8 , 
    R_65f_14874978 , 
    R_5df_13c24178 , 
    R_833_117f3dd8 , 
    R_a2a_14869bb8 , 
    R_1471_140adbb8 , 
    R_1049_11636138 , 
    R_e52_13d4e498 , 
    R_1668_13b909f8 , 
    R_15df_14b24c38 , 
    R_14fa_15ff7128 , 
    R_fc0_13beba98 , 
    R_8bc_14a0e338 , 
    R_9a1_123b5758 , 
    R_edb_17017048 , 
    R_1a0d_13ccaaf8 , 
    R_13ee_13d23398 , 
    R_dcf_13cccfd8 , 
    R_7b0_123bf4d8 , 
    R_aad_14873a78 , 
    R_10cc_13cd01d8 , 
    R_16eb_150e81f8 , 
    R_172d_13cda318 , 
    R_13ac_116343d8 , 
    R_110e_14a11998 , 
    R_19cb_13d3a758 , 
    R_aef_13d50dd8 , 
    R_76e_13bf8d38 , 
    R_d8d_13dd52b8 , 
    R_715_13b94ff8 , 
    R_1972_156aa918 , 
    R_1786_140b5778 , 
    R_d34_15ff3b68 , 
    R_1167_1587c7f8 , 
    R_1353_123c05b8 , 
    R_b48_15814378 , 
    R_17fb_11c6bd18 , 
    R_59e_13cd0098 , 
    R_cbf_15fed948 , 
    R_bbd_13b8f418 , 
    R_18fd_15882798 , 
    R_6a0_117edbb8 , 
    R_11dc_150db458 , 
    R_12de_117e9658 , 
    R_19db_123b8458 , 
    R_171d_13d45e78 , 
    R_10fe_117ebd18 , 
    R_adf_13ccfcd8 , 
    R_77e_123bcff8 , 
    R_d9d_12fc0298 , 
    R_13bc_13c07cf8 , 
    R_142a_14a0f2d8 , 
    R_1090_1486e7f8 , 
    R_e0b_156b7758 , 
    R_16af_1486be18 , 
    R_7ec_123b4038 , 
    R_1a49_13ccbb38 , 
    R_a71_117f59f8 , 
    R_15f2_13d4fe38 , 
    R_ec8_15883058 , 
    R_fd3_10088798 , 
    R_14e7_14b1ce98 , 
    R_9b4_13bf5b38 , 
    R_8a9_13c21298 , 
    R_ece_11634bf8 , 
    R_15ec_13d3f4d8 , 
    R_14ed_117f5f98 , 
    R_fcd_1580d258 , 
    R_8af_13ddfb78 , 
    R_9ae_140b18f8 , 
    R_1501_117f0a98 , 
    R_15d8_11c6ea18 , 
    R_fb9_15ff0be8 , 
    R_8c3_10081498 , 
    R_99a_15ffaaa8 , 
    R_ee2_13cd1b78 , 
    R_1712_11637178 , 
    R_10f3_14a19238 , 
    R_ad4_14a0a5f8 , 
    R_789_140b2cf8 , 
    R_da8_140b3838 , 
    R_13c7_13df0ed8 , 
    R_19e6_11636958 , 
    R_95d_117f8338 , 
    R_900_140b74d8 , 
    R_f1f_1587f1d8 , 
    R_153e_13d410f8 , 
    R_159b_1162f658 , 
    R_f7c_15ffc268 , 
    R_cc5_13b8c858 , 
    R_598_17015108 , 
    R_17f5_13c1c798 , 
    R_1903_1162d2b8 , 
    R_6a6_15816df8 , 
    R_bb7_14a17a78 , 
    R_12e4_13df4678 , 
    R_11d6_13cccf38 , 
    R_a4d_14a159f8 , 
    R_810_1007f918 , 
    R_106c_13cd4238 , 
    R_168b_13d20d78 , 
    R_144e_17019028 , 
    R_e2f_123b83b8 , 
    R_f66_1700e448 , 
    R_947_13cd36f8 , 
    R_916_12fbefd8 , 
    R_f35_13dd5fd8 , 
    R_1554_13c04918 , 
    R_1585_117efe18 , 
    R_16ff_13b95318 , 
    R_10e0_1580e478 , 
    R_ac1_13d23078 , 
    R_79c_1162d8f8 , 
    R_dbb_1580e018 , 
    R_13da_123c03d8 , 
    R_19f9_13cd81f8 , 
    R_a3f_13c012b8 , 
    R_81e_140b4cd8 , 
    R_105e_156ba278 , 
    R_145c_13ddc0b8 , 
    R_167d_124c5438 , 
    R_e3d_15889778 , 
    R_be0_117ea5f8 , 
    R_c9c_13b8ed38 , 
    R_11ff_14a17618 , 
    R_67d_156b7398 , 
    R_181e_13c04e18 , 
    R_18da_13cd38d8 , 
    R_5c1_13c0a818 , 
    R_12bb_13b8a918 , 
    R_ca4_156b1c18 , 
    R_bd8_117e87f8 , 
    R_685_13bf38d8 , 
    R_11f7_10080b38 , 
    R_18e2_13becfd8 , 
    R_1816_14b1ff58 , 
    R_12c3_10083478 , 
    R_5b9_140b2bb8 , 
    R_1630_123b9cb8 , 
    R_e8a_14b1db18 , 
    R_9f2_10089418 , 
    R_14a9_156acb78 , 
    R_1011_12fbe218 , 
    R_86b_124c4e98 , 
    R_1726_14869a78 , 
    R_19d2_13d533f8 , 
    R_1107_13df9038 , 
    R_ae8_13bef5f8 , 
    R_775_158109f8 , 
    R_d94_12fbf6b8 , 
    R_13b3_13d40158 , 
    R_1658_13bf9ff8 , 
    R_843_150e0458 , 
    R_1481_117e8e38 , 
    R_a1a_15fefd88 , 
    R_1039_13ddba78 , 
    R_e62_13c23098 , 
    R_1a0f_13c24038 , 
    R_13f0_11c6e338 , 
    R_dd1_13de4a38 , 
    R_7b2_13bf2898 , 
    R_aab_13c1cfb8 , 
    R_10ca_1700ac08 , 
    R_16e9_15ff3668 , 
    R_1793_150de018 , 
    R_708_14a0d258 , 
    R_1965_13ccb6d8 , 
    R_1174_11c6c358 , 
    R_d27_13dee138 , 
    R_b55_15ffb0e8 , 
    R_1346_13d3f2f8 , 
    R_e1f_123b6ab8 , 
    R_107c_117f4058 , 
    R_800_13d219f8 , 
    R_169b_150e49b8 , 
    R_1a5d_1486e398 , 
    R_143e_14a19f58 , 
    R_a5d_15880498 , 
    R_1a22_15810b38 , 
    R_1403_124c5398 , 
    R_de4_117f6498 , 
    R_7c5_15ffbe08 , 
    R_a98_1486db78 , 
    R_10b7_14a17578 , 
    R_16d6_14a10458 , 
    R_1a2d_13b8fcd8 , 
    R_140e_13def718 , 
    R_def_13d3eb78 , 
    R_7d0_156b2e38 , 
    R_a8d_11632678 , 
    R_10ac_156b5958 , 
    R_16cb_156b72f8 , 
    R_1634_17018c68 , 
    R_9f6_158867f8 , 
    R_e86_14a183d8 , 
    R_1015_14b1e6f8 , 
    R_867_15881398 , 
    R_14a5_11629ed8 , 
    R_e8e_150da878 , 
    R_9ee_13d54618 , 
    R_162c_13b96c18 , 
    R_14ad_12fbf618 , 
    R_86f_15ff83e8 , 
    R_100d_158136f8 , 
    R_189c_14a10c78 , 
    R_127d_11636318 , 
    R_c5e_15882a18 , 
    R_63f_156b5b38 , 
    R_5ff_13d40ab8 , 
    R_c1e_14a0b958 , 
    R_123d_13ddd5f8 , 
    R_185c_11630738 , 
    R_141e_13b90818 , 
    R_16bb_123b7d78 , 
    R_dff_117eeb58 , 
    R_7e0_13dfacf8 , 
    R_a7d_123b7af8 , 
    R_1a3d_156b9cd8 , 
    R_109c_13b98d38 , 
    R_cb9_150db638 , 
    R_bc3_156b6678 , 
    R_69a_13b8b6d8 , 
    R_18f7_13b90bd8 , 
    R_11e2_13d1e4d8 , 
    R_12d8_13d43718 , 
    R_1801_13c013f8 , 
    R_5a4_15ff7d08 , 
    R_13a5_13d45338 , 
    R_1115_11630b98 , 
    R_19c4_17016fa8 , 
    R_af6_117f49b8 , 
    R_767_117f2d98 , 
    R_d86_15fef7e8 , 
    R_1734_1580c718 , 
    R_836_123b33b8 , 
    R_a27_117ede38 , 
    R_1474_13c042d8 , 
    R_1046_123bc918 , 
    R_e55_124c3a98 , 
    R_1665_156ac678 , 
    R_122a_14a0b318 , 
    R_18af_11c6f7d8 , 
    R_1849_140b6358 , 
    R_1290_13dd8b98 , 
    R_c71_14a11e98 , 
    R_652_13d386d8 , 
    R_5ec_14868df8 , 
    R_c0b_13b8c038 , 
    R_574_13d4ec18 , 
    R_6ca_156b3f18 , 
    R_1308_117f2438 , 
    R_17d1_11c6fa58 , 
    R_b93_15881078 , 
    R_ce9_156b86f8 , 
    R_1927_123bb6f8 , 
    R_11b2_14a101d8 , 
    R_8f1_14a0fcd8 , 
    R_f10_156ab778 , 
    R_15aa_13c1f498 , 
    R_152f_158884b8 , 
    R_f8b_13dda218 , 
    R_96c_15ff4e28 , 
    R_948_15ff1728 , 
    R_915_158834b8 , 
    R_f34_123bd958 , 
    R_1553_1162fdd8 , 
    R_1586_13cd7938 , 
    R_f67_156b54f8 , 
    R_1701_117ee5b8 , 
    R_10e2_13b97cf8 , 
    R_ac3_13d41ff8 , 
    R_79a_13b8d758 , 
    R_db9_13d4e358 , 
    R_13d8_13c10178 , 
    R_19f7_123b4218 , 
    R_ec2_156acdf8 , 
    R_fd9_13cd6038 , 
    R_14e1_13d4fbb8 , 
    R_9ba_13d3b018 , 
    R_8a3_117f3298 , 
    R_15f8_150dd618 , 
    R_b1c_10084238 , 
    R_d60_1700c1e8 , 
    R_137f_13d27fd8 , 
    R_175a_15fedda8 , 
    R_199e_123b8d18 , 
    R_113b_11c703b8 , 
    R_741_156b0278 , 
    R_15e6_140b4238 , 
    R_14f3_10088a18 , 
    R_fc7_117e8c58 , 
    R_8b5_13ccefb8 , 
    R_9a8_14a19af8 , 
    R_ed4_150e1998 , 
    R_d68_15885b78 , 
    R_b14_11c6b8b8 , 
    R_1387_117eaf58 , 
    R_19a6_14a19738 , 
    R_1752_150e4738 , 
    R_749_123b2918 , 
    R_1133_1587e378 , 
    R_1417_15ff4428 , 
    R_df8_15888eb8 , 
    R_7d9_124c3098 , 
    R_a84_13b8b778 , 
    R_10a3_13c1e4f8 , 
    R_1a36_14b1b318 , 
    R_16c2_156b1e98 , 
    R_1a11_123b7b98 , 
    R_13f2_13de2738 , 
    R_dd3_14a19a58 , 
    R_7b4_15885a38 , 
    R_aa9_13cd5818 , 
    R_10c8_14a14058 , 
    R_16e7_117eea18 , 
    R_b27_10087e38 , 
    R_d55_117f0f98 , 
    R_1765_12fbdf98 , 
    R_1374_17015888 , 
    R_1146_123bed58 , 
    R_1993_13d53b78 , 
    R_736_15ff9108 , 
    R_56b_123b7558 , 
    R_6d3_1007e1f8 , 
    R_1311_10087a78 , 
    R_17c8_13d50a18 , 
    R_b8a_14b26858 , 
    R_cf2_14a17438 , 
    R_1930_13c083d8 , 
    R_11a9_117f1038 , 
    R_1638_15815818 , 
    R_9fa_123b77d8 , 
    R_e82_13df3ef8 , 
    R_1019_158858f8 , 
    R_863_13d47318 , 
    R_14a1_117ed938 , 
    R_eb2_11c6d2f8 , 
    R_fe9_1162ed98 , 
    R_14d1_1587ae58 , 
    R_9ca_1587bd58 , 
    R_893_13ccf238 , 
    R_1608_117f45f8 , 
    R_6f3_17012cc8 , 
    R_1189_13de2d78 , 
    R_1950_123b8098 , 
    R_d12_13cd6d58 , 
    R_b6a_140afff8 , 
    R_17a8_13d3cf58 , 
    R_1331_148755f8 , 
    R_e9f_17016288 , 
    R_9dd_156ab8b8 , 
    R_161b_13d3ca58 , 
    R_14be_13b98478 , 
    R_880_117ea2d8 , 
    R_ffc_13b8acd8 , 
    R_1789_13cca9b8 , 
    R_196f_13bf01d8 , 
    R_d31_156b13f8 , 
    R_116a_13c23e58 , 
    R_1350_11632498 , 
    R_b4b_156ad398 , 
    R_712_13b90d18 , 
    R_e92_117f2ed8 , 
    R_9ea_123b7e18 , 
    R_1628_123b7698 , 
    R_14b1_14a16e98 , 
    R_873_14a14238 , 
    R_1009_13b980b8 , 
    R_bf2_170099e8 , 
    R_12a9_1162d0d8 , 
    R_1211_150e5278 , 
    R_c8a_150e3798 , 
    R_1830_13bf6358 , 
    R_66b_150e1498 , 
    R_5d3_158808f8 , 
    R_18c8_13cd9f58 , 
    R_a42_15888198 , 
    R_81b_12fbec18 , 
    R_1061_13d3c558 , 
    R_1459_17016aa8 , 
    R_1680_1486aab8 , 
    R_e3a_123bb798 , 
    R_17ef_15889958 , 
    R_1909_15815e58 , 
    R_6ac_12fc1918 , 
    R_bb1_14874d38 , 
    R_12ea_13ddf358 , 
    R_11d0_170096c8 , 
    R_ccb_117ec038 , 
    R_592_13c23958 , 
    R_fee_14b29f58 , 
    R_ead_13c22378 , 
    R_9cf_1162e118 , 
    R_14cc_123c0b58 , 
    R_160d_123bff78 , 
    R_88e_123c0fb8 , 
    R_8ff_156b7c58 , 
    R_f1e_15880038 , 
    R_153d_15811218 , 
    R_159c_15815db8 , 
    R_f7d_13cd0778 , 
    R_95e_13b98018 , 
    R_189d_13cd3518 , 
    R_127e_13d4f118 , 
    R_c5f_12fbfa78 , 
    R_640_140b2258 , 
    R_5fe_15888558 , 
    R_c1d_13dfb1f8 , 
    R_123c_15fee708 , 
    R_185b_14b21538 , 
    R_15d1_123b63d8 , 
    R_fb2_15810818 , 
    R_8ca_15815bd8 , 
    R_993_11c6b598 , 
    R_ee9_1700fca8 , 
    R_1508_156b7898 , 
    R_121c_158871f8 , 
    R_129e_13d3cb98 , 
    R_183b_13c20bb8 , 
    R_c7f_13cd6ad8 , 
    R_660_156ba458 , 
    R_5de_123b7cd8 , 
    R_18bd_140b9878 , 
    R_bfd_11c6f238 , 
    R_16b4_117ead78 , 
    R_e06_1580ff58 , 
    R_7e7_15885858 , 
    R_1a44_1162c4f8 , 
    R_a76_13d38638 , 
    R_1095_156b0ef8 , 
    R_1425_13d571d8 , 
    R_8e5_150db318 , 
    R_15b6_1580e838 , 
    R_f04_15885038 , 
    R_f97_1700c288 , 
    R_1523_140b8e78 , 
    R_978_156b6498 , 
    R_914_13d54c58 , 
    R_f33_13d59258 , 
    R_1552_13ccfa58 , 
    R_1587_140aacd8 , 
    R_f68_140acb78 , 
    R_949_14b26a38 , 
    R_15c0_158147d8 , 
    R_8db_1580e158 , 
    R_fa1_1162ffb8 , 
    R_efa_13bf5818 , 
    R_982_13debcf8 , 
    R_1519_15813e78 , 
    R_164e_117eb138 , 
    R_148b_15886118 , 
    R_a10_13df0f78 , 
    R_e6c_15ff0d28 , 
    R_102f_123c08d8 , 
    R_84d_15feee88 , 
    R_1703_13c254d8 , 
    R_10e4_158894f8 , 
    R_ac5_15883558 , 
    R_798_123beb78 , 
    R_db7_14869938 , 
    R_13d6_156ae8d8 , 
    R_19f5_13d2c2b8 , 
    R_eb7_11c6d1b8 , 
    R_fe4_12fc21d8 , 
    R_14d6_1008b178 , 
    R_9c5_14b21d58 , 
    R_898_123b5c58 , 
    R_1603_14872fd8 , 
    R_1714_15889638 , 
    R_10f5_140b5f98 , 
    R_ad6_14873258 , 
    R_787_14a0e838 , 
    R_da6_13ddc158 , 
    R_13c5_15fee208 , 
    R_19e4_13de3a98 , 
    R_98b_13b8dcf8 , 
    R_ef1_13b924d8 , 
    R_8d2_156ad578 , 
    R_faa_156b0458 , 
    R_1510_13d1f0b8 , 
    R_15c9_13bf0b38 , 
    R_aa7_13d451f8 , 
    R_7b6_14a18018 , 
    R_dd5_124c5258 , 
    R_10c6_1700ff28 , 
    R_13f4_14a0b778 , 
    R_16e5_13c07ed8 , 
    R_1a13_117ef058 , 
    R_839_14b28f18 , 
    R_e58_158814d8 , 
    R_a24_123b5938 , 
    R_1043_14b26538 , 
    R_1477_117f0098 , 
    R_1662_13df1978 , 
    R_854_15ff3e88 , 
    R_e73_14b288d8 , 
    R_a09_123bb158 , 
    R_1028_117f4eb8 , 
    R_1492_13cd4378 , 
    R_1647_12fc19b8 , 
    R_be8_15ffcee8 , 
    R_5c9_14b27438 , 
    R_675_156aec98 , 
    R_c94_13b8fb98 , 
    R_1207_156b81f8 , 
    R_12b3_13ddf718 , 
    R_1826_140b01d8 , 
    R_18d2_13c290d8 , 
    R_cac_123c1058 , 
    R_5b1_13d28e38 , 
    R_68d_1700f2a8 , 
    R_bd0_13ccc538 , 
    R_11ef_117f3d38 , 
    R_12cb_123bfe38 , 
    R_180e_1580c7b8 , 
    R_18ea_14a115d8 , 
    R_d75_1486bc38 , 
    R_756_13b8ae18 , 
    R_b07_140aaa58 , 
    R_1126_156aaeb8 , 
    R_1394_15814878 , 
    R_1745_123b4cb8 , 
    R_19b3_123bc558 , 
    R_d7a_13b95ef8 , 
    R_75b_15814558 , 
    R_b02_14a13f18 , 
    R_1121_150e9c38 , 
    R_1399_158830f8 , 
    R_1740_13cd6fd8 , 
    R_19b8_15812c58 , 
    R_c0a_14a19ff8 , 
    R_5eb_15feeac8 , 
    R_653_123be358 , 
    R_c72_13df6fb8 , 
    R_1229_156b7938 , 
    R_1291_14a0d758 , 
    R_1848_14a197d8 , 
    R_18b0_15815a98 , 
    R_a96_150e8478 , 
    R_7c7_13d45c98 , 
    R_de6_13c05778 , 
    R_10b5_156ab6d8 , 
    R_1405_14a192d8 , 
    R_16d4_14868c18 , 
    R_1a24_116348d8 , 
    R_85f_13dd89b8 , 
    R_e7e_140ad6b8 , 
    R_9fe_13c02d98 , 
    R_101d_123b5d98 , 
    R_149d_156b8dd8 , 
    R_163c_1486a6f8 , 
    R_d9b_13d3dbd8 , 
    R_77c_116359b8 , 
    R_ae1_15fed768 , 
    R_1100_10085818 , 
    R_13ba_15881d98 , 
    R_171f_13bf08b8 , 
    R_19d9_1700c508 , 
    R_889_15ff9b08 , 
    R_9d4_11c6e6f8 , 
    R_ea8_13d1fe78 , 
    R_ff3_117efc38 , 
    R_14c7_140b4918 , 
    R_1612_13cd0278 , 
    R_582_14869118 , 
    R_cdb_14a0ae18 , 
    R_ba1_13d29338 , 
    R_6bc_13cd53b8 , 
    R_11c0_13deef98 , 
    R_12fa_11631638 , 
    R_17df_13cd0e58 , 
    R_1919_1587e2d8 , 
    R_e24_13ddcfb8 , 
    R_a58_14a18a18 , 
    R_805_1580a7d8 , 
    R_1077_11c6d898 , 
    R_1443_13d3f9d8 , 
    R_1696_156afd78 , 
    R_1a62_14b1b138 , 
    R_94a_156b24d8 , 
    R_f32_116350f8 , 
    R_913_100840f8 , 
    R_f69_117f0c78 , 
    R_1551_150dde38 , 
    R_1588_150e7d98 , 
    R_a50_13df7698 , 
    R_e2c_15881e38 , 
    R_80d_14a16a38 , 
    R_106f_156ad938 , 
    R_144b_1486ce58 , 
    R_168e_123bbc98 , 
    R_6fe_13bf5318 , 
    R_b5f_13cd4918 , 
    R_d1d_13def2b8 , 
    R_117e_14a0ccb8 , 
    R_133c_117f2938 , 
    R_179d_10085138 , 
    R_195b_14b1c8f8 , 
    R_cb3_1587b358 , 
    R_5aa_13dd5678 , 
    R_694_11636b38 , 
    R_bc9_124c3d18 , 
    R_11e8_13ccd258 , 
    R_12d2_123bdc78 , 
    R_1807_117ee298 , 
    R_18f1_156aba98 , 
    R_c1c_156ba3b8 , 
    R_5fd_14a10958 , 
    R_641_123b90d8 , 
    R_c60_158171b8 , 
    R_123b_1162cd18 , 
    R_127f_13b8a558 , 
    R_185a_15814cd8 , 
    R_189e_13bf8e78 , 
    R_877_13d3e498 , 
    R_9e6_14b28838 , 
    R_e96_156b4a58 , 
    R_1005_13c1edb8 , 
    R_14b5_15882018 , 
    R_1624_10086cb8 , 
    R_db5_117ece98 , 
    R_796_156b0138 , 
    R_ac7_148725d8 , 
    R_10e6_11630918 , 
    R_13d4_15882bf8 , 
    R_1705_10085db8 , 
    R_19f3_1008c618 , 
    R_96d_1162e7f8 , 
    R_f0f_13d3d9f8 , 
    R_8f0_13d29838 , 
    R_f8c_117f2578 , 
    R_152e_117f3f18 , 
    R_15ab_13ccc358 , 
    R_587_124c5118 , 
    R_cd6_13d39178 , 
    R_ba6_156ad9d8 , 
    R_6b7_13c0b718 , 
    R_11c5_13d39538 , 
    R_12f5_158104f8 , 
    R_17e4_156acf38 , 
    R_1914_10084f58 , 
    R_846_100885b8 , 
    R_e65_15810318 , 
    R_a17_13ccf878 , 
    R_1036_140b5278 , 
    R_1484_11c6b778 , 
    R_1655_1700cdc8 , 
    R_a45_17017188 , 
    R_e37_10083018 , 
    R_818_13b8dbb8 , 
    R_1064_1700d5e8 , 
    R_1456_13cd8518 , 
    R_1683_1587f6d8 , 
    R_57d_14b1ef18 , 
    R_ce0_1580ccb8 , 
    R_b9c_15884e58 , 
    R_6c1_156b1538 , 
    R_11bb_117ed2f8 , 
    R_12ff_17012408 , 
    R_17da_123bf398 , 
    R_191e_140b0c78 , 
    R_d58_13df39f8 , 
    R_b24_15815958 , 
    R_739_123c1698 , 
    R_1143_13cd7078 , 
    R_1377_158873d8 , 
    R_1762_140aef18 , 
    R_1996_156b4058 , 
    R_95f_13bf9918 , 
    R_f1d_15ff80c8 , 
    R_8fe_13d4f898 , 
    R_f7e_156b42d8 , 
    R_153c_13c1d698 , 
    R_159d_1162b198 , 
    R_aa5_156b4238 , 
    R_7b8_1162e9d8 , 
    R_dd7_140b62b8 , 
    R_10c4_12fc1878 , 
    R_13f6_1700d728 , 
    R_16e3_123b4d58 , 
    R_1a15_13d3e998 , 
    R_b0c_123c1878 , 
    R_d70_13b96038 , 
    R_751_13bf12b8 , 
    R_112b_13d5c3b8 , 
    R_138f_13df66f8 , 
    R_174a_13d24658 , 
    R_19ae_1587f818 , 
    R_a8b_117f7898 , 
    R_7d2_10082a78 , 
    R_df1_15884778 , 
    R_10aa_13c28458 , 
    R_1410_13cd5a98 , 
    R_16c9_13c03018 , 
    R_1a2f_15886b18 , 
    R_d7f_117f5ef8 , 
    R_760_13cce6f8 , 
    R_afd_156ae018 , 
    R_111c_13c0f138 , 
    R_139e_15ff9428 , 
    R_173b_13d23758 , 
    R_19bd_150e0c78 , 
    R_70f_14b26038 , 
    R_b4e_158835f8 , 
    R_d2e_15ff2d08 , 
    R_116d_14a0bc78 , 
    R_134d_13cd26b8 , 
    R_178c_13d39718 , 
    R_196c_117ef418 , 
    R_705_17018768 , 
    R_b58_12fc00b8 , 
    R_d24_13c0ca78 , 
    R_1177_13d5b558 , 
    R_1343_13d298d8 , 
    R_1796_156ae338 , 
    R_1962_13d5d218 , 
    R_c9d_13c00ef8 , 
    R_bdf_117f0638 , 
    R_5c0_117ea0f8 , 
    R_67e_14a0b8b8 , 
    R_11fe_124c36d8 , 
    R_12bc_13b981f8 , 
    R_181d_123ba758 , 
    R_18db_11c6d7f8 , 
    R_ebc_1580cfd8 , 
    R_89d_11c693d8 , 
    R_9c0_13d46b98 , 
    R_fdf_158176b8 , 
    R_14db_156b5e58 , 
    R_15fe_140b97d8 , 
    R_ee1_13d40c98 , 
    R_99b_156b3838 , 
    R_8c2_15813518 , 
    R_fba_140aebf8 , 
    R_1500_1700e8a8 , 
    R_15d9_13d53538 , 
    R_eda_13d57638 , 
    R_9a2_13c28bd8 , 
    R_8bb_13d43498 , 
    R_fc1_156b40f8 , 
    R_14f9_13cd6178 , 
    R_15e0_13cd0458 , 
    R_d8b_150dc7b8 , 
    R_76c_150e63f8 , 
    R_af1_13b8c3f8 , 
    R_1110_13d5cdb8 , 
    R_13aa_14b1d898 , 
    R_172f_11c6dbb8 , 
    R_19c9_1509b4f8 , 
    R_55a_158145f8 , 
    R_6e4_11630a58 , 
    R_b79_13ccfd78 , 
    R_d03_124c2eb8 , 
    R_1198_117f3b58 , 
    R_1322_15ff6ea8 , 
    R_17b7_15810bd8 , 
    R_1941_117ed4d8 , 
    R_6cf_1486c6d8 , 
    R_56f_14a0b598 , 
    R_cee_13cd9c38 , 
    R_b8e_150e97d8 , 
    R_11ad_13d569b8 , 
    R_130d_124c3818 , 
    R_17cc_117e9298 , 
    R_192c_13b94918 , 
    R_94b_100881f8 , 
    R_f31_13c231d8 , 
    R_912_11630f58 , 
    R_f6a_117ea058 , 
    R_1550_17014668 , 
    R_1589_123b7198 , 
    R_bd7_14a0ef18 , 
    R_ca5_1007eb58 , 
    R_5b8_170170e8 , 
    R_686_15810f98 , 
    R_11f6_14b22bb8 , 
    R_12c4_15ff0008 , 
    R_1815_156b1cb8 , 
    R_18e3_13ccb9f8 , 
    R_6e0_14a15f98 , 
    R_55e_148707d8 , 
    R_cff_14a0b458 , 
    R_b7d_156b6df8 , 
    R_119c_14872ad8 , 
    R_131e_13dd6e38 , 
    R_17bb_13bf1d58 , 
    R_193d_11c70638 , 
    R_d92_14b21358 , 
    R_773_117f54f8 , 
    R_aea_17012908 , 
    R_1109_15ff3de8 , 
    R_13b1_150dc358 , 
    R_1728_13d5beb8 , 
    R_19d0_14870af8 , 
    R_e12_13b8cc18 , 
    R_a6a_13d1d218 , 
    R_7f3_148688f8 , 
    R_1089_123b6838 , 
    R_1431_15812ed8 , 
    R_16a8_123bf118 , 
    R_1a50_117ed6b8 , 
    R_6f7_117e93d8 , 
    R_b66_14a0f238 , 
    R_d16_13c1b7f8 , 
    R_1185_13d1ecf8 , 
    R_1335_13bf1f38 , 
    R_17a4_14b1ea18 , 
    R_1954_15ff1ae8 , 
    R_e17_13df86d8 , 
    R_a65_14b22b18 , 
    R_7f8_1700bec8 , 
    R_1084_13d39038 , 
    R_1436_15fef608 , 
    R_16a3_15ff2768 , 
    R_1a55_123b5898 , 
    R_a21_1587bad8 , 
    R_83c_13cd7398 , 
    R_e5b_123bf898 , 
    R_1040_1008ac78 , 
    R_147a_13c04378 , 
    R_165f_13cd97d8 , 
    R_bfc_13d53cb8 , 
    R_5dd_123b45d8 , 
    R_661_13d3c2d8 , 
    R_c80_1008ca78 , 
    R_121b_14b24698 , 
    R_129f_1008b7b8 , 
    R_183a_156acc18 , 
    R_18be_14a0de38 , 
    R_c1b_123b48f8 , 
    R_5fc_140b3518 , 
    R_642_14a0d118 , 
    R_c61_13c06718 , 
    R_123a_15ffcf88 , 
    R_1280_14a106d8 , 
    R_1859_13d25378 , 
    R_189f_14a13c98 , 
    R_556_13d2a2d8 , 
    R_6e8_12fbf4d8 , 
    R_b75_156ae838 , 
    R_d07_156abe58 , 
    R_1194_1580f058 , 
    R_1326_11c684d8 , 
    R_17b3_13ddb4d8 , 
    R_1945_14b22898 , 
    R_bf1_13df18d8 , 
    R_5d2_10088f18 , 
    R_66c_123c06f8 , 
    R_c8b_13c0e5f8 , 
    R_1210_117f56d8 , 
    R_12aa_140afb98 , 
    R_182f_13d58998 , 
    R_18c9_11c6eb58 , 
    R_cc0_1580fcd8 , 
    R_59d_13df9d58 , 
    R_6a1_13cd9b98 , 
    R_bbc_13d4e678 , 
    R_11db_124c45d8 , 
    R_12df_13d27178 , 
    R_17fa_13beb8b8 , 
    R_18fe_1587ca78 , 
    R_d63_117f68f8 , 
    R_b19_158882d8 , 
    R_744_123bea38 , 
    R_1138_14869ed8 , 
    R_1382_13b8b958 , 
    R_1757_13de1978 , 
    R_19a1_123b3598 , 
    R_db3_14869898 , 
    R_794_17016788 , 
    R_ac9_15811cb8 , 
    R_10e8_140b1538 , 
    R_13d2_13c292b8 , 
    R_1707_13ddd9b8 , 
    R_19f1_13cce518 , 
    R_ecd_13d5b5f8 , 
    R_9af_1587fdb8 , 
    R_8ae_11631778 , 
    R_fce_13c051d8 , 
    R_14ec_156b01d8 , 
    R_15ed_1008af98 , 
    R_da4_13cd7438 , 
    R_785_116381b8 , 
    R_ad8_117f7a78 , 
    R_10f7_1587f598 , 
    R_13c3_13cd0b38 , 
    R_1716_123b6bf8 , 
    R_19e2_13d567d8 , 
    R_58c_1587fe58 , 
    R_cd1_1486dc18 , 
    R_bab_13df0e38 , 
    R_6b2_14867ef8 , 
    R_11ca_123bd9f8 , 
    R_12f0_158817f8 , 
    R_17e9_123bb5b8 , 
    R_190f_15881b18 , 
    R_979_117efcd8 , 
    R_f03_13c06f38 , 
    R_8e4_123b2b98 , 
    R_f98_13d588f8 , 
    R_1522_15817d98 , 
    R_15b7_11636bd8 , 
    R_c09_14a18bf8 , 
    R_5ea_1162b558 , 
    R_654_150e54f8 , 
    R_c73_15810958 , 
    R_1228_150e4ff8 , 
    R_1292_117e9fb8 , 
    R_1847_13d54898 , 
    R_18b1_1162ae78 , 
    R_ec7_10083838 , 
    R_8a8_140b6858 , 
    R_9b5_156b6038 , 
    R_fd4_13bef878 , 
    R_14e6_123be178 , 
    R_15f3_1580b958 , 
    R_6dc_13d56738 , 
    R_562_11630198 , 
    R_cfb_156b77f8 , 
    R_b81_14b23658 , 
    R_11a0_117f1a38 , 
    R_131a_13cd6678 , 
    R_17bf_1162eed8 , 
    R_1939_13b99198 , 
    R_85b_150e9ff8 , 
    R_e7a_13df06b8 , 
    R_a02_13d20378 , 
    R_1021_14873438 , 
    R_1499_13c056d8 , 
    R_1640_15816e98 , 
    R_6c6_14b27a78 , 
    R_578_13c06678 , 
    R_ce5_117e9518 , 
    R_b97_116328f8 , 
    R_11b6_123b6478 , 
    R_1304_150e5a98 , 
    R_17d5_13cd9eb8 , 
    R_1923_10086ad8 , 
    R_aa3_123ba9d8 , 
    R_7ba_17013308 , 
    R_dd9_1587f4f8 , 
    R_10c2_13de4358 , 
    R_13f8_14866c38 , 
    R_16e1_1587e058 , 
    R_1a17_13d3a398 , 
    R_ea3_117f04f8 , 
    R_884_124c4358 , 
    R_9d9_14a0c178 , 
    R_ff8_14a15098 , 
    R_14c2_13d50e78 , 
    R_1617_13de3e58 , 
    R_e0d_13c081f8 , 
    R_a6f_140ab4f8 , 
    R_7ee_117eb4f8 , 
    R_108e_117ecf38 , 
    R_142c_13d55f18 , 
    R_16ad_15885df8 , 
    R_1a4b_13d3a118 , 
    R_e01_13b8ca38 , 
    R_a7b_150e6f38 , 
    R_7e2_116332f8 , 
    R_109a_140adc58 , 
    R_1420_1580acd8 , 
    R_16b9_13b972f8 , 
    R_1a3f_13cd8f18 , 
    R_597_156aeab8 , 
    R_cc6_1486fd38 , 
    R_bb6_13d58fd8 , 
    R_6a7_140b7938 , 
    R_11d5_14871bd8 , 
    R_12e5_14b28bf8 , 
    R_17f4_156b4cd8 , 
    R_1904_140b9058 , 
    R_dfa_1486ff18 , 
    R_a82_116368b8 , 
    R_7db_150dd1b8 , 
    R_10a1_123b8598 , 
    R_1419_13df1b58 , 
    R_16c0_13b994b8 , 
    R_1a38_13ccab98 , 
    R_911_14b22078 , 
    R_94c_123bc7d8 , 
    R_f30_12fbf898 , 
    R_f6b_13c0a6d8 , 
    R_154f_1700ea88 , 
    R_158a_13c25758 , 
    R_d44_13b99418 , 
    R_b38_13d23618 , 
    R_725_13d4f618 , 
    R_1157_14a13298 , 
    R_1363_124c4718 , 
    R_1776_15882518 , 
    R_1982_15816fd8 , 
    R_983_1700b4c8 , 
    R_ef9_1007e338 , 
    R_8da_1587ba38 , 
    R_fa2_15ffaf08 , 
    R_1518_13c09ff8 , 
    R_15c1_13c1e138 , 
    R_d41_13bf8f18 , 
    R_722_14b26fd8 , 
    R_b3b_14a0f378 , 
    R_115a_156af9b8 , 
    R_1360_156aa5f8 , 
    R_1779_13dec3d8 , 
    R_197f_1700ba68 , 
    R_7fd_13d29658 , 
    R_e1c_156b8158 , 
    R_a60_124c2738 , 
    R_107f_13d55ab8 , 
    R_143b_13cd5458 , 
    R_169e_13d59618 , 
    R_1a5a_117ecd58 , 
    R_a94_158121b8 , 
    R_7c9_13c1bb18 , 
    R_de8_13df22d8 , 
    R_10b3_17011328 , 
    R_1407_140b9cd8 , 
    R_16d2_150e0098 , 
    R_1a26_14868678 , 
    R_e9a_14a0e1f8 , 
    R_87b_123b2e18 , 
    R_9e2_148680d8 , 
    R_1001_100877f8 , 
    R_14b9_150dda78 , 
    R_1620_117efff8 , 
    R_bc2_1580b098 , 
    R_cba_13c20118 , 
    R_5a3_13b98298 , 
    R_69b_13bf94b8 , 
    R_11e1_1486a798 , 
    R_12d9_123ba118 , 
    R_1800_15888378 , 
    R_18f8_156ac538 , 
    R_960_13ccf418 , 
    R_f1c_13df79b8 , 
    R_8fd_123b6fb8 , 
    R_f7f_140aa558 , 
    R_153b_117f5d18 , 
    R_159e_14871db8 , 
    R_d47_13d27998 , 
    R_b35_1587cc58 , 
    R_728_140ba318 , 
    R_1154_117e95b8 , 
    R_1366_17015568 , 
    R_1773_156ac2b8 , 
    R_1985_1162c3b8 , 
    R_b11_15883698 , 
    R_d6b_123b8958 , 
    R_74c_150e17b8 , 
    R_1130_13bef0f8 , 
    R_138a_13d25cd8 , 
    R_174f_13df2058 , 
    R_19a9_1486eed8 , 
    R_6ec_13c03b58 , 
    R_b71_140afd78 , 
    R_d0b_1587d158 , 
    R_1190_13c09198 , 
    R_132a_13d44bb8 , 
    R_17af_123b9d58 , 
    R_1949_140b51d8 , 
    R_815_158140f8 , 
    R_a48_13bed6b8 , 
    R_e34_13cd7e38 , 
    R_1067_13b93ab8 , 
    R_1453_15ff99c8 , 
    R_1686_1008c258 , 
    R_af8_148696b8 , 
    R_d84_156b3e78 , 
    R_765_13df9678 , 
    R_1117_140b2398 , 
    R_13a3_123bd598 , 
    R_1736_117f1218 , 
    R_19c2_14871098 , 
    R_d3e_14870198 , 
    R_71f_123b6e78 , 
    R_b3e_11631138 , 
    R_115d_1008bd58 , 
    R_135d_13cd9d78 , 
    R_177c_11629258 , 
    R_197c_13bec8f8 , 
    R_96e_1162bff8 , 
    R_f0e_17010f68 , 
    R_8ef_13dd96d8 , 
    R_f8d_13cd51d8 , 
    R_152d_13d1f8d8 , 
    R_15ac_12fc1418 , 
    R_ee8_13d55658 , 
    R_994_13c086f8 , 
    R_8c9_1162f838 , 
    R_fb3_11c6c7b8 , 
    R_1507_14b218f8 , 
    R_15d2_11c6e978 , 
    R_ed3_13b93018 , 
    R_9a9_140ac3f8 , 
    R_8b4_150e2e38 , 
    R_fc8_14875238 , 
    R_14f2_13cd1718 , 
    R_15e7_150e0e58 , 
    R_c1a_13d3c198 , 
    R_5fb_156b22f8 , 
    R_643_117ea698 , 
    R_c62_1162c598 , 
    R_1239_15817938 , 
    R_1281_158887d8 , 
    R_1858_13bea9b8 , 
    R_18a0_123bfcf8 , 
    R_98c_13c21f18 , 
    R_ef0_13d51418 , 
    R_8d1_12fc06f8 , 
    R_fab_14a127f8 , 
    R_150f_15817398 , 
    R_15ca_156b71b8 , 
    R_c95_123be2b8 , 
    R_be7_1162d858 , 
    R_5c8_15feeca8 , 
    R_676_13d37e18 , 
    R_1206_13ddcc98 , 
    R_12b4_10087938 , 
    R_1825_1486a298 , 
    R_18d3_17018f88 , 
    R_d5b_150e0958 , 
    R_b21_14b21e98 , 
    R_73c_13bec858 , 
    R_1140_13b98798 , 
    R_137a_13dd7018 , 
    R_175f_15ff7f88 , 
    R_1999_117f2118 , 
    R_d4a_13df40d8 , 
    R_b32_13c268d8 , 
    R_72b_11632c18 , 
    R_1151_11638898 , 
    R_1369_117f5138 , 
    R_1770_124c2a58 , 
    R_1988_150dfaf8 , 
    R_db1_13bf06d8 , 
    R_792_13ccb638 , 
    R_acb_13d2a378 , 
    R_10ea_13d2b598 , 
    R_13d0_1700b388 , 
    R_1709_1162a298 , 
    R_19ef_150de1f8 , 
    R_ae3_14b24738 , 
    R_d99_156abef8 , 
    R_77a_13c0f3b8 , 
    R_1102_11632358 , 
    R_13b8_13c29c18 , 
    R_1721_14870f58 , 
    R_19d7_13de38b8 , 
    R_6d8_1580ebf8 , 
    R_566_140b4f58 , 
    R_cf7_13d26778 , 
    R_b85_13df3958 , 
    R_11a4_140b1178 , 
    R_1316_13c24718 , 
    R_17c3_13df1e78 , 
    R_1935_14a13798 , 
    R_a0d_14a0f198 , 
    R_850_1700cbe8 , 
    R_e6f_117ee6f8 , 
    R_102c_156ae3d8 , 
    R_148e_17014208 , 
    R_164b_123b8638 , 
    R_f2f_13ccded8 , 
    R_910_158144b8 , 
    R_94d_13de1dd8 , 
    R_f6c_140aca38 , 
    R_154e_158131f8 , 
    R_158b_123b5078 , 
    R_70c_1162a338 , 
    R_b51_13df4c18 , 
    R_d2b_123bacf8 , 
    R_1170_13ddca18 , 
    R_134a_123bdb38 , 
    R_178f_14a0df78 , 
    R_1969_13c0e918 , 
    R_ec1_13c0ddd8 , 
    R_8a2_13dd9638 , 
    R_9bb_14a13d38 , 
    R_fda_14876098 , 
    R_14e0_117ea9b8 , 
    R_15f9_13d4fcf8 , 
    R_d3b_150e4a58 , 
    R_71c_150dba98 , 
    R_b41_100844b8 , 
    R_1160_14a16498 , 
    R_135a_156b8838 , 
    R_177f_13ccedd8 , 
    R_1979_156ad7f8 , 
    R_80a_11c686b8 , 
    R_a53_13d54ed8 , 
    R_e29_124c3138 , 
    R_1072_13d5c598 , 
    R_1448_156b5098 , 
    R_1691_13bf8478 , 
    R_1a67_13d3a898 , 
    R_aa1_13ccbd18 , 
    R_7bc_13ccc218 , 
    R_ddb_15812618 , 
    R_10c0_15816d58 , 
    R_13fa_14b29a58 , 
    R_16df_10084eb8 , 
    R_1a19_11c70a98 , 
    R_a1e_13de1338 , 
    R_83f_123bc5f8 , 
    R_e5e_13c25258 , 
    R_103d_123b2738 , 
    R_147d_13d53e98 , 
    R_165c_123b57f8 , 
    R_c74_14b242d8 , 
    R_c08_13ded7d8 , 
    R_5e9_15816178 , 
    R_655_13c026b8 , 
    R_1227_123b72d8 , 
    R_1293_1008c6b8 , 
    R_1846_13c22af8 , 
    R_18b2_150dd4d8 , 
    R_a14_11632038 , 
    R_849_123c1af8 , 
    R_e68_15887658 , 
    R_1033_13bf8518 , 
    R_1487_1007fc38 , 
    R_1652_11635418 , 
    R_68e_11630eb8 , 
    R_bcf_1486c4f8 , 
    R_cad_150e5c78 , 
    R_5b0_13d20c38 , 
    R_11ee_13df5938 , 
    R_12cc_156aee78 , 
    R_180d_13d29dd8 , 
    R_18eb_13cd2bb8 , 
    R_7e9_13b903b8 , 
    R_e08_14a11498 , 
    R_a74_13c02a78 , 
    R_1093_123bddb8 , 
    R_1427_1580dd98 , 
    R_16b2_123b89f8 , 
    R_1a46_150dff58 , 
    R_c81_140ac718 , 
    R_bfb_117e8f78 , 
    R_5dc_13cd21b8 , 
    R_662_11c6af58 , 
    R_121a_13dd6bb8 , 
    R_12a0_156af7d8 , 
    R_1839_10083a18 , 
    R_18bf_13cd63f8 , 
    R_d4d_14b1c218 , 
    R_b2f_14a168f8 , 
    R_72e_15885178 , 
    R_114e_14866878 , 
    R_136c_13d5ce58 , 
    R_176d_15883e18 , 
    R_198b_123ba938 , 
    R_bb0_11635198 , 
    R_6ad_14b295f8 , 
    R_591_123b56b8 , 
    R_ccc_13c02f78 , 
    R_11cf_13dedd78 , 
    R_12eb_156ab598 , 
    R_17ee_117f2a78 , 
    R_190a_1162b238 , 
    R_7d4_14a0fe18 , 
    R_df3_14b1e478 , 
    R_a89_13dd9278 , 
    R_10a8_13d52958 , 
    R_1412_11c6f198 , 
    R_16c7_13d27d58 , 
    R_1a31_140b9d78 , 
    R_c19_1700d408 , 
    R_5fa_13df88b8 , 
    R_644_13d23938 , 
    R_c63_1162e258 , 
    R_1238_13df9a38 , 
    R_1282_13c2acf8 , 
    R_1857_13cd2ed8 , 
    R_18a1_156aefb8 , 
    R_6f0_140ae658 , 
    R_b6d_123b4178 , 
    R_d0f_150df0f8 , 
    R_118c_14a17898 , 
    R_132e_13bed758 , 
    R_17ab_13cd0d18 , 
    R_194d_1008c438 , 
    R_802_13d3e5d8 , 
    R_e21_14a0aaf8 , 
    R_a5b_13bf7e38 , 
    R_107a_13d1ed98 , 
    R_1440_124c4d58 , 
    R_1699_140b0318 , 
    R_1a5f_124c5618 , 
    R_8fc_13bebd18 , 
    R_961_12fbe358 , 
    R_f1b_13ddafd8 , 
    R_f80_1486f478 , 
    R_153a_116341f8 , 
    R_159f_1008d338 , 
    R_ada_15812f78 , 
    R_da2_156b5ef8 , 
    R_783_123ba898 , 
    R_10f9_123b7a58 , 
    R_13c1_13d3bfb8 , 
    R_1718_156b8018 , 
    R_19e0_13dd4ef8 , 
    R_6cb_117f2258 , 
    R_573_1162dfd8 , 
    R_cea_13d5be18 , 
    R_b92_13c01998 , 
    R_11b1_1700a208 , 
    R_1309_117e8898 , 
    R_17d0_156b8d38 , 
    R_1928_14a0f738 , 
    R_eb1_156b8f18 , 
    R_892_11c69018 , 
    R_9cb_13bed1b8 , 
    R_fea_13d2b3b8 , 
    R_14d0_13ccf698 , 
    R_1609_13cd30b8 , 
    R_67f_13cd88d8 , 
    R_c9e_1580ee78 , 
    R_bde_123b3138 , 
    R_5bf_117f0b38 , 
    R_11fd_1162f3d8 , 
    R_12bd_13bf9698 , 
    R_181c_13bf7758 , 
    R_18dc_15817258 , 
    R_c8c_13b97258 , 
    R_bf0_13c26d38 , 
    R_5d1_14875af8 , 
    R_66d_1700eda8 , 
    R_120f_156b0a98 , 
    R_12ab_1486c278 , 
    R_182e_116366d8 , 
    R_18ca_11c708b8 , 
    R_f2e_13dddb98 , 
    R_90f_13b8e3d8 , 
    R_94e_117f3c98 , 
    R_f6d_13bf7a78 , 
    R_154d_13df8c78 , 
    R_158c_13d278f8 , 
    R_702_13de3598 , 
    R_b5b_13d45bf8 , 
    R_d21_156ac038 , 
    R_117a_14b292d8 , 
    R_1340_123bbab8 , 
    R_1799_13df1018 , 
    R_195f_13b92e38 , 
    R_d38_156afaf8 , 
    R_719_13d1d498 , 
    R_b44_13df7238 , 
    R_1163_13b91358 , 
    R_1357_13d5bcd8 , 
    R_1782_1486c138 , 
    R_1976_14b1de38 , 
    R_695_13b93b58 , 
    R_bc8_13dfb3d8 , 
    R_cb4_15817078 , 
    R_5a9_156b6998 , 
    R_11e7_13bf3298 , 
    R_12d3_14b28338 , 
    R_1806_123b6dd8 , 
    R_18f2_13d40338 , 
    R_a06_158876f8 , 
    R_857_14874dd8 , 
    R_e76_13bf0958 , 
    R_1025_13d59438 , 
    R_1495_14870238 , 
    R_1644_15ff4d88 , 
    R_6fb_156b9378 , 
    R_b62_123bb298 , 
    R_d1a_117ee1f8 , 
    R_1181_148748d8 , 
    R_1339_1580de38 , 
    R_17a0_13dd7478 , 
    R_1958_156ae5b8 , 
    R_97a_117eaff8 , 
    R_f02_13d538f8 , 
    R_8e3_13c107b8 , 
    R_f99_1580efb8 , 
    R_1521_148676d8 , 
    R_15b8_13b93e78 , 
    R_829_13b954f8 , 
    R_a34_156b03b8 , 
    R_e48_15813d38 , 
    R_1053_13cd3478 , 
    R_1467_13b8be58 , 
    R_1672_13cd1df8 , 
    R_e89_13de0078 , 
    R_9f3_156b0598 , 
    R_86a_13b94378 , 
    R_1012_123bf618 , 
    R_14a8_13becdf8 , 
    R_1631_1486c9f8 , 
    R_acd_1008bfd8 , 
    R_daf_123b59d8 , 
    R_790_13d2bd18 , 
    R_10ec_1700b6a8 , 
    R_13ce_13df2a58 , 
    R_170b_14b26178 , 
    R_19ed_148709b8 , 
    R_a31_13cd7d98 , 
    R_82c_140b1e98 , 
    R_e4b_116316d8 , 
    R_1050_13d3d138 , 
    R_146a_123bd318 , 
    R_166f_140ad118 , 
    R_eac_1007f418 , 
    R_88d_13bf99b8 , 
    R_9d0_17010748 , 
    R_fef_1580b138 , 
    R_14cb_13d44258 , 
    R_160e_11632a38 , 
    R_826_13c24cb8 , 
    R_a37_158112b8 , 
    R_e45_15fee168 , 
    R_1056_15fedc68 , 
    R_1464_13d3fa78 , 
    R_1675_14b28dd8 , 
    R_eb6_11c69518 , 
    R_897_11c69338 , 
    R_9c6_156ad258 , 
    R_fe5_14b1f4b8 , 
    R_14d5_14871a98 , 
    R_1604_13beed38 , 
    R_9ef_14a126b8 , 
    R_e8d_13c07578 , 
    R_86e_13ded738 , 
    R_100e_100810d8 , 
    R_14ac_13cce158 , 
    R_162d_13c0adb8 , 
    R_7cb_14a0acd8 , 
    R_dea_123c0798 , 
    R_a92_13d25238 , 
    R_10b1_13d55478 , 
    R_1409_1587f638 , 
    R_16d0_13c02ed8 , 
    R_1a28_14a12398 , 
    R_ee0_13d1ffb8 , 
    R_99c_14a0f418 , 
    R_8c1_14b25818 , 
    R_fbb_123b70f8 , 
    R_14ff_1580bf98 , 
    R_15da_140ba138 , 
    R_687_14b23fb8 , 
    R_bd6_13dd71f8 , 
    R_ca6_123bd098 , 
    R_5b7_117e8cf8 , 
    R_11f5_15815318 , 
    R_12c5_14a0f7d8 , 
    R_1814_170116e8 , 
    R_18e4_12fc1d78 , 
    R_812_12fc0018 , 
    R_a4b_13bf22f8 , 
    R_e31_13bee338 , 
    R_106a_13d56a58 , 
    R_1450_1580a738 , 
    R_1689_14a0c218 , 
    R_e85_156aa878 , 
    R_9f7_13d246f8 , 
    R_866_15ffb868 , 
    R_1016_156af698 , 
    R_14a4_11c6ec98 , 
    R_1635_15ff7588 , 
    R_8ee_140ae338 , 
    R_96f_13d3b8d8 , 
    R_f0d_13d4fa78 , 
    R_f8e_13d541b8 , 
    R_152c_156b2258 , 
    R_15ad_13d58218 , 
    R_9de_124c3458 , 
    R_e9e_123b9038 , 
    R_87f_117f0958 , 
    R_ffd_13c27f58 , 
    R_14bd_13cd71b8 , 
    R_161c_156b6178 , 
    R_aec_14866b98 , 
    R_d90_10081718 , 
    R_771_1007ee78 , 
    R_110b_14b24f58 , 
    R_13af_158110d8 , 
    R_172a_11c6feb8 , 
    R_19ce_11c6fc38 , 
    R_6d4_15ff47e8 , 
    R_56a_17018268 , 
    R_cf3_150e21b8 , 
    R_b89_13cd67b8 , 
    R_11a8_13c0ab38 , 
    R_1312_15881758 , 
    R_17c7_1580cf38 , 
    R_1931_11c6b4f8 , 
    R_7be_13d51918 , 
    R_ddd_10083fb8 , 
    R_a9f_140b7b18 , 
    R_10be_1162c138 , 
    R_13fc_13b967b8 , 
    R_16dd_15ffb728 , 
    R_1a1b_13d3ab18 , 
    R_a2e_1580aeb8 , 
    R_82f_14b26cb8 , 
    R_e4e_13dec798 , 
    R_104d_13de2af8 , 
    R_146d_156b1998 , 
    R_166c_117f5958 , 
    R_d50_156b51d8 , 
    R_b2c_12fc0478 , 
    R_731_15ffaa08 , 
    R_114b_13ddbed8 , 
    R_136f_11c6c718 , 
    R_176a_11628f38 , 
    R_198e_150e3518 , 
    R_ed9_15ff7948 , 
    R_9a3_13c1fad8 , 
    R_8ba_116386b8 , 
    R_fc2_1700f7a8 , 
    R_14f8_117f15d8 , 
    R_15e1_150dcd58 , 
    R_b16_13c1c1f8 , 
    R_d66_13b8b1d8 , 
    R_747_158864d8 , 
    R_1135_156b68f8 , 
    R_1385_1580b278 , 
    R_1754_156add98 , 
    R_19a4_13d4fd98 , 
    R_823_11c6f2d8 , 
    R_a3a_14871318 , 
    R_e42_156ade38 , 
    R_1059_13c0f318 , 
    R_1461_14a1a138 , 
    R_1678_14a0fd78 , 
    R_8d9_158837d8 , 
    R_984_15882d38 , 
    R_ef8_15816998 , 
    R_fa3_15815458 , 
    R_1517_156ad898 , 
    R_15c2_11630c38 , 
    R_af3_13beae18 , 
    R_d89_117e8938 , 
    R_76a_123bceb8 , 
    R_1112_13c20c58 , 
    R_13a8_117f4a58 , 
    R_1731_1008a818 , 
    R_19c7_13d38bd8 , 
    R_b04_156aed38 , 
    R_d78_13cd7758 , 
    R_759_11629938 , 
    R_1123_15ffb908 , 
    R_1397_13d37a58 , 
    R_1742_13d237f8 , 
    R_19b6_14b20778 , 
    R_c64_13c1fdf8 , 
    R_c18_12fc23b8 , 
    R_5f9_13b8f238 , 
    R_645_140b2118 , 
    R_1237_1162dad8 , 
    R_1283_14a18798 , 
    R_1856_117f4878 , 
    R_18a2_13d53998 , 
    R_f2d_100818f8 , 
    R_90e_11629898 , 
    R_94f_15888738 , 
    R_f6e_14a188d8 , 
    R_154c_14a147d8 , 
    R_158d_15ff0a08 , 
    R_9eb_117ef2d8 , 
    R_e91_1580e3d8 , 
    R_872_13c0c7f8 , 
    R_100a_117f81f8 , 
    R_14b0_124c2f58 , 
    R_1629_14a0b6d8 , 
    R_656_15886bb8 , 
    R_c75_156b0db8 , 
    R_c07_124c4cb8 , 
    R_5e8_1162f298 , 
    R_1226_13b8e018 , 
    R_1294_13b91ad8 , 
    R_1845_13cd83d8 , 
    R_18b3_13d1e118 , 
    R_ba0_156b4698 , 
    R_6bd_13c0ec38 , 
    R_581_13d1d8f8 , 
    R_cdc_13cd9378 , 
    R_11bf_123b6c98 , 
    R_12fb_150e3018 , 
    R_17de_14b20458 , 
    R_191a_123b2cd8 , 
    R_d5e_14a10278 , 
    R_b1e_13df7418 , 
    R_73f_1587b998 , 
    R_113d_13d58498 , 
    R_137d_14a11b78 , 
    R_175c_1587b218 , 
    R_199c_17017408 , 
    R_b09_15884f98 , 
    R_d73_1580b4f8 , 
    R_754_15811d58 , 
    R_1128_10084d78 , 
    R_1392_14a15db8 , 
    R_1747_17018588 , 
    R_19b1_13dd9f98 , 
    R_d35_14a11858 , 
    R_716_156b9c38 , 
    R_b47_140af4b8 , 
    R_1166_13ccdcf8 , 
    R_1354_13d41738 , 
    R_1785_1162d218 , 
    R_1973_14a18338 , 
    R_a2b_13c1e6d8 , 
    R_832_13df5c58 , 
    R_e51_156ab278 , 
    R_104a_14a108b8 , 
    R_1470_15887bf8 , 
    R_1669_158828d8 , 
    R_e81_1007dc58 , 
    R_9fb_1486fb58 , 
    R_862_156ab138 , 
    R_101a_13d5a798 , 
    R_14a0_13d38818 , 
    R_1639_1162abf8 , 
    R_ba5_140b4af8 , 
    R_6b8_1580d898 , 
    R_586_15ff8488 , 
    R_cd7_156b7e38 , 
    R_11c4_117ecad8 , 
    R_12f6_17015ba8 , 
    R_17e3_13c1dd78 , 
    R_1915_14a17f78 , 
    R_aff_140aba98 , 
    R_d7d_148714f8 , 
    R_75e_10084418 , 
    R_111e_11635918 , 
    R_139c_1580e0b8 , 
    R_173d_13deffd8 , 
    R_19bb_13df9df8 , 
    R_7dd_13d28898 , 
    R_dfc_156b9ff8 , 
    R_a80_13ddc8d8 , 
    R_109f_13cd2cf8 , 
    R_141b_12fc10f8 , 
    R_16be_13bf0098 , 
    R_1a3a_156b79d8 , 
    R_9d5_15ff1908 , 
    R_ea7_14a124d8 , 
    R_888_13deebd8 , 
    R_ff4_13cd7b18 , 
    R_14c6_13cd5d18 , 
    R_1613_123bc198 , 
    R_677_13c0c758 , 
    R_c96_13c0d838 , 
    R_be6_1162cf98 , 
    R_5c7_1162f1f8 , 
    R_1205_156b94b8 , 
    R_12b5_158816b8 , 
    R_1824_13c04f58 , 
    R_18d4_13beb958 , 
    R_f1a_124c4f38 , 
    R_8fb_13c1e9f8 , 
    R_962_14a15ef8 , 
    R_f81_1580d438 , 
    R_1539_14b267b8 , 
    R_15a0_15ff32a8 , 
    R_d28_156b3fb8 , 
    R_709_117ea4b8 , 
    R_b54_13c04c38 , 
    R_1173_15810778 , 
    R_1347_13dd5f38 , 
    R_1792_13d39858 , 
    R_1966_12fc2098 , 
    R_a1b_123c17d8 , 
    R_842_13bf4738 , 
    R_e61_13cd0958 , 
    R_103a_13ccdbb8 , 
    R_1480_117f1e98 , 
    R_1659_13c1fcb8 , 
    R_820_17013088 , 
    R_a3d_11c6bc78 , 
    R_e3f_123c0e78 , 
    R_105c_13dd87d8 , 
    R_145e_13d5a3d8 , 
    R_167b_14a19878 , 
    R_ebb_13def998 , 
    R_89c_1486e898 , 
    R_9c1_13cd04f8 , 
    R_fe0_15fee7a8 , 
    R_14da_13b95818 , 
    R_15ff_117f1538 , 
    R_8d0_13ccd078 , 
    R_98d_13cceab8 , 
    R_eef_15ff2308 , 
    R_fac_13df65b8 , 
    R_150e_13bed398 , 
    R_15cb_1580a558 , 
    R_663_13c24218 , 
    R_c82_11633bb8 , 
    R_bfa_117f1d58 , 
    R_5db_13c0d798 , 
    R_1219_156b0f98 , 
    R_12a1_15811e98 , 
    R_1838_123c2098 , 
    R_18c0_13ddb258 , 
    R_bbb_13c08dd8 , 
    R_6a2_14870cd8 , 
    R_59c_1700ffc8 , 
    R_cc1_13d5b0f8 , 
    R_11da_14b1dcf8 , 
    R_12e0_14b29c38 , 
    R_17f9_13ddb438 , 
    R_18ff_1162d538 , 
    R_ecc_123bde58 , 
    R_9b0_1587f458 , 
    R_8ad_10082e38 , 
    R_fcf_14a0e798 , 
    R_14eb_140ad258 , 
    R_15ee_117f3158 , 
    R_d13_13c25e38 , 
    R_6f4_156b4918 , 
    R_b69_11c6e8d8 , 
    R_1188_13cd35b8 , 
    R_1332_11637d58 , 
    R_17a7_117f6a38 , 
    R_1951_156b6b78 , 
    R_acf_13d503d8 , 
    R_dad_13cd3838 , 
    R_78e_13b929d8 , 
    R_10ee_1587c438 , 
    R_13cc_1587b3f8 , 
    R_170d_12fbf9d8 , 
    R_19eb_15ff53c8 , 
    R_8c8_12fbe038 , 
    R_ee7_13c03dd8 , 
    R_995_13d50518 , 
    R_fb4_156b0e58 , 
    R_1506_156b9e18 , 
    R_15d3_123b5ed8 , 
    R_b9b_13dfa118 , 
    R_6c2_14b1d618 , 
    R_57c_13d464b8 , 
    R_ce1_13d27358 , 
    R_11ba_13cda458 , 
    R_1300_13dec478 , 
    R_17d9_156af918 , 
    R_191f_14a0d578 , 
    R_7e4_117f6c18 , 
    R_e03_13b8c718 , 
    R_a79_13d52db8 , 
    R_1098_13cd2438 , 
    R_1422_13cd7f78 , 
    R_16b7_14b28518 , 
    R_1a41_150e4d78 , 
    R_ae5_17012048 , 
    R_d97_1162ab58 , 
    R_778_13d52098 , 
    R_1104_13dd7a18 , 
    R_13b6_14a17118 , 
    R_1723_13d50018 , 
    R_19d5_117edc58 , 
    R_d53_13c0ae58 , 
    R_b29_13b95c78 , 
    R_734_14a0f558 , 
    R_1148_117f6218 , 
    R_1372_11c6cd58 , 
    R_1767_11c691f8 , 
    R_1991_13cd58b8 , 
    R_f2c_15814d78 , 
    R_90d_158848b8 , 
    R_950_140b3798 , 
    R_f6f_14a1a318 , 
    R_154b_11632218 , 
    R_158e_14a0b1d8 , 
    R_ec6_13d37b98 , 
    R_8a7_1580e6f8 , 
    R_9b6_14a0cc18 , 
    R_fd5_1580cc18 , 
    R_14e5_13b8fd78 , 
    R_15f4_170165a8 , 
    R_7c0_100854f8 , 
    R_ddf_13b92898 , 
    R_a9d_1162c318 , 
    R_10bc_140b7d98 , 
    R_13fe_13cd60d8 , 
    R_16db_156aaf58 , 
    R_1a1d_13cd9ff8 , 
    R_7f5_13b9a1d8 , 
    R_e14_123bf078 , 
    R_a68_150dbbd8 , 
    R_1087_1587ad18 , 
    R_1433_13dd7978 , 
    R_16a6_13df8458 , 
    R_1a52_11c70778 , 
    R_646_156ad618 , 
    R_c65_10086538 , 
    R_c17_13ccb3b8 , 
    R_5f8_1580f418 , 
    R_1236_1587e558 , 
    R_1284_14a1a458 , 
    R_1855_10084a58 , 
    R_18a3_1700b1a8 , 
    R_69c_156b9058 , 
    R_bc1_13bee298 , 
    R_cbb_13ccbbd8 , 
    R_5a2_15813658 , 
    R_11e0_1587e878 , 
    R_12da_14b29d78 , 
    R_17ff_14a10b38 , 
    R_18f9_14a16718 , 
    R_adc_156ae6f8 , 
    R_da0_13bf5db8 , 
    R_781_13d42f98 , 
    R_10fb_10085778 , 
    R_13bf_123bf6b8 , 
    R_171a_150deb58 , 
    R_19de_117ef918 , 
    R_9e7_13d54578 , 
    R_e95_13d26ef8 , 
    R_876_13d41698 , 
    R_1006_13c08f18 , 
    R_14b4_1700e268 , 
    R_1625_13b96d58 , 
    R_807_13cd8478 , 
    R_e26_1700df48 , 
    R_a56_124c4ad8 , 
    R_1075_15883b98 , 
    R_1445_15880218 , 
    R_1694_13d218b8 , 
    R_1a64_13ccac38 , 
    R_a28_13cd9918 , 
    R_835_140b35b8 , 
    R_e54_14a179d8 , 
    R_1047_14b26df8 , 
    R_1473_156b60d8 , 
    R_1666_14a165d8 , 
    R_b0e_14a15818 , 
    R_d6e_14a0c998 , 
    R_74f_13c24678 , 
    R_112d_1162be18 , 
    R_138d_13b92258 , 
    R_174c_116339d8 , 
    R_19ac_14b1b4f8 , 
    R_bb5_13cd29d8 , 
    R_6a8_1162e618 , 
    R_596_13dd6398 , 
    R_cc7_123b4b78 , 
    R_11d4_15ff30c8 , 
    R_12e6_14a0ff58 , 
    R_17f3_13ddb578 , 
    R_1905_1486dfd8 , 
    R_baa_14a15278 , 
    R_6b3_17011288 , 
    R_58b_140b1c18 , 
    R_cd2_13d24dd8 , 
    R_11c9_14b25278 , 
    R_12f1_1587da18 , 
    R_17e8_1587c078 , 
    R_1910_12fc0978 , 
    R_66e_17014348 , 
    R_c8d_123b7ff8 , 
    R_bef_14a167b8 , 
    R_5d0_13c1db98 , 
    R_120e_13c0d518 , 
    R_12ac_13ccaf58 , 
    R_182d_140b0098 , 
    R_18cb_123b9e98 , 
    R_8b3_13c0d298 , 
    R_ed2_1580c538 , 
    R_9aa_124c51b8 , 
    R_fc9_13b8d118 , 
    R_14f1_150e8978 , 
    R_15e8_15884db8 , 
    R_8e2_13bf6858 , 
    R_97b_150e7a78 , 
    R_f01_14a13e78 , 
    R_f9a_116364f8 , 
    R_1520_1162d678 , 
    R_15b9_13d21a98 , 
    R_7fa_123bbbf8 , 
    R_e19_13d59ed8 , 
    R_a63_14a16678 , 
    R_1082_13c09d78 , 
    R_1438_13bf2398 , 
    R_16a1_14a16cb8 , 
    R_1a57_13c28a98 , 
    R_81d_1580d078 , 
    R_a40_123bcd78 , 
    R_e3c_117f2c58 , 
    R_105f_13de2558 , 
    R_145b_11633e38 , 
    R_167e_1486d858 , 
    R_7f0_13b90458 , 
    R_e0f_140ab138 , 
    R_a6d_117ee838 , 
    R_108c_13bf90f8 , 
    R_142e_11632538 , 
    R_16ab_140b8d38 , 
    R_1a4d_11c70bd8 , 
    R_7d6_14b1e3d8 , 
    R_df5_1580eab8 , 
    R_a87_14a10138 , 
    R_10a6_117efa58 , 
    R_1414_1162b9b8 , 
    R_16c5_14a10db8 , 
    R_1a33_1486ebb8 , 
    R_f0c_140b21b8 , 
    R_8ed_11636d18 , 
    R_970_13c0f818 , 
    R_f8f_11632fd8 , 
    R_152b_13beb778 , 
    R_15ae_123b2eb8 , 
    R_e6b_13b8ded8 , 
    R_a11_158133d8 , 
    R_84c_13bef918 , 
    R_1030_140b72f8 , 
    R_148a_140b0598 , 
    R_164f_13d52778 , 
    R_afa_123c0c98 , 
    R_d82_13cd1858 , 
    R_763_1580e298 , 
    R_1119_1587c118 , 
    R_13a1_158898b8 , 
    R_1738_11c6f878 , 
    R_19c0_1007ded8 , 
    R_e7d_15811538 , 
    R_9ff_13d245b8 , 
    R_85e_13cd3018 , 
    R_101e_13d5d8f8 , 
    R_149c_13d5a978 , 
    R_163d_13ccd438 , 
    R_b8d_156aae18 , 
    R_6d0_1162bb98 , 
    R_56e_10086e98 , 
    R_cef_14870eb8 , 
    R_11ac_13c24498 , 
    R_130e_14a17758 , 
    R_17cb_14a0e478 , 
    R_192d_123becb8 , 
    R_d32_13d20558 , 
    R_713_15882978 , 
    R_b4a_13d22cb8 , 
    R_1169_123b7c38 , 
    R_1351_14a14558 , 
    R_1788_13ccae18 , 
    R_1970_124c43f8 , 
    R_7cd_13d58df8 , 
    R_dec_156ae518 , 
    R_a90_13dd8058 , 
    R_10af_117f0818 , 
    R_140b_1580d1b8 , 
    R_16ce_117ebe58 , 
    R_1a2a_15810e58 , 
    R_e72_13c1e8b8 , 
    R_a0a_13d54438 , 
    R_853_123bd778 , 
    R_1029_13cd2898 , 
    R_1491_117f33d8 , 
    R_1648_15ff12c8 , 
    R_80f_13d449d8 , 
    R_a4e_13b8e798 , 
    R_e2e_13dd57b8 , 
    R_106d_13b8b598 , 
    R_144d_13cd65d8 , 
    R_168c_15ff1c28;
wire n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , 
     n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , 
     n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , 
     n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , 
     n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , 
     n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , 
     n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , 
     n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , 
     n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , 
     n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , 
     n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , 
     n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , 
     n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , 
     n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , 
     n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , 
     n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , 
     n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , 
     n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , 
     n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , 
     n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , 
     n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , 
     n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , 
     n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , 
     n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , 
     n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , 
     n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , 
     n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , 
     n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , 
     n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , 
     n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , 
     n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , 
     n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , 
     n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , 
     n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , 
     n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , 
     n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , 
     n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , 
     n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , 
     n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , 
     n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , 
     n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , 
     n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , 
     n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , 
     n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , 
     n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , 
     n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , 
     n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , 
     n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , 
     n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , 
     n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , 
     n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , 
     n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , 
     n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , 
     n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , 
     n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , 
     n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , 
     n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , 
     n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , 
     n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , 
     n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , 
     n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , 
     n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , 
     n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , 
     n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , 
     n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , 
     n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , 
     n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , 
     n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , 
     n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , 
     n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , 
     n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , 
     n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , 
     n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , 
     n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , 
     n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , 
     n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , 
     n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , 
     n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , 
     n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , 
     n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , 
     n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , 
     n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , 
     n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , 
     n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , 
     n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , 
     n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , 
     n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , 
     n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , 
     n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , 
     n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , 
     n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , 
     n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , 
     n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , 
     n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , 
     n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , 
     n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , 
     n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , 
     n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , 
     n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , 
     n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , 
     n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , 
     n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , 
     n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , 
     n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , 
     n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , 
     n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , 
     n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , 
     n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , 
     n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , 
     n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , 
     n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , 
     n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , 
     n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , 
     n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , 
     n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , 
     n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , 
     n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , 
     n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , 
     n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , 
     n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , 
     n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , 
     n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , 
     n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , 
     n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , 
     n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , 
     n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , 
     n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , 
     n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , 
     n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , 
     n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , 
     n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , 
     n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , 
     n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , 
     n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , 
     n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , 
     n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , 
     n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , 
     n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , 
     n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , 
     n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , 
     n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , 
     n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , 
     n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , 
     n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , 
     n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , 
     n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , 
     n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , 
     n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , 
     n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , 
     n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , 
     n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , 
     n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , 
     n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , 
     n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , 
     n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , 
     n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , 
     n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , 
     n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , 
     n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , 
     n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , 
     n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , 
     n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , 
     n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , 
     n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , 
     n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , 
     n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , 
     n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , 
     n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , 
     n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , 
     n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , 
     n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , 
     n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , 
     n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , 
     n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , 
     n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , 
     n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , 
     n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , 
     n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , 
     n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , 
     n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , 
     n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , 
     n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , 
     n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , 
     n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , 
     n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , 
     n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , 
     n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , 
     n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , 
     n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , 
     n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , 
     n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , 
     n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , 
     n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , 
     n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , 
     n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , 
     n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , 
     n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , 
     n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , 
     n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , 
     n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , 
     n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , 
     n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , 
     n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , 
     n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , 
     n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , 
     n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , 
     n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , 
     n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , 
     n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , 
     n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , 
     n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , 
     n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , 
     n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , 
     n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , 
     n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , 
     n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , 
     n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , 
     n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , 
     n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , 
     n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , 
     n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , 
     n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , 
     n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , 
     n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , 
     n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , 
     n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , 
     n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , 
     n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , 
     n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , 
     n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , 
     n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , 
     n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , 
     n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , 
     n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , 
     n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , 
     n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , 
     n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , 
     n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , 
     n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , 
     n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , 
     n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , 
     n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , 
     n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , 
     n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , 
     n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , 
     n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , 
     n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , 
     n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , 
     n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , 
     n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , 
     n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , 
     n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , 
     n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , 
     n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , 
     n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , 
     n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , 
     n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , 
     n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , 
     n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , 
     n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , 
     n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , 
     n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , 
     n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , 
     n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , 
     n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , 
     n16171 , n372368 , n372369 , n372370 , n372371 , n372372 , n372373 , n372374 , n372375 , n372376 , 
     n372377 , n372378 , n372379 , n372380 , n372381 , n372382 , n372383 , n372384 , n372385 , n372386 , 
     n372387 , n372388 , n372389 , n372390 , n372391 , n372392 , n372393 , n372394 , n372395 , n372396 , 
     n372397 , n372398 , n372399 , n372400 , n372401 , n372402 , n372403 , n372404 , n372405 , n372406 , 
     n372407 , n372408 , n372409 , n372410 , n372411 , n372412 , n372413 , n372414 , n372415 , n372416 , 
     n372417 , n372418 , n372419 , n372420 , n372421 , n372422 , n372423 , n372424 , n372425 , n372426 , 
     n372427 , n372428 , n372429 , n372430 , n372431 , n372432 , n372433 , n372434 , n372435 , n372436 , 
     n372437 , n372438 , n372439 , n372440 , n372441 , n372442 , n372443 , n372444 , n372445 , n372446 , 
     n372447 , n372448 , n372449 , n372450 , n372451 , n372452 , n372453 , n372454 , n372455 , n372456 , 
     n372457 , n372458 , n372459 , n372460 , n372461 , n372462 , n372463 , n372464 , n372465 , n372466 , 
     n372467 , n372468 , n372469 , n372470 , n372471 , n372472 , n372473 , n372474 , n372475 , n372476 , 
     n372477 , n372478 , n372479 , n372480 , n372481 , n372482 , n372483 , n372484 , n372485 , n372486 , 
     n372487 , n372488 , n372489 , n372490 , n372491 , n372492 , n372493 , n372494 , n372495 , n372496 , 
     n372497 , n372498 , n372499 , n372500 , n372501 , n372502 , n372503 , n372504 , n372505 , n372506 , 
     n372507 , n372508 , n372509 , n372510 , n372511 , n372512 , n372513 , n372514 , n372515 , n372516 , 
     n372517 , n372518 , n372519 , n372520 , n372521 , n372522 , n372523 , n372524 , n372525 , n372526 , 
     n372527 , n372528 , n372529 , n372530 , n372531 , n372532 , n372533 , n372534 , n372535 , n372536 , 
     n372537 , n372538 , n372539 , n372540 , n372541 , n372542 , n372543 , n372544 , n372545 , n372546 , 
     n372547 , n372548 , n372549 , n372550 , n372551 , n372552 , n372553 , n372554 , n372555 , n372556 , 
     n372557 , n372558 , n372559 , n372560 , n372561 , n372562 , n372563 , n372564 , n372565 , n372566 , 
     n372567 , n372568 , n372569 , n372570 , n372571 , n372572 , n372573 , n372574 , n372575 , n372576 , 
     n372577 , n372578 , n372579 , n372580 , n372581 , n372582 , n372583 , n372584 , n372585 , n372586 , 
     n372587 , n372588 , n372589 , n372590 , n372591 , n372592 , n372593 , n372594 , n372595 , n372596 , 
     n372597 , n372598 , n372599 , n372600 , n372601 , n372602 , n372603 , n372604 , n372605 , n372606 , 
     n372607 , n372608 , n372609 , n372610 , n372611 , n372612 , n372613 , n372614 , n372615 , n372616 , 
     n372617 , n372618 , n372619 , n372620 , n372621 , n372622 , n372623 , n372624 , n372625 , n372626 , 
     n372627 , n372628 , n372629 , n372630 , n372631 , n372632 , n372633 , n372634 , n372635 , n372636 , 
     n372637 , n372638 , n372639 , n372640 , n372641 , n372642 , n372643 , n372644 , n372645 , n372646 , 
     n372647 , n372648 , n372649 , n372650 , n372651 , n372652 , n372653 , n372654 , n372655 , n372656 , 
     n372657 , n372658 , n372659 , n372660 , n372661 , n372662 , n372663 , n372664 , n372665 , n372666 , 
     n372667 , n372668 , n372669 , n372670 , n372671 , n372672 , n372673 , n372674 , n372675 , n372676 , 
     n372677 , n372678 , n372679 , n372680 , n372681 , n372682 , n372683 , n372684 , n372685 , n372686 , 
     n372687 , n372688 , n372689 , n372690 , n372691 , n372692 , n372693 , n372694 , n372695 , n372696 , 
     n372697 , n372698 , n372699 , n372700 , n372701 , n372702 , n372703 , n372704 , n372705 , n372706 , 
     n372707 , n372708 , n372709 , n372710 , n372711 , n372712 , n372713 , n372714 , n372715 , n372716 , 
     n372717 , n372718 , n372719 , n372720 , n372721 , n372722 , n372723 , n372724 , n372725 , n372726 , 
     n372727 , n372728 , n372729 , n372730 , n372731 , n372732 , n372733 , n372734 , n372735 , n372736 , 
     n372737 , n372738 , n372739 , n372740 , n372741 , n372742 , n372743 , n372744 , n372745 , n372746 , 
     n372747 , n372748 , n372749 , n372750 , n372751 , n372752 , n372753 , n372754 , n372755 , n372756 , 
     n372757 , n372758 , n372759 , n372760 , n372761 , n372762 , n372763 , n372764 , n372765 , n372766 , 
     n372767 , n372768 , n372769 , n372770 , n372771 , n372772 , n372773 , n372774 , n372775 , n372776 , 
     n372777 , n372778 , n372779 , n372780 , n372781 , n372782 , n372783 , n372784 , n372785 , n372786 , 
     n372787 , n372788 , n372789 , n372790 , n372791 , n372792 , n372793 , n372794 , n372795 , n372796 , 
     n372797 , n372798 , n372799 , n372800 , n372801 , n372802 , n372803 , n372804 , n372805 , n372806 , 
     n372807 , n372808 , n372809 , n372810 , n372811 , n372812 , n372813 , n372814 , n372815 , n372816 , 
     n372817 , n372818 , n372819 , n372820 , n372821 , n372822 , n372823 , n372824 , n372825 , n372826 , 
     n372827 , n372828 , n372829 , n372830 , n372831 , n372832 , n372833 , n372834 , n372835 , n372836 , 
     n372837 , n372838 , n372839 , n372840 , n372841 , n372842 , n372843 , n372844 , n372845 , n372846 , 
     n372847 , n372848 , n372849 , n372850 , n372851 , n372852 , n372853 , n372854 , n372855 , n372856 , 
     n372857 , n372858 , n372859 , n372860 , n372861 , n372862 , n372863 , n372864 , n372865 , n372866 , 
     n372867 , n372868 , n372869 , n372870 , n372871 , n372872 , n372873 , n372874 , n372875 , n372876 , 
     n372877 , n372878 , n372879 , n372880 , n372881 , n372882 , n372883 , n372884 , n372885 , n372886 , 
     n372887 , n372888 , n372889 , n372890 , n372891 , n372892 , n372893 , n372894 , n372895 , n372896 , 
     n372897 , n372898 , n372899 , n372900 , n372901 , n372902 , n372903 , n372904 , n372905 , n372906 , 
     n372907 , n372908 , n372909 , n372910 , n372911 , n372912 , n372913 , n372914 , n372915 , n372916 , 
     n372917 , n372918 , n372919 , n372920 , n372921 , n372922 , n372923 , n372924 , n372925 , n372926 , 
     n372927 , n372928 , n372929 , n372930 , n372931 , n372932 , n372933 , n372934 , n372935 , n372936 , 
     n372937 , n372938 , n372939 , n372940 , n372941 , n372942 , n372943 , n372944 , n372945 , n372946 , 
     n372947 , n372948 , n372949 , n372950 , n372951 , n372952 , n372953 , n372954 , n372955 , n372956 , 
     n372957 , n372958 , n372959 , n372960 , n372961 , n372962 , n372963 , n372964 , n372965 , n372966 , 
     n372967 , n372968 , n372969 , n372970 , n372971 , n372972 , n372973 , n372974 , n372975 , n372976 , 
     n372977 , n372978 , n372979 , n372980 , n372981 , n372982 , n372983 , n372984 , n372985 , n372986 , 
     n372987 , n372988 , n372989 , n372990 , n372991 , n372992 , n372993 , n372994 , n372995 , n372996 , 
     n372997 , n372998 , n372999 , n373000 , n373001 , n373002 , n373003 , n373004 , n373005 , n373006 , 
     n373007 , n373008 , n373009 , n373010 , n373011 , n373012 , n373013 , n373014 , n373015 , n373016 , 
     n373017 , n373018 , n373019 , n373020 , n373021 , n373022 , n373023 , n373024 , n373025 , n373026 , 
     n373027 , n373028 , n373029 , n373030 , n373031 , n373032 , n373033 , n373034 , n373035 , n373036 , 
     n373037 , n373038 , n373039 , n373040 , n373041 , n373042 , n373043 , n373044 , n373045 , n373046 , 
     n373047 , n373048 , n373049 , n373050 , n373051 , n373052 , n373053 , n373054 , n373055 , n373056 , 
     n373057 , n373058 , n373059 , n373060 , n373061 , n373062 , n373063 , n373064 , n373065 , n373066 , 
     n373067 , n373068 , n373069 , n373070 , n373071 , n373072 , n373073 , n373074 , n373075 , n373076 , 
     n373077 , n373078 , n373079 , n373080 , n373081 , n373082 , n373083 , n373084 , n373085 , n373086 , 
     n373087 , n373088 , n373089 , n373090 , n373091 , n373092 , n373093 , n373094 , n373095 , n373096 , 
     n373097 , n373098 , n373099 , n373100 , n373101 , n373102 , n373103 , n373104 , n373105 , n373106 , 
     n373107 , n373108 , n373109 , n373110 , n373111 , n373112 , n373113 , n373114 , n373115 , n373116 , 
     n373117 , n373118 , n373119 , n373120 , n373121 , n373122 , n373123 , n373124 , n373125 , n373126 , 
     n373127 , n373128 , n373129 , n373130 , n373131 , n373132 , n373133 , n373134 , n373135 , n373136 , 
     n373137 , n373138 , n373139 , n373140 , n373141 , n373142 , n373143 , n373144 , n373145 , n373146 , 
     n373147 , n373148 , n373149 , n373150 , n373151 , n373152 , n373153 , n373154 , n373155 , n373156 , 
     n373157 , n373158 , n373159 , n373160 , n373161 , n373162 , n373163 , n373164 , n373165 , n373166 , 
     n373167 , n373168 , n373169 , n373170 , n373171 , n373172 , n373173 , n373174 , n373175 , n373176 , 
     n373177 , n373178 , n373179 , n373180 , n373181 , n373182 , n373183 , n373184 , n373185 , n373186 , 
     n373187 , n373188 , n373189 , n373190 , n373191 , n373192 , n373193 , n373194 , n373195 , n373196 , 
     n373197 , n373198 , n373199 , n373200 , n373201 , n373202 , n373203 , n373204 , n373205 , n373206 , 
     n373207 , n373208 , n373209 , n373210 , n373211 , n373212 , n373213 , n373214 , n373215 , n373216 , 
     n373217 , n373218 , n373219 , n373220 , n373221 , n373222 , n373223 , n373224 , n373225 , n373226 , 
     n373227 , n373228 , n373229 , n373230 , n373231 , n373232 , n373233 , n373234 , n373235 , n373236 , 
     n373237 , n373238 , n373239 , n373240 , n373241 , n373242 , n373243 , n373244 , n373245 , n373246 , 
     n373247 , n373248 , n373249 , n373250 , n373251 , n373252 , n373253 , n373254 , n373255 , n373256 , 
     n373257 , n373258 , n373259 , n373260 , n373261 , n373262 , n373263 , n373264 , n373265 , n373266 , 
     n373267 , n373268 , n373269 , n373270 , n373271 , n373272 , n373273 , n373274 , n373275 , n373276 , 
     n373277 , n373278 , n373279 , n373280 , n373281 , n373282 , n373283 , n373284 , n373285 , n373286 , 
     n373287 , n373288 , n373289 , n373290 , n373291 , n373292 , n373293 , n373294 , n373295 , n373296 , 
     n373297 , n373298 , n373299 , n373300 , n373301 , n373302 , n373303 , n373304 , n373305 , n373306 , 
     n373307 , n373308 , n373309 , n373310 , n373311 , n373312 , n373313 , n373314 , n373315 , n373316 , 
     n373317 , n373318 , n373319 , n373320 , n373321 , n373322 , n373323 , n373324 , n373325 , n373326 , 
     n373327 , n373328 , n373329 , n373330 , n373331 , n373332 , n373333 , n373334 , n373335 , n373336 , 
     n373337 , n373338 , n373339 , n373340 , n373341 , n373342 , n373343 , n373344 , n373345 , n373346 , 
     n373347 , n373348 , n373349 , n373350 , n373351 , n373352 , n373353 , n373354 , n373355 , n373356 , 
     n373357 , n373358 , n373359 , n373360 , n373361 , n373362 , n373363 , n373364 , n373365 , n373366 , 
     n373367 , n373368 , n373369 , n373370 , n373371 , n373372 , n373373 , n373374 , n373375 , n373376 , 
     n373377 , n373378 , n373379 , n373380 , n373381 , n373382 , n373383 , n373384 , n373385 , n373386 , 
     n373387 , n373388 , n373389 , n373390 , n373391 , n373392 , n373393 , n373394 , n373395 , n373396 , 
     n373397 , n373398 , n373399 , n373400 , n373401 , n373402 , n373403 , n373404 , n373405 , n373406 , 
     n373407 , n373408 , n373409 , n373410 , n373411 , n373412 , n373413 , n373414 , n373415 , n373416 , 
     n373417 , n373418 , n373419 , n373420 , n373421 , n373422 , n373423 , n373424 , n373425 , n373426 , 
     n373427 , n373428 , n373429 , n373430 , n373431 , n373432 , n373433 , n373434 , n373435 , n373436 , 
     n373437 , n373438 , n373439 , n373440 , n373441 , n373442 , n373443 , n373444 , n373445 , n373446 , 
     n373447 , n373448 , n373449 , n373450 , n373451 , n373452 , n373453 , n373454 , n373455 , n373456 , 
     n373457 , n373458 , n373459 , n373460 , n373461 , n373462 , n373463 , n373464 , n373465 , n373466 , 
     n373467 , n373468 , n373469 , n373470 , n373471 , n373472 , n373473 , n373474 , n373475 , n373476 , 
     n373477 , n373478 , n373479 , n373480 , n373481 , n373482 , n373483 , n373484 , n373485 , n373486 , 
     n373487 , n373488 , n373489 , n373490 , n373491 , n373492 , n373493 , n373494 , n373495 , n373496 , 
     n373497 , n373498 , n373499 , n373500 , n373501 , n373502 , n373503 , n373504 , n373505 , n373506 , 
     n373507 , n373508 , n373509 , n373510 , n373511 , n373512 , n373513 , n373514 , n373515 , n373516 , 
     n373517 , n373518 , n373519 , n373520 , n373521 , n373522 , n373523 , n373524 , n373525 , n373526 , 
     n373527 , n373528 , n373529 , n373530 , n373531 , n373532 , n373533 , n373534 , n373535 , n373536 , 
     n373537 , n373538 , n373539 , n373540 , n373541 , n373542 , n373543 , n373544 , n373545 , n373546 , 
     n373547 , n373548 , n373549 , n373550 , n373551 , n373552 , n373553 , n373554 , n373555 , n373556 , 
     n373557 , n373558 , n373559 , n373560 , n373561 , n373562 , n373563 , n373564 , n373565 , n373566 , 
     n373567 , n373568 , n373569 , n373570 , n373571 , n373572 , n373573 , n373574 , n373575 , n373576 , 
     n373577 , n373578 , n373579 , n373580 , n373581 , n373582 , n373583 , n373584 , n373585 , n373586 , 
     n373587 , n373588 , n373589 , n373590 , n373591 , n373592 , n373593 , n373594 , n373595 , n373596 , 
     n373597 , n373598 , n373599 , n373600 , n373601 , n373602 , n373603 , n373604 , n373605 , n373606 , 
     n373607 , n373608 , n373609 , n373610 , n373611 , n373612 , n373613 , n373614 , n373615 , n373616 , 
     n373617 , n373618 , n373619 , n373620 , n373621 , n373622 , n373623 , n373624 , n373625 , n373626 , 
     n373627 , n373628 , n373629 , n373630 , n373631 , n373632 , n373633 , n373634 , n373635 , n373636 , 
     n373637 , n373638 , n373639 , n373640 , n373641 , n373642 , n373643 , n373644 , n373645 , n373646 , 
     n373647 , n373648 , n373649 , n373650 , n373651 , n373652 , n373653 , n373654 , n373655 , n373656 , 
     n373657 , n373658 , n373659 , n373660 , n373661 , n373662 , n373663 , n373664 , n373665 , n373666 , 
     n373667 , n373668 , n373669 , n373670 , n373671 , n373672 , n373673 , n373674 , n373675 , n373676 , 
     n373677 , n373678 , n373679 , n373680 , n373681 , n373682 , n373683 , n373684 , n373685 , n373686 , 
     n373687 , n373688 , n373689 , n373690 , n373691 , n373692 , n373693 , n373694 , n17499 , n17500 , 
     n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , 
     n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , 
     n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , 
     n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , 
     n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , 
     n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , 
     n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , 
     n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , 
     n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , 
     n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , 
     n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , 
     n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , 
     n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , 
     n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , 
     n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , 
     n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , 
     n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , 
     n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , 
     n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , 
     n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , 
     n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , 
     n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , 
     n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , 
     n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , 
     n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , 
     n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , 
     n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , 
     n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , 
     n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , 
     n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , 
     n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , 
     n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , 
     n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , 
     n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , 
     n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , 
     n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , 
     n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , 
     n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , 
     n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , 
     n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , 
     n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , 
     n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , 
     n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , 
     n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , 
     n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , 
     n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , 
     n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , 
     n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , 
     n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , 
     n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , 
     n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , 
     n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , 
     n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , 
     n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , 
     n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , 
     n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , 
     n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , 
     n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , 
     n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , 
     n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , 
     n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , 
     n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , 
     n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , 
     n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , 
     n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , 
     n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , 
     n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , 
     n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , 
     n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , 
     n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , 
     n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , 
     n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , 
     n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , 
     n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , 
     n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , 
     n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , 
     n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , 
     n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , 
     n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , 
     n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , 
     n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , 
     n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , 
     n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , 
     n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , 
     n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , 
     n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , 
     n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , 
     n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , 
     n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , 
     n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , 
     n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , 
     n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , 
     n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , 
     n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , 
     n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , 
     n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , 
     n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , 
     n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , 
     n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , 
     n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , 
     n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , 
     n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , 
     n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , 
     n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , 
     n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , 
     n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , 
     n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , 
     n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , 
     n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , 
     n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , 
     n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , 
     n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , 
     n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , 
     n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , 
     n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , 
     n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , 
     n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , 
     n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , 
     n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , 
     n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , 
     n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , 
     n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , 
     n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , 
     n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , 
     n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , 
     n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , 
     n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , 
     n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , 
     n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , 
     n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , 
     n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , 
     n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , 
     n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , 
     n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , 
     n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , 
     n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , 
     n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , 
     n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , 
     n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , 
     n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , 
     n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , 
     n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , 
     n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , 
     n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , 
     n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , 
     n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , 
     n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , 
     n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , 
     n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , 
     n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , 
     n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , 
     n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , 
     n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , 
     n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , 
     n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , 
     n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , 
     n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , 
     n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , 
     n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , 
     n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , 
     n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , 
     n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , 
     n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , 
     n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , 
     n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , 
     n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , 
     n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , 
     n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , 
     n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , 
     n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , 
     n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , 
     n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , 
     n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , 
     n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , 
     n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , 
     n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , 
     n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , 
     n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , 
     n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , 
     n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , 
     n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , 
     n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , 
     n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , 
     n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , 
     n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , 
     n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , 
     n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , 
     n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , 
     n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , 
     n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , 
     n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , 
     n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , 
     n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , 
     n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , 
     n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , 
     n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , 
     n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , 
     n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , 
     n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , 
     n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , 
     n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , 
     n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , 
     n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , 
     n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , 
     n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , 
     n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , 
     n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , 
     n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , 
     n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , 
     n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , 
     n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , 
     n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , 
     n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , 
     n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , 
     n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , 
     n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , 
     n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , 
     n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , 
     n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , 
     n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , 
     n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , 
     n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , 
     n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , 
     n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , 
     n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , 
     n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , 
     n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , 
     n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , 
     n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , 
     n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , 
     n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , 
     n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , 
     n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , 
     n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , 
     n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , 
     n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , 
     n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , 
     n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , 
     n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , 
     n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , 
     n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , 
     n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , 
     n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , 
     n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , 
     n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , 
     n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , 
     n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , 
     n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , 
     n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , 
     n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , 
     n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , 
     n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , 
     n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , 
     n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , 
     n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , 
     n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , 
     n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , 
     n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , 
     n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , 
     n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , 
     n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , 
     n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , 
     n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , 
     n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , 
     n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , 
     n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , 
     n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , 
     n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , 
     n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , 
     n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , 
     n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , 
     n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , 
     n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , 
     n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , 
     n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , 
     n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , 
     n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , 
     n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , 
     n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , 
     n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , 
     n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , 
     n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , 
     n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , 
     n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , 
     n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , 
     n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , 
     n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , 
     n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , 
     n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , 
     n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , 
     n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , 
     n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , 
     n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , 
     n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , 
     n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , 
     n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , 
     n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , 
     n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , 
     n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , 
     n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , 
     n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , 
     n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , 
     n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , 
     n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , 
     n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , 
     n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , 
     n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , 
     n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , 
     n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , 
     n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , 
     n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , 
     n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , 
     n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , 
     n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , 
     n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , 
     n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , 
     n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , 
     n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , 
     n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , 
     n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , 
     n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , 
     n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , 
     n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , 
     n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , 
     n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , 
     n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , 
     n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , 
     n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , 
     n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , 
     n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , 
     n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , 
     n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , 
     n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , 
     n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , 
     n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , 
     n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , 
     n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , 
     n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , 
     n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , 
     n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , 
     n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , 
     n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , 
     n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , 
     n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , 
     n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , 
     n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , 
     n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , 
     n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , 
     n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , 
     n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , 
     n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , 
     n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , 
     n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , 
     n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , 
     n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , 
     n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , 
     n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , 
     n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , 
     n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , 
     n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , 
     n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , 
     n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , 
     n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , 
     n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , 
     n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , 
     n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , 
     n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , 
     n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , 
     n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , 
     n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , 
     n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , 
     n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , 
     n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , 
     n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , 
     n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , 
     n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , 
     n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , 
     n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , 
     n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , 
     n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , 
     n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , 
     n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , 
     n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , 
     n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , 
     n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , 
     n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , 
     n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , 
     n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , 
     n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , 
     n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , 
     n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , 
     n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , 
     n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , 
     n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , 
     n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , 
     n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , 
     n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , 
     n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , 
     n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , 
     n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , 
     n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , 
     n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , 
     n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , 
     n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , 
     n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , 
     n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , 
     n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , 
     n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , 
     n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , 
     n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , 
     n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , 
     n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , 
     n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , 
     n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , 
     n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , 
     n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , 
     n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , 
     n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , 
     n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , 
     n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , 
     n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , 
     n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , 
     n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , 
     n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , 
     n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , 
     n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , 
     n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , 
     n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , 
     n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , 
     n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , 
     n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , 
     n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , 
     n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , 
     n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , 
     n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , 
     n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , 
     n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , 
     n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , 
     n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , 
     n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , 
     n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , 
     n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , 
     n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , 
     n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , 
     n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , 
     n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , 
     n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , 
     n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , 
     n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , 
     n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , 
     n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , 
     n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , 
     n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , 
     n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , 
     n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , 
     n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , 
     n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , 
     n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , 
     n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , 
     n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , 
     n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , 
     n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , 
     n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , 
     n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , 
     n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , 
     n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , 
     n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , 
     n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , 
     n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , 
     n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , 
     n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , 
     n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , 
     n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , 
     n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , 
     n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , 
     n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , 
     n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , 
     n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , 
     n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , 
     n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , 
     n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , 
     n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , 
     n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , 
     n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , 
     n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , 
     n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , 
     n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , 
     n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , 
     n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , 
     n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , 
     n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , 
     n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , 
     n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , 
     n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , 
     n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , 
     n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , 
     n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , 
     n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , 
     n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , 
     n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , 
     n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , 
     n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , 
     n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , 
     n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , 
     n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , 
     n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , 
     n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , 
     n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , 
     n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , 
     n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , 
     n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , 
     n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , 
     n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , 
     n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , 
     n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , 
     n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , 
     n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , 
     n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , 
     n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , 
     n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , 
     n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , 
     n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , 
     n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , 
     n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , 
     n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , 
     n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , 
     n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , 
     n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , 
     n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , 
     n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , 
     n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , 
     n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , 
     n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , 
     n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , 
     n22841 , n22842 , n22843 , n379040 , n379041 , n379042 , n379043 , n379044 , n379045 , n379046 , 
     n379047 , n379048 , n379049 , n379050 , n379051 , n379052 , n379053 , n379054 , n379055 , n379056 , 
     n379057 , n379058 , n379059 , n379060 , n379061 , n379062 , n379063 , n379064 , n379065 , n379066 , 
     n379067 , n379068 , n379069 , n379070 , n379071 , n379072 , n379073 , n379074 , n379075 , n379076 , 
     n379077 , n379078 , n379079 , n379080 , n379081 , n379082 , n379083 , n379084 , n379085 , n379086 , 
     n379087 , n379088 , n379089 , n379090 , n379091 , n379092 , n379093 , n379094 , n379095 , n379096 , 
     n379097 , n379098 , n379099 , n379100 , n379101 , n379102 , n379103 , n379104 , n379105 , n379106 , 
     n379107 , n379108 , n379109 , n379110 , n379111 , n379112 , n379113 , n379114 , n379115 , n379116 , 
     n379117 , n379118 , n379119 , n379120 , n379121 , n379122 , n379123 , n379124 , n379125 , n379126 , 
     n379127 , n379128 , n379129 , n379130 , n379131 , n379132 , n379133 , n379134 , n379135 , n379136 , 
     n379137 , n379138 , n379139 , n379140 , n379141 , n379142 , n379143 , n379144 , n379145 , n379146 , 
     n379147 , n379148 , n379149 , n379150 , n379151 , n379152 , n379153 , n379154 , n379155 , n379156 , 
     n379157 , n379158 , n379159 , n379160 , n379161 , n379162 , n379163 , n379164 , n379165 , n379166 , 
     n379167 , n379168 , n379169 , n379170 , n379171 , n379172 , n379173 , n379174 , n379175 , n379176 , 
     n379177 , n379178 , n379179 , n379180 , n379181 , n379182 , n379183 , n379184 , n379185 , n379186 , 
     n379187 , n379188 , n379189 , n379190 , n379191 , n379192 , n379193 , n379194 , n379195 , n379196 , 
     n379197 , n379198 , n379199 , n379200 , n379201 , n379202 , n379203 , n379204 , n379205 , n379206 , 
     n379207 , n379208 , n379209 , n379210 , n379211 , n379212 , n379213 , n379214 , n379215 , n379216 , 
     n379217 , n379218 , n379219 , n379220 , n379221 , n379222 , n379223 , n379224 , n379225 , n379226 , 
     n379227 , n379228 , n379229 , n379230 , n379231 , n379232 , n379233 , n379234 , n379235 , n379236 , 
     n379237 , n379238 , n379239 , n379240 , n379241 , n379242 , n379243 , n379244 , n379245 , n379246 , 
     n379247 , n379248 , n379249 , n379250 , n379251 , n379252 , n379253 , n379254 , n379255 , n379256 , 
     n379257 , n379258 , n379259 , n379260 , n379261 , n379262 , n379263 , n379264 , n379265 , n379266 , 
     n379267 , n379268 , n379269 , n379270 , n379271 , n379272 , n379273 , n379274 , n379275 , n379276 , 
     n379277 , n379278 , n379279 , n379280 , n379281 , n379282 , n379283 , n379284 , n379285 , n379286 , 
     n379287 , n379288 , n379289 , n379290 , n379291 , n379292 , n379293 , n379294 , n379295 , n379296 , 
     n379297 , n379298 , n379299 , n379300 , n379301 , n379302 , n379303 , n379304 , n379305 , n379306 , 
     n379307 , n379308 , n379309 , n379310 , n379311 , n379312 , n379313 , n379314 , n379315 , n379316 , 
     n379317 , n379318 , n379319 , n379320 , n379321 , n379322 , n379323 , n379324 , n379325 , n379326 , 
     n379327 , n379328 , n379329 , n379330 , n379331 , n379332 , n379333 , n379334 , n379335 , n379336 , 
     n379337 , n379338 , n379339 , n379340 , n379341 , n379342 , n379343 , n379344 , n379345 , n379346 , 
     n379347 , n379348 , n379349 , n379350 , n379351 , n379352 , n379353 , n379354 , n379355 , n379356 , 
     n379357 , n379358 , n379359 , n379360 , n379361 , n379362 , n379363 , n379364 , n379365 , n379366 , 
     n379367 , n379368 , n379369 , n379370 , n379371 , n379372 , n379373 , n379374 , n379375 , n379376 , 
     n379377 , n379378 , n379379 , n379380 , n379381 , n379382 , n379383 , n379384 , n379385 , n379386 , 
     n379387 , n379388 , n379389 , n379390 , n379391 , n379392 , n379393 , n379394 , n379395 , n379396 , 
     n379397 , n379398 , n379399 , n379400 , n379401 , n379402 , n379403 , n379404 , n379405 , n379406 , 
     n379407 , n379408 , n379409 , n379410 , n379411 , n379412 , n379413 , n379414 , n379415 , n379416 , 
     n379417 , n379418 , n379419 , n379420 , n379421 , n379422 , n379423 , n379424 , n379425 , n379426 , 
     n379427 , n379428 , n379429 , n379430 , n379431 , n379432 , n379433 , n379434 , n379435 , n379436 , 
     n379437 , n379438 , n379439 , n379440 , n379441 , n379442 , n379443 , n379444 , n379445 , n379446 , 
     n379447 , n379448 , n379449 , n379450 , n379451 , n379452 , n379453 , n379454 , n379455 , n379456 , 
     n379457 , n379458 , n379459 , n379460 , n379461 , n379462 , n379463 , n379464 , n379465 , n379466 , 
     n379467 , n379468 , n379469 , n379470 , n379471 , n379472 , n379473 , n379474 , n379475 , n379476 , 
     n379477 , n379478 , n379479 , n379480 , n379481 , n379482 , n379483 , n379484 , n379485 , n379486 , 
     n379487 , n379488 , n379489 , n379490 , n379491 , n379492 , n379493 , n379494 , n379495 , n379496 , 
     n379497 , n379498 , n379499 , n379500 , n379501 , n379502 , n379503 , n379504 , n379505 , n379506 , 
     n379507 , n379508 , n379509 , n379510 , n379511 , n379512 , n379513 , n379514 , n379515 , n379516 , 
     n379517 , n379518 , n379519 , n379520 , n379521 , n379522 , n379523 , n379524 , n379525 , n379526 , 
     n379527 , n379528 , n379529 , n379530 , n379531 , n379532 , n379533 , n379534 , n379535 , n379536 , 
     n379537 , n379538 , n379539 , n379540 , n379541 , n379542 , n379543 , n379544 , n379545 , n379546 , 
     n379547 , n379548 , n379549 , n379550 , n379551 , n379552 , n379553 , n379554 , n379555 , n379556 , 
     n379557 , n379558 , n379559 , n379560 , n379561 , n379562 , n379563 , n379564 , n379565 , n379566 , 
     n379567 , n379568 , n379569 , n379570 , n379571 , n379572 , n379573 , n379574 , n379575 , n379576 , 
     n379577 , n379578 , n379579 , n379580 , n379581 , n379582 , n379583 , n379584 , n379585 , n379586 , 
     n379587 , n379588 , n379589 , n379590 , n379591 , n379592 , n379593 , n379594 , n379595 , n379596 , 
     n379597 , n379598 , n379599 , n379600 , n379601 , n379602 , n379603 , n379604 , n379605 , n379606 , 
     n379607 , n379608 , n379609 , n379610 , n379611 , n379612 , n379613 , n379614 , n379615 , n379616 , 
     n379617 , n379618 , n379619 , n379620 , n379621 , n379622 , n379623 , n379624 , n379625 , n379626 , 
     n379627 , n379628 , n379629 , n379630 , n379631 , n379632 , n379633 , n379634 , n379635 , n379636 , 
     n379637 , n379638 , n379639 , n379640 , n379641 , n379642 , n379643 , n379644 , n379645 , n379646 , 
     n379647 , n379648 , n379649 , n379650 , n379651 , n379652 , n379653 , n379654 , n379655 , n379656 , 
     n379657 , n379658 , n379659 , n379660 , n379661 , n379662 , n379663 , n379664 , n379665 , n379666 , 
     n379667 , n379668 , n379669 , n379670 , n379671 , n379672 , n379673 , n379674 , n379675 , n379676 , 
     n379677 , n379678 , n379679 , n379680 , n379681 , n379682 , n379683 , n379684 , n379685 , n379686 , 
     n379687 , n379688 , n379689 , n379690 , n379691 , n379692 , n379693 , n379694 , n379695 , n379696 , 
     n379697 , n379698 , n379699 , n379700 , n379701 , n379702 , n379703 , n379704 , n379705 , n379706 , 
     n379707 , n379708 , n379709 , n379710 , n379711 , n379712 , n379713 , n379714 , n379715 , n379716 , 
     n379717 , n379718 , n379719 , n379720 , n379721 , n379722 , n379723 , n379724 , n379725 , n379726 , 
     n379727 , n379728 , n379729 , n379730 , n379731 , n379732 , n379733 , n379734 , n379735 , n379736 , 
     n379737 , n379738 , n379739 , n379740 , n379741 , n379742 , n379743 , n379744 , n379745 , n379746 , 
     n379747 , n379748 , n379749 , n379750 , n379751 , n379752 , n379753 , n379754 , n379755 , n379756 , 
     n379757 , n379758 , n379759 , n379760 , n379761 , n379762 , n379763 , n379764 , n379765 , n379766 , 
     n379767 , n379768 , n379769 , n379770 , n379771 , n379772 , n379773 , n379774 , n379775 , n379776 , 
     n379777 , n379778 , n379779 , n379780 , n379781 , n379782 , n379783 , n379784 , n379785 , n379786 , 
     n379787 , n379788 , n379789 , n379790 , n379791 , n379792 , n379793 , n379794 , n379795 , n379796 , 
     n379797 , n379798 , n379799 , n379800 , n379801 , n379802 , n379803 , n379804 , n379805 , n379806 , 
     n379807 , n379808 , n379809 , n379810 , n379811 , n379812 , n379813 , n379814 , n379815 , n379816 , 
     n379817 , n379818 , n379819 , n379820 , n379821 , n379822 , n379823 , n379824 , n379825 , n379826 , 
     n379827 , n379828 , n379829 , n379830 , n379831 , n379832 , n379833 , n379834 , n379835 , n379836 , 
     n379837 , n379838 , n379839 , n379840 , n379841 , n379842 , n379843 , n379844 , n379845 , n379846 , 
     n379847 , n379848 , n379849 , n379850 , n379851 , n379852 , n379853 , n379854 , n379855 , n379856 , 
     n379857 , n379858 , n379859 , n379860 , n379861 , n379862 , n379863 , n379864 , n379865 , n379866 , 
     n379867 , n379868 , n379869 , n379870 , n379871 , n379872 , n379873 , n379874 , n379875 , n379876 , 
     n379877 , n379878 , n379879 , n379880 , n379881 , n379882 , n379883 , n379884 , n379885 , n379886 , 
     n379887 , n379888 , n379889 , n379890 , n379891 , n379892 , n379893 , n379894 , n379895 , n379896 , 
     n379897 , n379898 , n379899 , n379900 , n379901 , n379902 , n379903 , n379904 , n379905 , n379906 , 
     n379907 , n379908 , n379909 , n379910 , n379911 , n379912 , n379913 , n379914 , n379915 , n379916 , 
     n379917 , n379918 , n379919 , n379920 , n379921 , n379922 , n379923 , n379924 , n379925 , n379926 , 
     n379927 , n379928 , n379929 , n379930 , n379931 , n379932 , n379933 , n379934 , n379935 , n379936 , 
     n379937 , n379938 , n379939 , n379940 , n379941 , n379942 , n379943 , n379944 , n379945 , n379946 , 
     n379947 , n379948 , n379949 , n379950 , n379951 , n379952 , n379953 , n379954 , n379955 , n379956 , 
     n379957 , n379958 , n379959 , n379960 , n379961 , n379962 , n379963 , n379964 , n379965 , n379966 , 
     n379967 , n379968 , n379969 , n379970 , n379971 , n379972 , n379973 , n379974 , n379975 , n379976 , 
     n379977 , n379978 , n379979 , n379980 , n379981 , n379982 , n379983 , n379984 , n379985 , n379986 , 
     n379987 , n379988 , n379989 , n379990 , n379991 , n379992 , n379993 , n379994 , n379995 , n379996 , 
     n379997 , n379998 , n379999 , n380000 , n380001 , n380002 , n380003 , n380004 , n380005 , n380006 , 
     n380007 , n380008 , n380009 , n380010 , n380011 , n380012 , n380013 , n380014 , n380015 , n380016 , 
     n380017 , n380018 , n380019 , n380020 , n380021 , n380022 , n380023 , n380024 , n380025 , n380026 , 
     n380027 , n380028 , n380029 , n380030 , n380031 , n380032 , n380033 , n380034 , n380035 , n380036 , 
     n380037 , n380038 , n380039 , n380040 , n380041 , n380042 , n380043 , n380044 , n380045 , n380046 , 
     n380047 , n380048 , n380049 , n380050 , n380051 , n380052 , n380053 , n380054 , n380055 , n380056 , 
     n380057 , n380058 , n380059 , n380060 , n380061 , n380062 , n380063 , n380064 , n380065 , n380066 , 
     n380067 , n380068 , n380069 , n380070 , n380071 , n380072 , n380073 , n380074 , n380075 , n380076 , 
     n380077 , n380078 , n380079 , n380080 , n380081 , n380082 , n380083 , n380084 , n380085 , n380086 , 
     n380087 , n380088 , n380089 , n380090 , n380091 , n380092 , n380093 , n380094 , n380095 , n380096 , 
     n380097 , n380098 , n380099 , n380100 , n380101 , n380102 , n380103 , n380104 , n380105 , n380106 , 
     n380107 , n380108 , n380109 , n380110 , n380111 , n380112 , n380113 , n380114 , n380115 , n380116 , 
     n380117 , n380118 , n380119 , n380120 , n380121 , n380122 , n380123 , n380124 , n380125 , n380126 , 
     n380127 , n380128 , n380129 , n380130 , n380131 , n380132 , n380133 , n380134 , n380135 , n380136 , 
     n380137 , n380138 , n380139 , n380140 , n380141 , n380142 , n380143 , n380144 , n380145 , n380146 , 
     n380147 , n380148 , n380149 , n380150 , n380151 , n380152 , n380153 , n380154 , n380155 , n380156 , 
     n380157 , n380158 , n380159 , n380160 , n380161 , n380162 , n380163 , n380164 , n380165 , n380166 , 
     n380167 , n380168 , n380169 , n380170 , n380171 , n380172 , n380173 , n380174 , n380175 , n380176 , 
     n380177 , n380178 , n380179 , n380180 , n380181 , n380182 , n380183 , n380184 , n380185 , n380186 , 
     n380187 , n380188 , n380189 , n380190 , n380191 , n380192 , n380193 , n380194 , n380195 , n380196 , 
     n380197 , n380198 , n380199 , n380200 , n380201 , n380202 , n380203 , n380204 , n380205 , n380206 , 
     n380207 , n380208 , n380209 , n380210 , n380211 , n380212 , n380213 , n380214 , n380215 , n380216 , 
     n380217 , n380218 , n380219 , n380220 , n380221 , n380222 , n380223 , n380224 , n380225 , n380226 , 
     n380227 , n380228 , n380229 , n380230 , n380231 , n380232 , n380233 , n380234 , n380235 , n380236 , 
     n380237 , n380238 , n380239 , n380240 , n380241 , n380242 , n380243 , n380244 , n380245 , n380246 , 
     n380247 , n380248 , n380249 , n380250 , n380251 , n380252 , n380253 , n380254 , n380255 , n380256 , 
     n380257 , n380258 , n380259 , n380260 , n380261 , n380262 , n380263 , n380264 , n380265 , n380266 , 
     n380267 , n380268 , n380269 , n380270 , n380271 , n380272 , n380273 , n380274 , n380275 , n380276 , 
     n380277 , n380278 , n380279 , n380280 , n380281 , n380282 , n380283 , n380284 , n380285 , n380286 , 
     n380287 , n380288 , n380289 , n380290 , n380291 , n380292 , n380293 , n380294 , n380295 , n380296 , 
     n380297 , n380298 , n380299 , n380300 , n380301 , n380302 , n380303 , n380304 , n380305 , n380306 , 
     n380307 , n380308 , n380309 , n380310 , n380311 , n380312 , n380313 , n380314 , n380315 , n380316 , 
     n380317 , n380318 , n380319 , n380320 , n380321 , n380322 , n380323 , n380324 , n380325 , n380326 , 
     n380327 , n380328 , n380329 , n380330 , n380331 , n380332 , n380333 , n380334 , n380335 , n380336 , 
     n380337 , n380338 , n380339 , n380340 , n380341 , n380342 , n380343 , n380344 , n380345 , n380346 , 
     n380347 , n380348 , n380349 , n380350 , n380351 , n380352 , n380353 , n380354 , n380355 , n380356 , 
     n380357 , n380358 , n380359 , n380360 , n380361 , n380362 , n380363 , n380364 , n380365 , n380366 , 
     n380367 , n380368 , n380369 , n380370 , n380371 , n380372 , n380373 , n380374 , n380375 , n380376 , 
     n380377 , n380378 , n380379 , n380380 , n380381 , n380382 , n380383 , n380384 , n380385 , n380386 , 
     n380387 , n380388 , n380389 , n380390 , n380391 , n380392 , n380393 , n380394 , n380395 , n380396 , 
     n380397 , n380398 , n380399 , n380400 , n380401 , n380402 , n380403 , n380404 , n380405 , n380406 , 
     n380407 , n380408 , n380409 , n380410 , n380411 , n380412 , n380413 , n380414 , n380415 , n380416 , 
     n380417 , n380418 , n380419 , n380420 , n380421 , n380422 , n380423 , n380424 , n380425 , n380426 , 
     n380427 , n380428 , n380429 , n380430 , n380431 , n380432 , n380433 , n380434 , n380435 , n380436 , 
     n380437 , n380438 , n380439 , n380440 , n380441 , n380442 , n380443 , n380444 , n380445 , n380446 , 
     n380447 , n380448 , n380449 , n380450 , n380451 , n380452 , n380453 , n380454 , n380455 , n380456 , 
     n380457 , n380458 , n380459 , n380460 , n380461 , n380462 , n380463 , n380464 , n380465 , n380466 , 
     n380467 , n380468 , n380469 , n380470 , n380471 , n380472 , n380473 , n380474 , n380475 , n380476 , 
     n380477 , n380478 , n380479 , n380480 , n380481 , n380482 , n380483 , n380484 , n380485 , n380486 , 
     n380487 , n380488 , n380489 , n380490 , n380491 , n380492 , n380493 , n380494 , n380495 , n380496 , 
     n380497 , n380498 , n380499 , n380500 , n380501 , n380502 , n380503 , n380504 , n380505 , n380506 , 
     n380507 , n380508 , n380509 , n380510 , n380511 , n380512 , n380513 , n380514 , n380515 , n380516 , 
     n380517 , n380518 , n380519 , n380520 , n380521 , n380522 , n380523 , n380524 , n380525 , n380526 , 
     n380527 , n380528 , n380529 , n380530 , n380531 , n380532 , n380533 , n380534 , n380535 , n380536 , 
     n380537 , n380538 , n380539 , n380540 , n380541 , n380542 , n380543 , n380544 , n380545 , n380546 , 
     n380547 , n380548 , n380549 , n380550 , n380551 , n380552 , n380553 , n380554 , n380555 , n380556 , 
     n380557 , n380558 , n380559 , n380560 , n380561 , n380562 , n380563 , n380564 , n380565 , n380566 , 
     n380567 , n380568 , n380569 , n380570 , n380571 , n380572 , n380573 , n380574 , n380575 , n380576 , 
     n380577 , n380578 , n380579 , n380580 , n380581 , n380582 , n380583 , n380584 , n380585 , n380586 , 
     n380587 , n380588 , n380589 , n380590 , n380591 , n380592 , n380593 , n380594 , n380595 , n380596 , 
     n380597 , n380598 , n380599 , n380600 , n380601 , n380602 , n380603 , n380604 , n380605 , n380606 , 
     n380607 , n380608 , n380609 , n380610 , n380611 , n380612 , n380613 , n380614 , n380615 , n380616 , 
     n380617 , n380618 , n380619 , n380620 , n380621 , n380622 , n380623 , n380624 , n380625 , n380626 , 
     n380627 , n380628 , n380629 , n380630 , n380631 , n380632 , n380633 , n380634 , n380635 , n380636 , 
     n380637 , n380638 , n380639 , n380640 , n380641 , n380642 , n380643 , n380644 , n380645 , n380646 , 
     n380647 , n380648 , n380649 , n380650 , n380651 , n380652 , n380653 , n380654 , n380655 , n380656 , 
     n380657 , n380658 , n380659 , n380660 , n380661 , n380662 , n380663 , n380664 , n380665 , n380666 , 
     n380667 , n380668 , n380669 , n380670 , n380671 , n380672 , n380673 , n380674 , n380675 , n380676 , 
     n380677 , n380678 , n380679 , n380680 , n380681 , n380682 , n380683 , n380684 , n380685 , n380686 , 
     n380687 , n380688 , n380689 , n380690 , n380691 , n380692 , n380693 , n380694 , n380695 , n380696 , 
     n380697 , n380698 , n380699 , n380700 , n380701 , n380702 , n380703 , n380704 , n380705 , n380706 , 
     n380707 , n380708 , n380709 , n380710 , n380711 , n380712 , n380713 , n380714 , n380715 , n380716 , 
     n380717 , n380718 , n380719 , n380720 , n380721 , n380722 , n380723 , n380724 , n380725 , n380726 , 
     n380727 , n380728 , n380729 , n380730 , n380731 , n380732 , n380733 , n380734 , n380735 , n380736 , 
     n380737 , n380738 , n380739 , n380740 , n380741 , n380742 , n380743 , n380744 , n380745 , n380746 , 
     n380747 , n380748 , n380749 , n380750 , n380751 , n380752 , n380753 , n380754 , n380755 , n380756 , 
     n380757 , n380758 , n380759 , n380760 , n380761 , n380762 , n380763 , n380764 , n380765 , n380766 , 
     n380767 , n380768 , n380769 , n380770 , n380771 , n380772 , n380773 , n380774 , n380775 , n380776 , 
     n380777 , n380778 , n380779 , n380780 , n380781 , n380782 , n380783 , n380784 , n380785 , n380786 , 
     n380787 , n380788 , n380789 , n380790 , n380791 , n380792 , n380793 , n380794 , n380795 , n380796 , 
     n380797 , n380798 , n380799 , n380800 , n380801 , n380802 , n380803 , n380804 , n380805 , n380806 , 
     n380807 , n380808 , n380809 , n380810 , n380811 , n380812 , n380813 , n380814 , n380815 , n380816 , 
     n380817 , n380818 , n380819 , n380820 , n380821 , n380822 , n380823 , n380824 , n380825 , n380826 , 
     n380827 , n380828 , n380829 , n380830 , n380831 , n380832 , n380833 , n380834 , n380835 , n380836 , 
     n380837 , n380838 , n380839 , n380840 , n380841 , n380842 , n380843 , n380844 , n380845 , n380846 , 
     n380847 , n380848 , n380849 , n380850 , n380851 , n380852 , n380853 , n380854 , n380855 , n380856 , 
     n380857 , n380858 , n380859 , n380860 , n380861 , n380862 , n380863 , n380864 , n380865 , n380866 , 
     n380867 , n380868 , n380869 , n380870 , n380871 , n380872 , n380873 , n380874 , n380875 , n380876 , 
     n380877 , n380878 , n380879 , n380880 , n380881 , n380882 , n380883 , n380884 , n380885 , n380886 , 
     n380887 , n380888 , n380889 , n380890 , n380891 , n380892 , n380893 , n380894 , n380895 , n380896 , 
     n380897 , n380898 , n380899 , n380900 , n380901 , n380902 , n380903 , n380904 , n380905 , n380906 , 
     n380907 , n380908 , n380909 , n380910 , n380911 , n380912 , n380913 , n380914 , n380915 , n380916 , 
     n380917 , n380918 , n380919 , n380920 , n380921 , n380922 , n380923 , n380924 , n380925 , n380926 , 
     n380927 , n380928 , n380929 , n380930 , n380931 , n380932 , n380933 , n380934 , n380935 , n380936 , 
     n380937 , n380938 , n380939 , n380940 , n380941 , n380942 , n380943 , n380944 , n380945 , n380946 , 
     n380947 , n380948 , n380949 , n380950 , n380951 , n380952 , n380953 , n380954 , n380955 , n380956 , 
     n380957 , n380958 , n380959 , n380960 , n380961 , n380962 , n380963 , n380964 , n380965 , n380966 , 
     n380967 , n380968 , n380969 , n380970 , n380971 , n380972 , n380973 , n380974 , n380975 , n380976 , 
     n380977 , n380978 , n380979 , n380980 , n380981 , n380982 , n380983 , n380984 , n380985 , n380986 , 
     n380987 , n380988 , n380989 , n380990 , n380991 , n380992 , n380993 , n380994 , n380995 , n380996 , 
     n380997 , n380998 , n380999 , n381000 , n381001 , n381002 , n381003 , n381004 , n381005 , n381006 , 
     n381007 , n381008 , n381009 , n381010 , n381011 , n381012 , n381013 , n381014 , n381015 , n381016 , 
     n381017 , n381018 , n381019 , n381020 , n381021 , n381022 , n381023 , n381024 , n381025 , n381026 , 
     n381027 , n381028 , n381029 , n381030 , n381031 , n381032 , n381033 , n381034 , n381035 , n381036 , 
     n381037 , n381038 , n381039 , n381040 , n381041 , n381042 , n381043 , n381044 , n381045 , n381046 , 
     n381047 , n381048 , n381049 , n381050 , n381051 , n381052 , n381053 , n381054 , n381055 , n381056 , 
     n381057 , n381058 , n381059 , n381060 , n381061 , n381062 , n381063 , n381064 , n381065 , n381066 , 
     n381067 , n381068 , n381069 , n381070 , n381071 , n381072 , n381073 , n381074 , n381075 , n381076 , 
     n381077 , n381078 , n381079 , n381080 , n381081 , n381082 , n381083 , n381084 , n381085 , n381086 , 
     n381087 , n381088 , n381089 , n381090 , n381091 , n381092 , n381093 , n381094 , n381095 , n381096 , 
     n381097 , n381098 , n381099 , n381100 , n381101 , n381102 , n381103 , n381104 , n381105 , n381106 , 
     n381107 , n381108 , n381109 , n381110 , n381111 , n381112 , n381113 , n381114 , n381115 , n381116 , 
     n381117 , n381118 , n381119 , n381120 , n381121 , n381122 , n381123 , n381124 , n381125 , n381126 , 
     n381127 , n381128 , n381129 , n381130 , n381131 , n381132 , n381133 , n381134 , n381135 , n381136 , 
     n381137 , n381138 , n381139 , n381140 , n381141 , n381142 , n381143 , n381144 , n381145 , n381146 , 
     n381147 , n381148 , n381149 , n381150 , n381151 , n381152 , n381153 , n381154 , n381155 , n381156 , 
     n381157 , n381158 , n381159 , n381160 , n381161 , n381162 , n381163 , n381164 , n381165 , n381166 , 
     n381167 , n381168 , n381169 , n381170 , n381171 , n381172 , n381173 , n381174 , n381175 , n381176 , 
     n381177 , n381178 , n381179 , n381180 , n381181 , n381182 , n381183 , n381184 , n381185 , n381186 , 
     n381187 , n381188 , n381189 , n381190 , n381191 , n381192 , n381193 , n381194 , n381195 , n381196 , 
     n381197 , n381198 , n381199 , n381200 , n381201 , n381202 , n381203 , n381204 , n381205 , n381206 , 
     n381207 , n381208 , n381209 , n381210 , n381211 , n381212 , n381213 , n381214 , n381215 , n381216 , 
     n381217 , n381218 , n381219 , n381220 , n381221 , n381222 , n381223 , n381224 , n381225 , n381226 , 
     n381227 , n381228 , n381229 , n381230 , n381231 , n381232 , n381233 , n381234 , n381235 , n381236 , 
     n381237 , n381238 , n381239 , n381240 , n381241 , n381242 , n381243 , n381244 , n381245 , n381246 , 
     n381247 , n381248 , n381249 , n381250 , n381251 , n381252 , n381253 , n381254 , n381255 , n381256 , 
     n381257 , n381258 , n381259 , n381260 , n381261 , n381262 , n381263 , n381264 , n381265 , n381266 , 
     n381267 , n381268 , n381269 , n381270 , n381271 , n381272 , n381273 , n381274 , n381275 , n381276 , 
     n381277 , n381278 , n381279 , n381280 , n381281 , n381282 , n381283 , n381284 , n381285 , n381286 , 
     n381287 , n381288 , n381289 , n381290 , n381291 , n381292 , n381293 , n381294 , n381295 , n381296 , 
     n381297 , n381298 , n381299 , n381300 , n381301 , n381302 , n381303 , n381304 , n381305 , n381306 , 
     n381307 , n381308 , n381309 , n381310 , n381311 , n381312 , n381313 , n381314 , n381315 , n381316 , 
     n381317 , n381318 , n381319 , n381320 , n381321 , n381322 , n381323 , n381324 , n381325 , n381326 , 
     n381327 , n381328 , n381329 , n381330 , n381331 , n381332 , n381333 , n381334 , n381335 , n381336 , 
     n381337 , n381338 , n381339 , n381340 , n381341 , n381342 , n381343 , n381344 , n381345 , n381346 , 
     n381347 , n381348 , n381349 , n381350 , n381351 , n381352 , n381353 , n381354 , n381355 , n381356 , 
     n381357 , n381358 , n381359 , n381360 , n381361 , n381362 , n381363 , n381364 , n381365 , n381366 , 
     n381367 , n381368 , n381369 , n381370 , n381371 , n381372 , n381373 , n381374 , n381375 , n381376 , 
     n381377 , n381378 , n381379 , n381380 , n381381 , n381382 , n381383 , n381384 , n381385 , n381386 , 
     n381387 , n381388 , n381389 , n381390 , n381391 , n381392 , n381393 , n381394 , n381395 , n381396 , 
     n381397 , n381398 , n381399 , n381400 , n381401 , n381402 , n381403 , n381404 , n381405 , n381406 , 
     n381407 , n381408 , n381409 , n381410 , n381411 , n381412 , n381413 , n381414 , n381415 , n381416 , 
     n381417 , n381418 , n381419 , n381420 , n381421 , n381422 , n381423 , n381424 , n381425 , n381426 , 
     n381427 , n381428 , n381429 , n381430 , n381431 , n381432 , n381433 , n381434 , n381435 , n381436 , 
     n381437 , n381438 , n381439 , n381440 , n381441 , n381442 , n381443 , n381444 , n381445 , n381446 , 
     n381447 , n381448 , n381449 , n381450 , n381451 , n381452 , n381453 , n381454 , n381455 , n381456 , 
     n381457 , n381458 , n381459 , n381460 , n381461 , n381462 , n381463 , n381464 , n381465 , n381466 , 
     n381467 , n381468 , n381469 , n381470 , n381471 , n381472 , n381473 , n381474 , n381475 , n381476 , 
     n381477 , n381478 , n381479 , n381480 , n381481 , n381482 , n381483 , n381484 , n381485 , n381486 , 
     n381487 , n381488 , n381489 , n381490 , n381491 , n381492 , n381493 , n381494 , n381495 , n381496 , 
     n381497 , n381498 , n381499 , n381500 , n381501 , n381502 , n381503 , n381504 , n381505 , n381506 , 
     n381507 , n381508 , n381509 , n381510 , n381511 , n381512 , n381513 , n381514 , n381515 , n381516 , 
     n381517 , n381518 , n381519 , n381520 , n381521 , n381522 , n381523 , n381524 , n381525 , n381526 , 
     n381527 , n381528 , n381529 , n381530 , n381531 , n381532 , n381533 , n381534 , n381535 , n381536 , 
     n381537 , n381538 , n381539 , n381540 , n381541 , n381542 , n381543 , n381544 , n381545 , n381546 , 
     n381547 , n381548 , n381549 , n381550 , n381551 , n381552 , n381553 , n381554 , n381555 , n381556 , 
     n381557 , n381558 , n381559 , n381560 , n381561 , n381562 , n381563 , n381564 , n381565 , n381566 , 
     n381567 , n381568 , n381569 , n381570 , n381571 , n381572 , n381573 , n381574 , n381575 , n381576 , 
     n381577 , n381578 , n381579 , n381580 , n381581 , n381582 , n381583 , n381584 , n381585 , n381586 , 
     n381587 , n381588 , n381589 , n381590 , n381591 , n381592 , n381593 , n381594 , n381595 , n381596 , 
     n381597 , n381598 , n381599 , n381600 , n381601 , n381602 , n381603 , n381604 , n381605 , n381606 , 
     n381607 , n381608 , n381609 , n381610 , n381611 , n381612 , n381613 , n381614 , n381615 , n381616 , 
     n381617 , n381618 , n381619 , n381620 , n381621 , n381622 , n381623 , n381624 , n381625 , n381626 , 
     n381627 , n381628 , n381629 , n381630 , n381631 , n381632 , n381633 , n381634 , n381635 , n381636 , 
     n381637 , n381638 , n381639 , n381640 , n381641 , n381642 , n381643 , n381644 , n381645 , n381646 , 
     n381647 , n381648 , n381649 , n381650 , n381651 , n381652 , n381653 , n381654 , n381655 , n381656 , 
     n381657 , n381658 , n381659 , n381660 , n381661 , n381662 , n381663 , n381664 , n381665 , n381666 , 
     n381667 , n381668 , n381669 , n381670 , n381671 , n381672 , n381673 , n381674 , n381675 , n381676 , 
     n381677 , n381678 , n381679 , n381680 , n381681 , n381682 , n381683 , n381684 , n381685 , n381686 , 
     n381687 , n381688 , n381689 , n381690 , n381691 , n381692 , n381693 , n381694 , n381695 , n381696 , 
     n381697 , n381698 , n381699 , n381700 , n381701 , n381702 , n381703 , n381704 , n381705 , n381706 , 
     n381707 , n381708 , n381709 , n381710 , n381711 , n381712 , n381713 , n381714 , n381715 , n381716 , 
     n381717 , n381718 , n381719 , n381720 , n381721 , n381722 , n381723 , n381724 , n381725 , n381726 , 
     n381727 , n381728 , n381729 , n381730 , n381731 , n381732 , n381733 , n381734 , n381735 , n381736 , 
     n381737 , n381738 , n381739 , n381740 , n381741 , n381742 , n381743 , n381744 , n381745 , n381746 , 
     n381747 , n381748 , n381749 , n381750 , n381751 , n381752 , n381753 , n381754 , n381755 , n381756 , 
     n381757 , n381758 , n381759 , n381760 , n381761 , n381762 , n381763 , n381764 , n381765 , n381766 , 
     n381767 , n381768 , n381769 , n381770 , n381771 , n381772 , n381773 , n381774 , n381775 , n381776 , 
     n381777 , n381778 , n381779 , n381780 , n381781 , n381782 , n381783 , n381784 , n381785 , n381786 , 
     n381787 , n381788 , n381789 , n381790 , n381791 , n381792 , n381793 , n381794 , n381795 , n381796 , 
     n381797 , n381798 , n381799 , n381800 , n381801 , n381802 , n381803 , n381804 , n381805 , n381806 , 
     n381807 , n381808 , n381809 , n381810 , n381811 , n381812 , n381813 , n381814 , n381815 , n381816 , 
     n381817 , n381818 , n381819 , n381820 , n381821 , n381822 , n381823 , n381824 , n381825 , n381826 , 
     n381827 , n381828 , n381829 , n381830 , n381831 , n381832 , n381833 , n381834 , n381835 , n381836 , 
     n381837 , n381838 , n381839 , n381840 , n381841 , n381842 , n381843 , n381844 , n381845 , n381846 , 
     n381847 , n381848 , n381849 , n381850 , n381851 , n381852 , n381853 , n381854 , n381855 , n381856 , 
     n381857 , n381858 , n381859 , n381860 , n381861 , n381862 , n381863 , n381864 , n381865 , n381866 , 
     n381867 , n381868 , n381869 , n381870 , n381871 , n381872 , n381873 , n381874 , n381875 , n381876 , 
     n381877 , n381878 , n381879 , n381880 , n381881 , n381882 , n381883 , n381884 , n381885 , n381886 , 
     n381887 , n381888 , n381889 , n381890 , n381891 , n381892 , n381893 , n381894 , n381895 , n381896 , 
     n381897 , n381898 , n381899 , n381900 , n381901 , n381902 , n381903 , n381904 , n381905 , n381906 , 
     n381907 , n381908 , n381909 , n381910 , n381911 , n381912 , n381913 , n381914 , n381915 , n381916 , 
     n381917 , n381918 , n381919 , n381920 , n381921 , n381922 , n381923 , n381924 , n381925 , n381926 , 
     n381927 , n381928 , n381929 , n381930 , n381931 , n381932 , n381933 , n381934 , n381935 , n381936 , 
     n381937 , n381938 , n381939 , n381940 , n381941 , n381942 , n381943 , n381944 , n381945 , n381946 , 
     n381947 , n381948 , n381949 , n381950 , n381951 , n381952 , n381953 , n381954 , n381955 , n381956 , 
     n381957 , n381958 , n381959 , n381960 , n381961 , n381962 , n381963 , n381964 , n381965 , n381966 , 
     n381967 , n381968 , n381969 , n381970 , n381971 , n381972 , n381973 , n381974 , n381975 , n381976 , 
     n381977 , n381978 , n381979 , n381980 , n381981 , n381982 , n381983 , n381984 , n381985 , n381986 , 
     n381987 , n381988 , n381989 , n381990 , n381991 , n381992 , n381993 , n381994 , n381995 , n381996 , 
     n381997 , n381998 , n381999 , n382000 , n382001 , n382002 , n382003 , n382004 , n382005 , n382006 , 
     n382007 , n382008 , n382009 , n382010 , n382011 , n382012 , n382013 , n382014 , n382015 , n382016 , 
     n382017 , n382018 , n382019 , n382020 , n382021 , n382022 , n382023 , n382024 , n382025 , n382026 , 
     n382027 , n382028 , n382029 , n382030 , n382031 , n382032 , n382033 , n382034 , n382035 , n382036 , 
     n382037 , n382038 , n382039 , n382040 , n382041 , n382042 , n382043 , n382044 , n382045 , n382046 , 
     n382047 , n382048 , n382049 , n382050 , n382051 , n382052 , n382053 , n382054 , n382055 , n382056 , 
     n382057 , n382058 , n382059 , n382060 , n382061 , n382062 , n382063 , n382064 , n382065 , n382066 , 
     n382067 , n382068 , n382069 , n382070 , n382071 , n382072 , n382073 , n382074 , n382075 , n382076 , 
     n382077 , n382078 , n382079 , n382080 , n382081 , n382082 , n382083 , n382084 , n382085 , n382086 , 
     n382087 , n382088 , n382089 , n382090 , n382091 , n382092 , n382093 , n382094 , n382095 , n382096 , 
     n382097 , n382098 , n382099 , n382100 , n382101 , n382102 , n382103 , n382104 , n382105 , n382106 , 
     n382107 , n382108 , n382109 , n382110 , n382111 , n382112 , n382113 , n382114 , n382115 , n382116 , 
     n382117 , n382118 , n382119 , n382120 , n382121 , n382122 , n382123 , n382124 , n382125 , n382126 , 
     n382127 , n382128 , n382129 , n382130 , n382131 , n382132 , n382133 , n382134 , n382135 , n382136 , 
     n382137 , n382138 , n382139 , n382140 , n382141 , n382142 , n382143 , n382144 , n382145 , n382146 , 
     n382147 , n382148 , n382149 , n382150 , n382151 , n382152 , n382153 , n382154 , n382155 , n382156 , 
     n382157 , n382158 , n382159 , n382160 , n382161 , n382162 , n382163 , n382164 , n382165 , n382166 , 
     n382167 , n382168 , n382169 , n382170 , n382171 , n382172 , n382173 , n382174 , n382175 , n382176 , 
     n382177 , n382178 , n382179 , n382180 , n382181 , n382182 , n382183 , n382184 , n382185 , n382186 , 
     n382187 , n382188 , n382189 , n382190 , n382191 , n382192 , n382193 , n382194 , n382195 , n382196 , 
     n382197 , n382198 , n382199 , n382200 , n382201 , n382202 , n382203 , n382204 , n382205 , n382206 , 
     n382207 , n382208 , n382209 , n382210 , n382211 , n382212 , n382213 , n382214 , n382215 , n382216 , 
     n382217 , n382218 , n382219 , n382220 , n382221 , n382222 , n382223 , n382224 , n382225 , n382226 , 
     n382227 , n382228 , n382229 , n382230 , n382231 , n382232 , n382233 , n382234 , n382235 , n382236 , 
     n382237 , n382238 , n382239 , n382240 , n382241 , n382242 , n382243 , n382244 , n382245 , n382246 , 
     n382247 , n382248 , n382249 , n382250 , n382251 , n382252 , n382253 , n382254 , n382255 , n382256 , 
     n382257 , n382258 , n382259 , n382260 , n382261 , n382262 , n382263 , n382264 , n382265 , n382266 , 
     n382267 , n382268 , n382269 , n382270 , n382271 , n382272 , n382273 , n382274 , n382275 , n382276 , 
     n382277 , n382278 , n382279 , n382280 , n382281 , n382282 , n382283 , n382284 , n382285 , n382286 , 
     n382287 , n382288 , n382289 , n382290 , n382291 , n382292 , n382293 , n382294 , n382295 , n382296 , 
     n382297 , n382298 , n382299 , n382300 , n382301 , n382302 , n382303 , n382304 , n382305 , n382306 , 
     n382307 , n382308 , n382309 , n382310 , n382311 , n382312 , n382313 , n382314 , n382315 , n382316 , 
     n382317 , n382318 , n382319 , n382320 , n382321 , n382322 , n382323 , n382324 , n382325 , n382326 , 
     n382327 , n382328 , n382329 , n382330 , n382331 , n382332 , n382333 , n382334 , n382335 , n382336 , 
     n382337 , n382338 , n382339 , n382340 , n382341 , n382342 , n382343 , n382344 , n382345 , n382346 , 
     n382347 , n382348 , n382349 , n382350 , n382351 , n382352 , n382353 , n382354 , n382355 , n382356 , 
     n382357 , n382358 , n382359 , n382360 , n382361 , n382362 , n382363 , n382364 , n382365 , n382366 , 
     n382367 , n382368 , n382369 , n382370 , n382371 , n382372 , n382373 , n382374 , n382375 , n382376 , 
     n382377 , n382378 , n382379 , n382380 , n382381 , n382382 , n382383 , n382384 , n382385 , n382386 , 
     n382387 , n382388 , n382389 , n382390 , n382391 , n382392 , n382393 , n382394 , n382395 , n382396 , 
     n382397 , n382398 , n382399 , n382400 , n382401 , n382402 , n382403 , n382404 , n382405 , n382406 , 
     n382407 , n382408 , n382409 , n382410 , n382411 , n382412 , n382413 , n382414 , n382415 , n382416 , 
     n382417 , n382418 , n382419 , n382420 , n382421 , n382422 , n382423 , n382424 , n382425 , n382426 , 
     n382427 , n382428 , n382429 , n382430 , n382431 , n382432 , n382433 , n382434 , n382435 , n382436 , 
     n382437 , n382438 , n382439 , n382440 , n382441 , n382442 , n382443 , n382444 , n382445 , n382446 , 
     n382447 , n382448 , n382449 , n382450 , n382451 , n382452 , n382453 , n382454 , n382455 , n382456 , 
     n382457 , n382458 , n382459 , n382460 , n382461 , n382462 , n382463 , n382464 , n382465 , n382466 , 
     n382467 , n382468 , n382469 , n382470 , n382471 , n382472 , n382473 , n382474 , n382475 , n382476 , 
     n382477 , n382478 , n382479 , n382480 , n382481 , n382482 , n382483 , n382484 , n382485 , n382486 , 
     n382487 , n382488 , n382489 , n382490 , n382491 , n382492 , n382493 , n382494 , n382495 , n382496 , 
     n382497 , n382498 , n382499 , n382500 , n382501 , n382502 , n382503 , n382504 , n382505 , n382506 , 
     n382507 , n382508 , n382509 , n382510 , n382511 , n382512 , n382513 , n382514 , n382515 , n382516 , 
     n382517 , n382518 , n382519 , n382520 , n382521 , n382522 , n382523 , n382524 , n382525 , n382526 , 
     n382527 , n382528 , n382529 , n382530 , n382531 , n382532 , n382533 , n382534 , n382535 , n382536 , 
     n382537 , n382538 , n382539 , n382540 , n382541 , n382542 , n382543 , n382544 , n382545 , n382546 , 
     n382547 , n382548 , n382549 , n382550 , n382551 , n382552 , n382553 , n382554 , n382555 , n382556 , 
     n382557 , n382558 , n382559 , n382560 , n382561 , n382562 , n382563 , n382564 , n382565 , n382566 , 
     n382567 , n382568 , n382569 , n382570 , n382571 , n382572 , n382573 , n382574 , n382575 , n382576 , 
     n382577 , n382578 , n382579 , n382580 , n382581 , n382582 , n382583 , n382584 , n382585 , n382586 , 
     n382587 , n382588 , n382589 , n382590 , n382591 , n382592 , n382593 , n382594 , n382595 , n382596 , 
     n382597 , n382598 , n382599 , n382600 , n382601 , n382602 , n382603 , n382604 , n382605 , n382606 , 
     n382607 , n382608 , n382609 , n382610 , n382611 , n382612 , n382613 , n382614 , n382615 , n382616 , 
     n382617 , n382618 , n382619 , n382620 , n382621 , n382622 , n382623 , n382624 , n382625 , n382626 , 
     n382627 , n382628 , n382629 , n382630 , n382631 , n382632 , n382633 , n382634 , n382635 , n382636 , 
     n382637 , n382638 , n382639 , n382640 , n382641 , n382642 , n382643 , n382644 , n382645 , n382646 , 
     n382647 , n382648 , n382649 , n382650 , n382651 , n382652 , n382653 , n382654 , n382655 , n382656 , 
     n382657 , n382658 , n382659 , n382660 , n382661 , n382662 , n382663 , n382664 , n382665 , n382666 , 
     n382667 , n382668 , n382669 , n382670 , n382671 , n382672 , n382673 , n382674 , n382675 , n382676 , 
     n382677 , n382678 , n382679 , n382680 , n382681 , n382682 , n382683 , n382684 , n382685 , n382686 , 
     n382687 , n382688 , n382689 , n382690 , n382691 , n382692 , n382693 , n382694 , n382695 , n382696 , 
     n382697 , n382698 , n382699 , n382700 , n382701 , n382702 , n382703 , n382704 , n382705 , n382706 , 
     n382707 , n382708 , n382709 , n382710 , n382711 , n382712 , n382713 , n382714 , n382715 , n382716 , 
     n382717 , n382718 , n382719 , n382720 , n382721 , n382722 , n382723 , n382724 , n382725 , n382726 , 
     n382727 , n382728 , n382729 , n382730 , n382731 , n382732 , n382733 , n382734 , n382735 , n382736 , 
     n382737 , n382738 , n382739 , n382740 , n382741 , n382742 , n382743 , n382744 , n382745 , n382746 , 
     n382747 , n382748 , n382749 , n382750 , n382751 , n382752 , n382753 , n382754 , n382755 , n382756 , 
     n382757 , n382758 , n382759 , n382760 , n382761 , n382762 , n382763 , n382764 , n382765 , n382766 , 
     n382767 , n382768 , n382769 , n382770 , n382771 , n382772 , n382773 , n382774 , n382775 , n382776 , 
     n382777 , n382778 , n382779 , n382780 , n382781 , n382782 , n382783 , n382784 , n382785 , n382786 , 
     n382787 , n382788 , n382789 , n382790 , n382791 , n382792 , n382793 , n382794 , n382795 , n382796 , 
     n382797 , n382798 , n382799 , n382800 , n382801 , n382802 , n382803 , n382804 , n382805 , n382806 , 
     n382807 , n382808 , n382809 , n382810 , n382811 , n382812 , n382813 , n382814 , n382815 , n382816 , 
     n382817 , n382818 , n382819 , n382820 , n382821 , n382822 , n382823 , n382824 , n382825 , n382826 , 
     n382827 , n382828 , n382829 , n382830 , n382831 , n382832 , n382833 , n382834 , n382835 , n382836 , 
     n382837 , n382838 , n382839 , n382840 , n382841 , n382842 , n382843 , n382844 , n382845 , n382846 , 
     n382847 , n382848 , n382849 , n382850 , n382851 , n382852 , n382853 , n382854 , n382855 , n382856 , 
     n382857 , n382858 , n382859 , n382860 , n382861 , n382862 , n382863 , n382864 , n382865 , n382866 , 
     n382867 , n382868 , n382869 , n382870 , n382871 , n382872 , n382873 , n382874 , n382875 , n382876 , 
     n382877 , n382878 , n382879 , n382880 , n382881 , n382882 , n382883 , n382884 , n382885 , n382886 , 
     n382887 , n382888 , n382889 , n382890 , n382891 , n382892 , n382893 , n382894 , n382895 , n382896 , 
     n382897 , n382898 , n382899 , n382900 , n382901 , n382902 , n382903 , n382904 , n382905 , n382906 , 
     n382907 , n382908 , n382909 , n382910 , n382911 , n382912 , n382913 , n382914 , n382915 , n382916 , 
     n382917 , n382918 , n382919 , n382920 , n382921 , n382922 , n382923 , n382924 , n382925 , n382926 , 
     n382927 , n382928 , n382929 , n382930 , n382931 , n382932 , n382933 , n382934 , n382935 , n382936 , 
     n382937 , n382938 , n382939 , n382940 , n382941 , n382942 , n382943 , n382944 , n382945 , n382946 , 
     n382947 , n382948 , n382949 , n382950 , n382951 , n382952 , n382953 , n382954 , n382955 , n382956 , 
     n382957 , n382958 , n382959 , n382960 , n382961 , n382962 , n382963 , n382964 , n382965 , n382966 , 
     n382967 , n382968 , n382969 , n382970 , n382971 , n382972 , n382973 , n382974 , n382975 , n382976 , 
     n382977 , n382978 , n382979 , n382980 , n382981 , n382982 , n382983 , n382984 , n382985 , n382986 , 
     n382987 , n382988 , n382989 , n382990 , n382991 , n382992 , n382993 , n382994 , n382995 , n382996 , 
     n382997 , n382998 , n382999 , n383000 , n383001 , n383002 , n383003 , n383004 , n383005 , n383006 , 
     n383007 , n383008 , n383009 , n383010 , n383011 , n383012 , n383013 , n383014 , n383015 , n383016 , 
     n383017 , n383018 , n383019 , n383020 , n383021 , n383022 , n383023 , n383024 , n383025 , n383026 , 
     n383027 , n383028 , n383029 , n383030 , n383031 , n383032 , n383033 , n383034 , n383035 , n383036 , 
     n383037 , n383038 , n383039 , n383040 , n383041 , n383042 , n383043 , n383044 , n383045 , n383046 , 
     n383047 , n383048 , n383049 , n383050 , n383051 , n383052 , n383053 , n383054 , n383055 , n383056 , 
     n383057 , n383058 , n383059 , n383060 , n383061 , n383062 , n383063 , n383064 , n383065 , n383066 , 
     n383067 , n383068 , n383069 , n383070 , n383071 , n383072 , n383073 , n383074 , n383075 , n383076 , 
     n383077 , n383078 , n383079 , n383080 , n383081 , n383082 , n383083 , n383084 , n383085 , n383086 , 
     n383087 , n383088 , n383089 , n383090 , n383091 , n383092 , n383093 , n383094 , n383095 , n383096 , 
     n383097 , n383098 , n383099 , n383100 , n383101 , n383102 , n383103 , n383104 , n383105 , n383106 , 
     n383107 , n383108 , n383109 , n383110 , n383111 , n383112 , n383113 , n383114 , n383115 , n383116 , 
     n383117 , n383118 , n383119 , n383120 , n383121 , n383122 , n383123 , n383124 , n383125 , n383126 , 
     n383127 , n383128 , n383129 , n383130 , n383131 , n383132 , n383133 , n383134 , n383135 , n383136 , 
     n383137 , n383138 , n383139 , n383140 , n383141 , n383142 , n383143 , n383144 , n383145 , n383146 , 
     n383147 , n383148 , n383149 , n383150 , n383151 , n383152 , n383153 , n383154 , n383155 , n383156 , 
     n383157 , n383158 , n383159 , n383160 , n383161 , n383162 , n383163 , n383164 , n383165 , n383166 , 
     n383167 , n383168 , n383169 , n383170 , n383171 , n383172 , n383173 , n383174 , n383175 , n383176 , 
     n383177 , n383178 , n383179 , n383180 , n383181 , n383182 , n383183 , n383184 , n383185 , n383186 , 
     n383187 , n383188 , n383189 , n383190 , n383191 , n383192 , n383193 , n383194 , n383195 , n383196 , 
     n383197 , n383198 , n383199 , n383200 , n383201 , n383202 , n383203 , n383204 , n383205 , n383206 , 
     n383207 , n383208 , n383209 , n383210 , n383211 , n383212 , n383213 , n383214 , n383215 , n383216 , 
     n383217 , n383218 , n383219 , n383220 , n383221 , n383222 , n383223 , n383224 , n383225 , n383226 , 
     n383227 , n383228 , n383229 , n383230 , n383231 , n383232 , n383233 , n383234 , n383235 , n383236 , 
     n383237 , n383238 , n383239 , n383240 , n383241 , n383242 , n383243 , n383244 , n383245 , n383246 , 
     n383247 , n383248 , n383249 , n383250 , n383251 , n383252 , n383253 , n383254 , n383255 , n383256 , 
     n383257 , n383258 , n383259 , n383260 , n383261 , n383262 , n383263 , n383264 , n383265 , n383266 , 
     n383267 , n383268 , n383269 , n383270 , n383271 , n383272 , n383273 , n383274 , n383275 , n383276 , 
     n383277 , n383278 , n383279 , n383280 , n383281 , n383282 , n383283 , n383284 , n383285 , n383286 , 
     n383287 , n383288 , n383289 , n383290 , n383291 , n383292 , n383293 , n383294 , n383295 , n383296 , 
     n383297 , n383298 , n383299 , n383300 , n383301 , n383302 , n383303 , n383304 , n383305 , n383306 , 
     n383307 , n383308 , n383309 , n383310 , n383311 , n383312 , n383313 , n383314 , n383315 , n383316 , 
     n383317 , n383318 , n383319 , n383320 , n383321 , n383322 , n383323 , n383324 , n383325 , n383326 , 
     n383327 , n383328 , n383329 , n383330 , n383331 , n383332 , n383333 , n383334 , n383335 , n383336 , 
     n383337 , n383338 , n383339 , n383340 , n383341 , n383342 , n383343 , n383344 , n383345 , n383346 , 
     n383347 , n383348 , n383349 , n383350 , n383351 , n383352 , n383353 , n383354 , n383355 , n383356 , 
     n383357 , n383358 , n383359 , n383360 , n383361 , n383362 , n383363 , n383364 , n383365 , n383366 , 
     n383367 , n383368 , n383369 , n383370 , n383371 , n383372 , n383373 , n383374 , n383375 , n383376 , 
     n383377 , n383378 , n383379 , n383380 , n383381 , n383382 , n383383 , n383384 , n383385 , n383386 , 
     n383387 , n383388 , n383389 , n383390 , n383391 , n383392 , n383393 , n383394 , n383395 , n383396 , 
     n383397 , n383398 , n383399 , n383400 , n383401 , n383402 , n383403 , n383404 , n383405 , n383406 , 
     n383407 , n383408 , n383409 , n383410 , n383411 , n383412 , n383413 , n383414 , n383415 , n383416 , 
     n383417 , n383418 , n383419 , n383420 , n383421 , n383422 , n383423 , n383424 , n383425 , n383426 , 
     n383427 , n383428 , n383429 , n383430 , n383431 , n383432 , n383433 , n383434 , n383435 , n383436 , 
     n383437 , n383438 , n383439 , n383440 , n383441 , n383442 , n383443 , n383444 , n383445 , n383446 , 
     n383447 , n383448 , n383449 , n383450 , n383451 , n383452 , n383453 , n383454 , n383455 , n383456 , 
     n383457 , n383458 , n383459 , n383460 , n383461 , n383462 , n383463 , n383464 , n383465 , n383466 , 
     n383467 , n383468 , n383469 , n383470 , n383471 , n383472 , n383473 , n383474 , n383475 , n383476 , 
     n383477 , n383478 , n383479 , n383480 , n383481 , n383482 , n383483 , n383484 , n383485 , n383486 , 
     n383487 , n383488 , n383489 , n383490 , n383491 , n383492 , n383493 , n383494 , n383495 , n383496 , 
     n383497 , n383498 , n383499 , n383500 , n383501 , n383502 , n383503 , n383504 , n383505 , n383506 , 
     n383507 , n383508 , n383509 , n383510 , n383511 , n383512 , n383513 , n383514 , n383515 , n383516 , 
     n383517 , n383518 , n383519 , n383520 , n383521 , n383522 , n383523 , n383524 , n383525 , n383526 , 
     n383527 , n383528 , n383529 , n383530 , n383531 , n383532 , n383533 , n383534 , n383535 , n383536 , 
     n383537 , n383538 , n383539 , n383540 , n383541 , n383542 , n383543 , n383544 , n383545 , n383546 , 
     n383547 , n383548 , n383549 , n383550 , n383551 , n383552 , n383553 , n383554 , n383555 , n383556 , 
     n383557 , n383558 , n383559 , n383560 , n383561 , n383562 , n383563 , n383564 , n383565 , n383566 , 
     n383567 , n383568 , n383569 , n383570 , n383571 , n383572 , n383573 , n383574 , n383575 , n383576 , 
     n383577 , n383578 , n383579 , n383580 , n383581 , n383582 , n383583 , n383584 , n383585 , n383586 , 
     n383587 , n383588 , n383589 , n383590 , n383591 , n383592 , n383593 , n383594 , n383595 , n383596 , 
     n383597 , n383598 , n383599 , n383600 , n383601 , n383602 , n383603 , n383604 , n383605 , n383606 , 
     n383607 , n383608 , n383609 , n383610 , n383611 , n383612 , n383613 , n383614 , n383615 , n383616 , 
     n383617 , n383618 , n383619 , n383620 , n383621 , n383622 , n383623 , n383624 , n383625 , n383626 , 
     n383627 , n383628 , n383629 , n383630 , n383631 , n383632 , n383633 , n383634 , n383635 , n383636 , 
     n383637 , n383638 , n383639 , n383640 , n383641 , n383642 , n383643 , n383644 , n383645 , n383646 , 
     n383647 , n383648 , n383649 , n383650 , n383651 , n383652 , n383653 , n383654 , n383655 , n383656 , 
     n383657 , n383658 , n383659 , n383660 , n383661 , n383662 , n383663 , n383664 , n383665 , n383666 , 
     n383667 , n383668 , n383669 , n383670 , n383671 , n383672 , n383673 , n383674 , n383675 , n383676 , 
     n383677 , n383678 , n383679 , n383680 , n383681 , n383682 , n383683 , n383684 , n383685 , n383686 , 
     n383687 , n383688 , n383689 , n383690 , n383691 , n383692 , n383693 , n383694 , n383695 , n383696 , 
     n383697 , n383698 , n383699 , n383700 , n383701 , n383702 , n383703 , n383704 , n383705 , n383706 , 
     n383707 , n383708 , n383709 , n383710 , n383711 , n383712 , n383713 , n383714 , n383715 , n383716 , 
     n383717 , n383718 , n383719 , n383720 , n383721 , n383722 , n383723 , n383724 , n383725 , n383726 , 
     n383727 , n383728 , n383729 , n383730 , n383731 , n383732 , n383733 , n383734 , n383735 , n383736 , 
     n383737 , n383738 , n383739 , n383740 , n383741 , n383742 , n383743 , n383744 , n383745 , n383746 , 
     n383747 , n383748 , n383749 , n383750 , n383751 , n383752 , n383753 , n383754 , n383755 , n383756 , 
     n383757 , n383758 , n383759 , n383760 , n383761 , n383762 , n383763 , n383764 , n383765 , n383766 , 
     n383767 , n383768 , n383769 , n383770 , n383771 , n383772 , n383773 , n383774 , n383775 , n383776 , 
     n383777 , n383778 , n383779 , n383780 , n383781 , n383782 , n383783 , n383784 , n383785 , n383786 , 
     n383787 , n383788 , n383789 , n383790 , n383791 , n383792 , n383793 , n383794 , n383795 , n383796 , 
     n383797 , n383798 , n383799 , n383800 , n383801 , n383802 , n383803 , n383804 , n383805 , n383806 , 
     n383807 , n383808 , n383809 , n383810 , n383811 , n383812 , n383813 , n383814 , n383815 , n383816 , 
     n383817 , n383818 , n383819 , n383820 , n383821 , n383822 , n383823 , n383824 , n383825 , n383826 , 
     n383827 , n383828 , n383829 , n383830 , n383831 , n383832 , n383833 , n383834 , n383835 , n383836 , 
     n383837 , n383838 , n383839 , n383840 , n383841 , n383842 , n383843 , n383844 , n383845 , n383846 , 
     n383847 , n383848 , n383849 , n383850 , n383851 , n383852 , n383853 , n383854 , n383855 , n383856 , 
     n383857 , n383858 , n383859 , n383860 , n383861 , n383862 , n383863 , n383864 , n383865 , n383866 , 
     n383867 , n383868 , n383869 , n383870 , n383871 , n383872 , n383873 , n383874 , n383875 , n383876 , 
     n383877 , n383878 , n383879 , n383880 , n383881 , n383882 , n383883 , n383884 , n383885 , n383886 , 
     n383887 , n383888 , n383889 , n383890 , n383891 , n383892 , n383893 , n383894 , n383895 , n383896 , 
     n383897 , n383898 , n383899 , n383900 , n383901 , n383902 , n383903 , n383904 , n383905 , n383906 , 
     n383907 , n383908 , n383909 , n383910 , n383911 , n383912 , n383913 , n383914 , n383915 , n383916 , 
     n383917 , n383918 , n383919 , n383920 , n383921 , n383922 , n383923 , n383924 , n383925 , n383926 , 
     n383927 , n383928 , n383929 , n383930 , n383931 , n383932 , n383933 , n383934 , n383935 , n383936 , 
     n383937 , n383938 , n383939 , n383940 , n383941 , n383942 , n383943 , n383944 , n383945 , n383946 , 
     n383947 , n383948 , n383949 , n383950 , n383951 , n383952 , n383953 , n383954 , n383955 , n383956 , 
     n383957 , n383958 , n383959 , n383960 , n383961 , n383962 , n383963 , n383964 , n383965 , n383966 , 
     n383967 , n383968 , n383969 , n383970 , n383971 , n383972 , n383973 , n383974 , n383975 , n383976 , 
     n383977 , n383978 , n383979 , n383980 , n383981 , n383982 , n383983 , n383984 , n383985 , n383986 , 
     n383987 , n383988 , n383989 , n383990 , n383991 , n383992 , n383993 , n383994 , n383995 , n383996 , 
     n383997 , n383998 , n383999 , n384000 , n384001 , n384002 , n384003 , n384004 , n384005 , n384006 , 
     n384007 , n384008 , n384009 , n384010 , n384011 , n384012 , n384013 , n384014 , n384015 , n384016 , 
     n384017 , n384018 , n384019 , n384020 , n384021 , n384022 , n384023 , n384024 , n384025 , n384026 , 
     n384027 , n384028 , n384029 , n384030 , n384031 , n384032 , n384033 , n384034 , n384035 , n384036 , 
     n384037 , n384038 , n384039 , n384040 , n384041 , n384042 , n384043 , n384044 , n384045 , n384046 , 
     n384047 , n384048 , n384049 , n384050 , n384051 , n384052 , n384053 , n384054 , n384055 , n384056 , 
     n384057 , n384058 , n384059 , n384060 , n384061 , n384062 , n384063 , n384064 , n384065 , n384066 , 
     n384067 , n384068 , n384069 , n384070 , n384071 , n384072 , n384073 , n384074 , n384075 , n384076 , 
     n384077 , n384078 , n384079 , n384080 , n384081 , n384082 , n384083 , n384084 , n384085 , n384086 , 
     n384087 , n384088 , n384089 , n384090 , n384091 , n384092 , n384093 , n384094 , n384095 , n384096 , 
     n384097 , n384098 , n384099 , n384100 , n384101 , n384102 , n384103 , n384104 , n384105 , n384106 , 
     n384107 , n384108 , n384109 , n384110 , n384111 , n384112 , n384113 , n384114 , n384115 , n384116 , 
     n384117 , n384118 , n384119 , n384120 , n384121 , n384122 , n384123 , n384124 , n384125 , n384126 , 
     n384127 , n384128 , n384129 , n384130 , n384131 , n384132 , n384133 , n384134 , n384135 , n384136 , 
     n384137 , n384138 , n384139 , n384140 , n384141 , n384142 , n384143 , n384144 , n384145 , n384146 , 
     n384147 , n384148 , n384149 , n384150 , n384151 , n384152 , n384153 , n384154 , n384155 , n384156 , 
     n384157 , n384158 , n384159 , n384160 , n384161 , n384162 , n384163 , n384164 , n384165 , n384166 , 
     n384167 , n384168 , n384169 , n384170 , n384171 , n384172 , n384173 , n384174 , n384175 , n384176 , 
     n384177 , n384178 , n384179 , n384180 , n384181 , n384182 , n384183 , n384184 , n384185 , n384186 , 
     n384187 , n384188 , n384189 , n384190 , n384191 , n384192 , n384193 , n384194 , n384195 , n384196 , 
     n384197 , n384198 , n384199 , n384200 , n384201 , n384202 , n384203 , n384204 , n384205 , n384206 , 
     n384207 , n384208 , n384209 , n384210 , n384211 , n384212 , n384213 , n384214 , n384215 , n384216 , 
     n384217 , n384218 , n384219 , n384220 , n384221 , n384222 , n384223 , n384224 , n384225 , n384226 , 
     n384227 , n384228 , n384229 , n384230 , n384231 , n384232 , n384233 , n384234 , n384235 , n384236 , 
     n384237 , n384238 , n384239 , n384240 , n384241 , n384242 , n384243 , n384244 , n384245 , n384246 , 
     n384247 , n384248 , n384249 , n384250 , n384251 , n384252 , n384253 , n384254 , n384255 , n384256 , 
     n384257 , n384258 , n384259 , n384260 , n384261 , n384262 , n384263 , n384264 , n384265 , n384266 , 
     n384267 , n384268 , n384269 , n384270 , n384271 , n384272 , n384273 , n384274 , n384275 , n384276 , 
     n384277 , n384278 , n384279 , n384280 , n384281 , n384282 , n384283 , n384284 , n384285 , n384286 , 
     n384287 , n384288 , n384289 , n384290 , n384291 , n384292 , n384293 , n384294 , n384295 , n384296 , 
     n384297 , n384298 , n384299 , n384300 , n384301 , n384302 , n384303 , n384304 , n384305 , n384306 , 
     n384307 , n384308 , n384309 , n384310 , n384311 , n384312 , n384313 , n384314 , n384315 , n384316 , 
     n384317 , n384318 , n384319 , n384320 , n384321 , n384322 , n384323 , n384324 , n384325 , n384326 , 
     n384327 , n384328 , n384329 , n384330 , n384331 , n384332 , n384333 , n384334 , n384335 , n384336 , 
     n384337 , n384338 , n384339 , n384340 , n384341 , n384342 , n384343 , n384344 , n384345 , n384346 , 
     n384347 , n384348 , n384349 , n384350 , n384351 , n384352 , n384353 , n384354 , n384355 , n384356 , 
     n384357 , n384358 , n384359 , n384360 , n384361 , n384362 , n384363 , n384364 , n384365 , n384366 , 
     n384367 , n384368 , n384369 , n384370 , n384371 , n384372 , n384373 , n384374 , n384375 , n384376 , 
     n384377 , n384378 , n384379 , n384380 , n384381 , n384382 , n384383 , n384384 , n384385 , n384386 , 
     n384387 , n384388 , n384389 , n384390 , n384391 , n384392 , n384393 , n384394 , n384395 , n384396 , 
     n384397 , n384398 , n384399 , n384400 , n384401 , n384402 , n384403 , n384404 , n384405 , n384406 , 
     n384407 , n384408 , n384409 , n384410 , n384411 , n384412 , n384413 , n384414 , n384415 , n384416 , 
     n384417 , n384418 , n384419 , n384420 , n384421 , n384422 , n384423 , n384424 , n384425 , n384426 , 
     n384427 , n384428 , n384429 , n384430 , n384431 , n384432 , n384433 , n384434 , n384435 , n384436 , 
     n384437 , n384438 , n384439 , n384440 , n384441 , n384442 , n384443 , n384444 , n384445 , n384446 , 
     n384447 , n384448 , n384449 , n384450 , n384451 , n384452 , n384453 , n384454 , n384455 , n384456 , 
     n384457 , n384458 , n384459 , n384460 , n384461 , n384462 , n384463 , n384464 , n384465 , n384466 , 
     n384467 , n384468 , n384469 , n384470 , n384471 , n384472 , n384473 , n384474 , n384475 , n384476 , 
     n384477 , n384478 , n384479 , n384480 , n384481 , n384482 , n384483 , n384484 , n384485 , n384486 , 
     n384487 , n384488 , n384489 , n384490 , n384491 , n384492 , n384493 , n384494 , n384495 , n384496 , 
     n384497 , n384498 , n384499 , n384500 , n384501 , n384502 , n384503 , n384504 , n384505 , n384506 , 
     n384507 , n384508 , n384509 , n384510 , n384511 , n384512 , n384513 , n384514 , n384515 , n384516 , 
     n384517 , n384518 , n384519 , n384520 , n384521 , n384522 , n384523 , n384524 , n384525 , n384526 , 
     n384527 , n384528 , n384529 , n384530 , n384531 , n384532 , n384533 , n384534 , n384535 , n384536 , 
     n384537 , n384538 , n384539 , n384540 , n384541 , n384542 , n384543 , n384544 , n384545 , n384546 , 
     n384547 , n384548 , n384549 , n384550 , n384551 , n384552 , n384553 , n384554 , n384555 , n384556 , 
     n384557 , n384558 , n384559 , n384560 , n384561 , n384562 , n384563 , n384564 , n384565 , n384566 , 
     n384567 , n384568 , n384569 , n384570 , n384571 , n384572 , n384573 , n384574 , n384575 , n384576 , 
     n384577 , n384578 , n384579 , n384580 , n384581 , n384582 , n384583 , n384584 , n384585 , n384586 , 
     n384587 , n384588 , n384589 , n384590 , n384591 , n384592 , n384593 , n384594 , n384595 , n384596 , 
     n384597 , n384598 , n384599 , n384600 , n384601 , n384602 , n384603 , n384604 , n384605 , n384606 , 
     n384607 , n384608 , n384609 , n384610 , n384611 , n384612 , n384613 , n384614 , n384615 , n384616 , 
     n384617 , n384618 , n384619 , n384620 , n384621 , n384622 , n384623 , n384624 , n384625 , n384626 , 
     n384627 , n384628 , n384629 , n384630 , n384631 , n384632 , n384633 , n384634 , n384635 , n384636 , 
     n384637 , n384638 , n384639 , n384640 , n384641 , n384642 , n384643 , n384644 , n384645 , n384646 , 
     n384647 , n384648 , n384649 , n384650 , n384651 , n384652 , n384653 , n384654 , n384655 , n384656 , 
     n384657 , n384658 , n384659 , n384660 , n384661 , n384662 , n384663 , n384664 , n384665 , n384666 , 
     n384667 , n384668 , n384669 , n384670 , n384671 , n384672 , n384673 , n384674 , n384675 , n384676 , 
     n384677 , n384678 , n384679 , n384680 , n384681 , n384682 , n384683 , n384684 , n384685 , n384686 , 
     n384687 , n384688 , n384689 , n384690 , n384691 , n384692 , n384693 , n384694 , n384695 , n384696 , 
     n384697 , n384698 , n384699 , n384700 , n384701 , n384702 , n384703 , n384704 , n384705 , n384706 , 
     n384707 , n384708 , n384709 , n384710 , n384711 , n384712 , n384713 , n384714 , n384715 , n384716 , 
     n384717 , n384718 , n384719 , n384720 , n384721 , n384722 , n384723 , n384724 , n384725 , n384726 , 
     n384727 , n384728 , n384729 , n384730 , n384731 , n384732 , n384733 , n384734 , n384735 , n384736 , 
     n384737 , n384738 , n384739 , n384740 , n384741 , n384742 , n384743 , n384744 , n384745 , n384746 , 
     n384747 , n384748 , n384749 , n384750 , n384751 , n384752 , n384753 , n384754 , n384755 , n384756 , 
     n384757 , n384758 , n384759 , n384760 , n384761 , n384762 , n384763 , n384764 , n384765 , n384766 , 
     n384767 , n384768 , n384769 , n384770 , n384771 , n384772 , n384773 , n384774 , n384775 , n384776 , 
     n384777 , n384778 , n384779 , n384780 , n384781 , n384782 , n384783 , n384784 , n384785 , n384786 , 
     n384787 , n384788 , n384789 , n384790 , n384791 , n384792 , n384793 , n384794 , n384795 , n384796 , 
     n384797 , n384798 , n384799 , n384800 , n384801 , n384802 , n384803 , n384804 , n384805 , n384806 , 
     n384807 , n384808 , n384809 , n384810 , n384811 , n384812 , n384813 , n384814 , n384815 , n384816 , 
     n384817 , n384818 , n384819 , n384820 , n384821 , n384822 , n384823 , n384824 , n384825 , n384826 , 
     n384827 , n384828 , n384829 , n384830 , n384831 , n384832 , n384833 , n384834 , n384835 , n384836 , 
     n384837 , n384838 , n384839 , n384840 , n384841 , n384842 , n384843 , n384844 , n384845 , n384846 , 
     n384847 , n384848 , n384849 , n384850 , n384851 , n384852 , n384853 , n384854 , n384855 , n384856 , 
     n384857 , n384858 , n384859 , n384860 , n384861 , n384862 , n384863 , n384864 , n384865 , n384866 , 
     n384867 , n384868 , n384869 , n384870 , n384871 , n384872 , n384873 , n384874 , n384875 , n384876 , 
     n384877 , n384878 , n384879 , n384880 , n384881 , n384882 , n384883 , n384884 , n384885 , n384886 , 
     n384887 , n384888 , n384889 , n384890 , n384891 , n384892 , n384893 , n384894 , n384895 , n384896 , 
     n384897 , n384898 , n384899 , n384900 , n384901 , n384902 , n384903 , n384904 , n384905 , n384906 , 
     n384907 , n384908 , n384909 , n384910 , n384911 , n384912 , n384913 , n384914 , n384915 , n384916 , 
     n384917 , n384918 , n384919 , n384920 , n384921 , n384922 , n384923 , n384924 , n384925 , n384926 , 
     n384927 , n384928 , n384929 , n384930 , n384931 , n384932 , n384933 , n384934 , n384935 , n384936 , 
     n384937 , n384938 , n384939 , n384940 , n384941 , n384942 , n384943 , n384944 , n384945 , n384946 , 
     n384947 , n384948 , n384949 , n384950 , n384951 , n384952 , n384953 , n384954 , n384955 , n384956 , 
     n384957 , n384958 , n384959 , n384960 , n384961 , n384962 , n384963 , n384964 , n384965 , n384966 , 
     n384967 , n384968 , n384969 , n384970 , n384971 , n384972 , n384973 , n384974 , n384975 , n384976 , 
     n384977 , n384978 , n384979 , n384980 , n384981 , n384982 , n384983 , n384984 , n384985 , n384986 , 
     n384987 , n384988 , n384989 , n384990 , n384991 , n384992 , n384993 , n384994 , n384995 , n384996 , 
     n384997 , n384998 , n384999 , n385000 , n385001 , n385002 , n385003 , n385004 , n385005 , n385006 , 
     n385007 , n385008 , n385009 , n385010 , n385011 , n385012 , n385013 , n385014 , n385015 , n385016 , 
     n385017 , n385018 , n385019 , n385020 , n385021 , n385022 , n385023 , n385024 , n385025 , n385026 , 
     n385027 , n385028 , n385029 , n385030 , n385031 , n385032 , n385033 , n385034 , n385035 , n385036 , 
     n385037 , n385038 , n385039 , n385040 , n385041 , n385042 , n385043 , n385044 , n385045 , n385046 , 
     n385047 , n385048 , n385049 , n385050 , n385051 , n385052 , n385053 , n385054 , n385055 , n385056 , 
     n385057 , n385058 , n385059 , n385060 , n385061 , n385062 , n385063 , n385064 , n385065 , n385066 , 
     n385067 , n385068 , n385069 , n385070 , n385071 , n385072 , n385073 , n385074 , n385075 , n385076 , 
     n385077 , n385078 , n385079 , n385080 , n385081 , n385082 , n385083 , n385084 , n385085 , n385086 , 
     n385087 , n385088 , n385089 , n385090 , n385091 , n385092 , n385093 , n385094 , n385095 , n385096 , 
     n385097 , n385098 , n385099 , n385100 , n385101 , n385102 , n385103 , n385104 , n385105 , n385106 , 
     n385107 , n385108 , n385109 , n385110 , n385111 , n385112 , n385113 , n385114 , n385115 , n385116 , 
     n385117 , n385118 , n385119 , n385120 , n385121 , n385122 , n385123 , n385124 , n385125 , n385126 , 
     n385127 , n385128 , n385129 , n385130 , n385131 , n385132 , n385133 , n385134 , n385135 , n385136 , 
     n385137 , n385138 , n385139 , n385140 , n385141 , n385142 , n385143 , n385144 , n385145 , n385146 , 
     n385147 , n385148 , n385149 , n385150 , n385151 , n385152 , n385153 , n385154 , n385155 , n385156 , 
     n385157 , n385158 , n385159 , n385160 , n385161 , n385162 , n385163 , n385164 , n385165 , n385166 , 
     n385167 , n385168 , n385169 , n385170 , n385171 , n385172 , n385173 , n385174 , n385175 , n385176 , 
     n385177 , n385178 , n385179 , n385180 , n385181 , n385182 , n385183 , n385184 , n385185 , n385186 , 
     n385187 , n385188 , n385189 , n385190 , n385191 , n385192 , n385193 , n385194 , n385195 , n385196 , 
     n385197 , n385198 , n385199 , n385200 , n385201 , n385202 , n385203 , n385204 , n385205 , n385206 , 
     n385207 , n385208 , n385209 , n385210 , n385211 , n385212 , n385213 , n385214 , n385215 , n385216 , 
     n385217 , n385218 , n385219 , n385220 , n385221 , n385222 , n385223 , n385224 , n385225 , n385226 , 
     n385227 , n385228 , n385229 , n385230 , n385231 , n385232 , n385233 , n385234 , n385235 , n385236 , 
     n385237 , n385238 , n385239 , n385240 , n385241 , n385242 , n385243 , n385244 , n385245 , n385246 , 
     n385247 , n385248 , n385249 , n385250 , n385251 , n385252 , n385253 , n385254 , n385255 , n385256 , 
     n385257 , n385258 , n385259 , n385260 , n385261 , n385262 , n385263 , n385264 , n385265 , n385266 , 
     n385267 , n385268 , n385269 , n385270 , n385271 , n385272 , n385273 , n385274 , n385275 , n385276 , 
     n385277 , n385278 , n385279 , n385280 , n385281 , n385282 , n385283 , n385284 , n385285 , n385286 , 
     n385287 , n385288 , n385289 , n385290 , n385291 , n385292 , n385293 , n385294 , n385295 , n385296 , 
     n385297 , n385298 , n385299 , n385300 , n385301 , n385302 , n385303 , n385304 , n385305 , n385306 , 
     n385307 , n385308 , n385309 , n385310 , n385311 , n385312 , n385313 , n385314 , n385315 , n385316 , 
     n385317 , n385318 , n385319 , n385320 , n385321 , n385322 , n385323 , n385324 , n385325 , n385326 , 
     n385327 , n385328 , n385329 , n385330 , n385331 , n385332 , n385333 , n385334 , n385335 , n385336 , 
     n385337 , n385338 , n385339 , n385340 , n385341 , n385342 , n385343 , n385344 , n385345 , n385346 , 
     n385347 , n385348 , n385349 , n385350 , n385351 , n385352 , n385353 , n385354 , n385355 , n385356 , 
     n385357 , n385358 , n385359 , n385360 , n385361 , n385362 , n385363 , n385364 , n385365 , n385366 , 
     n385367 , n385368 , n385369 , n385370 , n385371 , n385372 , n385373 , n385374 , n385375 , n385376 , 
     n385377 , n385378 , n385379 , n385380 , n385381 , n385382 , n385383 , n385384 , n385385 , n385386 , 
     n385387 , n385388 , n385389 , n385390 , n385391 , n385392 , n385393 , n385394 , n385395 , n385396 , 
     n385397 , n385398 , n385399 , n385400 , n385401 , n385402 , n385403 , n385404 , n385405 , n385406 , 
     n385407 , n385408 , n385409 , n385410 , n385411 , n385412 , n385413 , n385414 , n385415 , n385416 , 
     n385417 , n385418 , n385419 , n385420 , n385421 , n385422 , n385423 , n385424 , n385425 , n385426 , 
     n385427 , n385428 , n385429 , n385430 , n385431 , n385432 , n385433 , n385434 , n385435 , n385436 , 
     n385437 , n385438 , n385439 , n385440 , n385441 , n385442 , n385443 , n385444 , n385445 , n385446 , 
     n385447 , n385448 , n385449 , n385450 , n385451 , n385452 , n385453 , n385454 , n385455 , n385456 , 
     n385457 , n385458 , n385459 , n385460 , n385461 , n385462 , n385463 , n385464 , n385465 , n385466 , 
     n385467 , n385468 , n385469 , n385470 , n385471 , n385472 , n385473 , n385474 , n385475 , n385476 , 
     n385477 , n385478 , n385479 , n385480 , n385481 , n385482 , n385483 , n385484 , n385485 , n385486 , 
     n385487 , n385488 , n385489 , n385490 , n385491 , n385492 , n385493 , n385494 , n385495 , n385496 , 
     n385497 , n385498 , n385499 , n385500 , n385501 , n385502 , n385503 , n385504 , n385505 , n385506 , 
     n385507 , n385508 , n385509 , n385510 , n385511 , n385512 , n385513 , n385514 , n385515 , n385516 , 
     n385517 , n385518 , n385519 , n385520 , n385521 , n385522 , n385523 , n385524 , n385525 , n385526 , 
     n385527 , n385528 , n385529 , n385530 , n385531 , n385532 , n385533 , n385534 , n385535 , n385536 , 
     n385537 , n385538 , n385539 , n385540 , n385541 , n385542 , n385543 , n385544 , n385545 , n385546 , 
     n385547 , n385548 , n385549 , n385550 , n385551 , n385552 , n385553 , n385554 , n385555 , n385556 , 
     n385557 , n385558 , n385559 , n385560 , n385561 , n385562 , n385563 , n385564 , n385565 , n385566 , 
     n385567 , n385568 , n385569 , n385570 , n385571 , n385572 , n385573 , n385574 , n385575 , n385576 , 
     n385577 , n385578 , n385579 , n385580 , n385581 , n385582 , n385583 , n385584 , n385585 , n385586 , 
     n385587 , n385588 , n385589 , n385590 , n385591 , n385592 , n385593 , n385594 , n385595 , n385596 , 
     n385597 , n385598 , n385599 , n385600 , n385601 , n385602 , n385603 , n385604 , n385605 , n385606 , 
     n385607 , n385608 , n385609 , n385610 , n385611 , n385612 , n385613 , n385614 , n385615 , n385616 , 
     n385617 , n385618 , n385619 , n385620 , n385621 , n385622 , n385623 , n385624 , n385625 , n385626 , 
     n385627 , n385628 , n385629 , n385630 , n385631 , n385632 , n385633 , n385634 , n385635 , n385636 , 
     n385637 , n385638 , n385639 , n385640 , n385641 , n385642 , n385643 , n385644 , n385645 , n385646 , 
     n385647 , n385648 , n385649 , n385650 , n385651 , n385652 , n385653 , n385654 , n385655 , n385656 , 
     n385657 , n385658 , n385659 , n385660 , n385661 , n385662 , n385663 , n385664 , n385665 , n385666 , 
     n385667 , n385668 , n385669 , n385670 , n385671 , n385672 , n385673 , n385674 , n385675 , n385676 , 
     n385677 , n385678 , n385679 , n385680 , n385681 , n385682 , n385683 , n385684 , n385685 , n385686 , 
     n385687 , n385688 , n385689 , n385690 , n385691 , n385692 , n385693 , n385694 , n385695 , n385696 , 
     n385697 , n385698 , n385699 , n385700 , n385701 , n385702 , n385703 , n385704 , n385705 , n385706 , 
     n385707 , n385708 , n385709 , n385710 , n385711 , n385712 , n385713 , n385714 , n385715 , n385716 , 
     n385717 , n385718 , n385719 , n385720 , n385721 , n385722 , n385723 , n385724 , n385725 , n385726 , 
     n385727 , n385728 , n385729 , n385730 , n385731 , n385732 , n385733 , n385734 , n385735 , n385736 , 
     n385737 , n385738 , n385739 , n385740 , n385741 , n385742 , n385743 , n385744 , n385745 , n385746 , 
     n385747 , n385748 , n385749 , n385750 , n385751 , n385752 , n385753 , n385754 , n385755 , n385756 , 
     n385757 , n385758 , n385759 , n385760 , n385761 , n385762 , n385763 , n385764 , n385765 , n385766 , 
     n385767 , n385768 , n385769 , n385770 , n385771 , n385772 , n385773 , n385774 , n385775 , n385776 , 
     n385777 , n385778 , n385779 , n385780 , n385781 , n385782 , n385783 , n385784 , n385785 , n385786 , 
     n385787 , n385788 , n385789 , n385790 , n385791 , n385792 , n385793 , n385794 , n385795 , n385796 , 
     n385797 , n385798 , n385799 , n385800 , n385801 , n385802 , n385803 , n385804 , n385805 , n385806 , 
     n385807 , n385808 , n385809 , n385810 , n385811 , n385812 , n385813 , n385814 , n385815 , n385816 , 
     n385817 , n385818 , n385819 , n385820 , n385821 , n385822 , n385823 , n385824 , n385825 , n385826 , 
     n385827 , n385828 , n385829 , n385830 , n385831 , n385832 , n385833 , n385834 , n385835 , n385836 , 
     n385837 , n385838 , n385839 , n385840 , n385841 , n385842 , n385843 , n385844 , n385845 , n385846 , 
     n385847 , n385848 , n385849 , n385850 , n385851 , n385852 , n385853 , n385854 , n385855 , n385856 , 
     n385857 , n385858 , n385859 , n385860 , n385861 , n385862 , n385863 , n385864 , n385865 , n385866 , 
     n385867 , n385868 , n385869 , n385870 , n385871 , n385872 , n385873 , n385874 , n385875 , n385876 , 
     n385877 , n385878 , n385879 , n385880 , n385881 , n385882 , n385883 , n385884 , n385885 , n385886 , 
     n385887 , n385888 , n385889 , n385890 , n385891 , n385892 , n385893 , n385894 , n385895 , n385896 , 
     n385897 , n385898 , n385899 , n385900 , n385901 , n385902 , n385903 , n385904 , n385905 , n385906 , 
     n385907 , n385908 , n385909 , n385910 , n385911 , n385912 , n385913 , n385914 , n385915 , n385916 , 
     n385917 , n385918 , n385919 , n385920 , n385921 , n385922 , n385923 , n385924 , n385925 , n385926 , 
     n385927 , n385928 , n385929 , n385930 , n385931 , n385932 , n385933 , n385934 , n385935 , n385936 , 
     n385937 , n385938 , n385939 , n385940 , n385941 , n385942 , n385943 , n385944 , n385945 , n385946 , 
     n385947 , n385948 , n385949 , n385950 , n385951 , n385952 , n385953 , n385954 , n385955 , n385956 , 
     n385957 , n385958 , n385959 , n385960 , n385961 , n385962 , n385963 , n385964 , n385965 , n385966 , 
     n385967 , n385968 , n385969 , n385970 , n385971 , n385972 , n385973 , n385974 , n385975 , n385976 , 
     n385977 , n385978 , n385979 , n385980 , n385981 , n385982 , n385983 , n385984 , n385985 , n385986 , 
     n385987 , n385988 , n385989 , n385990 , n385991 , n385992 , n385993 , n385994 , n385995 , n385996 , 
     n385997 , n385998 , n385999 , n386000 , n386001 , n386002 , n386003 , n386004 , n386005 , n386006 , 
     n386007 , n386008 , n386009 , n386010 , n386011 , n386012 , n386013 , n386014 , n386015 , n386016 , 
     n386017 , n386018 , n386019 , n386020 , n386021 , n386022 , n386023 , n386024 , n386025 , n386026 , 
     n386027 , n386028 , n386029 , n386030 , n386031 , n386032 , n386033 , n386034 , n386035 , n386036 , 
     n386037 , n386038 , n386039 , n386040 , n386041 , n386042 , n386043 , n386044 , n386045 , n386046 , 
     n386047 , n386048 , n386049 , n386050 , n386051 , n386052 , n386053 , n386054 , n386055 , n386056 , 
     n386057 , n386058 , n386059 , n386060 , n386061 , n386062 , n386063 , n386064 , n386065 , n386066 , 
     n386067 , n386068 , n386069 , n386070 , n386071 , n386072 , n386073 , n386074 , n386075 , n386076 , 
     n386077 , n386078 , n386079 , n386080 , n386081 , n386082 , n386083 , n386084 , n386085 , n386086 , 
     n386087 , n386088 , n386089 , n386090 , n386091 , n386092 , n386093 , n386094 , n386095 , n386096 , 
     n386097 , n386098 , n386099 , n386100 , n386101 , n386102 , n386103 , n386104 , n386105 , n386106 , 
     n386107 , n386108 , n386109 , n386110 , n386111 , n386112 , n386113 , n386114 , n386115 , n386116 , 
     n386117 , n386118 , n386119 , n386120 , n386121 , n386122 , n386123 , n386124 , n386125 , n386126 , 
     n386127 , n386128 , n386129 , n386130 , n386131 , n386132 , n386133 , n386134 , n386135 , n386136 , 
     n386137 , n386138 , n386139 , n386140 , n386141 , n386142 , n386143 , n386144 , n386145 , n386146 , 
     n386147 , n386148 , n386149 , n386150 , n386151 , n386152 , n386153 , n386154 , n386155 , n386156 , 
     n386157 , n386158 , n386159 , n386160 , n386161 , n386162 , n386163 , n386164 , n386165 , n386166 , 
     n386167 , n386168 , n386169 , n386170 , n386171 , n386172 , n386173 , n386174 , n386175 , n386176 , 
     n386177 , n386178 , n386179 , n386180 , n386181 , n386182 , n386183 , n386184 , n386185 , n386186 , 
     n386187 , n386188 , n386189 , n386190 , n386191 , n386192 , n386193 , n386194 , n386195 , n386196 , 
     n386197 , n386198 , n386199 , n386200 , n386201 , n386202 , n386203 , n386204 , n386205 , n386206 , 
     n386207 , n386208 , n386209 , n386210 , n386211 , n386212 , n386213 , n386214 , n386215 , n386216 , 
     n386217 , n386218 , n386219 , n386220 , n386221 , n386222 , n386223 , n386224 , n386225 , n386226 , 
     n386227 , n386228 , n386229 , n386230 , n386231 , n386232 , n386233 , n386234 , n386235 , n386236 , 
     n386237 , n386238 , n386239 , n386240 , n386241 , n386242 , n386243 , n386244 , n386245 , n386246 , 
     n386247 , n386248 , n386249 , n386250 , n386251 , n386252 , n386253 , n386254 , n386255 , n386256 , 
     n386257 , n386258 , n386259 , n386260 , n386261 , n386262 , n386263 , n386264 , n386265 , n386266 , 
     n386267 , n386268 , n386269 , n386270 , n386271 , n386272 , n386273 , n386274 , n386275 , n386276 , 
     n386277 , n386278 , n386279 , n386280 , n386281 , n386282 , n386283 , n386284 , n386285 , n386286 , 
     n386287 , n386288 , n386289 , n386290 , n386291 , n386292 , n386293 , n386294 , n386295 , n386296 , 
     n386297 , n386298 , n386299 , n386300 , n386301 , n386302 , n386303 , n386304 , n386305 , n386306 , 
     n386307 , n386308 , n386309 , n386310 , n386311 , n386312 , n386313 , n386314 , n386315 , n386316 , 
     n386317 , n386318 , n386319 , n386320 , n386321 , n386322 , n386323 , n386324 , n386325 , n386326 , 
     n386327 , n386328 , n386329 , n386330 , n386331 , n386332 , n386333 , n386334 , n386335 , n386336 , 
     n386337 , n386338 , n386339 , n386340 , n386341 , n386342 , n386343 , n386344 , n386345 , n386346 , 
     n386347 , n386348 , n386349 , n386350 , n386351 , n386352 , n386353 , n386354 , n386355 , n386356 , 
     n386357 , n386358 , n386359 , n386360 , n386361 , n386362 , n386363 , n386364 , n386365 , n386366 , 
     n386367 , n386368 , n386369 , n386370 , n386371 , n386372 , n386373 , n386374 , n386375 , n386376 , 
     n386377 , n386378 , n386379 , n386380 , n386381 , n386382 , n386383 , n386384 , n386385 , n386386 , 
     n386387 , n386388 , n386389 , n386390 , n386391 , n386392 , n386393 , n386394 , n386395 , n386396 , 
     n386397 , n386398 , n386399 , n386400 , n386401 , n386402 , n386403 , n386404 , n386405 , n386406 , 
     n386407 , n386408 , n386409 , n386410 , n386411 , n386412 , n386413 , n386414 , n386415 , n386416 , 
     n386417 , n386418 , n386419 , n386420 , n386421 , n386422 , n386423 , n386424 , n386425 , n386426 , 
     n386427 , n386428 , n386429 , n386430 , n386431 , n386432 , n386433 , n386434 , n386435 , n386436 , 
     n386437 , n386438 , n386439 , n386440 , n386441 , n386442 , n386443 , n386444 , n386445 , n386446 , 
     n386447 , n386448 , n386449 , n386450 , n386451 , n386452 , n386453 , n386454 , n386455 , n386456 , 
     n386457 , n386458 , n386459 , n386460 , n386461 , n386462 , n386463 , n386464 , n386465 , n386466 , 
     n386467 , n386468 , n386469 , n386470 , n386471 , n386472 , n386473 , n386474 , n386475 , n386476 , 
     n386477 , n386478 , n386479 , n386480 , n386481 , n386482 , n386483 , n386484 , n386485 , n386486 , 
     n386487 , n386488 , n386489 , n386490 , n386491 , n386492 , n386493 , n386494 , n386495 , n386496 , 
     n386497 , n386498 , n386499 , n386500 , n386501 , n386502 , n386503 , n386504 , n386505 , n386506 , 
     n386507 , n386508 , n386509 , n386510 , n386511 , n386512 , n386513 , n386514 , n386515 , n386516 , 
     n386517 , n386518 , n386519 , n386520 , n386521 , n386522 , n386523 , n386524 , n386525 , n386526 , 
     n386527 , n386528 , n386529 , n386530 , n386531 , n386532 , n386533 , n386534 , n386535 , n386536 , 
     n386537 , n386538 , n386539 , n386540 , n386541 , n386542 , n386543 , n386544 , n386545 , n386546 , 
     n386547 , n386548 , n386549 , n386550 , n386551 , n386552 , n386553 , n386554 , n386555 , n386556 , 
     n386557 , n386558 , n386559 , n386560 , n386561 , n386562 , n386563 , n386564 , n386565 , n386566 , 
     n386567 , n386568 , n386569 , n386570 , n386571 , n386572 , n386573 , n386574 , n386575 , n386576 , 
     n386577 , n386578 , n386579 , n386580 , n386581 , n386582 , n386583 , n386584 , n386585 , n386586 , 
     n386587 , n386588 , n386589 , n386590 , n386591 , n386592 , n386593 , n386594 , n386595 , n386596 , 
     n386597 , n386598 , n386599 , n386600 , n386601 , n386602 , n386603 , n386604 , n386605 , n386606 , 
     n386607 , n386608 , n386609 , n386610 , n386611 , n386612 , n386613 , n386614 , n386615 , n386616 , 
     n386617 , n386618 , n386619 , n386620 , n386621 , n386622 , n386623 , n386624 , n386625 , n386626 , 
     n386627 , n386628 , n386629 , n386630 , n386631 , n386632 , n386633 , n386634 , n386635 , n386636 , 
     n386637 , n386638 , n386639 , n386640 , n386641 , n386642 , n386643 , n386644 , n386645 , n386646 , 
     n386647 , n386648 , n386649 , n386650 , n386651 , n386652 , n386653 , n386654 , n386655 , n386656 , 
     n386657 , n386658 , n386659 , n386660 , n386661 , n386662 , n386663 , n386664 , n386665 , n386666 , 
     n386667 , n386668 , n386669 , n386670 , n386671 , n386672 , n386673 , n386674 , n386675 , n386676 , 
     n386677 , n386678 , n386679 , n386680 , n386681 , n386682 , n386683 , n386684 , n386685 , n386686 , 
     n386687 , n386688 , n386689 , n386690 , n386691 , n386692 , n386693 , n386694 , n386695 , n386696 , 
     n386697 , n386698 , n386699 , n386700 , n386701 , n386702 , n386703 , n386704 , n386705 , n386706 , 
     n386707 , n386708 , n386709 , n386710 , n386711 , n386712 , n386713 , n386714 , n386715 , n386716 , 
     n386717 , n386718 , n386719 , n386720 , n386721 , n386722 , n386723 , n386724 , n386725 , n386726 , 
     n386727 , n386728 , n386729 , n386730 , n386731 , n386732 , n386733 , n386734 , n386735 , n386736 , 
     n386737 , n386738 , n386739 , n386740 , n386741 , n386742 , n386743 , n386744 , n386745 , n386746 , 
     n386747 , n386748 , n386749 , n386750 , n386751 , n386752 , n386753 , n386754 , n386755 , n386756 , 
     n386757 , n386758 , n386759 , n386760 , n386761 , n386762 , n386763 , n386764 , n386765 , n386766 , 
     n386767 , n386768 , n386769 , n386770 , n386771 , n386772 , n386773 , n386774 , n386775 , n386776 , 
     n386777 , n386778 , n386779 , n386780 , n386781 , n386782 , n386783 , n386784 , n386785 , n386786 , 
     n386787 , n386788 , n386789 , n386790 , n386791 , n386792 , n386793 , n386794 , n386795 , n386796 , 
     n386797 , n386798 , n386799 , n386800 , n386801 , n386802 , n386803 , n386804 , n386805 , n386806 , 
     n386807 , n386808 , n386809 , n386810 , n386811 , n386812 , n386813 , n386814 , n386815 , n386816 , 
     n386817 , n386818 , n386819 , n386820 , n386821 , n386822 , n386823 , n386824 , n386825 , n386826 , 
     n386827 , n386828 , n386829 , n386830 , n386831 , n386832 , n386833 , n386834 , n386835 , n386836 , 
     n386837 , n386838 , n386839 , n386840 , n386841 , n386842 , n386843 , n386844 , n386845 , n386846 , 
     n386847 , n386848 , n386849 , n386850 , n386851 , n386852 , n386853 , n386854 , n386855 , n386856 , 
     n386857 , n386858 , n386859 , n386860 , n386861 , n386862 , n386863 , n386864 , n386865 , n386866 , 
     n386867 , n386868 , n386869 , n386870 , n386871 , n386872 , n386873 , n386874 , n386875 , n386876 , 
     n386877 , n386878 , n386879 , n386880 , n386881 , n386882 , n386883 , n386884 , n386885 , n386886 , 
     n386887 , n386888 , n386889 , n386890 , n386891 , n386892 , n386893 , n386894 , n386895 , n386896 , 
     n386897 , n386898 , n386899 , n386900 , n386901 , n386902 , n386903 , n386904 , n386905 , n386906 , 
     n386907 , n386908 , n386909 , n386910 , n386911 , n386912 , n386913 , n386914 , n386915 , n386916 , 
     n386917 , n386918 , n386919 , n386920 , n386921 , n386922 , n386923 , n386924 , n386925 , n386926 , 
     n386927 , n386928 , n386929 , n386930 , n386931 , n386932 , n386933 , n386934 , n386935 , n386936 , 
     n386937 , n386938 , n386939 , n386940 , n386941 , n386942 , n386943 , n386944 , n386945 , n386946 , 
     n386947 , n386948 , n386949 , n386950 , n386951 , n386952 , n386953 , n386954 , n386955 , n386956 , 
     n386957 , n386958 , n386959 , n386960 , n386961 , n386962 , n386963 , n386964 , n386965 , n386966 , 
     n386967 , n386968 , n386969 , n386970 , n386971 , n386972 , n386973 , n386974 , n386975 , n386976 , 
     n386977 , n386978 , n386979 , n386980 , n386981 , n386982 , n386983 , n386984 , n386985 , n386986 , 
     n386987 , n386988 , n386989 , n386990 , n386991 , n386992 , n386993 , n386994 , n386995 , n386996 , 
     n386997 , n386998 , n386999 , n387000 , n387001 , n387002 , n387003 , n387004 , n387005 , n387006 , 
     n387007 , n387008 , n387009 , n387010 , n387011 , n387012 , n387013 , n387014 , n387015 , n387016 , 
     n387017 , n387018 , n387019 , n387020 , n387021 , n387022 , n387023 , n387024 , n387025 , n387026 , 
     n387027 , n387028 , n387029 , n387030 , n387031 , n387032 , n387033 , n387034 , n387035 , n387036 , 
     n387037 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , 
     n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , 
     n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , 
     n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , 
     n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , 
     n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , 
     n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , 
     n30911 , n30912 , n30913 , n387110 , n387111 , n387112 , n387113 , n387114 , n387115 , n387116 , 
     n387117 , n387118 , n387119 , n387120 , n387121 , n387122 , n387123 , n387124 , n387125 , n387126 , 
     n387127 , n387128 , n387129 , n387130 , n387131 , n387132 , n387133 , n387134 , n387135 , n387136 , 
     n387137 , n387138 , n387139 , n387140 , n387141 , n387142 , n387143 , n387144 , n387145 , n387146 , 
     n387147 , n387148 , n387149 , n387150 , n387151 , n387152 , n387153 , n387154 , n387155 , n387156 , 
     n387157 , n387158 , n387159 , n387160 , n387161 , n387162 , n387163 , n387164 , n387165 , n387166 , 
     n387167 , n387168 , n387169 , n387170 , n387171 , n387172 , n387173 , n387174 , n387175 , n387176 , 
     n387177 , n387178 , n387179 , n387180 , n387181 , n387182 , n30987 , n30988 , n30989 , n30990 , 
     n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , 
     n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , 
     n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , 
     n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , 
     n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , 
     n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , 
     n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , 
     n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , 
     n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , 
     n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , 
     n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , 
     n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , 
     n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , 
     n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , 
     n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , 
     n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , 
     n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , 
     n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , 
     n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , 
     n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , 
     n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , 
     n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , 
     n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , 
     n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , 
     n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , 
     n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , 
     n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , 
     n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , 
     n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , 
     n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , 
     n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , 
     n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , 
     n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , 
     n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , 
     n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , 
     n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , 
     n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , 
     n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , 
     n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , 
     n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , 
     n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , 
     n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , 
     n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , 
     n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , 
     n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , 
     n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , 
     n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , 
     n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , 
     n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , 
     n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , 
     n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , 
     n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , 
     n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , 
     n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , 
     n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , 
     n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , 
     n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , 
     n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , 
     n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , 
     n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , 
     n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , 
     n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , 
     n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , 
     n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , 
     n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , 
     n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , 
     n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , 
     n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , 
     n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , 
     n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , 
     n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , 
     n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , 
     n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , 
     n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , 
     n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , 
     n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , 
     n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , 
     n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , 
     n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , 
     n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , 
     n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , 
     n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , 
     n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , 
     n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , 
     n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , 
     n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , 
     n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , 
     n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , 
     n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , 
     n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , 
     n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , 
     n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , 
     n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , 
     n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , 
     n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , 
     n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , 
     n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , 
     n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , 
     n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , 
     n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , 
     n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , 
     n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , 
     n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , 
     n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , 
     n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , 
     n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , 
     n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , 
     n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , 
     n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , 
     n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , 
     n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , 
     n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , 
     n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , 
     n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , 
     n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , 
     n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , 
     n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , 
     n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , 
     n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , 
     n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , 
     n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , 
     n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , 
     n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , 
     n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , 
     n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , 
     n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , 
     n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , 
     n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , 
     n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , 
     n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , 
     n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , 
     n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , 
     n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , 
     n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , 
     n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , 
     n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , 
     n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , 
     n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , 
     n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , 
     n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , 
     n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , 
     n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , 
     n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , 
     n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , 
     n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , 
     n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , 
     n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , 
     n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , 
     n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , 
     n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , 
     n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , 
     n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , 
     n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , 
     n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , 
     n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , 
     n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , 
     n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , 
     n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , 
     n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , 
     n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , 
     n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , 
     n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , 
     n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , 
     n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , 
     n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , 
     n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , 
     n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , 
     n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , 
     n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , 
     n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , 
     n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , 
     n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , 
     n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , 
     n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , 
     n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , 
     n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , 
     n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , 
     n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , 
     n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , 
     n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , 
     n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , 
     n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , 
     n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , 
     n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , 
     n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , 
     n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , 
     n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , 
     n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , 
     n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , 
     n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , 
     n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , 
     n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , 
     n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , 
     n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , 
     n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , 
     n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , 
     n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , 
     n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , 
     n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , 
     n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , 
     n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , 
     n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , 
     n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , 
     n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , 
     n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , 
     n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , 
     n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , 
     n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , 
     n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , 
     n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , 
     n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , 
     n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , 
     n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , 
     n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , 
     n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , 
     n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , 
     n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , 
     n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , 
     n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , 
     n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , 
     n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , 
     n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , 
     n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , 
     n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , 
     n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , 
     n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , 
     n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , 
     n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , 
     n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , 
     n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , 
     n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , 
     n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , 
     n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , 
     n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , 
     n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , 
     n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , 
     n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , 
     n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , 
     n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , 
     n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , 
     n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , 
     n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , 
     n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , 
     n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , 
     n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , 
     n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , 
     n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , 
     n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , 
     n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , 
     n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , 
     n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , 
     n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , 
     n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , 
     n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , 
     n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , 
     n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , 
     n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , 
     n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , 
     n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , 
     n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , 
     n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , 
     n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , 
     n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , 
     n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , 
     n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , 
     n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , 
     n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , 
     n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , 
     n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , 
     n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , 
     n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , 
     n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , 
     n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , 
     n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , 
     n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , 
     n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , 
     n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , 
     n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , 
     n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , 
     n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , 
     n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , 
     n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , 
     n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , 
     n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , 
     n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , 
     n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , 
     n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , 
     n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , 
     n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , 
     n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , 
     n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , 
     n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , 
     n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , 
     n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , 
     n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , 
     n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , 
     n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , 
     n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , 
     n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , 
     n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , 
     n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , 
     n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , 
     n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , 
     n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , 
     n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , 
     n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , 
     n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , 
     n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , 
     n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , 
     n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , 
     n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , 
     n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , 
     n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , 
     n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , 
     n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , 
     n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , 
     n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , 
     n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , 
     n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , 
     n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , 
     n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , 
     n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , 
     n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , 
     n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , 
     n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , 
     n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , 
     n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , 
     n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , 
     n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , 
     n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , 
     n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , 
     n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , 
     n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , 
     n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , 
     n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , 
     n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , 
     n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , 
     n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , 
     n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , 
     n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , 
     n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , 
     n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , 
     n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , 
     n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , 
     n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , 
     n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , 
     n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , 
     n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , 
     n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , 
     n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , 
     n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , 
     n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , 
     n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , 
     n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , 
     n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , 
     n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , 
     n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , 
     n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , 
     n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , 
     n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , 
     n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , 
     n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , 
     n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , 
     n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , 
     n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , 
     n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , 
     n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , 
     n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , 
     n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , 
     n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , 
     n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , 
     n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , 
     n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , 
     n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , 
     n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , 
     n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , 
     n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , 
     n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , 
     n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , 
     n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , 
     n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , 
     n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , 
     n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , 
     n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , 
     n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , 
     n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , 
     n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , 
     n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , 
     n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , 
     n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , 
     n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , 
     n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , 
     n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , 
     n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , 
     n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , 
     n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , 
     n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , 
     n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , 
     n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , 
     n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , 
     n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , 
     n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , 
     n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , 
     n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , 
     n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , 
     n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , 
     n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , 
     n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , 
     n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , 
     n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , 
     n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , 
     n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , 
     n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , 
     n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , 
     n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , 
     n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , 
     n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , 
     n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , 
     n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , 
     n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , 
     n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , 
     n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , 
     n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , 
     n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , 
     n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , 
     n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , 
     n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , 
     n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , 
     n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , 
     n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , 
     n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , 
     n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , 
     n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , 
     n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , 
     n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , 
     n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , 
     n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , 
     n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , 
     n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , 
     n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , 
     n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , 
     n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , 
     n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , 
     n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , 
     n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , 
     n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , 
     n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , 
     n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , 
     n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , 
     n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , 
     n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , 
     n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , 
     n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , 
     n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , 
     n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , 
     n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , 
     n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , 
     n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , 
     n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , 
     n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , 
     n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , 
     n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , 
     n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , 
     n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , 
     n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , 
     n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , 
     n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , 
     n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , 
     n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , 
     n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , 
     n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , 
     n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , 
     n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , 
     n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , 
     n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , 
     n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , 
     n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , 
     n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , 
     n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , 
     n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , 
     n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , 
     n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , 
     n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , 
     n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , 
     n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , 
     n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , 
     n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , 
     n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , 
     n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , 
     n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , 
     n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , 
     n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , 
     n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , 
     n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , 
     n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , 
     n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , 
     n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , 
     n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , 
     n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , 
     n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , 
     n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , 
     n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , 
     n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , 
     n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , 
     n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , 
     n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , 
     n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , 
     n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , 
     n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , 
     n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , 
     n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , 
     n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , 
     n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , 
     n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , 
     n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , 
     n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , 
     n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , 
     n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , 
     n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , 
     n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , 
     n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , 
     n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , 
     n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , 
     n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , 
     n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , 
     n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , 
     n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , 
     n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , 
     n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , 
     n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , 
     n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , 
     n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , 
     n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , 
     n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , 
     n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , 
     n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , 
     n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , 
     n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , 
     n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , 
     n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , 
     n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , 
     n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , 
     n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , 
     n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , 
     n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , 
     n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , 
     n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , 
     n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , 
     n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , 
     n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , 
     n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , 
     n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , 
     n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , 
     n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , 
     n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , 
     n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , 
     n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , 
     n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , 
     n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , 
     n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , 
     n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , 
     n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , 
     n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , 
     n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , 
     n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , 
     n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , 
     n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , 
     n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , 
     n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , 
     n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , 
     n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , 
     n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , 
     n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , 
     n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , 
     n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , 
     n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , 
     n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , 
     n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , 
     n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , 
     n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , 
     n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , 
     n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , 
     n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , 
     n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , 
     n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , 
     n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , 
     n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , 
     n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , 
     n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , 
     n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , 
     n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , 
     n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , 
     n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , 
     n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , 
     n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , 
     n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , 
     n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , 
     n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , 
     n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , 
     n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , 
     n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , 
     n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , 
     n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , 
     n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , 
     n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , 
     n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , 
     n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , 
     n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , 
     n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , 
     n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , 
     n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , 
     n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , 
     n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , 
     n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , 
     n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , 
     n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , 
     n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , 
     n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , 
     n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , 
     n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , 
     n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , 
     n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , 
     n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , 
     n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , 
     n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , 
     n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , 
     n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , 
     n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , 
     n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , 
     n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , 
     n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , 
     n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , 
     n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , 
     n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , 
     n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , 
     n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , 
     n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , 
     n37361 , n37362 , n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , 
     n37371 , n37372 , n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , 
     n37381 , n37382 , n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , 
     n37391 , n37392 , n37393 , n37394 , n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , 
     n37401 , n37402 , n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , 
     n37411 , n37412 , n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , 
     n37421 , n37422 , n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , 
     n37431 , n37432 , n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , 
     n37441 , n37442 , n37443 , n37444 , n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , 
     n37451 , n37452 , n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , 
     n37461 , n37462 , n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , 
     n37471 , n37472 , n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , 
     n37481 , n37482 , n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , 
     n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , 
     n37501 , n37502 , n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , 
     n37511 , n37512 , n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , 
     n37521 , n37522 , n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , 
     n37531 , n37532 , n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , 
     n37541 , n37542 , n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , 
     n37551 , n37552 , n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , 
     n37561 , n37562 , n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , 
     n37571 , n37572 , n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , 
     n37581 , n37582 , n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , 
     n37591 , n37592 , n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , 
     n37601 , n37602 , n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , 
     n37611 , n37612 , n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , 
     n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , 
     n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , 
     n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , 
     n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , 
     n37661 , n37662 , n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , 
     n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , 
     n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , 
     n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , 
     n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , 
     n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , 
     n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , 
     n37731 , n37732 , n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , 
     n37741 , n37742 , n37743 , n37744 , n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , 
     n37751 , n37752 , n37753 , n37754 , n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , 
     n37761 , n37762 , n37763 , n37764 , n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , 
     n37771 , n37772 , n37773 , n37774 , n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , 
     n37781 , n37782 , n37783 , n37784 , n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , 
     n37791 , n37792 , n37793 , n37794 , n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , 
     n37801 , n37802 , n37803 , n37804 , n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , 
     n37811 , n37812 , n37813 , n37814 , n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , 
     n37821 , n37822 , n37823 , n37824 , n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , 
     n37831 , n37832 , n37833 , n37834 , n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , 
     n37841 , n37842 , n37843 , n37844 , n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , 
     n37851 , n37852 , n37853 , n37854 , n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , 
     n37861 , n37862 , n37863 , n37864 , n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , 
     n37871 , n37872 , n37873 , n37874 , n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , 
     n37881 , n37882 , n37883 , n37884 , n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , 
     n37891 , n37892 , n37893 , n37894 , n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , 
     n37901 , n37902 , n37903 , n37904 , n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , 
     n37911 , n37912 , n37913 , n37914 , n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , 
     n37921 , n37922 , n37923 , n37924 , n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , 
     n37931 , n37932 , n37933 , n37934 , n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , 
     n37941 , n37942 , n37943 , n37944 , n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , 
     n37951 , n37952 , n37953 , n37954 , n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , 
     n37961 , n37962 , n37963 , n37964 , n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , 
     n37971 , n37972 , n37973 , n37974 , n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , 
     n37981 , n37982 , n37983 , n37984 , n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , 
     n37991 , n37992 , n37993 , n37994 , n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , 
     n38001 , n38002 , n38003 , n38004 , n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , 
     n38011 , n38012 , n38013 , n38014 , n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , 
     n38021 , n38022 , n38023 , n38024 , n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , 
     n38031 , n38032 , n38033 , n38034 , n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , 
     n38041 , n38042 , n38043 , n38044 , n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , 
     n38051 , n38052 , n38053 , n38054 , n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , 
     n38061 , n38062 , n38063 , n38064 , n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , 
     n38071 , n38072 , n38073 , n38074 , n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , 
     n38081 , n38082 , n38083 , n38084 , n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , 
     n38091 , n38092 , n38093 , n38094 , n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , 
     n38101 , n38102 , n38103 , n38104 , n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , 
     n38111 , n38112 , n38113 , n38114 , n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , 
     n38121 , n38122 , n38123 , n38124 , n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , 
     n38131 , n38132 , n38133 , n38134 , n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , 
     n38141 , n38142 , n38143 , n38144 , n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , 
     n38151 , n38152 , n38153 , n38154 , n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , 
     n38161 , n38162 , n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , 
     n38171 , n38172 , n38173 , n38174 , n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , 
     n38181 , n38182 , n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , 
     n38191 , n38192 , n38193 , n38194 , n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , 
     n38201 , n38202 , n38203 , n38204 , n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , 
     n38211 , n38212 , n38213 , n38214 , n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , 
     n38221 , n38222 , n38223 , n38224 , n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , 
     n38231 , n38232 , n38233 , n38234 , n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , 
     n38241 , n38242 , n38243 , n38244 , n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , 
     n38251 , n38252 , n38253 , n38254 , n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , 
     n38261 , n38262 , n38263 , n38264 , n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , 
     n38271 , n38272 , n38273 , n38274 , n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , 
     n38281 , n38282 , n38283 , n38284 , n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , 
     n38291 , n38292 , n38293 , n38294 , n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , 
     n38301 , n38302 , n38303 , n38304 , n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , 
     n38311 , n38312 , n38313 , n38314 , n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , 
     n38321 , n38322 , n38323 , n38324 , n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , 
     n38331 , n38332 , n38333 , n38334 , n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , 
     n38341 , n38342 , n38343 , n38344 , n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , 
     n38351 , n38352 , n38353 , n38354 , n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , 
     n38361 , n38362 , n38363 , n38364 , n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , 
     n38371 , n38372 , n38373 , n38374 , n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , 
     n38381 , n38382 , n38383 , n38384 , n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , 
     n38391 , n38392 , n38393 , n38394 , n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , 
     n38401 , n38402 , n38403 , n38404 , n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , 
     n38411 , n38412 , n38413 , n38414 , n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , 
     n38421 , n38422 , n38423 , n38424 , n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , 
     n38431 , n38432 , n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , 
     n38441 , n38442 , n38443 , n38444 , n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , 
     n38451 , n38452 , n38453 , n38454 , n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , 
     n38461 , n38462 , n38463 , n38464 , n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , 
     n38471 , n38472 , n38473 , n38474 , n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , 
     n38481 , n38482 , n38483 , n38484 , n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , 
     n38491 , n38492 , n38493 , n38494 , n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , 
     n38501 , n38502 , n38503 , n38504 , n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , 
     n38511 , n38512 , n38513 , n38514 , n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , 
     n38521 , n38522 , n38523 , n38524 , n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , 
     n38531 , n38532 , n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , 
     n38541 , n38542 , n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , 
     n38551 , n38552 , n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , 
     n38561 , n38562 , n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , 
     n38571 , n38572 , n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , 
     n38581 , n38582 , n38583 , n38584 , n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , 
     n38591 , n38592 , n38593 , n38594 , n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , 
     n38601 , n38602 , n38603 , n38604 , n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , 
     n38611 , n38612 , n38613 , n38614 , n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , 
     n38621 , n38622 , n38623 , n38624 , n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , 
     n38631 , n38632 , n38633 , n38634 , n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , 
     n38641 , n38642 , n38643 , n38644 , n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , 
     n38651 , n38652 , n38653 , n38654 , n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , 
     n38661 , n38662 , n38663 , n38664 , n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , 
     n38671 , n38672 , n38673 , n38674 , n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , 
     n38681 , n38682 , n38683 , n38684 , n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , 
     n38691 , n38692 , n38693 , n38694 , n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , 
     n38701 , n38702 , n38703 , n38704 , n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , 
     n38711 , n38712 , n38713 , n38714 , n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , 
     n38721 , n38722 , n38723 , n38724 , n38725 , n38726 , n38727 , n38728 , n38729 , n38730 , 
     n38731 , n38732 , n38733 , n38734 , n38735 , n38736 , n38737 , n38738 , n38739 , n38740 , 
     n38741 , n38742 , n38743 , n38744 , n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , 
     n38751 , n38752 , n38753 , n38754 , n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , 
     n38761 , n38762 , n38763 , n38764 , n38765 , n38766 , n38767 , n38768 , n38769 , n38770 , 
     n38771 , n38772 , n38773 , n38774 , n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , 
     n38781 , n38782 , n38783 , n38784 , n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , 
     n38791 , n38792 , n38793 , n38794 , n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , 
     n38801 , n38802 , n38803 , n38804 , n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , 
     n38811 , n38812 , n38813 , n38814 , n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , 
     n38821 , n38822 , n38823 , n38824 , n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , 
     n38831 , n38832 , n38833 , n38834 , n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , 
     n38841 , n38842 , n38843 , n38844 , n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , 
     n38851 , n38852 , n38853 , n38854 , n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , 
     n38861 , n38862 , n38863 , n38864 , n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , 
     n38871 , n38872 , n38873 , n38874 , n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , 
     n38881 , n38882 , n38883 , n38884 , n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , 
     n38891 , n38892 , n38893 , n38894 , n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , 
     n38901 , n38902 , n38903 , n38904 , n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , 
     n38911 , n38912 , n38913 , n38914 , n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , 
     n38921 , n38922 , n38923 , n38924 , n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , 
     n38931 , n38932 , n38933 , n38934 , n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , 
     n38941 , n38942 , n38943 , n38944 , n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , 
     n38951 , n38952 , n38953 , n38954 , n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , 
     n38961 , n38962 , n38963 , n38964 , n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , 
     n38971 , n38972 , n38973 , n38974 , n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , 
     n38981 , n38982 , n38983 , n38984 , n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , 
     n38991 , n38992 , n38993 , n38994 , n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , 
     n39001 , n39002 , n39003 , n39004 , n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , 
     n39011 , n39012 , n39013 , n39014 , n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , 
     n39021 , n39022 , n39023 , n39024 , n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , 
     n39031 , n39032 , n39033 , n39034 , n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , 
     n39041 , n39042 , n39043 , n39044 , n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , 
     n39051 , n39052 , n39053 , n39054 , n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , 
     n39061 , n39062 , n39063 , n39064 , n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , 
     n39071 , n39072 , n39073 , n39074 , n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , 
     n39081 , n39082 , n39083 , n39084 , n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , 
     n39091 , n39092 , n39093 , n39094 , n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , 
     n39101 , n39102 , n39103 , n39104 , n39105 , n39106 , n39107 , n39108 , n39109 , n39110 , 
     n39111 , n39112 , n39113 , n39114 , n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , 
     n39121 , n39122 , n39123 , n39124 , n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , 
     n39131 , n39132 , n39133 , n39134 , n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , 
     n39141 , n39142 , n39143 , n39144 , n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , 
     n39151 , n39152 , n39153 , n39154 , n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , 
     n39161 , n39162 , n39163 , n39164 , n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , 
     n39171 , n39172 , n39173 , n39174 , n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , 
     n39181 , n39182 , n39183 , n39184 , n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , 
     n39191 , n39192 , n39193 , n39194 , n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , 
     n39201 , n39202 , n39203 , n39204 , n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , 
     n39211 , n39212 , n39213 , n39214 , n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , 
     n39221 , n39222 , n39223 , n39224 , n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , 
     n39231 , n39232 , n39233 , n39234 , n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , 
     n39241 , n39242 , n39243 , n39244 , n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , 
     n39251 , n39252 , n39253 , n39254 , n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , 
     n39261 , n39262 , n39263 , n39264 , n39265 , n39266 , n39267 , n39268 , n39269 , n39270 , 
     n39271 , n39272 , n39273 , n39274 , n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , 
     n39281 , n39282 , n39283 , n39284 , n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , 
     n39291 , n39292 , n39293 , n39294 , n39295 , n39296 , n39297 , n39298 , n39299 , n39300 , 
     n39301 , n39302 , n39303 , n39304 , n39305 , n39306 , n39307 , n39308 , n39309 , n39310 , 
     n39311 , n39312 , n39313 , n39314 , n39315 , n39316 , n39317 , n39318 , n39319 , n39320 , 
     n39321 , n39322 , n39323 , n39324 , n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , 
     n39331 , n39332 , n39333 , n39334 , n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , 
     n39341 , n39342 , n39343 , n39344 , n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , 
     n39351 , n39352 , n39353 , n39354 , n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , 
     n39361 , n39362 , n39363 , n39364 , n39365 , n39366 , n39367 , n39368 , n39369 , n39370 , 
     n39371 , n39372 , n39373 , n39374 , n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , 
     n39381 , n39382 , n39383 , n39384 , n39385 , n39386 , n39387 , n39388 , n39389 , n39390 , 
     n39391 , n39392 , n39393 , n39394 , n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , 
     n39401 , n39402 , n39403 , n39404 , n39405 , n39406 , n39407 , n39408 , n39409 , n39410 , 
     n39411 , n39412 , n39413 , n39414 , n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , 
     n39421 , n39422 , n39423 , n39424 , n39425 , n39426 , n39427 , n39428 , n39429 , n39430 , 
     n39431 , n39432 , n39433 , n39434 , n39435 , n39436 , n39437 , n39438 , n39439 , n39440 , 
     n39441 , n39442 , n39443 , n39444 , n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , 
     n39451 , n39452 , n39453 , n39454 , n39455 , n39456 , n39457 , n39458 , n39459 , n39460 , 
     n39461 , n39462 , n39463 , n39464 , n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , 
     n39471 , n39472 , n39473 , n39474 , n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , 
     n39481 , n39482 , n39483 , n39484 , n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , 
     n39491 , n39492 , n39493 , n39494 , n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , 
     n39501 , n39502 , n39503 , n39504 , n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , 
     n39511 , n39512 , n39513 , n39514 , n39515 , n39516 , n39517 , n39518 , n39519 , n39520 , 
     n39521 , n39522 , n39523 , n39524 , n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , 
     n39531 , n39532 , n39533 , n39534 , n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , 
     n39541 , n39542 , n39543 , n39544 , n39545 , n39546 , n39547 , n39548 , n39549 , n39550 , 
     n39551 , n39552 , n39553 , n39554 , n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , 
     n39561 , n39562 , n39563 , n39564 , n39565 , n39566 , n39567 , n39568 , n39569 , n39570 , 
     n39571 , n39572 , n39573 , n39574 , n39575 , n39576 , n39577 , n39578 , n39579 , n39580 , 
     n39581 , n39582 , n39583 , n39584 , n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , 
     n39591 , n39592 , n39593 , n39594 , n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , 
     n39601 , n39602 , n39603 , n39604 , n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , 
     n39611 , n39612 , n39613 , n39614 , n39615 , n39616 , n39617 , n39618 , n39619 , n39620 , 
     n39621 , n39622 , n39623 , n39624 , n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , 
     n39631 , n39632 , n39633 , n39634 , n39635 , n39636 , n39637 , n39638 , n39639 , n39640 , 
     n39641 , n39642 , n39643 , n39644 , n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , 
     n39651 , n39652 , n39653 , n39654 , n39655 , n39656 , n39657 , n39658 , n39659 , n39660 , 
     n39661 , n39662 , n39663 , n39664 , n39665 , n39666 , n39667 , n39668 , n39669 , n39670 , 
     n39671 , n39672 , n39673 , n39674 , n39675 , n39676 , n39677 , n39678 , n39679 , n39680 , 
     n39681 , n39682 , n39683 , n39684 , n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , 
     n39691 , n39692 , n39693 , n39694 , n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , 
     n39701 , n39702 , n39703 , n39704 , n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , 
     n39711 , n39712 , n39713 , n39714 , n39715 , n39716 , n39717 , n39718 , n39719 , n39720 , 
     n39721 , n39722 , n39723 , n39724 , n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , 
     n39731 , n39732 , n39733 , n39734 , n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , 
     n39741 , n39742 , n39743 , n39744 , n39745 , n39746 , n39747 , n39748 , n39749 , n39750 , 
     n39751 , n39752 , n39753 , n39754 , n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , 
     n39761 , n39762 , n39763 , n39764 , n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , 
     n39771 , n39772 , n39773 , n39774 , n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , 
     n39781 , n39782 , n39783 , n39784 , n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , 
     n39791 , n39792 , n39793 , n39794 , n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , 
     n39801 , n39802 , n39803 , n39804 , n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , 
     n39811 , n39812 , n39813 , n39814 , n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , 
     n39821 , n39822 , n39823 , n39824 , n39825 , n39826 , n39827 , n39828 , n39829 , n39830 , 
     n39831 , n39832 , n39833 , n39834 , n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , 
     n39841 , n39842 , n39843 , n39844 , n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , 
     n39851 , n39852 , n39853 , n39854 , n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , 
     n39861 , n39862 , n39863 , n39864 , n39865 , n39866 , n39867 , n39868 , n39869 , n39870 , 
     n39871 , n39872 , n39873 , n39874 , n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , 
     n39881 , n39882 , n39883 , n39884 , n39885 , n39886 , n39887 , n39888 , n39889 , n39890 , 
     n39891 , n39892 , n39893 , n39894 , n39895 , n39896 , n39897 , n39898 , n39899 , n39900 , 
     n39901 , n39902 , n39903 , n39904 , n39905 , n39906 , n39907 , n39908 , n39909 , n39910 , 
     n39911 , n39912 , n39913 , n39914 , n39915 , n39916 , n39917 , n39918 , n39919 , n39920 , 
     n39921 , n39922 , n39923 , n39924 , n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , 
     n39931 , n39932 , n39933 , n39934 , n39935 , n39936 , n39937 , n39938 , n39939 , n39940 , 
     n39941 , n39942 , n39943 , n39944 , n39945 , n39946 , n39947 , n39948 , n39949 , n39950 , 
     n39951 , n39952 , n39953 , n39954 , n39955 , n39956 , n39957 , n39958 , n39959 , n39960 , 
     n39961 , n39962 , n39963 , n39964 , n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , 
     n39971 , n39972 , n39973 , n39974 , n39975 , n39976 , n39977 , n39978 , n39979 , n39980 , 
     n39981 , n39982 , n39983 , n39984 , n39985 , n39986 , n39987 , n39988 , n39989 , n39990 , 
     n39991 , n39992 , n39993 , n39994 , n39995 , n39996 , n39997 , n39998 , n39999 , n40000 , 
     n40001 , n40002 , n40003 , n40004 , n40005 , n40006 , n40007 , n40008 , n40009 , n40010 , 
     n40011 , n40012 , n40013 , n40014 , n40015 , n40016 , n40017 , n40018 , n40019 , n40020 , 
     n40021 , n40022 , n40023 , n40024 , n40025 , n40026 , n40027 , n40028 , n40029 , n40030 , 
     n40031 , n40032 , n40033 , n40034 , n40035 , n40036 , n40037 , n40038 , n40039 , n40040 , 
     n40041 , n40042 , n40043 , n40044 , n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , 
     n40051 , n40052 , n40053 , n40054 , n40055 , n40056 , n40057 , n40058 , n40059 , n40060 , 
     n40061 , n40062 , n40063 , n40064 , n40065 , n40066 , n40067 , n40068 , n40069 , n40070 , 
     n40071 , n40072 , n40073 , n40074 , n40075 , n40076 , n40077 , n40078 , n40079 , n40080 , 
     n40081 , n40082 , n40083 , n40084 , n40085 , n40086 , n40087 , n40088 , n40089 , n40090 , 
     n40091 , n40092 , n40093 , n40094 , n40095 , n40096 , n40097 , n40098 , n40099 , n40100 , 
     n40101 , n40102 , n40103 , n40104 , n40105 , n40106 , n40107 , n40108 , n40109 , n40110 , 
     n40111 , n40112 , n40113 , n40114 , n40115 , n40116 , n40117 , n40118 , n40119 , n40120 , 
     n40121 , n40122 , n40123 , n40124 , n40125 , n40126 , n40127 , n40128 , n40129 , n40130 , 
     n40131 , n40132 , n40133 , n40134 , n40135 , n40136 , n40137 , n40138 , n40139 , n40140 , 
     n40141 , n40142 , n40143 , n40144 , n40145 , n40146 , n40147 , n40148 , n40149 , n40150 , 
     n40151 , n40152 , n40153 , n40154 , n40155 , n40156 , n40157 , n40158 , n40159 , n40160 , 
     n40161 , n40162 , n40163 , n40164 , n40165 , n40166 , n40167 , n40168 , n40169 , n40170 , 
     n40171 , n40172 , n40173 , n40174 , n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , 
     n40181 , n40182 , n40183 , n40184 , n40185 , n40186 , n40187 , n40188 , n40189 , n40190 , 
     n40191 , n40192 , n40193 , n40194 , n40195 , n40196 , n40197 , n40198 , n40199 , n40200 , 
     n40201 , n40202 , n40203 , n40204 , n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , 
     n40211 , n40212 , n40213 , n40214 , n40215 , n40216 , n40217 , n40218 , n40219 , n40220 , 
     n40221 , n40222 , n40223 , n40224 , n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , 
     n40231 , n40232 , n40233 , n40234 , n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , 
     n40241 , n40242 , n40243 , n40244 , n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , 
     n40251 , n40252 , n40253 , n40254 , n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , 
     n40261 , n40262 , n40263 , n40264 , n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , 
     n40271 , n40272 , n40273 , n40274 , n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , 
     n40281 , n40282 , n40283 , n40284 , n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , 
     n40291 , n40292 , n40293 , n40294 , n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , 
     n40301 , n40302 , n40303 , n40304 , n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , 
     n40311 , n40312 , n40313 , n40314 , n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , 
     n40321 , n40322 , n40323 , n40324 , n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , 
     n40331 , n40332 , n40333 , n40334 , n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , 
     n40341 , n40342 , n40343 , n40344 , n40345 , n40346 , n40347 , n40348 , n40349 , n40350 , 
     n40351 , n40352 , n40353 , n40354 , n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , 
     n40361 , n40362 , n40363 , n40364 , n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , 
     n40371 , n40372 , n40373 , n40374 , n40375 , n40376 , n40377 , n40378 , n40379 , n40380 , 
     n40381 , n40382 , n40383 , n40384 , n40385 , n40386 , n40387 , n40388 , n40389 , n40390 , 
     n40391 , n40392 , n40393 , n40394 , n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , 
     n40401 , n40402 , n40403 , n40404 , n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , 
     n40411 , n40412 , n40413 , n40414 , n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , 
     n40421 , n40422 , n40423 , n40424 , n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , 
     n40431 , n40432 , n40433 , n40434 , n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , 
     n40441 , n40442 , n40443 , n40444 , n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , 
     n40451 , n40452 , n40453 , n40454 , n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , 
     n40461 , n40462 , n40463 , n40464 , n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , 
     n40471 , n40472 , n40473 , n40474 , n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , 
     n40481 , n40482 , n40483 , n40484 , n40485 , n40486 , n40487 , n40488 , n40489 , n40490 , 
     n40491 , n40492 , n40493 , n40494 , n40495 , n40496 , n40497 , n40498 , n40499 , n40500 , 
     n40501 , n40502 , n40503 , n40504 , n40505 , n40506 , n40507 , n40508 , n40509 , n40510 , 
     n40511 , n40512 , n40513 , n40514 , n40515 , n40516 , n40517 , n40518 , n40519 , n40520 , 
     n40521 , n40522 , n40523 , n40524 , n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , 
     n40531 , n40532 , n40533 , n40534 , n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , 
     n40541 , n40542 , n40543 , n40544 , n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , 
     n40551 , n40552 , n40553 , n40554 , n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , 
     n40561 , n40562 , n40563 , n40564 , n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , 
     n40571 , n40572 , n40573 , n40574 , n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , 
     n40581 , n40582 , n40583 , n40584 , n40585 , n40586 , n40587 , n40588 , n40589 , n40590 , 
     n40591 , n40592 , n40593 , n40594 , n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , 
     n40601 , n40602 , n40603 , n40604 , n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , 
     n40611 , n40612 , n40613 , n40614 , n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , 
     n40621 , n40622 , n40623 , n40624 , n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , 
     n40631 , n40632 , n40633 , n40634 , n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , 
     n40641 , n40642 , n40643 , n40644 , n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , 
     n40651 , n40652 , n40653 , n40654 , n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , 
     n40661 , n40662 , n40663 , n40664 , n40665 , n40666 , n40667 , n40668 , n40669 , n40670 , 
     n40671 , n40672 , n40673 , n40674 , n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , 
     n40681 , n40682 , n40683 , n40684 , n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , 
     n40691 , n40692 , n40693 , n40694 , n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , 
     n40701 , n40702 , n40703 , n40704 , n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , 
     n40711 , n40712 , n40713 , n40714 , n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , 
     n40721 , n40722 , n40723 , n40724 , n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , 
     n40731 , n40732 , n40733 , n40734 , n40735 , n40736 , n40737 , n40738 , n40739 , n40740 , 
     n40741 , n40742 , n40743 , n40744 , n40745 , n40746 , n40747 , n40748 , n40749 , n40750 , 
     n40751 , n40752 , n40753 , n40754 , n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , 
     n40761 , n40762 , n40763 , n40764 , n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , 
     n40771 , n40772 , n40773 , n40774 , n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , 
     n40781 , n40782 , n40783 , n40784 , n40785 , n40786 , n40787 , n40788 , n40789 , n40790 , 
     n40791 , n40792 , n40793 , n40794 , n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , 
     n40801 , n40802 , n40803 , n40804 , n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , 
     n40811 , n40812 , n40813 , n40814 , n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , 
     n40821 , n40822 , n40823 , n40824 , n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , 
     n40831 , n40832 , n40833 , n40834 , n40835 , n40836 , n40837 , n40838 , n40839 , n40840 , 
     n40841 , n40842 , n40843 , n40844 , n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , 
     n40851 , n40852 , n40853 , n40854 , n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , 
     n40861 , n40862 , n40863 , n40864 , n40865 , n40866 , n40867 , n40868 , n40869 , n40870 , 
     n40871 , n40872 , n40873 , n40874 , n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , 
     n40881 , n40882 , n40883 , n40884 , n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , 
     n40891 , n40892 , n40893 , n40894 , n40895 , n40896 , n40897 , n40898 , n40899 , n40900 , 
     n40901 , n40902 , n40903 , n40904 , n40905 , n40906 , n40907 , n40908 , n40909 , n40910 , 
     n40911 , n40912 , n40913 , n40914 , n40915 , n40916 , n40917 , n40918 , n40919 , n40920 , 
     n40921 , n40922 , n40923 , n40924 , n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , 
     n40931 , n40932 , n40933 , n40934 , n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , 
     n40941 , n40942 , n40943 , n40944 , n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , 
     n40951 , n40952 , n40953 , n40954 , n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , 
     n40961 , n40962 , n40963 , n40964 , n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , 
     n40971 , n40972 , n40973 , n40974 , n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , 
     n40981 , n40982 , n40983 , n40984 , n40985 , n40986 , n40987 , n40988 , n40989 , n40990 , 
     n40991 , n40992 , n40993 , n40994 , n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , 
     n41001 , n41002 , n41003 , n41004 , n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , 
     n41011 , n41012 , n41013 , n41014 , n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , 
     n41021 , n41022 , n41023 , n41024 , n41025 , n41026 , n41027 , n41028 , n41029 , n41030 , 
     n41031 , n41032 , n41033 , n41034 , n41035 , n41036 , n41037 , n41038 , n41039 , n41040 , 
     n41041 , n41042 , n41043 , n41044 , n41045 , n41046 , n41047 , n41048 , n41049 , n41050 , 
     n41051 , n41052 , n41053 , n41054 , n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , 
     n41061 , n41062 , n41063 , n41064 , n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , 
     n41071 , n41072 , n41073 , n41074 , n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , 
     n41081 , n41082 , n41083 , n41084 , n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , 
     n41091 , n41092 , n41093 , n41094 , n41095 , n41096 , n41097 , n41098 , n41099 , n41100 , 
     n41101 , n41102 , n41103 , n41104 , n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , 
     n41111 , n41112 , n41113 , n41114 , n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , 
     n41121 , n41122 , n41123 , n41124 , n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , 
     n41131 , n41132 , n41133 , n41134 , n41135 , n41136 , n41137 , n41138 , n41139 , n41140 , 
     n41141 , n41142 , n41143 , n41144 , n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , 
     n41151 , n41152 , n41153 , n41154 , n41155 , n41156 , n41157 , n41158 , n41159 , n41160 , 
     n41161 , n41162 , n41163 , n41164 , n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , 
     n41171 , n41172 , n41173 , n41174 , n41175 , n41176 , n41177 , n41178 , n41179 , n41180 , 
     n41181 , n41182 , n41183 , n41184 , n41185 , n41186 , n41187 , n41188 , n41189 , n41190 , 
     n41191 , n41192 , n41193 , n41194 , n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , 
     n41201 , n41202 , n41203 , n41204 , n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , 
     n41211 , n41212 , n41213 , n41214 , n41215 , n41216 , n41217 , n41218 , n41219 , n41220 , 
     n41221 , n41222 , n41223 , n41224 , n41225 , n41226 , n41227 , n41228 , n41229 , n41230 , 
     n41231 , n41232 , n41233 , n41234 , n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , 
     n41241 , n41242 , n41243 , n41244 , n41245 , n41246 , n41247 , n41248 , n41249 , n41250 , 
     n41251 , n41252 , n41253 , n41254 , n41255 , n41256 , n41257 , n41258 , n41259 , n41260 , 
     n41261 , n41262 , n41263 , n41264 , n41265 , n41266 , n41267 , n41268 , n41269 , n41270 , 
     n41271 , n41272 , n41273 , n41274 , n41275 , n41276 , n41277 , n41278 , n41279 , n41280 , 
     n41281 , n41282 , n41283 , n41284 , n41285 , n41286 , n41287 , n41288 , n41289 , n41290 , 
     n41291 , n41292 , n41293 , n41294 , n41295 , n41296 , n41297 , n41298 , n41299 , n41300 , 
     n41301 , n41302 , n41303 , n41304 , n41305 , n41306 , n41307 , n41308 , n41309 , n41310 , 
     n41311 , n41312 , n41313 , n41314 , n41315 , n41316 , n41317 , n41318 , n41319 , n41320 , 
     n41321 , n41322 , n41323 , n41324 , n41325 , n41326 , n41327 , n41328 , n41329 , n41330 , 
     n41331 , n41332 , n41333 , n41334 , n41335 , n41336 , n41337 , n41338 , n41339 , n41340 , 
     n41341 , n41342 , n41343 , n41344 , n41345 , n41346 , n41347 , n41348 , n41349 , n41350 , 
     n41351 , n41352 , n41353 , n41354 , n41355 , n41356 , n41357 , n41358 , n41359 , n41360 , 
     n41361 , n41362 , n41363 , n41364 , n41365 , n41366 , n41367 , n41368 , n41369 , n41370 , 
     n41371 , n41372 , n41373 , n41374 , n41375 , n41376 , n41377 , n41378 , n41379 , n41380 , 
     n41381 , n41382 , n41383 , n41384 , n41385 , n41386 , n41387 , n41388 , n41389 , n41390 , 
     n41391 , n41392 , n41393 , n41394 , n41395 , n41396 , n41397 , n41398 , n41399 , n41400 , 
     n41401 , n41402 , n41403 , n41404 , n41405 , n41406 , n41407 , n41408 , n41409 , n41410 , 
     n41411 , n41412 , n41413 , n41414 , n41415 , n41416 , n41417 , n41418 , n41419 , n41420 , 
     n41421 , n41422 , n41423 , n41424 , n41425 , n41426 , n41427 , n41428 , n41429 , n41430 , 
     n41431 , n41432 , n41433 , n41434 , n41435 , n41436 , n41437 , n41438 , n41439 , n41440 , 
     n41441 , n41442 , n41443 , n41444 , n41445 , n41446 , n41447 , n41448 , n41449 , n41450 , 
     n41451 , n41452 , n41453 , n41454 , n41455 , n41456 , n41457 , n41458 , n41459 , n41460 , 
     n41461 , n41462 , n41463 , n41464 , n41465 , n41466 , n41467 , n41468 , n41469 , n41470 , 
     n41471 , n41472 , n41473 , n41474 , n41475 , n41476 , n41477 , n41478 , n41479 , n41480 , 
     n41481 , n41482 , n41483 , n41484 , n41485 , n41486 , n41487 , n41488 , n41489 , n41490 , 
     n41491 , n41492 , n41493 , n41494 , n41495 , n41496 , n41497 , n41498 , n41499 , n41500 , 
     n41501 , n41502 , n41503 , n41504 , n41505 , n41506 , n41507 , n41508 , n41509 , n41510 , 
     n41511 , n41512 , n41513 , n41514 , n41515 , n41516 , n41517 , n41518 , n41519 , n41520 , 
     n41521 , n41522 , n41523 , n41524 , n41525 , n41526 , n41527 , n41528 , n41529 , n41530 , 
     n41531 , n41532 , n41533 , n41534 , n41535 , n41536 , n41537 , n41538 , n41539 , n41540 , 
     n41541 , n41542 , n41543 , n41544 , n41545 , n41546 , n41547 , n41548 , n41549 , n41550 , 
     n41551 , n41552 , n41553 , n41554 , n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , 
     n41561 , n41562 , n41563 , n41564 , n41565 , n41566 , n41567 , n41568 , n41569 , n41570 , 
     n41571 , n41572 , n41573 , n41574 , n41575 , n41576 , n41577 , n41578 , n41579 , n41580 , 
     n41581 , n41582 , n41583 , n41584 , n41585 , n41586 , n41587 , n41588 , n41589 , n41590 , 
     n41591 , n41592 , n41593 , n41594 , n41595 , n41596 , n41597 , n41598 , n41599 , n41600 , 
     n41601 , n41602 , n41603 , n41604 , n41605 , n41606 , n41607 , n41608 , n41609 , n41610 , 
     n41611 , n41612 , n41613 , n41614 , n41615 , n41616 , n41617 , n41618 , n41619 , n41620 , 
     n41621 , n41622 , n41623 , n41624 , n41625 , n41626 , n41627 , n41628 , n41629 , n41630 , 
     n41631 , n41632 , n41633 , n41634 , n41635 , n41636 , n41637 , n41638 , n41639 , n41640 , 
     n41641 , n41642 , n41643 , n41644 , n41645 , n41646 , n41647 , n41648 , n41649 , n41650 , 
     n41651 , n41652 , n41653 , n41654 , n41655 , n41656 , n41657 , n41658 , n41659 , n41660 , 
     n41661 , n41662 , n41663 , n41664 , n41665 , n41666 , n41667 , n41668 , n41669 , n41670 , 
     n41671 , n41672 , n41673 , n41674 , n41675 , n41676 , n41677 , n41678 , n41679 , n41680 , 
     n41681 , n41682 , n41683 , n41684 , n41685 , n41686 , n41687 , n41688 , n41689 , n41690 , 
     n41691 , n41692 , n41693 , n41694 , n41695 , n41696 , n41697 , n41698 , n41699 , n41700 , 
     n41701 , n41702 , n41703 , n41704 , n41705 , n41706 , n41707 , n41708 , n41709 , n41710 , 
     n41711 , n41712 , n41713 , n41714 , n41715 , n41716 , n41717 , n41718 , n41719 , n41720 , 
     n41721 , n41722 , n41723 , n41724 , n41725 , n41726 , n41727 , n41728 , n41729 , n41730 , 
     n41731 , n41732 , n41733 , n41734 , n41735 , n41736 , n41737 , n41738 , n41739 , n41740 , 
     n41741 , n41742 , n41743 , n41744 , n41745 , n41746 , n41747 , n41748 , n41749 , n41750 , 
     n41751 , n41752 , n41753 , n41754 , n41755 , n41756 , n41757 , n41758 , n41759 , n41760 , 
     n41761 , n41762 , n41763 , n41764 , n41765 , n41766 , n41767 , n41768 , n41769 , n41770 , 
     n41771 , n41772 , n41773 , n41774 , n41775 , n41776 , n41777 , n41778 , n41779 , n41780 , 
     n41781 , n41782 , n41783 , n41784 , n41785 , n41786 , n41787 , n41788 , n41789 , n41790 , 
     n41791 , n41792 , n41793 , n41794 , n41795 , n41796 , n41797 , n41798 , n41799 , n41800 , 
     n41801 , n41802 , n41803 , n41804 , n41805 , n41806 , n41807 , n41808 , n41809 , n41810 , 
     n41811 , n41812 , n41813 , n41814 , n41815 , n41816 , n41817 , n41818 , n41819 , n41820 , 
     n41821 , n41822 , n41823 , n41824 , n41825 , n41826 , n41827 , n41828 , n41829 , n41830 , 
     n41831 , n41832 , n41833 , n41834 , n41835 , n41836 , n41837 , n41838 , n41839 , n41840 , 
     n41841 , n41842 , n41843 , n41844 , n41845 , n41846 , n41847 , n41848 , n41849 , n41850 , 
     n41851 , n41852 , n41853 , n41854 , n41855 , n41856 , n41857 , n41858 , n41859 , n41860 , 
     n41861 , n41862 , n41863 , n41864 , n41865 , n41866 , n41867 , n41868 , n41869 , n41870 , 
     n41871 , n41872 , n41873 , n41874 , n41875 , n41876 , n41877 , n41878 , n41879 , n41880 , 
     n41881 , n41882 , n41883 , n41884 , n41885 , n41886 , n41887 , n41888 , n41889 , n41890 , 
     n41891 , n41892 , n41893 , n41894 , n41895 , n41896 , n41897 , n41898 , n41899 , n41900 , 
     n41901 , n41902 , n41903 , n41904 , n41905 , n41906 , n41907 , n41908 , n41909 , n41910 , 
     n41911 , n41912 , n41913 , n41914 , n41915 , n41916 , n41917 , n41918 , n41919 , n41920 , 
     n41921 , n41922 , n41923 , n41924 , n41925 , n41926 , n41927 , n41928 , n41929 , n41930 , 
     n41931 , n41932 , n41933 , n41934 , n41935 , n41936 , n41937 , n41938 , n41939 , n41940 , 
     n41941 , n41942 , n41943 , n41944 , n41945 , n41946 , n41947 , n41948 , n41949 , n41950 , 
     n41951 , n41952 , n41953 , n41954 , n41955 , n41956 , n41957 , n41958 , n41959 , n41960 , 
     n41961 , n41962 , n41963 , n41964 , n41965 , n41966 , n41967 , n41968 , n41969 , n41970 , 
     n41971 , n41972 , n41973 , n41974 , n41975 , n41976 , n41977 , n41978 , n41979 , n41980 , 
     n41981 , n41982 , n41983 , n41984 , n41985 , n41986 , n41987 , n41988 , n41989 , n41990 , 
     n41991 , n41992 , n41993 , n41994 , n41995 , n41996 , n41997 , n41998 , n41999 , n42000 , 
     n42001 , n42002 , n42003 , n42004 , n42005 , n42006 , n42007 , n42008 , n42009 , n42010 , 
     n42011 , n42012 , n42013 , n42014 , n42015 , n42016 , n42017 , n42018 , n42019 , n42020 , 
     n42021 , n42022 , n42023 , n42024 , n42025 , n42026 , n42027 , n42028 , n42029 , n42030 , 
     n42031 , n42032 , n42033 , n42034 , n42035 , n42036 , n42037 , n42038 , n42039 , n42040 , 
     n42041 , n42042 , n42043 , n42044 , n42045 , n42046 , n42047 , n42048 , n42049 , n42050 , 
     n42051 , n42052 , n42053 , n42054 , n42055 , n42056 , n42057 , n42058 , n42059 , n42060 , 
     n42061 , n42062 , n42063 , n42064 , n42065 , n42066 , n42067 , n42068 , n42069 , n42070 , 
     n42071 , n42072 , n42073 , n42074 , n42075 , n42076 , n42077 , n42078 , n42079 , n42080 , 
     n42081 , n42082 , n42083 , n42084 , n42085 , n42086 , n42087 , n42088 , n42089 , n42090 , 
     n42091 , n42092 , n42093 , n42094 , n42095 , n42096 , n42097 , n42098 , n42099 , n42100 , 
     n42101 , n42102 , n42103 , n42104 , n42105 , n42106 , n42107 , n42108 , n42109 , n42110 , 
     n42111 , n42112 , n42113 , n42114 , n42115 , n42116 , n42117 , n42118 , n42119 , n42120 , 
     n42121 , n42122 , n42123 , n42124 , n42125 , n42126 , n42127 , n42128 , n42129 , n42130 , 
     n42131 , n42132 , n42133 , n42134 , n42135 , n42136 , n42137 , n42138 , n42139 , n42140 , 
     n42141 , n42142 , n42143 , n42144 , n42145 , n42146 , n42147 , n42148 , n42149 , n42150 , 
     n42151 , n42152 , n42153 , n42154 , n42155 , n42156 , n42157 , n42158 , n42159 , n42160 , 
     n42161 , n42162 , n42163 , n42164 , n42165 , n42166 , n42167 , n42168 , n42169 , n42170 , 
     n42171 , n42172 , n42173 , n42174 , n42175 , n42176 , n42177 , n42178 , n42179 , n42180 , 
     n42181 , n42182 , n42183 , n42184 , n42185 , n42186 , n42187 , n42188 , n42189 , n42190 , 
     n42191 , n42192 , n42193 , n42194 , n42195 , n42196 , n42197 , n42198 , n42199 , n42200 , 
     n42201 , n42202 , n42203 , n42204 , n42205 , n42206 , n42207 , n42208 , n42209 , n42210 , 
     n42211 , n42212 , n42213 , n42214 , n42215 , n42216 , n42217 , n42218 , n42219 , n42220 , 
     n42221 , n42222 , n42223 , n42224 , n42225 , n42226 , n42227 , n42228 , n42229 , n42230 , 
     n42231 , n42232 , n42233 , n42234 , n42235 , n42236 , n42237 , n42238 , n42239 , n42240 , 
     n42241 , n42242 , n42243 , n42244 , n42245 , n42246 , n42247 , n42248 , n42249 , n42250 , 
     n42251 , n42252 , n42253 , n42254 , n42255 , n42256 , n42257 , n42258 , n42259 , n42260 , 
     n42261 , n42262 , n42263 , n42264 , n42265 , n42266 , n42267 , n42268 , n42269 , n42270 , 
     n42271 , n42272 , n42273 , n42274 , n42275 , n42276 , n42277 , n42278 , n42279 , n42280 , 
     n42281 , n42282 , n42283 , n42284 , n42285 , n42286 , n42287 , n42288 , n42289 , n42290 , 
     n42291 , n42292 , n42293 , n42294 , n42295 , n42296 , n42297 , n42298 , n42299 , n42300 , 
     n42301 , n42302 , n42303 , n42304 , n42305 , n42306 , n42307 , n42308 , n42309 , n42310 , 
     n42311 , n42312 , n42313 , n42314 , n42315 , n42316 , n42317 , n42318 , n42319 , n42320 , 
     n42321 , n42322 , n42323 , n42324 , n42325 , n42326 , n42327 , n42328 , n42329 , n42330 , 
     n42331 , n42332 , n42333 , n42334 , n42335 , n42336 , n42337 , n42338 , n42339 , n42340 , 
     n42341 , n42342 , n42343 , n42344 , n42345 , n42346 , n42347 , n42348 , n42349 , n42350 , 
     n42351 , n42352 , n42353 , n42354 , n42355 , n42356 , n42357 , n42358 , n42359 , n42360 , 
     n42361 , n42362 , n42363 , n42364 , n42365 , n42366 , n42367 , n42368 , n42369 , n42370 , 
     n42371 , n42372 , n42373 , n42374 , n42375 , n42376 , n42377 , n42378 , n42379 , n42380 , 
     n42381 , n42382 , n42383 , n42384 , n42385 , n42386 , n42387 , n42388 , n42389 , n42390 , 
     n42391 , n42392 , n42393 , n42394 , n42395 , n42396 , n42397 , n42398 , n42399 , n42400 , 
     n42401 , n42402 , n42403 , n42404 , n42405 , n42406 , n42407 , n42408 , n42409 , n42410 , 
     n42411 , n42412 , n42413 , n42414 , n42415 , n42416 , n42417 , n42418 , n42419 , n42420 , 
     n42421 , n42422 , n42423 , n42424 , n42425 , n42426 , n42427 , n42428 , n42429 , n42430 , 
     n42431 , n42432 , n42433 , n42434 , n42435 , n42436 , n42437 , n42438 , n42439 , n42440 , 
     n42441 , n42442 , n42443 , n42444 , n42445 , n42446 , n42447 , n42448 , n42449 , n42450 , 
     n42451 , n42452 , n42453 , n42454 , n42455 , n42456 , n42457 , n42458 , n42459 , n42460 , 
     n42461 , n42462 , n42463 , n42464 , n42465 , n42466 , n42467 , n42468 , n42469 , n42470 , 
     n42471 , n42472 , n42473 , n42474 , n42475 , n42476 , n42477 , n42478 , n42479 , n42480 , 
     n42481 , n42482 , n42483 , n42484 , n42485 , n42486 , n42487 , n42488 , n42489 , n42490 , 
     n42491 , n42492 , n42493 , n42494 , n42495 , n42496 , n42497 , n42498 , n42499 , n42500 , 
     n42501 , n42502 , n42503 , n42504 , n42505 , n42506 , n42507 , n42508 , n42509 , n42510 , 
     n42511 , n42512 , n42513 , n42514 , n42515 , n42516 , n42517 , n42518 , n42519 , n42520 , 
     n42521 , n42522 , n42523 , n42524 , n42525 , n42526 , n42527 , n42528 , n42529 , n42530 , 
     n42531 , n42532 , n42533 , n42534 , n42535 , n42536 , n42537 , n42538 , n42539 , n42540 , 
     n42541 , n42542 , n42543 , n42544 , n42545 , n42546 , n42547 , n42548 , n42549 , n42550 , 
     n42551 , n42552 , n42553 , n42554 , n42555 , n42556 , n42557 , n42558 , n42559 , n42560 , 
     n42561 , n42562 , n42563 , n42564 , n42565 , n42566 , n42567 , n42568 , n42569 , n42570 , 
     n42571 , n42572 , n42573 , n42574 , n42575 , n42576 , n42577 , n42578 , n42579 , n42580 , 
     n42581 , n42582 , n42583 , n42584 , n42585 , n42586 , n42587 , n42588 , n42589 , n42590 , 
     n42591 , n42592 , n42593 , n42594 , n42595 , n42596 , n42597 , n42598 , n42599 , n42600 , 
     n42601 , n42602 , n42603 , n42604 , n42605 , n42606 , n42607 , n42608 , n42609 , n42610 , 
     n42611 , n42612 , n42613 , n42614 , n42615 , n42616 , n42617 , n42618 , n42619 , n42620 , 
     n42621 , n42622 , n42623 , n42624 , n42625 , n42626 , n42627 , n42628 , n42629 , n42630 , 
     n42631 , n42632 , n42633 , n42634 , n42635 , n42636 , n42637 , n42638 , n42639 , n42640 , 
     n42641 , n42642 , n42643 , n42644 , n42645 , n42646 , n42647 , n42648 , n42649 , n42650 , 
     n42651 , n42652 , n42653 , n42654 , n42655 , n42656 , n42657 , n42658 , n42659 , n42660 , 
     n42661 , n42662 , n42663 , n42664 , n42665 , n42666 , n42667 , n42668 , n42669 , n42670 , 
     n42671 , n42672 , n42673 , n42674 , n42675 , n42676 , n42677 , n42678 , n42679 , n42680 , 
     n42681 , n42682 , n42683 , n42684 , n42685 , n42686 , n42687 , n42688 , n42689 , n42690 , 
     n42691 , n42692 , n42693 , n42694 , n42695 , n42696 , n42697 , n42698 , n42699 , n42700 , 
     n42701 , n42702 , n42703 , n42704 , n42705 , n42706 , n42707 , n42708 , n42709 , n42710 , 
     n42711 , n42712 , n42713 , n42714 , n42715 , n42716 , n42717 , n42718 , n42719 , n42720 , 
     n42721 , n42722 , n42723 , n42724 , n42725 , n42726 , n42727 , n42728 , n42729 , n42730 , 
     n42731 , n42732 , n42733 , n42734 , n42735 , n42736 , n42737 , n42738 , n42739 , n42740 , 
     n42741 , n42742 , n42743 , n42744 , n42745 , n42746 , n42747 , n42748 , n42749 , n42750 , 
     n42751 , n42752 , n42753 , n42754 , n42755 , n42756 , n42757 , n42758 , n42759 , n42760 , 
     n42761 , n42762 , n42763 , n42764 , n42765 , n42766 , n42767 , n42768 , n42769 , n42770 , 
     n42771 , n42772 , n42773 , n42774 , n42775 , n42776 , n42777 , n42778 , n42779 , n42780 , 
     n42781 , n42782 , n42783 , n42784 , n42785 , n42786 , n42787 , n42788 , n42789 , n42790 , 
     n42791 , n42792 , n42793 , n42794 , n42795 , n42796 , n42797 , n42798 , n42799 , n42800 , 
     n42801 , n42802 , n42803 , n42804 , n42805 , n42806 , n42807 , n42808 , n42809 , n42810 , 
     n42811 , n42812 , n42813 , n42814 , n42815 , n42816 , n42817 , n42818 , n42819 , n42820 , 
     n42821 , n42822 , n42823 , n42824 , n42825 , n42826 , n42827 , n42828 , n42829 , n42830 , 
     n42831 , n42832 , n42833 , n42834 , n42835 , n42836 , n42837 , n42838 , n42839 , n42840 , 
     n42841 , n42842 , n42843 , n42844 , n42845 , n42846 , n42847 , n42848 , n42849 , n42850 , 
     n42851 , n42852 , n42853 , n42854 , n42855 , n42856 , n42857 , n42858 , n42859 , n42860 , 
     n42861 , n42862 , n42863 , n42864 , n42865 , n42866 , n42867 , n42868 , n42869 , n42870 , 
     n42871 , n42872 , n42873 , n42874 , n42875 , n42876 , n42877 , n42878 , n42879 , n42880 , 
     n42881 , n42882 , n42883 , n42884 , n42885 , n42886 , n42887 , n42888 , n42889 , n42890 , 
     n42891 , n42892 , n42893 , n42894 , n42895 , n42896 , n42897 , n42898 , n42899 , n42900 , 
     n42901 , n42902 , n42903 , n42904 , n42905 , n42906 , n42907 , n42908 , n42909 , n42910 , 
     n42911 , n42912 , n42913 , n42914 , n42915 , n42916 , n42917 , n42918 , n42919 , n42920 , 
     n42921 , n42922 , n42923 , n42924 , n42925 , n42926 , n42927 , n42928 , n42929 , n42930 , 
     n42931 , n42932 , n42933 , n42934 , n42935 , n42936 , n42937 , n42938 , n42939 , n42940 , 
     n42941 , n42942 , n42943 , n42944 , n42945 , n42946 , n42947 , n42948 , n42949 , n42950 , 
     n42951 , n42952 , n42953 , n42954 , n42955 , n42956 , n42957 , n42958 , n42959 , n42960 , 
     n42961 , n42962 , n42963 , n42964 , n42965 , n42966 , n42967 , n42968 , n42969 , n42970 , 
     n42971 , n42972 , n42973 , n42974 , n42975 , n42976 , n42977 , n42978 , n42979 , n42980 , 
     n42981 , n42982 , n42983 , n42984 , n42985 , n42986 , n42987 , n42988 , n42989 , n42990 , 
     n42991 , n42992 , n42993 , n42994 , n42995 , n42996 , n42997 , n42998 , n42999 , n43000 , 
     n43001 , n43002 , n43003 , n43004 , n43005 , n43006 , n43007 , n43008 , n43009 , n43010 , 
     n43011 , n43012 , n43013 , n43014 , n43015 , n43016 , n43017 , n43018 , n43019 , n43020 , 
     n43021 , n43022 , n43023 , n43024 , n43025 , n43026 , n43027 , n43028 , n43029 , n43030 , 
     n43031 , n43032 , n43033 , n43034 , n43035 , n43036 , n43037 , n43038 , n43039 , n43040 , 
     n43041 , n43042 , n43043 , n43044 , n43045 , n43046 , n43047 , n43048 , n43049 , n43050 , 
     n43051 , n43052 , n43053 , n43054 , n43055 , n43056 , n43057 , n43058 , n43059 , n43060 , 
     n43061 , n43062 , n43063 , n43064 , n43065 , n43066 , n43067 , n43068 , n43069 , n43070 , 
     n43071 , n43072 , n43073 , n43074 , n43075 , n43076 , n43077 , n43078 , n43079 , n43080 , 
     n43081 , n43082 , n43083 , n43084 , n43085 , n43086 , n43087 , n43088 , n43089 , n43090 , 
     n43091 , n43092 , n43093 , n43094 , n43095 , n43096 , n43097 , n43098 , n43099 , n43100 , 
     n43101 , n43102 , n43103 , n43104 , n43105 , n43106 , n43107 , n43108 , n43109 , n43110 , 
     n43111 , n43112 , n43113 , n43114 , n43115 , n43116 , n43117 , n43118 , n43119 , n43120 , 
     n43121 , n43122 , n43123 , n43124 , n43125 , n43126 , n43127 , n43128 , n43129 , n43130 , 
     n43131 , n43132 , n43133 , n43134 , n43135 , n43136 , n43137 , n43138 , n43139 , n43140 , 
     n43141 , n43142 , n43143 , n43144 , n43145 , n43146 , n43147 , n43148 , n43149 , n43150 , 
     n43151 , n43152 , n43153 , n43154 , n43155 , n43156 , n43157 , n43158 , n43159 , n43160 , 
     n43161 , n43162 , n43163 , n43164 , n43165 , n43166 , n43167 , n43168 , n43169 , n43170 , 
     n43171 , n43172 , n43173 , n43174 , n43175 , n43176 , n43177 , n43178 , n43179 , n43180 , 
     n43181 , n43182 , n43183 , n43184 , n43185 , n43186 , n43187 , n43188 , n43189 , n43190 , 
     n43191 , n43192 , n43193 , n43194 , n43195 , n43196 , n43197 , n43198 , n43199 , n43200 , 
     n43201 , n43202 , n43203 , n43204 , n43205 , n43206 , n43207 , n43208 , n43209 , n43210 , 
     n43211 , n43212 , n43213 , n43214 , n43215 , n43216 , n43217 , n43218 , n43219 , n43220 , 
     n43221 , n43222 , n43223 , n43224 , n43225 , n43226 , n43227 , n43228 , n43229 , n43230 , 
     n43231 , n43232 , n43233 , n43234 , n43235 , n43236 , n43237 , n43238 , n43239 , n43240 , 
     n43241 , n43242 , n43243 , n43244 , n43245 , n43246 , n43247 , n43248 , n43249 , n43250 , 
     n43251 , n43252 , n43253 , n43254 , n43255 , n43256 , n43257 , n43258 , n43259 , n43260 , 
     n43261 , n43262 , n43263 , n43264 , n43265 , n43266 , n43267 , n43268 , n43269 , n43270 , 
     n43271 , n43272 , n43273 , n43274 , n43275 , n43276 , n43277 , n43278 , n43279 , n43280 , 
     n43281 , n43282 , n43283 , n43284 , n43285 , n43286 , n43287 , n43288 , n43289 , n43290 , 
     n43291 , n43292 , n43293 , n43294 , n43295 , n43296 , n43297 , n43298 , n43299 , n43300 , 
     n43301 , n43302 , n43303 , n43304 , n43305 , n43306 , n43307 , n43308 , n43309 , n43310 , 
     n43311 , n43312 , n43313 , n43314 , n43315 , n43316 , n43317 , n43318 , n43319 , n43320 , 
     n43321 , n43322 , n43323 , n43324 , n43325 , n43326 , n43327 , n43328 , n43329 , n43330 , 
     n43331 , n43332 , n43333 , n43334 , n43335 , n43336 , n43337 , n43338 , n43339 , n43340 , 
     n43341 , n43342 , n43343 , n43344 , n43345 , n43346 , n43347 , n43348 , n43349 , n43350 , 
     n43351 , n43352 , n43353 , n43354 , n43355 , n43356 , n43357 , n43358 , n43359 , n43360 , 
     n43361 , n43362 , n43363 , n43364 , n43365 , n43366 , n43367 , n43368 , n43369 , n43370 , 
     n43371 , n43372 , n43373 , n43374 , n43375 , n43376 , n43377 , n43378 , n43379 , n43380 , 
     n43381 , n43382 , n43383 , n43384 , n43385 , n43386 , n43387 , n43388 , n43389 , n43390 , 
     n43391 , n43392 , n43393 , n43394 , n43395 , n43396 , n43397 , n43398 , n43399 , n43400 , 
     n43401 , n43402 , n43403 , n43404 , n43405 , n43406 , n43407 , n43408 , n43409 , n43410 , 
     n43411 , n43412 , n43413 , n43414 , n43415 , n43416 , n43417 , n43418 , n43419 , n43420 , 
     n43421 , n43422 , n43423 , n43424 , n43425 , n43426 , n43427 , n43428 , n43429 , n43430 , 
     n43431 , n43432 , n43433 , n43434 , n43435 , n43436 , n43437 , n43438 , n43439 , n43440 , 
     n43441 , n43442 , n43443 , n43444 , n43445 , n43446 , n43447 , n43448 , n43449 , n43450 , 
     n43451 , n43452 , n43453 , n43454 , n43455 , n43456 , n43457 , n43458 , n43459 , n43460 , 
     n43461 , n43462 , n43463 , n43464 , n43465 , n43466 , n43467 , n43468 , n43469 , n43470 , 
     n43471 , n43472 , n43473 , n43474 , n43475 , n43476 , n43477 , n43478 , n43479 , n43480 , 
     n43481 , n43482 , n43483 , n43484 , n43485 , n43486 , n43487 , n43488 , n43489 , n43490 , 
     n43491 , n43492 , n43493 , n43494 , n43495 , n43496 , n43497 , n43498 , n43499 , n43500 , 
     n43501 , n43502 , n43503 , n43504 , n43505 , n43506 , n43507 , n43508 , n43509 , n43510 , 
     n43511 , n43512 , n43513 , n43514 , n43515 , n43516 , n43517 , n43518 , n43519 , n43520 , 
     n43521 , n43522 , n43523 , n43524 , n43525 , n43526 , n43527 , n43528 , n43529 , n43530 , 
     n43531 , n43532 , n43533 , n43534 , n43535 , n43536 , n43537 , n43538 , n43539 , n43540 , 
     n43541 , n43542 , n43543 , n43544 , n43545 , n43546 , n43547 , n43548 , n43549 , n43550 , 
     n43551 , n43552 , n43553 , n43554 , n43555 , n43556 , n43557 , n43558 , n43559 , n43560 , 
     n43561 , n43562 , n43563 , n43564 , n43565 , n43566 , n43567 , n43568 , n43569 , n43570 , 
     n43571 , n43572 , n43573 , n43574 , n43575 , n43576 , n43577 , n43578 , n43579 , n43580 , 
     n43581 , n43582 , n43583 , n43584 , n43585 , n43586 , n43587 , n43588 , n43589 , n43590 , 
     n43591 , n43592 , n43593 , n43594 , n43595 , n43596 , n43597 , n43598 , n43599 , n43600 , 
     n43601 , n43602 , n43603 , n43604 , n43605 , n43606 , n43607 , n43608 , n43609 , n43610 , 
     n43611 , n43612 , n43613 , n43614 , n43615 , n43616 , n43617 , n43618 , n43619 , n43620 , 
     n43621 , n43622 , n43623 , n43624 , n43625 , n43626 , n43627 , n43628 , n43629 , n43630 , 
     n43631 , n43632 , n43633 , n43634 , n43635 , n43636 , n43637 , n43638 , n43639 , n43640 , 
     n43641 , n43642 , n43643 , n43644 , n43645 , n43646 , n43647 , n43648 , n43649 , n43650 , 
     n43651 , n43652 , n43653 , n43654 , n43655 , n43656 , n43657 , n43658 , n43659 , n43660 , 
     n43661 , n43662 , n43663 , n43664 , n43665 , n43666 , n43667 , n43668 , n43669 , n43670 , 
     n43671 , n43672 , n43673 , n43674 , n43675 , n43676 , n43677 , n43678 , n43679 , n43680 , 
     n43681 , n43682 , n43683 , n43684 , n43685 , n43686 , n43687 , n43688 , n43689 , n43690 , 
     n43691 , n43692 , n43693 , n43694 , n43695 , n43696 , n43697 , n43698 , n43699 , n43700 , 
     n43701 , n43702 , n43703 , n43704 , n43705 , n43706 , n43707 , n43708 , n43709 , n43710 , 
     n43711 , n43712 , n43713 , n43714 , n43715 , n43716 , n43717 , n43718 , n43719 , n43720 , 
     n43721 , n43722 , n43723 , n43724 , n43725 , n43726 , n43727 , n43728 , n43729 , n43730 , 
     n43731 , n43732 , n43733 , n43734 , n43735 , n43736 , n43737 , n43738 , n43739 , n43740 , 
     n43741 , n43742 , n43743 , n43744 , n43745 , n43746 , n43747 , n43748 , n43749 , n43750 , 
     n43751 , n43752 , n43753 , n43754 , n43755 , n43756 , n43757 , n43758 , n43759 , n43760 , 
     n43761 , n43762 , n43763 , n43764 , n43765 , n43766 , n43767 , n43768 , n43769 , n43770 , 
     n43771 , n43772 , n43773 , n43774 , n43775 , n43776 , n43777 , n43778 , n43779 , n43780 , 
     n43781 , n43782 , n43783 , n43784 , n43785 , n43786 , n43787 , n43788 , n43789 , n43790 , 
     n43791 , n43792 , n43793 , n43794 , n43795 , n43796 , n43797 , n43798 , n43799 , n43800 , 
     n43801 , n43802 , n43803 , n43804 , n43805 , n43806 , n43807 , n43808 , n43809 , n43810 , 
     n43811 , n43812 , n43813 , n43814 , n43815 , n43816 , n43817 , n43818 , n43819 , n43820 , 
     n43821 , n43822 , n43823 , n43824 , n43825 , n43826 , n43827 , n43828 , n43829 , n43830 , 
     n43831 , n43832 , n43833 , n43834 , n43835 , n43836 , n43837 , n43838 , n43839 , n43840 , 
     n43841 , n43842 , n43843 , n43844 , n43845 , n43846 , n43847 , n43848 , n43849 , n43850 , 
     n43851 , n43852 , n43853 , n43854 , n43855 , n43856 , n43857 , n43858 , n43859 , n43860 , 
     n43861 , n43862 , n43863 , n43864 , n43865 , n43866 , n43867 , n43868 , n43869 , n43870 , 
     n43871 , n43872 , n43873 , n43874 , n43875 , n43876 , n43877 , n43878 , n43879 , n43880 , 
     n43881 , n43882 , n43883 , n43884 , n43885 , n43886 , n43887 , n43888 , n43889 , n43890 , 
     n43891 , n43892 , n43893 , n43894 , n43895 , n43896 , n43897 , n43898 , n43899 , n43900 , 
     n43901 , n43902 , n43903 , n43904 , n43905 , n43906 , n43907 , n43908 , n43909 , n43910 , 
     n43911 , n43912 , n43913 , n43914 , n43915 , n43916 , n43917 , n43918 , n43919 , n43920 , 
     n43921 , n43922 , n43923 , n43924 , n43925 , n43926 , n43927 , n43928 , n43929 , n43930 , 
     n43931 , n43932 , n43933 , n43934 , n43935 , n43936 , n43937 , n43938 , n43939 , n43940 , 
     n43941 , n43942 , n43943 , n43944 , n43945 , n43946 , n43947 , n43948 , n43949 , n43950 , 
     n43951 , n43952 , n43953 , n43954 , n43955 , n43956 , n43957 , n43958 , n43959 , n43960 , 
     n43961 , n43962 , n43963 , n43964 , n43965 , n43966 , n43967 , n43968 , n43969 , n43970 , 
     n43971 , n43972 , n43973 , n43974 , n43975 , n43976 , n43977 , n43978 , n43979 , n43980 , 
     n43981 , n43982 , n43983 , n43984 , n43985 , n43986 , n43987 , n43988 , n43989 , n43990 , 
     n43991 , n43992 , n43993 , n43994 , n43995 , n43996 , n43997 , n43998 , n43999 , n44000 , 
     n44001 , n44002 , n44003 , n44004 , n44005 , n44006 , n44007 , n44008 , n44009 , n44010 , 
     n44011 , n44012 , n44013 , n44014 , n44015 , n44016 , n44017 , n44018 , n44019 , n44020 , 
     n44021 , n44022 , n44023 , n44024 , n44025 , n44026 , n44027 , n44028 , n44029 , n44030 , 
     n44031 , n44032 , n44033 , n44034 , n44035 , n44036 , n44037 , n44038 , n44039 , n44040 , 
     n44041 , n44042 , n44043 , n44044 , n44045 , n44046 , n44047 , n44048 , n44049 , n44050 , 
     n44051 , n44052 , n44053 , n44054 , n44055 , n44056 , n44057 , n44058 , n44059 , n44060 , 
     n44061 , n44062 , n44063 , n44064 , n44065 , n44066 , n44067 , n44068 , n44069 , n44070 , 
     n44071 , n44072 , n44073 , n44074 , n44075 , n44076 , n44077 , n44078 , n44079 , n44080 , 
     n44081 , n44082 , n44083 , n44084 , n44085 , n44086 , n44087 , n44088 , n44089 , n44090 , 
     n44091 , n44092 , n44093 , n44094 , n44095 , n44096 , n44097 , n44098 , n44099 , n44100 , 
     n44101 , n44102 , n44103 , n44104 , n44105 , n44106 , n44107 , n44108 , n44109 , n44110 , 
     n44111 , n44112 , n44113 , n44114 , n44115 , n44116 , n44117 , n44118 , n44119 , n44120 , 
     n44121 , n44122 , n44123 , n44124 , n44125 , n44126 , n44127 , n44128 , n44129 , n44130 , 
     n44131 , n44132 , n44133 , n44134 , n44135 , n44136 , n44137 , n44138 , n44139 , n44140 , 
     n44141 , n44142 , n44143 , n44144 , n44145 , n44146 , n44147 , n44148 , n44149 , n44150 , 
     n44151 , n44152 , n44153 , n44154 , n44155 , n44156 , n44157 , n44158 , n44159 , n44160 , 
     n44161 , n44162 , n44163 , n44164 , n44165 , n44166 , n44167 , n44168 , n44169 , n44170 , 
     n44171 , n44172 , n44173 , n44174 , n44175 , n44176 , n44177 , n44178 , n44179 , n44180 , 
     n44181 , n44182 , n44183 , n44184 , n44185 , n44186 , n44187 , n44188 , n44189 , n44190 , 
     n44191 , n44192 , n44193 , n44194 , n44195 , n44196 , n44197 , n44198 , n44199 , n44200 , 
     n44201 , n44202 , n44203 , n44204 , n44205 , n44206 , n44207 , n44208 , n44209 , n44210 , 
     n44211 , n44212 , n44213 , n44214 , n44215 , n44216 , n44217 , n44218 , n44219 , n44220 , 
     n44221 , n44222 , n44223 , n44224 , n44225 , n44226 , n44227 , n44228 , n44229 , n44230 , 
     n44231 , n44232 , n44233 , n44234 , n44235 , n44236 , n44237 , n44238 , n44239 , n44240 , 
     n44241 , n44242 , n44243 , n44244 , n44245 , n44246 , n44247 , n44248 , n44249 , n44250 , 
     n44251 , n44252 , n44253 , n44254 , n44255 , n44256 , n44257 , n44258 , n44259 , n44260 , 
     n44261 , n44262 , n44263 , n44264 , n44265 , n44266 , n44267 , n44268 , n44269 , n44270 , 
     n44271 , n44272 , n44273 , n44274 , n44275 , n44276 , n44277 , n44278 , n44279 , n44280 , 
     n44281 , n44282 , n44283 , n44284 , n44285 , n44286 , n44287 , n44288 , n44289 , n44290 , 
     n44291 , n44292 , n44293 , n44294 , n44295 , n44296 , n44297 , n44298 , n44299 , n44300 , 
     n44301 , n44302 , n44303 , n44304 , n44305 , n44306 , n44307 , n44308 , n44309 , n44310 , 
     n44311 , n44312 , n44313 , n44314 , n44315 , n44316 , n44317 , n44318 , n44319 , n44320 , 
     n44321 , n44322 , n44323 , n44324 , n44325 , n44326 , n44327 , n44328 , n44329 , n44330 , 
     n44331 , n44332 , n44333 , n44334 , n44335 , n44336 , n44337 , n44338 , n44339 , n44340 , 
     n44341 , n44342 , n44343 , n44344 , n44345 , n44346 , n44347 , n44348 , n44349 , n44350 , 
     n44351 , n44352 , n44353 , n44354 , n44355 , n44356 , n44357 , n44358 , n44359 , n44360 , 
     n44361 , n44362 , n44363 , n44364 , n44365 , n44366 , n44367 , n44368 , n44369 , n44370 , 
     n44371 , n44372 , n44373 , n44374 , n44375 , n44376 , n44377 , n44378 , n44379 , n44380 , 
     n44381 , n44382 , n44383 , n44384 , n44385 , n44386 , n44387 , n44388 , n44389 , n44390 , 
     n44391 , n44392 , n44393 , n44394 , n44395 , n44396 , n44397 , n44398 , n44399 , n44400 , 
     n44401 , n44402 , n44403 , n44404 , n44405 , n44406 , n44407 , n44408 , n44409 , n44410 , 
     n44411 , n44412 , n44413 , n44414 , n44415 , n44416 , n44417 , n44418 , n44419 , n44420 , 
     n44421 , n44422 , n44423 , n44424 , n44425 , n44426 , n44427 , n44428 , n44429 , n44430 , 
     n44431 , n44432 , n44433 , n44434 , n44435 , n44436 , n44437 , n44438 , n44439 , n44440 , 
     n44441 , n44442 , n44443 , n44444 , n44445 , n44446 , n44447 , n44448 , n44449 , n44450 , 
     n44451 , n44452 , n44453 , n44454 , n44455 , n44456 , n44457 , n44458 , n44459 , n44460 , 
     n44461 , n44462 , n44463 , n44464 , n44465 , n44466 , n44467 , n44468 , n44469 , n44470 , 
     n44471 , n44472 , n44473 , n44474 , n44475 , n44476 , n44477 , n44478 , n44479 , n44480 , 
     n44481 , n44482 , n44483 , n44484 , n44485 , n44486 , n44487 , n44488 , n44489 , n44490 , 
     n44491 , n44492 , n44493 , n44494 , n44495 , n44496 , n44497 , n44498 , n44499 , n44500 , 
     n44501 , n44502 , n44503 , n44504 , n44505 , n44506 , n44507 , n44508 , n44509 , n44510 , 
     n44511 , n44512 , n44513 , n44514 , n44515 , n44516 , n44517 , n44518 , n44519 , n44520 , 
     n44521 , n44522 , n44523 , n44524 , n44525 , n44526 , n44527 , n44528 , n44529 , n44530 , 
     n44531 , n44532 , n44533 , n44534 , n44535 , n44536 , n44537 , n44538 , n44539 , n44540 , 
     n44541 , n44542 , n44543 , n44544 , n44545 , n44546 , n44547 , n44548 , n44549 , n44550 , 
     n44551 , n44552 , n44553 , n44554 , n44555 , n44556 , n44557 , n44558 , n44559 , n44560 , 
     n44561 , n44562 , n44563 , n44564 , n44565 , n44566 , n44567 , n44568 , n44569 , n44570 , 
     n44571 , n44572 , n44573 , n44574 , n44575 , n44576 , n44577 , n44578 , n44579 , n44580 , 
     n44581 , n44582 , n44583 , n44584 , n44585 , n44586 , n44587 , n44588 , n44589 , n44590 , 
     n44591 , n44592 , n44593 , n44594 , n44595 , n44596 , n44597 , n44598 , n44599 , n44600 , 
     n44601 , n44602 , n44603 , n44604 , n44605 , n44606 , n44607 , n44608 , n44609 , n44610 , 
     n44611 , n44612 , n44613 , n44614 , n44615 , n44616 , n44617 , n44618 , n44619 , n44620 , 
     n44621 , n44622 , n44623 , n44624 , n44625 , n44626 , n44627 , n44628 , n44629 , n44630 , 
     n44631 , n44632 , n44633 , n44634 , n44635 , n44636 , n44637 , n44638 , n44639 , n44640 , 
     n44641 , n44642 , n44643 , n44644 , n44645 , n44646 , n44647 , n44648 , n44649 , n44650 , 
     n44651 , n44652 , n44653 , n44654 , n44655 , n44656 , n44657 , n44658 , n44659 , n44660 , 
     n44661 , n44662 , n44663 , n44664 , n44665 , n44666 , n44667 , n44668 , n44669 , n44670 , 
     n44671 , n44672 , n44673 , n44674 , n44675 , n44676 , n44677 , n44678 , n44679 , n44680 , 
     n44681 , n44682 , n44683 , n44684 , n44685 , n44686 , n44687 , n44688 , n44689 , n44690 , 
     n44691 , n44692 , n44693 , n44694 , n44695 , n44696 , n44697 , n44698 , n44699 , n44700 , 
     n44701 , n44702 , n44703 , n44704 , n44705 , n44706 , n44707 , n44708 , n44709 , n44710 , 
     n44711 , n44712 , n44713 , n44714 , n44715 , n44716 , n44717 , n44718 , n44719 , n44720 , 
     n44721 , n44722 , n44723 , n44724 , n44725 , n44726 , n44727 , n44728 , n44729 , n44730 , 
     n44731 , n44732 , n44733 , n44734 , n44735 , n44736 , n44737 , n44738 , n44739 , n44740 , 
     n44741 , n44742 , n44743 , n44744 , n44745 , n44746 , n44747 , n44748 , n44749 , n44750 , 
     n44751 , n44752 , n44753 , n44754 , n44755 , n44756 , n44757 , n44758 , n44759 , n44760 , 
     n44761 , n44762 , n44763 , n44764 , n44765 , n44766 , n44767 , n44768 , n44769 , n44770 , 
     n44771 , n44772 , n44773 , n44774 , n44775 , n44776 , n44777 , n44778 , n44779 , n44780 , 
     n44781 , n44782 , n44783 , n44784 , n44785 , n44786 , n44787 , n44788 , n44789 , n44790 , 
     n44791 , n44792 , n44793 , n44794 , n44795 , n44796 , n44797 , n44798 , n44799 , n44800 , 
     n44801 , n44802 , n44803 , n44804 , n44805 , n44806 , n44807 , n44808 , n44809 , n44810 , 
     n44811 , n44812 , n44813 , n44814 , n44815 , n44816 , n44817 , n44818 , n44819 , n44820 , 
     n44821 , n44822 , n44823 , n44824 , n44825 , n44826 , n44827 , n44828 , n44829 , n44830 , 
     n44831 , n44832 , n44833 , n44834 , n44835 , n44836 , n44837 , n44838 , n44839 , n44840 , 
     n44841 , n44842 , n44843 , n44844 , n44845 , n44846 , n44847 , n44848 , n44849 , n44850 , 
     n44851 , n44852 , n44853 , n44854 , n44855 , n44856 , n44857 , n44858 , n44859 , n44860 , 
     n44861 , n44862 , n44863 , n44864 , n44865 , n44866 , n44867 , n44868 , n44869 , n44870 , 
     n44871 , n44872 , n44873 , n44874 , n44875 , n44876 , n44877 , n44878 , n44879 , n44880 , 
     n44881 , n44882 , n44883 , n44884 , n44885 , n44886 , n44887 , n44888 , n44889 , n44890 , 
     n44891 , n44892 , n44893 , n44894 , n44895 , n44896 , n44897 , n44898 , n44899 , n44900 , 
     n44901 , n44902 , n44903 , n44904 , n44905 , n44906 , n44907 , n44908 , n44909 , n44910 , 
     n44911 , n44912 , n44913 , n44914 , n44915 , n44916 , n44917 , n44918 , n44919 , n44920 , 
     n44921 , n44922 , n44923 , n44924 , n44925 , n44926 , n44927 , n44928 , n44929 , n44930 , 
     n44931 , n44932 , n44933 , n44934 , n44935 , n44936 , n44937 , n44938 , n44939 , n44940 , 
     n44941 , n44942 , n44943 , n44944 , n44945 , n44946 , n44947 , n44948 , n44949 , n44950 , 
     n44951 , n44952 , n44953 , n44954 , n44955 , n44956 , n44957 , n44958 , n44959 , n44960 , 
     n44961 , n44962 , n44963 , n44964 , n44965 , n44966 , n44967 , n44968 , n44969 , n44970 , 
     n44971 , n44972 , n44973 , n44974 , n44975 , n44976 , n44977 , n44978 , n44979 , n44980 , 
     n44981 , n44982 , n44983 , n44984 , n44985 , n44986 , n44987 , n44988 , n44989 , n44990 , 
     n44991 , n44992 , n44993 , n44994 , n44995 , n44996 , n44997 , n44998 , n44999 , n45000 , 
     n45001 , n45002 , n45003 , n45004 , n45005 , n45006 , n45007 , n45008 , n45009 , n45010 , 
     n45011 , n45012 , n45013 , n45014 , n45015 , n45016 , n45017 , n45018 , n45019 , n45020 , 
     n45021 , n45022 , n45023 , n45024 , n45025 , n45026 , n45027 , n45028 , n45029 , n45030 , 
     n45031 , n45032 , n45033 , n45034 , n45035 , n45036 , n45037 , n45038 , n45039 , n45040 , 
     n45041 , n45042 , n45043 , n45044 , n45045 , n45046 , n45047 , n45048 , n45049 , n45050 , 
     n45051 , n45052 , n45053 , n45054 , n45055 , n45056 , n45057 , n45058 , n45059 , n45060 , 
     n45061 , n45062 , n45063 , n45064 , n45065 , n45066 , n45067 , n45068 , n45069 , n45070 , 
     n45071 , n45072 , n45073 , n45074 , n45075 , n45076 , n45077 , n45078 , n45079 , n45080 , 
     n45081 , n45082 , n45083 , n45084 , n45085 , n45086 , n45087 , n45088 , n45089 , n45090 , 
     n45091 , n45092 , n45093 , n45094 , n45095 , n45096 , n45097 , n45098 , n45099 , n45100 , 
     n45101 , n45102 , n45103 , n45104 , n45105 , n45106 , n45107 , n45108 , n45109 , n45110 , 
     n45111 , n45112 , n45113 , n45114 , n45115 , n45116 , n45117 , n45118 , n45119 , n45120 , 
     n45121 , n45122 , n45123 , n45124 , n45125 , n45126 , n45127 , n45128 , n45129 , n45130 , 
     n45131 , n45132 , n45133 , n45134 , n45135 , n45136 , n45137 , n45138 , n45139 , n45140 , 
     n45141 , n45142 , n45143 , n45144 , n45145 , n45146 , n45147 , n45148 , n45149 , n45150 , 
     n45151 , n45152 , n45153 , n45154 , n45155 , n45156 , n45157 , n45158 , n45159 , n45160 , 
     n45161 , n45162 , n45163 , n45164 , n45165 , n45166 , n45167 , n45168 , n45169 , n45170 , 
     n45171 , n45172 , n45173 , n45174 , n45175 , n45176 , n45177 , n45178 , n45179 , n45180 , 
     n45181 , n45182 , n45183 , n45184 , n45185 , n45186 , n45187 , n45188 , n45189 , n45190 , 
     n45191 , n45192 , n45193 , n45194 , n45195 , n45196 , n45197 , n45198 , n45199 , n45200 , 
     n45201 , n45202 , n45203 , n45204 , n45205 , n45206 , n45207 , n45208 , n45209 , n45210 , 
     n45211 , n45212 , n45213 , n45214 , n45215 , n45216 , n45217 , n45218 , n45219 , n45220 , 
     n45221 , n45222 , n45223 , n45224 , n45225 , n45226 , n45227 , n45228 , n45229 , n45230 , 
     n45231 , n45232 , n45233 , n45234 , n45235 , n45236 , n45237 , n45238 , n45239 , n45240 , 
     n45241 , n45242 , n45243 , n45244 , n45245 , n45246 , n45247 , n45248 , n45249 , n45250 , 
     n45251 , n45252 , n45253 , n45254 , n45255 , n45256 , n45257 , n45258 , n45259 , n45260 , 
     n45261 , n45262 , n45263 , n45264 , n45265 , n45266 , n45267 , n45268 , n45269 , n45270 , 
     n45271 , n45272 , n45273 , n45274 , n45275 , n45276 , n45277 , n45278 , n45279 , n45280 , 
     n45281 , n45282 , n45283 , n45284 , n45285 , n45286 , n45287 , n45288 , n45289 , n45290 , 
     n45291 , n45292 , n45293 , n45294 , n45295 , n45296 , n45297 , n45298 , n45299 , n45300 , 
     n45301 , n45302 , n45303 , n45304 , n45305 , n45306 , n45307 , n45308 , n45309 , n45310 , 
     n45311 , n45312 , n45313 , n45314 , n45315 , n45316 , n45317 , n45318 , n45319 , n45320 , 
     n45321 , n45322 , n45323 , n45324 , n45325 , n45326 , n45327 , n45328 , n45329 , n45330 , 
     n45331 , n45332 , n45333 , n45334 , n45335 , n45336 , n45337 , n45338 , n45339 , n45340 , 
     n45341 , n45342 , n45343 , n45344 , n45345 , n45346 , n45347 , n45348 , n45349 , n45350 , 
     n45351 , n45352 , n45353 , n45354 , n45355 , n45356 , n45357 , n45358 , n45359 , n45360 , 
     n45361 , n45362 , n45363 , n45364 , n45365 , n45366 , n45367 , n45368 , n45369 , n45370 , 
     n45371 , n45372 , n45373 , n45374 , n45375 , n45376 , n45377 , n45378 , n45379 , n45380 , 
     n45381 , n45382 , n45383 , n45384 , n45385 , n45386 , n45387 , n45388 , n45389 , n45390 , 
     n45391 , n45392 , n45393 , n45394 , n45395 , n45396 , n45397 , n45398 , n45399 , n45400 , 
     n45401 , n45402 , n45403 , n45404 , n45405 , n45406 , n45407 , n45408 , n45409 , n45410 , 
     n45411 , n45412 , n45413 , n45414 , n45415 , n45416 , n45417 , n45418 , n45419 , n45420 , 
     n45421 , n45422 , n45423 , n45424 , n45425 , n45426 , n45427 , n45428 , n45429 , n45430 , 
     n45431 , n45432 , n45433 , n45434 , n45435 , n45436 , n45437 , n45438 , n45439 , n45440 , 
     n45441 , n45442 , n45443 , n45444 , n45445 , n45446 , n45447 , n45448 , n45449 , n45450 , 
     n45451 , n45452 , n45453 , n45454 , n45455 , n45456 , n45457 , n45458 , n45459 , n45460 , 
     n45461 , n45462 , n45463 , n45464 , n45465 , n45466 , n45467 , n45468 , n45469 , n45470 , 
     n45471 , n45472 , n45473 , n45474 , n45475 , n45476 , n45477 , n45478 , n45479 , n45480 , 
     n45481 , n45482 , n45483 , n45484 , n45485 , n45486 , n45487 , n45488 , n45489 , n45490 , 
     n45491 , n45492 , n45493 , n45494 , n45495 , n45496 , n45497 , n45498 , n45499 , n45500 , 
     n45501 , n45502 , n45503 , n45504 , n45505 , n45506 , n45507 , n45508 , n45509 , n45510 , 
     n45511 , n45512 , n45513 , n45514 , n45515 , n45516 , n45517 , n45518 , n45519 , n45520 , 
     n45521 , n45522 , n45523 , n45524 , n45525 , n45526 , n45527 , n45528 , n45529 , n45530 , 
     n45531 , n45532 , n45533 , n45534 , n45535 , n45536 , n45537 , n45538 , n45539 , n45540 , 
     n45541 , n45542 , n45543 , n45544 , n45545 , n45546 , n45547 , n45548 , n45549 , n45550 , 
     n45551 , n45552 , n45553 , n45554 , n45555 , n45556 , n45557 , n45558 , n45559 , n45560 , 
     n45561 , n45562 , n45563 , n45564 , n45565 , n45566 , n45567 , n45568 , n45569 , n45570 , 
     n45571 , n45572 , n45573 , n45574 , n45575 , n45576 , n45577 , n45578 , n45579 , n45580 , 
     n45581 , n45582 , n45583 , n45584 , n45585 , n45586 , n45587 , n45588 , n45589 , n45590 , 
     n45591 , n45592 , n45593 , n45594 , n45595 , n45596 , n45597 , n45598 , n45599 , n45600 , 
     n45601 , n45602 , n45603 , n45604 , n45605 , n45606 , n45607 , n45608 , n45609 , n45610 , 
     n45611 , n45612 , n45613 , n45614 , n45615 , n45616 , n45617 , n45618 , n45619 , n45620 , 
     n45621 , n45622 , n45623 , n45624 , n45625 , n45626 , n45627 , n45628 , n45629 , n45630 , 
     n45631 , n45632 , n45633 , n45634 , n45635 , n45636 , n45637 , n45638 , n45639 , n45640 , 
     n45641 , n45642 , n45643 , n45644 , n45645 , n45646 , n45647 , n45648 , n45649 , n45650 , 
     n45651 , n45652 , n45653 , n45654 , n45655 , n45656 , n45657 , n45658 , n45659 , n45660 , 
     n45661 , n45662 , n45663 , n45664 , n45665 , n45666 , n45667 , n45668 , n45669 , n45670 , 
     n45671 , n45672 , n45673 , n45674 , n45675 , n45676 , n45677 , n45678 , n45679 , n45680 , 
     n45681 , n45682 , n45683 , n45684 , n45685 , n45686 , n45687 , n45688 , n45689 , n45690 , 
     n45691 , n45692 , n45693 , n45694 , n45695 , n45696 , n45697 , n45698 , n45699 , n45700 , 
     n45701 , n45702 , n45703 , n45704 , n45705 , n45706 , n45707 , n45708 , n45709 , n45710 , 
     n45711 , n45712 , n45713 , n45714 , n45715 , n45716 , n45717 , n45718 , n45719 , n45720 , 
     n45721 , n45722 , n45723 , n45724 , n45725 , n45726 , n45727 , n45728 , n45729 , n45730 , 
     n45731 , n45732 , n45733 , n45734 , n45735 , n45736 , n45737 , n45738 , n45739 , n45740 , 
     n45741 , n45742 , n45743 , n45744 , n45745 , n45746 , n45747 , n45748 , n45749 , n45750 , 
     n45751 , n45752 , n45753 , n45754 , n45755 , n45756 , n45757 , n45758 , n45759 , n45760 , 
     n45761 , n45762 , n45763 , n45764 , n45765 , n45766 , n45767 , n45768 , n45769 , n45770 , 
     n45771 , n45772 , n45773 , n45774 , n45775 , n45776 , n45777 , n45778 , n45779 , n45780 , 
     n45781 , n45782 , n45783 , n45784 , n45785 , n45786 , n45787 , n45788 , n45789 , n45790 , 
     n45791 , n45792 , n45793 , n45794 , n45795 , n45796 , n45797 , n45798 , n45799 , n45800 , 
     n45801 , n45802 , n45803 , n45804 , n45805 , n45806 , n45807 , n45808 , n45809 , n45810 , 
     n45811 , n45812 , n45813 , n45814 , n45815 , n45816 , n45817 , n45818 , n45819 , n45820 , 
     n45821 , n45822 , n45823 , n45824 , n45825 , n45826 , n45827 , n45828 , n45829 , n45830 , 
     n45831 , n45832 , n45833 , n45834 , n45835 , n45836 , n45837 , n45838 , n45839 , n45840 , 
     n45841 , n45842 , n45843 , n45844 , n45845 , n45846 , n45847 , n45848 , n45849 , n45850 , 
     n45851 , n45852 , n45853 , n45854 , n45855 , n45856 , n45857 , n45858 , n45859 , n45860 , 
     n45861 , n45862 , n45863 , n45864 , n45865 , n45866 , n45867 , n45868 , n45869 , n45870 , 
     n45871 , n45872 , n45873 , n45874 , n45875 , n45876 , n45877 , n45878 , n45879 , n45880 , 
     n45881 , n45882 , n45883 , n45884 , n45885 , n45886 , n45887 , n45888 , n45889 , n45890 , 
     n45891 , n45892 , n45893 , n45894 , n45895 , n45896 , n45897 , n45898 , n45899 , n45900 , 
     n45901 , n45902 , n45903 , n45904 , n45905 , n45906 , n45907 , n45908 , n45909 , n45910 , 
     n45911 , n45912 , n45913 , n45914 , n45915 , n45916 , n45917 , n45918 , n45919 , n45920 , 
     n45921 , n45922 , n45923 , n45924 , n45925 , n45926 , n45927 , n45928 , n45929 , n45930 , 
     n45931 , n45932 , n45933 , n45934 , n45935 , n45936 , n45937 , n45938 , n45939 , n45940 , 
     n45941 , n45942 , n45943 , n45944 , n45945 , n45946 , n45947 , n45948 , n45949 , n45950 , 
     n45951 , n45952 , n45953 , n45954 , n45955 , n45956 , n45957 , n45958 , n45959 , n45960 , 
     n45961 , n45962 , n45963 , n45964 , n45965 , n45966 , n45967 , n45968 , n45969 , n45970 , 
     n45971 , n45972 , n45973 , n45974 , n45975 , n45976 , n45977 , n45978 , n45979 , n45980 , 
     n45981 , n45982 , n45983 , n45984 , n45985 , n45986 , n45987 , n45988 , n45989 , n45990 , 
     n45991 , n45992 , n45993 , n45994 , n45995 , n45996 , n45997 , n45998 , n45999 , n46000 , 
     n46001 , n46002 , n46003 , n46004 , n46005 , n46006 , n46007 , n46008 , n46009 , n46010 , 
     n46011 , n46012 , n46013 , n46014 , n46015 , n46016 , n46017 , n46018 , n46019 , n46020 , 
     n46021 , n46022 , n46023 , n46024 , n46025 , n46026 , n46027 , n46028 , n46029 , n46030 , 
     n46031 , n46032 , n46033 , n46034 , n46035 , n46036 , n46037 , n46038 , n46039 , n46040 , 
     n46041 , n46042 , n46043 , n46044 , n46045 , n46046 , n46047 , n46048 , n46049 , n46050 , 
     n46051 , n46052 , n46053 , n46054 , n46055 , n46056 , n46057 , n46058 , n46059 , n46060 , 
     n46061 , n46062 , n46063 , n46064 , n46065 , n46066 , n46067 , n46068 , n46069 , n46070 , 
     n46071 , n46072 , n46073 , n46074 , n46075 , n46076 , n46077 , n46078 , n46079 , n46080 , 
     n46081 , n46082 , n46083 , n46084 , n46085 , n46086 , n46087 , n46088 , n46089 , n46090 , 
     n46091 , n46092 , n46093 , n46094 , n46095 , n46096 , n46097 , n46098 , n46099 , n46100 , 
     n46101 , n46102 , n46103 , n46104 , n46105 , n46106 , n46107 , n46108 , n46109 , n46110 , 
     n46111 , n46112 , n46113 , n46114 , n46115 , n46116 , n46117 , n46118 , n46119 , n46120 , 
     n46121 , n46122 , n46123 , n46124 , n46125 , n46126 , n46127 , n46128 , n46129 , n46130 , 
     n46131 , n46132 , n46133 , n46134 , n46135 , n46136 , n46137 , n46138 , n46139 , n46140 , 
     n46141 , n46142 , n46143 , n46144 , n46145 , n46146 , n46147 , n46148 , n46149 , n46150 , 
     n46151 , n46152 , n46153 , n46154 , n46155 , n46156 , n46157 , n46158 , n46159 , n46160 , 
     n46161 , n46162 , n46163 , n46164 , n46165 , n46166 , n46167 , n46168 , n46169 , n46170 , 
     n46171 , n46172 , n46173 , n46174 , n46175 , n46176 , n46177 , n46178 , n46179 , n46180 , 
     n46181 , n46182 , n46183 , n46184 , n46185 , n46186 , n46187 , n46188 , n46189 , n46190 , 
     n46191 , n46192 , n46193 , n46194 , n46195 , n46196 , n46197 , n46198 , n46199 , n46200 , 
     n46201 , n46202 , n46203 , n46204 , n46205 , n46206 , n46207 , n46208 , n46209 , n46210 , 
     n46211 , n46212 , n46213 , n46214 , n46215 , n46216 , n46217 , n46218 , n46219 , n46220 , 
     n46221 , n46222 , n46223 , n46224 , n46225 , n46226 , n46227 , n46228 , n46229 , n46230 , 
     n46231 , n46232 , n46233 , n46234 , n46235 , n46236 , n46237 , n46238 , n46239 , n46240 , 
     n46241 , n46242 , n46243 , n46244 , n46245 , n46246 , n46247 , n46248 , n46249 , n46250 , 
     n46251 , n46252 , n46253 , n46254 , n46255 , n46256 , n46257 , n46258 , n46259 , n46260 , 
     n46261 , n46262 , n46263 , n46264 , n46265 , n46266 , n46267 , n46268 , n46269 , n46270 , 
     n46271 , n46272 , n46273 , n46274 , n46275 , n46276 , n46277 , n46278 , n46279 , n46280 , 
     n46281 , n46282 , n46283 , n46284 , n46285 , n46286 , n46287 , n46288 , n46289 , n46290 , 
     n46291 , n46292 , n46293 , n46294 , n46295 , n46296 , n46297 , n46298 , n46299 , n46300 , 
     n46301 , n46302 , n46303 , n46304 , n46305 , n46306 , n46307 , n46308 , n46309 , n46310 , 
     n46311 , n46312 , n46313 , n46314 , n46315 , n46316 , n46317 , n46318 , n46319 , n46320 , 
     n46321 , n46322 , n46323 , n46324 , n46325 , n46326 , n46327 , n46328 , n46329 , n46330 , 
     n46331 , n46332 , n46333 , n46334 , n46335 , n46336 , n46337 , n46338 , n46339 , n46340 , 
     n46341 , n46342 , n46343 , n46344 , n46345 , n46346 , n46347 , n46348 , n46349 , n46350 , 
     n46351 , n46352 , n46353 , n46354 , n46355 , n46356 , n46357 , n46358 , n46359 , n46360 , 
     n46361 , n46362 , n46363 , n46364 , n46365 , n46366 , n46367 , n46368 , n46369 , n46370 , 
     n46371 , n46372 , n46373 , n46374 , n46375 , n46376 , n46377 , n46378 , n46379 , n46380 , 
     n46381 , n46382 , n46383 , n46384 , n46385 , n46386 , n46387 , n46388 , n46389 , n46390 , 
     n46391 , n46392 , n46393 , n46394 , n46395 , n46396 , n46397 , n46398 , n46399 , n46400 , 
     n46401 , n46402 , n46403 , n46404 , n46405 , n46406 , n46407 , n46408 , n46409 , n46410 , 
     n46411 , n46412 , n46413 , n46414 , n46415 , n46416 , n46417 , n46418 , n46419 , n46420 , 
     n46421 , n46422 , n46423 , n46424 , n46425 , n46426 , n46427 , n46428 , n46429 , n46430 , 
     n46431 , n46432 , n46433 , n46434 , n46435 , n46436 , n46437 , n46438 , n46439 , n46440 , 
     n46441 , n46442 , n46443 , n46444 , n46445 , n46446 , n46447 , n46448 , n46449 , n46450 , 
     n46451 , n46452 , n46453 , n46454 , n46455 , n46456 , n46457 , n46458 , n46459 , n46460 , 
     n46461 , n46462 , n46463 , n46464 , n46465 , n46466 , n46467 , n46468 , n46469 , n46470 , 
     n46471 , n46472 , n46473 , n46474 , n46475 , n46476 , n46477 , n46478 , n46479 , n46480 , 
     n46481 , n46482 , n46483 , n46484 , n46485 , n46486 , n46487 , n46488 , n46489 , n46490 , 
     n46491 , n46492 , n46493 , n46494 , n46495 , n46496 , n46497 , n46498 , n46499 , n46500 , 
     n46501 , n46502 , n46503 , n46504 , n46505 , n46506 , n46507 , n46508 , n46509 , n46510 , 
     n46511 , n46512 , n46513 , n46514 , n46515 , n46516 , n46517 , n46518 , n46519 , n46520 , 
     n46521 , n46522 , n46523 , n46524 , n46525 , n46526 , n46527 , n46528 , n46529 , n46530 , 
     n46531 , n46532 , n46533 , n46534 , n46535 , n46536 , n46537 , n46538 , n46539 , n46540 , 
     n46541 , n46542 , n46543 , n46544 , n46545 , n46546 , n46547 , n46548 , n46549 , n46550 , 
     n46551 , n46552 , n46553 , n46554 , n46555 , n46556 , n46557 , n46558 , n46559 , n46560 , 
     n46561 , n46562 , n46563 , n46564 , n46565 , n46566 , n46567 , n46568 , n46569 , n46570 , 
     n46571 , n46572 , n46573 , n46574 , n46575 , n46576 , n46577 , n46578 , n46579 , n46580 , 
     n46581 , n46582 , n46583 , n46584 , n46585 , n46586 , n46587 , n46588 , n46589 , n46590 , 
     n46591 , n46592 , n46593 , n46594 , n46595 , n46596 , n46597 , n46598 , n46599 , n46600 , 
     n46601 , n46602 , n46603 , n46604 , n46605 , n46606 , n46607 , n46608 , n46609 , n46610 , 
     n46611 , n46612 , n46613 , n46614 , n46615 , n46616 , n46617 , n46618 , n46619 , n46620 , 
     n46621 , n46622 , n46623 , n46624 , n46625 , n46626 , n46627 , n46628 , n46629 , n46630 , 
     n46631 , n46632 , n46633 , n46634 , n46635 , n46636 , n46637 , n46638 , n46639 , n46640 , 
     n46641 , n46642 , n46643 , n46644 , n46645 , n46646 , n46647 , n46648 , n46649 , n46650 , 
     n46651 , n46652 , n46653 , n46654 , n46655 , n46656 , n46657 , n46658 , n46659 , n46660 , 
     n46661 , n46662 , n46663 , n46664 , n46665 , n46666 , n46667 , n46668 , n46669 , n46670 , 
     n46671 , n46672 , n46673 , n46674 , n46675 , n46676 , n46677 , n46678 , n46679 , n46680 , 
     n46681 , n46682 , n46683 , n46684 , n46685 , n46686 , n46687 , n46688 , n46689 , n46690 , 
     n46691 , n46692 , n46693 , n46694 , n46695 , n46696 , n46697 , n46698 , n46699 , n46700 , 
     n46701 , n46702 , n46703 , n46704 , n46705 , n46706 , n46707 , n46708 , n46709 , n46710 , 
     n46711 , n46712 , n46713 , n46714 , n46715 , n46716 , n46717 , n46718 , n46719 , n46720 , 
     n46721 , n46722 , n46723 , n46724 , n46725 , n46726 , n46727 , n46728 , n46729 , n46730 , 
     n46731 , n46732 , n46733 , n46734 , n46735 , n46736 , n46737 , n46738 , n46739 , n46740 , 
     n46741 , n46742 , n46743 , n46744 , n46745 , n46746 , n46747 , n46748 , n46749 , n46750 , 
     n46751 , n46752 , n46753 , n46754 , n46755 , n46756 , n46757 , n46758 , n46759 , n46760 , 
     n46761 , n46762 , n46763 , n46764 , n46765 , n46766 , n46767 , n46768 , n46769 , n46770 , 
     n46771 , n46772 , n46773 , n46774 , n46775 , n46776 , n46777 , n46778 , n46779 , n46780 , 
     n46781 , n46782 , n46783 , n46784 , n46785 , n46786 , n46787 , n46788 , n46789 , n46790 , 
     n46791 , n46792 , n46793 , n46794 , n46795 , n46796 , n46797 , n46798 , n46799 , n46800 , 
     n46801 , n46802 , n46803 , n46804 , n46805 , n46806 , n46807 , n46808 , n46809 , n46810 , 
     n46811 , n46812 , n46813 , n46814 , n46815 , n46816 , n46817 , n46818 , n46819 , n46820 , 
     n46821 , n46822 , n46823 , n46824 , n46825 , n46826 , n46827 , n46828 , n46829 , n46830 , 
     n46831 , n46832 , n46833 , n46834 , n46835 , n46836 , n46837 , n46838 , n46839 , n46840 , 
     n46841 , n46842 , n46843 , n46844 , n46845 , n46846 , n46847 , n46848 , n46849 , n46850 , 
     n46851 , n46852 , n46853 , n46854 , n46855 , n46856 , n46857 , n46858 , n46859 , n46860 , 
     n46861 , n46862 , n46863 , n46864 , n46865 , n46866 , n46867 , n46868 , n46869 , n46870 , 
     n46871 , n46872 , n46873 , n46874 , n46875 , n46876 , n46877 , n46878 , n46879 , n46880 , 
     n46881 , n46882 , n46883 , n46884 , n46885 , n46886 , n46887 , n46888 , n46889 , n46890 , 
     n46891 , n46892 , n46893 , n46894 , n46895 , n46896 , n46897 , n46898 , n46899 , n46900 , 
     n46901 , n46902 , n46903 , n46904 , n46905 , n46906 , n46907 , n46908 , n46909 , n46910 , 
     n46911 , n46912 , n46913 , n46914 , n46915 , n46916 , n46917 , n46918 , n46919 , n46920 , 
     n46921 , n46922 , n46923 , n46924 , n46925 , n46926 , n46927 , n46928 , n46929 , n46930 , 
     n46931 , n46932 , n46933 , n46934 , n46935 , n46936 , n46937 , n46938 , n46939 , n46940 , 
     n46941 , n46942 , n46943 , n46944 , n46945 , n46946 , n46947 , n46948 , n46949 , n46950 , 
     n46951 , n46952 , n46953 , n46954 , n46955 , n46956 , n46957 , n46958 , n46959 , n46960 , 
     n46961 , n46962 , n46963 , n46964 , n46965 , n46966 , n46967 , n46968 , n46969 , n46970 , 
     n46971 , n46972 , n46973 , n46974 , n46975 , n46976 , n46977 , n46978 , n46979 , n46980 , 
     n46981 , n46982 , n46983 , n46984 , n46985 , n46986 , n46987 , n46988 , n46989 , n46990 , 
     n46991 , n46992 , n46993 , n46994 , n46995 , n46996 , n46997 , n46998 , n46999 , n47000 , 
     n47001 , n47002 , n47003 , n47004 , n47005 , n47006 , n47007 , n47008 , n47009 , n47010 , 
     n47011 , n47012 , n47013 , n47014 , n47015 , n47016 , n47017 , n47018 , n47019 , n47020 , 
     n47021 , n47022 , n47023 , n47024 , n47025 , n47026 , n47027 , n47028 , n47029 , n47030 , 
     n47031 , n47032 , n47033 , n47034 , n47035 , n47036 , n47037 , n47038 , n47039 , n47040 , 
     n47041 , n47042 , n47043 , n47044 , n47045 , n47046 , n47047 , n47048 , n47049 , n47050 , 
     n47051 , n47052 , n47053 , n47054 , n47055 , n47056 , n47057 , n47058 , n47059 , n47060 , 
     n47061 , n47062 , n47063 , n47064 , n47065 , n47066 , n47067 , n47068 , n47069 , n47070 , 
     n47071 , n47072 , n47073 , n47074 , n47075 , n47076 , n47077 , n47078 , n47079 , n47080 , 
     n47081 , n47082 , n47083 , n47084 , n47085 , n47086 , n47087 , n47088 , n47089 , n47090 , 
     n47091 , n47092 , n47093 , n47094 , n47095 , n47096 , n47097 , n47098 , n47099 , n47100 , 
     n47101 , n47102 , n47103 , n47104 , n47105 , n47106 , n47107 , n47108 , n47109 , n47110 , 
     n47111 , n47112 , n47113 , n47114 , n47115 , n47116 , n47117 , n47118 , n47119 , n47120 , 
     n47121 , n47122 , n47123 , n47124 , n47125 , n47126 , n47127 , n47128 , n47129 , n47130 , 
     n47131 , n47132 , n47133 , n47134 , n47135 , n47136 , n47137 , n47138 , n47139 , n47140 , 
     n47141 , n47142 , n47143 , n47144 , n47145 , n47146 , n47147 , n47148 , n47149 , n47150 , 
     n47151 , n47152 , n47153 , n47154 , n47155 , n47156 , n47157 , n47158 , n47159 , n47160 , 
     n47161 , n47162 , n47163 , n47164 , n47165 , n47166 , n47167 , n47168 , n47169 , n47170 , 
     n47171 , n47172 , n47173 , n47174 , n47175 , n47176 , n47177 , n47178 , n47179 , n47180 , 
     n47181 , n47182 , n47183 , n47184 , n47185 , n47186 , n47187 , n47188 , n47189 , n47190 , 
     n47191 , n47192 , n47193 , n47194 , n47195 , n47196 , n47197 , n47198 , n47199 , n47200 , 
     n47201 , n47202 , n47203 , n47204 , n47205 , n47206 , n47207 , n47208 , n47209 , n47210 , 
     n47211 , n47212 , n47213 , n47214 , n47215 , n47216 , n47217 , n47218 , n47219 , n47220 , 
     n47221 , n47222 , n47223 , n47224 , n47225 , n47226 , n47227 , n47228 , n47229 , n47230 , 
     n47231 , n47232 , n47233 , n47234 , n47235 , n47236 , n47237 , n47238 , n47239 , n47240 , 
     n47241 , n47242 , n47243 , n47244 , n47245 , n47246 , n47247 , n47248 , n47249 , n47250 , 
     n47251 , n47252 , n47253 , n47254 , n47255 , n47256 , n47257 , n47258 , n47259 , n47260 , 
     n47261 , n47262 , n47263 , n47264 , n47265 , n47266 , n47267 , n47268 , n47269 , n47270 , 
     n47271 , n47272 , n47273 , n47274 , n47275 , n47276 , n47277 , n47278 , n47279 , n47280 , 
     n47281 , n47282 , n47283 , n47284 , n47285 , n47286 , n47287 , n47288 , n47289 , n47290 , 
     n47291 , n47292 , n47293 , n47294 , n47295 , n47296 , n47297 , n47298 , n47299 , n47300 , 
     n47301 , n47302 , n47303 , n47304 , n47305 , n47306 , n47307 , n47308 , n47309 , n47310 , 
     n47311 , n47312 , n47313 , n47314 , n47315 , n47316 , n47317 , n47318 , n47319 , n47320 , 
     n47321 , n47322 , n47323 , n47324 , n47325 , n47326 , n47327 , n47328 , n47329 , n47330 , 
     n47331 , n47332 , n47333 , n47334 , n47335 , n47336 , n47337 , n47338 , n47339 , n47340 , 
     n47341 , n47342 , n47343 , n47344 , n47345 , n47346 , n47347 , n47348 , n47349 , n47350 , 
     n47351 , n47352 , n47353 , n47354 , n47355 , n47356 , n47357 , n47358 , n47359 , n47360 , 
     n47361 , n47362 , n47363 , n47364 , n47365 , n47366 , n47367 , n47368 , n47369 , n47370 , 
     n47371 , n47372 , n47373 , n47374 , n47375 , n47376 , n47377 , n47378 , n47379 , n47380 , 
     n47381 , n47382 , n47383 , n47384 , n47385 , n47386 , n47387 , n47388 , n47389 , n47390 , 
     n47391 , n47392 , n47393 , n47394 , n47395 , n47396 , n47397 , n47398 , n47399 , n47400 , 
     n47401 , n47402 , n47403 , n47404 , n47405 , n47406 , n47407 , n47408 , n47409 , n47410 , 
     n47411 , n47412 , n47413 , n47414 , n47415 , n47416 , n47417 , n47418 , n47419 , n47420 , 
     n47421 , n47422 , n47423 , n47424 , n47425 , n47426 , n47427 , n47428 , n47429 , n47430 , 
     n47431 , n47432 , n47433 , n47434 , n47435 , n47436 , n47437 , n47438 , n47439 , n47440 , 
     n47441 , n47442 , n47443 , n47444 , n47445 , n47446 , n47447 , n47448 , n47449 , n47450 , 
     n47451 , n47452 , n47453 , n47454 , n47455 , n47456 , n47457 , n47458 , n47459 , n47460 , 
     n47461 , n47462 , n47463 , n47464 , n47465 , n47466 , n47467 , n47468 , n47469 , n47470 , 
     n47471 , n47472 , n47473 , n47474 , n47475 , n47476 , n47477 , n47478 , n47479 , n47480 , 
     n47481 , n47482 , n47483 , n47484 , n47485 , n47486 , n47487 , n47488 , n47489 , n47490 , 
     n47491 , n47492 , n47493 , n47494 , n47495 , n47496 , n47497 , n47498 , n47499 , n47500 , 
     n47501 , n47502 , n47503 , n47504 , n47505 , n47506 , n47507 , n47508 , n47509 , n47510 , 
     n47511 , n47512 , n47513 , n47514 , n47515 , n47516 , n47517 , n47518 , n47519 , n47520 , 
     n47521 , n47522 , n47523 , n47524 , n47525 , n47526 , n47527 , n47528 , n47529 , n47530 , 
     n47531 , n47532 , n47533 , n47534 , n47535 , n47536 , n47537 , n47538 , n47539 , n47540 , 
     n47541 , n47542 , n47543 , n47544 , n47545 , n47546 , n47547 , n47548 , n47549 , n47550 , 
     n47551 , n47552 , n47553 , n47554 , n47555 , n47556 , n47557 , n47558 , n47559 , n47560 , 
     n47561 , n47562 , n47563 , n47564 , n47565 , n47566 , n47567 , n47568 , n47569 , n47570 , 
     n47571 , n47572 , n47573 , n47574 , n47575 , n47576 , n47577 , n47578 , n47579 , n47580 , 
     n47581 , n47582 , n47583 , n47584 , n47585 , n47586 , n47587 , n47588 , n47589 , n47590 , 
     n47591 , n47592 , n47593 , n47594 , n47595 , n47596 , n47597 , n47598 , n47599 , n47600 , 
     n47601 , n47602 , n47603 , n47604 , n47605 , n47606 , n47607 , n47608 , n47609 , n47610 , 
     n47611 , n47612 , n47613 , n47614 , n47615 , n47616 , n47617 , n47618 , n47619 , n47620 , 
     n47621 , n47622 , n47623 , n47624 , n47625 , n47626 , n47627 , n47628 , n47629 , n47630 , 
     n47631 , n47632 , n47633 , n47634 , n47635 , n47636 , n47637 , n47638 , n47639 , n47640 , 
     n47641 , n47642 , n47643 , n47644 , n47645 , n47646 , n47647 , n47648 , n47649 , n47650 , 
     n47651 , n47652 , n47653 , n47654 , n47655 , n47656 , n47657 , n47658 , n47659 , n47660 , 
     n47661 , n47662 , n47663 , n47664 , n47665 , n47666 , n47667 , n47668 , n47669 , n47670 , 
     n47671 , n47672 , n47673 , n47674 , n47675 , n47676 , n47677 , n47678 , n47679 , n47680 , 
     n47681 , n47682 , n47683 , n47684 , n47685 , n47686 , n47687 , n47688 , n47689 , n47690 , 
     n47691 , n47692 , n47693 , n47694 , n47695 , n47696 , n47697 , n47698 , n47699 , n47700 , 
     n47701 , n47702 , n47703 , n47704 , n47705 , n47706 , n47707 , n47708 , n47709 , n47710 , 
     n47711 , n47712 , n47713 , n47714 , n47715 , n47716 , n47717 , n47718 , n47719 , n47720 , 
     n47721 , n47722 , n47723 , n47724 , n47725 , n47726 , n47727 , n47728 , n47729 , n47730 , 
     n47731 , n47732 , n47733 , n47734 , n47735 , n47736 , n47737 , n47738 , n47739 , n47740 , 
     n47741 , n47742 , n47743 , n47744 , n47745 , n47746 , n47747 , n47748 , n47749 , n47750 , 
     n47751 , n47752 , n47753 , n47754 , n47755 , n47756 , n47757 , n47758 , n47759 , n47760 , 
     n47761 , n47762 , n47763 , n47764 , n47765 , n47766 , n47767 , n47768 , n47769 , n47770 , 
     n47771 , n47772 , n47773 , n47774 , n47775 , n47776 , n47777 , n47778 , n47779 , n47780 , 
     n47781 , n47782 , n47783 , n47784 , n47785 , n47786 , n47787 , n47788 , n47789 , n47790 , 
     n47791 , n47792 , n47793 , n47794 , n47795 , n47796 , n47797 , n47798 , n47799 , n47800 , 
     n47801 , n47802 , n47803 , n47804 , n47805 , n47806 , n47807 , n47808 , n47809 , n47810 , 
     n47811 , n47812 , n47813 , n47814 , n47815 , n47816 , n47817 , n47818 , n47819 , n47820 , 
     n47821 , n47822 , n47823 , n47824 , n47825 , n47826 , n47827 , n47828 , n47829 , n47830 , 
     n47831 , n47832 , n47833 , n47834 , n47835 , n47836 , n47837 , n47838 , n47839 , n47840 , 
     n47841 , n47842 , n47843 , n47844 , n47845 , n47846 , n47847 , n47848 , n47849 , n47850 , 
     n47851 , n47852 , n47853 , n47854 , n47855 , n47856 , n47857 , n47858 , n47859 , n47860 , 
     n47861 , n47862 , n47863 , n47864 , n47865 , n47866 , n47867 , n47868 , n47869 , n47870 , 
     n47871 , n47872 , n47873 , n47874 , n47875 , n47876 , n47877 , n47878 , n47879 , n47880 , 
     n47881 , n47882 , n47883 , n47884 , n47885 , n47886 , n47887 , n47888 , n47889 , n47890 , 
     n47891 , n47892 , n47893 , n47894 , n47895 , n47896 , n47897 , n47898 , n47899 , n47900 , 
     n47901 , n47902 , n47903 , n47904 , n47905 , n47906 , n47907 , n47908 , n47909 , n47910 , 
     n47911 , n47912 , n47913 , n47914 , n47915 , n47916 , n47917 , n47918 , n47919 , n47920 , 
     n47921 , n47922 , n47923 , n47924 , n47925 , n47926 , n47927 , n47928 , n47929 , n47930 , 
     n47931 , n47932 , n47933 , n47934 , n47935 , n47936 , n47937 , n47938 , n47939 , n47940 , 
     n47941 , n47942 , n47943 , n47944 , n47945 , n47946 , n47947 , n47948 , n47949 , n47950 , 
     n47951 , n47952 , n47953 , n47954 , n47955 , n47956 , n47957 , n47958 , n47959 , n47960 , 
     n47961 , n47962 , n47963 , n47964 , n47965 , n47966 , n47967 , n47968 , n47969 , n47970 , 
     n47971 , n47972 , n47973 , n47974 , n47975 , n47976 , n47977 , n47978 , n47979 , n47980 , 
     n47981 , n47982 , n47983 , n47984 , n47985 , n47986 , n47987 , n47988 , n47989 , n47990 , 
     n47991 , n47992 , n47993 , n47994 , n47995 , n47996 , n47997 , n47998 , n47999 , n48000 , 
     n48001 , n48002 , n48003 , n48004 , n48005 , n48006 , n48007 , n48008 , n48009 , n48010 , 
     n48011 , n48012 , n48013 , n48014 , n48015 , n48016 , n48017 , n48018 , n48019 , n48020 , 
     n48021 , n48022 , n48023 , n48024 , n48025 , n48026 , n48027 , n48028 , n48029 , n48030 , 
     n48031 , n48032 , n48033 , n48034 , n48035 , n48036 , n48037 , n48038 , n48039 , n48040 , 
     n48041 , n48042 , n48043 , n48044 , n48045 , n48046 , n48047 , n48048 , n48049 , n48050 , 
     n48051 , n48052 , n48053 , n48054 , n48055 , n48056 , n48057 , n48058 , n48059 , n48060 , 
     n48061 , n48062 , n48063 , n48064 , n48065 , n48066 , n48067 , n48068 , n48069 , n48070 , 
     n48071 , n48072 , n48073 , n48074 , n48075 , n48076 , n48077 , n48078 , n48079 , n48080 , 
     n48081 , n48082 , n48083 , n48084 , n48085 , n48086 , n48087 , n48088 , n48089 , n48090 , 
     n48091 , n48092 , n48093 , n48094 , n48095 , n48096 , n48097 , n48098 , n48099 , n48100 , 
     n48101 , n48102 , n48103 , n48104 , n48105 , n48106 , n48107 , n48108 , n48109 , n48110 , 
     n48111 , n48112 , n48113 , n48114 , n48115 , n48116 , n48117 , n48118 , n48119 , n48120 , 
     n48121 , n48122 , n48123 , n48124 , n48125 , n48126 , n48127 , n48128 , n48129 , n48130 , 
     n48131 , n48132 , n48133 , n48134 , n48135 , n48136 , n48137 , n48138 , n48139 , n48140 , 
     n48141 , n48142 , n48143 , n48144 , n48145 , n48146 , n48147 , n48148 , n48149 , n48150 , 
     n48151 , n48152 , n48153 , n48154 , n48155 , n48156 , n48157 , n48158 , n48159 , n48160 , 
     n48161 , n48162 , n48163 , n48164 , n48165 , n48166 , n48167 , n48168 , n48169 , n48170 , 
     n48171 , n48172 , n48173 , n48174 , n48175 , n48176 , n48177 , n48178 , n48179 , n48180 , 
     n48181 , n48182 , n48183 , n48184 , n48185 , n48186 , n48187 , n48188 , n48189 , n48190 , 
     n48191 , n48192 , n48193 , n48194 , n48195 , n48196 , n48197 , n48198 , n48199 , n48200 , 
     n48201 , n48202 , n48203 , n48204 , n48205 , n48206 , n48207 , n48208 , n48209 , n48210 , 
     n48211 , n48212 , n48213 , n48214 , n48215 , n48216 , n48217 , n48218 , n48219 , n48220 , 
     n48221 , n48222 , n48223 , n48224 , n48225 , n48226 , n48227 , n48228 , n48229 , n48230 , 
     n48231 , n48232 , n48233 , n48234 , n48235 , n48236 , n48237 , n48238 , n48239 , n48240 , 
     n48241 , n48242 , n48243 , n48244 , n48245 , n48246 , n48247 , n48248 , n48249 , n48250 , 
     n48251 , n48252 , n48253 , n48254 , n48255 , n48256 , n48257 , n48258 , n48259 , n48260 , 
     n48261 , n48262 , n48263 , n48264 , n48265 , n48266 , n48267 , n48268 , n48269 , n48270 , 
     n48271 , n48272 , n48273 , n48274 , n48275 , n48276 , n48277 , n48278 , n48279 , n48280 , 
     n48281 , n48282 , n48283 , n48284 , n48285 , n48286 , n48287 , n48288 , n48289 , n48290 , 
     n48291 , n48292 , n48293 , n48294 , n48295 , n48296 , n48297 , n48298 , n48299 , n48300 , 
     n48301 , n48302 , n48303 , n48304 , n48305 , n48306 , n48307 , n48308 , n48309 , n48310 , 
     n48311 , n48312 , n48313 , n48314 , n48315 , n48316 , n48317 , n48318 , n48319 , n48320 , 
     n48321 , n48322 , n48323 , n48324 , n48325 , n48326 , n48327 , n48328 , n48329 , n48330 , 
     n48331 , n48332 , n48333 , n48334 , n48335 , n48336 , n48337 , n48338 , n48339 , n48340 , 
     n48341 , n48342 , n48343 , n48344 , n48345 , n48346 , n48347 , n48348 , n48349 , n48350 , 
     n48351 , n48352 , n48353 , n48354 , n48355 , n48356 , n48357 , n48358 , n48359 , n48360 , 
     n48361 , n48362 , n48363 , n48364 , n48365 , n48366 , n48367 , n48368 , n48369 , n48370 , 
     n48371 , n48372 , n48373 , n48374 , n48375 , n48376 , n48377 , n48378 , n48379 , n48380 , 
     n48381 , n48382 , n48383 , n48384 , n48385 , n48386 , n48387 , n48388 , n48389 , n48390 , 
     n48391 , n48392 , n48393 , n48394 , n48395 , n48396 , n48397 , n48398 , n48399 , n48400 , 
     n48401 , n48402 , n48403 , n48404 , n48405 , n48406 , n48407 , n48408 , n48409 , n48410 , 
     n48411 , n48412 , n48413 , n48414 , n48415 , n48416 , n48417 , n48418 , n48419 , n48420 , 
     n48421 , n48422 , n48423 , n48424 , n48425 , n48426 , n48427 , n48428 , n48429 , n48430 , 
     n48431 , n48432 , n48433 , n48434 , n48435 , n48436 , n48437 , n48438 , n48439 , n48440 , 
     n48441 , n48442 , n48443 , n48444 , n48445 , n48446 , n48447 , n48448 , n48449 , n48450 , 
     n48451 , n48452 , n48453 , n48454 , n48455 , n48456 , n48457 , n48458 , n48459 , n48460 , 
     n48461 , n48462 , n48463 , n48464 , n48465 , n48466 , n48467 , n48468 , n48469 , n48470 , 
     n48471 , n48472 , n48473 , n48474 , n48475 , n48476 , n48477 , n48478 , n48479 , n48480 , 
     n48481 , n48482 , n48483 , n48484 , n48485 , n48486 , n48487 , n48488 , n48489 , n48490 , 
     n48491 , n48492 , n48493 , n48494 , n48495 , n48496 , n48497 , n48498 , n48499 , n48500 , 
     n48501 , n48502 , n48503 , n48504 , n48505 , n48506 , n48507 , n48508 , n48509 , n48510 , 
     n48511 , n48512 , n48513 , n48514 , n48515 , n48516 , n48517 , n48518 , n48519 , n48520 , 
     n48521 , n48522 , n48523 , n48524 , n48525 , n48526 , n48527 , n48528 , n48529 , n48530 , 
     n48531 , n48532 , n48533 , n48534 , n48535 , n48536 , n48537 , n48538 , n48539 , n48540 , 
     n48541 , n48542 , n48543 , n48544 , n48545 , n48546 , n48547 , n48548 , n48549 , n48550 , 
     n48551 , n48552 , n48553 , n48554 , n48555 , n48556 , n48557 , n48558 , n48559 , n48560 , 
     n48561 , n48562 , n48563 , n48564 , n48565 , n48566 , n48567 , n48568 , n48569 , n48570 , 
     n48571 , n48572 , n48573 , n48574 , n48575 , n48576 , n48577 , n48578 , n48579 , n48580 , 
     n48581 , n48582 , n48583 , n48584 , n48585 , n48586 , n48587 , n48588 , n48589 , n48590 , 
     n48591 , n48592 , n48593 , n48594 , n48595 , n48596 , n48597 , n48598 , n48599 , n48600 , 
     n48601 , n48602 , n48603 , n48604 , n48605 , n48606 , n48607 , n48608 , n48609 , n48610 , 
     n48611 , n48612 , n48613 , n48614 , n48615 , n48616 , n48617 , n48618 , n48619 , n48620 , 
     n48621 , n48622 , n48623 , n48624 , n48625 , n48626 , n48627 , n48628 , n48629 , n48630 , 
     n48631 , n48632 , n48633 , n48634 , n48635 , n48636 , n48637 , n48638 , n48639 , n48640 , 
     n48641 , n48642 , n48643 , n48644 , n48645 , n48646 , n48647 , n48648 , n48649 , n48650 , 
     n48651 , n48652 , n48653 , n48654 , n48655 , n48656 , n48657 , n48658 , n48659 , n48660 , 
     n48661 , n48662 , n48663 , n48664 , n48665 , n48666 , n48667 , n48668 , n48669 , n48670 , 
     n48671 , n48672 , n48673 , n48674 , n48675 , n48676 , n48677 , n48678 , n48679 , n48680 , 
     n48681 , n48682 , n48683 , n48684 , n48685 , n48686 , n48687 , n48688 , n48689 , n48690 , 
     n48691 , n48692 , n48693 , n48694 , n48695 , n48696 , n48697 , n48698 , n48699 , n48700 , 
     n48701 , n48702 , n48703 , n48704 , n48705 , n48706 , n48707 , n48708 , n48709 , n48710 , 
     n48711 , n48712 , n48713 , n48714 , n48715 , n48716 , n48717 , n48718 , n48719 , n48720 , 
     n48721 , n48722 , n48723 , n48724 , n48725 , n48726 , n48727 , n48728 , n48729 , n48730 , 
     n48731 , n48732 , n48733 , n48734 , n48735 , n48736 , n48737 , n48738 , n48739 , n48740 , 
     n48741 , n48742 , n48743 , n48744 , n48745 , n48746 , n48747 , n48748 , n48749 , n48750 , 
     n48751 , n48752 , n48753 , n48754 , n48755 , n48756 , n48757 , n48758 , n48759 , n48760 , 
     n48761 , n48762 , n48763 , n48764 , n48765 , n48766 , n48767 , n48768 , n48769 , n48770 , 
     n48771 , n48772 , n48773 , n48774 , n48775 , n48776 , n48777 , n48778 , n48779 , n48780 , 
     n48781 , n48782 , n48783 , n48784 , n48785 , n48786 , n48787 , n48788 , n48789 , n48790 , 
     n48791 , n48792 , n48793 , n48794 , n48795 , n48796 , n48797 , n48798 , n48799 , n48800 , 
     n48801 , n48802 , n48803 , n48804 , n48805 , n48806 , n48807 , n48808 , n48809 , n48810 , 
     n48811 , n48812 , n48813 , n48814 , n48815 , n48816 , n48817 , n48818 , n48819 , n48820 , 
     n48821 , n48822 , n48823 , n48824 , n48825 , n48826 , n48827 , n48828 , n48829 , n48830 , 
     n48831 , n48832 , n48833 , n48834 , n48835 , n48836 , n48837 , n48838 , n48839 , n48840 , 
     n48841 , n48842 , n48843 , n48844 , n48845 , n48846 , n48847 , n48848 , n48849 , n48850 , 
     n48851 , n48852 , n48853 , n48854 , n48855 , n48856 , n48857 , n48858 , n48859 , n48860 , 
     n48861 , n48862 , n48863 , n48864 , n48865 , n48866 , n48867 , n48868 , n48869 , n48870 , 
     n48871 , n48872 , n48873 , n48874 , n48875 , n48876 , n48877 , n48878 , n48879 , n48880 , 
     n48881 , n48882 , n48883 , n48884 , n48885 , n48886 , n48887 , n48888 , n48889 , n48890 , 
     n48891 , n48892 , n48893 , n48894 , n48895 , n48896 , n48897 , n48898 , n48899 , n48900 , 
     n48901 , n48902 , n48903 , n48904 , n48905 , n48906 , n48907 , n48908 , n48909 , n48910 , 
     n48911 , n48912 , n48913 , n48914 , n48915 , n48916 , n48917 , n48918 , n48919 , n48920 , 
     n48921 , n48922 , n48923 , n48924 , n48925 , n48926 , n48927 , n48928 , n48929 , n48930 , 
     n48931 , n48932 , n48933 , n48934 , n48935 , n48936 , n48937 , n48938 , n48939 , n48940 , 
     n48941 , n48942 , n48943 , n48944 , n48945 , n48946 , n48947 , n48948 , n48949 , n48950 , 
     n48951 , n48952 , n48953 , n48954 , n48955 , n48956 , n48957 , n48958 , n48959 , n48960 , 
     n48961 , n48962 , n48963 , n48964 , n48965 , n48966 , n48967 , n48968 , n48969 , n48970 , 
     n48971 , n48972 , n48973 , n48974 , n48975 , n48976 , n48977 , n48978 , n48979 , n48980 , 
     n48981 , n48982 , n48983 , n48984 , n48985 , n48986 , n48987 , n48988 , n48989 , n48990 , 
     n48991 , n48992 , n48993 , n48994 , n48995 , n48996 , n48997 , n48998 , n48999 , n49000 , 
     n49001 , n49002 , n49003 , n49004 , n49005 , n49006 , n49007 , n49008 , n49009 , n49010 , 
     n49011 , n49012 , n49013 , n49014 , n49015 , n49016 , n49017 , n49018 , n49019 , n49020 , 
     n49021 , n49022 , n49023 , n49024 , n49025 , n49026 , n49027 , n49028 , n49029 , n49030 , 
     n49031 , n49032 , n49033 , n49034 , n49035 , n49036 , n49037 , n49038 , n49039 , n49040 , 
     n49041 , n49042 , n49043 , n49044 , n49045 , n49046 , n49047 , n49048 , n49049 , n49050 , 
     n49051 , n49052 , n49053 , n49054 , n49055 , n49056 , n49057 , n49058 , n49059 , n49060 , 
     n49061 , n49062 , n49063 , n49064 , n49065 , n49066 , n49067 , n49068 , n49069 , n49070 , 
     n49071 , n49072 , n49073 , n49074 , n49075 , n49076 , n49077 , n49078 , n49079 , n49080 , 
     n49081 , n49082 , n49083 , n49084 , n49085 , n49086 , n49087 , n49088 , n49089 , n49090 , 
     n49091 , n49092 , n49093 , n49094 , n49095 , n49096 , n49097 , n49098 , n49099 , n49100 , 
     n49101 , n49102 , n49103 , n49104 , n49105 , n49106 , n49107 , n49108 , n49109 , n49110 , 
     n49111 , n49112 , n49113 , n49114 , n49115 , n49116 , n49117 , n49118 , n49119 , n49120 , 
     n49121 , n49122 , n49123 , n49124 , n49125 , n49126 , n49127 , n49128 , n49129 , n49130 , 
     n49131 , n49132 , n49133 , n49134 , n49135 , n49136 , n49137 , n49138 , n49139 , n49140 , 
     n49141 , n49142 , n49143 , n49144 , n49145 , n49146 , n49147 , n49148 , n49149 , n49150 , 
     n49151 , n49152 , n49153 , n49154 , n49155 , n49156 , n49157 , n49158 , n49159 , n49160 , 
     n49161 , n49162 , n49163 , n49164 , n49165 , n49166 , n49167 , n49168 , n49169 , n49170 , 
     n49171 , n49172 , n49173 , n49174 , n49175 , n49176 , n49177 , n49178 , n49179 , n49180 , 
     n49181 , n49182 , n49183 , n49184 , n49185 , n49186 , n49187 , n49188 , n49189 , n49190 , 
     n49191 , n49192 , n49193 , n49194 , n49195 , n49196 , n49197 , n49198 , n49199 , n49200 , 
     n49201 , n49202 , n49203 , n49204 , n49205 , n49206 , n49207 , n49208 , n49209 , n49210 , 
     n49211 , n49212 , n49213 , n49214 , n49215 , n49216 , n49217 , n49218 , n49219 , n49220 , 
     n49221 , n49222 , n49223 , n49224 , n49225 , n49226 , n49227 , n49228 , n49229 , n49230 , 
     n49231 , n49232 , n49233 , n49234 , n49235 , n49236 , n49237 , n49238 , n49239 , n49240 , 
     n49241 , n49242 , n49243 , n49244 , n49245 , n49246 , n49247 , n49248 , n49249 , n49250 , 
     n49251 , n49252 , n49253 , n49254 , n49255 , n49256 , n49257 , n49258 , n49259 , n49260 , 
     n49261 , n49262 , n49263 , n49264 , n49265 , n49266 , n49267 , n49268 , n49269 , n49270 , 
     n49271 , n49272 , n49273 , n49274 , n49275 , n49276 , n49277 , n49278 , n49279 , n49280 , 
     n49281 , n49282 , n49283 , n49284 , n49285 , n49286 , n49287 , n49288 , n49289 , n49290 , 
     n49291 , n49292 , n49293 , n49294 , n49295 , n49296 , n49297 , n49298 , n49299 , n49300 , 
     n49301 , n49302 , n49303 , n49304 , n49305 , n49306 , n49307 , n49308 , n49309 , n49310 , 
     n49311 , n49312 , n49313 , n49314 , n49315 , n49316 , n49317 , n49318 , n49319 , n49320 , 
     n49321 , n49322 , n49323 , n49324 , n49325 , n49326 , n49327 , n49328 , n49329 , n49330 , 
     n49331 , n49332 , n49333 , n49334 , n49335 , n49336 , n49337 , n49338 , n49339 , n49340 , 
     n49341 , n49342 , n49343 , n49344 , n49345 , n49346 , n49347 , n49348 , n49349 , n49350 , 
     n49351 , n49352 , n49353 , n49354 , n49355 , n49356 , n49357 , n49358 , n49359 , n49360 , 
     n49361 , n49362 , n49363 , n49364 , n49365 , n49366 , n49367 , n49368 , n49369 , n49370 , 
     n49371 , n49372 , n49373 , n49374 , n49375 , n49376 , n49377 , n49378 , n49379 , n49380 , 
     n49381 , n49382 , n49383 , n49384 , n49385 , n49386 , n49387 , n49388 , n49389 , n49390 , 
     n49391 , n49392 , n49393 , n49394 , n49395 , n49396 , n49397 , n49398 , n49399 , n49400 , 
     n49401 , n49402 , n49403 , n49404 , n49405 , n49406 , n49407 , n49408 , n49409 , n49410 , 
     n49411 , n49412 , n49413 , n49414 , n49415 , n49416 , n49417 , n49418 , n49419 , n49420 , 
     n49421 , n49422 , n49423 , n49424 , n49425 , n49426 , n49427 , n49428 , n49429 , n49430 , 
     n49431 , n49432 , n49433 , n49434 , n49435 , n49436 , n49437 , n49438 , n49439 , n49440 , 
     n49441 , n49442 , n49443 , n49444 , n49445 , n49446 , n49447 , n49448 , n49449 , n49450 , 
     n49451 , n49452 , n49453 , n49454 , n49455 , n49456 , n49457 , n49458 , n49459 , n49460 , 
     n49461 , n49462 , n49463 , n49464 , n49465 , n49466 , n49467 , n49468 , n49469 , n49470 , 
     n49471 , n49472 , n49473 , n49474 , n49475 , n49476 , n49477 , n49478 , n49479 , n49480 , 
     n49481 , n49482 , n49483 , n49484 , n49485 , n49486 , n49487 , n49488 , n49489 , n49490 , 
     n49491 , n49492 , n49493 , n49494 , n49495 , n49496 , n49497 , n49498 , n49499 , n49500 , 
     n49501 , n49502 , n49503 , n49504 , n49505 , n49506 , n49507 , n49508 , n49509 , n49510 , 
     n49511 , n49512 , n49513 , n49514 , n49515 , n49516 , n49517 , n49518 , n49519 , n49520 , 
     n49521 , n49522 , n49523 , n49524 , n49525 , n49526 , n49527 , n49528 , n49529 , n49530 , 
     n49531 , n49532 , n49533 , n49534 , n49535 , n49536 , n49537 , n49538 , n49539 , n49540 , 
     n49541 , n49542 , n49543 , n49544 , n49545 , n49546 , n49547 , n49548 , n49549 , n49550 , 
     n49551 , n49552 , n49553 , n49554 , n49555 , n49556 , n49557 , n49558 , n49559 , n49560 , 
     n49561 , n49562 , n49563 , n49564 , n49565 , n49566 , n49567 , n49568 , n49569 , n49570 , 
     n49571 , n49572 , n49573 , n49574 , n49575 , n49576 , n49577 , n49578 , n49579 , n49580 , 
     n49581 , n49582 , n49583 , n49584 , n49585 , n49586 , n49587 , n49588 , n49589 , n49590 , 
     n49591 , n49592 , n49593 , n49594 , n49595 , n49596 , n49597 , n49598 , n49599 , n49600 , 
     n49601 , n49602 , n49603 , n49604 , n49605 , n49606 , n49607 , n49608 , n49609 , n49610 , 
     n49611 , n49612 , n49613 , n49614 , n49615 , n49616 , n49617 , n49618 , n49619 , n49620 , 
     n49621 , n49622 , n49623 , n49624 , n49625 , n49626 , n49627 , n49628 , n49629 , n49630 , 
     n49631 , n49632 , n49633 , n49634 , n49635 , n49636 , n49637 , n49638 , n49639 , n49640 , 
     n49641 , n49642 , n49643 , n49644 , n49645 , n49646 , n49647 , n49648 , n49649 , n49650 , 
     n49651 , n49652 , n49653 , n49654 , n49655 , n49656 , n49657 , n49658 , n49659 , n49660 , 
     n49661 , n49662 , n49663 , n49664 , n49665 , n49666 , n49667 , n49668 , n49669 , n49670 , 
     n49671 , n49672 , n49673 , n49674 , n49675 , n49676 , n49677 , n49678 , n49679 , n49680 , 
     n49681 , n49682 , n49683 , n49684 , n49685 , n49686 , n49687 , n49688 , n49689 , n49690 , 
     n49691 , n49692 , n49693 , n49694 , n49695 , n49696 , n49697 , n49698 , n49699 , n49700 , 
     n49701 , n49702 , n49703 , n49704 , n49705 , n49706 , n49707 , n49708 , n49709 , n49710 , 
     n49711 , n49712 , n49713 , n49714 , n49715 , n49716 , n49717 , n49718 , n49719 , n49720 , 
     n49721 , n49722 , n49723 , n49724 , n49725 , n49726 , n49727 , n49728 , n49729 , n49730 , 
     n49731 , n49732 , n49733 , n49734 , n49735 , n49736 , n49737 , n49738 , n49739 , n49740 , 
     n49741 , n49742 , n49743 , n49744 , n49745 , n49746 , n49747 , n49748 , n49749 , n49750 , 
     n49751 , n49752 , n49753 , n49754 , n49755 , n49756 , n49757 , n49758 , n49759 , n49760 , 
     n49761 , n49762 , n49763 , n49764 , n49765 , n49766 , n49767 , n49768 , n49769 , n49770 , 
     n49771 , n49772 , n49773 , n49774 , n49775 , n49776 , n49777 , n49778 , n49779 , n49780 , 
     n49781 , n49782 , n49783 , n49784 , n49785 , n49786 , n49787 , n49788 , n49789 , n49790 , 
     n49791 , n49792 , n49793 , n49794 , n49795 , n49796 , n49797 , n49798 , n49799 , n49800 , 
     n49801 , n49802 , n49803 , n49804 , n49805 , n49806 , n49807 , n49808 , n49809 , n49810 , 
     n49811 , n49812 , n49813 , n49814 , n49815 , n49816 , n49817 , n49818 , n49819 , n49820 , 
     n49821 , n49822 , n49823 , n49824 , n49825 , n49826 , n49827 , n49828 , n49829 , n49830 , 
     n49831 , n49832 , n49833 , n49834 , n49835 , n49836 , n49837 , n49838 , n49839 , n49840 , 
     n49841 , n49842 , n49843 , n49844 , n49845 , n49846 , n49847 , n49848 , n49849 , n49850 , 
     n49851 , n49852 , n49853 , n49854 , n49855 , n49856 , n49857 , n49858 , n49859 , n49860 , 
     n49861 , n49862 , n49863 , n49864 , n49865 , n49866 , n49867 , n49868 , n49869 , n49870 , 
     n49871 , n49872 , n49873 , n49874 , n49875 , n49876 , n49877 , n49878 , n49879 , n49880 , 
     n49881 , n49882 , n49883 , n49884 , n49885 , n49886 , n49887 , n49888 , n49889 , n49890 , 
     n49891 , n49892 , n49893 , n49894 , n49895 , n49896 , n49897 , n49898 , n49899 , n49900 , 
     n49901 , n49902 , n49903 , n49904 , n49905 , n49906 , n49907 , n49908 , n49909 , n49910 , 
     n49911 , n49912 , n49913 , n49914 , n49915 , n49916 , n49917 , n49918 , n49919 , n49920 , 
     n49921 , n49922 , n49923 , n49924 , n49925 , n49926 , n49927 , n49928 , n49929 , n49930 , 
     n49931 , n49932 , n49933 , n49934 , n49935 , n49936 , n49937 , n49938 , n49939 , n49940 , 
     n49941 , n49942 , n49943 , n49944 , n49945 , n49946 , n49947 , n49948 , n49949 , n49950 , 
     n49951 , n49952 , n49953 , n49954 , n49955 , n49956 , n49957 , n49958 , n49959 , n49960 , 
     n49961 , n49962 , n49963 , n49964 , n49965 , n49966 , n49967 , n49968 , n49969 , n49970 , 
     n49971 , n49972 , n49973 , n49974 , n49975 , n49976 , n49977 , n49978 , n49979 , n49980 , 
     n49981 , n49982 , n49983 , n49984 , n49985 , n49986 , n49987 , n49988 , n49989 , n49990 , 
     n49991 , n49992 , n49993 , n49994 , n49995 , n49996 , n49997 , n49998 , n49999 , n50000 , 
     n50001 , n50002 , n50003 , n50004 , n50005 , n50006 , n50007 , n50008 , n50009 , n50010 , 
     n50011 , n50012 , n50013 , n50014 , n50015 , n50016 , n50017 , n50018 , n50019 , n50020 , 
     n50021 , n50022 , n50023 , n50024 , n50025 , n50026 , n50027 , n50028 , n50029 , n50030 , 
     n50031 , n50032 , n50033 , n50034 , n50035 , n50036 , n50037 , n50038 , n50039 , n50040 , 
     n50041 , n50042 , n50043 , n50044 , n50045 , n50046 , n50047 , n50048 , n50049 , n50050 , 
     n50051 , n50052 , n50053 , n50054 , n50055 , n50056 , n50057 , n50058 , n50059 , n50060 , 
     n50061 , n50062 , n50063 , n50064 , n50065 , n50066 , n50067 , n50068 , n50069 , n50070 , 
     n50071 , n50072 , n50073 , n50074 , n50075 , n50076 , n50077 , n50078 , n50079 , n50080 , 
     n50081 , n50082 , n50083 , n50084 , n50085 , n50086 , n50087 , n50088 , n50089 , n50090 , 
     n50091 , n50092 , n50093 , n50094 , n50095 , n50096 , n50097 , n50098 , n50099 , n50100 , 
     n50101 , n50102 , n50103 , n50104 , n50105 , n50106 , n50107 , n50108 , n50109 , n50110 , 
     n50111 , n50112 , n50113 , n50114 , n50115 , n50116 , n50117 , n50118 , n50119 , n50120 , 
     n50121 , n50122 , n50123 , n50124 , n50125 , n50126 , n50127 , n50128 , n50129 , n50130 , 
     n50131 , n50132 , n50133 , n50134 , n50135 , n50136 , n50137 , n50138 , n50139 , n50140 , 
     n50141 , n50142 , n50143 , n50144 , n50145 , n50146 , n50147 , n50148 , n50149 , n50150 , 
     n50151 , n50152 , n50153 , n50154 , n50155 , n50156 , n50157 , n50158 , n50159 , n50160 , 
     n50161 , n50162 , n50163 , n50164 , n50165 , n50166 , n50167 , n50168 , n50169 , n50170 , 
     n50171 , n50172 , n50173 , n50174 , n50175 , n50176 , n50177 , n50178 , n50179 , n50180 , 
     n50181 , n50182 , n50183 , n50184 , n50185 , n50186 , n50187 , n50188 , n50189 , n50190 , 
     n50191 , n50192 , n50193 , n50194 , n50195 , n50196 , n50197 , n50198 , n50199 , n50200 , 
     n50201 , n50202 , n50203 , n50204 , n50205 , n50206 , n50207 , n50208 , n50209 , n50210 , 
     n50211 , n50212 , n50213 , n50214 , n50215 , n50216 , n50217 , n50218 , n50219 , n50220 , 
     n50221 , n50222 , n50223 , n50224 , n50225 , n50226 , n50227 , n50228 , n50229 , n50230 , 
     n50231 , n50232 , n50233 , n50234 , n50235 , n50236 , n50237 , n50238 , n50239 , n50240 , 
     n50241 , n50242 , n50243 , n50244 , n50245 , n50246 , n50247 , n50248 , n50249 , n50250 , 
     n50251 , n50252 , n50253 , n50254 , n50255 , n50256 , n50257 , n50258 , n50259 , n50260 , 
     n50261 , n50262 , n50263 , n50264 , n50265 , n50266 , n50267 , n50268 , n50269 , n50270 , 
     n50271 , n50272 , n50273 , n50274 , n50275 , n50276 , n50277 , n50278 , n50279 , n50280 , 
     n50281 , n50282 , n50283 , n50284 , n50285 , n50286 , n50287 , n50288 , n50289 , n50290 , 
     n50291 , n50292 , n50293 , n50294 , n50295 , n50296 , n50297 , n50298 , n50299 , n50300 , 
     n50301 , n50302 , n50303 , n50304 , n50305 , n50306 , n50307 , n50308 , n50309 , n50310 , 
     n50311 , n50312 , n50313 , n50314 , n50315 , n50316 , n50317 , n50318 , n50319 , n50320 , 
     n50321 , n50322 , n50323 , n50324 , n50325 , n50326 , n50327 , n50328 , n50329 , n50330 , 
     n50331 , n50332 , n50333 , n50334 , n50335 , n50336 , n50337 , n50338 , n50339 , n50340 , 
     n50341 , n50342 , n50343 , n50344 , n50345 , n50346 , n50347 , n50348 , n50349 , n50350 , 
     n50351 , n50352 , n50353 , n50354 , n50355 , n50356 , n50357 , n50358 , n50359 , n50360 , 
     n50361 , n50362 , n50363 , n50364 , n50365 , n50366 , n50367 , n50368 , n50369 , n50370 , 
     n50371 , n50372 , n50373 , n50374 , n50375 , n50376 , n50377 , n50378 , n50379 , n50380 , 
     n50381 , n50382 , n50383 , n50384 , n50385 , n50386 , n50387 , n50388 , n50389 , n50390 , 
     n50391 , n50392 , n50393 , n50394 , n50395 , n50396 , n50397 , n50398 , n50399 , n50400 , 
     n50401 , n50402 , n50403 , n50404 , n50405 , n50406 , n50407 , n50408 , n50409 , n50410 , 
     n50411 , n50412 , n50413 , n50414 , n50415 , n50416 , n50417 , n50418 , n50419 , n50420 , 
     n50421 , n50422 , n50423 , n50424 , n50425 , n50426 , n50427 , n50428 , n50429 , n50430 , 
     n50431 , n50432 , n50433 , n50434 , n50435 , n50436 , n50437 , n50438 , n50439 , n50440 , 
     n50441 , n50442 , n50443 , n50444 , n50445 , n50446 , n50447 , n50448 , n50449 , n50450 , 
     n50451 , n50452 , n50453 , n50454 , n50455 , n50456 , n50457 , n50458 , n50459 , n50460 , 
     n50461 , n50462 , n50463 , n50464 , n50465 , n50466 , n50467 , n50468 , n50469 , n50470 , 
     n50471 , n50472 , n50473 , n50474 , n50475 , n50476 , n50477 , n50478 , n50479 , n50480 , 
     n50481 , n50482 , n50483 , n50484 , n50485 , n50486 , n50487 , n50488 , n50489 , n50490 , 
     n50491 , n50492 , n50493 , n50494 , n50495 , n50496 , n50497 , n50498 , n50499 , n50500 , 
     n50501 , n50502 , n50503 , n50504 , n50505 , n50506 , n50507 , n50508 , n50509 , n50510 , 
     n50511 , n50512 , n50513 , n50514 , n50515 , n50516 , n50517 , n50518 , n50519 , n50520 , 
     n50521 , n50522 , n50523 , n50524 , n50525 , n50526 , n50527 , n50528 , n50529 , n50530 , 
     n50531 , n50532 , n50533 , n50534 , n50535 , n50536 , n50537 , n50538 , n50539 , n50540 , 
     n50541 , n50542 , n50543 , n50544 , n50545 , n50546 , n50547 , n50548 , n50549 , n50550 , 
     n50551 , n50552 , n50553 , n50554 , n50555 , n50556 , n50557 , n50558 , n50559 , n50560 , 
     n50561 , n50562 , n50563 , n50564 , n50565 , n50566 , n50567 , n50568 , n50569 , n50570 , 
     n50571 , n50572 , n50573 , n50574 , n50575 , n50576 , n50577 , n50578 , n50579 , n50580 , 
     n50581 , n50582 , n50583 , n50584 , n50585 , n50586 , n50587 , n50588 , n50589 , n50590 , 
     n50591 , n50592 , n50593 , n50594 , n50595 , n50596 , n50597 , n50598 , n50599 , n50600 , 
     n50601 , n50602 , n50603 , n50604 , n50605 , n50606 , n50607 , n50608 , n50609 , n50610 , 
     n50611 , n50612 , n50613 , n50614 , n50615 , n50616 , n50617 , n50618 , n50619 , n50620 , 
     n50621 , n50622 , n50623 , n50624 , n50625 , n50626 , n50627 , n50628 , n50629 , n50630 , 
     n50631 , n50632 , n50633 , n50634 , n50635 , n50636 , n50637 , n50638 , n50639 , n50640 , 
     n50641 , n50642 , n50643 , n50644 , n50645 , n50646 , n50647 , n50648 , n50649 , n50650 , 
     n50651 , n50652 , n50653 , n50654 , n50655 , n50656 , n50657 , n50658 , n50659 , n50660 , 
     n50661 , n50662 , n50663 , n50664 , n50665 , n50666 , n50667 , n50668 , n50669 , n50670 , 
     n50671 , n50672 , n50673 , n50674 , n50675 , n50676 , n50677 , n50678 , n50679 , n50680 , 
     n50681 , n50682 , n50683 , n50684 , n50685 , n50686 , n50687 , n50688 , n50689 , n50690 , 
     n50691 , n50692 , n50693 , n50694 , n50695 , n50696 , n50697 , n50698 , n50699 , n50700 , 
     n50701 , n50702 , n50703 , n50704 , n50705 , n50706 , n50707 , n50708 , n50709 , n50710 , 
     n50711 , n50712 , n50713 , n50714 , n50715 , n50716 , n50717 , n50718 , n50719 , n50720 , 
     n50721 , n50722 , n50723 , n50724 , n50725 , n50726 , n50727 , n50728 , n50729 , n50730 , 
     n50731 , n50732 , n50733 , n50734 , n50735 , n50736 , n50737 , n50738 , n50739 , n50740 , 
     n50741 , n50742 , n50743 , n50744 , n50745 , n50746 , n50747 , n50748 , n50749 , n50750 , 
     n50751 , n50752 , n50753 , n50754 , n50755 , n50756 , n50757 , n50758 , n50759 , n50760 , 
     n50761 , n50762 , n50763 , n50764 , n50765 , n50766 , n50767 , n50768 , n50769 , n50770 , 
     n50771 , n50772 , n50773 , n50774 , n50775 , n50776 , n50777 , n50778 , n50779 , n50780 , 
     n50781 , n50782 , n50783 , n50784 , n50785 , n50786 , n50787 , n50788 , n50789 , n50790 , 
     n50791 , n50792 , n50793 , n50794 , n50795 , n50796 , n50797 , n50798 , n50799 , n50800 , 
     n50801 , n50802 , n50803 , n50804 , n50805 , n50806 , n50807 , n50808 , n50809 , n50810 , 
     n50811 , n50812 , n50813 , n50814 , n50815 , n50816 , n50817 , n50818 , n50819 , n50820 , 
     n50821 , n50822 , n50823 , n50824 , n50825 , n50826 , n50827 , n50828 , n50829 , n50830 , 
     n50831 , n50832 , n50833 , n50834 , n50835 , n50836 , n50837 , n50838 , n50839 , n50840 , 
     n50841 , n50842 , n50843 , n50844 , n50845 , n50846 , n50847 , n50848 , n50849 , n50850 , 
     n50851 , n50852 , n50853 , n50854 , n50855 , n50856 , n50857 , n50858 , n50859 , n50860 , 
     n50861 , n50862 , n50863 , n50864 , n50865 , n50866 , n50867 , n50868 , n50869 , n50870 , 
     n50871 , n50872 , n50873 , n50874 , n50875 , n50876 , n50877 , n50878 , n50879 , n50880 , 
     n50881 , n50882 , n50883 , n50884 , n50885 , n50886 , n50887 , n50888 , n50889 , n50890 , 
     n50891 , n50892 , n50893 , n50894 , n50895 , n50896 , n50897 , n50898 , n50899 , n50900 , 
     n50901 , n50902 , n50903 , n50904 , n50905 , n50906 , n50907 , n50908 , n50909 , n50910 , 
     n50911 , n50912 , n50913 , n50914 , n50915 , n50916 , n50917 , n50918 , n50919 , n50920 , 
     n50921 , n50922 , n50923 , n50924 , n50925 , n50926 , n50927 , n50928 , n50929 , n50930 , 
     n50931 , n50932 , n50933 , n50934 , n50935 , n50936 , n50937 , n50938 , n50939 , n50940 , 
     n50941 , n50942 , n50943 , n50944 , n50945 , n50946 , n50947 , n50948 , n50949 , n50950 , 
     n50951 , n50952 , n50953 , n50954 , n50955 , n50956 , n50957 , n50958 , n50959 , n50960 , 
     n50961 , n50962 , n50963 , n50964 , n50965 , n50966 , n50967 , n50968 , n50969 , n50970 , 
     n50971 , n50972 , n50973 , n50974 , n50975 , n50976 , n50977 , n50978 , n50979 , n50980 , 
     n50981 , n50982 , n50983 , n50984 , n50985 , n50986 , n50987 , n50988 , n50989 , n50990 , 
     n50991 , n50992 , n50993 , n50994 , n50995 , n50996 , n50997 , n50998 , n50999 , n51000 , 
     n51001 , n51002 , n51003 , n51004 , n51005 , n51006 , n51007 , n51008 , n51009 , n51010 , 
     n51011 , n51012 , n51013 , n51014 , n51015 , n51016 , n51017 , n51018 , n51019 , n51020 , 
     n51021 , n51022 , n51023 , n51024 , n51025 , n51026 , n51027 , n51028 , n51029 , n51030 , 
     n51031 , n51032 , n51033 , n51034 , n51035 , n51036 , n51037 , n51038 , n51039 , n51040 , 
     n51041 , n51042 , n51043 , n51044 , n51045 , n51046 , n51047 , n51048 , n51049 , n51050 , 
     n51051 , n51052 , n51053 , n51054 , n51055 , n51056 , n51057 , n51058 , n51059 , n51060 , 
     n51061 , n51062 , n51063 , n51064 , n51065 , n51066 , n51067 , n51068 , n51069 , n51070 , 
     n51071 , n51072 , n51073 , n51074 , n51075 , n51076 , n51077 , n51078 , n51079 , n51080 , 
     n51081 , n51082 , n51083 , n51084 , n51085 , n51086 , n51087 , n51088 , n51089 , n51090 , 
     n51091 , n51092 , n51093 , n51094 , n51095 , n51096 , n51097 , n51098 , n51099 , n51100 , 
     n51101 , n51102 , n51103 , n51104 , n51105 , n51106 , n51107 , n51108 , n51109 , n51110 , 
     n51111 , n51112 , n51113 , n51114 , n51115 , n51116 , n51117 , n51118 , n51119 , n51120 , 
     n51121 , n51122 , n51123 , n51124 , n51125 , n51126 , n51127 , n51128 , n51129 , n51130 , 
     n51131 , n51132 , n51133 , n51134 , n51135 , n51136 , n51137 , n51138 , n51139 , n51140 , 
     n51141 , n51142 , n51143 , n51144 , n51145 , n51146 , n51147 , n51148 , n51149 , n51150 , 
     n51151 , n51152 , n51153 , n51154 , n51155 , n51156 , n51157 , n51158 , n51159 , n51160 , 
     n51161 , n51162 , n51163 , n51164 , n51165 , n51166 , n51167 , n51168 , n51169 , n51170 , 
     n51171 , n51172 , n51173 , n51174 , n51175 , n51176 , n51177 , n51178 , n51179 , n51180 , 
     n51181 , n51182 , n51183 , n51184 , n51185 , n51186 , n51187 , n51188 , n51189 , n51190 , 
     n51191 , n51192 , n51193 , n51194 , n51195 , n51196 , n51197 , n51198 , n51199 , n51200 , 
     n51201 , n51202 , n51203 , n51204 , n51205 , n51206 , n51207 , n51208 , n51209 , n51210 , 
     n51211 , n51212 , n51213 , n51214 , n51215 , n51216 , n51217 , n51218 , n51219 , n51220 , 
     n51221 , n51222 , n51223 , n51224 , n51225 , n51226 , n51227 , n51228 , n51229 , n51230 , 
     n51231 , n51232 , n51233 , n51234 , n51235 , n51236 , n51237 , n51238 , n51239 , n51240 , 
     n51241 , n51242 , n51243 , n51244 , n51245 , n51246 , n51247 , n51248 , n51249 , n51250 , 
     n51251 , n51252 , n51253 , n51254 , n51255 , n51256 , n51257 , n51258 , n51259 , n51260 , 
     n51261 , n51262 , n51263 , n51264 , n51265 , n51266 , n51267 , n51268 , n51269 , n51270 , 
     n51271 , n51272 , n51273 , n51274 , n51275 , n51276 , n51277 , n51278 , n51279 , n51280 , 
     n51281 , n51282 , n51283 , n51284 , n51285 , n51286 , n51287 , n51288 , n51289 , n51290 , 
     n51291 , n51292 , n51293 , n51294 , n51295 , n51296 , n51297 , n51298 , n51299 , n51300 , 
     n51301 , n51302 , n51303 , n51304 , n51305 , n51306 , n51307 , n51308 , n51309 , n51310 , 
     n51311 , n51312 , n51313 , n51314 , n51315 , n51316 , n51317 , n51318 , n51319 , n51320 , 
     n51321 , n51322 , n51323 , n51324 , n51325 , n51326 , n51327 , n51328 , n51329 , n51330 , 
     n51331 , n51332 , n51333 , n51334 , n51335 , n51336 , n51337 , n51338 , n51339 , n51340 , 
     n51341 , n51342 , n51343 , n51344 , n51345 , n51346 , n51347 , n51348 , n51349 , n51350 , 
     n51351 , n51352 , n51353 , n51354 , n51355 , n51356 , n51357 , n51358 , n51359 , n51360 , 
     n51361 , n51362 , n51363 , n51364 , n51365 , n51366 , n51367 , n51368 , n51369 , n51370 , 
     n51371 , n51372 , n51373 , n51374 , n51375 , n51376 , n51377 , n51378 , n51379 , n51380 , 
     n51381 , n51382 , n51383 , n51384 , n51385 , n51386 , n51387 , n51388 , n51389 , n51390 , 
     n51391 , n51392 , n51393 , n51394 , n51395 , n51396 , n51397 , n51398 , n51399 , n51400 , 
     n51401 , n51402 , n51403 , n51404 , n51405 , n51406 , n51407 , n51408 , n51409 , n51410 , 
     n51411 , n51412 , n51413 , n51414 , n51415 , n51416 , n51417 , n51418 , n51419 , n51420 , 
     n51421 , n51422 , n51423 , n51424 , n51425 , n51426 , n51427 , n51428 , n51429 , n51430 , 
     n51431 , n51432 , n51433 , n51434 , n51435 , n51436 , n51437 , n51438 , n51439 , n51440 , 
     n51441 , n51442 , n51443 , n51444 , n51445 , n51446 , n51447 , n51448 , n51449 , n51450 , 
     n51451 , n51452 , n51453 , n51454 , n51455 , n51456 , n51457 , n51458 , n51459 , n51460 , 
     n51461 , n51462 , n51463 , n51464 , n51465 , n51466 , n51467 , n51468 , n51469 , n51470 , 
     n51471 , n51472 , n51473 , n51474 , n51475 , n51476 , n51477 , n51478 , n51479 , n51480 , 
     n51481 , n51482 , n51483 , n51484 , n51485 , n51486 , n51487 , n51488 , n51489 , n51490 , 
     n51491 , n51492 , n51493 , n51494 , n51495 , n51496 , n51497 , n51498 , n51499 , n51500 , 
     n51501 , n51502 , n51503 , n51504 , n51505 , n51506 , n51507 , n51508 , n51509 , n51510 , 
     n51511 , n51512 , n51513 , n51514 , n51515 , n51516 , n51517 , n51518 , n51519 , n51520 , 
     n51521 , n51522 , n51523 , n51524 , n51525 , n51526 , n51527 , n51528 , n51529 , n51530 , 
     n51531 , n51532 , n51533 , n51534 , n51535 , n51536 , n51537 , n51538 , n51539 , n51540 , 
     n51541 , n51542 , n51543 , n51544 , n51545 , n51546 , n51547 , n51548 , n51549 , n51550 , 
     n51551 , n51552 , n51553 , n51554 , n51555 , n51556 , n51557 , n51558 , n51559 , n51560 , 
     n51561 , n51562 , n51563 , n51564 , n51565 , n51566 , n51567 , n51568 , n51569 , n51570 , 
     n51571 , n51572 , n51573 , n51574 , n51575 , n51576 , n51577 , n51578 , n51579 , n51580 , 
     n51581 , n51582 , n51583 , n51584 , n51585 , n51586 , n51587 , n51588 , n51589 , n51590 , 
     n51591 , n51592 , n51593 , n51594 , n51595 , n51596 , n51597 , n51598 , n51599 , n51600 , 
     n51601 , n51602 , n51603 , n51604 , n51605 , n51606 , n51607 , n51608 , n51609 , n51610 , 
     n51611 , n51612 , n51613 , n51614 , n51615 , n51616 , n51617 , n51618 , n51619 , n51620 , 
     n51621 , n51622 , n51623 , n51624 , n51625 , n51626 , n51627 , n51628 , n51629 , n51630 , 
     n51631 , n51632 , n51633 , n51634 , n51635 , n51636 , n51637 , n51638 , n51639 , n51640 , 
     n51641 , n51642 , n51643 , n51644 , n51645 , n51646 , n51647 , n51648 , n51649 , n51650 , 
     n51651 , n51652 , n51653 , n51654 , n51655 , n51656 , n51657 , n51658 , n51659 , n51660 , 
     n51661 , n51662 , n51663 , n51664 , n51665 , n51666 , n51667 , n51668 , n51669 , n51670 , 
     n51671 , n51672 , n51673 , n51674 , n51675 , n51676 , n51677 , n51678 , n51679 , n51680 , 
     n51681 , n51682 , n51683 , n51684 , n51685 , n51686 , n51687 , n51688 , n51689 , n51690 , 
     n51691 , n51692 , n51693 , n51694 , n51695 , n51696 , n51697 , n51698 , n51699 , n51700 , 
     n51701 , n51702 , n51703 , n51704 , n51705 , n51706 , n51707 , n51708 , n51709 , n51710 , 
     n51711 , n51712 , n51713 , n51714 , n51715 , n51716 , n51717 , n51718 , n51719 , n51720 , 
     n51721 , n51722 , n51723 , n51724 , n51725 , n51726 , n51727 , n51728 , n51729 , n51730 , 
     n51731 , n51732 , n51733 , n51734 , n51735 , n51736 , n51737 , n51738 , n51739 , n51740 , 
     n51741 , n51742 , n51743 , n51744 , n51745 , n51746 , n51747 , n51748 , n51749 , n51750 , 
     n51751 , n51752 , n51753 , n51754 , n51755 , n51756 , n51757 , n51758 , n51759 , n51760 , 
     n51761 , n51762 , n51763 , n51764 , n51765 , n51766 , n51767 , n51768 , n51769 , n51770 , 
     n51771 , n51772 , n51773 , n51774 , n51775 , n51776 , n51777 , n51778 , n51779 , n51780 , 
     n51781 , n51782 , n51783 , n51784 , n51785 , n51786 , n51787 , n51788 , n51789 , n51790 , 
     n51791 , n51792 , n51793 , n51794 , n51795 , n51796 , n51797 , n51798 , n51799 , n51800 , 
     n51801 , n51802 , n51803 , n51804 , n51805 , n51806 , n51807 , n51808 , n51809 , n51810 , 
     n51811 , n51812 , n51813 , n51814 , n51815 , n51816 , n51817 , n51818 , n51819 , n51820 , 
     n51821 , n51822 , n51823 , n51824 , n51825 , n51826 , n51827 , n51828 , n51829 , n51830 , 
     n51831 , n51832 , n51833 , n51834 , n51835 , n51836 , n51837 , n51838 , n51839 , n51840 , 
     n51841 , n51842 , n51843 , n51844 , n51845 , n51846 , n51847 , n51848 , n51849 , n51850 , 
     n51851 , n51852 , n51853 , n51854 , n51855 , n51856 , n51857 , n51858 , n51859 , n51860 , 
     n51861 , n51862 , n51863 , n51864 , n51865 , n51866 , n51867 , n51868 , n51869 , n51870 , 
     n51871 , n51872 , n51873 , n51874 , n51875 , n51876 , n51877 , n51878 , n51879 , n51880 , 
     n51881 , n51882 , n51883 , n51884 , n51885 , n51886 , n51887 , n51888 , n51889 , n51890 , 
     n51891 , n51892 , n51893 , n51894 , n51895 , n51896 , n51897 , n51898 , n51899 , n51900 , 
     n51901 , n51902 , n51903 , n51904 , n51905 , n51906 , n51907 , n51908 , n51909 , n51910 , 
     n51911 , n51912 , n51913 , n51914 , n51915 , n51916 , n51917 , n51918 , n51919 , n51920 , 
     n51921 , n51922 , n51923 , n51924 , n51925 , n51926 , n51927 , n51928 , n51929 , n51930 , 
     n51931 , n51932 , n51933 , n51934 , n51935 , n51936 , n51937 , n51938 , n51939 , n51940 , 
     n51941 , n51942 , n51943 , n51944 , n51945 , n51946 , n51947 , n51948 , n51949 , n51950 , 
     n51951 , n51952 , n51953 , n51954 , n51955 , n51956 , n51957 , n51958 , n51959 , n51960 , 
     n51961 , n51962 , n51963 , n51964 , n51965 , n51966 , n51967 , n51968 , n51969 , n51970 , 
     n51971 , n51972 , n51973 , n51974 , n51975 , n51976 , n51977 , n51978 , n51979 , n51980 , 
     n51981 , n51982 , n51983 , n51984 , n51985 , n51986 , n51987 , n51988 , n51989 , n51990 , 
     n51991 , n51992 , n51993 , n51994 , n51995 , n51996 , n51997 , n51998 , n51999 , n52000 , 
     n52001 , n52002 , n52003 , n52004 , n52005 , n52006 , n52007 , n52008 , n52009 , n52010 , 
     n52011 , n52012 , n52013 , n52014 , n52015 , n52016 , n52017 , n52018 , n52019 , n52020 , 
     n52021 , n52022 , n52023 , n52024 , n52025 , n52026 , n52027 , n52028 , n52029 , n52030 , 
     n52031 , n52032 , n52033 , n52034 , n52035 , n52036 , n52037 , n52038 , n52039 , n52040 , 
     n52041 , n52042 , n52043 , n52044 , n52045 , n52046 , n52047 , n52048 , n52049 , n52050 , 
     n52051 , n52052 , n52053 , n52054 , n52055 , n52056 , n52057 , n52058 , n52059 , n52060 , 
     n52061 , n52062 , n52063 , n52064 , n52065 , n52066 , n52067 , n52068 , n52069 , n52070 , 
     n52071 , n52072 , n52073 , n52074 , n52075 , n52076 , n52077 , n52078 , n52079 , n52080 , 
     n52081 , n52082 , n52083 , n52084 , n52085 , n52086 , n52087 , n52088 , n52089 , n52090 , 
     n52091 , n52092 , n52093 , n52094 , n52095 , n52096 , n52097 , n52098 , n52099 , n52100 , 
     n52101 , n52102 , n52103 , n52104 , n52105 , n52106 , n52107 , n52108 , n52109 , n52110 , 
     n52111 , n52112 , n52113 , n52114 , n52115 , n52116 , n52117 , n52118 , n52119 , n52120 , 
     n52121 , n52122 , n52123 , n52124 , n52125 , n52126 , n52127 , n52128 , n52129 , n52130 , 
     n52131 , n52132 , n52133 , n52134 , n52135 , n52136 , n52137 , n52138 , n52139 , n52140 , 
     n52141 , n52142 , n52143 , n52144 , n52145 , n52146 , n52147 , n52148 , n52149 , n52150 , 
     n52151 , n52152 , n52153 , n52154 , n52155 , n52156 , n52157 , n52158 , n52159 , n52160 , 
     n52161 , n52162 , n52163 , n52164 , n52165 , n52166 , n52167 , n52168 , n52169 , n52170 , 
     n52171 , n52172 , n52173 , n52174 , n52175 , n52176 , n52177 , n52178 , n52179 , n52180 , 
     n52181 , n52182 , n52183 , n52184 , n52185 , n52186 , n52187 , n52188 , n52189 , n52190 , 
     n52191 , n52192 , n52193 , n52194 , n52195 , n52196 , n52197 , n52198 , n52199 , n52200 , 
     n52201 , n52202 , n52203 , n52204 , n52205 , n52206 , n52207 , n52208 , n52209 , n52210 , 
     n52211 , n52212 , n52213 , n52214 , n52215 , n52216 , n52217 , n52218 , n52219 , n52220 , 
     n52221 , n52222 , n52223 , n52224 , n52225 , n52226 , n52227 , n52228 , n52229 , n52230 , 
     n52231 , n52232 , n52233 , n52234 , n52235 , n52236 , n52237 , n52238 , n52239 , n52240 , 
     n52241 , n52242 , n52243 , n52244 , n52245 , n52246 , n52247 , n52248 , n52249 , n52250 , 
     n52251 , n52252 , n52253 , n52254 , n52255 , n52256 , n52257 , n52258 , n52259 , n52260 , 
     n52261 , n52262 , n52263 , n52264 , n52265 , n52266 , n52267 , n52268 , n52269 , n52270 , 
     n52271 , n52272 , n52273 , n52274 , n52275 , n52276 , n52277 , n52278 , n52279 , n52280 , 
     n52281 , n52282 , n52283 , n52284 , n52285 , n52286 , n52287 , n52288 , n52289 , n52290 , 
     n52291 , n52292 , n52293 , n52294 , n52295 , n52296 , n52297 , n52298 , n52299 , n52300 , 
     n52301 , n52302 , n52303 , n52304 , n52305 , n52306 , n52307 , n52308 , n52309 , n52310 , 
     n52311 , n52312 , n52313 , n52314 , n52315 , n52316 , n52317 , n52318 , n52319 , n52320 , 
     n52321 , n52322 , n52323 , n52324 , n52325 , n52326 , n52327 , n52328 , n52329 , n52330 , 
     n52331 , n52332 , n52333 , n52334 , n52335 , n52336 , n52337 , n52338 , n52339 , n52340 , 
     n52341 , n52342 , n52343 , n52344 , n52345 , n52346 , n52347 , n52348 , n52349 , n52350 , 
     n52351 , n52352 , n52353 , n52354 , n52355 , n52356 , n52357 , n52358 , n52359 , n52360 , 
     n52361 , n52362 , n52363 , n52364 , n52365 , n52366 , n52367 , n52368 , n52369 , n52370 , 
     n52371 , n52372 , n52373 , n52374 , n52375 , n52376 , n52377 , n52378 , n52379 , n52380 , 
     n52381 , n52382 , n52383 , n52384 , n52385 , n52386 , n52387 , n52388 , n52389 , n52390 , 
     n52391 , n52392 , n52393 , n52394 , n52395 , n52396 , n52397 , n52398 , n52399 , n52400 , 
     n52401 , n52402 , n52403 , n52404 , n52405 , n52406 , n52407 , n52408 , n52409 , n52410 , 
     n52411 , n52412 , n52413 , n52414 , n52415 , n52416 , n52417 , n52418 , n52419 , n52420 , 
     n52421 , n52422 , n52423 , n52424 , n52425 , n52426 , n52427 , n52428 , n52429 , n52430 , 
     n52431 , n52432 , n52433 , n52434 , n52435 , n52436 , n52437 , n52438 , n52439 , n52440 , 
     n52441 , n52442 , n52443 , n52444 , n52445 , n52446 , n52447 , n52448 , n52449 , n52450 , 
     n52451 , n52452 , n52453 , n52454 , n52455 , n52456 , n52457 , n52458 , n52459 , n52460 , 
     n52461 , n52462 , n52463 , n52464 , n52465 , n52466 , n52467 , n52468 , n52469 , n52470 , 
     n52471 , n52472 , n52473 , n52474 , n52475 , n52476 , n52477 , n52478 , n52479 , n52480 , 
     n52481 , n52482 , n52483 , n52484 , n52485 , n52486 , n52487 , n52488 , n52489 , n52490 , 
     n52491 , n52492 , n52493 , n52494 , n52495 , n52496 , n52497 , n52498 , n52499 , n52500 , 
     n52501 , n52502 , n52503 , n52504 , n52505 , n52506 , n52507 , n52508 , n52509 , n52510 , 
     n52511 , n52512 , n52513 , n52514 , n52515 , n52516 , n52517 , n52518 , n52519 , n52520 , 
     n52521 , n52522 , n52523 , n52524 , n52525 , n52526 , n52527 , n52528 , n52529 , n52530 , 
     n52531 , n52532 , n52533 , n52534 , n52535 , n52536 , n52537 , n52538 , n52539 , n52540 , 
     n52541 , n52542 , n52543 , n52544 , n52545 , n52546 , n52547 , n52548 , n52549 , n52550 , 
     n52551 , n52552 , n52553 , n52554 , n52555 , n52556 , n52557 , n52558 , n52559 , n52560 , 
     n52561 , n52562 , n52563 , n52564 , n52565 , n52566 , n52567 , n52568 , n52569 , n52570 , 
     n52571 , n52572 , n52573 , n52574 , n52575 , n52576 , n52577 , n52578 , n52579 , n52580 , 
     n52581 , n52582 , n52583 , n52584 , n52585 , n52586 , n52587 , n52588 , n52589 , n52590 , 
     n52591 , n52592 , n52593 , n52594 , n52595 , n52596 , n52597 , n52598 , n52599 , n52600 , 
     n52601 , n52602 , n52603 , n52604 , n52605 , n52606 , n52607 , n52608 , n52609 , n52610 , 
     n52611 , n52612 , n52613 , n52614 , n52615 , n52616 , n52617 , n52618 , n52619 , n52620 , 
     n52621 , n52622 , n52623 , n52624 , n52625 , n52626 , n52627 , n52628 , n52629 , n52630 , 
     n52631 , n52632 , n52633 , n52634 , n52635 , n52636 , n52637 , n52638 , n52639 , n52640 , 
     n52641 , n52642 , n52643 , n52644 , n52645 , n52646 , n52647 , n52648 , n52649 , n52650 , 
     n52651 , n52652 , n52653 , n52654 , n52655 , n52656 , n52657 , n52658 , n52659 , n52660 , 
     n52661 , n52662 , n52663 , n52664 , n52665 , n52666 , n52667 , n52668 , n52669 , n52670 , 
     n52671 , n52672 , n52673 , n52674 , n52675 , n52676 , n52677 , n52678 , n52679 , n52680 , 
     n52681 , n52682 , n52683 , n52684 , n52685 , n52686 , n52687 , n52688 , n52689 , n52690 , 
     n52691 , n52692 , n52693 , n52694 , n52695 , n52696 , n52697 , n52698 , n52699 , n52700 , 
     n52701 , n52702 , n52703 , n52704 , n52705 , n52706 , n52707 , n52708 , n52709 , n52710 , 
     n52711 , n52712 , n52713 , n52714 , n52715 , n52716 , n52717 , n52718 , n52719 , n52720 , 
     n52721 , n52722 , n52723 , n52724 , n52725 , n52726 , n52727 , n52728 , n52729 , n52730 , 
     n52731 , n52732 , n52733 , n52734 , n52735 , n52736 , n52737 , n52738 , n52739 , n52740 , 
     n52741 , n52742 , n52743 , n52744 , n52745 , n52746 , n52747 , n52748 , n52749 , n52750 , 
     n52751 , n52752 , n52753 , n52754 , n52755 , n52756 , n52757 , n52758 , n52759 , n52760 , 
     n52761 , n52762 , n52763 , n52764 , n52765 , n52766 , n52767 , n52768 , n52769 , n52770 , 
     n52771 , n52772 , n52773 , n52774 , n52775 , n52776 , n52777 , n52778 , n52779 , n52780 , 
     n52781 , n52782 , n52783 , n52784 , n52785 , n52786 , n52787 , n52788 , n52789 , n52790 , 
     n52791 , n52792 , n52793 , n52794 , n52795 , n52796 , n52797 , n52798 , n52799 , n52800 , 
     n52801 , n52802 , n52803 , n52804 , n52805 , n52806 , n52807 , n52808 , n52809 , n52810 , 
     n52811 , n52812 , n52813 , n52814 , n52815 , n52816 , n52817 , n52818 , n52819 , n52820 , 
     n52821 , n52822 , n52823 , n52824 , n52825 , n52826 , n52827 , n52828 , n52829 , n52830 , 
     n52831 , n52832 , n52833 , n52834 , n52835 , n52836 , n52837 , n52838 , n52839 , n52840 , 
     n52841 , n52842 , n52843 , n52844 , n52845 , n52846 , n52847 , n52848 , n52849 , n52850 , 
     n52851 , n52852 , n52853 , n52854 , n52855 , n52856 , n52857 , n52858 , n52859 , n52860 , 
     n52861 , n52862 , n52863 , n52864 , n52865 , n52866 , n52867 , n52868 , n52869 , n52870 , 
     n52871 , n52872 , n52873 , n52874 , n52875 , n52876 , n52877 , n52878 , n52879 , n52880 , 
     n52881 , n52882 , n52883 , n52884 , n52885 , n52886 , n52887 , n52888 , n52889 , n52890 , 
     n52891 , n52892 , n52893 , n52894 , n52895 , n52896 , n52897 , n52898 , n52899 , n52900 , 
     n52901 , n52902 , n52903 , n52904 , n52905 , n52906 , n52907 , n52908 , n52909 , n52910 , 
     n52911 , n52912 , n52913 , n52914 , n52915 , n52916 , n52917 , n52918 , n52919 , n52920 , 
     n52921 , n52922 , n52923 , n52924 , n52925 , n52926 , n52927 , n52928 , n52929 , n52930 , 
     n52931 , n52932 , n52933 , n52934 , n52935 , n52936 , n52937 , n52938 , n52939 , n52940 , 
     n52941 , n52942 , n52943 , n52944 , n52945 , n52946 , n52947 , n52948 , n52949 , n52950 , 
     n52951 , n52952 , n52953 , n52954 , n52955 , n52956 , n52957 , n52958 , n52959 , n52960 , 
     n52961 , n52962 , n52963 , n52964 , n52965 , n52966 , n52967 , n52968 , n52969 , n52970 , 
     n52971 , n52972 , n52973 , n52974 , n52975 , n52976 , n52977 , n52978 , n52979 , n52980 , 
     n52981 , n52982 , n52983 , n52984 , n52985 , n52986 , n52987 , n52988 , n52989 , n52990 , 
     n52991 , n52992 , n52993 , n52994 , n52995 , n52996 , n52997 , n52998 , n52999 , n53000 , 
     n53001 , n53002 , n53003 , n53004 , n53005 , n53006 , n53007 , n53008 , n53009 , n53010 , 
     n53011 , n53012 , n53013 , n53014 , n53015 , n53016 , n53017 , n53018 , n53019 , n53020 , 
     n53021 , n53022 , n53023 , n53024 , n53025 , n53026 , n53027 , n53028 , n53029 , n53030 , 
     n53031 , n53032 , n53033 , n53034 , n53035 , n53036 , n53037 , n53038 , n53039 , n53040 , 
     n53041 , n53042 , n53043 , n53044 , n53045 , n53046 , n53047 , n53048 , n53049 , n53050 , 
     n53051 , n53052 , n53053 , n53054 , n53055 , n53056 , n53057 , n53058 , n53059 , n53060 , 
     n53061 , n53062 , n53063 , n53064 , n53065 , n53066 , n53067 , n53068 , n53069 , n53070 , 
     n53071 , n53072 , n53073 , n53074 , n53075 , n53076 , n53077 , n53078 , n53079 , n53080 , 
     n53081 , n53082 , n53083 , n53084 , n53085 , n53086 , n53087 , n53088 , n53089 , n53090 , 
     n53091 , n53092 , n53093 , n53094 , n53095 , n53096 , n53097 , n53098 , n53099 , n53100 , 
     n53101 , n53102 , n53103 , n53104 , n53105 , n53106 , n53107 , n53108 , n53109 , n53110 , 
     n53111 , n53112 , n53113 , n53114 , n53115 , n53116 , n53117 , n53118 , n53119 , n53120 , 
     n53121 , n53122 , n53123 , n53124 , n53125 , n53126 , n53127 , n53128 , n53129 , n53130 , 
     n53131 , n53132 , n53133 , n53134 , n53135 , n53136 , n53137 , n53138 , n53139 , n53140 , 
     n53141 , n53142 , n53143 , n53144 , n53145 , n53146 , n53147 , n53148 , n53149 , n53150 , 
     n53151 , n53152 , n53153 , n53154 , n53155 , n53156 , n53157 , n53158 , n53159 , n53160 , 
     n53161 , n53162 , n53163 , n53164 , n53165 , n53166 , n53167 , n53168 , n53169 , n53170 , 
     n53171 , n53172 , n53173 , n53174 , n53175 , n53176 , n53177 , n53178 , n53179 , n53180 , 
     n53181 , n53182 , n53183 , n53184 , n53185 , n53186 , n53187 , n53188 , n53189 , n53190 , 
     n53191 , n53192 , n53193 , n53194 , n53195 , n53196 , n53197 , n53198 , n53199 , n53200 , 
     n53201 , n53202 , n53203 , n53204 , n53205 , n53206 , n53207 , n53208 , n53209 , n53210 , 
     n53211 , n53212 , n53213 , n53214 , n53215 , n53216 , n53217 , n53218 , n53219 , n53220 , 
     n53221 , n53222 , n53223 , n53224 , n53225 , n53226 , n53227 , n53228 , n53229 , n53230 , 
     n53231 , n53232 , n53233 , n53234 , n53235 , n53236 , n53237 , n53238 , n53239 , n53240 , 
     n53241 , n53242 , n53243 , n53244 , n53245 , n53246 , n53247 , n53248 , n53249 , n53250 , 
     n53251 , n53252 , n53253 , n53254 , n53255 , n53256 , n53257 , n53258 , n53259 , n53260 , 
     n53261 , n53262 , n53263 , n53264 , n53265 , n53266 , n53267 , n53268 , n53269 , n53270 , 
     n53271 , n53272 , n53273 , n53274 , n53275 , n53276 , n53277 , n53278 , n53279 , n53280 , 
     n53281 , n53282 , n53283 , n53284 , n53285 , n53286 , n53287 , n53288 , n53289 , n53290 , 
     n53291 , n53292 , n53293 , n53294 , n53295 , n53296 , n53297 , n53298 , n53299 , n53300 , 
     n53301 , n53302 , n53303 , n53304 , n53305 , n53306 , n53307 , n53308 , n53309 , n53310 , 
     n53311 , n53312 , n53313 , n53314 , n53315 , n53316 , n53317 , n53318 , n53319 , n53320 , 
     n53321 , n53322 , n53323 , n53324 , n53325 , n53326 , n53327 , n53328 , n53329 , n53330 , 
     n53331 , n53332 , n53333 , n53334 , n53335 , n53336 , n53337 , n53338 , n53339 , n53340 , 
     n53341 , n53342 , n53343 , n53344 , n53345 , n53346 , n53347 , n53348 , n53349 , n53350 , 
     n53351 , n53352 , n53353 , n53354 , n53355 , n53356 , n53357 , n53358 , n53359 , n53360 , 
     n53361 , n53362 , n53363 , n53364 , n53365 , n53366 , n53367 , n53368 , n53369 , n53370 , 
     n53371 , n53372 , n53373 , n53374 , n53375 , n53376 , n53377 , n53378 , n53379 , n53380 , 
     n53381 , n53382 , n53383 , n53384 , n53385 , n53386 , n53387 , n53388 , n53389 , n53390 , 
     n53391 , n53392 , n53393 , n53394 , n53395 , n53396 , n53397 , n53398 , n53399 , n53400 , 
     n53401 , n53402 , n53403 , n53404 , n53405 , n53406 , n53407 , n53408 , n53409 , n53410 , 
     n53411 , n53412 , n53413 , n53414 , n53415 , n53416 , n53417 , n53418 , n53419 , n53420 , 
     n53421 , n53422 , n53423 , n53424 , n53425 , n53426 , n53427 , n53428 , n53429 , n53430 , 
     n53431 , n53432 , n53433 , n53434 , n53435 , n53436 , n53437 , n53438 , n53439 , n53440 , 
     n53441 , n53442 , n53443 , n53444 , n53445 , n53446 , n53447 , n53448 , n53449 , n53450 , 
     n53451 , n53452 , n53453 , n53454 , n53455 , n53456 , n53457 , n53458 , n53459 , n53460 , 
     n53461 , n53462 , n53463 , n53464 , n53465 , n53466 , n53467 , n53468 , n53469 , n53470 , 
     n53471 , n53472 , n53473 , n53474 , n53475 , n53476 , n53477 , n53478 , n53479 , n53480 , 
     n53481 , n53482 , n53483 , n53484 , n53485 , n53486 , n53487 , n53488 , n53489 , n53490 , 
     n53491 , n53492 , n53493 , n53494 , n53495 , n53496 , n53497 , n53498 , n53499 , n53500 , 
     n53501 , n53502 , n53503 , n53504 , n53505 , n53506 , n53507 , n53508 , n53509 , n53510 , 
     n53511 , n53512 , n53513 , n53514 , n53515 , n53516 , n53517 , n53518 , n53519 , n53520 , 
     n53521 , n53522 , n53523 , n53524 , n53525 , n53526 , n53527 , n53528 , n53529 , n53530 , 
     n53531 , n53532 , n53533 , n53534 , n53535 , n53536 , n53537 , n53538 , n53539 , n53540 , 
     n53541 , n53542 , n53543 , n53544 , n53545 , n53546 , n53547 , n53548 , n53549 , n53550 , 
     n53551 , n53552 , n53553 , n53554 , n53555 , n53556 , n53557 , n53558 , n53559 , n53560 , 
     n53561 , n53562 , n53563 , n53564 , n53565 , n53566 , n53567 , n53568 , n53569 , n53570 , 
     n53571 , n53572 , n53573 , n53574 , n53575 , n53576 , n53577 , n53578 , n53579 , n53580 , 
     n53581 , n53582 , n53583 , n53584 , n53585 , n53586 , n53587 , n53588 , n53589 , n53590 , 
     n53591 , n53592 , n53593 , n53594 , n53595 , n53596 , n53597 , n53598 , n53599 , n53600 , 
     n53601 , n53602 , n53603 , n53604 , n53605 , n53606 , n53607 , n53608 , n53609 , n53610 , 
     n53611 , n53612 , n53613 , n53614 , n53615 , n53616 , n53617 , n53618 , n53619 , n53620 , 
     n53621 , n53622 , n53623 , n53624 , n53625 , n53626 , n53627 , n53628 , n53629 , n53630 , 
     n53631 , n53632 , n53633 , n53634 , n53635 , n53636 , n53637 , n53638 , n53639 , n53640 , 
     n53641 , n53642 , n53643 , n53644 , n53645 , n53646 , n53647 , n53648 , n53649 , n53650 , 
     n53651 , n53652 , n53653 , n53654 , n53655 , n53656 , n53657 , n53658 , n53659 , n53660 , 
     n53661 , n53662 , n53663 , n53664 , n53665 , n53666 , n53667 , n53668 , n53669 , n53670 , 
     n53671 , n53672 , n53673 , n53674 , n53675 , n53676 , n53677 , n53678 , n53679 , n53680 , 
     n53681 , n53682 , n53683 , n53684 , n53685 , n53686 , n53687 , n53688 , n53689 , n53690 , 
     n53691 , n53692 , n53693 , n53694 , n53695 , n53696 , n53697 , n53698 , n53699 , n53700 , 
     n53701 , n53702 , n53703 , n53704 , n53705 , n53706 , n53707 , n53708 , n53709 , n53710 , 
     n53711 , n53712 , n53713 , n53714 , n53715 , n53716 , n53717 , n53718 , n53719 , n53720 , 
     n53721 , n53722 , n53723 , n53724 , n53725 , n53726 , n53727 , n53728 , n53729 , n53730 , 
     n53731 , n53732 , n53733 , n53734 , n53735 , n53736 , n53737 , n53738 , n53739 , n53740 , 
     n53741 , n53742 , n53743 , n53744 , n53745 , n53746 , n53747 , n53748 , n53749 , n53750 , 
     n53751 , n53752 , n53753 , n53754 , n53755 , n53756 , n53757 , n53758 , n53759 , n53760 , 
     n53761 , n53762 , n53763 , n53764 , n53765 , n53766 , n53767 , n53768 , n53769 , n53770 , 
     n53771 , n53772 , n53773 , n53774 , n53775 , n53776 , n53777 , n53778 , n53779 , n53780 , 
     n53781 , n53782 , n53783 , n53784 , n53785 , n53786 , n53787 , n53788 , n53789 , n53790 , 
     n53791 , n53792 , n53793 , n53794 , n53795 , n53796 , n53797 , n53798 , n53799 , n53800 , 
     n53801 , n53802 , n53803 , n53804 , n53805 , n53806 , n53807 , n53808 , n53809 , n53810 , 
     n53811 , n53812 , n53813 , n53814 , n53815 , n53816 , n53817 , n53818 , n53819 , n53820 , 
     n53821 , n53822 , n53823 , n53824 , n53825 , n53826 , n53827 , n53828 , n53829 , n53830 , 
     n53831 , n53832 , n53833 , n53834 , n53835 , n53836 , n53837 , n53838 , n53839 , n53840 , 
     n53841 , n53842 , n53843 , n53844 , n53845 , n53846 , n53847 , n53848 , n53849 , n53850 , 
     n53851 , n53852 , n53853 , n53854 , n53855 , n53856 , n53857 , n53858 , n53859 , n53860 , 
     n53861 , n53862 , n53863 , n53864 , n53865 , n53866 , n53867 , n53868 , n53869 , n53870 , 
     n53871 , n53872 , n53873 , n53874 , n53875 , n53876 , n53877 , n53878 , n53879 , n53880 , 
     n53881 , n53882 , n53883 , n53884 , n53885 , n53886 , n53887 , n53888 , n53889 , n53890 , 
     n53891 , n53892 , n53893 , n53894 , n53895 , n53896 , n53897 , n53898 , n53899 , n53900 , 
     n53901 , n53902 , n53903 , n53904 , n53905 , n53906 , n53907 , n53908 , n53909 , n53910 , 
     n53911 , n53912 , n53913 , n53914 , n53915 , n53916 , n53917 , n53918 , n53919 , n53920 , 
     n53921 , n53922 , n53923 , n53924 , n53925 , n53926 , n53927 , n53928 , n53929 , n53930 , 
     n53931 , n53932 , n53933 , n53934 , n53935 , n53936 , n53937 , n53938 , n53939 , n53940 , 
     n53941 , n53942 , n53943 , n53944 , n53945 , n53946 , n53947 , n53948 , n53949 , n53950 , 
     n53951 , n53952 , n53953 , n53954 , n53955 , n53956 , n53957 , n53958 , n53959 , n53960 , 
     n53961 , n53962 , n53963 , n53964 , n53965 , n53966 , n53967 , n53968 , n53969 , n53970 , 
     n53971 , n53972 , n53973 , n53974 , n53975 , n53976 , n53977 , n53978 , n53979 , n53980 , 
     n53981 , n53982 , n53983 , n53984 , n53985 , n53986 , n53987 , n53988 , n53989 , n53990 , 
     n53991 , n53992 , n53993 , n53994 , n53995 , n53996 , n53997 , n53998 , n53999 , n54000 , 
     n54001 , n54002 , n54003 , n54004 , n54005 , n54006 , n54007 , n54008 , n54009 , n54010 , 
     n54011 , n54012 , n54013 , n54014 , n54015 , n54016 , n54017 , n54018 , n54019 , n54020 , 
     n54021 , n54022 , n54023 , n54024 , n54025 , n54026 , n54027 , n54028 , n54029 , n54030 , 
     n54031 , n54032 , n54033 , n54034 , n54035 , n54036 , n54037 , n54038 , n54039 , n54040 , 
     n54041 , n54042 , n54043 , n54044 , n54045 , n54046 , n54047 , n54048 , n54049 , n54050 , 
     n54051 , n54052 , n54053 , n54054 , n54055 , n54056 , n54057 , n54058 , n54059 , n54060 , 
     n54061 , n54062 , n54063 , n54064 , n54065 , n54066 , n54067 , n54068 , n54069 , n54070 , 
     n54071 , n54072 , n54073 , n54074 , n54075 , n54076 , n54077 , n54078 , n54079 , n54080 , 
     n54081 , n54082 , n54083 , n54084 , n54085 , n54086 , n54087 , n54088 , n54089 , n54090 , 
     n54091 , n54092 , n54093 , n54094 , n54095 , n54096 , n54097 , n54098 , n54099 , n54100 , 
     n54101 , n54102 , n54103 , n54104 , n54105 , n54106 , n54107 , n54108 , n54109 , n54110 , 
     n54111 , n54112 , n54113 , n54114 , n54115 , n54116 , n54117 , n54118 , n54119 , n54120 , 
     n54121 , n54122 , n54123 , n54124 , n54125 , n54126 , n54127 , n54128 , n54129 , n54130 , 
     n54131 , n54132 , n54133 , n54134 , n54135 , n54136 , n54137 , n54138 , n54139 , n54140 , 
     n54141 , n54142 , n54143 , n54144 , n54145 , n54146 , n54147 , n54148 , n54149 , n54150 , 
     n54151 , n54152 , n54153 , n54154 , n54155 , n54156 , n54157 , n54158 , n54159 , n54160 , 
     n54161 , n54162 , n54163 , n54164 , n54165 , n54166 , n54167 , n54168 , n54169 , n54170 , 
     n54171 , n54172 , n54173 , n54174 , n54175 , n54176 , n54177 , n54178 , n54179 , n54180 , 
     n54181 , n54182 , n54183 , n54184 , n54185 , n54186 , n54187 , n54188 , n54189 , n54190 , 
     n54191 , n54192 , n54193 , n54194 , n54195 , n54196 , n54197 , n54198 , n54199 , n54200 , 
     n54201 , n54202 , n54203 , n54204 , n54205 , n54206 , n54207 , n54208 , n54209 , n54210 , 
     n54211 , n54212 , n54213 , n54214 , n54215 , n54216 , n54217 , n54218 , n54219 , n54220 , 
     n54221 , n54222 , n54223 , n54224 , n54225 , n54226 , n54227 , n54228 , n54229 , n54230 , 
     n54231 , n54232 , n54233 , n54234 , n54235 , n54236 , n54237 , n54238 , n54239 , n54240 , 
     n54241 , n54242 , n54243 , n54244 , n54245 , n54246 , n54247 , n54248 , n54249 , n54250 , 
     n54251 , n54252 , n54253 , n54254 , n54255 , n54256 , n54257 , n54258 , n54259 , n54260 , 
     n54261 , n54262 , n54263 , n54264 , n54265 , n54266 , n54267 , n54268 , n54269 , n54270 , 
     n54271 , n54272 , n54273 , n54274 , n54275 , n54276 , n54277 , n54278 , n54279 , n54280 , 
     n54281 , n54282 , n54283 , n54284 , n54285 , n54286 , n54287 , n54288 , n54289 , n54290 , 
     n54291 , n54292 , n54293 , n54294 , n54295 , n54296 , n54297 , n54298 , n54299 , n54300 , 
     n54301 , n54302 , n54303 , n54304 , n54305 , n54306 , n54307 , n54308 , n54309 , n54310 , 
     n54311 , n54312 , n54313 , n54314 , n54315 , n54316 , n54317 , n54318 , n54319 , n54320 , 
     n54321 , n54322 , n54323 , n54324 , n54325 , n54326 , n54327 , n54328 , n54329 , n54330 , 
     n54331 , n54332 , n54333 , n54334 , n54335 , n54336 , n54337 , n54338 , n54339 , n54340 , 
     n54341 , n54342 , n54343 , n54344 , n54345 , n54346 , n54347 , n54348 , n54349 , n54350 , 
     n54351 , n54352 , n54353 , n54354 , n54355 , n54356 , n54357 , n54358 , n54359 , n54360 , 
     n54361 , n54362 , n54363 , n54364 , n54365 , n54366 , n54367 , n54368 , n54369 , n54370 , 
     n54371 , n54372 , n54373 , n54374 , n54375 , n54376 , n54377 , n54378 , n54379 , n54380 , 
     n54381 , n54382 , n54383 , n54384 , n54385 , n54386 , n54387 , n54388 , n54389 , n54390 , 
     n54391 , n54392 , n54393 , n54394 , n54395 , n54396 , n54397 , n54398 , n54399 , n54400 , 
     n54401 , n54402 , n54403 , n54404 , n54405 , n54406 , n54407 , n54408 , n54409 , n54410 , 
     n54411 , n54412 , n54413 , n54414 , n54415 , n54416 , n54417 , n54418 , n54419 , n54420 , 
     n54421 , n54422 , n54423 , n54424 , n54425 , n54426 , n54427 , n54428 , n54429 , n54430 , 
     n54431 , n54432 , n54433 , n54434 , n54435 , n54436 , n54437 , n54438 , n54439 , n54440 , 
     n54441 , n54442 , n54443 , n54444 , n54445 , n54446 , n54447 , n54448 , n54449 , n54450 , 
     n54451 , n54452 , n54453 , n54454 , n54455 , n54456 , n54457 , n54458 , n54459 , n54460 , 
     n54461 , n54462 , n54463 , n54464 , n54465 , n54466 , n54467 , n54468 , n54469 , n54470 , 
     n54471 , n54472 , n54473 , n54474 , n54475 , n54476 , n54477 , n54478 , n54479 , n54480 , 
     n54481 , n54482 , n54483 , n54484 , n54485 , n54486 , n54487 , n54488 , n54489 , n54490 , 
     n54491 , n54492 , n54493 , n54494 , n54495 , n54496 , n54497 , n54498 , n54499 , n54500 , 
     n54501 , n54502 , n54503 , n54504 , n54505 , n54506 , n54507 , n54508 , n54509 , n54510 , 
     n54511 , n54512 , n54513 , n54514 , n54515 , n54516 , n54517 , n54518 , n54519 , n54520 , 
     n54521 , n54522 , n54523 , n54524 , n54525 , n54526 , n54527 , n54528 , n54529 , n54530 , 
     n54531 , n54532 , n54533 , n54534 , n54535 , n54536 , n54537 , n54538 , n54539 , n54540 , 
     n54541 , n54542 , n54543 , n54544 , n54545 , n54546 , n54547 , n54548 , n54549 , n54550 , 
     n54551 , n54552 , n54553 , n54554 , n54555 , n54556 , n54557 , n54558 , n54559 , n54560 , 
     n54561 , n54562 , n54563 , n54564 , n54565 , n54566 , n54567 , n54568 , n54569 , n54570 , 
     n54571 , n54572 , n54573 , n54574 , n54575 , n54576 , n54577 , n54578 , n54579 , n54580 , 
     n54581 , n54582 , n54583 , n54584 , n54585 , n54586 , n54587 , n54588 , n54589 , n54590 , 
     n54591 , n54592 , n54593 , n54594 , n54595 , n54596 , n54597 , n54598 , n54599 , n54600 , 
     n54601 , n54602 , n54603 , n54604 , n54605 , n54606 , n54607 , n54608 , n54609 , n54610 , 
     n54611 , n54612 , n54613 , n54614 , n54615 , n54616 , n54617 , n54618 , n54619 , n54620 , 
     n54621 , n54622 , n54623 , n54624 , n54625 , n54626 , n54627 , n54628 , n54629 , n54630 , 
     n54631 , n54632 , n54633 , n54634 , n54635 , n54636 , n54637 , n54638 , n54639 , n54640 , 
     n54641 , n54642 , n54643 , n54644 , n54645 , n54646 , n54647 , n54648 , n54649 , n54650 , 
     n54651 , n54652 , n54653 , n54654 , n54655 , n54656 , n54657 , n54658 , n54659 , n54660 , 
     n54661 , n54662 , n54663 , n54664 , n54665 , n54666 , n54667 , n54668 , n54669 , n54670 , 
     n54671 , n54672 , n54673 , n54674 , n54675 , n54676 , n54677 , n54678 , n54679 , n54680 , 
     n54681 , n54682 , n54683 , n54684 , n54685 , n54686 , n54687 , n54688 , n54689 , n54690 , 
     n54691 , n54692 , n54693 , n54694 , n54695 , n54696 , n54697 , n54698 , n54699 , n54700 , 
     n54701 , n54702 , n54703 , n54704 , n54705 , n54706 , n54707 , n54708 , n54709 , n54710 , 
     n54711 , n54712 , n54713 , n54714 , n54715 , n54716 , n54717 , n54718 , n54719 , n54720 , 
     n54721 , n54722 , n54723 , n54724 , n54725 , n54726 , n54727 , n54728 , n54729 , n54730 , 
     n54731 , n54732 , n54733 , n54734 , n54735 , n54736 , n54737 , n54738 , n54739 , n54740 , 
     n54741 , n54742 , n54743 , n54744 , n54745 , n54746 , n54747 , n54748 , n54749 , n54750 , 
     n54751 , n54752 , n54753 , n54754 , n54755 , n54756 , n54757 , n54758 , n54759 , n54760 , 
     n54761 , n54762 , n54763 , n54764 , n54765 , n54766 , n54767 , n54768 , n54769 , n54770 , 
     n54771 , n54772 , n54773 , n54774 , n54775 , n54776 , n54777 , n54778 , n54779 , n54780 , 
     n54781 , n54782 , n54783 , n54784 , n54785 , n54786 , n54787 , n54788 , n54789 , n54790 , 
     n54791 , n54792 , n54793 , n54794 , n54795 , n54796 , n54797 , n54798 , n54799 , n54800 , 
     n54801 , n54802 , n54803 , n54804 , n54805 , n54806 , n54807 , n54808 , n54809 , n54810 , 
     n54811 , n54812 , n54813 , n54814 , n54815 , n54816 , n54817 , n54818 , n54819 , n54820 , 
     n54821 , n54822 , n54823 , n54824 , n54825 , n54826 , n54827 , n54828 , n54829 , n54830 , 
     n54831 , n54832 , n54833 , n54834 , n54835 , n54836 , n54837 , n54838 , n54839 , n54840 , 
     n54841 , n54842 , n54843 , n54844 , n54845 , n54846 , n54847 , n54848 , n54849 , n54850 , 
     n54851 , n54852 , n54853 , n54854 , n54855 , n54856 , n54857 , n54858 , n54859 , n54860 , 
     n54861 , n54862 , n54863 , n54864 , n54865 , n54866 , n54867 , n54868 , n54869 , n54870 , 
     n54871 , n54872 , n54873 , n54874 , n54875 , n54876 , n54877 , n54878 , n54879 , n54880 , 
     n54881 , n54882 , n54883 , n54884 , n54885 , n54886 , n54887 , n54888 , n54889 , n54890 , 
     n54891 , n54892 , n54893 , n54894 , n54895 , n54896 , n54897 , n54898 , n54899 , n54900 , 
     n54901 , n54902 , n54903 , n54904 , n54905 , n54906 , n54907 , n54908 , n54909 , n54910 , 
     n54911 , n54912 , n54913 , n54914 , n54915 , n54916 , n54917 , n54918 , n54919 , n54920 , 
     n54921 , n54922 , n54923 , n54924 , n54925 , n54926 , n54927 , n54928 , n54929 , n54930 , 
     n54931 , n54932 , n54933 , n54934 , n54935 , n54936 , n54937 , n54938 , n54939 , n54940 , 
     n54941 , n54942 , n54943 , n54944 , n54945 , n54946 , n54947 , n54948 , n54949 , n54950 , 
     n54951 , n54952 , n54953 , n54954 , n54955 , n54956 , n54957 , n54958 , n54959 , n54960 , 
     n54961 , n54962 , n54963 , n54964 , n54965 , n54966 , n54967 , n54968 , n54969 , n54970 , 
     n54971 , n54972 , n54973 , n54974 , n54975 , n54976 , n54977 , n54978 , n54979 , n54980 , 
     n54981 , n54982 , n54983 , n54984 , n54985 , n54986 , n54987 , n54988 , n54989 , n54990 , 
     n54991 , n54992 , n54993 , n54994 , n54995 , n54996 , n54997 , n54998 , n54999 , n55000 , 
     n55001 , n55002 , n55003 , n55004 , n55005 , n55006 , n55007 , n55008 , n55009 , n55010 , 
     n55011 , n55012 , n55013 , n55014 , n55015 , n55016 , n55017 , n55018 , n55019 , n55020 , 
     n55021 , n55022 , n55023 , n55024 , n55025 , n55026 , n55027 , n55028 , n55029 , n55030 , 
     n55031 , n55032 , n55033 , n55034 , n55035 , n55036 , n55037 , n55038 , n55039 , n55040 , 
     n55041 , n55042 , n55043 , n55044 , n55045 , n55046 , n55047 , n55048 , n55049 , n55050 , 
     n55051 , n55052 , n55053 , n55054 , n55055 , n55056 , n55057 , n55058 , n55059 , n55060 , 
     n55061 , n55062 , n55063 , n55064 , n55065 , n55066 , n55067 , n55068 , n55069 , n55070 , 
     n55071 , n55072 , n55073 , n55074 , n55075 , n55076 , n55077 , n55078 , n55079 , n55080 , 
     n55081 , n55082 , n55083 , n55084 , n55085 , n55086 , n55087 , n55088 , n55089 , n55090 , 
     n55091 , n55092 , n55093 , n55094 , n55095 , n55096 , n55097 , n55098 , n55099 , n55100 , 
     n55101 , n55102 , n55103 , n55104 , n55105 , n55106 , n55107 , n55108 , n55109 , n55110 , 
     n55111 , n55112 , n55113 , n55114 , n55115 , n55116 , n55117 , n55118 , n55119 , n55120 , 
     n55121 , n55122 , n55123 , n55124 , n55125 , n55126 , n55127 , n55128 , n55129 , n55130 , 
     n55131 , n55132 , n55133 , n55134 , n55135 , n55136 , n55137 , n55138 , n55139 , n55140 , 
     n55141 , n55142 , n55143 , n55144 , n55145 , n55146 , n55147 , n55148 , n55149 , n55150 , 
     n55151 , n55152 , n55153 , n55154 , n55155 , n55156 , n55157 , n55158 , n55159 , n55160 , 
     n55161 , n55162 , n55163 , n55164 , n55165 , n55166 , n55167 , n55168 , n55169 , n55170 , 
     n55171 , n55172 , n55173 , n55174 , n55175 , n55176 , n55177 , n55178 , n55179 , n55180 , 
     n55181 , n55182 , n55183 , n55184 , n55185 , n55186 , n55187 , n55188 , n55189 , n55190 , 
     n55191 , n55192 , n55193 , n55194 , n55195 , n55196 , n55197 , n55198 , n55199 , n55200 , 
     n55201 , n55202 , n55203 , n55204 , n55205 , n55206 , n55207 , n55208 , n55209 , n55210 , 
     n55211 , n55212 , n55213 , n55214 , n55215 , n55216 , n55217 , n55218 , n55219 , n55220 , 
     n55221 , n55222 , n55223 , n55224 , n55225 , n55226 , n55227 , n55228 , n55229 , n55230 , 
     n55231 , n55232 , n55233 , n55234 , n55235 , n55236 , n55237 , n55238 , n55239 , n55240 , 
     n55241 , n55242 , n55243 , n55244 , n55245 , n55246 , n55247 , n55248 , n55249 , n55250 , 
     n55251 , n55252 , n55253 , n55254 , n55255 , n55256 , n55257 , n55258 , n55259 , n55260 , 
     n55261 , n55262 , n55263 , n55264 , n55265 , n55266 , n55267 , n55268 , n55269 , n55270 , 
     n55271 , n55272 , n55273 , n55274 , n55275 , n55276 , n55277 , n55278 , n55279 , n55280 , 
     n55281 , n55282 , n55283 , n55284 , n55285 , n55286 , n55287 , n55288 , n55289 , n55290 , 
     n55291 , n55292 , n55293 , n55294 , n55295 , n55296 , n55297 , n55298 , n55299 , n55300 , 
     n55301 , n55302 , n55303 , n55304 , n55305 , n55306 , n55307 , n55308 , n55309 , n55310 , 
     n55311 , n55312 , n55313 , n55314 , n55315 , n55316 , n55317 , n55318 , n55319 , n55320 , 
     n55321 , n55322 , n55323 , n55324 , n55325 , n55326 , n55327 , n55328 , n55329 , n55330 , 
     n55331 , n55332 , n55333 , n55334 , n55335 , n55336 , n55337 , n55338 , n55339 , n55340 , 
     n55341 , n55342 , n55343 , n55344 , n55345 , n55346 , n55347 , n55348 , n55349 , n55350 , 
     n55351 , n55352 , n55353 , n55354 , n55355 , n55356 , n55357 , n55358 , n55359 , n55360 , 
     n55361 , n55362 , n55363 , n55364 , n55365 , n55366 , n55367 , n55368 , n55369 , n55370 , 
     n55371 , n55372 , n55373 , n55374 , n55375 , n55376 , n55377 , n55378 , n55379 , n55380 , 
     n55381 , n55382 , n55383 , n55384 , n55385 , n55386 , n55387 , n55388 , n55389 , n55390 , 
     n55391 , n55392 , n55393 , n55394 , n55395 , n55396 , n55397 , n55398 , n55399 , n55400 , 
     n55401 , n55402 , n55403 , n55404 , n55405 , n55406 , n55407 , n55408 , n55409 , n55410 , 
     n55411 , n55412 , n55413 , n55414 , n55415 , n55416 , n55417 , n55418 , n55419 , n55420 , 
     n55421 , n55422 , n55423 , n55424 , n55425 , n55426 , n55427 , n55428 , n55429 , n55430 , 
     n55431 , n55432 , n55433 , n55434 , n55435 , n55436 , n55437 , n55438 , n55439 , n55440 , 
     n55441 , n55442 , n55443 , n55444 , n55445 , n55446 , n55447 , n55448 , n55449 , n55450 , 
     n55451 , n55452 , n55453 , n55454 , n55455 , n55456 , n55457 , n55458 , n55459 , n55460 , 
     n55461 , n55462 , n55463 , n55464 , n55465 , n55466 , n55467 , n55468 , n55469 , n55470 , 
     n55471 , n55472 , n55473 , n55474 , n55475 , n55476 , n55477 , n55478 , n55479 , n55480 , 
     n55481 , n55482 , n55483 , n55484 , n55485 , n55486 , n55487 , n55488 , n55489 , n55490 , 
     n55491 , n55492 , n55493 , n55494 , n55495 , n55496 , n55497 , n55498 , n55499 , n55500 , 
     n55501 , n55502 , n55503 , n55504 , n55505 , n55506 , n55507 , n55508 , n55509 , n55510 , 
     n55511 , n55512 , n55513 , n55514 , n55515 , n55516 , n55517 , n55518 , n55519 , n55520 , 
     n55521 , n55522 , n55523 , n55524 , n55525 , n55526 , n55527 , n55528 , n55529 , n55530 , 
     n55531 , n55532 , n55533 , n55534 , n55535 , n55536 , n55537 , n55538 , n55539 , n55540 , 
     n55541 , n55542 , n55543 , n55544 , n55545 , n55546 , n55547 , n55548 , n55549 , n55550 , 
     n55551 , n55552 , n55553 , n55554 , n55555 , n55556 , n55557 , n55558 , n55559 , n55560 , 
     n55561 , n55562 , n55563 , n55564 , n55565 , n55566 , n55567 , n55568 , n55569 , n55570 , 
     n55571 , n55572 , n55573 , n55574 , n55575 , n55576 , n55577 , n55578 , n55579 , n55580 , 
     n55581 , n55582 , n55583 , n55584 , n55585 , n55586 , n55587 , n55588 , n55589 , n55590 , 
     n55591 , n55592 , n55593 , n55594 , n55595 , n55596 , n55597 , n55598 , n55599 , n55600 , 
     n55601 , n55602 , n55603 , n55604 , n55605 , n55606 , n55607 , n55608 , n55609 , n55610 , 
     n55611 , n55612 , n55613 , n55614 , n55615 , n55616 , n55617 , n55618 , n55619 , n55620 , 
     n55621 , n55622 , n55623 , n55624 , n55625 , n55626 , n55627 , n55628 , n55629 , n55630 , 
     n55631 , n55632 , n55633 , n55634 , n55635 , n55636 , n55637 , n55638 , n55639 , n55640 , 
     n55641 , n55642 , n55643 , n55644 , n55645 , n55646 , n55647 , n55648 , n55649 , n55650 , 
     n55651 , n55652 , n55653 , n55654 , n55655 , n55656 , n55657 , n55658 , n55659 , n55660 , 
     n55661 , n55662 , n55663 , n55664 , n55665 , n55666 , n55667 , n55668 , n55669 , n55670 , 
     n55671 , n55672 , n55673 , n55674 , n55675 , n55676 , n55677 , n55678 , n55679 , n55680 , 
     n55681 , n55682 , n55683 , n55684 , n55685 , n55686 , n55687 , n55688 , n55689 , n55690 , 
     n55691 , n55692 , n55693 , n55694 , n55695 , n55696 , n55697 , n55698 , n55699 , n55700 , 
     n55701 , n55702 , n55703 , n55704 , n55705 , n55706 , n55707 , n55708 , n55709 , n55710 , 
     n55711 , n55712 , n55713 , n55714 , n55715 , n55716 , n55717 , n55718 , n55719 , n55720 , 
     n55721 , n55722 , n55723 , n55724 , n55725 , n55726 , n55727 , n55728 , n55729 , n55730 , 
     n55731 , n55732 , n55733 , n55734 , n55735 , n55736 , n55737 , n55738 , n55739 , n55740 , 
     n55741 , n55742 , n55743 , n55744 , n55745 , n55746 , n55747 , n55748 , n55749 , n55750 , 
     n55751 , n55752 , n55753 , n55754 , n55755 , n55756 , n55757 , n55758 , n55759 , n55760 , 
     n55761 , n55762 , n55763 , n55764 , n55765 , n55766 , n55767 , n55768 , n55769 , n55770 , 
     n55771 , n55772 , n55773 , n55774 , n55775 , n55776 , n55777 , n55778 , n55779 , n55780 , 
     n55781 , n55782 , n55783 , n55784 , n55785 , n55786 , n55787 , n55788 , n55789 , n55790 , 
     n55791 , n55792 , n55793 , n55794 , n55795 , n55796 , n55797 , n55798 , n55799 , n55800 , 
     n55801 , n55802 , n55803 , n55804 , n55805 , n55806 , n55807 , n55808 , n55809 , n55810 , 
     n55811 , n55812 , n55813 , n55814 , n55815 , n55816 , n55817 , n55818 , n55819 , n55820 , 
     n55821 , n55822 , n55823 , n55824 , n55825 , n55826 , n55827 , n55828 , n55829 , n55830 , 
     n55831 , n55832 , n55833 , n55834 , n55835 , n55836 , n55837 , n55838 , n55839 , n55840 , 
     n55841 , n55842 , n55843 , n55844 , n55845 , n55846 , n55847 , n55848 , n55849 , n55850 , 
     n55851 , n55852 , n55853 , n55854 , n55855 , n55856 , n55857 , n55858 , n55859 , n55860 , 
     n55861 , n55862 , n55863 , n55864 , n55865 , n55866 , n55867 , n55868 , n55869 , n55870 , 
     n55871 , n55872 , n55873 , n55874 , n55875 , n55876 , n55877 , n55878 , n55879 , n55880 , 
     n55881 , n55882 , n55883 , n55884 , n55885 , n55886 , n55887 , n55888 , n55889 , n55890 , 
     n55891 , n55892 , n55893 , n55894 , n55895 , n55896 , n55897 , n55898 , n55899 , n55900 , 
     n55901 , n55902 , n55903 , n55904 , n55905 , n55906 , n55907 , n55908 , n55909 , n55910 , 
     n55911 , n55912 , n55913 , n55914 , n55915 , n55916 , n55917 , n55918 , n55919 , n55920 , 
     n55921 , n55922 , n55923 , n55924 , n55925 , n55926 , n55927 , n55928 , n55929 , n55930 , 
     n55931 , n55932 , n55933 , n55934 , n55935 , n55936 , n55937 , n55938 , n55939 , n55940 , 
     n55941 , n55942 , n55943 , n55944 , n55945 , n55946 , n55947 , n55948 , n55949 , n55950 , 
     n55951 , n55952 , n55953 , n55954 , n55955 , n55956 , n55957 , n55958 , n55959 , n55960 , 
     n55961 , n55962 , n55963 , n55964 , n55965 , n55966 , n55967 , n55968 , n55969 , n55970 , 
     n55971 , n55972 , n55973 , n55974 , n55975 , n55976 , n55977 , n55978 , n55979 , n55980 , 
     n55981 , n55982 , n55983 , n55984 , n55985 , n55986 , n55987 , n55988 , n55989 , n55990 , 
     n55991 , n55992 , n55993 , n55994 , n55995 , n55996 , n55997 , n55998 , n55999 , n56000 , 
     n56001 , n56002 , n56003 , n56004 , n56005 , n56006 , n56007 , n56008 , n56009 , n56010 , 
     n56011 , n56012 , n56013 , n56014 , n56015 , n56016 , n56017 , n56018 , n56019 , n56020 , 
     n56021 , n56022 , n56023 , n56024 , n56025 , n56026 , n56027 , n56028 , n56029 , n56030 , 
     n56031 , n56032 , n56033 , n56034 , n56035 , n56036 , n56037 , n56038 , n56039 , n56040 , 
     n56041 , n56042 , n56043 , n56044 , n56045 , n56046 , n56047 , n56048 , n56049 , n56050 , 
     n56051 , n56052 , n56053 , n56054 , n56055 , n56056 , n56057 , n56058 , n56059 , n56060 , 
     n56061 , n56062 , n56063 , n56064 , n56065 , n56066 , n56067 , n56068 , n56069 , n56070 , 
     n56071 , n56072 , n56073 , n56074 , n56075 , n56076 , n56077 , n56078 , n56079 , n56080 , 
     n56081 , n56082 , n56083 , n56084 , n56085 , n56086 , n56087 , n56088 , n56089 , n56090 , 
     n56091 , n56092 , n56093 , n56094 , n56095 , n56096 , n56097 , n56098 , n56099 , n56100 , 
     n56101 , n56102 , n56103 , n56104 , n56105 , n56106 , n56107 , n56108 , n56109 , n56110 , 
     n56111 , n56112 , n56113 , n56114 , n56115 , n56116 , n56117 , n56118 , n56119 , n56120 , 
     n56121 , n56122 , n56123 , n56124 , n56125 , n56126 , n56127 , n56128 , n56129 , n56130 , 
     n56131 , n56132 , n56133 , n56134 , n56135 , n56136 , n56137 , n56138 , n56139 , n56140 , 
     n56141 , n56142 , n56143 , n56144 , n56145 , n56146 , n56147 , n56148 , n56149 , n56150 , 
     n56151 , n56152 , n56153 , n56154 , n56155 , n56156 , n56157 , n56158 , n56159 , n56160 , 
     n56161 , n56162 , n56163 , n56164 , n56165 , n56166 , n56167 , n56168 , n56169 , n56170 , 
     n56171 , n56172 , n56173 , n56174 , n56175 , n56176 , n56177 , n56178 , n56179 , n56180 , 
     n56181 , n56182 , n56183 , n56184 , n56185 , n56186 , n56187 , n56188 , n56189 , n56190 , 
     n56191 , n56192 , n56193 , n56194 , n56195 , n56196 , n56197 , n56198 , n56199 , n56200 , 
     n56201 , n56202 , n56203 , n56204 , n56205 , n56206 , n56207 , n56208 , n56209 , n56210 , 
     n56211 , n56212 , n56213 , n56214 , n56215 , n56216 , n56217 , n56218 , n56219 , n56220 , 
     n56221 , n56222 , n56223 , n56224 , n56225 , n56226 , n56227 , n56228 , n56229 , n56230 , 
     n56231 , n56232 , n56233 , n56234 , n56235 , n56236 , n56237 , n56238 , n56239 , n56240 , 
     n56241 , n56242 , n56243 , n56244 , n56245 , n56246 , n56247 , n56248 , n56249 , n56250 , 
     n56251 , n56252 , n56253 , n56254 , n56255 , n56256 , n56257 , n56258 , n56259 , n56260 , 
     n56261 , n56262 , n56263 , n56264 , n56265 , n56266 , n56267 , n56268 , n56269 , n56270 , 
     n56271 , n56272 , n56273 , n56274 , n56275 , n56276 , n56277 , n56278 , n56279 , n56280 , 
     n56281 , n56282 , n56283 , n56284 , n56285 , n56286 , n56287 , n56288 , n56289 , n56290 , 
     n56291 , n56292 , n56293 , n56294 , n56295 , n56296 , n56297 , n56298 , n56299 , n56300 , 
     n56301 , n56302 , n56303 , n56304 , n56305 , n56306 , n56307 , n56308 , n56309 , n56310 , 
     n56311 , n56312 , n56313 , n56314 , n56315 , n56316 , n56317 , n56318 , n56319 , n56320 , 
     n56321 , n56322 , n56323 , n56324 , n56325 , n56326 , n56327 , n56328 , n56329 , n56330 , 
     n56331 , n56332 , n56333 , n56334 , n56335 , n56336 , n56337 , n56338 , n56339 , n56340 , 
     n56341 , n56342 , n56343 , n56344 , n56345 , n56346 , n56347 , n56348 , n56349 , n56350 , 
     n56351 , n56352 , n56353 , n56354 , n56355 , n56356 , n56357 , n56358 , n56359 , n56360 , 
     n56361 , n56362 , n56363 , n56364 , n56365 , n56366 , n56367 , n56368 , n56369 , n56370 , 
     n56371 , n56372 , n56373 , n56374 , n56375 , n56376 , n56377 , n56378 , n56379 , n56380 , 
     n56381 , n56382 , n56383 , n56384 , n56385 , n56386 , n56387 , n56388 , n56389 , n56390 , 
     n56391 , n56392 , n56393 , n56394 , n56395 , n56396 , n56397 , n56398 , n56399 , n56400 , 
     n56401 , n56402 , n56403 , n56404 , n56405 , n56406 , n56407 , n56408 , n56409 , n56410 , 
     n56411 , n56412 , n56413 , n56414 , n56415 , n56416 , n56417 , n56418 , n56419 , n56420 , 
     n56421 , n56422 , n56423 , n56424 , n56425 , n56426 , n56427 , n56428 , n56429 , n56430 , 
     n56431 , n56432 , n56433 , n56434 , n56435 , n56436 , n56437 , n56438 , n56439 , n56440 , 
     n56441 , n56442 , n56443 , n56444 , n56445 , n56446 , n56447 , n56448 , n56449 , n56450 , 
     n56451 , n56452 , n56453 , n56454 , n56455 , n56456 , n56457 , n56458 , n56459 , n56460 , 
     n56461 , n56462 , n56463 , n56464 , n56465 , n56466 , n56467 , n56468 , n56469 , n56470 , 
     n56471 , n56472 , n56473 , n56474 , n56475 , n56476 , n56477 , n56478 , n56479 , n56480 , 
     n56481 , n56482 , n56483 , n56484 , n56485 , n56486 , n56487 , n56488 , n56489 , n56490 , 
     n56491 , n56492 , n56493 , n56494 , n56495 , n56496 , n56497 , n56498 , n56499 , n56500 , 
     n56501 , n56502 , n56503 , n56504 , n56505 , n56506 , n56507 , n56508 , n56509 , n56510 , 
     n56511 , n56512 , n56513 , n56514 , n56515 , n56516 , n56517 , n56518 , n56519 , n56520 , 
     n56521 , n56522 , n56523 , n56524 , n56525 , n56526 , n56527 , n56528 , n56529 , n56530 , 
     n56531 , n56532 , n56533 , n56534 , n56535 , n56536 , n56537 , n56538 , n56539 , n56540 , 
     n56541 , n56542 , n56543 , n56544 , n56545 , n56546 , n56547 , n56548 , n56549 , n56550 , 
     n56551 , n56552 , n56553 , n56554 , n56555 , n56556 , n56557 , n56558 , n56559 , n56560 , 
     n56561 , n56562 , n56563 , n56564 , n56565 , n56566 , n56567 , n56568 , n56569 , n56570 , 
     n56571 , n56572 , n56573 , n56574 , n56575 , n56576 , n56577 , n56578 , n56579 , n56580 , 
     n56581 , n56582 , n56583 , n56584 , n56585 , n56586 , n56587 , n56588 , n56589 , n56590 , 
     n56591 , n56592 , n56593 , n56594 , n56595 , n56596 , n56597 , n56598 , n56599 , n56600 , 
     n56601 , n56602 , n56603 , n56604 , n56605 , n56606 , n56607 , n56608 , n56609 , n56610 , 
     n56611 , n56612 , n56613 , n56614 , n56615 , n56616 , n56617 , n56618 , n56619 , n56620 , 
     n56621 , n56622 , n56623 , n56624 , n56625 , n56626 , n56627 , n56628 , n56629 , n56630 , 
     n56631 , n56632 , n56633 , n56634 , n56635 , n56636 , n56637 , n56638 , n56639 , n56640 , 
     n56641 , n56642 , n56643 , n56644 , n56645 , n56646 , n56647 , n56648 , n56649 , n56650 , 
     n56651 , n56652 , n56653 , n56654 , n56655 , n56656 , n56657 , n56658 , n56659 , n56660 , 
     n56661 , n56662 , n56663 , n56664 , n56665 , n56666 , n56667 , n56668 , n56669 , n56670 , 
     n56671 , n56672 , n56673 , n56674 , n56675 , n56676 , n56677 , n56678 , n56679 , n56680 , 
     n56681 , n56682 , n56683 , n56684 , n56685 , n56686 , n56687 , n56688 , n56689 , n56690 , 
     n56691 , n56692 , n56693 , n56694 , n56695 , n56696 , n56697 , n56698 , n56699 , n56700 , 
     n56701 , n56702 , n56703 , n56704 , n56705 , n56706 , n56707 , n56708 , n56709 , n56710 , 
     n56711 , n56712 , n56713 , n56714 , n56715 , n56716 , n56717 , n56718 , n56719 , n56720 , 
     n56721 , n56722 , n56723 , n56724 , n56725 , n56726 , n56727 , n56728 , n56729 , n56730 , 
     n56731 , n56732 , n56733 , n56734 , n56735 , n56736 , n56737 , n56738 , n56739 , n56740 , 
     n56741 , n56742 , n56743 , n56744 , n56745 , n56746 , n56747 , n56748 , n56749 , n56750 , 
     n56751 , n56752 , n56753 , n56754 , n56755 , n56756 , n56757 , n56758 , n56759 , n56760 , 
     n56761 , n56762 , n56763 , n56764 , n56765 , n56766 , n56767 , n56768 , n56769 , n56770 , 
     n56771 , n56772 , n56773 , n56774 , n56775 , n56776 , n56777 , n56778 , n56779 , n56780 , 
     n56781 , n56782 , n56783 , n56784 , n56785 , n56786 , n56787 , n56788 , n56789 , n56790 , 
     n56791 , n56792 , n56793 , n56794 , n56795 , n56796 , n56797 , n56798 , n56799 , n56800 , 
     n56801 , n56802 , n56803 , n56804 , n56805 , n56806 , n56807 , n56808 , n56809 , n56810 , 
     n56811 , n56812 , n56813 , n56814 , n56815 , n56816 , n56817 , n56818 , n56819 , n56820 , 
     n56821 , n56822 , n56823 , n56824 , n56825 , n56826 , n56827 , n56828 , n56829 , n56830 , 
     n56831 , n56832 , n56833 , n56834 , n56835 , n56836 , n56837 , n56838 , n56839 , n56840 , 
     n56841 , n56842 , n56843 , n56844 , n56845 , n56846 , n56847 , n56848 , n56849 , n56850 , 
     n56851 , n56852 , n56853 , n56854 , n56855 , n56856 , n56857 , n56858 , n56859 , n56860 , 
     n56861 , n56862 , n56863 , n56864 , n56865 , n56866 , n56867 , n56868 , n56869 , n56870 , 
     n56871 , n56872 , n56873 , n56874 , n56875 , n56876 , n56877 , n56878 , n56879 , n56880 , 
     n56881 , n56882 , n56883 , n56884 , n56885 , n56886 , n56887 , n56888 , n56889 , n56890 , 
     n56891 , n56892 , n56893 , n56894 , n56895 , n56896 , n56897 , n56898 , n56899 , n56900 , 
     n56901 , n56902 , n56903 , n56904 , n56905 , n56906 , n56907 , n56908 , n56909 , n56910 , 
     n56911 , n56912 , n56913 , n56914 , n56915 , n56916 , n56917 , n56918 , n56919 , n56920 , 
     n56921 , n56922 , n56923 , n56924 , n56925 , n56926 , n56927 , n56928 , n56929 , n56930 , 
     n56931 , n56932 , n56933 , n56934 , n56935 , n56936 , n56937 , n56938 , n56939 , n56940 , 
     n56941 , n56942 , n56943 , n56944 , n56945 , n56946 , n56947 , n56948 , n56949 , n56950 , 
     n56951 , n56952 , n56953 , n56954 , n56955 , n56956 , n56957 , n56958 , n56959 , n56960 , 
     n56961 , n56962 , n56963 , n56964 , n56965 , n56966 , n56967 , n56968 , n56969 , n56970 , 
     n56971 , n56972 , n56973 , n56974 , n56975 , n56976 , n56977 , n56978 , n56979 , n56980 , 
     n56981 , n56982 , n56983 , n56984 , n56985 , n56986 , n56987 , n56988 , n56989 , n56990 , 
     n56991 , n56992 , n56993 , n56994 , n56995 , n56996 , n56997 , n56998 , n56999 , n57000 , 
     n57001 , n57002 , n57003 , n57004 , n57005 , n57006 , n57007 , n57008 , n57009 , n57010 , 
     n57011 , n57012 , n57013 , n57014 , n57015 , n57016 , n57017 , n57018 , n57019 , n57020 , 
     n57021 , n57022 , n57023 , n57024 , n57025 , n57026 , n57027 , n57028 , n57029 , n57030 , 
     n57031 , n57032 , n57033 , n57034 , n57035 , n57036 , n57037 , n57038 , n57039 , n57040 , 
     n57041 , n57042 , n57043 , n57044 , n57045 , n57046 , n57047 , n57048 , n57049 , n57050 , 
     n57051 , n57052 , n57053 , n57054 , n57055 , n57056 , n57057 , n57058 , n57059 , n57060 , 
     n57061 , n57062 , n57063 , n57064 , n57065 , n57066 , n57067 , n57068 , n57069 , n57070 , 
     n57071 , n57072 , n57073 , n57074 , n57075 , n57076 , n57077 , n57078 , n57079 , n57080 , 
     n57081 , n57082 , n57083 , n57084 , n57085 , n57086 , n57087 , n57088 , n57089 , n57090 , 
     n57091 , n57092 , n57093 , n57094 , n57095 , n57096 , n57097 , n57098 , n57099 , n57100 , 
     n57101 , n57102 , n57103 , n57104 , n57105 , n57106 , n57107 , n57108 , n57109 , n57110 , 
     n57111 , n57112 , n57113 , n57114 , n57115 , n57116 , n57117 , n57118 , n57119 , n57120 , 
     n57121 , n57122 , n57123 , n57124 , n57125 , n57126 , n57127 , n57128 , n57129 , n57130 , 
     n57131 , n57132 , n57133 , n57134 , n57135 , n57136 , n57137 , n57138 , n57139 , n57140 , 
     n57141 , n57142 , n57143 , n57144 , n57145 , n57146 , n57147 , n57148 , n57149 , n57150 , 
     n57151 , n57152 , n57153 , n57154 , n57155 , n57156 , n57157 , n57158 , n57159 , n57160 , 
     n57161 , n57162 , n57163 , n57164 , n57165 , n57166 , n57167 , n57168 , n57169 , n57170 , 
     n57171 , n57172 , n57173 , n57174 , n57175 , n57176 , n57177 , n57178 , n57179 , n57180 , 
     n57181 , n57182 , n57183 , n57184 , n57185 , n57186 , n57187 , n57188 , n57189 , n57190 , 
     n57191 , n57192 , n57193 , n57194 , n57195 , n57196 , n57197 , n57198 , n57199 , n57200 , 
     n57201 , n57202 , n57203 , n57204 , n57205 , n57206 , n57207 , n57208 , n57209 , n57210 , 
     n57211 , n57212 , n57213 , n57214 , n57215 , n57216 , n57217 , n57218 , n57219 , n57220 , 
     n57221 , n57222 , n57223 , n57224 , n57225 , n57226 , n57227 , n57228 , n57229 , n57230 , 
     n57231 , n57232 , n57233 , n57234 , n57235 , n57236 , n57237 , n57238 , n57239 , n57240 , 
     n57241 , n57242 , n57243 , n57244 , n57245 , n57246 , n57247 , n57248 , n57249 , n57250 , 
     n57251 , n57252 , n57253 , n57254 , n57255 , n57256 , n57257 , n57258 , n57259 , n57260 , 
     n57261 , n57262 , n57263 , n57264 , n57265 , n57266 , n57267 , n57268 , n57269 , n57270 , 
     n57271 , n57272 , n57273 , n57274 , n57275 , n57276 , n57277 , n57278 , n57279 , n57280 , 
     n57281 , n57282 , n57283 , n57284 , n57285 , n57286 , n57287 , n57288 , n57289 , n57290 , 
     n57291 , n57292 , n57293 , n57294 , n57295 , n57296 , n57297 , n57298 , n57299 , n57300 , 
     n57301 , n57302 , n57303 , n57304 , n57305 , n57306 , n57307 , n57308 , n57309 , n57310 , 
     n57311 , n57312 , n57313 , n57314 , n57315 , n57316 , n57317 , n57318 , n57319 , n57320 , 
     n57321 , n57322 , n57323 , n57324 , n57325 , n57326 , n57327 , n57328 , n57329 , n57330 , 
     n57331 , n57332 , n57333 , n57334 , n57335 , n57336 , n57337 , n57338 , n57339 , n57340 , 
     n57341 , n57342 , n57343 , n57344 , n57345 , n57346 , n57347 , n57348 , n57349 , n57350 , 
     n57351 , n57352 , n57353 , n57354 , n57355 , n57356 , n57357 , n57358 , n57359 , n57360 , 
     n57361 , n57362 , n57363 , n57364 , n57365 , n57366 , n57367 , n57368 , n57369 , n57370 , 
     n57371 , n57372 , n57373 , n57374 , n57375 , n57376 , n57377 , n57378 , n57379 , n57380 , 
     n57381 , n57382 , n57383 , n57384 , n57385 , n57386 , n57387 , n57388 , n57389 , n57390 , 
     n57391 , n57392 , n57393 , n57394 , n57395 , n57396 , n57397 , n57398 , n57399 , n57400 , 
     n57401 , n57402 , n57403 , n57404 , n57405 , n57406 , n57407 , n57408 , n57409 , n57410 , 
     n57411 , n57412 , n57413 , n57414 , n57415 , n57416 , n57417 , n57418 , n57419 , n57420 , 
     n57421 , n57422 , n57423 , n57424 , n57425 , n57426 , n57427 , n57428 , n57429 , n57430 , 
     n57431 , n57432 , n57433 , n57434 , n57435 , n57436 , n57437 , n57438 , n57439 , n57440 , 
     n57441 , n57442 , n57443 , n57444 , n57445 , n57446 , n57447 , n57448 , n57449 , n57450 , 
     n57451 , n57452 , n57453 , n57454 , n57455 , n57456 , n57457 , n57458 , n57459 , n57460 , 
     n57461 , n57462 , n57463 , n57464 , n57465 , n57466 , n57467 , n57468 , n57469 , n57470 , 
     n57471 , n57472 , n57473 , n57474 , n57475 , n57476 , n57477 , n57478 , n57479 , n57480 , 
     n57481 , n57482 , n57483 , n57484 , n57485 , n57486 , n57487 , n57488 , n57489 , n57490 , 
     n57491 , n57492 , n57493 , n57494 , n57495 , n57496 , n57497 , n57498 , n57499 , n57500 , 
     n57501 , n57502 , n57503 , n57504 , n57505 , n57506 , n57507 , n57508 , n57509 , n57510 , 
     n57511 , n57512 , n57513 , n57514 , n57515 , n57516 , n57517 , n57518 , n57519 , n57520 , 
     n57521 , n57522 , n57523 , n57524 , n57525 , n57526 , n57527 , n57528 , n57529 , n57530 , 
     n57531 , n57532 , n57533 , n57534 , n57535 , n57536 , n57537 , n57538 , n57539 , n57540 , 
     n57541 , n57542 , n57543 , n57544 , n57545 , n57546 , n57547 , n57548 , n57549 , n57550 , 
     n57551 , n57552 , n57553 , n57554 , n57555 , n57556 , n57557 , n57558 ;
buf ( RI15b3e9d0_1 , n0 );
buf ( RI15b51198_632 , n4 );
buf ( RI15b51210_633 , n5 );
buf ( RI15b51120_631 , n2 );
buf ( RI15b51288_634 , n3 );
buf ( RI15b54690_745 , n150 );
buf ( RI15b56760_815 , n187 );
buf ( RI15b567d8_816 , n186 );
buf ( RI15b566e8_814 , n188 );
buf ( RI15b570c0_835 , n168 );
buf ( RI15b57138_836 , n167 );
buf ( RI15b571b0_837 , n166 );
buf ( RI15b57228_838 , n165 );
buf ( RI15b572a0_839 , n164 );
buf ( RI15b57318_840 , n163 );
buf ( RI15b57390_841 , n162 );
buf ( RI15b57408_842 , n161 );
buf ( RI15b56850_817 , n1 );
buf ( RI15b568c8_818 , n185 );
buf ( RI15b56940_819 , n184 );
buf ( RI15b569b8_820 , n183 );
buf ( RI15b56a30_821 , n182 );
buf ( RI15b56aa8_822 , n181 );
buf ( RI15b56b20_823 , n180 );
buf ( RI15b56b98_824 , n179 );
buf ( RI15b56c10_825 , n178 );
buf ( RI15b56c88_826 , n177 );
buf ( RI15b56d00_827 , n176 );
buf ( RI15b56d78_828 , n175 );
buf ( RI15b56df0_829 , n174 );
buf ( RI15b56e68_830 , n173 );
buf ( RI15b56ee0_831 , n172 );
buf ( RI15b56f58_832 , n171 );
buf ( RI15b56fd0_833 , n170 );
buf ( RI15b57048_834 , n169 );
buf ( RI15b57480_843 , n160 );
buf ( RI15b574f8_844 , n159 );
buf ( RI15b57570_845 , n158 );
buf ( RI15b4d340_499 , n60 );
buf ( RI15b50e50_625 , n15 );
buf ( RI15b50ec8_626 , n13 );
buf ( RI15b50f40_627 , n11 );
buf ( RI15b50fb8_628 , n9 );
buf ( RI15b51030_629 , n7 );
buf ( RI15b4dac0_515 , n58 );
buf ( RI15b4e9c0_547 , n54 );
buf ( RI15b4ed80_555 , n53 );
buf ( RI15b4fc80_587 , n49 );
buf ( RI15b4e600_539 , n55 );
buf ( RI15b4c800_475 , n63 );
buf ( RI15b4d700_507 , n59 );
buf ( RI15b4c440_467 , n64 );
buf ( RI15b4cbc0_483 , n62 );
buf ( RI15b4cf80_491 , n61 );
buf ( RI15b4f140_563 , n52 );
buf ( RI15b4f8c0_579 , n50 );
buf ( RI15b4e240_531 , n56 );
buf ( RI15b4f500_571 , n51 );
buf ( RI15b4de80_523 , n57 );
buf ( RI15b4d3b8_500 , n76 );
buf ( RI15b4db38_516 , n74 );
buf ( RI15b4ea38_548 , n70 );
buf ( RI15b4edf8_556 , n69 );
buf ( RI15b4fcf8_588 , n65 );
buf ( RI15b4e678_540 , n71 );
buf ( RI15b4c878_476 , n79 );
buf ( RI15b4d778_508 , n75 );
buf ( RI15b4cc38_484 , n78 );
buf ( RI15b4c4b8_468 , n80 );
buf ( RI15b4cff8_492 , n77 );
buf ( RI15b4f1b8_564 , n68 );
buf ( RI15b4f938_580 , n66 );
buf ( RI15b4e2b8_532 , n72 );
buf ( RI15b4f578_572 , n67 );
buf ( RI15b4def8_524 , n73 );
buf ( RI15b4d598_504 , n140 );
buf ( RI15b4dd18_520 , n138 );
buf ( RI15b4ec18_552 , n134 );
buf ( RI15b4efd8_560 , n133 );
buf ( RI15b4fed8_592 , n129 );
buf ( RI15b4e858_544 , n135 );
buf ( RI15b4ca58_480 , n143 );
buf ( RI15b4d958_512 , n139 );
buf ( RI15b4ce18_488 , n142 );
buf ( RI15b4c698_472 , n144 );
buf ( RI15b4d1d8_496 , n141 );
buf ( RI15b4f398_568 , n132 );
buf ( RI15b4fb18_584 , n130 );
buf ( RI15b4e498_536 , n136 );
buf ( RI15b4f758_576 , n131 );
buf ( RI15b4e0d8_528 , n137 );
buf ( RI15b4d4a8_502 , n108 );
buf ( RI15b4dc28_518 , n106 );
buf ( RI15b4eb28_550 , n102 );
buf ( RI15b4eee8_558 , n101 );
buf ( RI15b4fde8_590 , n97 );
buf ( RI15b4c968_478 , n111 );
buf ( RI15b4d868_510 , n107 );
buf ( RI15b4cd28_486 , n110 );
buf ( RI15b4c5a8_470 , n112 );
buf ( RI15b4d0e8_494 , n109 );
buf ( RI15b4e768_542 , n103 );
buf ( RI15b4f2a8_566 , n100 );
buf ( RI15b4fa28_582 , n98 );
buf ( RI15b4e3a8_534 , n104 );
buf ( RI15b4f668_574 , n99 );
buf ( RI15b4dfe8_526 , n105 );
buf ( RI15b4d430_501 , n92 );
buf ( RI15b4dbb0_517 , n90 );
buf ( RI15b4eab0_549 , n86 );
buf ( RI15b4ee70_557 , n85 );
buf ( RI15b4fd70_589 , n81 );
buf ( RI15b4c8f0_477 , n95 );
buf ( RI15b4d7f0_509 , n91 );
buf ( RI15b4d070_493 , n93 );
buf ( RI15b4e6f0_541 , n87 );
buf ( RI15b4c530_469 , n96 );
buf ( RI15b4ccb0_485 , n94 );
buf ( RI15b4f230_565 , n84 );
buf ( RI15b4f9b0_581 , n82 );
buf ( RI15b4e330_533 , n88 );
buf ( RI15b4f5f0_573 , n83 );
buf ( RI15b4df70_525 , n89 );
buf ( RI15b4d520_503 , n124 );
buf ( RI15b4dca0_519 , n122 );
buf ( RI15b4eba0_551 , n118 );
buf ( RI15b4ef60_559 , n117 );
buf ( RI15b4fe60_591 , n113 );
buf ( RI15b4e7e0_543 , n119 );
buf ( RI15b4c9e0_479 , n127 );
buf ( RI15b4d8e0_511 , n123 );
buf ( RI15b4cda0_487 , n126 );
buf ( RI15b4c620_471 , n128 );
buf ( RI15b4d160_495 , n125 );
buf ( RI15b4f320_567 , n116 );
buf ( RI15b4faa0_583 , n114 );
buf ( RI15b4e420_535 , n120 );
buf ( RI15b4f6e0_575 , n115 );
buf ( RI15b4e060_527 , n121 );
buf ( RI15b4c788_474 , n47 );
buf ( RI15b4cf08_490 , n45 );
buf ( RI15b4d688_506 , n43 );
buf ( RI15b4c3c8_466 , n48 );
buf ( RI15b4cb48_482 , n46 );
buf ( RI15b4f0c8_562 , n36 );
buf ( RI15b4e588_538 , n39 );
buf ( RI15b4f848_578 , n34 );
buf ( RI15b4f488_570 , n35 );
buf ( RI15b4de08_522 , n41 );
buf ( RI15b4e1c8_530 , n40 );
buf ( RI15b4d2c8_498 , n44 );
buf ( RI15b4ed08_554 , n37 );
buf ( RI15b4fc08_586 , n33 );
buf ( RI15b4e948_546 , n38 );
buf ( RI15b4da48_514 , n42 );
buf ( RI15b4d250_497 , n28 );
buf ( RI15b4d9d0_513 , n26 );
buf ( RI15b4e8d0_545 , n22 );
buf ( RI15b4ec90_553 , n21 );
buf ( RI15b4fb90_585 , n17 );
buf ( RI15b4e510_537 , n23 );
buf ( RI15b4c710_473 , n31 );
buf ( RI15b4d610_505 , n27 );
buf ( RI15b4cad0_481 , n30 );
buf ( RI15b4c350_465 , n32 );
buf ( RI15b4ce90_489 , n29 );
buf ( RI15b4f050_561 , n20 );
buf ( RI15b4f7d0_577 , n18 );
buf ( RI15b4e150_529 , n24 );
buf ( RI15b4f410_569 , n19 );
buf ( RI15b4dd90_521 , n25 );
buf ( RI15b4c1e8_462 , n10 );
buf ( RI15b4c0f8_460 , n14 );
buf ( RI15b4c170_461 , n12 );
buf ( RI15b4c260_463 , n8 );
buf ( RI15b4c2d8_464 , n6 );
buf ( RI15b667c8_1362 , n148 );
buf ( RI15b66840_1363 , n149 );
buf ( RI15b557e8_782 , n157 );
buf ( RI15b55860_783 , n156 );
buf ( RI15b558d8_784 , n155 );
buf ( RI15b56670_813 , n154 );
buf ( RI15b547f8_748 , n146 );
buf ( RI15b54870_749 , n147 );
buf ( RI15b54780_747 , n145 );
buf ( RI15b55950_785 , n151 );
buf ( RI15b57750_849 , n16 );
buf ( RI15b57660_847 , n153 );
buf ( RI15b576d8_848 , n152 );
buf ( RI15b3ea48_2 , n189 );
buf ( RI15b5c4a8_1014 , n207 );
buf ( RI15b5c520_1015 , n206 );
buf ( RI15b5c598_1016 , n205 );
buf ( RI15b5c430_1013 , n208 );
buf ( RI15b5c610_1017 , n204 );
buf ( RI15b5c688_1018 , n203 );
buf ( RI15b5c700_1019 , n202 );
buf ( RI15b5c778_1020 , n201 );
buf ( RI15b5d2b8_1044 , n199 );
buf ( RI15b5d330_1045 , n197 );
buf ( RI15b5d420_1047 , n193 );
buf ( RI15b5d3a8_1046 , n195 );
buf ( RI15b5b440_979 , n214 );
buf ( RI15b5b080_971 , n215 );
buf ( RI15b5a900_955 , n217 );
buf ( RI15b5acc0_963 , n216 );
buf ( RI15b5b800_987 , n213 );
buf ( RI15b5bbc0_995 , n212 );
buf ( RI15b5bf80_1003 , n211 );
buf ( RI15b5c340_1011 , n210 );
buf ( RI15b59a00_923 , n221 );
buf ( RI15b59dc0_931 , n220 );
buf ( RI15b5a180_939 , n219 );
buf ( RI15b5a540_947 , n218 );
buf ( RI15b59640_915 , n222 );
buf ( RI15b59280_907 , n223 );
buf ( RI15b58b00_891 , n225 );
buf ( RI15b58ec0_899 , n224 );
buf ( RI15b5b008_970 , n231 );
buf ( RI15b5b3c8_978 , n230 );
buf ( RI15b5a4c8_946 , n234 );
buf ( RI15b5a108_938 , n235 );
buf ( RI15b5a888_954 , n233 );
buf ( RI15b5ac48_962 , n232 );
buf ( RI15b59988_922 , n237 );
buf ( RI15b59d48_930 , n236 );
buf ( RI15b5bf08_1002 , n227 );
buf ( RI15b5c2c8_1010 , n226 );
buf ( RI15b595c8_914 , n238 );
buf ( RI15b59208_906 , n239 );
buf ( RI15b58a88_890 , n241 );
buf ( RI15b58e48_898 , n240 );
buf ( RI15b5b788_986 , n229 );
buf ( RI15b5bb48_994 , n228 );
buf ( RI15b5be18_1000 , n259 );
buf ( RI15b5c1d8_1008 , n258 );
buf ( RI15b59118_904 , n271 );
buf ( RI15b594d8_912 , n270 );
buf ( RI15b5a798_952 , n265 );
buf ( RI15b5ab58_960 , n264 );
buf ( RI15b59898_920 , n269 );
buf ( RI15b59c58_928 , n268 );
buf ( RI15b5b2d8_976 , n262 );
buf ( RI15b5af18_968 , n263 );
buf ( RI15b5a3d8_944 , n266 );
buf ( RI15b5a018_936 , n267 );
buf ( RI15b58998_888 , n273 );
buf ( RI15b58d58_896 , n272 );
buf ( RI15b5b698_984 , n261 );
buf ( RI15b5ba58_992 , n260 );
buf ( RI15b59820_919 , n285 );
buf ( RI15b59be0_927 , n284 );
buf ( RI15b5b260_975 , n278 );
buf ( RI15b5aea0_967 , n279 );
buf ( RI15b5a360_943 , n282 );
buf ( RI15b59fa0_935 , n283 );
buf ( RI15b5a720_951 , n281 );
buf ( RI15b5aae0_959 , n280 );
buf ( RI15b58920_887 , n289 );
buf ( RI15b58ce0_895 , n288 );
buf ( RI15b5c160_1007 , n274 );
buf ( RI15b5bda0_999 , n275 );
buf ( RI15b5b620_983 , n277 );
buf ( RI15b5b9e0_991 , n276 );
buf ( RI15b59460_911 , n286 );
buf ( RI15b590a0_903 , n287 );
buf ( RI15b5ae28_966 , n295 );
buf ( RI15b5b1e8_974 , n294 );
buf ( RI15b5c0e8_1006 , n290 );
buf ( RI15b5bd28_998 , n291 );
buf ( RI15b5b5a8_982 , n293 );
buf ( RI15b5b968_990 , n292 );
buf ( RI15b593e8_910 , n302 );
buf ( RI15b59028_902 , n303 );
buf ( RI15b5a6a8_950 , n297 );
buf ( RI15b5a2e8_942 , n298 );
buf ( RI15b59f28_934 , n299 );
buf ( RI15b5aa68_958 , n296 );
buf ( RI15b588a8_886 , n305 );
buf ( RI15b58c68_894 , n304 );
buf ( RI15b597a8_918 , n301 );
buf ( RI15b59b68_926 , n300 );
buf ( RI15b5b170_973 , n310 );
buf ( RI15b5adb0_965 , n311 );
buf ( RI15b59370_909 , n318 );
buf ( RI15b58fb0_901 , n319 );
buf ( RI15b5c070_1005 , n306 );
buf ( RI15b5bcb0_997 , n307 );
buf ( RI15b5a270_941 , n314 );
buf ( RI15b59eb0_933 , n315 );
buf ( RI15b5a630_949 , n313 );
buf ( RI15b58830_885 , n321 );
buf ( RI15b58bf0_893 , n320 );
buf ( RI15b5a9f0_957 , n312 );
buf ( RI15b5b530_981 , n309 );
buf ( RI15b59730_917 , n317 );
buf ( RI15b59af0_925 , n316 );
buf ( RI15b5b8f0_989 , n308 );
buf ( RI15b5bff8_1004 , n322 );
buf ( RI15b5bc38_996 , n323 );
buf ( RI15b592f8_908 , n334 );
buf ( RI15b58f38_900 , n335 );
buf ( RI15b5b0f8_972 , n326 );
buf ( RI15b5ad38_964 , n327 );
buf ( RI15b5a1f8_940 , n330 );
buf ( RI15b59e38_932 , n331 );
buf ( RI15b5a5b8_948 , n329 );
buf ( RI15b596b8_916 , n333 );
buf ( RI15b5b4b8_980 , n325 );
buf ( RI15b5a978_956 , n328 );
buf ( RI15b587b8_884 , n337 );
buf ( RI15b59a78_924 , n332 );
buf ( RI15b5b878_988 , n324 );
buf ( RI15b58b78_892 , n336 );
buf ( RI15b5c3b8_1012 , n209 );
buf ( RI15b5c250_1009 , n242 );
buf ( RI15b5be90_1001 , n243 );
buf ( RI15b5b350_977 , n246 );
buf ( RI15b5af90_969 , n247 );
buf ( RI15b5a810_953 , n249 );
buf ( RI15b5abd0_961 , n248 );
buf ( RI15b5b710_985 , n245 );
buf ( RI15b5bad0_993 , n244 );
buf ( RI15b5a450_945 , n250 );
buf ( RI15b5a090_937 , n251 );
buf ( RI15b59550_913 , n254 );
buf ( RI15b59190_905 , n255 );
buf ( RI15b58a10_889 , n257 );
buf ( RI15b58dd0_897 , n256 );
buf ( RI15b59910_921 , n253 );
buf ( RI15b59cd0_929 , n252 );
buf ( RI15b5d498_1048 , n191 );
buf ( RI15b5d588_1050 , n338 );
buf ( RI15b5d6f0_1053 , n339 );
buf ( RI15b5d600_1051 , n340 );
buf ( RI15b5d678_1052 , n341 );
buf ( RI15b58740_883 , n190 );
buf ( RI15b586c8_882 , n192 );
buf ( RI15b58650_881 , n194 );
buf ( RI15b58560_879 , n198 );
buf ( RI15b585d8_880 , n196 );
buf ( RI15b63e10_1273 , n350 );
buf ( RI15b62f10_1241 , n200 );
buf ( RI15b62c40_1235 , n347 );
buf ( RI15b62cb8_1236 , n346 );
buf ( RI15b62d30_1237 , n345 );
buf ( RI15b62da8_1238 , n344 );
buf ( RI15b62e20_1239 , n343 );
buf ( RI15b62e98_1240 , n342 );
buf ( RI15b62bc8_1234 , n348 );
buf ( RI15b606c0_1155 , n349 );
buf ( RI15b4a370_397 , n590 );
buf ( RI15b4a3e8_398 , n589 );
buf ( RI15b4a460_399 , n588 );
buf ( RI15b4a4d8_400 , n587 );
buf ( RI15b4a550_401 , n586 );
buf ( RI15b4a5c8_402 , n585 );
buf ( RI15b4a640_403 , n584 );
buf ( RI15b4a6b8_404 , n583 );
buf ( RI15b4a730_405 , n582 );
buf ( RI15b4a7a8_406 , n581 );
buf ( RI15b4a820_407 , n580 );
buf ( RI15b4a898_408 , n579 );
buf ( RI15b4a910_409 , n578 );
buf ( RI15b4a988_410 , n577 );
buf ( RI15b4a2f8_396 , n591 );
buf ( RI15b4aa00_411 , n576 );
buf ( RI15b4aa78_412 , n575 );
buf ( RI15b4aaf0_413 , n574 );
buf ( RI15b4ab68_414 , n573 );
buf ( RI15b4abe0_415 , n572 );
buf ( RI15b4ac58_416 , n571 );
buf ( RI15b4acd0_417 , n570 );
buf ( RI15b4ad48_418 , n569 );
buf ( RI15b4adc0_419 , n568 );
buf ( RI15b4ae38_420 , n567 );
buf ( RI15b4aeb0_421 , n566 );
buf ( RI15b4af28_422 , n565 );
buf ( RI15b4afa0_423 , n564 );
buf ( RI15b4b018_424 , n563 );
buf ( RI15b4a280_395 , n592 );
buf ( RI15b44d30_213 , n354 );
buf ( RI15b44cb8_212 , n352 );
buf ( RI15b44da8_214 , n355 );
buf ( RI15b44e20_215 , n353 );
buf ( RI15b47df0_317 , n500 );
buf ( RI15b4b090_425 , n351 );
buf ( RI15b4b108_426 , n562 );
buf ( RI15b4a0a0_391 , n533 );
buf ( RI15b49380_363 , n561 );
buf ( RI15b493f8_364 , n560 );
buf ( RI15b49470_365 , n559 );
buf ( RI15b494e8_366 , n558 );
buf ( RI15b49560_367 , n557 );
buf ( RI15b495d8_368 , n556 );
buf ( RI15b49650_369 , n555 );
buf ( RI15b496c8_370 , n554 );
buf ( RI15b49740_371 , n553 );
buf ( RI15b497b8_372 , n552 );
buf ( RI15b49830_373 , n551 );
buf ( RI15b498a8_374 , n550 );
buf ( RI15b49920_375 , n549 );
buf ( RI15b49998_376 , n548 );
buf ( RI15b49a10_377 , n547 );
buf ( RI15b49a88_378 , n546 );
buf ( RI15b49b00_379 , n545 );
buf ( RI15b49b78_380 , n544 );
buf ( RI15b49bf0_381 , n543 );
buf ( RI15b49c68_382 , n542 );
buf ( RI15b49ce0_383 , n541 );
buf ( RI15b49d58_384 , n540 );
buf ( RI15b49dd0_385 , n539 );
buf ( RI15b49e48_386 , n538 );
buf ( RI15b49ec0_387 , n537 );
buf ( RI15b49f38_388 , n536 );
buf ( RI15b49fb0_389 , n535 );
buf ( RI15b4a028_390 , n534 );
buf ( RI15b4a118_392 , n532 );
buf ( RI15b42918_136 , n403 );
buf ( RI15b449e8_206 , n365 );
buf ( RI15b44a60_207 , n363 );
buf ( RI15b44b50_209 , n359 );
buf ( RI15b44ad8_208 , n361 );
buf ( RI15b44bc8_210 , n357 );
buf ( RI15b41298_88 , n409 );
buf ( RI15b40ed8_80 , n410 );
buf ( RI15b41658_96 , n408 );
buf ( RI15b40758_64 , n412 );
buf ( RI15b41a18_104 , n407 );
buf ( RI15b42198_120 , n405 );
buf ( RI15b42558_128 , n404 );
buf ( RI15b42cd8_144 , n402 );
buf ( RI15b43098_152 , n401 );
buf ( RI15b43458_160 , n400 );
buf ( RI15b43818_168 , n399 );
buf ( RI15b41dd8_112 , n406 );
buf ( RI15b40b18_72 , n411 );
buf ( RI15b40398_56 , n413 );
buf ( RI15b3ffd8_48 , n414 );
buf ( RI15b432f0_157 , n481 );
buf ( RI15b42f30_149 , n482 );
buf ( RI15b43a70_173 , n479 );
buf ( RI15b436b0_165 , n480 );
buf ( RI15b42030_117 , n486 );
buf ( RI15b40d70_77 , n491 );
buf ( RI15b405f0_61 , n493 );
buf ( RI15b40230_53 , n494 );
buf ( RI15b42b70_141 , n483 );
buf ( RI15b414f0_93 , n489 );
buf ( RI15b41130_85 , n490 );
buf ( RI15b418b0_101 , n488 );
buf ( RI15b409b0_69 , n492 );
buf ( RI15b41c70_109 , n487 );
buf ( RI15b423f0_125 , n485 );
buf ( RI15b427b0_133 , n484 );
buf ( RI15b43110_153 , n417 );
buf ( RI15b42d50_145 , n418 );
buf ( RI15b43890_169 , n415 );
buf ( RI15b434d0_161 , n416 );
buf ( RI15b41e50_113 , n422 );
buf ( RI15b40b90_73 , n427 );
buf ( RI15b40410_57 , n429 );
buf ( RI15b40050_49 , n430 );
buf ( RI15b42990_137 , n419 );
buf ( RI15b41310_89 , n425 );
buf ( RI15b40f50_81 , n426 );
buf ( RI15b416d0_97 , n424 );
buf ( RI15b407d0_65 , n428 );
buf ( RI15b41a90_105 , n423 );
buf ( RI15b42210_121 , n421 );
buf ( RI15b425d0_129 , n420 );
buf ( RI15b42828_134 , n371 );
buf ( RI15b411a8_86 , n377 );
buf ( RI15b40de8_78 , n378 );
buf ( RI15b41568_94 , n376 );
buf ( RI15b40668_62 , n380 );
buf ( RI15b41928_102 , n375 );
buf ( RI15b420a8_118 , n373 );
buf ( RI15b42468_126 , n372 );
buf ( RI15b42be8_142 , n370 );
buf ( RI15b42fa8_150 , n369 );
buf ( RI15b43368_158 , n368 );
buf ( RI15b43728_166 , n367 );
buf ( RI15b41ce8_110 , n374 );
buf ( RI15b40a28_70 , n379 );
buf ( RI15b402a8_54 , n381 );
buf ( RI15b3fee8_46 , n382 );
buf ( RI15b42a08_138 , n435 );
buf ( RI15b41388_90 , n441 );
buf ( RI15b40fc8_82 , n442 );
buf ( RI15b41748_98 , n440 );
buf ( RI15b40848_66 , n444 );
buf ( RI15b41b08_106 , n439 );
buf ( RI15b42288_122 , n437 );
buf ( RI15b42648_130 , n436 );
buf ( RI15b42dc8_146 , n434 );
buf ( RI15b43188_154 , n433 );
buf ( RI15b43548_162 , n432 );
buf ( RI15b43908_170 , n431 );
buf ( RI15b41ec8_114 , n438 );
buf ( RI15b40c08_74 , n443 );
buf ( RI15b400c8_50 , n446 );
buf ( RI15b40488_58 , n445 );
buf ( RI15b428a0_135 , n387 );
buf ( RI15b41220_87 , n393 );
buf ( RI15b40e60_79 , n394 );
buf ( RI15b415e0_95 , n392 );
buf ( RI15b406e0_63 , n396 );
buf ( RI15b419a0_103 , n391 );
buf ( RI15b42120_119 , n389 );
buf ( RI15b424e0_127 , n388 );
buf ( RI15b42c60_143 , n386 );
buf ( RI15b43020_151 , n385 );
buf ( RI15b433e0_159 , n384 );
buf ( RI15b437a0_167 , n383 );
buf ( RI15b41d60_111 , n390 );
buf ( RI15b40aa0_71 , n395 );
buf ( RI15b3ff60_47 , n398 );
buf ( RI15b40320_55 , n397 );
buf ( RI15b42e40_147 , n450 );
buf ( RI15b43200_155 , n449 );
buf ( RI15b43980_171 , n447 );
buf ( RI15b435c0_163 , n448 );
buf ( RI15b41f40_115 , n454 );
buf ( RI15b40c80_75 , n459 );
buf ( RI15b40500_59 , n461 );
buf ( RI15b40140_51 , n462 );
buf ( RI15b41b80_107 , n455 );
buf ( RI15b42300_123 , n453 );
buf ( RI15b426c0_131 , n452 );
buf ( RI15b41400_91 , n457 );
buf ( RI15b42a80_139 , n451 );
buf ( RI15b417c0_99 , n456 );
buf ( RI15b408c0_67 , n460 );
buf ( RI15b41040_83 , n458 );
buf ( RI15b42af8_140 , n467 );
buf ( RI15b41478_92 , n473 );
buf ( RI15b410b8_84 , n474 );
buf ( RI15b41838_100 , n472 );
buf ( RI15b40938_68 , n476 );
buf ( RI15b41bf8_108 , n471 );
buf ( RI15b42378_124 , n469 );
buf ( RI15b42738_132 , n468 );
buf ( RI15b42eb8_148 , n466 );
buf ( RI15b43278_156 , n465 );
buf ( RI15b43638_164 , n464 );
buf ( RI15b439f8_172 , n463 );
buf ( RI15b41fb8_116 , n470 );
buf ( RI15b40cf8_76 , n475 );
buf ( RI15b40578_60 , n477 );
buf ( RI15b401b8_52 , n478 );
buf ( RI15b3fd80_43 , n360 );
buf ( RI15b3fc90_41 , n364 );
buf ( RI15b3fd08_42 , n362 );
buf ( RI15b3fe70_45 , n356 );
buf ( RI15b3fdf8_44 , n358 );
buf ( RI15b3fba0_39 , n499 );
buf ( RI15b668b8_1364 , n498 );
buf ( RI15b4a208_394 , n531 );
buf ( RI15b48390_329 , n496 );
buf ( RI15b48408_330 , n497 );
buf ( RI15b48318_328 , n495 );
buf ( RI15b4a190_393 , n501 );
buf ( RI15b4b2e8_430 , n528 );
buf ( RI15b4b1f8_428 , n530 );
buf ( RI15b4b270_429 , n529 );
buf ( RI15b4b360_431 , n527 );
buf ( RI15b4b3d8_432 , n526 );
buf ( RI15b4b450_433 , n525 );
buf ( RI15b4b4c8_434 , n524 );
buf ( RI15b4b540_435 , n523 );
buf ( RI15b4b5b8_436 , n522 );
buf ( RI15b4b630_437 , n521 );
buf ( RI15b4b6a8_438 , n520 );
buf ( RI15b4b720_439 , n519 );
buf ( RI15b4b798_440 , n518 );
buf ( RI15b4b888_442 , n516 );
buf ( RI15b4b810_441 , n517 );
buf ( RI15b4b900_443 , n515 );
buf ( RI15b4b978_444 , n514 );
buf ( RI15b4b9f0_445 , n513 );
buf ( RI15b4ba68_446 , n512 );
buf ( RI15b4bae0_447 , n511 );
buf ( RI15b4bb58_448 , n510 );
buf ( RI15b4bbd0_449 , n509 );
buf ( RI15b4bc48_450 , n508 );
buf ( RI15b4bcc0_451 , n507 );
buf ( RI15b4bd38_452 , n506 );
buf ( RI15b4bdb0_453 , n505 );
buf ( RI15b4be28_454 , n504 );
buf ( RI15b4bea0_455 , n503 );
buf ( RI15b4bf18_456 , n502 );
buf ( RI15b4bf90_457 , n366 );
buf ( RI15b508b0_613 , n594 );
buf ( RI15b4ffc8_594 , n613 );
buf ( RI15b50040_595 , n612 );
buf ( RI15b500b8_596 , n611 );
buf ( RI15b50130_597 , n610 );
buf ( RI15b501a8_598 , n609 );
buf ( RI15b50220_599 , n608 );
buf ( RI15b50298_600 , n607 );
buf ( RI15b50310_601 , n606 );
buf ( RI15b50388_602 , n605 );
buf ( RI15b50400_603 , n604 );
buf ( RI15b50478_604 , n603 );
buf ( RI15b504f0_605 , n602 );
buf ( RI15b50568_606 , n601 );
buf ( RI15b505e0_607 , n600 );
buf ( RI15b50658_608 , n599 );
buf ( RI15b506d0_609 , n598 );
buf ( RI15b50748_610 , n597 );
buf ( RI15b507c0_611 , n596 );
buf ( RI15b50838_612 , n595 );
buf ( RI15b4ff50_593 , n614 );
buf ( RI15b50928_614 , n593 );
buf ( RI15b57fc0_867 , n615 );
buf ( RI15b577c8_850 , n630 );
buf ( RI15b57840_851 , n629 );
buf ( RI15b578b8_852 , n628 );
buf ( RI15b57930_853 , n627 );
buf ( RI15b579a8_854 , n626 );
buf ( RI15b57a20_855 , n625 );
buf ( RI15b57a98_856 , n624 );
buf ( RI15b57b10_857 , n623 );
buf ( RI15b57b88_858 , n622 );
buf ( RI15b57c00_859 , n621 );
buf ( RI15b57c78_860 , n620 );
buf ( RI15b57cf0_861 , n619 );
buf ( RI15b57de0_863 , n616 );
buf ( RI15b559c8_786 , n643 );
buf ( RI15b55a40_787 , n642 );
buf ( RI15b55ab8_788 , n641 );
buf ( RI15b55b30_789 , n640 );
buf ( RI15b55ba8_790 , n639 );
buf ( RI15b55c20_791 , n638 );
buf ( RI15b55c98_792 , n637 );
buf ( RI15b55d10_793 , n636 );
buf ( RI15b55d88_794 , n635 );
buf ( RI15b55e00_795 , n634 );
buf ( RI15b55e78_796 , n633 );
buf ( RI15b55ef0_797 , n632 );
buf ( RI15b55f68_798 , n631 );
buf ( RI15b55fe0_799 , n617 );
buf ( RI15b57d68_862 , n618 );
buf ( RI15b66408_1354 , n667 );
buf ( RI15b65850_1329 , n644 );
buf ( RI15b658c8_1330 , n646 );
buf ( RI15b65940_1331 , n647 );
buf ( RI15b659b8_1332 , n648 );
buf ( RI15b65a30_1333 , n649 );
buf ( RI15b65aa8_1334 , n650 );
buf ( RI15b65b20_1335 , n651 );
buf ( RI15b65b98_1336 , n652 );
buf ( RI15b65c10_1337 , n661 );
buf ( RI15b65c88_1338 , n660 );
buf ( RI15b65d00_1339 , n659 );
buf ( RI15b65d78_1340 , n658 );
buf ( RI15b65df0_1341 , n657 );
buf ( RI15b65e68_1342 , n656 );
buf ( RI15b65ee0_1343 , n655 );
buf ( RI15b65f58_1344 , n654 );
buf ( RI15b65fd0_1345 , n653 );
buf ( RI15b66048_1346 , n675 );
buf ( RI15b660c0_1347 , n674 );
buf ( RI15b66138_1348 , n673 );
buf ( RI15b661b0_1349 , n672 );
buf ( RI15b66228_1350 , n671 );
buf ( RI15b662a0_1351 , n670 );
buf ( RI15b66318_1352 , n669 );
buf ( RI15b66390_1353 , n668 );
buf ( RI15b66480_1355 , n666 );
buf ( RI15b666d8_1360 , n645 );
buf ( RI15b664f8_1356 , n665 );
buf ( RI15b66570_1357 , n664 );
buf ( RI15b3fb28_38 , n682 );
buf ( RI15b66750_1361 , n681 );
buf ( RI15b60be8_1166 , n678 );
buf ( RI15b60c60_1167 , n679 );
buf ( RI15b60cd8_1168 , n680 );
buf ( RI15b63a50_1265 , n677 );
buf ( RI15b61c50_1201 , n683 );
buf ( RI15b62b50_1233 , n676 );
buf ( RI15b56058_800 , n709 );
buf ( RI15b560d0_801 , n708 );
buf ( RI15b56148_802 , n707 );
buf ( RI15b561c0_803 , n706 );
buf ( RI15b56238_804 , n705 );
buf ( RI15b562b0_805 , n704 );
buf ( RI15b56328_806 , n703 );
buf ( RI15b563a0_807 , n702 );
buf ( RI15b56418_808 , n701 );
buf ( RI15b56490_809 , n700 );
buf ( RI15b56508_810 , n699 );
buf ( RI15b56580_811 , n698 );
buf ( RI15b565f8_812 , n697 );
buf ( RI15b58470_877 , n684 );
buf ( RI15b583f8_876 , n685 );
buf ( RI15b57e58_864 , n696 );
buf ( RI15b57ed0_865 , n695 );
buf ( RI15b57f48_866 , n694 );
buf ( RI15b58038_868 , n693 );
buf ( RI15b580b0_869 , n692 );
buf ( RI15b58128_870 , n691 );
buf ( RI15b581a0_871 , n690 );
buf ( RI15b58218_872 , n689 );
buf ( RI15b58290_873 , n688 );
buf ( RI15b58308_874 , n687 );
buf ( RI15b58380_875 , n686 );
buf ( RI15b60648_1154 , n711 );
buf ( RI15b605d0_1153 , n710 );
buf ( RI15b47d78_316 , n715 );
buf ( RI15b47d00_315 , n714 );
buf ( RI15b541e0_735 , n713 );
buf ( RI15b54168_734 , n712 );
buf ( RI15b450f0_221 , n717 );
buf ( RI15b51558_640 , n716 );
buf ( RI15b4c008_458 , n718 );
buf ( RI15b63d98_1272 , n719 );
buf ( RI15b575e8_846 , n720 );
buf ( RI15b63ac8_1266 , n722 );
buf ( RI15b648d8_1296 , n721 );
buf ( RI15b63b40_1267 , n749 );
buf ( RI15b64860_1295 , n723 );
buf ( RI15b63c30_1269 , n747 );
buf ( RI15b63ca8_1270 , n746 );
buf ( RI15b63bb8_1268 , n748 );
buf ( RI15b63e88_1274 , n744 );
buf ( RI15b63f00_1275 , n743 );
buf ( RI15b63d20_1271 , n745 );
buf ( RI15b63f78_1276 , n742 );
buf ( RI15b63ff0_1277 , n741 );
buf ( RI15b64068_1278 , n740 );
buf ( RI15b640e0_1279 , n739 );
buf ( RI15b64158_1280 , n738 );
buf ( RI15b641d0_1281 , n737 );
buf ( RI15b64248_1282 , n736 );
buf ( RI15b642c0_1283 , n735 );
buf ( RI15b64338_1284 , n734 );
buf ( RI15b643b0_1285 , n733 );
buf ( RI15b64428_1286 , n732 );
buf ( RI15b644a0_1287 , n731 );
buf ( RI15b64518_1288 , n730 );
buf ( RI15b64590_1289 , n729 );
buf ( RI15b64608_1290 , n728 );
buf ( RI15b64680_1291 , n727 );
buf ( RI15b646f8_1292 , n726 );
buf ( RI15b64770_1293 , n725 );
buf ( RI15b647e8_1294 , n724 );
buf ( RI15b5d948_1058 , n750 );
buf ( RI15b484f8_332 , n754 );
buf ( RI15b467e8_270 , n751 );
buf ( RI15b5e5f0_1085 , n769 );
buf ( RI15b5ddf8_1068 , n780 );
buf ( RI15b5de70_1069 , n781 );
buf ( RI15b5dee8_1070 , n782 );
buf ( RI15b5df60_1071 , n783 );
buf ( RI15b5dfd8_1072 , n784 );
buf ( RI15b5e050_1073 , n785 );
buf ( RI15b5e0c8_1074 , n786 );
buf ( RI15b5e140_1075 , n787 );
buf ( RI15b5da38_1060 , n772 );
buf ( RI15b5dab0_1061 , n773 );
buf ( RI15b5db28_1062 , n774 );
buf ( RI15b5dba0_1063 , n775 );
buf ( RI15b5e398_1080 , n792 );
buf ( RI15b5e410_1081 , n793 );
buf ( RI15b5e488_1082 , n794 );
buf ( RI15b5e500_1083 , n795 );
buf ( RI15b5dc18_1064 , n776 );
buf ( RI15b5dc90_1065 , n777 );
buf ( RI15b5dd08_1066 , n778 );
buf ( RI15b5dd80_1067 , n779 );
buf ( RI15b5e1b8_1076 , n788 );
buf ( RI15b5e230_1077 , n789 );
buf ( RI15b5e2a8_1078 , n790 );
buf ( RI15b5e320_1079 , n791 );
buf ( RI15b5e578_1084 , n796 );
buf ( RI15b5d9c0_1059 , n771 );
buf ( RI15b5e668_1086 , n797 );
buf ( RI15b5e6e0_1087 , n770 );
buf ( RI15b657d8_1328 , n801 );
buf ( RI15b3eac0_3 , n800 );
buf ( RI15b64ab8_1300 , n807 );
buf ( RI15b3f7e0_31 , n806 );
buf ( RI15b64b30_1301 , n809 );
buf ( RI15b3f768_30 , n808 );
buf ( RI15b64ba8_1302 , n811 );
buf ( RI15b3f6f0_29 , n810 );
buf ( RI15b649c8_1298 , n803 );
buf ( RI15b3f8d0_33 , n802 );
buf ( RI15b64950_1297 , n799 );
buf ( RI15b3f948_34 , n798 );
buf ( RI15b64a40_1299 , n805 );
buf ( RI15b3f858_32 , n804 );
buf ( RI15b64c20_1303 , n813 );
buf ( RI15b3f678_28 , n812 );
buf ( RI15b64c98_1304 , n815 );
buf ( RI15b3f600_27 , n814 );
buf ( RI15b64d10_1305 , n833 );
buf ( RI15b3f588_26 , n832 );
buf ( RI15b64d88_1306 , n831 );
buf ( RI15b3f510_25 , n830 );
buf ( RI15b64e00_1307 , n829 );
buf ( RI15b3f498_24 , n828 );
buf ( RI15b64e78_1308 , n827 );
buf ( RI15b3f420_23 , n826 );
buf ( RI15b64ef0_1309 , n825 );
buf ( RI15b3f3a8_22 , n824 );
buf ( RI15b64f68_1310 , n823 );
buf ( RI15b3f330_21 , n822 );
buf ( RI15b64fe0_1311 , n821 );
buf ( RI15b3f2b8_20 , n820 );
buf ( RI15b65058_1312 , n819 );
buf ( RI15b3f240_19 , n818 );
buf ( RI15b650d0_1313 , n817 );
buf ( RI15b3f1c8_18 , n816 );
buf ( RI15b65148_1314 , n861 );
buf ( RI15b3f150_17 , n860 );
buf ( RI15b65328_1318 , n853 );
buf ( RI15b3ef70_13 , n852 );
buf ( RI15b65238_1316 , n857 );
buf ( RI15b3f060_15 , n856 );
buf ( RI15b652b0_1317 , n855 );
buf ( RI15b3efe8_14 , n854 );
buf ( RI15b651c0_1315 , n859 );
buf ( RI15b3f0d8_16 , n858 );
buf ( RI15b65490_1321 , n847 );
buf ( RI15b3ee08_10 , n846 );
buf ( RI15b65508_1322 , n845 );
buf ( RI15b3ed90_9 , n844 );
buf ( RI15b3eef8_12 , n850 );
buf ( RI15b653a0_1319 , n851 );
buf ( RI15b65418_1320 , n849 );
buf ( RI15b3ee80_11 , n848 );
buf ( RI15b65580_1323 , n843 );
buf ( RI15b655f8_1324 , n841 );
buf ( RI15b3eca0_7 , n840 );
buf ( RI15b3ed18_8 , n842 );
buf ( RI15b3ec28_6 , n838 );
buf ( RI15b65670_1325 , n839 );
buf ( RI15b656e8_1326 , n837 );
buf ( RI15b3ebb0_5 , n836 );
buf ( RI15b65760_1327 , n835 );
buf ( RI15b3eb38_4 , n834 );
buf ( RI15b5c7f0_1021 , n863 );
buf ( RI15b62f88_1242 , n862 );
buf ( RI15b479b8_308 , n864 );
buf ( RI15b665e8_1358 , n663 );
buf ( RI15b47b98_312 , n865 );
buf ( RI15b523e0_671 , n868 );
buf ( RI15b51300_635 , n871 );
buf ( RI15b51378_636 , n872 );
buf ( RI15b513f0_637 , n873 );
buf ( RI15b51468_638 , n874 );
buf ( RI15b52368_670 , n869 );
buf ( RI15b522f0_669 , n870 );
buf ( RI15b52458_672 , n867 );
buf ( RI15b52278_668 , n866 );
buf ( RI15b534c0_707 , n875 );
buf ( RI15b515d0_641 , n895 );
buf ( RI15b51648_642 , n896 );
buf ( RI15b516c0_643 , n897 );
buf ( RI15b51738_644 , n898 );
buf ( RI15b517b0_645 , n899 );
buf ( RI15b51828_646 , n900 );
buf ( RI15b518a0_647 , n901 );
buf ( RI15b51918_648 , n902 );
buf ( RI15b52110_665 , n919 );
buf ( RI15b52188_666 , n920 );
buf ( RI15b514e0_639 , n894 );
buf ( RI15b52200_667 , n921 );
buf ( RI15b51990_649 , n903 );
buf ( RI15b51a08_650 , n904 );
buf ( RI15b51a80_651 , n905 );
buf ( RI15b51af8_652 , n906 );
buf ( RI15b51b70_653 , n907 );
buf ( RI15b51be8_654 , n908 );
buf ( RI15b51c60_655 , n909 );
buf ( RI15b51cd8_656 , n910 );
buf ( RI15b51d50_657 , n911 );
buf ( RI15b51dc8_658 , n912 );
buf ( RI15b51e40_659 , n913 );
buf ( RI15b51eb8_660 , n914 );
buf ( RI15b51f30_661 , n915 );
buf ( RI15b51fa8_662 , n916 );
buf ( RI15b52020_663 , n917 );
buf ( RI15b52098_664 , n918 );
buf ( RI15b548e8_750 , n877 );
buf ( RI15b54b40_755 , n883 );
buf ( RI15b54bb8_756 , n884 );
buf ( RI15b54960_751 , n879 );
buf ( RI15b549d8_752 , n880 );
buf ( RI15b54a50_753 , n881 );
buf ( RI15b54ac8_754 , n882 );
buf ( RI15b55770_781 , n878 );
buf ( RI15b54c30_757 , n885 );
buf ( RI15b54ca8_758 , n886 );
buf ( RI15b52f98_696 , n876 );
buf ( RI15b509a0_615 , n925 );
buf ( RI15b50a18_616 , n924 );
buf ( RI15b50a90_617 , n923 );
buf ( RI15b50b08_618 , n922 );
buf ( RI15b46e00_283 , n926 );
buf ( RI15b48480_331 , n752 );
buf ( RI15b486d8_336 , n758 );
buf ( RI15b48570_333 , n755 );
buf ( RI15b48750_337 , n759 );
buf ( RI15b488b8_340 , n762 );
buf ( RI15b48a20_343 , n765 );
buf ( RI15b48930_341 , n763 );
buf ( RI15b48a98_344 , n766 );
buf ( RI15b48660_335 , n757 );
buf ( RI15b485e8_334 , n756 );
buf ( RI15b48840_339 , n761 );
buf ( RI15b487c8_338 , n760 );
buf ( RI15b489a8_342 , n764 );
buf ( RI15b48b10_345 , n767 );
buf ( RI15b49308_362 , n753 );
buf ( RI15b48228_326 , n928 );
buf ( RI15b482a0_327 , n929 );
buf ( RI15b4b180_427 , n927 );
buf ( RI15b45348_226 , n930 );
buf ( RI15b4c080_459 , n931 );
buf ( RI15b54d20_759 , n887 );
buf ( RI15b54d98_760 , n888 );
buf ( RI15b54e10_761 , n889 );
buf ( RI15b54e88_762 , n890 );
buf ( RI15b54f00_763 , n891 );
buf ( RI15b54f78_764 , n892 );
buf ( RI15b54ff0_765 , n893 );
buf ( RI15b55068_766 , n945 );
buf ( RI15b550e0_767 , n944 );
buf ( RI15b55158_768 , n943 );
buf ( RI15b551d0_769 , n942 );
buf ( RI15b55248_770 , n941 );
buf ( RI15b552c0_771 , n940 );
buf ( RI15b55338_772 , n939 );
buf ( RI15b553b0_773 , n938 );
buf ( RI15b554a0_775 , n936 );
buf ( RI15b55428_774 , n937 );
buf ( RI15b55518_776 , n935 );
buf ( RI15b55590_777 , n934 );
buf ( RI15b55608_778 , n933 );
buf ( RI15b55680_779 , n932 );
buf ( RI15b52908_682 , n946 );
buf ( RI15b53f10_729 , n947 );
buf ( RI15b556f8_780 , n948 );
buf ( RI15b52b60_687 , n949 );
buf ( RI15b61cc8_1202 , n952 );
buf ( RI15b62ad8_1232 , n951 );
buf ( RI15b61d40_1203 , n950 );
buf ( RI15b63528_1254 , n963 );
buf ( RI15b635a0_1255 , n962 );
buf ( RI15b63618_1256 , n961 );
buf ( RI15b63690_1257 , n960 );
buf ( RI15b63708_1258 , n959 );
buf ( RI15b63780_1259 , n958 );
buf ( RI15b637f8_1260 , n957 );
buf ( RI15b63870_1261 , n956 );
buf ( RI15b638e8_1262 , n955 );
buf ( RI15b63960_1263 , n954 );
buf ( RI15b63168_1246 , n971 );
buf ( RI15b631e0_1247 , n970 );
buf ( RI15b63258_1248 , n969 );
buf ( RI15b632d0_1249 , n968 );
buf ( RI15b63348_1250 , n967 );
buf ( RI15b633c0_1251 , n966 );
buf ( RI15b63438_1252 , n965 );
buf ( RI15b63000_1243 , n974 );
buf ( RI15b63078_1244 , n973 );
buf ( RI15b630f0_1245 , n972 );
buf ( RI15b634b0_1253 , n964 );
buf ( RI15b639d8_1264 , n953 );
buf ( RI15b60d50_1169 , n977 );
buf ( RI15b60fa8_1174 , n983 );
buf ( RI15b61020_1175 , n984 );
buf ( RI15b60dc8_1170 , n979 );
buf ( RI15b60e40_1171 , n980 );
buf ( RI15b60eb8_1172 , n981 );
buf ( RI15b60f30_1173 , n982 );
buf ( RI15b61bd8_1200 , n978 );
buf ( RI15b61098_1176 , n985 );
buf ( RI15b61110_1177 , n986 );
buf ( RI15b61188_1178 , n987 );
buf ( RI15b61200_1179 , n988 );
buf ( RI15b61278_1180 , n989 );
buf ( RI15b612f0_1181 , n990 );
buf ( RI15b61368_1182 , n991 );
buf ( RI15b5fdd8_1136 , n976 );
buf ( RI15b5f658_1120 , n975 );
buf ( RI15b66660_1359 , n662 );
buf ( RI15b62100_1211 , n994 );
buf ( RI15b61db8_1204 , n1001 );
buf ( RI15b61e30_1205 , n1000 );
buf ( RI15b61ea8_1206 , n999 );
buf ( RI15b61f20_1207 , n998 );
buf ( RI15b61f98_1208 , n997 );
buf ( RI15b62010_1209 , n996 );
buf ( RI15b62088_1210 , n995 );
buf ( RI15b45438_228 , n1002 );
buf ( RI15b477d8_304 , n1003 );
buf ( RI15b5c868_1022 , n1019 );
buf ( RI15b5c8e0_1023 , n1018 );
buf ( RI15b5c958_1024 , n1017 );
buf ( RI15b5c9d0_1025 , n1016 );
buf ( RI15b5ca48_1026 , n1015 );
buf ( RI15b5cac0_1027 , n1014 );
buf ( RI15b5cb38_1028 , n1013 );
buf ( RI15b5cbb0_1029 , n1012 );
buf ( RI15b5cc28_1030 , n1011 );
buf ( RI15b5cca0_1031 , n1010 );
buf ( RI15b5cd18_1032 , n1009 );
buf ( RI15b5cd90_1033 , n1008 );
buf ( RI15b5ce08_1034 , n1007 );
buf ( RI15b5ce80_1035 , n1006 );
buf ( RI15b5cef8_1036 , n1005 );
buf ( RI15b5cf70_1037 , n1004 );
buf ( RI15b5f388_1114 , n1020 );
buf ( RI15b3f9c0_35 , n1022 );
buf ( RI15b60738_1156 , n1021 );
buf ( RI15b3fa38_36 , n1023 );
buf ( RI15b5e848_1090 , n1025 );
buf ( RI15b60828_1158 , n1024 );
buf ( RI15b470d0_289 , n1027 );
buf ( RI15b46950_273 , n1026 );
buf ( RI15b43bd8_176 , n1055 );
buf ( RI15b43c50_177 , n1054 );
buf ( RI15b43cc8_178 , n1053 );
buf ( RI15b43b60_175 , n1056 );
buf ( RI15b43d40_179 , n1052 );
buf ( RI15b43db8_180 , n1051 );
buf ( RI15b43e30_181 , n1050 );
buf ( RI15b43ea8_182 , n1049 );
buf ( RI15b43f20_183 , n1048 );
buf ( RI15b43f98_184 , n1047 );
buf ( RI15b44010_185 , n1046 );
buf ( RI15b44268_190 , n1041 );
buf ( RI15b44088_186 , n1045 );
buf ( RI15b44100_187 , n1044 );
buf ( RI15b44178_188 , n1043 );
buf ( RI15b441f0_189 , n1042 );
buf ( RI15b43ae8_174 , n1057 );
buf ( RI15b442e0_191 , n1040 );
buf ( RI15b44358_192 , n1039 );
buf ( RI15b443d0_193 , n1038 );
buf ( RI15b445b0_197 , n1034 );
buf ( RI15b44448_194 , n1037 );
buf ( RI15b444c0_195 , n1036 );
buf ( RI15b44538_196 , n1035 );
buf ( RI15b44628_198 , n1033 );
buf ( RI15b446a0_199 , n1032 );
buf ( RI15b44718_200 , n1031 );
buf ( RI15b44790_201 , n1030 );
buf ( RI15b44808_202 , n1029 );
buf ( RI15b44880_203 , n1028 );
buf ( RI15b62178_1212 , n1078 );
buf ( RI15b621f0_1213 , n1077 );
buf ( RI15b62268_1214 , n1076 );
buf ( RI15b622e0_1215 , n1075 );
buf ( RI15b62358_1216 , n1074 );
buf ( RI15b623d0_1217 , n1073 );
buf ( RI15b62448_1218 , n1072 );
buf ( RI15b624c0_1219 , n1071 );
buf ( RI15b62538_1220 , n1070 );
buf ( RI15b625b0_1221 , n1069 );
buf ( RI15b62628_1222 , n1068 );
buf ( RI15b626a0_1223 , n1067 );
buf ( RI15b62718_1224 , n1066 );
buf ( RI15b62790_1225 , n1065 );
buf ( RI15b62808_1226 , n1064 );
buf ( RI15b62880_1227 , n1063 );
buf ( RI15b628f8_1228 , n1062 );
buf ( RI15b62970_1229 , n1061 );
buf ( RI15b629e8_1230 , n1060 );
buf ( RI15b62a60_1231 , n1059 );
buf ( RI15b613e0_1183 , n992 );
buf ( RI15b5cfe8_1038 , n1084 );
buf ( RI15b5d060_1039 , n1083 );
buf ( RI15b5d0d8_1040 , n1082 );
buf ( RI15b5d150_1041 , n1081 );
buf ( RI15b5d1c8_1042 , n1080 );
buf ( RI15b45618_232 , n1085 );
buf ( RI15b53538_708 , n1094 );
buf ( RI15b5d768_1054 , n1090 );
buf ( RI15b5d7e0_1055 , n1091 );
buf ( RI15b5d858_1056 , n1092 );
buf ( RI15b5d8d0_1057 , n1093 );
buf ( RI15b5e758_1088 , n1089 );
buf ( RI15b5e7d0_1089 , n1088 );
buf ( RI15b5e8c0_1091 , n1087 );
buf ( RI15b5f9a0_1127 , n1095 );
buf ( RI15b615c0_1187 , n1110 );
buf ( RI15b61458_1184 , n993 );
buf ( RI15b614d0_1185 , n1097 );
buf ( RI15b61548_1186 , n1111 );
buf ( RI15b61638_1188 , n1109 );
buf ( RI15b616b0_1189 , n1108 );
buf ( RI15b61728_1190 , n1107 );
buf ( RI15b617a0_1191 , n1106 );
buf ( RI15b5ec08_1098 , n1096 );
buf ( RI15b526b0_677 , n1112 );
buf ( RI15b46ba8_278 , n1115 );
buf ( RI15b53f88_730 , n1117 );
buf ( RI15b603f0_1149 , n1118 );
buf ( RI15b45d98_248 , n1119 );
buf ( RI15b475f8_300 , n1126 );
buf ( RI15b3fab0_37 , n1127 );
buf ( RI15b45168_222 , n1128 );
buf ( RI15b542d0_737 , n1129 );
buf ( RI15b45ac8_242 , n1130 );
buf ( RI15b527a0_679 , n1131 );
buf ( RI15b53808_714 , n1133 );
buf ( RI15b53088_698 , n1132 );
buf ( RI15b61818_1192 , n1105 );
buf ( RI15b61890_1193 , n1104 );
buf ( RI15b61908_1194 , n1103 );
buf ( RI15b61980_1195 , n1102 );
buf ( RI15b619f8_1196 , n1101 );
buf ( RI15b60468_1150 , n1135 );
buf ( RI15b5ee60_1103 , n1134 );
buf ( RI15b54618_744 , n1136 );
buf ( RI15b54708_746 , n1137 );
buf ( RI15b46fe0_287 , n1138 );
buf ( RI15b60918_1160 , n1139 );
buf ( RI15b48b88_346 , n768 );
buf ( RI15b48c00_347 , n1143 );
buf ( RI15b48c78_348 , n1157 );
buf ( RI15b48cf0_349 , n1156 );
buf ( RI15b48d68_350 , n1155 );
buf ( RI15b48de0_351 , n1154 );
buf ( RI15b48e58_352 , n1153 );
buf ( RI15b48ed0_353 , n1152 );
buf ( RI15b48f48_354 , n1151 );
buf ( RI15b48fc0_355 , n1150 );
buf ( RI15b490b0_357 , n1148 );
buf ( RI15b49128_358 , n1147 );
buf ( RI15b49038_356 , n1149 );
buf ( RI15b49290_361 , n1144 );
buf ( RI15b491a0_359 , n1146 );
buf ( RI15b49218_360 , n1145 );
buf ( RI15b460e0_255 , n1141 );
buf ( RI15b476e8_302 , n1142 );
buf ( RI15b53c40_723 , n1159 );
buf ( RI15b52638_676 , n1158 );
buf ( RI15b45f78_252 , n1162 );
buf ( RI15b45e88_250 , n1164 );
buf ( RI15b45f00_251 , n1163 );
buf ( RI15b45ff0_253 , n1161 );
buf ( RI15b44e98_216 , n1165 );
buf ( RI15b44f10_217 , n1166 );
buf ( RI15b44f88_218 , n1167 );
buf ( RI15b45000_219 , n1168 );
buf ( RI15b54258_736 , n1169 );
buf ( RI15b53b50_721 , n1170 );
buf ( RI15b53da8_726 , n1172 );
buf ( RI15b5f220_1111 , n1174 );
buf ( RI15b47328_294 , n1175 );
buf ( RI15b45a50_241 , n1176 );
buf ( RI15b584e8_878 , n1177 );
buf ( RI15b535b0_709 , n1180 );
buf ( RI15b52e30_693 , n1179 );
buf ( RI15b53e20_727 , n1181 );
buf ( RI15b60288_1146 , n1182 );
buf ( RI15b3fc18_40 , n1183 );
buf ( RI15b608a0_1159 , n1186 );
buf ( RI15b45780_235 , n1187 );
buf ( RI15b52cc8_690 , n1114 );
buf ( RI15b525c0_675 , n1188 );
buf ( RI15b47418_296 , n1189 );
buf ( RI15b50b80_619 , n1125 );
buf ( RI15b50bf8_620 , n1124 );
buf ( RI15b50c70_621 , n1123 );
buf ( RI15b50ce8_622 , n1122 );
buf ( RI15b44c40_211 , n1191 );
buf ( RI15b46a40_275 , n1192 );
buf ( RI15b60af8_1164 , n1193 );
buf ( RI15b47f58_320 , n1194 );
buf ( RI15b53718_712 , n1195 );
buf ( RI15b5fb80_1131 , n1196 );
buf ( RI15b45d20_247 , n1198 );
buf ( RI15b52f20_695 , n1199 );
buf ( RI15b47ee0_319 , n1200 );
buf ( RI15b543c0_739 , n1201 );
buf ( RI15b61a70_1197 , n1100 );
buf ( RI15b61ae8_1198 , n1099 );
buf ( RI15b5ef50_1105 , n1202 );
buf ( RI15b5ec80_1099 , n1203 );
buf ( RI15b50d60_623 , n1121 );
buf ( RI15b50dd8_624 , n1120 );
buf ( RI15b53448_706 , n1204 );
buf ( RI15b54000_731 , n1206 );
buf ( RI15b529f8_684 , n1205 );
buf ( RI15b5f838_1124 , n1207 );
buf ( RI15b5f0b8_1108 , n1171 );
buf ( RI15b53880_715 , n1208 );
buf ( RI15b5fce8_1134 , n1209 );
buf ( RI15b46d10_281 , n1210 );
buf ( RI15b52890_681 , n1211 );
buf ( RI15b5fd60_1135 , n1213 );
buf ( RI15b5f5e0_1119 , n1212 );
buf ( RI15b454b0_229 , n1214 );
buf ( RI15b46860_271 , n1215 );
buf ( RI15b540f0_733 , n1218 );
buf ( RI15b60558_1152 , n1219 );
buf ( RI15b47490_297 , n1220 );
buf ( RI15b471c0_291 , n1221 );
buf ( RI15b47238_292 , n1222 );
buf ( RI15b539e8_718 , n1224 );
buf ( RI15b53268_702 , n1223 );
buf ( RI15b5f130_1109 , n1225 );
buf ( RI15b5fb08_1130 , n1226 );
buf ( RI15b607b0_1157 , n1227 );
buf ( RI15b544b0_741 , n1228 );
buf ( RI15b604e0_1151 , n1230 );
buf ( RI15b5eed8_1104 , n1229 );
buf ( RI15b510a8_630 , n1231 );
buf ( RI15b5d240_1043 , n1178 );
buf ( RI15b463b0_261 , n1232 );
buf ( RI15b46428_262 , n1233 );
buf ( RI15b5f298_1112 , n1234 );
buf ( RI15b47a30_309 , n1236 );
buf ( RI15b53bc8_722 , n1237 );
buf ( RI15b46338_260 , n1238 );
buf ( RI15b47c10_313 , n1239 );
buf ( RI15b48048_322 , n1240 );
buf ( RI15b464a0_263 , n1241 );
buf ( RI15b5ecf8_1100 , n1242 );
buf ( RI15b53628_710 , n1244 );
buf ( RI15b52ea8_694 , n1243 );
buf ( RI15b47850_305 , n1245 );
buf ( RI15b47670_301 , n1247 );
buf ( RI15b46068_254 , n1246 );
buf ( RI15b524d0_673 , n1248 );
buf ( RI15b52ae8_686 , n1250 );
buf ( RI15b451e0_223 , n1251 );
buf ( RI15b52548_674 , n1252 );
buf ( RI15b60030_1141 , n1253 );
buf ( RI15b457f8_236 , n1254 );
buf ( RI15b60990_1161 , n1255 );
buf ( RI15b53ad8_720 , n1256 );
buf ( RI15b5ff40_1139 , n1257 );
buf ( RI15b45528_230 , n1258 );
buf ( RI15b5fa18_1128 , n1259 );
buf ( RI15b53358_704 , n1260 );
buf ( RI15b5f7c0_1123 , n1261 );
buf ( RI15b462c0_259 , n1262 );
buf ( RI15b453c0_227 , n1263 );
buf ( RI15b45870_237 , n1264 );
buf ( RI15b46518_264 , n1265 );
buf ( RI15b47058_288 , n1266 );
buf ( RI15b60b70_1165 , n1267 );
buf ( RI15b45bb8_244 , n1268 );
buf ( RI15b533d0_705 , n1269 );
buf ( RI15b47e68_318 , n1270 );
buf ( RI15b44970_205 , n1184 );
buf ( RI15b53100_699 , n1113 );
buf ( RI15b47fd0_321 , n1271 );
buf ( RI15b5f568_1118 , n1272 );
buf ( RI15b480c0_323 , n1273 );
buf ( RI15b45960_239 , n1274 );
buf ( RI15b52980_683 , n1275 );
buf ( RI15b53cb8_724 , n1276 );
buf ( RI15b60120_1143 , n1277 );
buf ( RI15b5f4f0_1117 , n1278 );
buf ( RI15b46248_258 , n1279 );
buf ( RI15b46590_265 , n1281 );
buf ( RI15b5fe50_1137 , n1282 );
buf ( RI15b52c50_689 , n1086 );
buf ( RI15b47aa8_310 , n1283 );
buf ( RI15b47b20_311 , n1284 );
buf ( RI15b61b60_1199 , n1098 );
buf ( RI15b5efc8_1106 , n1285 );
buf ( RI15b468d8_272 , n1160 );
buf ( RI15b60378_1148 , n1286 );
buf ( RI15b5ed70_1101 , n1287 );
buf ( RI15b5f6d0_1121 , n1079 );
buf ( RI15b46c20_279 , n1288 );
buf ( RI15b5d510_1049 , n1289 );
buf ( RI15b46ab8_276 , n1216 );
buf ( RI15b45258_224 , n1290 );
buf ( RI15b46f68_286 , n1291 );
buf ( RI15b461d0_257 , n1292 );
buf ( RI15b472b0_293 , n1293 );
buf ( RI15b5f928_1126 , n1294 );
buf ( RI15b5f1a8_1110 , n1235 );
buf ( RI15b536a0_711 , n1295 );
buf ( RI15b45b40_243 , n1296 );
buf ( RI15b48138_324 , n1297 );
buf ( RI15b5f400_1115 , n1298 );
buf ( RI15b46b30_277 , n1299 );
buf ( RI15b46608_266 , n1300 );
buf ( RI15b45690_233 , n1301 );
buf ( RI15b53790_713 , n1302 );
buf ( RI15b5fbf8_1132 , n1303 );
buf ( RI15b54078_732 , n1304 );
buf ( RI15b46e78_284 , n1280 );
buf ( RI15b46c98_280 , n1305 );
buf ( RI15b53e98_728 , n1306 );
buf ( RI15b455a0_231 , n1307 );
buf ( RI15b47940_307 , n1308 );
buf ( RI15b45e10_249 , n1309 );
buf ( RI15b5fa90_1129 , n1310 );
buf ( RI15b5f310_1113 , n1190 );
buf ( RI15b54348_738 , n1311 );
buf ( RI15b60a08_1162 , n1312 );
buf ( RI15b60210_1145 , n1314 );
buf ( RI15b478c8_306 , n1315 );
buf ( RI15b47c88_314 , n1316 );
buf ( RI15b46680_267 , n1317 );
buf ( RI15b46158_256 , n1318 );
buf ( RI15b5fc70_1133 , n1319 );
buf ( RI15b53a60_719 , n1320 );
buf ( RI15b532e0_703 , n1058 );
buf ( RI15b538f8_716 , n1321 );
buf ( RI15b5eb18_1096 , n1322 );
buf ( RI15b52728_678 , n1324 );
buf ( RI15b600a8_1142 , n1326 );
buf ( RI15b5eaa0_1095 , n1325 );
buf ( RI15b5ede8_1102 , n1327 );
buf ( RI15b5f040_1107 , n1323 );
buf ( RI15b5eb90_1097 , n1328 );
buf ( RI15b60198_1144 , n1329 );
buf ( RI15b481b0_325 , n1330 );
buf ( RI15b545a0_743 , n1331 );
buf ( RI15b452d0_225 , n1332 );
buf ( RI15b46d88_282 , n1333 );
buf ( RI15b5ea28_1094 , n1334 );
buf ( RI15b54438_740 , n1335 );
buf ( RI15b47508_298 , n1336 );
buf ( RI15b466f8_268 , n1337 );
buf ( RI15b53178_700 , n1249 );
buf ( RI15b47148_290 , n1338 );
buf ( RI15b469c8_274 , n1173 );
buf ( RI15b458e8_238 , n1339 );
buf ( RI15b448f8_204 , n1185 );
buf ( RI15b52a70_685 , n1340 );
buf ( RI15b52818_680 , n1341 );
buf ( RI15b5ffb8_1140 , n1343 );
buf ( RI15b5e9b0_1093 , n1342 );
buf ( RI15b5f8b0_1125 , n1344 );
buf ( RI15b531f0_701 , n1313 );
buf ( RI15b46ef0_285 , n1345 );
buf ( RI15b45ca8_246 , n1346 );
buf ( RI15b52bd8_688 , n1116 );
buf ( RI15b53970_717 , n1347 );
buf ( RI15b52db8_692 , n1197 );
buf ( RI15b47580_299 , n1348 );
buf ( RI15b5e938_1092 , n1350 );
buf ( RI15b45078_220 , n1351 );
buf ( RI15b60300_1147 , n1352 );
buf ( RI15b60a80_1163 , n1354 );
buf ( RI15b5f478_1116 , n1217 );
buf ( RI15b473a0_295 , n1355 );
buf ( RI15b47760_303 , n1356 );
buf ( RI15b5fec8_1138 , n1358 );
buf ( RI15b5f748_1122 , n1357 );
buf ( RI15b45c30_245 , n1359 );
buf ( RI15b46770_269 , n1353 );
buf ( RI15b53010_697 , n1349 );
buf ( RI15b53d30_725 , n1360 );
buf ( RI15b52d40_691 , n1140 );
buf ( RI15b45708_234 , n1361 );
buf ( RI15b54528_742 , n1362 );
buf ( RI15b459d8_240 , n1363 );
buf ( n1364 , R_187c_13cca558 );
buf ( n1365 , R_125d_156aaaf8 );
buf ( n1366 , R_c3e_13d2c178 );
buf ( n1367 , R_61f_117eb278 );
buf ( n1368 , R_187d_117f5b38 );
buf ( n1369 , R_125e_13b8fe18 );
buf ( n1370 , R_c3f_123b4358 );
buf ( n1371 , R_187b_13ccb278 );
buf ( n1372 , R_620_13dfb518 );
buf ( n1373 , R_125c_15816b78 );
buf ( n1374 , R_c3d_13c22918 );
buf ( n1375 , R_61e_14a0c538 );
buf ( n1376 , R_5e7_10080958 );
buf ( n1377 , R_c06_170189e8 );
buf ( n1378 , R_18b4_1162f978 );
buf ( n1379 , R_1225_13c08298 );
buf ( n1380 , R_1844_117ef378 );
buf ( n1381 , R_1295_123bcf58 );
buf ( n1382 , R_c76_15ff42e8 );
buf ( n1383 , R_657_13bf5c78 );
buf ( n1384 , R_187e_140ac0d8 );
buf ( n1385 , R_125f_13c0f638 );
buf ( n1386 , R_c40_1580a9b8 );
buf ( n1387 , R_621_11c70318 );
buf ( n1388 , R_187a_13ddd2d8 );
buf ( n1389 , R_61d_123b84f8 );
buf ( n1390 , R_125b_1162bf58 );
buf ( n1391 , R_c3c_15ff9928 );
buf ( n1392 , R_12be_13ccf378 );
buf ( n1393 , R_5be_11c6a738 );
buf ( n1394 , R_bdd_17016508 );
buf ( n1395 , R_c9f_11636598 );
buf ( n1396 , R_11fc_13ddf7b8 );
buf ( n1397 , R_680_10085638 );
buf ( n1398 , R_181b_13d430d8 );
buf ( n1399 , R_18dd_13c062b8 );
buf ( n1400 , R_180c_156b4eb8 );
buf ( n1401 , R_12cd_13d535d8 );
buf ( n1402 , R_5af_1700c3c8 );
buf ( n1403 , R_cae_14a14ff8 );
buf ( n1404 , R_bce_15ff4608 );
buf ( n1405 , R_68f_13befcd8 );
buf ( n1406 , R_18ec_13d204b8 );
buf ( n1407 , R_11ed_116361d8 );
buf ( n1408 , R_187f_15811038 );
buf ( n1409 , R_1260_13d3b6f8 );
buf ( n1410 , R_c41_14a0bef8 );
buf ( n1411 , R_622_123b3bd8 );
buf ( n1412 , R_61c_13d56378 );
buf ( n1413 , R_c3b_150e7c58 );
buf ( n1414 , R_1879_15ff5c88 );
buf ( n1415 , R_125a_13bf58b8 );
buf ( n1416 , R_f82_13c1cd38 );
buf ( n1417 , R_963_13c209d8 );
buf ( n1418 , R_8fa_117ec678 );
buf ( n1419 , R_f19_15ff0648 );
buf ( n1420 , R_1538_13d29bf8 );
buf ( n1421 , R_15a1_150e22f8 );
buf ( n1422 , R_158f_13cd9058 );
buf ( n1423 , R_f70_17015608 );
buf ( n1424 , R_951_156b2578 );
buf ( n1425 , R_90c_13c0e0f8 );
buf ( n1426 , R_f2b_140b8838 );
buf ( n1427 , R_154a_1587f278 );
buf ( n1428 , R_1880_13c22738 );
buf ( n1429 , R_1261_13ccc0d8 );
buf ( n1430 , R_c42_117eb818 );
buf ( n1431 , R_623_140b3158 );
buf ( n1432 , R_61b_11c70458 );
buf ( n1433 , R_c3a_13b96218 );
buf ( n1434 , R_1259_13d23578 );
buf ( n1435 , R_1878_1162da38 );
buf ( n1436 , R_ce6_14875d78 );
buf ( n1437 , R_1924_13d1df38 );
buf ( n1438 , R_11b5_13d56f58 );
buf ( n1439 , R_577_1162c818 );
buf ( n1440 , R_6c7_10082438 );
buf ( n1441 , R_17d4_13cda278 );
buf ( n1442 , R_1305_10081fd8 );
buf ( n1443 , R_b96_15812b18 );
buf ( n1444 , R_1881_156b0638 );
buf ( n1445 , R_1262_12fc1698 );
buf ( n1446 , R_c43_140b0138 );
buf ( n1447 , R_624_13d421d8 );
buf ( n1448 , R_61a_14b2a318 );
buf ( n1449 , R_c39_117eaeb8 );
buf ( n1450 , R_1258_117e8618 );
buf ( n1451 , R_1877_1162cdb8 );
buf ( n1452 , R_119b_15ffa3c8 );
buf ( n1453 , R_55d_13b8e5b8 );
buf ( n1454 , R_131f_158106d8 );
buf ( n1455 , R_6e1_13c0fb38 );
buf ( n1456 , R_17ba_15fed6c8 );
buf ( n1457 , R_b7c_13b96e98 );
buf ( n1458 , R_193e_123b6018 );
buf ( n1459 , R_d00_117ec358 );
buf ( n1460 , R_1323_13d5b878 );
buf ( n1461 , R_6e5_15ff5328 );
buf ( n1462 , R_559_13c024d8 );
buf ( n1463 , R_1197_13bf4918 );
buf ( n1464 , R_1942_11c6dd98 );
buf ( n1465 , R_d04_14a16df8 );
buf ( n1466 , R_17b6_13dec158 );
buf ( n1467 , R_b78_13c10c18 );
buf ( n1468 , R_13ca_13d2c718 );
buf ( n1469 , R_19e9_13bf62b8 );
buf ( n1470 , R_170f_150defb8 );
buf ( n1471 , R_10f0_140b1ad8 );
buf ( n1472 , R_ad1_11c6ac38 );
buf ( n1473 , R_78c_13d5d3f8 );
buf ( n1474 , R_dab_140b3dd8 );
buf ( n1475 , R_883_13b936f8 );
buf ( n1476 , R_ff9_11631958 );
buf ( n1477 , R_ea2_150dd758 );
buf ( n1478 , R_9da_13cd8018 );
buf ( n1479 , R_1618_117f3658 );
buf ( n1480 , R_14c1_123ba4d8 );
buf ( n1481 , R_b5e_14a0f918 );
buf ( n1482 , R_179c_123bb018 );
buf ( n1483 , R_133d_13cd4e18 );
buf ( n1484 , R_6ff_14a0a918 );
buf ( n1485 , R_195c_150ddf78 );
buf ( n1486 , R_117d_123b8c78 );
buf ( n1487 , R_d1e_124c2cd8 );
buf ( n1488 , R_5f7_12fbf758 );
buf ( n1489 , R_c16_13df9858 );
buf ( n1490 , R_1235_15880cb8 );
buf ( n1491 , R_1854_1580fd78 );
buf ( n1492 , R_18a4_13bf2d98 );
buf ( n1493 , R_1285_100890f8 );
buf ( n1494 , R_c66_13bed2f8 );
buf ( n1495 , R_647_13d51af8 );
buf ( n1496 , R_1882_13d1fbf8 );
buf ( n1497 , R_1263_123be498 );
buf ( n1498 , R_c44_13c229b8 );
buf ( n1499 , R_625_13c1e638 );
buf ( n1500 , R_619_156b6718 );
buf ( n1501 , R_c38_117efd78 );
buf ( n1502 , R_1257_14a0f0f8 );
buf ( n1503 , R_1876_15ffcb28 );
buf ( n1504 , R_985_1587c4d8 );
buf ( n1505 , R_1516_12fc1eb8 );
buf ( n1506 , R_15c3_13c02078 );
buf ( n1507 , R_8d8_13d22fd8 );
buf ( n1508 , R_fa4_13d1e898 );
buf ( n1509 , R_ef7_1162bd78 );
buf ( n1510 , R_1663_124c2698 );
buf ( n1511 , R_838_1580b8b8 );
buf ( n1512 , R_a25_13bf4ff8 );
buf ( n1513 , R_1476_1486bd78 );
buf ( n1514 , R_1044_13d57818 );
buf ( n1515 , R_e57_13b8f738 );
buf ( n1516 , R_15fa_13c0bb78 );
buf ( n1517 , R_ec0_13c1bf78 );
buf ( n1518 , R_fdb_15ff7308 );
buf ( n1519 , R_14df_14a0cdf8 );
buf ( n1520 , R_9bc_15812758 );
buf ( n1521 , R_8a1_13d21818 );
buf ( n1522 , R_1883_13d41058 );
buf ( n1523 , R_1264_13c02758 );
buf ( n1524 , R_c45_13d24c98 );
buf ( n1525 , R_626_123b86d8 );
buf ( n1526 , R_618_1587ea58 );
buf ( n1527 , R_c37_13c0bfd8 );
buf ( n1528 , R_1256_13d54258 );
buf ( n1529 , R_1875_158179d8 );
buf ( n1530 , R_1145_13b98658 );
buf ( n1531 , R_737_116313b8 );
buf ( n1532 , R_b26_1486a518 );
buf ( n1533 , R_d56_117e9d38 );
buf ( n1534 , R_1764_13ccf7d8 );
buf ( n1535 , R_1375_13c275f8 );
buf ( n1536 , R_1994_123bac58 );
buf ( n1537 , R_143d_13bf2258 );
buf ( n1538 , R_a5e_1587ed78 );
buf ( n1539 , R_e1e_13c1bbb8 );
buf ( n1540 , R_107d_15888418 );
buf ( n1541 , R_7ff_13cd45f8 );
buf ( n1542 , R_169c_15885fd8 );
buf ( n1543 , R_1a5c_13de04d8 );
buf ( n1544 , R_1a48_13c1ff38 );
buf ( n1545 , R_a72_1486d358 );
buf ( n1546 , R_1429_13d23438 );
buf ( n1547 , R_1091_14a11d58 );
buf ( n1548 , R_e0a_13bfa3b8 );
buf ( n1549 , R_16b0_140aae18 );
buf ( n1550 , R_7eb_123b8278 );
buf ( n1551 , R_12c6_13cd49b8 );
buf ( n1552 , R_5b6_117f1f38 );
buf ( n1553 , R_ca7_140b4418 );
buf ( n1554 , R_bd5_13d51698 );
buf ( n1555 , R_688_13b99af8 );
buf ( n1556 , R_11f4_13d1e6b8 );
buf ( n1557 , R_18e5_13d45658 );
buf ( n1558 , R_1813_13d29c98 );
buf ( n1559 , R_16d9_14a17cf8 );
buf ( n1560 , R_1a1f_11c70958 );
buf ( n1561 , R_1400_14b29b98 );
buf ( n1562 , R_de1_13cd0638 );
buf ( n1563 , R_7c2_15ffa508 );
buf ( n1564 , R_a9b_100865d8 );
buf ( n1565 , R_10ba_15881938 );
buf ( n1566 , R_1805_14b271b8 );
buf ( n1567 , R_5a8_123b8318 );
buf ( n1568 , R_cb5_170107e8 );
buf ( n1569 , R_bc7_13c2a758 );
buf ( n1570 , R_696_10082ed8 );
buf ( n1571 , R_18f3_15ffc628 );
buf ( n1572 , R_11e6_14b222f8 );
buf ( n1573 , R_12d4_11634d38 );
buf ( n1574 , R_119f_156b4738 );
buf ( n1575 , R_561_1162a658 );
buf ( n1576 , R_6dd_117f36f8 );
buf ( n1577 , R_131b_15ff76c8 );
buf ( n1578 , R_17be_15816538 );
buf ( n1579 , R_b80_13cd8338 );
buf ( n1580 , R_cfc_1700d2c8 );
buf ( n1581 , R_193a_15885718 );
buf ( n1582 , R_5da_13df70f8 );
buf ( n1583 , R_18c1_11c6f738 );
buf ( n1584 , R_bf9_13d28ed8 );
buf ( n1585 , R_12a2_13bf2578 );
buf ( n1586 , R_1218_13d28078 );
buf ( n1587 , R_c83_13d59f78 );
buf ( n1588 , R_1837_13deb9d8 );
buf ( n1589 , R_664_123b47b8 );
buf ( n1590 , R_e39_156b3518 );
buf ( n1591 , R_a43_14b1feb8 );
buf ( n1592 , R_81a_13cceb58 );
buf ( n1593 , R_1062_117eedd8 );
buf ( n1594 , R_1458_13df07f8 );
buf ( n1595 , R_1681_140b99b8 );
buf ( n1596 , R_1327_124c2b98 );
buf ( n1597 , R_6e9_156b3158 );
buf ( n1598 , R_555_13d59b18 );
buf ( n1599 , R_1193_13b97438 );
buf ( n1600 , R_1946_14a16858 );
buf ( n1601 , R_d08_13d59938 );
buf ( n1602 , R_b74_123c0478 );
buf ( n1603 , R_17b2_13cd6498 );
buf ( n1604 , R_113a_117eb458 );
buf ( n1605 , R_742_14a129d8 );
buf ( n1606 , R_b1b_11629758 );
buf ( n1607 , R_d61_11633618 );
buf ( n1608 , R_1380_15887338 );
buf ( n1609 , R_1759_14874518 );
buf ( n1610 , R_199f_13d3c9b8 );
buf ( n1611 , R_1884_13cd1c18 );
buf ( n1612 , R_1265_156b0818 );
buf ( n1613 , R_c46_1580b598 );
buf ( n1614 , R_627_117efb98 );
buf ( n1615 , R_617_158807b8 );
buf ( n1616 , R_c36_156b63f8 );
buf ( n1617 , R_1255_1580dbb8 );
buf ( n1618 , R_1874_13df9c18 );
buf ( n1619 , R_87a_13c286d8 );
buf ( n1620 , R_1002_14a17938 );
buf ( n1621 , R_e99_123ba258 );
buf ( n1622 , R_9e3_170110a8 );
buf ( n1623 , R_1621_117eacd8 );
buf ( n1624 , R_14b8_123b31d8 );
buf ( n1625 , R_edf_117f5bd8 );
buf ( n1626 , R_14fe_13d55518 );
buf ( n1627 , R_15db_117f7258 );
buf ( n1628 , R_fbc_13beb9f8 );
buf ( n1629 , R_8c0_11631ef8 );
buf ( n1630 , R_99d_13cd4d78 );
buf ( n1631 , R_845_15888918 );
buf ( n1632 , R_1656_117f4af8 );
buf ( n1633 , R_1483_13d53d58 );
buf ( n1634 , R_a18_12fbdef8 );
buf ( n1635 , R_e64_14875058 );
buf ( n1636 , R_1037_15815098 );
buf ( n1637 , R_d8e_11630878 );
buf ( n1638 , R_172c_13d39d58 );
buf ( n1639 , R_13ad_14a12618 );
buf ( n1640 , R_19cc_13cda1d8 );
buf ( n1641 , R_110d_13dd5cb8 );
buf ( n1642 , R_aee_117e9478 );
buf ( n1643 , R_76f_117f4378 );
buf ( n1644 , R_ccd_13b8c8f8 );
buf ( n1645 , R_590_13dd64d8 );
buf ( n1646 , R_17ed_156b36f8 );
buf ( n1647 , R_190b_14872038 );
buf ( n1648 , R_6ae_156ab958 );
buf ( n1649 , R_baf_1700cd28 );
buf ( n1650 , R_12ec_124c3778 );
buf ( n1651 , R_11ce_11c6cad8 );
buf ( n1652 , R_17a3_150e7398 );
buf ( n1653 , R_1336_148754b8 );
buf ( n1654 , R_6f8_13c1c018 );
buf ( n1655 , R_1184_150e6498 );
buf ( n1656 , R_1955_14b235b8 );
buf ( n1657 , R_d17_14b27398 );
buf ( n1658 , R_b65_13dde318 );
buf ( n1659 , R_1885_1486cdb8 );
buf ( n1660 , R_1266_14a12438 );
buf ( n1661 , R_c47_100803b8 );
buf ( n1662 , R_628_117eb098 );
buf ( n1663 , R_616_170152e8 );
buf ( n1664 , R_c35_123b88b8 );
buf ( n1665 , R_1254_150e59f8 );
buf ( n1666 , R_1873_12fc2278 );
buf ( n1667 , R_74a_1008cb18 );
buf ( n1668 , R_1132_15880e98 );
buf ( n1669 , R_d69_14b23158 );
buf ( n1670 , R_b13_140b3d38 );
buf ( n1671 , R_1388_140aaf58 );
buf ( n1672 , R_19a7_140b9b98 );
buf ( n1673 , R_1751_1007feb8 );
buf ( n1674 , R_b57_13ccd6b8 );
buf ( n1675 , R_1344_117f3018 );
buf ( n1676 , R_1795_1008b678 );
buf ( n1677 , R_706_1580bd18 );
buf ( n1678 , R_1963_13d1f478 );
buf ( n1679 , R_1176_17015b08 );
buf ( n1680 , R_d25_15882298 );
buf ( n1681 , R_1590_150e4b98 );
buf ( n1682 , R_f71_124c4998 );
buf ( n1683 , R_952_14b26e98 );
buf ( n1684 , R_90b_13d41af8 );
buf ( n1685 , R_f2a_1162a158 );
buf ( n1686 , R_1549_1587ff98 );
buf ( n1687 , R_5c6_15816218 );
buf ( n1688 , R_12b6_1587db58 );
buf ( n1689 , R_be5_140b5818 );
buf ( n1690 , R_c97_156b09f8 );
buf ( n1691 , R_1204_13c23b38 );
buf ( n1692 , R_678_15884ef8 );
buf ( n1693 , R_1823_13d53df8 );
buf ( n1694 , R_18d5_11636098 );
buf ( n1695 , R_ed8_117e9c98 );
buf ( n1696 , R_15e2_14a140f8 );
buf ( n1697 , R_14f7_13b965d8 );
buf ( n1698 , R_fc3_14b27e38 );
buf ( n1699 , R_8b9_14875e18 );
buf ( n1700 , R_9a4_117ee018 );
buf ( n1701 , R_1a04_13c22b98 );
buf ( n1702 , R_13e5_13de07f8 );
buf ( n1703 , R_16f4_123b9fd8 );
buf ( n1704 , R_dc6_14873f78 );
buf ( n1705 , R_10d5_13b94a58 );
buf ( n1706 , R_7a7_116355f8 );
buf ( n1707 , R_ab6_15814e18 );
buf ( n1708 , R_1886_11638c58 );
buf ( n1709 , R_1267_14b23f18 );
buf ( n1710 , R_c48_13bf5e58 );
buf ( n1711 , R_629_150e7e38 );
buf ( n1712 , R_615_13c1d7d8 );
buf ( n1713 , R_c34_15ff1228 );
buf ( n1714 , R_1253_13d222b8 );
buf ( n1715 , R_1872_13ccb4f8 );
buf ( n1716 , R_16f6_116389d8 );
buf ( n1717 , R_10d7_156b5778 );
buf ( n1718 , R_ab8_156ac8f8 );
buf ( n1719 , R_1a02_13cd8298 );
buf ( n1720 , R_13e3_14a0a7d8 );
buf ( n1721 , R_7a5_13d456f8 );
buf ( n1722 , R_dc4_11634b58 );
buf ( n1723 , R_b4d_1700f208 );
buf ( n1724 , R_710_156ac718 );
buf ( n1725 , R_178b_1580ca38 );
buf ( n1726 , R_196d_117eb8b8 );
buf ( n1727 , R_d2f_13dedf58 );
buf ( n1728 , R_116c_140b8338 );
buf ( n1729 , R_134e_13d282f8 );
buf ( n1730 , R_1a06_1486e1b8 );
buf ( n1731 , R_13e7_116377b8 );
buf ( n1732 , R_dc8_1162b058 );
buf ( n1733 , R_7a9_123bd458 );
buf ( n1734 , R_16f2_158857b8 );
buf ( n1735 , R_ab4_12fbed58 );
buf ( n1736 , R_10d3_158899f8 );
buf ( n1737 , R_85a_156b1a38 );
buf ( n1738 , R_1498_15811c18 );
buf ( n1739 , R_1641_150db8b8 );
buf ( n1740 , R_a03_123bd818 );
buf ( n1741 , R_e79_13cd8658 );
buf ( n1742 , R_1022_11c6cf38 );
buf ( n1743 , R_150d_14b21678 );
buf ( n1744 , R_15cc_14a0ba98 );
buf ( n1745 , R_8cf_13ded9b8 );
buf ( n1746 , R_fad_140ac038 );
buf ( n1747 , R_eee_11632e98 );
buf ( n1748 , R_98e_12fbecb8 );
buf ( n1749 , R_13bd_13df6c98 );
buf ( n1750 , R_19dc_156b6858 );
buf ( n1751 , R_171c_117ecb78 );
buf ( n1752 , R_10fd_117eef18 );
buf ( n1753 , R_ade_13dd7658 );
buf ( n1754 , R_77f_117f4558 );
buf ( n1755 , R_d9e_13ddc3d8 );
buf ( n1756 , R_16f8_14a0e018 );
buf ( n1757 , R_10d9_123b9538 );
buf ( n1758 , R_aba_13c29678 );
buf ( n1759 , R_7a3_13ccb138 );
buf ( n1760 , R_dc2_158108b8 );
buf ( n1761 , R_13e1_156b8478 );
buf ( n1762 , R_1a00_123b7f58 );
buf ( n1763 , R_971_13df5618 );
buf ( n1764 , R_8ec_123bbd38 );
buf ( n1765 , R_15af_14866eb8 );
buf ( n1766 , R_f0b_13cd72f8 );
buf ( n1767 , R_f90_15812438 );
buf ( n1768 , R_152a_13df8818 );
buf ( n1769 , R_c15_15fee528 );
buf ( n1770 , R_1234_15ff9e28 );
buf ( n1771 , R_1853_13dd8738 );
buf ( n1772 , R_18a5_170177c8 );
buf ( n1773 , R_1286_124c4858 );
buf ( n1774 , R_c67_13ccba98 );
buf ( n1775 , R_648_15814058 );
buf ( n1776 , R_5f6_13cce018 );
buf ( n1777 , R_c05_14866d78 );
buf ( n1778 , R_18b5_10087cf8 );
buf ( n1779 , R_1224_13ccff58 );
buf ( n1780 , R_1296_13dda7b8 );
buf ( n1781 , R_1843_1580a878 );
buf ( n1782 , R_c77_13d523b8 );
buf ( n1783 , R_658_140ae1f8 );
buf ( n1784 , R_5e6_13d46698 );
buf ( n1785 , R_1a08_14b1b958 );
buf ( n1786 , R_13e9_13d22358 );
buf ( n1787 , R_dca_14b297d8 );
buf ( n1788 , R_7ab_15887ab8 );
buf ( n1789 , R_ab2_13df75f8 );
buf ( n1790 , R_10d1_13d55d38 );
buf ( n1791 , R_16f0_14b1e978 );
buf ( n1792 , R_d87_123bae38 );
buf ( n1793 , R_1733_15ff79e8 );
buf ( n1794 , R_13a6_156b1718 );
buf ( n1795 , R_1114_13d46ff8 );
buf ( n1796 , R_19c5_13bf6ad8 );
buf ( n1797 , R_af5_13c1b6b8 );
buf ( n1798 , R_768_158896d8 );
buf ( n1799 , R_964_123c1f58 );
buf ( n1800 , R_8f9_117ee658 );
buf ( n1801 , R_f18_14a19d78 );
buf ( n1802 , R_1537_117e9b58 );
buf ( n1803 , R_15a2_13ccce98 );
buf ( n1804 , R_f83_14a0e978 );
buf ( n1805 , R_1887_17018da8 );
buf ( n1806 , R_1268_13d38278 );
buf ( n1807 , R_c49_123b36d8 );
buf ( n1808 , R_62a_13d42278 );
buf ( n1809 , R_614_13c2a258 );
buf ( n1810 , R_c33_150e7bb8 );
buf ( n1811 , R_1252_116378f8 );
buf ( n1812 , R_1871_13defad8 );
buf ( n1813 , R_11a3_13c1be38 );
buf ( n1814 , R_565_13ddbb18 );
buf ( n1815 , R_6d9_11636818 );
buf ( n1816 , R_1317_1580c5d8 );
buf ( n1817 , R_17c2_13c03518 );
buf ( n1818 , R_b84_156b5278 );
buf ( n1819 , R_cf8_15881a78 );
buf ( n1820 , R_1936_13d2a558 );
buf ( n1821 , R_13b4_156abb38 );
buf ( n1822 , R_19d3_13bf92d8 );
buf ( n1823 , R_1725_13cd9a58 );
buf ( n1824 , R_1106_14b1c718 );
buf ( n1825 , R_ae7_13cd22f8 );
buf ( n1826 , R_776_14873bb8 );
buf ( n1827 , R_d95_15815778 );
buf ( n1828 , R_feb_1486c818 );
buf ( n1829 , R_eb0_13d53498 );
buf ( n1830 , R_14cf_14b1bd18 );
buf ( n1831 , R_9cc_158172f8 );
buf ( n1832 , R_160a_17010ce8 );
buf ( n1833 , R_891_13b8ab98 );
buf ( n1834 , R_132b_1007f7d8 );
buf ( n1835 , R_6ed_140b6538 );
buf ( n1836 , R_118f_14b1ee78 );
buf ( n1837 , R_194a_13d2ae18 );
buf ( n1838 , R_d0c_13dee8b8 );
buf ( n1839 , R_b70_13d20f58 );
buf ( n1840 , R_17ae_13d29a18 );
buf ( n1841 , R_1a3c_13b95278 );
buf ( n1842 , R_109d_10084878 );
buf ( n1843 , R_141d_13d441b8 );
buf ( n1844 , R_16bc_14a0bdb8 );
buf ( n1845 , R_dfe_15ff38e8 );
buf ( n1846 , R_7df_1587d338 );
buf ( n1847 , R_a7e_14a0bb38 );
buf ( n1848 , R_151f_12fbe998 );
buf ( n1849 , R_97c_13d528b8 );
buf ( n1850 , R_15ba_1008b0d8 );
buf ( n1851 , R_8e1_15889818 );
buf ( n1852 , R_f00_17017ae8 );
buf ( n1853 , R_f9b_13b974d8 );
buf ( n1854 , R_16fa_14b299b8 );
buf ( n1855 , R_10db_13cd6cb8 );
buf ( n1856 , R_abc_15882b58 );
buf ( n1857 , R_7a1_15ffcd08 );
buf ( n1858 , R_dc0_117f53b8 );
buf ( n1859 , R_13df_156b9238 );
buf ( n1860 , R_19fe_13c01fd8 );
buf ( n1861 , R_5cf_124c4678 );
buf ( n1862 , R_12ad_13cca878 );
buf ( n1863 , R_bee_156ac498 );
buf ( n1864 , R_c8e_156b6cb8 );
buf ( n1865 , R_120d_123be218 );
buf ( n1866 , R_66f_13df8d18 );
buf ( n1867 , R_182c_13b90598 );
buf ( n1868 , R_18cc_170190c8 );
buf ( n1869 , R_1505_13d27858 );
buf ( n1870 , R_15d4_13d3a078 );
buf ( n1871 , R_fb5_13c265b8 );
buf ( n1872 , R_8c7_13ccf738 );
buf ( n1873 , R_996_13cd1498 );
buf ( n1874 , R_ee6_156ae158 );
buf ( n1875 , R_1a0a_140b9238 );
buf ( n1876 , R_13eb_150e7438 );
buf ( n1877 , R_dcc_15815c78 );
buf ( n1878 , R_7ad_1008c078 );
buf ( n1879 , R_ab0_11629618 );
buf ( n1880 , R_10cf_1580df78 );
buf ( n1881 , R_16ee_123bf758 );
buf ( n1882 , R_1660_13dd6258 );
buf ( n1883 , R_83b_117f03b8 );
buf ( n1884 , R_a22_156b92d8 );
buf ( n1885 , R_1479_13ddc518 );
buf ( n1886 , R_1041_14a0db18 );
buf ( n1887 , R_e5a_11633118 );
buf ( n1888 , R_1711_11c69d38 );
buf ( n1889 , R_10f2_1486ad38 );
buf ( n1890 , R_ad3_13d5a5b8 );
buf ( n1891 , R_78a_13dfa2f8 );
buf ( n1892 , R_da9_123bc9b8 );
buf ( n1893 , R_13c8_11628e98 );
buf ( n1894 , R_19e7_14a10098 );
buf ( n1895 , R_eb5_13cd9cd8 );
buf ( n1896 , R_fe6_13df1d38 );
buf ( n1897 , R_14d4_13c27a58 );
buf ( n1898 , R_9c7_140af5f8 );
buf ( n1899 , R_896_123b6658 );
buf ( n1900 , R_1605_156b1b78 );
buf ( n1901 , R_1888_1580c858 );
buf ( n1902 , R_1269_13b99c38 );
buf ( n1903 , R_c4a_14a0cb78 );
buf ( n1904 , R_62b_1162a1f8 );
buf ( n1905 , R_613_124c47b8 );
buf ( n1906 , R_c32_14b23518 );
buf ( n1907 , R_1251_13d3fed8 );
buf ( n1908 , R_1870_13b92bb8 );
buf ( n1909 , R_16cc_156ba318 );
buf ( n1910 , R_1a2c_156b08b8 );
buf ( n1911 , R_140d_11638258 );
buf ( n1912 , R_dee_13c0e058 );
buf ( n1913 , R_7cf_123bbe78 );
buf ( n1914 , R_a8e_170160a8 );
buf ( n1915 , R_10ad_10082618 );
buf ( n1916 , R_11b0_13b99f58 );
buf ( n1917 , R_572_140ab458 );
buf ( n1918 , R_6cc_117e8a78 );
buf ( n1919 , R_130a_13dda498 );
buf ( n1920 , R_17cf_13d389f8 );
buf ( n1921 , R_b91_14b1f418 );
buf ( n1922 , R_ceb_13d56d78 );
buf ( n1923 , R_1929_13cd4af8 );
buf ( n1924 , R_f72_13c2a1b8 );
buf ( n1925 , R_953_14b20a98 );
buf ( n1926 , R_90a_156ae658 );
buf ( n1927 , R_f29_11630698 );
buf ( n1928 , R_1548_140ac538 );
buf ( n1929 , R_1591_13c25618 );
buf ( n1930 , R_16fc_156b9a58 );
buf ( n1931 , R_10dd_13d551f8 );
buf ( n1932 , R_abe_14a15958 );
buf ( n1933 , R_79f_140af7d8 );
buf ( n1934 , R_dbe_13cd4c38 );
buf ( n1935 , R_13dd_15884b38 );
buf ( n1936 , R_19fc_13b96fd8 );
buf ( n1937 , R_ff0_123b3b38 );
buf ( n1938 , R_eab_11634518 );
buf ( n1939 , R_9d1_13d4ed58 );
buf ( n1940 , R_14ca_11631e58 );
buf ( n1941 , R_160f_170102e8 );
buf ( n1942 , R_88c_116319f8 );
buf ( n1943 , R_e36_13c05b38 );
buf ( n1944 , R_a46_11637e98 );
buf ( n1945 , R_817_116294d8 );
buf ( n1946 , R_1065_13c0b218 );
buf ( n1947 , R_1455_117ef238 );
buf ( n1948 , R_1684_13dd5ad8 );
buf ( n1949 , R_e2b_13d28578 );
buf ( n1950 , R_a51_11630ff8 );
buf ( n1951 , R_80c_13d2acd8 );
buf ( n1952 , R_1070_150e2d98 );
buf ( n1953 , R_1a69_11c6fe18 );
buf ( n1954 , R_168f_13d295b8 );
buf ( n1955 , R_144a_1580c678 );
buf ( n1956 , R_1a0c_13ccacd8 );
buf ( n1957 , R_13ed_13cd4ff8 );
buf ( n1958 , R_dce_14871f98 );
buf ( n1959 , R_7af_11633578 );
buf ( n1960 , R_aae_15814238 );
buf ( n1961 , R_10cd_13d20878 );
buf ( n1962 , R_16ec_13df6a18 );
buf ( n1963 , R_1889_13bf9c38 );
buf ( n1964 , R_126a_15886a78 );
buf ( n1965 , R_c4b_13cd76b8 );
buf ( n1966 , R_62c_10086038 );
buf ( n1967 , R_612_10088dd8 );
buf ( n1968 , R_c31_13b90778 );
buf ( n1969 , R_1250_13d58c18 );
buf ( n1970 , R_186f_1162dcb8 );
buf ( n1971 , R_1a21_150e5598 );
buf ( n1972 , R_1402_140b1cb8 );
buf ( n1973 , R_de3_140b0778 );
buf ( n1974 , R_7c4_13cd5138 );
buf ( n1975 , R_a99_13cd0a98 );
buf ( n1976 , R_10b8_13bea7d8 );
buf ( n1977 , R_16d7_15888a58 );
buf ( n1978 , R_b23_1587bc18 );
buf ( n1979 , R_d59_14868cb8 );
buf ( n1980 , R_1378_14b28158 );
buf ( n1981 , R_1761_11631f98 );
buf ( n1982 , R_1997_13d45158 );
buf ( n1983 , R_1142_117f06d8 );
buf ( n1984 , R_73a_13de1158 );
buf ( n1985 , R_1a35_1486d7b8 );
buf ( n1986 , R_16c3_13c01498 );
buf ( n1987 , R_1416_1162ee38 );
buf ( n1988 , R_df7_117f35b8 );
buf ( n1989 , R_7d8_156abc78 );
buf ( n1990 , R_a85_17014168 );
buf ( n1991 , R_10a4_1486b0f8 );
buf ( n1992 , R_a59_14a1a1d8 );
buf ( n1993 , R_e23_13df5f78 );
buf ( n1994 , R_1078_1580f558 );
buf ( n1995 , R_804_156b6f38 );
buf ( n1996 , R_1697_13d59d98 );
buf ( n1997 , R_1a61_14a195f8 );
buf ( n1998 , R_1442_14a18c98 );
buf ( n1999 , R_1096_13dd6f78 );
buf ( n2000 , R_1424_13b906d8 );
buf ( n2001 , R_16b5_13c045f8 );
buf ( n2002 , R_e05_140ad938 );
buf ( n2003 , R_7e6_1486dd58 );
buf ( n2004 , R_a77_100895f8 );
buf ( n2005 , R_1a43_170104c8 );
buf ( n2006 , R_15ef_15889318 );
buf ( n2007 , R_ecb_13df7198 );
buf ( n2008 , R_14ea_13cd2078 );
buf ( n2009 , R_fd0_13cd59f8 );
buf ( n2010 , R_8ac_15889278 );
buf ( n2011 , R_9b1_1008a3b8 );
buf ( n2012 , R_cc2_14a11218 );
buf ( n2013 , R_17f8_13c28d18 );
buf ( n2014 , R_59b_15812bb8 );
buf ( n2015 , R_1900_1486c318 );
buf ( n2016 , R_6a3_11c69658 );
buf ( n2017 , R_bba_13deb7f8 );
buf ( n2018 , R_12e1_123bbf18 );
buf ( n2019 , R_11d9_14a18518 );
buf ( n2020 , R_1125_124c3e58 );
buf ( n2021 , R_d76_156b6218 );
buf ( n2022 , R_b06_14b24af8 );
buf ( n2023 , R_1395_13c0d978 );
buf ( n2024 , R_19b4_14a10598 );
buf ( n2025 , R_1744_11c6e3d8 );
buf ( n2026 , R_757_13d3ceb8 );
buf ( n2027 , R_16fe_123b51b8 );
buf ( n2028 , R_10df_156b31f8 );
buf ( n2029 , R_ac0_123c19b8 );
buf ( n2030 , R_79d_13ddd698 );
buf ( n2031 , R_dbc_13d207d8 );
buf ( n2032 , R_13db_13d412d8 );
buf ( n2033 , R_19fa_140afeb8 );
buf ( n2034 , R_188a_14a0dd98 );
buf ( n2035 , R_126b_170193e8 );
buf ( n2036 , R_c4c_14874a18 );
buf ( n2037 , R_62d_123c23b8 );
buf ( n2038 , R_611_156aa558 );
buf ( n2039 , R_c30_13cd8158 );
buf ( n2040 , R_124f_13cd9418 );
buf ( n2041 , R_186e_1162cb38 );
buf ( n2042 , R_1233_13d5c318 );
buf ( n2043 , R_1852_11635698 );
buf ( n2044 , R_18a6_15885218 );
buf ( n2045 , R_1287_13c29e98 );
buf ( n2046 , R_c68_12fc1cd8 );
buf ( n2047 , R_649_150e1f38 );
buf ( n2048 , R_5f5_13bf7398 );
buf ( n2049 , R_c14_13defe98 );
buf ( n2050 , R_18c2_13d5d998 );
buf ( n2051 , R_bf8_13bf77f8 );
buf ( n2052 , R_12a3_14b20278 );
buf ( n2053 , R_1217_123bdd18 );
buf ( n2054 , R_c84_123bee98 );
buf ( n2055 , R_1836_14a16038 );
buf ( n2056 , R_665_117eefb8 );
buf ( n2057 , R_5d9_15fed588 );
buf ( n2058 , R_84f_1587bdf8 );
buf ( n2059 , R_148d_156b2d98 );
buf ( n2060 , R_164c_156b65d8 );
buf ( n2061 , R_a0e_13cd5098 );
buf ( n2062 , R_e6e_13c1e818 );
buf ( n2063 , R_102d_14a14878 );
buf ( n2064 , R_d7b_1007dbb8 );
buf ( n2065 , R_1120_13cd3158 );
buf ( n2066 , R_139a_12fbf398 );
buf ( n2067 , R_b01_1587af98 );
buf ( n2068 , R_19b9_116327b8 );
buf ( n2069 , R_75c_13d54b18 );
buf ( n2070 , R_173f_14a0d1b8 );
buf ( n2071 , R_ca0_117f3978 );
buf ( n2072 , R_bdc_14867a98 );
buf ( n2073 , R_11fb_13d26638 );
buf ( n2074 , R_681_13c02c58 );
buf ( n2075 , R_18de_1162c638 );
buf ( n2076 , R_181a_15887fb8 );
buf ( n2077 , R_12bf_12fbe3f8 );
buf ( n2078 , R_5bd_123b9678 );
buf ( n2079 , R_1a0e_1486b698 );
buf ( n2080 , R_13ef_156ba1d8 );
buf ( n2081 , R_dd0_12fc0798 );
buf ( n2082 , R_7b1_14a13478 );
buf ( n2083 , R_aac_116311d8 );
buf ( n2084 , R_10cb_150dccb8 );
buf ( n2085 , R_16ea_140b6cb8 );
buf ( n2086 , R_ffe_13ccf198 );
buf ( n2087 , R_e9d_13d27038 );
buf ( n2088 , R_9df_14a17398 );
buf ( n2089 , R_161d_13b962b8 );
buf ( n2090 , R_14bc_117f0598 );
buf ( n2091 , R_87e_140b08b8 );
buf ( n2092 , R_5a1_13d446b8 );
buf ( n2093 , R_cbc_12fc1b98 );
buf ( n2094 , R_bc0_13dfb338 );
buf ( n2095 , R_69d_11c69798 );
buf ( n2096 , R_18fa_140b5098 );
buf ( n2097 , R_11df_15880998 );
buf ( n2098 , R_12db_156b4af8 );
buf ( n2099 , R_17fe_1580f5f8 );
buf ( n2100 , R_191b_13c25f78 );
buf ( n2101 , R_580_1162b4b8 );
buf ( n2102 , R_6be_158101d8 );
buf ( n2103 , R_17dd_14872358 );
buf ( n2104 , R_12fc_15813dd8 );
buf ( n2105 , R_b9f_140b49b8 );
buf ( n2106 , R_cdd_13bf42d8 );
buf ( n2107 , R_11be_150e4378 );
buf ( n2108 , R_eba_13d29158 );
buf ( n2109 , R_fe1_13d2bef8 );
buf ( n2110 , R_14d9_13c21338 );
buf ( n2111 , R_9c2_116297f8 );
buf ( n2112 , R_89b_117ed118 );
buf ( n2113 , R_1600_117e96f8 );
buf ( n2114 , R_585_14a19b98 );
buf ( n2115 , R_1916_150e99b8 );
buf ( n2116 , R_17e2_123c1d78 );
buf ( n2117 , R_6b9_150dc998 );
buf ( n2118 , R_ba4_13c04d78 );
buf ( n2119 , R_12f7_117f4ff8 );
buf ( n2120 , R_11c3_117ee158 );
buf ( n2121 , R_cd8_150deab8 );
buf ( n2122 , R_15c4_13d46e18 );
buf ( n2123 , R_8d7_13de10b8 );
buf ( n2124 , R_fa5_13df4858 );
buf ( n2125 , R_ef6_13c1f358 );
buf ( n2126 , R_986_11631278 );
buf ( n2127 , R_1515_13ccb8b8 );
buf ( n2128 , R_11a7_123b9b78 );
buf ( n2129 , R_569_12fbfd98 );
buf ( n2130 , R_6d5_14b25958 );
buf ( n2131 , R_1313_1587dab8 );
buf ( n2132 , R_17c6_13d290b8 );
buf ( n2133 , R_b88_14a0d9d8 );
buf ( n2134 , R_cf4_13bea558 );
buf ( n2135 , R_1932_13cd1538 );
buf ( n2136 , R_1778_11631598 );
buf ( n2137 , R_d42_1580f918 );
buf ( n2138 , R_1159_148722b8 );
buf ( n2139 , R_1361_14a18658 );
buf ( n2140 , R_b3a_11637678 );
buf ( n2141 , R_1980_15883a58 );
buf ( n2142 , R_723_14a0aeb8 );
buf ( n2143 , R_ec5_123c1eb8 );
buf ( n2144 , R_fd6_15ff7448 );
buf ( n2145 , R_14e4_14a121b8 );
buf ( n2146 , R_9b7_117eaaf8 );
buf ( n2147 , R_8a6_156b3018 );
buf ( n2148 , R_15f5_140ade38 );
buf ( n2149 , R_d45_117f4418 );
buf ( n2150 , R_1775_140b5d18 );
buf ( n2151 , R_1364_13c1d918 );
buf ( n2152 , R_1156_15ff6fe8 );
buf ( n2153 , R_1983_100863f8 );
buf ( n2154 , R_726_13d39498 );
buf ( n2155 , R_b37_10089b98 );
buf ( n2156 , R_15e9_11636db8 );
buf ( n2157 , R_14f0_13b92398 );
buf ( n2158 , R_fca_156b44b8 );
buf ( n2159 , R_8b2_11629078 );
buf ( n2160 , R_9ab_14866698 );
buf ( n2161 , R_ed1_158870b8 );
buf ( n2162 , R_1632_117f1178 );
buf ( n2163 , R_9f4_1486d2b8 );
buf ( n2164 , R_e88_124c4498 );
buf ( n2165 , R_1013_14a135b8 );
buf ( n2166 , R_14a7_15814af8 );
buf ( n2167 , R_869_14a19e18 );
buf ( n2168 , R_132f_13c0b8f8 );
buf ( n2169 , R_6f1_150df878 );
buf ( n2170 , R_118b_14b27618 );
buf ( n2171 , R_194e_14b236f8 );
buf ( n2172 , R_d10_123b2d78 );
buf ( n2173 , R_b6c_123b8138 );
buf ( n2174 , R_17aa_13dfac58 );
buf ( n2175 , R_188b_117e9978 );
buf ( n2176 , R_126c_1580edd8 );
buf ( n2177 , R_c4d_13d24b58 );
buf ( n2178 , R_62e_13bf7438 );
buf ( n2179 , R_610_14a186f8 );
buf ( n2180 , R_c2f_14a0c038 );
buf ( n2181 , R_124e_117ee338 );
buf ( n2182 , R_186d_15fee348 );
buf ( n2183 , R_e8c_1587e738 );
buf ( n2184 , R_162e_123b25f8 );
buf ( n2185 , R_9f0_140abe58 );
buf ( n2186 , R_14ab_13dd50d8 );
buf ( n2187 , R_86d_14a18dd8 );
buf ( n2188 , R_100f_13d5dad8 );
buf ( n2189 , R_8f8_15ff8668 );
buf ( n2190 , R_f17_14a18e78 );
buf ( n2191 , R_1536_14a0dc58 );
buf ( n2192 , R_15a3_12fc08d8 );
buf ( n2193 , R_f84_117e8d98 );
buf ( n2194 , R_965_140b2578 );
buf ( n2195 , R_d71_14b23018 );
buf ( n2196 , R_b0b_13c21e78 );
buf ( n2197 , R_1390_17016a08 );
buf ( n2198 , R_19af_11636458 );
buf ( n2199 , R_1749_117ec178 );
buf ( n2200 , R_752_15ff64a8 );
buf ( n2201 , R_112a_1587e0f8 );
buf ( n2202 , R_18b6_13bf3018 );
buf ( n2203 , R_1223_13dd8418 );
buf ( n2204 , R_1297_13b99738 );
buf ( n2205 , R_1842_123b43f8 );
buf ( n2206 , R_c78_15887018 );
buf ( n2207 , R_659_123b34f8 );
buf ( n2208 , R_5e5_13df0578 );
buf ( n2209 , R_c04_13cd6f38 );
buf ( n2210 , R_954_17014988 );
buf ( n2211 , R_909_13d3efd8 );
buf ( n2212 , R_f28_13bf6fd8 );
buf ( n2213 , R_1547_13df7b98 );
buf ( n2214 , R_1592_156b9918 );
buf ( n2215 , R_f73_13d22a38 );
buf ( n2216 , R_70d_13beb098 );
buf ( n2217 , R_178e_13c1cb58 );
buf ( n2218 , R_196a_156b6d58 );
buf ( n2219 , R_d2c_14a0ec98 );
buf ( n2220 , R_116f_13d3e7b8 );
buf ( n2221 , R_134b_15ff6cc8 );
buf ( n2222 , R_b50_15815598 );
buf ( n2223 , R_caf_156adc58 );
buf ( n2224 , R_bcd_1162baf8 );
buf ( n2225 , R_690_13c1e098 );
buf ( n2226 , R_18ed_124c3278 );
buf ( n2227 , R_11ec_1008d0b8 );
buf ( n2228 , R_12ce_13c071b8 );
buf ( n2229 , R_180b_1008abd8 );
buf ( n2230 , R_5ae_13cd7ed8 );
buf ( n2231 , R_177b_1007d6b8 );
buf ( n2232 , R_d3f_13cd10d8 );
buf ( n2233 , R_115c_150e8f18 );
buf ( n2234 , R_135e_11c696f8 );
buf ( n2235 , R_b3d_13dddeb8 );
buf ( n2236 , R_720_13d395d8 );
buf ( n2237 , R_197d_14a15458 );
buf ( n2238 , R_1700_140ae8d8 );
buf ( n2239 , R_10e1_13c07758 );
buf ( n2240 , R_ac2_156ad2f8 );
buf ( n2241 , R_79b_15886398 );
buf ( n2242 , R_dba_116373f8 );
buf ( n2243 , R_13d9_14a14378 );
buf ( n2244 , R_19f8_117ef558 );
buf ( n2245 , R_595_13def178 );
buf ( n2246 , R_17f2_1580c998 );
buf ( n2247 , R_1906_13ccad78 );
buf ( n2248 , R_6a9_15ff4ba8 );
buf ( n2249 , R_bb4_117f4d78 );
buf ( n2250 , R_12e7_13cd42d8 );
buf ( n2251 , R_11d3_1162b0f8 );
buf ( n2252 , R_cc8_123b7738 );
buf ( n2253 , R_d48_13c21c98 );
buf ( n2254 , R_1772_14a16998 );
buf ( n2255 , R_1367_15880858 );
buf ( n2256 , R_1153_117f1678 );
buf ( n2257 , R_1986_11c6c038 );
buf ( n2258 , R_729_117f72f8 );
buf ( n2259 , R_b34_158825b8 );
buf ( n2260 , R_ff5_13c2a618 );
buf ( n2261 , R_ea6_150dd7f8 );
buf ( n2262 , R_9d6_13c01f38 );
buf ( n2263 , R_14c5_14a0e518 );
buf ( n2264 , R_1614_156b2b18 );
buf ( n2265 , R_887_14a18298 );
buf ( n2266 , R_848_13ddf218 );
buf ( n2267 , R_1653_14869438 );
buf ( n2268 , R_1486_156afe18 );
buf ( n2269 , R_a15_1700ed08 );
buf ( n2270 , R_e67_117f4e18 );
buf ( n2271 , R_1034_156ac5d8 );
buf ( n2272 , R_8eb_150db1d8 );
buf ( n2273 , R_15b0_1580bdb8 );
buf ( n2274 , R_f0a_14a0ce98 );
buf ( n2275 , R_f91_117f6f38 );
buf ( n2276 , R_1529_123bca58 );
buf ( n2277 , R_972_13ccc038 );
buf ( n2278 , R_1a10_123b4718 );
buf ( n2279 , R_13f1_13d24298 );
buf ( n2280 , R_dd2_14a19198 );
buf ( n2281 , R_7b3_13c07938 );
buf ( n2282 , R_aaa_13b8cfd8 );
buf ( n2283 , R_10c9_15812a78 );
buf ( n2284 , R_16e8_13cd8d38 );
buf ( n2285 , R_d64_15ff5968 );
buf ( n2286 , R_b18_117f40f8 );
buf ( n2287 , R_1383_13c2a438 );
buf ( n2288 , R_19a2_117f01d8 );
buf ( n2289 , R_1756_123c0f18 );
buf ( n2290 , R_1137_13d20ff8 );
buf ( n2291 , R_745_13c1d5f8 );
buf ( n2292 , R_1636_14b22618 );
buf ( n2293 , R_9f8_13decdd8 );
buf ( n2294 , R_e84_14875b98 );
buf ( n2295 , R_1017_13d3bbf8 );
buf ( n2296 , R_865_13d4e7b8 );
buf ( n2297 , R_14a3_11c6d078 );
buf ( n2298 , R_83e_13d43ad8 );
buf ( n2299 , R_a1f_13d22d58 );
buf ( n2300 , R_147c_1580d398 );
buf ( n2301 , R_103e_13d57958 );
buf ( n2302 , R_e5d_1486ddf8 );
buf ( n2303 , R_165d_13bec038 );
buf ( n2304 , R_1494_117f6718 );
buf ( n2305 , R_1645_11c6c178 );
buf ( n2306 , R_a07_14b251d8 );
buf ( n2307 , R_e75_1580a5f8 );
buf ( n2308 , R_1026_158103b8 );
buf ( n2309 , R_856_13cd2a78 );
buf ( n2310 , R_188c_13d39ad8 );
buf ( n2311 , R_126d_11636638 );
buf ( n2312 , R_c4e_13c0fe58 );
buf ( n2313 , R_62f_116305f8 );
buf ( n2314 , R_60f_13bf44b8 );
buf ( n2315 , R_c2e_156b6c18 );
buf ( n2316 , R_124d_123b5438 );
buf ( n2317 , R_186c_15817758 );
buf ( n2318 , R_57b_12fc1f58 );
buf ( n2319 , R_6c3_14a11718 );
buf ( n2320 , R_17d8_13bf24d8 );
buf ( n2321 , R_1301_13ccee78 );
buf ( n2322 , R_b9a_140b40f8 );
buf ( n2323 , R_ce2_156b49b8 );
buf ( n2324 , R_11b9_13d5d5d8 );
buf ( n2325 , R_1920_117ea198 );
buf ( n2326 , R_1713_14a0f878 );
buf ( n2327 , R_10f4_13de4c18 );
buf ( n2328 , R_ad5_117ed1b8 );
buf ( n2329 , R_788_117e8ed8 );
buf ( n2330 , R_da7_11635ff8 );
buf ( n2331 , R_13c6_123c10f8 );
buf ( n2332 , R_19e5_1580eb58 );
buf ( n2333 , R_e90_11637038 );
buf ( n2334 , R_9ec_117eb958 );
buf ( n2335 , R_162a_117ec0d8 );
buf ( n2336 , R_14af_156abdb8 );
buf ( n2337 , R_871_1587f138 );
buf ( n2338 , R_100b_11631d18 );
buf ( n2339 , R_111b_1580faf8 );
buf ( n2340 , R_139f_150df058 );
buf ( n2341 , R_afc_117f8158 );
buf ( n2342 , R_19be_13ccfff8 );
buf ( n2343 , R_761_12fbf078 );
buf ( n2344 , R_173a_156b5a98 );
buf ( n2345 , R_d80_13c1d418 );
buf ( n2346 , R_58a_13ddaf38 );
buf ( n2347 , R_1911_124c4038 );
buf ( n2348 , R_17e7_15883198 );
buf ( n2349 , R_6b4_15881bb8 );
buf ( n2350 , R_ba9_13d5c958 );
buf ( n2351 , R_12f2_17013c68 );
buf ( n2352 , R_11c8_11634fb8 );
buf ( n2353 , R_cd3_13c06178 );
buf ( n2354 , R_6fc_13de34f8 );
buf ( n2355 , R_1180_13ddc298 );
buf ( n2356 , R_1959_14a14698 );
buf ( n2357 , R_d1b_13cd9558 );
buf ( n2358 , R_b61_13d22538 );
buf ( n2359 , R_179f_150e5818 );
buf ( n2360 , R_133a_13d57138 );
buf ( n2361 , R_be4_15817bb8 );
buf ( n2362 , R_c98_13dec298 );
buf ( n2363 , R_1203_1587d978 );
buf ( n2364 , R_679_123b7918 );
buf ( n2365 , R_1822_117e9018 );
buf ( n2366 , R_18d6_13c2ad98 );
buf ( n2367 , R_5c5_1162b5f8 );
buf ( n2368 , R_12b7_117f83d8 );
buf ( n2369 , R_ca8_14a11038 );
buf ( n2370 , R_bd4_11637ad8 );
buf ( n2371 , R_689_158869d8 );
buf ( n2372 , R_11f3_116300f8 );
buf ( n2373 , R_18e6_156b1678 );
buf ( n2374 , R_1812_11c6f558 );
buf ( n2375 , R_12c7_13b97c58 );
buf ( n2376 , R_5b5_11637fd8 );
buf ( n2377 , R_177e_14b1a738 );
buf ( n2378 , R_d3c_13b8b278 );
buf ( n2379 , R_115f_156ac7b8 );
buf ( n2380 , R_135b_13d38b38 );
buf ( n2381 , R_b40_158142d8 );
buf ( n2382 , R_71d_13c1ea98 );
buf ( n2383 , R_197a_13c0a318 );
buf ( n2384 , R_e16_17018088 );
buf ( n2385 , R_1085_13c03e78 );
buf ( n2386 , R_7f7_15888b98 );
buf ( n2387 , R_16a4_158821f8 );
buf ( n2388 , R_1a54_13de0438 );
buf ( n2389 , R_1435_10082258 );
buf ( n2390 , R_a66_15882838 );
buf ( n2391 , R_703_14867bd8 );
buf ( n2392 , R_1960_1162c958 );
buf ( n2393 , R_1179_13d3c7d8 );
buf ( n2394 , R_d22_13d599d8 );
buf ( n2395 , R_b5a_13bf68f8 );
buf ( n2396 , R_1341_13d458d8 );
buf ( n2397 , R_1798_1700e9e8 );
buf ( n2398 , R_171e_13df60b8 );
buf ( n2399 , R_10ff_13ddcab8 );
buf ( n2400 , R_ae0_14a11f38 );
buf ( n2401 , R_77d_13d27df8 );
buf ( n2402 , R_d9c_13ccd4d8 );
buf ( n2403 , R_13bb_1587d478 );
buf ( n2404 , R_19da_13dd5a38 );
buf ( n2405 , R_108a_1486e938 );
buf ( n2406 , R_e11_13cd8c98 );
buf ( n2407 , R_16a9_14a130b8 );
buf ( n2408 , R_7f2_156b2938 );
buf ( n2409 , R_1a4f_13d3a618 );
buf ( n2410 , R_a6b_13b8e1f8 );
buf ( n2411 , R_1430_13dd84b8 );
buf ( n2412 , R_d4b_117f6178 );
buf ( n2413 , R_176f_13d447f8 );
buf ( n2414 , R_136a_13c26838 );
buf ( n2415 , R_1150_15ff71c8 );
buf ( n2416 , R_1989_13ccbc78 );
buf ( n2417 , R_72c_10083c98 );
buf ( n2418 , R_b31_13d44c58 );
buf ( n2419 , R_814_13d51eb8 );
buf ( n2420 , R_1068_1580ea18 );
buf ( n2421 , R_1687_123b81d8 );
buf ( n2422 , R_1452_13df0938 );
buf ( n2423 , R_e33_14a0c3f8 );
buf ( n2424 , R_a49_14a0eb58 );
buf ( n2425 , R_1851_13d5b058 );
buf ( n2426 , R_18a7_13b96858 );
buf ( n2427 , R_1288_13c1daf8 );
buf ( n2428 , R_c69_156af738 );
buf ( n2429 , R_64a_11629438 );
buf ( n2430 , R_5f4_140b13f8 );
buf ( n2431 , R_c13_1162db78 );
buf ( n2432 , R_1232_156aaa58 );
buf ( n2433 , R_15bb_117f3338 );
buf ( n2434 , R_8e0_14a0f698 );
buf ( n2435 , R_f9c_14a104f8 );
buf ( n2436 , R_eff_13d381d8 );
buf ( n2437 , R_151e_15883af8 );
buf ( n2438 , R_97d_14a16178 );
buf ( n2439 , R_1702_13cd9198 );
buf ( n2440 , R_10e3_117f2f78 );
buf ( n2441 , R_ac4_1700f028 );
buf ( n2442 , R_799_13d5a018 );
buf ( n2443 , R_db8_150e6998 );
buf ( n2444 , R_13d7_14b1d1b8 );
buf ( n2445 , R_19f6_1580aa58 );
buf ( n2446 , R_14fd_156b56d8 );
buf ( n2447 , R_15dc_123bfd98 );
buf ( n2448 , R_fbd_14a0b098 );
buf ( n2449 , R_8bf_14875f58 );
buf ( n2450 , R_99e_15ff9388 );
buf ( n2451 , R_ede_11634338 );
buf ( n2452 , R_188d_17018e48 );
buf ( n2453 , R_126e_150e04f8 );
buf ( n2454 , R_c4f_15814918 );
buf ( n2455 , R_630_13d25558 );
buf ( n2456 , R_60e_13cd3d38 );
buf ( n2457 , R_c2d_1580aaf8 );
buf ( n2458 , R_124c_13d40018 );
buf ( n2459 , R_186b_13d42bd8 );
buf ( n2460 , R_1a23_13d52458 );
buf ( n2461 , R_1404_1486a8d8 );
buf ( n2462 , R_de5_11633a78 );
buf ( n2463 , R_7c6_156b9738 );
buf ( n2464 , R_a97_13c05e58 );
buf ( n2465 , R_10b6_124c3638 );
buf ( n2466 , R_16d5_123bc4b8 );
buf ( n2467 , R_bed_13b90db8 );
buf ( n2468 , R_c8f_117ef4b8 );
buf ( n2469 , R_120c_13ddcd38 );
buf ( n2470 , R_670_13ccfaf8 );
buf ( n2471 , R_182b_13cd80b8 );
buf ( n2472 , R_18cd_13c1ca18 );
buf ( n2473 , R_5ce_14b1ded8 );
buf ( n2474 , R_12ae_13c1f178 );
buf ( n2475 , R_bc6_13cd7bb8 );
buf ( n2476 , R_697_13bf83d8 );
buf ( n2477 , R_18f4_15881cf8 );
buf ( n2478 , R_11e5_1162add8 );
buf ( n2479 , R_12d5_17015928 );
buf ( n2480 , R_1804_150e44b8 );
buf ( n2481 , R_5a7_12fbe178 );
buf ( n2482 , R_cb6_1162e398 );
buf ( n2483 , R_110f_15887518 );
buf ( n2484 , R_19ca_156b8a18 );
buf ( n2485 , R_af0_17012a48 );
buf ( n2486 , R_76d_156b1df8 );
buf ( n2487 , R_d8c_15814b98 );
buf ( n2488 , R_172e_117ed438 );
buf ( n2489 , R_13ab_13b99878 );
buf ( n2490 , R_1a12_13d52ef8 );
buf ( n2491 , R_13f3_156b74d8 );
buf ( n2492 , R_dd4_140ac5d8 );
buf ( n2493 , R_7b5_13c1f718 );
buf ( n2494 , R_aa8_14a0ea18 );
buf ( n2495 , R_10c7_13df2c38 );
buf ( n2496 , R_16e6_156b9eb8 );
buf ( n2497 , R_15cd_13cd86f8 );
buf ( n2498 , R_8ce_13d1e2f8 );
buf ( n2499 , R_fae_13bf6df8 );
buf ( n2500 , R_eed_15812578 );
buf ( n2501 , R_98f_117f62b8 );
buf ( n2502 , R_150c_15ff3848 );
buf ( n2503 , R_908_123c0658 );
buf ( n2504 , R_f27_13cd08b8 );
buf ( n2505 , R_1546_14a18f18 );
buf ( n2506 , R_1593_13d58e98 );
buf ( n2507 , R_f74_158805d8 );
buf ( n2508 , R_955_1580f0f8 );
buf ( n2509 , R_d5c_1580ed38 );
buf ( n2510 , R_137b_13d5cc78 );
buf ( n2511 , R_175e_15813478 );
buf ( n2512 , R_199a_117e8b18 );
buf ( n2513 , R_113f_123b3098 );
buf ( n2514 , R_73d_13c220f8 );
buf ( n2515 , R_b20_13c06c18 );
buf ( n2516 , R_163a_13d3ddb8 );
buf ( n2517 , R_9fc_14a0b818 );
buf ( n2518 , R_e80_11633ed8 );
buf ( n2519 , R_101b_123b6518 );
buf ( n2520 , R_861_124c3bd8 );
buf ( n2521 , R_149f_123b5e38 );
buf ( n2522 , R_1080_14a149b8 );
buf ( n2523 , R_7fc_13d3f258 );
buf ( n2524 , R_169f_124c2d78 );
buf ( n2525 , R_1a59_117eded8 );
buf ( n2526 , R_143a_14a0edd8 );
buf ( n2527 , R_a61_1700dd68 );
buf ( n2528 , R_e1b_13cd1178 );
buf ( n2529 , R_140f_117f1cb8 );
buf ( n2530 , R_df0_13c09cd8 );
buf ( n2531 , R_7d1_14b28978 );
buf ( n2532 , R_a8c_123c0338 );
buf ( n2533 , R_10ab_13df0398 );
buf ( n2534 , R_16ca_13d52f98 );
buf ( n2535 , R_1a2e_13c22698 );
buf ( n2536 , R_b10_14b21fd8 );
buf ( n2537 , R_138b_156b0318 );
buf ( n2538 , R_19aa_14a194b8 );
buf ( n2539 , R_174e_15811a38 );
buf ( n2540 , R_74d_117f0e58 );
buf ( n2541 , R_112f_156aac38 );
buf ( n2542 , R_d6c_156b62b8 );
buf ( n2543 , R_1781_1162d5d8 );
buf ( n2544 , R_d39_15811b78 );
buf ( n2545 , R_1162_124c2558 );
buf ( n2546 , R_1358_156b8e78 );
buf ( n2547 , R_b43_13c06858 );
buf ( n2548 , R_71a_117ee798 );
buf ( n2549 , R_1977_15880b78 );
buf ( n2550 , R_1108_13ccfb98 );
buf ( n2551 , R_ae9_1580cd58 );
buf ( n2552 , R_774_1700a7a8 );
buf ( n2553 , R_d93_13cce0b8 );
buf ( n2554 , R_13b2_15886898 );
buf ( n2555 , R_1727_14870e18 );
buf ( n2556 , R_19d1_123b5b18 );
buf ( n2557 , R_188e_11c6a698 );
buf ( n2558 , R_126f_14b23c98 );
buf ( n2559 , R_c50_13d471d8 );
buf ( n2560 , R_631_13ddd7d8 );
buf ( n2561 , R_60d_117f3a18 );
buf ( n2562 , R_c2c_13d2c498 );
buf ( n2563 , R_124b_156b97d8 );
buf ( n2564 , R_186a_13ddb118 );
buf ( n2565 , R_fdc_1162ca98 );
buf ( n2566 , R_14de_13c202f8 );
buf ( n2567 , R_9bd_11632cb8 );
buf ( n2568 , R_8a0_13bf81f8 );
buf ( n2569 , R_15fb_123ba078 );
buf ( n2570 , R_ebf_13b91678 );
buf ( n2571 , R_e94_148719f8 );
buf ( n2572 , R_9e8_15ff97e8 );
buf ( n2573 , R_1626_13de2918 );
buf ( n2574 , R_14b3_13dde9f8 );
buf ( n2575 , R_875_156aea18 );
buf ( n2576 , R_1007_15881578 );
buf ( n2577 , R_14f6_11638938 );
buf ( n2578 , R_fc4_1580d578 );
buf ( n2579 , R_8b8_123ba2f8 );
buf ( n2580 , R_9a5_117ecc18 );
buf ( n2581 , R_ed7_14a0da78 );
buf ( n2582 , R_15e3_123c0158 );
buf ( n2583 , R_e0c_1700d0e8 );
buf ( n2584 , R_16ae_123b38b8 );
buf ( n2585 , R_7ed_117ef738 );
buf ( n2586 , R_1a4a_12fc1c38 );
buf ( n2587 , R_a70_150dbc78 );
buf ( n2588 , R_142b_15889bd8 );
buf ( n2589 , R_108f_13de36d8 );
buf ( n2590 , R_d4e_11c6b6d8 );
buf ( n2591 , R_176c_13ddfcb8 );
buf ( n2592 , R_136d_11634dd8 );
buf ( n2593 , R_114d_158861b8 );
buf ( n2594 , R_198c_13d53a38 );
buf ( n2595 , R_72f_11637498 );
buf ( n2596 , R_b2e_170098a8 );
buf ( n2597 , R_8f7_13b8e298 );
buf ( n2598 , R_f16_1587d838 );
buf ( n2599 , R_1535_13ded2d8 );
buf ( n2600 , R_15a4_1162bcd8 );
buf ( n2601 , R_f85_170174a8 );
buf ( n2602 , R_966_156acd58 );
buf ( n2603 , R_12a4_13cd0db8 );
buf ( n2604 , R_1216_13c26518 );
buf ( n2605 , R_c85_13d505b8 );
buf ( n2606 , R_1835_13b8eb58 );
buf ( n2607 , R_666_13cd8798 );
buf ( n2608 , R_5d8_14a11fd8 );
buf ( n2609 , R_18c3_156b8c98 );
buf ( n2610 , R_bf7_156b4418 );
buf ( n2611 , R_15d5_117ed898 );
buf ( n2612 , R_fb6_14b24558 );
buf ( n2613 , R_8c6_13d442f8 );
buf ( n2614 , R_997_123bb478 );
buf ( n2615 , R_ee5_14a14af8 );
buf ( n2616 , R_1504_13d553d8 );
buf ( n2617 , R_6d1_158167b8 );
buf ( n2618 , R_130f_156ab4f8 );
buf ( n2619 , R_17ca_150df9b8 );
buf ( n2620 , R_b8c_124c3ef8 );
buf ( n2621 , R_cf0_11c6a878 );
buf ( n2622 , R_192e_150e8a18 );
buf ( n2623 , R_11ab_13d29d38 );
buf ( n2624 , R_56d_156b76b8 );
buf ( n2625 , R_1704_13bf4238 );
buf ( n2626 , R_10e5_14871778 );
buf ( n2627 , R_ac6_1587bcb8 );
buf ( n2628 , R_797_14b1c178 );
buf ( n2629 , R_db6_13ddd058 );
buf ( n2630 , R_13d5_1587c618 );
buf ( n2631 , R_19f4_150e3ab8 );
buf ( n2632 , R_1298_156b1d58 );
buf ( n2633 , R_1841_13d2c538 );
buf ( n2634 , R_c79_156b5598 );
buf ( n2635 , R_65a_14874ab8 );
buf ( n2636 , R_5e4_13bf0278 );
buf ( n2637 , R_c03_14a0d2f8 );
buf ( n2638 , R_18b7_13ccd1b8 );
buf ( n2639 , R_1222_14b1acd8 );
buf ( n2640 , R_1073_14b20f98 );
buf ( n2641 , R_809_13d3e678 );
buf ( n2642 , R_1a66_123b6158 );
buf ( n2643 , R_1692_117f31f8 );
buf ( n2644 , R_1447_13b93338 );
buf ( n2645 , R_e28_156abbd8 );
buf ( n2646 , R_a54_13cce838 );
buf ( n2647 , R_1054_13bf8ab8 );
buf ( n2648 , R_1466_13d5abf8 );
buf ( n2649 , R_1673_1580e798 );
buf ( n2650 , R_e47_1587b178 );
buf ( n2651 , R_a35_117f5db8 );
buf ( n2652 , R_828_10081f38 );
buf ( n2653 , R_1469_1587ee18 );
buf ( n2654 , R_1051_11635c38 );
buf ( n2655 , R_e4a_11629118 );
buf ( n2656 , R_1670_1007f238 );
buf ( n2657 , R_82b_13cd7258 );
buf ( n2658 , R_a32_1486afb8 );
buf ( n2659 , R_1187_117f4198 );
buf ( n2660 , R_1952_14a0c0d8 );
buf ( n2661 , R_d14_13dee778 );
buf ( n2662 , R_b68_10089d78 );
buf ( n2663 , R_17a6_15811f38 );
buf ( n2664 , R_1333_117f21b8 );
buf ( n2665 , R_6f5_13d43678 );
buf ( n2666 , R_6c8_1580d758 );
buf ( n2667 , R_1306_1580d938 );
buf ( n2668 , R_17d3_13d3a578 );
buf ( n2669 , R_b95_117f7618 );
buf ( n2670 , R_ce7_13d27218 );
buf ( n2671 , R_1925_15ff0328 );
buf ( n2672 , R_11b4_13b8ec98 );
buf ( n2673 , R_576_13d2bf98 );
buf ( n2674 , R_e00_13cd8bf8 );
buf ( n2675 , R_7e1_150e4058 );
buf ( n2676 , R_a7c_156b7118 );
buf ( n2677 , R_1a3e_14a0b278 );
buf ( n2678 , R_109b_123bd4f8 );
buf ( n2679 , R_141f_1008c578 );
buf ( n2680 , R_16ba_156b6e98 );
buf ( n2681 , R_188f_156b5458 );
buf ( n2682 , R_1270_14a103b8 );
buf ( n2683 , R_c51_11630af8 );
buf ( n2684 , R_632_13ccde38 );
buf ( n2685 , R_60c_13dd9c78 );
buf ( n2686 , R_c2b_14b23478 );
buf ( n2687 , R_124a_140b7898 );
buf ( n2688 , R_1869_14b29cd8 );
buf ( n2689 , R_1a14_117ebbd8 );
buf ( n2690 , R_13f5_13cd8a18 );
buf ( n2691 , R_dd6_13de0d98 );
buf ( n2692 , R_7b7_15816a38 );
buf ( n2693 , R_aa6_13d28c58 );
buf ( n2694 , R_10c5_11632998 );
buf ( n2695 , R_16e4_10087078 );
buf ( n2696 , R_190c_13d1d998 );
buf ( n2697 , R_6af_124c33b8 );
buf ( n2698 , R_bae_1587b5d8 );
buf ( n2699 , R_12ed_14a176b8 );
buf ( n2700 , R_11cd_13cd27f8 );
buf ( n2701 , R_cce_116331b8 );
buf ( n2702 , R_58f_156b9558 );
buf ( n2703 , R_17ec_13dd7fb8 );
buf ( n2704 , R_1057_123bd278 );
buf ( n2705 , R_1463_124c4b78 );
buf ( n2706 , R_1676_140ae6f8 );
buf ( n2707 , R_e44_148741f8 );
buf ( n2708 , R_a38_150dc3f8 );
buf ( n2709 , R_825_123b3278 );
buf ( n2710 , R_18a8_1580c8f8 );
buf ( n2711 , R_1289_13c09738 );
buf ( n2712 , R_c6a_15811fd8 );
buf ( n2713 , R_64b_1007d938 );
buf ( n2714 , R_5f3_116307d8 );
buf ( n2715 , R_c12_1162cc78 );
buf ( n2716 , R_1231_13dee9f8 );
buf ( n2717 , R_1850_1587f778 );
buf ( n2718 , R_146c_14872f38 );
buf ( n2719 , R_104e_1580f7d8 );
buf ( n2720 , R_e4d_14b20d18 );
buf ( n2721 , R_166d_13d20058 );
buf ( n2722 , R_82e_1580f2d8 );
buf ( n2723 , R_a2f_123b3db8 );
buf ( n2724 , R_19c3_116340b8 );
buf ( n2725 , R_af7_13cd2d98 );
buf ( n2726 , R_766_13c07618 );
buf ( n2727 , R_1735_13bf9f58 );
buf ( n2728 , R_d85_13dd7518 );
buf ( n2729 , R_13a4_150ea138 );
buf ( n2730 , R_1116_13c02438 );
buf ( n2731 , R_df9_13dd9458 );
buf ( n2732 , R_7da_14a16fd8 );
buf ( n2733 , R_a83_13b9a278 );
buf ( n2734 , R_10a2_123b3d18 );
buf ( n2735 , R_1a37_1587f958 );
buf ( n2736 , R_16c1_13d3d458 );
buf ( n2737 , R_1418_13d2b1d8 );
buf ( n2738 , R_ea1_156b5c78 );
buf ( n2739 , R_9db_13c05bd8 );
buf ( n2740 , R_1619_15888d78 );
buf ( n2741 , R_14c0_17012fe8 );
buf ( n2742 , R_882_13dee458 );
buf ( n2743 , R_ffa_11c68f78 );
buf ( n2744 , R_1967_15ff9608 );
buf ( n2745 , R_1172_170122c8 );
buf ( n2746 , R_d29_13bed898 );
buf ( n2747 , R_1348_156b1178 );
buf ( n2748 , R_b53_1162fe78 );
buf ( n2749 , R_1791_15ff73a8 );
buf ( n2750 , R_70a_13dee818 );
buf ( n2751 , R_8ea_13b91c18 );
buf ( n2752 , R_15b1_140b0d18 );
buf ( n2753 , R_f09_13d4f9d8 );
buf ( n2754 , R_f92_13b99238 );
buf ( n2755 , R_1528_13cca918 );
buf ( n2756 , R_973_12fc1738 );
buf ( n2757 , R_907_13d1cef8 );
buf ( n2758 , R_f26_13d51378 );
buf ( n2759 , R_1545_13ddab78 );
buf ( n2760 , R_1594_123b52f8 );
buf ( n2761 , R_f75_1587ec38 );
buf ( n2762 , R_956_117f3bf8 );
buf ( n2763 , R_a1c_13d42098 );
buf ( n2764 , R_147f_15ffd208 );
buf ( n2765 , R_103b_12fbfbb8 );
buf ( n2766 , R_e60_13b98dd8 );
buf ( n2767 , R_165a_156b9418 );
buf ( n2768 , R_841_13de1e78 );
buf ( n2769 , R_1715_13c03ab8 );
buf ( n2770 , R_10f6_1587fc78 );
buf ( n2771 , R_ad7_11c6aaf8 );
buf ( n2772 , R_786_13bf7938 );
buf ( n2773 , R_da5_13c24c18 );
buf ( n2774 , R_13c4_156adbb8 );
buf ( n2775 , R_19e3_13b8b4f8 );
buf ( n2776 , R_15c5_13cce478 );
buf ( n2777 , R_8d6_14a156d8 );
buf ( n2778 , R_fa6_13ccd7f8 );
buf ( n2779 , R_ef5_13c0f8b8 );
buf ( n2780 , R_987_148737f8 );
buf ( n2781 , R_1514_13d4ea38 );
buf ( n2782 , R_d36_13cd2938 );
buf ( n2783 , R_1165_1700dae8 );
buf ( n2784 , R_1355_13c0e2d8 );
buf ( n2785 , R_b46_12fbedf8 );
buf ( n2786 , R_717_13c1ebd8 );
buf ( n2787 , R_1974_13b938d8 );
buf ( n2788 , R_1784_14b1b3b8 );
buf ( n2789 , R_156d_13b91d58 );
buf ( n2790 , R_f4e_13d2bb38 );
buf ( n2791 , R_156c_1486f8d8 );
buf ( n2792 , R_92f_1587e418 );
buf ( n2793 , R_f4d_158174d8 );
buf ( n2794 , R_92e_15880df8 );
buf ( n2795 , R_156e_13bee0b8 );
buf ( n2796 , R_f4f_13d1f298 );
buf ( n2797 , R_930_117f5818 );
buf ( n2798 , R_156b_13cd6a38 );
buf ( n2799 , R_f4c_13d4edf8 );
buf ( n2800 , R_92d_13b93838 );
buf ( n2801 , R_156f_1700c828 );
buf ( n2802 , R_f50_13d5d038 );
buf ( n2803 , R_931_1007f198 );
buf ( n2804 , R_92c_13bef238 );
buf ( n2805 , R_156a_14a0d7f8 );
buf ( n2806 , R_f4b_1162df38 );
buf ( n2807 , R_682_13dd6a78 );
buf ( n2808 , R_11fa_12fbfe38 );
buf ( n2809 , R_18df_1162e1b8 );
buf ( n2810 , R_1819_117f44b8 );
buf ( n2811 , R_12c0_156b3478 );
buf ( n2812 , R_5bc_150db098 );
buf ( n2813 , R_ca1_15888af8 );
buf ( n2814 , R_bdb_123b9178 );
buf ( n2815 , R_1890_13c0a4f8 );
buf ( n2816 , R_1271_13cd3e78 );
buf ( n2817 , R_c52_11629cf8 );
buf ( n2818 , R_633_1587c6b8 );
buf ( n2819 , R_60b_17014c08 );
buf ( n2820 , R_c2a_13c01d58 );
buf ( n2821 , R_1249_150de798 );
buf ( n2822 , R_1868_13cd62b8 );
buf ( n2823 , R_105a_14a112b8 );
buf ( n2824 , R_1460_158862f8 );
buf ( n2825 , R_1679_13cd44b8 );
buf ( n2826 , R_e41_14a14e18 );
buf ( n2827 , R_a3b_13cd1998 );
buf ( n2828 , R_822_117e9158 );
buf ( n2829 , R_1570_13d44118 );
buf ( n2830 , R_f51_13ccb778 );
buf ( n2831 , R_932_15810d18 );
buf ( n2832 , R_92b_14a180b8 );
buf ( n2833 , R_f4a_1162c8b8 );
buf ( n2834 , R_1569_13bede38 );
buf ( n2835 , R_163e_12fc0338 );
buf ( n2836 , R_a00_13df4df8 );
buf ( n2837 , R_e7c_13c08798 );
buf ( n2838 , R_101f_117ed9d8 );
buf ( n2839 , R_85d_117f4738 );
buf ( n2840 , R_149b_13cd1038 );
buf ( n2841 , R_146f_117f47d8 );
buf ( n2842 , R_104b_158885f8 );
buf ( n2843 , R_e50_12fbe858 );
buf ( n2844 , R_166a_1587c938 );
buf ( n2845 , R_831_156b2398 );
buf ( n2846 , R_a2c_11c701d8 );
buf ( n2847 , R_801_150e6e98 );
buf ( n2848 , R_169a_13b94878 );
buf ( n2849 , R_1a5e_1162d3f8 );
buf ( n2850 , R_143f_13b8c218 );
buf ( n2851 , R_a5c_13b8c178 );
buf ( n2852 , R_e20_13ddd0f8 );
buf ( n2853 , R_107b_156b2118 );
buf ( n2854 , R_d51_13df3b38 );
buf ( n2855 , R_1769_14b21038 );
buf ( n2856 , R_1370_13cd2618 );
buf ( n2857 , R_114a_13c218d8 );
buf ( n2858 , R_198f_13d28bb8 );
buf ( n2859 , R_732_13d55fb8 );
buf ( n2860 , R_b2b_13ccd2f8 );
buf ( n2861 , R_1571_1580af58 );
buf ( n2862 , R_f52_12fc1ff8 );
buf ( n2863 , R_933_14868718 );
buf ( n2864 , R_92a_13c01a38 );
buf ( n2865 , R_f49_13d4f4d8 );
buf ( n2866 , R_1568_1580c218 );
buf ( n2867 , R_1706_15814eb8 );
buf ( n2868 , R_10e7_14a160d8 );
buf ( n2869 , R_ac8_156afa58 );
buf ( n2870 , R_795_14a12b18 );
buf ( n2871 , R_db4_117edd98 );
buf ( n2872 , R_13d3_13b90f98 );
buf ( n2873 , R_19f2_12fbf258 );
buf ( n2874 , R_17b9_156b0b38 );
buf ( n2875 , R_193f_13d3aa78 );
buf ( n2876 , R_b7b_13befeb8 );
buf ( n2877 , R_d01_140ab318 );
buf ( n2878 , R_119a_13b8a5f8 );
buf ( n2879 , R_1320_14b27f78 );
buf ( n2880 , R_55c_11630e18 );
buf ( n2881 , R_6e2_158149b8 );
buf ( n2882 , R_106b_117f3518 );
buf ( n2883 , R_168a_117eb598 );
buf ( n2884 , R_144f_14b26718 );
buf ( n2885 , R_e30_123b3e58 );
buf ( n2886 , R_a4c_170172c8 );
buf ( n2887 , R_811_15882478 );
buf ( n2888 , R_1406_148665f8 );
buf ( n2889 , R_de7_1007fcd8 );
buf ( n2890 , R_7c8_156b7f78 );
buf ( n2891 , R_a95_117f6cb8 );
buf ( n2892 , R_10b4_13d3d598 );
buf ( n2893 , R_16d3_1700be28 );
buf ( n2894 , R_1a25_13b9a318 );
buf ( n2895 , R_1572_156b67b8 );
buf ( n2896 , R_f53_123c01f8 );
buf ( n2897 , R_934_156b0958 );
buf ( n2898 , R_929_13d5bf58 );
buf ( n2899 , R_f48_13c256b8 );
buf ( n2900 , R_1567_13b91e98 );
buf ( n2901 , R_1943_11c70598 );
buf ( n2902 , R_d05_13c0cd98 );
buf ( n2903 , R_b77_13d415f8 );
buf ( n2904 , R_17b5_14a12118 );
buf ( n2905 , R_1324_15887298 );
buf ( n2906 , R_6e6_13becb78 );
buf ( n2907 , R_558_116299d8 );
buf ( n2908 , R_1196_13d4f398 );
buf ( n2909 , R_e98_13d433f8 );
buf ( n2910 , R_9e4_13cccdf8 );
buf ( n2911 , R_1622_13c044b8 );
buf ( n2912 , R_14b7_13d21318 );
buf ( n2913 , R_879_15884c78 );
buf ( n2914 , R_1003_124c39f8 );
buf ( n2915 , R_1a16_1486b418 );
buf ( n2916 , R_13f7_13d24338 );
buf ( n2917 , R_dd8_1587fd18 );
buf ( n2918 , R_7b9_13c0f458 );
buf ( n2919 , R_aa4_13c1d0f8 );
buf ( n2920 , R_10c3_13ccbef8 );
buf ( n2921 , R_16e2_140b6df8 );
buf ( n2922 , R_1573_14a0c498 );
buf ( n2923 , R_f54_11632858 );
buf ( n2924 , R_935_150e5318 );
buf ( n2925 , R_928_156aab98 );
buf ( n2926 , R_f47_13cd9238 );
buf ( n2927 , R_1566_123b2a58 );
buf ( n2928 , R_a0b_11637858 );
buf ( n2929 , R_e71_14b21a38 );
buf ( n2930 , R_102a_11c6ccb8 );
buf ( n2931 , R_852_14b1d938 );
buf ( n2932 , R_1490_13bf8158 );
buf ( n2933 , R_1649_13dd4f98 );
buf ( n2934 , R_a12_1008b358 );
buf ( n2935 , R_e6a_156b7a78 );
buf ( n2936 , R_1031_14b25778 );
buf ( n2937 , R_84b_156ad1b8 );
buf ( n2938 , R_1650_13dd4e58 );
buf ( n2939 , R_1489_13c21978 );
buf ( n2940 , R_7e8_1486a0b8 );
buf ( n2941 , R_1a45_1162e2f8 );
buf ( n2942 , R_a75_156b0778 );
buf ( n2943 , R_1426_11637718 );
buf ( n2944 , R_1094_13d28398 );
buf ( n2945 , R_16b3_117efeb8 );
buf ( n2946 , R_e07_13d453d8 );
buf ( n2947 , R_17bd_1162b918 );
buf ( n2948 , R_b7f_14a0be58 );
buf ( n2949 , R_cfd_13d1d038 );
buf ( n2950 , R_193b_13d39f38 );
buf ( n2951 , R_119e_13c1bcf8 );
buf ( n2952 , R_560_12fbf118 );
buf ( n2953 , R_6de_13cd4058 );
buf ( n2954 , R_131c_13c245d8 );
buf ( n2955 , R_1891_123b9858 );
buf ( n2956 , R_1272_13dd9ef8 );
buf ( n2957 , R_c53_15ff5148 );
buf ( n2958 , R_634_11631818 );
buf ( n2959 , R_60a_156b2758 );
buf ( n2960 , R_c29_13cd0598 );
buf ( n2961 , R_1248_12fbfcf8 );
buf ( n2962 , R_1867_14a0ded8 );
buf ( n2963 , R_9cd_13d1f518 );
buf ( n2964 , R_14ce_1008b5d8 );
buf ( n2965 , R_160b_14b24cd8 );
buf ( n2966 , R_890_11628df8 );
buf ( n2967 , R_fec_13ccc5d8 );
buf ( n2968 , R_eaf_13d5baf8 );
buf ( n2969 , R_15bc_15889138 );
buf ( n2970 , R_8df_11637358 );
buf ( n2971 , R_f9d_158889b8 );
buf ( n2972 , R_efe_11632b78 );
buf ( n2973 , R_97e_13c29718 );
buf ( n2974 , R_151d_1700bc48 );
buf ( n2975 , R_ae2_123bdef8 );
buf ( n2976 , R_77b_17011828 );
buf ( n2977 , R_d9a_13c047d8 );
buf ( n2978 , R_13b9_15ffc948 );
buf ( n2979 , R_19d8_14870b98 );
buf ( n2980 , R_1720_156b9198 );
buf ( n2981 , R_1101_140b7398 );
buf ( n2982 , R_1202_15881898 );
buf ( n2983 , R_67a_13de2878 );
buf ( n2984 , R_1821_117f1c18 );
buf ( n2985 , R_18d7_1580f378 );
buf ( n2986 , R_5c4_14868fd8 );
buf ( n2987 , R_12b8_11631b38 );
buf ( n2988 , R_be3_13de2198 );
buf ( n2989 , R_c99_13c029d8 );
buf ( n2990 , R_fd1_13c1d058 );
buf ( n2991 , R_14e9_14868538 );
buf ( n2992 , R_9b2_1580b6d8 );
buf ( n2993 , R_8ab_14a0fc38 );
buf ( n2994 , R_15f0_140ae3d8 );
buf ( n2995 , R_eca_14a11df8 );
buf ( n2996 , R_1574_13cd7cf8 );
buf ( n2997 , R_f55_14b1ac38 );
buf ( n2998 , R_936_140acf38 );
buf ( n2999 , R_927_124c4178 );
buf ( n3000 , R_f46_14a0af58 );
buf ( n3001 , R_1565_1700e808 );
buf ( n3002 , R_14d3_1580e5b8 );
buf ( n3003 , R_9c8_15fef248 );
buf ( n3004 , R_895_13d532b8 );
buf ( n3005 , R_1606_1007ef18 );
buf ( n3006 , R_eb4_117eda78 );
buf ( n3007 , R_fe7_1162ba58 );
buf ( n3008 , R_8f6_156b7b18 );
buf ( n3009 , R_f15_158819d8 );
buf ( n3010 , R_15a5_158168f8 );
buf ( n3011 , R_1534_123b9c18 );
buf ( n3012 , R_f86_13c1ce78 );
buf ( n3013 , R_967_11c68938 );
buf ( n3014 , R_1901_15817ed8 );
buf ( n3015 , R_6a4_1162c1d8 );
buf ( n3016 , R_bb9_156ab1d8 );
buf ( n3017 , R_12e2_11636a98 );
buf ( n3018 , R_11d8_156aa738 );
buf ( n3019 , R_cc3_15887c98 );
buf ( n3020 , R_59a_117f76b8 );
buf ( n3021 , R_17f7_117e9838 );
buf ( n3022 , R_105d_123b4998 );
buf ( n3023 , R_145d_123bec18 );
buf ( n3024 , R_167c_140b6178 );
buf ( n3025 , R_e3e_150da7d8 );
buf ( n3026 , R_a3e_11635cd8 );
buf ( n3027 , R_81f_156b45f8 );
buf ( n3028 , R_120b_13def358 );
buf ( n3029 , R_671_140b4058 );
buf ( n3030 , R_182a_117ef698 );
buf ( n3031 , R_18ce_156b4e18 );
buf ( n3032 , R_5cd_14a185b8 );
buf ( n3033 , R_12af_15ff69a8 );
buf ( n3034 , R_bec_124c2878 );
buf ( n3035 , R_c90_117eb778 );
buf ( n3036 , R_1386_14a0c7b8 );
buf ( n3037 , R_19a5_1008a598 );
buf ( n3038 , R_1753_13cd1218 );
buf ( n3039 , R_748_13d3b518 );
buf ( n3040 , R_1134_1580ad78 );
buf ( n3041 , R_d67_13d3caf8 );
buf ( n3042 , R_b15_156b2078 );
buf ( n3043 , R_128a_15880718 );
buf ( n3044 , R_c6b_14a13518 );
buf ( n3045 , R_64c_148739d8 );
buf ( n3046 , R_5f2_13dd5538 );
buf ( n3047 , R_c11_15ff5aa8 );
buf ( n3048 , R_1230_124c42b8 );
buf ( n3049 , R_184f_1587fa98 );
buf ( n3050 , R_18a9_11c6f918 );
buf ( n3051 , R_bbf_1587ddd8 );
buf ( n3052 , R_69e_123b5bb8 );
buf ( n3053 , R_18fb_13df16f8 );
buf ( n3054 , R_11de_10089058 );
buf ( n3055 , R_12dc_13c0bc18 );
buf ( n3056 , R_17fd_13d408d8 );
buf ( n3057 , R_5a0_11631db8 );
buf ( n3058 , R_cbd_14872df8 );
buf ( n3059 , R_691_15883378 );
buf ( n3060 , R_18ee_14a171b8 );
buf ( n3061 , R_11eb_13d4f078 );
buf ( n3062 , R_12cf_158850d8 );
buf ( n3063 , R_180a_13d3fc58 );
buf ( n3064 , R_5ad_14a0c2b8 );
buf ( n3065 , R_cb0_13de1658 );
buf ( n3066 , R_bcc_13df1f18 );
buf ( n3067 , R_1472_13d3c698 );
buf ( n3068 , R_1048_13df8bd8 );
buf ( n3069 , R_e53_10087b18 );
buf ( n3070 , R_1667_13beaf58 );
buf ( n3071 , R_834_15888698 );
buf ( n3072 , R_a29_13de0618 );
buf ( n3073 , R_1575_13d42598 );
buf ( n3074 , R_f56_13c0c578 );
buf ( n3075 , R_937_15886c58 );
buf ( n3076 , R_926_158846d8 );
buf ( n3077 , R_f45_13d4f438 );
buf ( n3078 , R_1564_1587b038 );
buf ( n3079 , R_906_14a145f8 );
buf ( n3080 , R_f25_13d24e78 );
buf ( n3081 , R_1544_124c4fd8 );
buf ( n3082 , R_1595_14b1f698 );
buf ( n3083 , R_f76_117f6fd8 );
buf ( n3084 , R_957_15888878 );
buf ( n3085 , R_c7a_140ac998 );
buf ( n3086 , R_65b_1580b778 );
buf ( n3087 , R_5e3_117eba98 );
buf ( n3088 , R_c02_123b2f58 );
buf ( n3089 , R_18b8_12fc05b8 );
buf ( n3090 , R_1221_15812cf8 );
buf ( n3091 , R_1299_14b1fc38 );
buf ( n3092 , R_1840_13d549d8 );
buf ( n3093 , R_1947_156ac3f8 );
buf ( n3094 , R_d09_150dd438 );
buf ( n3095 , R_b73_117f7938 );
buf ( n3096 , R_17b1_14a0dcf8 );
buf ( n3097 , R_1328_13d2aeb8 );
buf ( n3098 , R_6ea_123bbb58 );
buf ( n3099 , R_1192_1587dbf8 );
buf ( n3100 , R_137e_13c27738 );
buf ( n3101 , R_175b_15883ff8 );
buf ( n3102 , R_199d_1008a6d8 );
buf ( n3103 , R_113c_13d20eb8 );
buf ( n3104 , R_740_13bf6b78 );
buf ( n3105 , R_b1d_123c1918 );
buf ( n3106 , R_d5f_15888c38 );
buf ( n3107 , R_fcb_13def8f8 );
buf ( n3108 , R_8b1_170124a8 );
buf ( n3109 , R_9ac_14a190f8 );
buf ( n3110 , R_ed0_13d23d98 );
buf ( n3111 , R_15ea_1580e658 );
buf ( n3112 , R_14ef_123bead8 );
buf ( n3113 , R_d33_123bd8b8 );
buf ( n3114 , R_1168_156b6fd8 );
buf ( n3115 , R_1352_13c10b78 );
buf ( n3116 , R_b49_14a158b8 );
buf ( n3117 , R_714_1587c898 );
buf ( n3118 , R_1971_13ddfe98 );
buf ( n3119 , R_1787_1486e2f8 );
buf ( n3120 , R_68a_14a15b38 );
buf ( n3121 , R_11f2_1162a6f8 );
buf ( n3122 , R_18e7_13c08c98 );
buf ( n3123 , R_1811_117e9a18 );
buf ( n3124 , R_12c8_140aa878 );
buf ( n3125 , R_5b4_140b2a78 );
buf ( n3126 , R_ca9_15887e78 );
buf ( n3127 , R_bd3_13c0e9b8 );
buf ( n3128 , R_195d_15884818 );
buf ( n3129 , R_117c_14874838 );
buf ( n3130 , R_d1f_1007f698 );
buf ( n3131 , R_b5d_123bb8d8 );
buf ( n3132 , R_133e_13d55dd8 );
buf ( n3133 , R_179b_12fbde58 );
buf ( n3134 , R_700_13cd9878 );
buf ( n3135 , R_1576_1700c6e8 );
buf ( n3136 , R_f57_14a14198 );
buf ( n3137 , R_938_13bedc58 );
buf ( n3138 , R_925_13df1338 );
buf ( n3139 , R_f44_156b99b8 );
buf ( n3140 , R_1563_158841d8 );
buf ( n3141 , R_c86_14a12e38 );
buf ( n3142 , R_1834_13cd3f18 );
buf ( n3143 , R_667_1486b558 );
buf ( n3144 , R_5d7_156b0c78 );
buf ( n3145 , R_18c4_11c709f8 );
buf ( n3146 , R_bf6_11c6f378 );
buf ( n3147 , R_12a5_1162d718 );
buf ( n3148 , R_1215_117f51d8 );
buf ( n3149 , R_1892_13d3b1f8 );
buf ( n3150 , R_1273_13dd5c18 );
buf ( n3151 , R_c54_13becd58 );
buf ( n3152 , R_635_13d2c678 );
buf ( n3153 , R_609_1580ef18 );
buf ( n3154 , R_c28_140ba098 );
buf ( n3155 , R_1247_13ccda78 );
buf ( n3156 , R_1866_13bf9eb8 );
buf ( n3157 , R_9d2_13ccb958 );
buf ( n3158 , R_14c9_117f80b8 );
buf ( n3159 , R_1610_1700a988 );
buf ( n3160 , R_88b_1587e5f8 );
buf ( n3161 , R_ff1_13b8bd18 );
buf ( n3162 , R_eaa_13dd6618 );
buf ( n3163 , R_1708_11630558 );
buf ( n3164 , R_10e9_123c2138 );
buf ( n3165 , R_aca_14a131f8 );
buf ( n3166 , R_793_12fc2138 );
buf ( n3167 , R_db2_123b68d8 );
buf ( n3168 , R_13d1_156ac998 );
buf ( n3169 , R_19f0_13d47138 );
buf ( n3170 , R_7d3_13dd99f8 );
buf ( n3171 , R_a8a_150e0ef8 );
buf ( n3172 , R_10a9_1486ae78 );
buf ( n3173 , R_16c8_13dfaed8 );
buf ( n3174 , R_1a30_14a19698 );
buf ( n3175 , R_1411_13dfa438 );
buf ( n3176 , R_df2_150e09f8 );
buf ( n3177 , R_14e3_11634838 );
buf ( n3178 , R_9b8_13d43b78 );
buf ( n3179 , R_8a5_13bee798 );
buf ( n3180 , R_15f6_117f0458 );
buf ( n3181 , R_ec4_11c68a78 );
buf ( n3182 , R_fd7_116387f8 );
buf ( n3183 , R_17c1_13d57d18 );
buf ( n3184 , R_b83_13bedd98 );
buf ( n3185 , R_cf9_1587d798 );
buf ( n3186 , R_1937_150e3c98 );
buf ( n3187 , R_11a2_13c05138 );
buf ( n3188 , R_564_15815278 );
buf ( n3189 , R_6da_13c00f98 );
buf ( n3190 , R_1318_1008a9f8 );
buf ( n3191 , R_faf_158866b8 );
buf ( n3192 , R_8cd_15ff2ee8 );
buf ( n3193 , R_eec_117f7078 );
buf ( n3194 , R_990_11633c58 );
buf ( n3195 , R_150b_13cd8dd8 );
buf ( n3196 , R_15ce_13df0898 );
buf ( n3197 , R_1766_116318b8 );
buf ( n3198 , R_1373_15810598 );
buf ( n3199 , R_1147_13b8d438 );
buf ( n3200 , R_1992_13b8d1b8 );
buf ( n3201 , R_735_13cd4cd8 );
buf ( n3202 , R_b28_1162fab8 );
buf ( n3203 , R_d54_150e15d8 );
buf ( n3204 , R_1577_13d44ed8 );
buf ( n3205 , R_f58_13d3e178 );
buf ( n3206 , R_939_123b2878 );
buf ( n3207 , R_924_140b7118 );
buf ( n3208 , R_f43_140aeab8 );
buf ( n3209 , R_1562_100874d8 );
buf ( n3210 , R_17ce_13d50b58 );
buf ( n3211 , R_b90_14a17e38 );
buf ( n3212 , R_cec_156b8fb8 );
buf ( n3213 , R_192a_13df93f8 );
buf ( n3214 , R_11af_156b2a78 );
buf ( n3215 , R_571_13b96ad8 );
buf ( n3216 , R_6cd_150dc5d8 );
buf ( n3217 , R_130b_14b1eab8 );
buf ( n3218 , R_19b7_117f7758 );
buf ( n3219 , R_75a_150de5b8 );
buf ( n3220 , R_1741_100824d8 );
buf ( n3221 , R_d79_1008a638 );
buf ( n3222 , R_1122_150e9a58 );
buf ( n3223 , R_1398_10083978 );
buf ( n3224 , R_b03_158129d8 );
buf ( n3225 , R_14d8_13cd4698 );
buf ( n3226 , R_9c3_13befa58 );
buf ( n3227 , R_89a_117edb18 );
buf ( n3228 , R_1601_13d272b8 );
buf ( n3229 , R_eb9_11638438 );
buf ( n3230 , R_fe2_13defdf8 );
buf ( n3231 , R_13f9_1580cb78 );
buf ( n3232 , R_dda_117f7118 );
buf ( n3233 , R_7bb_13bf54f8 );
buf ( n3234 , R_aa2_12fc1a58 );
buf ( n3235 , R_10c1_13b901d8 );
buf ( n3236 , R_16e0_158811b8 );
buf ( n3237 , R_1a18_156b8bf8 );
buf ( n3238 , R_fbe_13cd90f8 );
buf ( n3239 , R_8be_13df3278 );
buf ( n3240 , R_99f_123b6b58 );
buf ( n3241 , R_edd_13b99cd8 );
buf ( n3242 , R_15dd_156aef18 );
buf ( n3243 , R_14fc_140b09f8 );
buf ( n3244 , R_19b2_150e0318 );
buf ( n3245 , R_1746_123b75f8 );
buf ( n3246 , R_755_14a13338 );
buf ( n3247 , R_1127_13de3318 );
buf ( n3248 , R_d74_17011d28 );
buf ( n3249 , R_b08_150dce98 );
buf ( n3250 , R_1393_11c68c58 );
buf ( n3251 , R_1956_15813158 );
buf ( n3252 , R_d18_156b9698 );
buf ( n3253 , R_b64_156b3a18 );
buf ( n3254 , R_17a2_117e8758 );
buf ( n3255 , R_1337_13d20af8 );
buf ( n3256 , R_6f9_17012b88 );
buf ( n3257 , R_1183_1580f698 );
buf ( n3258 , R_bb3_17013d08 );
buf ( n3259 , R_12e8_14b1e158 );
buf ( n3260 , R_11d2_124c3318 );
buf ( n3261 , R_cc9_11c6e018 );
buf ( n3262 , R_594_13cd9698 );
buf ( n3263 , R_17f1_13c0bdf8 );
buf ( n3264 , R_1907_13ccaa58 );
buf ( n3265 , R_6aa_13de4038 );
buf ( n3266 , R_ba3_13cd5bd8 );
buf ( n3267 , R_12f8_13cd2758 );
buf ( n3268 , R_11c2_13c1fc18 );
buf ( n3269 , R_cd9_14b1f878 );
buf ( n3270 , R_584_12fc0bf8 );
buf ( n3271 , R_1917_13d21f98 );
buf ( n3272 , R_17e1_13d37878 );
buf ( n3273 , R_6ba_11637b78 );
buf ( n3274 , R_8e9_13cd6b78 );
buf ( n3275 , R_15b2_117f08b8 );
buf ( n3276 , R_f08_156b5db8 );
buf ( n3277 , R_f93_13b92758 );
buf ( n3278 , R_1527_13ccaeb8 );
buf ( n3279 , R_974_13c0c2f8 );
buf ( n3280 , R_ad9_150e2a78 );
buf ( n3281 , R_784_13dfa4d8 );
buf ( n3282 , R_da3_14a0cd58 );
buf ( n3283 , R_13c2_13d2a4b8 );
buf ( n3284 , R_19e1_1700c5a8 );
buf ( n3285 , R_1717_13df61f8 );
buf ( n3286 , R_10f8_156b7258 );
buf ( n3287 , R_1578_123bab18 );
buf ( n3288 , R_f59_13c10358 );
buf ( n3289 , R_93a_1486f978 );
buf ( n3290 , R_923_11632178 );
buf ( n3291 , R_f42_14b1f9b8 );
buf ( n3292 , R_1561_13bf4a58 );
buf ( n3293 , R_1060_13c0b358 );
buf ( n3294 , R_145a_14a12bb8 );
buf ( n3295 , R_167f_14a19378 );
buf ( n3296 , R_e3b_13dd7f18 );
buf ( n3297 , R_a41_14a10d18 );
buf ( n3298 , R_81c_13bf79d8 );
buf ( n3299 , R_12fd_1007d9d8 );
buf ( n3300 , R_b9e_123ba618 );
buf ( n3301 , R_cde_13d39218 );
buf ( n3302 , R_11bd_11c6dcf8 );
buf ( n3303 , R_191c_1580c038 );
buf ( n3304 , R_57f_158160d8 );
buf ( n3305 , R_6bf_13df4e98 );
buf ( n3306 , R_17dc_15ff5508 );
buf ( n3307 , R_1893_117f0d18 );
buf ( n3308 , R_1274_156b1218 );
buf ( n3309 , R_c55_13cce338 );
buf ( n3310 , R_636_123c1238 );
buf ( n3311 , R_608_13d58678 );
buf ( n3312 , R_c27_13bf2a78 );
buf ( n3313 , R_1246_14b229d8 );
buf ( n3314 , R_1865_156b4d78 );
buf ( n3315 , R_772_11634a18 );
buf ( n3316 , R_d91_13c0fdb8 );
buf ( n3317 , R_13b0_1486d0d8 );
buf ( n3318 , R_1729_123b6338 );
buf ( n3319 , R_19cf_11c70c78 );
buf ( n3320 , R_110a_156b12b8 );
buf ( n3321 , R_aeb_11638758 );
buf ( n3322 , R_e78_117ef0f8 );
buf ( n3323 , R_1023_15ff3ac8 );
buf ( n3324 , R_859_13c0f098 );
buf ( n3325 , R_1497_116337f8 );
buf ( n3326 , R_1642_1162e578 );
buf ( n3327 , R_a04_13c22e18 );
buf ( n3328 , R_76b_13ddaad8 );
buf ( n3329 , R_d8a_10085458 );
buf ( n3330 , R_1730_11c6fd78 );
buf ( n3331 , R_13a9_15887978 );
buf ( n3332 , R_1111_11629c58 );
buf ( n3333 , R_19c8_123b61f8 );
buf ( n3334 , R_af2_11635558 );
buf ( n3335 , R_1045_13c2abb8 );
buf ( n3336 , R_e56_13c1f0d8 );
buf ( n3337 , R_1664_1700d9a8 );
buf ( n3338 , R_837_13d43c18 );
buf ( n3339 , R_a26_13c28c78 );
buf ( n3340 , R_1475_123b8bd8 );
buf ( n3341 , R_e63_156b1358 );
buf ( n3342 , R_1038_10085f98 );
buf ( n3343 , R_1657_13cd2c58 );
buf ( n3344 , R_844_117f3ab8 );
buf ( n3345 , R_1482_140b29d8 );
buf ( n3346 , R_a19_156ad4d8 );
buf ( n3347 , R_18f5_1587d518 );
buf ( n3348 , R_11e4_158159f8 );
buf ( n3349 , R_12d6_11c6c5d8 );
buf ( n3350 , R_1803_123b54d8 );
buf ( n3351 , R_5a6_13ccf5f8 );
buf ( n3352 , R_cb7_1162c458 );
buf ( n3353 , R_bc5_14a0c5d8 );
buf ( n3354 , R_698_14a0feb8 );
buf ( n3355 , R_194b_15882658 );
buf ( n3356 , R_d0d_1580bef8 );
buf ( n3357 , R_b6f_117eb638 );
buf ( n3358 , R_17ad_156b4f58 );
buf ( n3359 , R_132c_158823d8 );
buf ( n3360 , R_6ee_14a0faf8 );
buf ( n3361 , R_118e_156ab3b8 );
buf ( n3362 , R_75f_14870918 );
buf ( n3363 , R_173c_123b9218 );
buf ( n3364 , R_d7e_11634018 );
buf ( n3365 , R_111d_13beeb58 );
buf ( n3366 , R_139d_100868f8 );
buf ( n3367 , R_afe_15ff7ee8 );
buf ( n3368 , R_19bc_17010248 );
buf ( n3369 , R_1175_11634c98 );
buf ( n3370 , R_d26_1587cf78 );
buf ( n3371 , R_b56_13c236d8 );
buf ( n3372 , R_1345_13cd4738 );
buf ( n3373 , R_1794_15813338 );
buf ( n3374 , R_707_13d580d8 );
buf ( n3375 , R_1964_13d42b38 );
buf ( n3376 , R_f24_13b92938 );
buf ( n3377 , R_1543_15ff0828 );
buf ( n3378 , R_1596_15ff8a28 );
buf ( n3379 , R_f77_158124d8 );
buf ( n3380 , R_958_13df5bb8 );
buf ( n3381 , R_905_13d4f758 );
buf ( n3382 , R_1579_13b8d078 );
buf ( n3383 , R_f5a_15884d18 );
buf ( n3384 , R_93b_1580c3f8 );
buf ( n3385 , R_922_140af198 );
buf ( n3386 , R_f41_156b7cf8 );
buf ( n3387 , R_1560_14a14cd8 );
buf ( n3388 , R_c6c_14b20318 );
buf ( n3389 , R_64d_13ccebf8 );
buf ( n3390 , R_5f1_15814c38 );
buf ( n3391 , R_c10_15817898 );
buf ( n3392 , R_122f_13d22038 );
buf ( n3393 , R_184e_14b1b8b8 );
buf ( n3394 , R_18aa_11638b18 );
buf ( n3395 , R_128b_1587eaf8 );
buf ( n3396 , R_1695_14a12ed8 );
buf ( n3397 , R_1a63_1486ec58 );
buf ( n3398 , R_1444_15ff0788 );
buf ( n3399 , R_a57_13d5aa18 );
buf ( n3400 , R_e25_14a17078 );
buf ( n3401 , R_1076_1587b678 );
buf ( n3402 , R_806_14a0bd18 );
buf ( n3403 , R_fb7_15887158 );
buf ( n3404 , R_8c5_1008b2b8 );
buf ( n3405 , R_998_13d573b8 );
buf ( n3406 , R_ee4_15ff7da8 );
buf ( n3407 , R_1503_150daf58 );
buf ( n3408 , R_15d6_117ed398 );
buf ( n3409 , R_7ca_150de978 );
buf ( n3410 , R_a93_156af4b8 );
buf ( n3411 , R_10b2_100826b8 );
buf ( n3412 , R_16d1_156b27f8 );
buf ( n3413 , R_1a27_13cd2118 );
buf ( n3414 , R_1408_1587fbd8 );
buf ( n3415 , R_de9_13cd12b8 );
buf ( n3416 , R_9e0_15ffc9e8 );
buf ( n3417 , R_161e_123b8a98 );
buf ( n3418 , R_14bb_10081cb8 );
buf ( n3419 , R_87d_123b9498 );
buf ( n3420 , R_fff_12fbe5d8 );
buf ( n3421 , R_e9c_13df34f8 );
buf ( n3422 , R_ba8_123c12d8 );
buf ( n3423 , R_12f3_11634f18 );
buf ( n3424 , R_11c7_17013b28 );
buf ( n3425 , R_cd4_13c2b018 );
buf ( n3426 , R_589_14a19058 );
buf ( n3427 , R_1912_156aacd8 );
buf ( n3428 , R_17e6_140b2758 );
buf ( n3429 , R_6b5_1587d658 );
buf ( n3430 , R_f14_13d26458 );
buf ( n3431 , R_15a6_1162eb18 );
buf ( n3432 , R_1533_14b268f8 );
buf ( n3433 , R_f87_11637998 );
buf ( n3434 , R_968_13d2b958 );
buf ( n3435 , R_8f5_13bebe58 );
buf ( n3436 , R_8d5_150e1c18 );
buf ( n3437 , R_fa7_12fbff78 );
buf ( n3438 , R_ef4_1162ea78 );
buf ( n3439 , R_988_15814198 );
buf ( n3440 , R_1513_13c06498 );
buf ( n3441 , R_15c6_12fbf2f8 );
buf ( n3442 , R_8b7_15ffa468 );
buf ( n3443 , R_9a6_13d46058 );
buf ( n3444 , R_ed6_13d57598 );
buf ( n3445 , R_15e4_156aeb58 );
buf ( n3446 , R_14f5_13c29178 );
buf ( n3447 , R_fc5_13b8d258 );
buf ( n3448 , R_acc_13df8638 );
buf ( n3449 , R_791_13d42818 );
buf ( n3450 , R_db0_13bf9418 );
buf ( n3451 , R_13cf_123c2318 );
buf ( n3452 , R_19ee_11630cd8 );
buf ( n3453 , R_170a_13d25698 );
buf ( n3454 , R_10eb_13debbb8 );
buf ( n3455 , R_19ad_1587f9f8 );
buf ( n3456 , R_174b_15ff3528 );
buf ( n3457 , R_750_1008c9d8 );
buf ( n3458 , R_112c_13c015d8 );
buf ( n3459 , R_d6f_117eae18 );
buf ( n3460 , R_b0d_13d41c38 );
buf ( n3461 , R_138e_158113f8 );
buf ( n3462 , R_168d_156b2f78 );
buf ( n3463 , R_144c_14a0dbb8 );
buf ( n3464 , R_e2d_1587d3d8 );
buf ( n3465 , R_a4f_15814418 );
buf ( n3466 , R_80e_156ac218 );
buf ( n3467 , R_106e_14a15318 );
buf ( n3468 , R_157a_156b4198 );
buf ( n3469 , R_f5b_1162d7b8 );
buf ( n3470 , R_93c_13b933d8 );
buf ( n3471 , R_921_15813298 );
buf ( n3472 , R_f40_13cd1fd8 );
buf ( n3473 , R_155f_148745b8 );
buf ( n3474 , R_1275_13d26bd8 );
buf ( n3475 , R_c56_12fbf438 );
buf ( n3476 , R_637_14b20db8 );
buf ( n3477 , R_607_15886258 );
buf ( n3478 , R_c26_13d3ac58 );
buf ( n3479 , R_1245_13d261d8 );
buf ( n3480 , R_1864_13ddb2f8 );
buf ( n3481 , R_1894_13cd6998 );
buf ( n3482 , R_9d7_1580ac38 );
buf ( n3483 , R_1615_150e0598 );
buf ( n3484 , R_14c4_15ffa148 );
buf ( n3485 , R_886_156aa9b8 );
buf ( n3486 , R_ff6_13d424f8 );
buf ( n3487 , R_ea5_13d23b18 );
buf ( n3488 , R_1a51_13cda098 );
buf ( n3489 , R_a69_123b4f38 );
buf ( n3490 , R_1432_14b1d258 );
buf ( n3491 , R_1088_13bec3f8 );
buf ( n3492 , R_e13_140ab1d8 );
buf ( n3493 , R_16a7_156afb98 );
buf ( n3494 , R_7f4_14b238d8 );
buf ( n3495 , R_17c5_12fc1058 );
buf ( n3496 , R_b87_140b0db8 );
buf ( n3497 , R_cf5_156ab818 );
buf ( n3498 , R_1933_11633258 );
buf ( n3499 , R_11a6_13c243f8 );
buf ( n3500 , R_568_13ccd9d8 );
buf ( n3501 , R_6d6_13ccc498 );
buf ( n3502 , R_1314_13b93158 );
buf ( n3503 , R_a81_11c6b098 );
buf ( n3504 , R_10a0_148694d8 );
buf ( n3505 , R_1a39_150e4cd8 );
buf ( n3506 , R_16bf_13d3e8f8 );
buf ( n3507 , R_141a_13ccc678 );
buf ( n3508 , R_dfb_123b4c18 );
buf ( n3509 , R_7dc_14b22578 );
buf ( n3510 , R_116b_13ddcb58 );
buf ( n3511 , R_134f_14b1c7b8 );
buf ( n3512 , R_b4c_13d41eb8 );
buf ( n3513 , R_711_140b8798 );
buf ( n3514 , R_178a_13b96538 );
buf ( n3515 , R_196e_150e3658 );
buf ( n3516 , R_d30_13df5118 );
buf ( n3517 , R_b99_13df2ff8 );
buf ( n3518 , R_ce3_10088b58 );
buf ( n3519 , R_11b8_156b8798 );
buf ( n3520 , R_1921_13b91df8 );
buf ( n3521 , R_57a_13ccb818 );
buf ( n3522 , R_6c4_15887798 );
buf ( n3523 , R_17d7_11c6faf8 );
buf ( n3524 , R_1302_12fbe8f8 );
buf ( n3525 , R_65c_117f0278 );
buf ( n3526 , R_5e2_117ef198 );
buf ( n3527 , R_c01_13df0118 );
buf ( n3528 , R_18b9_13ded058 );
buf ( n3529 , R_1220_117f77f8 );
buf ( n3530 , R_129a_14a10ef8 );
buf ( n3531 , R_183f_140b7f78 );
buf ( n3532 , R_c7b_1580c178 );
buf ( n3533 , R_7bd_12fc1558 );
buf ( n3534 , R_aa0_11c6be58 );
buf ( n3535 , R_10bf_13df54d8 );
buf ( n3536 , R_16de_13de3138 );
buf ( n3537 , R_1a1a_156b8ab8 );
buf ( n3538 , R_13fb_156b4b98 );
buf ( n3539 , R_ddc_11632df8 );
buf ( n3540 , R_a7a_11c6b1d8 );
buf ( n3541 , R_1a40_140b6d58 );
buf ( n3542 , R_1099_116354b8 );
buf ( n3543 , R_1421_117ef7d8 );
buf ( n3544 , R_16b8_13d3ea38 );
buf ( n3545 , R_e02_15ff37a8 );
buf ( n3546 , R_7e3_15812118 );
buf ( n3547 , R_1a56_13bf0818 );
buf ( n3548 , R_1437_123bad98 );
buf ( n3549 , R_a64_13beb318 );
buf ( n3550 , R_e18_156afc38 );
buf ( n3551 , R_1083_123c0a18 );
buf ( n3552 , R_7f9_156b30b8 );
buf ( n3553 , R_16a2_150e9418 );
buf ( n3554 , R_18e0_13c201b8 );
buf ( n3555 , R_1818_140b47d8 );
buf ( n3556 , R_12c1_123bb838 );
buf ( n3557 , R_5bb_156b5638 );
buf ( n3558 , R_ca2_13dd9d18 );
buf ( n3559 , R_bda_13b985b8 );
buf ( n3560 , R_683_11634478 );
buf ( n3561 , R_11f9_13ccd938 );
buf ( n3562 , R_157b_1486f0b8 );
buf ( n3563 , R_f5c_13de2378 );
buf ( n3564 , R_93d_117f0ef8 );
buf ( n3565 , R_920_13df90d8 );
buf ( n3566 , R_f3f_13bf1a38 );
buf ( n3567 , R_155e_123c0d38 );
buf ( n3568 , R_8de_13d4e0d8 );
buf ( n3569 , R_f9e_13b8a738 );
buf ( n3570 , R_efd_123bfed8 );
buf ( n3571 , R_97f_123c21d8 );
buf ( n3572 , R_151c_13d5c4f8 );
buf ( n3573 , R_15bd_13df43f8 );
buf ( n3574 , R_1763_13d44618 );
buf ( n3575 , R_1995_17017548 );
buf ( n3576 , R_1144_17018948 );
buf ( n3577 , R_738_1700bce8 );
buf ( n3578 , R_b25_1162ad38 );
buf ( n3579 , R_d57_13c242b8 );
buf ( n3580 , R_1376_117f5098 );
buf ( n3581 , R_9be_140aaaf8 );
buf ( n3582 , R_89f_156b2ed8 );
buf ( n3583 , R_15fc_13c28db8 );
buf ( n3584 , R_ebe_13cd5c78 );
buf ( n3585 , R_fdd_1162dd58 );
buf ( n3586 , R_14dd_123b8db8 );
buf ( n3587 , R_14aa_13c0f9f8 );
buf ( n3588 , R_86c_13df77d8 );
buf ( n3589 , R_1010_15884278 );
buf ( n3590 , R_e8b_15880ad8 );
buf ( n3591 , R_162f_15ff7808 );
buf ( n3592 , R_9f1_123be718 );
buf ( n3593 , R_1457_13d54758 );
buf ( n3594 , R_1682_1587fb38 );
buf ( n3595 , R_e38_150debf8 );
buf ( n3596 , R_a44_1580d618 );
buf ( n3597 , R_819_14873898 );
buf ( n3598 , R_1063_13cd8978 );
buf ( n3599 , R_1a4c_156b8b58 );
buf ( n3600 , R_a6e_117ec3f8 );
buf ( n3601 , R_142d_14b1c998 );
buf ( n3602 , R_108d_14a0a878 );
buf ( n3603 , R_e0e_156b9f58 );
buf ( n3604 , R_16ac_13bf1218 );
buf ( n3605 , R_7ef_1700c788 );
buf ( n3606 , R_1014_13c079d8 );
buf ( n3607 , R_868_1587de78 );
buf ( n3608 , R_14a6_10081998 );
buf ( n3609 , R_1633_117e9ab8 );
buf ( n3610 , R_9f5_13d25c38 );
buf ( n3611 , R_e87_15ff9ce8 );
buf ( n3612 , R_1829_123b40d8 );
buf ( n3613 , R_18cf_13ded238 );
buf ( n3614 , R_5cc_156aa698 );
buf ( n3615 , R_12b0_14a177f8 );
buf ( n3616 , R_beb_13cca738 );
buf ( n3617 , R_c91_15ff1cc8 );
buf ( n3618 , R_120a_13cd9738 );
buf ( n3619 , R_672_13c06fd8 );
buf ( n3620 , R_779_13cd2258 );
buf ( n3621 , R_d98_13b958b8 );
buf ( n3622 , R_13b7_1700e308 );
buf ( n3623 , R_19d6_117ecfd8 );
buf ( n3624 , R_1722_123b5a78 );
buf ( n3625 , R_1103_117f7bb8 );
buf ( n3626 , R_ae4_11634ab8 );
buf ( n3627 , R_c57_15814f58 );
buf ( n3628 , R_638_14a151d8 );
buf ( n3629 , R_606_13d50838 );
buf ( n3630 , R_c25_10083bf8 );
buf ( n3631 , R_1244_13ddb898 );
buf ( n3632 , R_1863_123b9f38 );
buf ( n3633 , R_1895_13df3a98 );
buf ( n3634 , R_1276_123bda98 );
buf ( n3635 , R_1042_13cd6718 );
buf ( n3636 , R_e59_1587dd38 );
buf ( n3637 , R_1661_13de0758 );
buf ( n3638 , R_83a_13d21598 );
buf ( n3639 , R_a23_14869cf8 );
buf ( n3640 , R_1478_13cd7618 );
buf ( n3641 , R_668_11c6aff8 );
buf ( n3642 , R_5d6_13d24158 );
buf ( n3643 , R_18c5_123b5f78 );
buf ( n3644 , R_bf5_123ba7f8 );
buf ( n3645 , R_12a6_148674f8 );
buf ( n3646 , R_1214_15886cf8 );
buf ( n3647 , R_c87_13c21bf8 );
buf ( n3648 , R_1833_117f3838 );
buf ( n3649 , R_1820_14872a38 );
buf ( n3650 , R_18d8_13b8ef18 );
buf ( n3651 , R_5c3_10080778 );
buf ( n3652 , R_12b9_140abb38 );
buf ( n3653 , R_be2_13b98338 );
buf ( n3654 , R_c9a_13cd1f38 );
buf ( n3655 , R_1201_15ff65e8 );
buf ( n3656 , R_67b_13c02bb8 );
buf ( n3657 , R_1542_14a19cd8 );
buf ( n3658 , R_1597_117ee478 );
buf ( n3659 , R_f78_156af198 );
buf ( n3660 , R_959_11631bd8 );
buf ( n3661 , R_904_13bebbd8 );
buf ( n3662 , R_f23_13c2b338 );
buf ( n3663 , R_157c_14a0eab8 );
buf ( n3664 , R_f5d_15817c58 );
buf ( n3665 , R_93e_13cd6858 );
buf ( n3666 , R_91f_117f7d98 );
buf ( n3667 , R_f3e_1700a708 );
buf ( n3668 , R_155d_1700fa28 );
buf ( n3669 , R_764_150dee78 );
buf ( n3670 , R_1737_13cd6538 );
buf ( n3671 , R_d83_150dc678 );
buf ( n3672 , R_1118_13cce3d8 );
buf ( n3673 , R_13a2_13df95d8 );
buf ( n3674 , R_af9_14b1bc78 );
buf ( n3675 , R_19c1_15811358 );
buf ( n3676 , R_14ae_14b22438 );
buf ( n3677 , R_870_158800d8 );
buf ( n3678 , R_100c_14b1bef8 );
buf ( n3679 , R_e8f_13c27cd8 );
buf ( n3680 , R_9ed_150e3a18 );
buf ( n3681 , R_162b_13d24478 );
buf ( n3682 , R_64e_12fbeb78 );
buf ( n3683 , R_5f0_13d25738 );
buf ( n3684 , R_c0f_1587ef58 );
buf ( n3685 , R_122e_14a181f8 );
buf ( n3686 , R_184d_1486ac98 );
buf ( n3687 , R_18ab_13bf9d78 );
buf ( n3688 , R_128c_11c6a378 );
buf ( n3689 , R_c6d_13d3be78 );
buf ( n3690 , R_d11_117f09f8 );
buf ( n3691 , R_b6b_13c0e878 );
buf ( n3692 , R_17a9_15ff62c8 );
buf ( n3693 , R_1330_1580d6b8 );
buf ( n3694 , R_6f2_123ba398 );
buf ( n3695 , R_118a_13c1eef8 );
buf ( n3696 , R_194f_13c0e738 );
buf ( n3697 , R_1758_14a14eb8 );
buf ( n3698 , R_19a0_13c204d8 );
buf ( n3699 , R_1139_117ef878 );
buf ( n3700 , R_743_13d5a478 );
buf ( n3701 , R_b1a_13c01038 );
buf ( n3702 , R_d62_15811df8 );
buf ( n3703 , R_1381_123b3a98 );
buf ( n3704 , R_e6d_123b7238 );
buf ( n3705 , R_102e_150ddd98 );
buf ( n3706 , R_84e_15883418 );
buf ( n3707 , R_164d_14a0c678 );
buf ( n3708 , R_148c_1580e8d8 );
buf ( n3709 , R_a0f_15ffbae8 );
buf ( n3710 , R_12ee_13d3d958 );
buf ( n3711 , R_11cc_14a11a38 );
buf ( n3712 , R_ccf_15812258 );
buf ( n3713 , R_58e_150e4558 );
buf ( n3714 , R_17eb_150e6538 );
buf ( n3715 , R_190d_14b294b8 );
buf ( n3716 , R_6b0_14a172f8 );
buf ( n3717 , R_bad_15883c38 );
buf ( n3718 , R_1018_13d2a878 );
buf ( n3719 , R_864_13c09238 );
buf ( n3720 , R_14a2_13cd9e18 );
buf ( n3721 , R_1637_1162fbf8 );
buf ( n3722 , R_9f9_156b7438 );
buf ( n3723 , R_e83_15886438 );
buf ( n3724 , R_1a5b_13df6158 );
buf ( n3725 , R_143c_15ff2a88 );
buf ( n3726 , R_a5f_13df1518 );
buf ( n3727 , R_e1d_13c288b8 );
buf ( n3728 , R_107e_13c1c298 );
buf ( n3729 , R_7fe_117f30b8 );
buf ( n3730 , R_169d_156abf98 );
buf ( n3731 , R_15b3_13cd6e98 );
buf ( n3732 , R_f07_13b953b8 );
buf ( n3733 , R_f94_13d25198 );
buf ( n3734 , R_1526_1486bf58 );
buf ( n3735 , R_975_13d529f8 );
buf ( n3736 , R_8e8_117f0bd8 );
buf ( n3737 , R_78f_1162c9f8 );
buf ( n3738 , R_dae_11c6d578 );
buf ( n3739 , R_13cd_14a162b8 );
buf ( n3740 , R_19ec_15814738 );
buf ( n3741 , R_170c_13ccdd98 );
buf ( n3742 , R_10ed_15882dd8 );
buf ( n3743 , R_ace_15885cb8 );
buf ( n3744 , R_157d_13cd56d8 );
buf ( n3745 , R_f5e_140b53b8 );
buf ( n3746 , R_93f_13d57778 );
buf ( n3747 , R_91e_15886f78 );
buf ( n3748 , R_f3d_11634798 );
buf ( n3749 , R_155c_156adf78 );
buf ( n3750 , R_782_15ffd168 );
buf ( n3751 , R_da1_14b290f8 );
buf ( n3752 , R_13c0_117f6b78 );
buf ( n3753 , R_19df_117eb318 );
buf ( n3754 , R_1719_13c1f8f8 );
buf ( n3755 , R_10fa_13decd38 );
buf ( n3756 , R_adb_17014708 );
buf ( n3757 , R_a88_13cd40f8 );
buf ( n3758 , R_10a7_117eb1d8 );
buf ( n3759 , R_16c6_158880f8 );
buf ( n3760 , R_1a32_15818018 );
buf ( n3761 , R_1413_13d57ef8 );
buf ( n3762 , R_df4_17013f88 );
buf ( n3763 , R_7d5_15889098 );
buf ( n3764 , R_639_13df0cf8 );
buf ( n3765 , R_605_14b1c3f8 );
buf ( n3766 , R_c24_11632d58 );
buf ( n3767 , R_1243_158151d8 );
buf ( n3768 , R_1862_140b94b8 );
buf ( n3769 , R_1896_13c0a598 );
buf ( n3770 , R_1277_13c27378 );
buf ( n3771 , R_c58_13dddc38 );
buf ( n3772 , R_15a7_17013448 );
buf ( n3773 , R_1532_156b4ff8 );
buf ( n3774 , R_f88_13d225d8 );
buf ( n3775 , R_969_13cce298 );
buf ( n3776 , R_8f4_156b9af8 );
buf ( n3777 , R_f13_13c2b478 );
buf ( n3778 , R_1750_14a13018 );
buf ( n3779 , R_74b_123b9998 );
buf ( n3780 , R_1131_13d21c78 );
buf ( n3781 , R_d6a_13c0c118 );
buf ( n3782 , R_b12_1587bb78 );
buf ( n3783 , R_1389_13c2a4d8 );
buf ( n3784 , R_19a8_124c5578 );
buf ( n3785 , R_a9e_13de43f8 );
buf ( n3786 , R_10bd_1162e6b8 );
buf ( n3787 , R_16dc_14b1f058 );
buf ( n3788 , R_1a1c_13cda138 );
buf ( n3789 , R_13fd_14a0e0b8 );
buf ( n3790 , R_dde_15ffc448 );
buf ( n3791 , R_7bf_123bb0b8 );
buf ( n3792 , R_1027_13c277d8 );
buf ( n3793 , R_855_14a117b8 );
buf ( n3794 , R_1493_13bee3d8 );
buf ( n3795 , R_1646_13ccbdb8 );
buf ( n3796 , R_a08_15ffa5a8 );
buf ( n3797 , R_e74_123b4678 );
buf ( n3798 , R_12d0_14a11cb8 );
buf ( n3799 , R_1809_13d4f7f8 );
buf ( n3800 , R_5ac_11c6e838 );
buf ( n3801 , R_cb1_13d2c998 );
buf ( n3802 , R_bcb_1007e3d8 );
buf ( n3803 , R_692_1587be98 );
buf ( n3804 , R_18ef_13d28758 );
buf ( n3805 , R_11ea_1580f238 );
buf ( n3806 , R_991_1007ff58 );
buf ( n3807 , R_eeb_12fbe0d8 );
buf ( n3808 , R_150a_14a0b3b8 );
buf ( n3809 , R_15cf_10085958 );
buf ( n3810 , R_fb0_117f5318 );
buf ( n3811 , R_8cc_13bf3338 );
buf ( n3812 , R_ce8_11c6a7d8 );
buf ( n3813 , R_1926_116372b8 );
buf ( n3814 , R_11b3_13cd3fb8 );
buf ( n3815 , R_575_15817438 );
buf ( n3816 , R_6c9_13dee318 );
buf ( n3817 , R_1307_15ff2da8 );
buf ( n3818 , R_17d2_156b8978 );
buf ( n3819 , R_b94_1587e198 );
buf ( n3820 , R_1810_117f12b8 );
buf ( n3821 , R_12c9_17017868 );
buf ( n3822 , R_5b3_123baa78 );
buf ( n3823 , R_caa_15fedbc8 );
buf ( n3824 , R_bd2_1580d9d8 );
buf ( n3825 , R_68b_13ddf038 );
buf ( n3826 , R_11f1_13c2a938 );
buf ( n3827 , R_18e8_123bd638 );
buf ( n3828 , R_157e_13dee278 );
buf ( n3829 , R_f5f_1162d038 );
buf ( n3830 , R_940_1486f838 );
buf ( n3831 , R_91d_14b1cdf8 );
buf ( n3832 , R_f3c_148682b8 );
buf ( n3833 , R_155b_12fc0158 );
buf ( n3834 , R_14b2_15ff2628 );
buf ( n3835 , R_874_123c0298 );
buf ( n3836 , R_1008_1587dc98 );
buf ( n3837 , R_e93_13cd4878 );
buf ( n3838 , R_9e9_123b4498 );
buf ( n3839 , R_1627_156b7578 );
buf ( n3840 , R_cf1_124c34f8 );
buf ( n3841 , R_192f_14a12cf8 );
buf ( n3842 , R_11aa_117e9bf8 );
buf ( n3843 , R_56c_140ab598 );
buf ( n3844 , R_6d2_1162ec58 );
buf ( n3845 , R_1310_13ddf538 );
buf ( n3846 , R_17c9_11638578 );
buf ( n3847 , R_b8b_13df36d8 );
buf ( n3848 , R_a91_13ccfeb8 );
buf ( n3849 , R_10b0_117ea418 );
buf ( n3850 , R_16cf_11c6b138 );
buf ( n3851 , R_1a29_13d384f8 );
buf ( n3852 , R_140a_140aa5f8 );
buf ( n3853 , R_deb_140b71b8 );
buf ( n3854 , R_7cc_13cd94b8 );
buf ( n3855 , R_1a47_100862b8 );
buf ( n3856 , R_a73_123be538 );
buf ( n3857 , R_1428_13dde3b8 );
buf ( n3858 , R_1092_15ff41a8 );
buf ( n3859 , R_e09_15887a18 );
buf ( n3860 , R_16b1_13c0c258 );
buf ( n3861 , R_7ea_11c6e518 );
buf ( n3862 , R_e66_170138a8 );
buf ( n3863 , R_1035_1162a478 );
buf ( n3864 , R_847_14a15a98 );
buf ( n3865 , R_1654_1580fff8 );
buf ( n3866 , R_1485_117f6358 );
buf ( n3867 , R_a16_14b25638 );
buf ( n3868 , R_b60_13b97b18 );
buf ( n3869 , R_179e_156b3c98 );
buf ( n3870 , R_133b_13ddde18 );
buf ( n3871 , R_6fd_156b8338 );
buf ( n3872 , R_117f_13cd7578 );
buf ( n3873 , R_195a_150e1218 );
buf ( n3874 , R_d1c_13d3fd98 );
buf ( n3875 , R_134c_14a11ad8 );
buf ( n3876 , R_b4f_12fbee98 );
buf ( n3877 , R_70e_124c25f8 );
buf ( n3878 , R_178d_11638a78 );
buf ( n3879 , R_196b_1580a918 );
buf ( n3880 , R_d2d_13cd54f8 );
buf ( n3881 , R_116e_117ebb38 );
buf ( n3882 , R_5e1_14b286f8 );
buf ( n3883 , R_c00_150df558 );
buf ( n3884 , R_18ba_11638bb8 );
buf ( n3885 , R_121f_13dfa1b8 );
buf ( n3886 , R_129b_13cd3298 );
buf ( n3887 , R_183e_1587c398 );
buf ( n3888 , R_c7c_11c6a558 );
buf ( n3889 , R_65d_13cd74d8 );
buf ( n3890 , R_9b3_13df8138 );
buf ( n3891 , R_8aa_13dd9a98 );
buf ( n3892 , R_15f1_156b5d18 );
buf ( n3893 , R_ec9_1587c1b8 );
buf ( n3894 , R_fd2_13c05098 );
buf ( n3895 , R_14e8_1700a528 );
buf ( n3896 , R_11dd_14875918 );
buf ( n3897 , R_12dd_14a0e158 );
buf ( n3898 , R_17fc_11635eb8 );
buf ( n3899 , R_59f_14a14c38 );
buf ( n3900 , R_cbe_116357d8 );
buf ( n3901 , R_bbe_15881438 );
buf ( n3902 , R_18fc_17009bc8 );
buf ( n3903 , R_69f_13d56b98 );
buf ( n3904 , R_1598_13cd92d8 );
buf ( n3905 , R_f79_13bf2e38 );
buf ( n3906 , R_95a_13d37698 );
buf ( n3907 , R_903_117ec7b8 );
buf ( n3908 , R_f22_14a13978 );
buf ( n3909 , R_1541_15886758 );
buf ( n3910 , R_12e3_17014028 );
buf ( n3911 , R_11d7_1587d5b8 );
buf ( n3912 , R_cc4_13bead78 );
buf ( n3913 , R_599_150dcf38 );
buf ( n3914 , R_17f6_117f1498 );
buf ( n3915 , R_1902_14b1af58 );
buf ( n3916 , R_6a5_13df56b8 );
buf ( n3917 , R_bb8_124c3b38 );
buf ( n3918 , R_14bf_150dd938 );
buf ( n3919 , R_881_150db278 );
buf ( n3920 , R_ffb_15813ab8 );
buf ( n3921 , R_ea0_13b95778 );
buf ( n3922 , R_9dc_15ff19a8 );
buf ( n3923 , R_161a_14b23bf8 );
buf ( n3924 , R_1454_123b4538 );
buf ( n3925 , R_e35_11c70098 );
buf ( n3926 , R_a47_1486f3d8 );
buf ( n3927 , R_816_13c06cb8 );
buf ( n3928 , R_1066_13bee838 );
buf ( n3929 , R_1685_15ff1d68 );
buf ( n3930 , R_8b0_15813c98 );
buf ( n3931 , R_9ad_13de0bb8 );
buf ( n3932 , R_ecf_13c26798 );
buf ( n3933 , R_15eb_140b6498 );
buf ( n3934 , R_14ee_13d5a298 );
buf ( n3935 , R_fcc_150e33d8 );
buf ( n3936 , R_101c_11c6ce98 );
buf ( n3937 , R_860_14a17b18 );
buf ( n3938 , R_149e_11c6edd8 );
buf ( n3939 , R_163b_13c04b98 );
buf ( n3940 , R_9fd_117ebf98 );
buf ( n3941 , R_e7f_117f6038 );
buf ( n3942 , R_604_15811718 );
buf ( n3943 , R_c23_123bfc58 );
buf ( n3944 , R_1242_10080c78 );
buf ( n3945 , R_1861_12fbf7f8 );
buf ( n3946 , R_1897_13d3d1d8 );
buf ( n3947 , R_1278_117f4f58 );
buf ( n3948 , R_c59_116304b8 );
buf ( n3949 , R_63a_13c0a278 );
buf ( n3950 , R_b59_15feff68 );
buf ( n3951 , R_1342_148716d8 );
buf ( n3952 , R_1797_117f7e38 );
buf ( n3953 , R_704_123b2ff8 );
buf ( n3954 , R_1961_1162de98 );
buf ( n3955 , R_1178_13cd24d8 );
buf ( n3956 , R_d23_11c68618 );
buf ( n3957 , R_157f_13b8ce98 );
buf ( n3958 , R_f60_140af9b8 );
buf ( n3959 , R_941_13df8b38 );
buf ( n3960 , R_91c_13df6d38 );
buf ( n3961 , R_f3b_15810c78 );
buf ( n3962 , R_155a_15882338 );
buf ( n3963 , R_e5c_117f6df8 );
buf ( n3964 , R_165e_117edf78 );
buf ( n3965 , R_83d_13c24ad8 );
buf ( n3966 , R_a20_15883738 );
buf ( n3967 , R_147b_1700f5c8 );
buf ( n3968 , R_103f_123b9ad8 );
buf ( n3969 , R_5ef_1162a018 );
buf ( n3970 , R_c0e_158802b8 );
buf ( n3971 , R_122d_150e4eb8 );
buf ( n3972 , R_184c_14a19418 );
buf ( n3973 , R_18ac_117f13f8 );
buf ( n3974 , R_128d_123b2af8 );
buf ( n3975 , R_c6e_15ff6408 );
buf ( n3976 , R_64f_13bf1ad8 );
buf ( n3977 , R_9a0_13dd6078 );
buf ( n3978 , R_edc_123be678 );
buf ( n3979 , R_15de_15ff2268 );
buf ( n3980 , R_14fb_13c29038 );
buf ( n3981 , R_fbf_150e4f58 );
buf ( n3982 , R_8bd_13cd5ef8 );
buf ( n3983 , R_1998_14b279d8 );
buf ( n3984 , R_1141_1580bbd8 );
buf ( n3985 , R_73b_14a15638 );
buf ( n3986 , R_b22_13cce8d8 );
buf ( n3987 , R_d5a_13bf6178 );
buf ( n3988 , R_1379_123bdbd8 );
buf ( n3989 , R_1760_117f7f78 );
buf ( n3990 , R_1981_1587b7b8 );
buf ( n3991 , R_b39_15ffae68 );
buf ( n3992 , R_724_117ec8f8 );
buf ( n3993 , R_1777_1587ccf8 );
buf ( n3994 , R_d43_13beedd8 );
buf ( n3995 , R_1362_150dfcd8 );
buf ( n3996 , R_1158_13bf0f98 );
buf ( n3997 , R_770_15888058 );
buf ( n3998 , R_d8f_11629f78 );
buf ( n3999 , R_13ae_13bf3478 );
buf ( n4000 , R_172b_156b88d8 );
buf ( n4001 , R_19cd_117ed578 );
buf ( n4002 , R_110c_15810458 );
buf ( n4003 , R_aed_14a0e298 );
buf ( n4004 , R_1449_14b26678 );
buf ( n4005 , R_e2a_13c29858 );
buf ( n4006 , R_a52_140af378 );
buf ( n4007 , R_80b_158154f8 );
buf ( n4008 , R_1071_123c1378 );
buf ( n4009 , R_1a68_117ed618 );
buf ( n4010 , R_1690_13c216f8 );
buf ( n4011 , R_ef3_13cd06d8 );
buf ( n4012 , R_989_13c068f8 );
buf ( n4013 , R_1512_1162e078 );
buf ( n4014 , R_15c7_13d3c4b8 );
buf ( n4015 , R_8d4_123c1738 );
buf ( n4016 , R_fa8_123be858 );
buf ( n4017 , R_1984_1162e438 );
buf ( n4018 , R_727_1700aca8 );
buf ( n4019 , R_b36_123bb338 );
buf ( n4020 , R_d46_13cd3338 );
buf ( n4021 , R_1774_13c26c98 );
buf ( n4022 , R_1365_150db818 );
buf ( n4023 , R_1155_17012868 );
buf ( n4024 , R_b3c_13cd4eb8 );
buf ( n4025 , R_721_156b7d98 );
buf ( n4026 , R_197e_13d5c8b8 );
buf ( n4027 , R_177a_123c1418 );
buf ( n4028 , R_d40_11635af8 );
buf ( n4029 , R_115b_123bf2f8 );
buf ( n4030 , R_135f_11c6da78 );
buf ( n4031 , R_894_1587b2b8 );
buf ( n4032 , R_1607_123bd138 );
buf ( n4033 , R_eb3_123b5cf8 );
buf ( n4034 , R_fe8_15816678 );
buf ( n4035 , R_14d2_11636e58 );
buf ( n4036 , R_9c9_13cce798 );
buf ( n4037 , R_160c_117f74d8 );
buf ( n4038 , R_88f_13c0d338 );
buf ( n4039 , R_fed_12fc1198 );
buf ( n4040 , R_eae_13cd1d58 );
buf ( n4041 , R_9ce_1162c6d8 );
buf ( n4042 , R_14cd_10081178 );
buf ( n4043 , R_dac_14a109f8 );
buf ( n4044 , R_13cb_13ccf0f8 );
buf ( n4045 , R_19ea_11629b18 );
buf ( n4046 , R_170e_1580e338 );
buf ( n4047 , R_10ef_14a199b8 );
buf ( n4048 , R_ad0_123b65b8 );
buf ( n4049 , R_78d_15817618 );
buf ( n4050 , R_999_1008a138 );
buf ( n4051 , R_ee3_158135b8 );
buf ( n4052 , R_1502_117ea238 );
buf ( n4053 , R_15d7_11c6ab98 );
buf ( n4054 , R_fb8_156b7bb8 );
buf ( n4055 , R_8c4_117f8018 );
buf ( n4056 , R_efc_12fc14b8 );
buf ( n4057 , R_980_13d2b9f8 );
buf ( n4058 , R_151b_14a153b8 );
buf ( n4059 , R_15be_11629bb8 );
buf ( n4060 , R_8dd_13d1dcb8 );
buf ( n4061 , R_f9f_13bf1858 );
buf ( n4062 , R_8a4_13cd4418 );
buf ( n4063 , R_15f7_117ea878 );
buf ( n4064 , R_ec3_14a15e58 );
buf ( n4065 , R_fd8_117f1718 );
buf ( n4066 , R_14e2_13ddc478 );
buf ( n4067 , R_9b9_1008a458 );
buf ( n4068 , R_1580_123b3958 );
buf ( n4069 , R_f61_14867318 );
buf ( n4070 , R_942_140b3a18 );
buf ( n4071 , R_91b_156b0d18 );
buf ( n4072 , R_f3a_1007f4b8 );
buf ( n4073 , R_1559_13c234f8 );
buf ( n4074 , R_1441_13ded378 );
buf ( n4075 , R_a5a_13c097d8 );
buf ( n4076 , R_e22_117eccb8 );
buf ( n4077 , R_1079_13beb6d8 );
buf ( n4078 , R_803_140b8158 );
buf ( n4079 , R_1698_15811998 );
buf ( n4080 , R_1a60_14b1b778 );
buf ( n4081 , R_1987_140b7cf8 );
buf ( n4082 , R_72a_158127f8 );
buf ( n4083 , R_b33_13d2aaf8 );
buf ( n4084 , R_d49_15811678 );
buf ( n4085 , R_1771_17009c68 );
buf ( n4086 , R_1368_1587e9b8 );
buf ( n4087 , R_1152_13c0bd58 );
buf ( n4088 , R_5d5_123be038 );
buf ( n4089 , R_18c6_13d3a1b8 );
buf ( n4090 , R_bf4_1587cb18 );
buf ( n4091 , R_12a7_15817cf8 );
buf ( n4092 , R_1213_140ad078 );
buf ( n4093 , R_c88_17017cc8 );
buf ( n4094 , R_1832_123bc2d8 );
buf ( n4095 , R_669_116322b8 );
buf ( n4096 , R_769_150da558 );
buf ( n4097 , R_d88_117f22f8 );
buf ( n4098 , R_1732_123b2558 );
buf ( n4099 , R_13a7_13c08ab8 );
buf ( n4100 , R_1113_123c1e18 );
buf ( n4101 , R_19c6_13cd18f8 );
buf ( n4102 , R_af4_1580feb8 );
buf ( n4103 , R_b3f_13c22198 );
buf ( n4104 , R_71e_140aec98 );
buf ( n4105 , R_197b_123c14b8 );
buf ( n4106 , R_177d_17012728 );
buf ( n4107 , R_d3d_13c053b8 );
buf ( n4108 , R_115e_15885c18 );
buf ( n4109 , R_135c_13cda3b8 );
buf ( n4110 , R_12d7_13cd2578 );
buf ( n4111 , R_1802_13d3fbb8 );
buf ( n4112 , R_5a5_13d375f8 );
buf ( n4113 , R_cb8_11c6c218 );
buf ( n4114 , R_bc4_14b2a138 );
buf ( n4115 , R_699_15888ff8 );
buf ( n4116 , R_18f6_124c27d8 );
buf ( n4117 , R_11e3_1162fa18 );
buf ( n4118 , R_b67_13cd4f58 );
buf ( n4119 , R_17a5_116334d8 );
buf ( n4120 , R_1334_13cd5598 );
buf ( n4121 , R_6f6_117f1858 );
buf ( n4122 , R_1186_11635d78 );
buf ( n4123 , R_1953_117eb6d8 );
buf ( n4124 , R_d15_123b5578 );
buf ( n4125 , R_603_13ddbe38 );
buf ( n4126 , R_c22_117f71b8 );
buf ( n4127 , R_1241_1162a5b8 );
buf ( n4128 , R_1860_13ccdf78 );
buf ( n4129 , R_1898_11c6bb38 );
buf ( n4130 , R_1279_15887478 );
buf ( n4131 , R_c5a_14a16538 );
buf ( n4132 , R_63b_15883cd8 );
buf ( n4133 , R_10bb_1587d8d8 );
buf ( n4134 , R_16da_124c3db8 );
buf ( n4135 , R_1a1e_11c6ed38 );
buf ( n4136 , R_13ff_17012c28 );
buf ( n4137 , R_de0_13d3abb8 );
buf ( n4138 , R_7c1_156b3bf8 );
buf ( n4139 , R_a9c_1162e4d8 );
buf ( n4140 , R_18d0_117f1358 );
buf ( n4141 , R_5cb_12fc0d38 );
buf ( n4142 , R_12b1_124c38b8 );
buf ( n4143 , R_bea_13ccb098 );
buf ( n4144 , R_c92_150e3838 );
buf ( n4145 , R_1209_14a0aa58 );
buf ( n4146 , R_673_14a13fb8 );
buf ( n4147 , R_1828_1580ab98 );
buf ( n4148 , R_14b6_1587d1f8 );
buf ( n4149 , R_878_13c100d8 );
buf ( n4150 , R_1004_156ab318 );
buf ( n4151 , R_e97_14866918 );
buf ( n4152 , R_9e5_1587d6f8 );
buf ( n4153 , R_1623_13b96178 );
buf ( n4154 , R_11d1_1162f6f8 );
buf ( n4155 , R_cca_117eebf8 );
buf ( n4156 , R_593_117ee0b8 );
buf ( n4157 , R_17f0_100833d8 );
buf ( n4158 , R_1908_1162f5b8 );
buf ( n4159 , R_6ab_13ccbe58 );
buf ( n4160 , R_bb2_15810278 );
buf ( n4161 , R_12e9_13d26818 );
buf ( n4162 , R_f89_13d51738 );
buf ( n4163 , R_96a_1587c258 );
buf ( n4164 , R_8f3_10082b18 );
buf ( n4165 , R_f12_1162b2d8 );
buf ( n4166 , R_15a8_14b25db8 );
buf ( n4167 , R_1531_13c0ac78 );
buf ( n4168 , R_12c2_13d4e2b8 );
buf ( n4169 , R_5ba_13b94d78 );
buf ( n4170 , R_ca3_13ddaa38 );
buf ( n4171 , R_bd9_13d54398 );
buf ( n4172 , R_684_117f5a98 );
buf ( n4173 , R_11f8_13bf1538 );
buf ( n4174 , R_18e1_17010388 );
buf ( n4175 , R_1817_1580f9b8 );
buf ( n4176 , R_a7f_117ebc78 );
buf ( n4177 , R_1a3b_13d275d8 );
buf ( n4178 , R_109e_14a11538 );
buf ( n4179 , R_16bd_117eb9f8 );
buf ( n4180 , R_141c_123b3f98 );
buf ( n4181 , R_dfd_1700cf08 );
buf ( n4182 , R_7de_15881ed8 );
buf ( n4183 , R_f95_13d51058 );
buf ( n4184 , R_1525_140b5598 );
buf ( n4185 , R_976_140b2f78 );
buf ( n4186 , R_8e7_13dd8ff8 );
buf ( n4187 , R_15b4_13dee598 );
buf ( n4188 , R_f06_14b29238 );
buf ( n4189 , R_899_13d5a8d8 );
buf ( n4190 , R_1602_13c28ef8 );
buf ( n4191 , R_eb8_13c1c0b8 );
buf ( n4192 , R_fe3_13ccb598 );
buf ( n4193 , R_14d7_14a0fb98 );
buf ( n4194 , R_9c4_123c1a58 );
buf ( n4195 , R_1599_13bf40f8 );
buf ( n4196 , R_f7a_13d510f8 );
buf ( n4197 , R_95b_15813838 );
buf ( n4198 , R_902_14a0aff8 );
buf ( n4199 , R_f21_15812398 );
buf ( n4200 , R_1540_14871458 );
buf ( n4201 , R_1321_156b1038 );
buf ( n4202 , R_1199_13cd3bf8 );
buf ( n4203 , R_6e3_140b27f8 );
buf ( n4204 , R_55b_13d54f78 );
buf ( n4205 , R_1940_117ed758 );
buf ( n4206 , R_17b8_14b1ca38 );
buf ( n4207 , R_d02_14b21998 );
buf ( n4208 , R_b7a_140b8298 );
buf ( n4209 , R_ed5_123b27d8 );
buf ( n4210 , R_15e5_13d3e0d8 );
buf ( n4211 , R_14f4_1580cad8 );
buf ( n4212 , R_fc6_117f2078 );
buf ( n4213 , R_8b6_12fbe7b8 );
buf ( n4214 , R_9a7_13dd6118 );
buf ( n4215 , R_d96_13c23778 );
buf ( n4216 , R_13b5_124c31d8 );
buf ( n4217 , R_19d4_123b6798 );
buf ( n4218 , R_1724_117edcf8 );
buf ( n4219 , R_1105_158130b8 );
buf ( n4220 , R_ae6_14873e38 );
buf ( n4221 , R_777_17012228 );
buf ( n4222 , R_1581_10080458 );
buf ( n4223 , R_f62_13ccaff8 );
buf ( n4224 , R_943_156b21b8 );
buf ( n4225 , R_91a_13d23e38 );
buf ( n4226 , R_f39_117f5778 );
buf ( n4227 , R_1558_15ffb2c8 );
buf ( n4228 , R_88a_15880c18 );
buf ( n4229 , R_ff2_13d42638 );
buf ( n4230 , R_ea9_15810ef8 );
buf ( n4231 , R_9d3_12fc1e18 );
buf ( n4232 , R_14c8_13d50d38 );
buf ( n4233 , R_1611_13df2b98 );
buf ( n4234 , R_5c2_150db138 );
buf ( n4235 , R_12ba_158138d8 );
buf ( n4236 , R_be1_10082898 );
buf ( n4237 , R_c9b_13b977f8 );
buf ( n4238 , R_1200_13d3d778 );
buf ( n4239 , R_67c_13dec978 );
buf ( n4240 , R_181f_156b4558 );
buf ( n4241 , R_18d9_117f3e78 );
buf ( n4242 , R_1743_15ff3488 );
buf ( n4243 , R_758_13cd0ef8 );
buf ( n4244 , R_1124_14a17d98 );
buf ( n4245 , R_d77_14a0ca38 );
buf ( n4246 , R_1396_156ace98 );
buf ( n4247 , R_b05_13d37d78 );
buf ( n4248 , R_19b5_13cd3c98 );
buf ( n4249 , R_d9f_1580b818 );
buf ( n4250 , R_13be_156af5f8 );
buf ( n4251 , R_19dd_13d56238 );
buf ( n4252 , R_171b_14a0ac38 );
buf ( n4253 , R_10fc_13d52c78 );
buf ( n4254 , R_add_17015ce8 );
buf ( n4255 , R_780_13cd31f8 );
buf ( n4256 , R_198a_12fc1af8 );
buf ( n4257 , R_72d_13d467d8 );
buf ( n4258 , R_b30_156ac358 );
buf ( n4259 , R_d4c_11633d98 );
buf ( n4260 , R_176e_12fbe678 );
buf ( n4261 , R_136b_15810638 );
buf ( n4262 , R_114f_123ba1b8 );
buf ( n4263 , R_119d_123ba578 );
buf ( n4264 , R_55f_13cce658 );
buf ( n4265 , R_6df_13bf5ef8 );
buf ( n4266 , R_131d_14a11c18 );
buf ( n4267 , R_17bc_15886d98 );
buf ( n4268 , R_b7e_123b7eb8 );
buf ( n4269 , R_cfe_123b7418 );
buf ( n4270 , R_193c_123b6298 );
buf ( n4271 , R_b42_116296b8 );
buf ( n4272 , R_71b_13cd8fb8 );
buf ( n4273 , R_1978_1587e698 );
buf ( n4274 , R_1780_1587b718 );
buf ( n4275 , R_d3a_117f6678 );
buf ( n4276 , R_1161_13beb3b8 );
buf ( n4277 , R_1359_11c6d9d8 );
buf ( n4278 , R_1325_156ac178 );
buf ( n4279 , R_6e7_15882fb8 );
buf ( n4280 , R_557_15885f38 );
buf ( n4281 , R_1195_116363b8 );
buf ( n4282 , R_1944_124c2918 );
buf ( n4283 , R_d06_13dde818 );
buf ( n4284 , R_b76_13d41b98 );
buf ( n4285 , R_17b4_13d29ab8 );
buf ( n4286 , R_1020_117ed258 );
buf ( n4287 , R_85c_1580fc38 );
buf ( n4288 , R_149a_13bf0ef8 );
buf ( n4289 , R_163f_13de4218 );
buf ( n4290 , R_a01_156b1498 );
buf ( n4291 , R_e7b_1486b738 );
buf ( n4292 , R_11c1_123b5618 );
buf ( n4293 , R_cda_156b9878 );
buf ( n4294 , R_1918_15880f38 );
buf ( n4295 , R_583_13cccb78 );
buf ( n4296 , R_17e0_14a15d18 );
buf ( n4297 , R_6bb_117f2398 );
buf ( n4298 , R_ba2_14a0e5b8 );
buf ( n4299 , R_12f9_13d5c9f8 );
buf ( n4300 , R_5ee_12fc0c98 );
buf ( n4301 , R_c0d_13b93fb8 );
buf ( n4302 , R_122c_14b217b8 );
buf ( n4303 , R_18ad_13cd6358 );
buf ( n4304 , R_184b_1486d3f8 );
buf ( n4305 , R_128e_13b91a38 );
buf ( n4306 , R_c6f_150e83d8 );
buf ( n4307 , R_650_116346f8 );
buf ( n4308 , R_5e0_13df04d8 );
buf ( n4309 , R_bff_123b92b8 );
buf ( n4310 , R_18bb_11c6f698 );
buf ( n4311 , R_121e_14b1d438 );
buf ( n4312 , R_129c_1007ebf8 );
buf ( n4313 , R_183d_15882e78 );
buf ( n4314 , R_c7d_13c108f8 );
buf ( n4315 , R_65e_13d43998 );
buf ( n4316 , R_75d_156ad118 );
buf ( n4317 , R_173e_148678b8 );
buf ( n4318 , R_d7c_123be998 );
buf ( n4319 , R_111f_14a110d8 );
buf ( n4320 , R_139b_156b35b8 );
buf ( n4321 , R_b00_13ccf558 );
buf ( n4322 , R_19ba_17014d48 );
buf ( n4323 , R_a78_13cd1cb8 );
buf ( n4324 , R_1a42_15817118 );
buf ( n4325 , R_1097_13d240b8 );
buf ( n4326 , R_1423_13c05a98 );
buf ( n4327 , R_16b6_140aab98 );
buf ( n4328 , R_e04_156b17b8 );
buf ( n4329 , R_7e5_14b1e798 );
buf ( n4330 , R_746_170166e8 );
buf ( n4331 , R_1136_13d56558 );
buf ( n4332 , R_d65_1008bb78 );
buf ( n4333 , R_b17_123bcc38 );
buf ( n4334 , R_1384_140b3298 );
buf ( n4335 , R_19a3_117eaa58 );
buf ( n4336 , R_1755_10087258 );
buf ( n4337 , R_c21_1700d4a8 );
buf ( n4338 , R_1240_11630238 );
buf ( n4339 , R_185f_13bf7118 );
buf ( n4340 , R_1899_156b1fd8 );
buf ( n4341 , R_127a_14b28298 );
buf ( n4342 , R_c5b_13d26278 );
buf ( n4343 , R_63c_1587b538 );
buf ( n4344 , R_602_156afff8 );
buf ( n4345 , R_753_116336b8 );
buf ( n4346 , R_1129_13ccc3f8 );
buf ( n4347 , R_d72_13b95e58 );
buf ( n4348 , R_b0a_156ad438 );
buf ( n4349 , R_1391_15886578 );
buf ( n4350 , R_19b0_17014a28 );
buf ( n4351 , R_1748_117eeab8 );
buf ( n4352 , R_e32_13c05c78 );
buf ( n4353 , R_a4a_117e8bb8 );
buf ( n4354 , R_813_11631318 );
buf ( n4355 , R_1069_116369f8 );
buf ( n4356 , R_1688_156b6a38 );
buf ( n4357 , R_1451_150e6b78 );
buf ( n4358 , R_cdf_150dfa58 );
buf ( n4359 , R_11bc_11c6a9b8 );
buf ( n4360 , R_191d_13c10678 );
buf ( n4361 , R_57e_1162f338 );
buf ( n4362 , R_6c0_13b98c98 );
buf ( n4363 , R_17db_117f6858 );
buf ( n4364 , R_12fe_116291b8 );
buf ( n4365 , R_b9d_14872678 );
buf ( n4366 , R_1349_13d26db8 );
buf ( n4367 , R_b52_1162a978 );
buf ( n4368 , R_1790_117e9798 );
buf ( n4369 , R_70b_17018808 );
buf ( n4370 , R_1968_13bf0318 );
buf ( n4371 , R_d2a_15fef568 );
buf ( n4372 , R_1171_117f5278 );
buf ( n4373 , R_192b_11633cf8 );
buf ( n4374 , R_11ae_123bc238 );
buf ( n4375 , R_570_117ec218 );
buf ( n4376 , R_6ce_13dee1d8 );
buf ( n4377 , R_130c_15ff67c8 );
buf ( n4378 , R_17cd_13b91858 );
buf ( n4379 , R_b8f_14b25b38 );
buf ( n4380 , R_ced_14a0a558 );
buf ( n4381 , R_1582_150e7ed8 );
buf ( n4382 , R_f63_13cca7d8 );
buf ( n4383 , R_944_13d1fab8 );
buf ( n4384 , R_919_123bdf98 );
buf ( n4385 , R_f38_13d26958 );
buf ( n4386 , R_1557_14a16c18 );
buf ( n4387 , R_10ae_123b9358 );
buf ( n4388 , R_16cd_117eee78 );
buf ( n4389 , R_1a2b_140accb8 );
buf ( n4390 , R_140c_11c6f058 );
buf ( n4391 , R_ded_14a14738 );
buf ( n4392 , R_7ce_13d45d38 );
buf ( n4393 , R_a8f_17014de8 );
buf ( n4394 , R_10a5_13d564b8 );
buf ( n4395 , R_16c4_1580f878 );
buf ( n4396 , R_1a34_14a19558 );
buf ( n4397 , R_1415_158165d8 );
buf ( n4398 , R_df6_156b2bb8 );
buf ( n4399 , R_7d7_13c29998 );
buf ( n4400 , R_a86_123bc0f8 );
buf ( n4401 , R_165b_13de0898 );
buf ( n4402 , R_840_156b26b8 );
buf ( n4403 , R_a1d_14a15778 );
buf ( n4404 , R_147e_11638078 );
buf ( n4405 , R_103c_140b0ef8 );
buf ( n4406 , R_e5f_150e3d38 );
buf ( n4407 , R_11c6_13def038 );
buf ( n4408 , R_cd5_13cd09f8 );
buf ( n4409 , R_588_13de09d8 );
buf ( n4410 , R_1913_13beef18 );
buf ( n4411 , R_17e5_150de518 );
buf ( n4412 , R_6b6_13d519b8 );
buf ( n4413 , R_ba7_13d2ca38 );
buf ( n4414 , R_12f4_11c6ca38 );
buf ( n4415 , R_19e8_15888e18 );
buf ( n4416 , R_1710_13bf6718 );
buf ( n4417 , R_10f1_124c52f8 );
buf ( n4418 , R_ad2_156b8658 );
buf ( n4419 , R_78b_1162ddf8 );
buf ( n4420 , R_daa_1008ced8 );
buf ( n4421 , R_13c9_13de18d8 );
buf ( n4422 , R_11a1_117e91f8 );
buf ( n4423 , R_563_13d1ea78 );
buf ( n4424 , R_6db_13dd91d8 );
buf ( n4425 , R_1319_117f10d8 );
buf ( n4426 , R_17c0_15ff4888 );
buf ( n4427 , R_b82_13beff58 );
buf ( n4428 , R_cfa_14b21ad8 );
buf ( n4429 , R_1938_13df6ab8 );
buf ( n4430 , R_82a_14a0cfd8 );
buf ( n4431 , R_a33_11c70278 );
buf ( n4432 , R_1468_158803f8 );
buf ( n4433 , R_1052_117f42d8 );
buf ( n4434 , R_1671_13dd6898 );
buf ( n4435 , R_e49_15ff8f28 );
buf ( n4436 , R_1329_14a16ad8 );
buf ( n4437 , R_6eb_13d45b58 );
buf ( n4438 , R_1191_15881618 );
buf ( n4439 , R_1948_13c26a18 );
buf ( n4440 , R_d0a_158820b8 );
buf ( n4441 , R_b72_13c103f8 );
buf ( n4442 , R_17b0_13decf18 );
buf ( n4443 , R_a36_13b92438 );
buf ( n4444 , R_827_123b8f98 );
buf ( n4445 , R_1055_11635738 );
buf ( n4446 , R_1465_14a18ab8 );
buf ( n4447 , R_1674_11636c78 );
buf ( n4448 , R_e46_15884098 );
buf ( n4449 , R_851_11635238 );
buf ( n4450 , R_148f_13df4358 );
buf ( n4451 , R_164a_13c1e318 );
buf ( n4452 , R_a0c_100899b8 );
buf ( n4453 , R_e70_117ec538 );
buf ( n4454 , R_102b_13d38d18 );
buf ( n4455 , R_198d_156b4378 );
buf ( n4456 , R_730_123bb518 );
buf ( n4457 , R_b2d_124c29b8 );
buf ( n4458 , R_d4f_13cd15d8 );
buf ( n4459 , R_176b_150e5bd8 );
buf ( n4460 , R_136e_15ff6b88 );
buf ( n4461 , R_114c_140b06d8 );
buf ( n4462 , R_16f5_13d39b78 );
buf ( n4463 , R_1a03_14b23338 );
buf ( n4464 , R_10d6_150df4b8 );
buf ( n4465 , R_13e4_13cd99b8 );
buf ( n4466 , R_ab7_1700b748 );
buf ( n4467 , R_dc5_15ff3f28 );
buf ( n4468 , R_7a6_150dad78 );
buf ( n4469 , R_1a05_1162d498 );
buf ( n4470 , R_13e6_1486e578 );
buf ( n4471 , R_dc7_13cd2398 );
buf ( n4472 , R_16f3_10088bf8 );
buf ( n4473 , R_7a8_13beac38 );
buf ( n4474 , R_10d4_13d1de98 );
buf ( n4475 , R_ab5_13df25f8 );
buf ( n4476 , R_82d_13c24b78 );
buf ( n4477 , R_a30_117ef9b8 );
buf ( n4478 , R_146b_150da9b8 );
buf ( n4479 , R_104f_170118c8 );
buf ( n4480 , R_e4c_13ddfd58 );
buf ( n4481 , R_166e_123be3f8 );
buf ( n4482 , R_73e_15883878 );
buf ( n4483 , R_b1f_11631098 );
buf ( n4484 , R_d5d_11636778 );
buf ( n4485 , R_137c_11634e78 );
buf ( n4486 , R_175d_13df13d8 );
buf ( n4487 , R_199b_150dc8f8 );
buf ( n4488 , R_113e_10081ad8 );
buf ( n4489 , R_b45_13cce978 );
buf ( n4490 , R_718_123b4fd8 );
buf ( n4491 , R_1975_13deedb8 );
buf ( n4492 , R_1783_15817e38 );
buf ( n4493 , R_d37_13d26d18 );
buf ( n4494 , R_1164_13df29b8 );
buf ( n4495 , R_1356_15884958 );
buf ( n4496 , R_16f7_140b9558 );
buf ( n4497 , R_10d8_13d55158 );
buf ( n4498 , R_ab9_14a16358 );
buf ( n4499 , R_1a01_14a0bf98 );
buf ( n4500 , R_7a4_13cca698 );
buf ( n4501 , R_13e2_13d50338 );
buf ( n4502 , R_dc3_13d5b918 );
buf ( n4503 , R_1509_13c080b8 );
buf ( n4504 , R_15d0_13d5d7b8 );
buf ( n4505 , R_fb1_17011fa8 );
buf ( n4506 , R_8cb_1162afb8 );
buf ( n4507 , R_992_158117b8 );
buf ( n4508 , R_eea_158843b8 );
buf ( n4509 , R_1a07_15817f78 );
buf ( n4510 , R_13e8_13d57458 );
buf ( n4511 , R_dc9_13dedb98 );
buf ( n4512 , R_7aa_14a113f8 );
buf ( n4513 , R_ab3_13ccea18 );
buf ( n4514 , R_16f1_13c2b298 );
buf ( n4515 , R_10d2_14a0f4b8 );
buf ( n4516 , R_84a_1700eee8 );
buf ( n4517 , R_1651_100849b8 );
buf ( n4518 , R_1488_15811858 );
buf ( n4519 , R_a13_117f7ed8 );
buf ( n4520 , R_e69_14b24ff8 );
buf ( n4521 , R_1032_15884638 );
buf ( n4522 , R_1434_15884a98 );
buf ( n4523 , R_a67_1587c9d8 );
buf ( n4524 , R_e15_117f6538 );
buf ( n4525 , R_1086_158844f8 );
buf ( n4526 , R_16a5_1587d018 );
buf ( n4527 , R_7f6_14a10318 );
buf ( n4528 , R_1a53_11c70b38 );
buf ( n4529 , R_f7b_13c24f38 );
buf ( n4530 , R_95c_13b8ad78 );
buf ( n4531 , R_901_15ff0dc8 );
buf ( n4532 , R_f20_11633078 );
buf ( n4533 , R_153f_140abef8 );
buf ( n4534 , R_159a_13d58d58 );
buf ( n4535 , R_1a20_117f5638 );
buf ( n4536 , R_1401_14a19918 );
buf ( n4537 , R_de2_123bef38 );
buf ( n4538 , R_7c3_14a0f058 );
buf ( n4539 , R_a9a_15816f38 );
buf ( n4540 , R_10b9_15ff6908 );
buf ( n4541 , R_16d8_14b209f8 );
buf ( n4542 , R_1583_13b8ba98 );
buf ( n4543 , R_f64_123b9718 );
buf ( n4544 , R_945_123bcaf8 );
buf ( n4545 , R_918_13c20ed8 );
buf ( n4546 , R_f37_158875b8 );
buf ( n4547 , R_1556_140b5db8 );
buf ( n4548 , R_a39_17016d28 );
buf ( n4549 , R_824_140b4b98 );
buf ( n4550 , R_1058_13b8c7b8 );
buf ( n4551 , R_1462_13d228f8 );
buf ( n4552 , R_1677_1008aef8 );
buf ( n4553 , R_e43_140ab8b8 );
buf ( n4554 , R_123f_12fc2458 );
buf ( n4555 , R_185e_100815d8 );
buf ( n4556 , R_189a_15ff14a8 );
buf ( n4557 , R_127b_13de1a18 );
buf ( n4558 , R_c5c_140b8518 );
buf ( n4559 , R_63d_13df0438 );
buf ( n4560 , R_601_14a12c58 );
buf ( n4561 , R_c20_1486b7d8 );
buf ( n4562 , R_15fd_156b4c38 );
buf ( n4563 , R_ebd_117f1ad8 );
buf ( n4564 , R_fde_13d429f8 );
buf ( n4565 , R_14dc_13ddc5b8 );
buf ( n4566 , R_9bf_15ff2128 );
buf ( n4567 , R_89e_123bbdd8 );
buf ( n4568 , R_16f9_13cd6218 );
buf ( n4569 , R_10da_14a0d4d8 );
buf ( n4570 , R_abb_14b262b8 );
buf ( n4571 , R_7a2_13de1fb8 );
buf ( n4572 , R_dc1_13c211f8 );
buf ( n4573 , R_13e0_1486e4d8 );
buf ( n4574 , R_19ff_123b42b8 );
buf ( n4575 , R_1739_15ff78a8 );
buf ( n4576 , R_d81_140ad4d8 );
buf ( n4577 , R_111a_13d42ef8 );
buf ( n4578 , R_13a0_117f2bb8 );
buf ( n4579 , R_afb_13bf4af8 );
buf ( n4580 , R_19bf_117f5e58 );
buf ( n4581 , R_762_156b33d8 );
buf ( n4582 , R_1a09_1162d358 );
buf ( n4583 , R_13ea_1580dc58 );
buf ( n4584 , R_dcb_1162f798 );
buf ( n4585 , R_7ac_13c08838 );
buf ( n4586 , R_ab1_150e1b78 );
buf ( n4587 , R_10d0_150e7938 );
buf ( n4588 , R_16ef_14a136f8 );
buf ( n4589 , R_a6c_123b7378 );
buf ( n4590 , R_142f_117f79d8 );
buf ( n4591 , R_108b_156b83d8 );
buf ( n4592 , R_e10_14a0b4f8 );
buf ( n4593 , R_16aa_150e47d8 );
buf ( n4594 , R_7f1_123bc378 );
buf ( n4595 , R_1a4e_123b60b8 );
buf ( n4596 , R_5b2_1486f018 );
buf ( n4597 , R_cab_15fee028 );
buf ( n4598 , R_bd1_1587dfb8 );
buf ( n4599 , R_68c_123c1b98 );
buf ( n4600 , R_11f0_13cd3a18 );
buf ( n4601 , R_18e9_13b98a18 );
buf ( n4602 , R_180f_13c1cbf8 );
buf ( n4603 , R_12ca_14a13dd8 );
buf ( n4604 , R_1000_13d4e858 );
buf ( n4605 , R_e9b_13cd5f98 );
buf ( n4606 , R_9e1_13bea878 );
buf ( n4607 , R_161f_10080098 );
buf ( n4608 , R_14ba_1580ba98 );
buf ( n4609 , R_87c_13dee6d8 );
buf ( n4610 , R_830_1008cc58 );
buf ( n4611 , R_a2d_13d43f38 );
buf ( n4612 , R_146e_17010ba8 );
buf ( n4613 , R_104c_13d1f658 );
buf ( n4614 , R_e4f_13ccef18 );
buf ( n4615 , R_166b_116345b8 );
buf ( n4616 , R_ff7_13c0cf78 );
buf ( n4617 , R_ea4_117ea738 );
buf ( n4618 , R_9d8_156b6ad8 );
buf ( n4619 , R_1616_17009da8 );
buf ( n4620 , R_14c3_116384d8 );
buf ( n4621 , R_885_13de02f8 );
buf ( n4622 , R_11b7_11c6de38 );
buf ( n4623 , R_1922_13c26018 );
buf ( n4624 , R_579_13d5d358 );
buf ( n4625 , R_6c5_13d59398 );
buf ( n4626 , R_17d6_11c6d258 );
buf ( n4627 , R_1303_156b3d38 );
buf ( n4628 , R_b98_14b1aeb8 );
buf ( n4629 , R_ce4_117f17b8 );
buf ( n4630 , R_96b_15816c18 );
buf ( n4631 , R_8f2_158891d8 );
buf ( n4632 , R_f11_124c3598 );
buf ( n4633 , R_15a9_1007e0b8 );
buf ( n4634 , R_1530_13c1c5b8 );
buf ( n4635 , R_f8a_1580da78 );
buf ( n4636 , R_5ab_13d20b98 );
buf ( n4637 , R_cb2_15883eb8 );
buf ( n4638 , R_bca_1162ecf8 );
buf ( n4639 , R_693_1580e978 );
buf ( n4640 , R_18f0_14868178 );
buf ( n4641 , R_11e9_12fc0518 );
buf ( n4642 , R_12d1_15ff4388 );
buf ( n4643 , R_1808_117ec998 );
buf ( n4644 , R_112e_124c40d8 );
buf ( n4645 , R_d6d_10080278 );
buf ( n4646 , R_b0f_150e1e98 );
buf ( n4647 , R_138c_14a12938 );
buf ( n4648 , R_19ab_1486d5d8 );
buf ( n4649 , R_174d_13c05318 );
buf ( n4650 , R_74e_117e9dd8 );
buf ( n4651 , R_5d4_1587e918 );
buf ( n4652 , R_18c7_117ed7f8 );
buf ( n4653 , R_bf3_158826f8 );
buf ( n4654 , R_12a8_140b92d8 );
buf ( n4655 , R_1212_13debed8 );
buf ( n4656 , R_c89_15886078 );
buf ( n4657 , R_1831_13b99eb8 );
buf ( n4658 , R_66a_117f7c58 );
buf ( n4659 , R_16fb_13d39a38 );
buf ( n4660 , R_10dc_140acad8 );
buf ( n4661 , R_abd_12fbf938 );
buf ( n4662 , R_7a0_1162cef8 );
buf ( n4663 , R_dbf_13d1dd58 );
buf ( n4664 , R_13de_13bf51d8 );
buf ( n4665 , R_19fd_13c22cd8 );
buf ( n4666 , R_a62_11630378 );
buf ( n4667 , R_e1a_13d29f18 );
buf ( n4668 , R_1081_156ae298 );
buf ( n4669 , R_7fb_13c27c38 );
buf ( n4670 , R_16a0_1007f9b8 );
buf ( n4671 , R_1a58_123b6a18 );
buf ( n4672 , R_1439_11637c18 );
buf ( n4673 , R_1511_1162c778 );
buf ( n4674 , R_15c8_10085a98 );
buf ( n4675 , R_8d3_15fefba8 );
buf ( n4676 , R_fa9_150dc218 );
buf ( n4677 , R_ef2_13d3af78 );
buf ( n4678 , R_98a_11629578 );
buf ( n4679 , R_151a_15ff8d48 );
buf ( n4680 , R_15bf_15ff4f68 );
buf ( n4681 , R_8dc_13dd7b58 );
buf ( n4682 , R_fa0_1162a838 );
buf ( n4683 , R_efb_13ccc2b8 );
buf ( n4684 , R_981_156acad8 );
buf ( n4685 , R_133f_11636ef8 );
buf ( n4686 , R_179a_13ccf918 );
buf ( n4687 , R_701_13dd6438 );
buf ( n4688 , R_195e_15817578 );
buf ( n4689 , R_117b_156b5f98 );
buf ( n4690 , R_d20_1162aa18 );
buf ( n4691 , R_b5c_116370d8 );
buf ( n4692 , R_c0c_13d3f7f8 );
buf ( n4693 , R_122b_117ec498 );
buf ( n4694 , R_18ae_13d39998 );
buf ( n4695 , R_184a_124c54d8 );
buf ( n4696 , R_128f_123b97b8 );
buf ( n4697 , R_c70_15885998 );
buf ( n4698 , R_651_14a122f8 );
buf ( n4699 , R_5ed_13cccad8 );
buf ( n4700 , R_1a0b_1486ee38 );
buf ( n4701 , R_13ec_117f2758 );
buf ( n4702 , R_dcd_13d1e438 );
buf ( n4703 , R_7ae_13d3c058 );
buf ( n4704 , R_aaf_140af698 );
buf ( n4705 , R_10ce_11637538 );
buf ( n4706 , R_16ed_156af558 );
buf ( n4707 , R_a55_12fbef38 );
buf ( n4708 , R_e27_13d405b8 );
buf ( n4709 , R_1074_14b1a878 );
buf ( n4710 , R_808_13c22c38 );
buf ( n4711 , R_1693_13cd4558 );
buf ( n4712 , R_1a65_1587f8b8 );
buf ( n4713 , R_1446_1587eff8 );
buf ( n4714 , R_a3c_150e6038 );
buf ( n4715 , R_821_117f1b78 );
buf ( n4716 , R_105b_13cd2f78 );
buf ( n4717 , R_145f_13b8d398 );
buf ( n4718 , R_167a_13df45d8 );
buf ( n4719 , R_e40_13c26f18 );
buf ( n4720 , R_1584_1580b318 );
buf ( n4721 , R_f65_13d3b5b8 );
buf ( n4722 , R_946_14a10a98 );
buf ( n4723 , R_917_117f5458 );
buf ( n4724 , R_f36_14a118f8 );
buf ( n4725 , R_1555_15815638 );
buf ( n4726 , R_cd0_117f6d58 );
buf ( n4727 , R_58d_1587f3b8 );
buf ( n4728 , R_17ea_15ffadc8 );
buf ( n4729 , R_190e_13bf3d38 );
buf ( n4730 , R_6b1_15ffc808 );
buf ( n4731 , R_bac_13c0a098 );
buf ( n4732 , R_12ef_14b277f8 );
buf ( n4733 , R_11cb_15ff6f48 );
buf ( n4734 , R_977_1580b1d8 );
buf ( n4735 , R_8e6_1580c0d8 );
buf ( n4736 , R_15b5_14866f58 );
buf ( n4737 , R_f05_123b8ef8 );
buf ( n4738 , R_f96_15885538 );
buf ( n4739 , R_1524_1162d178 );
buf ( n4740 , R_11a5_156b5138 );
buf ( n4741 , R_567_13bf17b8 );
buf ( n4742 , R_6d7_12fc12d8 );
buf ( n4743 , R_1315_123b2698 );
buf ( n4744 , R_17c4_13ccc718 );
buf ( n4745 , R_b86_123b9a38 );
buf ( n4746 , R_cf6_14b29738 );
buf ( n4747 , R_1934_123bf7f8 );
buf ( n4748 , R_1338_116375d8 );
buf ( n4749 , R_6fa_13bec218 );
buf ( n4750 , R_1182_13c1c658 );
buf ( n4751 , R_1957_13d3ec18 );
buf ( n4752 , R_d19_13def3f8 );
buf ( n4753 , R_b63_15ffbb88 );
buf ( n4754 , R_17a1_117f24d8 );
buf ( n4755 , R_132d_1587ce38 );
buf ( n4756 , R_6ef_158893b8 );
buf ( n4757 , R_118d_124c3958 );
buf ( n4758 , R_194c_1587cbb8 );
buf ( n4759 , R_d0e_13c10998 );
buf ( n4760 , R_b6e_117ef5f8 );
buf ( n4761 , R_17ac_1486cb38 );
buf ( n4762 , R_12b2_156ab458 );
buf ( n4763 , R_be9_14867638 );
buf ( n4764 , R_c93_14a12258 );
buf ( n4765 , R_1208_13bec358 );
buf ( n4766 , R_674_123c0018 );
buf ( n4767 , R_1827_13c01b78 );
buf ( n4768 , R_18d1_117e98d8 );
buf ( n4769 , R_5ca_13ccca38 );
buf ( n4770 , R_16fd_13bf4378 );
buf ( n4771 , R_10de_140b68f8 );
buf ( n4772 , R_abf_13befd78 );
buf ( n4773 , R_79e_15817b18 );
buf ( n4774 , R_dbd_117f2b18 );
buf ( n4775 , R_13dc_13d1ce58 );
buf ( n4776 , R_19fb_150e3978 );
buf ( n4777 , R_858_150dae18 );
buf ( n4778 , R_1496_13b8b098 );
buf ( n4779 , R_1643_1162c278 );
buf ( n4780 , R_a05_117f4cd8 );
buf ( n4781 , R_e77_1486b878 );
buf ( n4782 , R_1024_11635058 );
buf ( n4783 , R_733_10086998 );
buf ( n4784 , R_b2a_150dd2f8 );
buf ( n4785 , R_d52_1580c498 );
buf ( n4786 , R_1768_15813b58 );
buf ( n4787 , R_1371_156b10d8 );
buf ( n4788 , R_1149_156aff58 );
buf ( n4789 , R_1990_117f1df8 );
buf ( n4790 , R_185d_1162a0b8 );
buf ( n4791 , R_189b_123bccd8 );
buf ( n4792 , R_127c_1580f198 );
buf ( n4793 , R_c5d_13bf88d8 );
buf ( n4794 , R_63e_170163c8 );
buf ( n4795 , R_600_150e8798 );
buf ( n4796 , R_c1f_117ebdb8 );
buf ( n4797 , R_123e_13ccb318 );
buf ( n4798 , R_bfe_17018b28 );
buf ( n4799 , R_18bc_123b9df8 );
buf ( n4800 , R_121d_11632718 );
buf ( n4801 , R_129d_117f6998 );
buf ( n4802 , R_183c_14b21498 );
buf ( n4803 , R_c7e_14a0d6b8 );
buf ( n4804 , R_65f_14874978 );
buf ( n4805 , R_5df_13c24178 );
buf ( n4806 , R_833_117f3dd8 );
buf ( n4807 , R_a2a_14869bb8 );
buf ( n4808 , R_1471_140adbb8 );
buf ( n4809 , R_1049_11636138 );
buf ( n4810 , R_e52_13d4e498 );
buf ( n4811 , R_1668_13b909f8 );
buf ( n4812 , R_15df_14b24c38 );
buf ( n4813 , R_14fa_15ff7128 );
buf ( n4814 , R_fc0_13beba98 );
buf ( n4815 , R_8bc_14a0e338 );
buf ( n4816 , R_9a1_123b5758 );
buf ( n4817 , R_edb_17017048 );
buf ( n4818 , R_1a0d_13ccaaf8 );
buf ( n4819 , R_13ee_13d23398 );
buf ( n4820 , R_dcf_13cccfd8 );
buf ( n4821 , R_7b0_123bf4d8 );
buf ( n4822 , R_aad_14873a78 );
buf ( n4823 , R_10cc_13cd01d8 );
buf ( n4824 , R_16eb_150e81f8 );
buf ( n4825 , R_172d_13cda318 );
buf ( n4826 , R_13ac_116343d8 );
buf ( n4827 , R_110e_14a11998 );
buf ( n4828 , R_19cb_13d3a758 );
buf ( n4829 , R_aef_13d50dd8 );
buf ( n4830 , R_76e_13bf8d38 );
buf ( n4831 , R_d8d_13dd52b8 );
buf ( n4832 , R_715_13b94ff8 );
buf ( n4833 , R_1972_156aa918 );
buf ( n4834 , R_1786_140b5778 );
buf ( n4835 , R_d34_15ff3b68 );
buf ( n4836 , R_1167_1587c7f8 );
buf ( n4837 , R_1353_123c05b8 );
buf ( n4838 , R_b48_15814378 );
buf ( n4839 , R_17fb_11c6bd18 );
buf ( n4840 , R_59e_13cd0098 );
buf ( n4841 , R_cbf_15fed948 );
buf ( n4842 , R_bbd_13b8f418 );
buf ( n4843 , R_18fd_15882798 );
buf ( n4844 , R_6a0_117edbb8 );
buf ( n4845 , R_11dc_150db458 );
buf ( n4846 , R_12de_117e9658 );
buf ( n4847 , R_19db_123b8458 );
buf ( n4848 , R_171d_13d45e78 );
buf ( n4849 , R_10fe_117ebd18 );
buf ( n4850 , R_adf_13ccfcd8 );
buf ( n4851 , R_77e_123bcff8 );
buf ( n4852 , R_d9d_12fc0298 );
buf ( n4853 , R_13bc_13c07cf8 );
buf ( n4854 , R_142a_14a0f2d8 );
buf ( n4855 , R_1090_1486e7f8 );
buf ( n4856 , R_e0b_156b7758 );
buf ( n4857 , R_16af_1486be18 );
buf ( n4858 , R_7ec_123b4038 );
buf ( n4859 , R_1a49_13ccbb38 );
buf ( n4860 , R_a71_117f59f8 );
buf ( n4861 , R_15f2_13d4fe38 );
buf ( n4862 , R_ec8_15883058 );
buf ( n4863 , R_fd3_10088798 );
buf ( n4864 , R_14e7_14b1ce98 );
buf ( n4865 , R_9b4_13bf5b38 );
buf ( n4866 , R_8a9_13c21298 );
buf ( n4867 , R_ece_11634bf8 );
buf ( n4868 , R_15ec_13d3f4d8 );
buf ( n4869 , R_14ed_117f5f98 );
buf ( n4870 , R_fcd_1580d258 );
buf ( n4871 , R_8af_13ddfb78 );
buf ( n4872 , R_9ae_140b18f8 );
buf ( n4873 , R_1501_117f0a98 );
buf ( n4874 , R_15d8_11c6ea18 );
buf ( n4875 , R_fb9_15ff0be8 );
buf ( n4876 , R_8c3_10081498 );
buf ( n4877 , R_99a_15ffaaa8 );
buf ( n4878 , R_ee2_13cd1b78 );
buf ( n4879 , R_1712_11637178 );
buf ( n4880 , R_10f3_14a19238 );
buf ( n4881 , R_ad4_14a0a5f8 );
buf ( n4882 , R_789_140b2cf8 );
buf ( n4883 , R_da8_140b3838 );
buf ( n4884 , R_13c7_13df0ed8 );
buf ( n4885 , R_19e6_11636958 );
buf ( n4886 , R_95d_117f8338 );
buf ( n4887 , R_900_140b74d8 );
buf ( n4888 , R_f1f_1587f1d8 );
buf ( n4889 , R_153e_13d410f8 );
buf ( n4890 , R_159b_1162f658 );
buf ( n4891 , R_f7c_15ffc268 );
buf ( n4892 , R_cc5_13b8c858 );
buf ( n4893 , R_598_17015108 );
buf ( n4894 , R_17f5_13c1c798 );
buf ( n4895 , R_1903_1162d2b8 );
buf ( n4896 , R_6a6_15816df8 );
buf ( n4897 , R_bb7_14a17a78 );
buf ( n4898 , R_12e4_13df4678 );
buf ( n4899 , R_11d6_13cccf38 );
buf ( n4900 , R_a4d_14a159f8 );
buf ( n4901 , R_810_1007f918 );
buf ( n4902 , R_106c_13cd4238 );
buf ( n4903 , R_168b_13d20d78 );
buf ( n4904 , R_144e_17019028 );
buf ( n4905 , R_e2f_123b83b8 );
buf ( n4906 , R_f66_1700e448 );
buf ( n4907 , R_947_13cd36f8 );
buf ( n4908 , R_916_12fbefd8 );
buf ( n4909 , R_f35_13dd5fd8 );
buf ( n4910 , R_1554_13c04918 );
buf ( n4911 , R_1585_117efe18 );
buf ( n4912 , R_16ff_13b95318 );
buf ( n4913 , R_10e0_1580e478 );
buf ( n4914 , R_ac1_13d23078 );
buf ( n4915 , R_79c_1162d8f8 );
buf ( n4916 , R_dbb_1580e018 );
buf ( n4917 , R_13da_123c03d8 );
buf ( n4918 , R_19f9_13cd81f8 );
buf ( n4919 , R_a3f_13c012b8 );
buf ( n4920 , R_81e_140b4cd8 );
buf ( n4921 , R_105e_156ba278 );
buf ( n4922 , R_145c_13ddc0b8 );
buf ( n4923 , R_167d_124c5438 );
buf ( n4924 , R_e3d_15889778 );
buf ( n4925 , R_be0_117ea5f8 );
buf ( n4926 , R_c9c_13b8ed38 );
buf ( n4927 , R_11ff_14a17618 );
buf ( n4928 , R_67d_156b7398 );
buf ( n4929 , R_181e_13c04e18 );
buf ( n4930 , R_18da_13cd38d8 );
buf ( n4931 , R_5c1_13c0a818 );
buf ( n4932 , R_12bb_13b8a918 );
buf ( n4933 , R_ca4_156b1c18 );
buf ( n4934 , R_bd8_117e87f8 );
buf ( n4935 , R_685_13bf38d8 );
buf ( n4936 , R_11f7_10080b38 );
buf ( n4937 , R_18e2_13becfd8 );
buf ( n4938 , R_1816_14b1ff58 );
buf ( n4939 , R_12c3_10083478 );
buf ( n4940 , R_5b9_140b2bb8 );
buf ( n4941 , R_1630_123b9cb8 );
buf ( n4942 , R_e8a_14b1db18 );
buf ( n4943 , R_9f2_10089418 );
buf ( n4944 , R_14a9_156acb78 );
buf ( n4945 , R_1011_12fbe218 );
buf ( n4946 , R_86b_124c4e98 );
buf ( n4947 , R_1726_14869a78 );
buf ( n4948 , R_19d2_13d533f8 );
buf ( n4949 , R_1107_13df9038 );
buf ( n4950 , R_ae8_13bef5f8 );
buf ( n4951 , R_775_158109f8 );
buf ( n4952 , R_d94_12fbf6b8 );
buf ( n4953 , R_13b3_13d40158 );
buf ( n4954 , R_1658_13bf9ff8 );
buf ( n4955 , R_843_150e0458 );
buf ( n4956 , R_1481_117e8e38 );
buf ( n4957 , R_a1a_15fefd88 );
buf ( n4958 , R_1039_13ddba78 );
buf ( n4959 , R_e62_13c23098 );
buf ( n4960 , R_1a0f_13c24038 );
buf ( n4961 , R_13f0_11c6e338 );
buf ( n4962 , R_dd1_13de4a38 );
buf ( n4963 , R_7b2_13bf2898 );
buf ( n4964 , R_aab_13c1cfb8 );
buf ( n4965 , R_10ca_1700ac08 );
buf ( n4966 , R_16e9_15ff3668 );
buf ( n4967 , R_1793_150de018 );
buf ( n4968 , R_708_14a0d258 );
buf ( n4969 , R_1965_13ccb6d8 );
buf ( n4970 , R_1174_11c6c358 );
buf ( n4971 , R_d27_13dee138 );
buf ( n4972 , R_b55_15ffb0e8 );
buf ( n4973 , R_1346_13d3f2f8 );
buf ( n4974 , R_e1f_123b6ab8 );
buf ( n4975 , R_107c_117f4058 );
buf ( n4976 , R_800_13d219f8 );
buf ( n4977 , R_169b_150e49b8 );
buf ( n4978 , R_1a5d_1486e398 );
buf ( n4979 , R_143e_14a19f58 );
buf ( n4980 , R_a5d_15880498 );
buf ( n4981 , R_1a22_15810b38 );
buf ( n4982 , R_1403_124c5398 );
buf ( n4983 , R_de4_117f6498 );
buf ( n4984 , R_7c5_15ffbe08 );
buf ( n4985 , R_a98_1486db78 );
buf ( n4986 , R_10b7_14a17578 );
buf ( n4987 , R_16d6_14a10458 );
buf ( n4988 , R_1a2d_13b8fcd8 );
buf ( n4989 , R_140e_13def718 );
buf ( n4990 , R_def_13d3eb78 );
buf ( n4991 , R_7d0_156b2e38 );
buf ( n4992 , R_a8d_11632678 );
buf ( n4993 , R_10ac_156b5958 );
buf ( n4994 , R_16cb_156b72f8 );
buf ( n4995 , R_1634_17018c68 );
buf ( n4996 , R_9f6_158867f8 );
buf ( n4997 , R_e86_14a183d8 );
buf ( n4998 , R_1015_14b1e6f8 );
buf ( n4999 , R_867_15881398 );
buf ( n5000 , R_14a5_11629ed8 );
buf ( n5001 , R_e8e_150da878 );
buf ( n5002 , R_9ee_13d54618 );
buf ( n5003 , R_162c_13b96c18 );
buf ( n5004 , R_14ad_12fbf618 );
buf ( n5005 , R_86f_15ff83e8 );
buf ( n5006 , R_100d_158136f8 );
buf ( n5007 , R_189c_14a10c78 );
buf ( n5008 , R_127d_11636318 );
buf ( n5009 , R_c5e_15882a18 );
buf ( n5010 , R_63f_156b5b38 );
buf ( n5011 , R_5ff_13d40ab8 );
buf ( n5012 , R_c1e_14a0b958 );
buf ( n5013 , R_123d_13ddd5f8 );
buf ( n5014 , R_185c_11630738 );
buf ( n5015 , R_141e_13b90818 );
buf ( n5016 , R_16bb_123b7d78 );
buf ( n5017 , R_dff_117eeb58 );
buf ( n5018 , R_7e0_13dfacf8 );
buf ( n5019 , R_a7d_123b7af8 );
buf ( n5020 , R_1a3d_156b9cd8 );
buf ( n5021 , R_109c_13b98d38 );
buf ( n5022 , R_cb9_150db638 );
buf ( n5023 , R_bc3_156b6678 );
buf ( n5024 , R_69a_13b8b6d8 );
buf ( n5025 , R_18f7_13b90bd8 );
buf ( n5026 , R_11e2_13d1e4d8 );
buf ( n5027 , R_12d8_13d43718 );
buf ( n5028 , R_1801_13c013f8 );
buf ( n5029 , R_5a4_15ff7d08 );
buf ( n5030 , R_13a5_13d45338 );
buf ( n5031 , R_1115_11630b98 );
buf ( n5032 , R_19c4_17016fa8 );
buf ( n5033 , R_af6_117f49b8 );
buf ( n5034 , R_767_117f2d98 );
buf ( n5035 , R_d86_15fef7e8 );
buf ( n5036 , R_1734_1580c718 );
buf ( n5037 , R_836_123b33b8 );
buf ( n5038 , R_a27_117ede38 );
buf ( n5039 , R_1474_13c042d8 );
buf ( n5040 , R_1046_123bc918 );
buf ( n5041 , R_e55_124c3a98 );
buf ( n5042 , R_1665_156ac678 );
buf ( n5043 , R_122a_14a0b318 );
buf ( n5044 , R_18af_11c6f7d8 );
buf ( n5045 , R_1849_140b6358 );
buf ( n5046 , R_1290_13dd8b98 );
buf ( n5047 , R_c71_14a11e98 );
buf ( n5048 , R_652_13d386d8 );
buf ( n5049 , R_5ec_14868df8 );
buf ( n5050 , R_c0b_13b8c038 );
buf ( n5051 , R_574_13d4ec18 );
buf ( n5052 , R_6ca_156b3f18 );
buf ( n5053 , R_1308_117f2438 );
buf ( n5054 , R_17d1_11c6fa58 );
buf ( n5055 , R_b93_15881078 );
buf ( n5056 , R_ce9_156b86f8 );
buf ( n5057 , R_1927_123bb6f8 );
buf ( n5058 , R_11b2_14a101d8 );
buf ( n5059 , R_8f1_14a0fcd8 );
buf ( n5060 , R_f10_156ab778 );
buf ( n5061 , R_15aa_13c1f498 );
buf ( n5062 , R_152f_158884b8 );
buf ( n5063 , R_f8b_13dda218 );
buf ( n5064 , R_96c_15ff4e28 );
buf ( n5065 , R_948_15ff1728 );
buf ( n5066 , R_915_158834b8 );
buf ( n5067 , R_f34_123bd958 );
buf ( n5068 , R_1553_1162fdd8 );
buf ( n5069 , R_1586_13cd7938 );
buf ( n5070 , R_f67_156b54f8 );
buf ( n5071 , R_1701_117ee5b8 );
buf ( n5072 , R_10e2_13b97cf8 );
buf ( n5073 , R_ac3_13d41ff8 );
buf ( n5074 , R_79a_13b8d758 );
buf ( n5075 , R_db9_13d4e358 );
buf ( n5076 , R_13d8_13c10178 );
buf ( n5077 , R_19f7_123b4218 );
buf ( n5078 , R_ec2_156acdf8 );
buf ( n5079 , R_fd9_13cd6038 );
buf ( n5080 , R_14e1_13d4fbb8 );
buf ( n5081 , R_9ba_13d3b018 );
buf ( n5082 , R_8a3_117f3298 );
buf ( n5083 , R_15f8_150dd618 );
buf ( n5084 , R_b1c_10084238 );
buf ( n5085 , R_d60_1700c1e8 );
buf ( n5086 , R_137f_13d27fd8 );
buf ( n5087 , R_175a_15fedda8 );
buf ( n5088 , R_199e_123b8d18 );
buf ( n5089 , R_113b_11c703b8 );
buf ( n5090 , R_741_156b0278 );
buf ( n5091 , R_15e6_140b4238 );
buf ( n5092 , R_14f3_10088a18 );
buf ( n5093 , R_fc7_117e8c58 );
buf ( n5094 , R_8b5_13ccefb8 );
buf ( n5095 , R_9a8_14a19af8 );
buf ( n5096 , R_ed4_150e1998 );
buf ( n5097 , R_d68_15885b78 );
buf ( n5098 , R_b14_11c6b8b8 );
buf ( n5099 , R_1387_117eaf58 );
buf ( n5100 , R_19a6_14a19738 );
buf ( n5101 , R_1752_150e4738 );
buf ( n5102 , R_749_123b2918 );
buf ( n5103 , R_1133_1587e378 );
buf ( n5104 , R_1417_15ff4428 );
buf ( n5105 , R_df8_15888eb8 );
buf ( n5106 , R_7d9_124c3098 );
buf ( n5107 , R_a84_13b8b778 );
buf ( n5108 , R_10a3_13c1e4f8 );
buf ( n5109 , R_1a36_14b1b318 );
buf ( n5110 , R_16c2_156b1e98 );
buf ( n5111 , R_1a11_123b7b98 );
buf ( n5112 , R_13f2_13de2738 );
buf ( n5113 , R_dd3_14a19a58 );
buf ( n5114 , R_7b4_15885a38 );
buf ( n5115 , R_aa9_13cd5818 );
buf ( n5116 , R_10c8_14a14058 );
buf ( n5117 , R_16e7_117eea18 );
buf ( n5118 , R_b27_10087e38 );
buf ( n5119 , R_d55_117f0f98 );
buf ( n5120 , R_1765_12fbdf98 );
buf ( n5121 , R_1374_17015888 );
buf ( n5122 , R_1146_123bed58 );
buf ( n5123 , R_1993_13d53b78 );
buf ( n5124 , R_736_15ff9108 );
buf ( n5125 , R_56b_123b7558 );
buf ( n5126 , R_6d3_1007e1f8 );
buf ( n5127 , R_1311_10087a78 );
buf ( n5128 , R_17c8_13d50a18 );
buf ( n5129 , R_b8a_14b26858 );
buf ( n5130 , R_cf2_14a17438 );
buf ( n5131 , R_1930_13c083d8 );
buf ( n5132 , R_11a9_117f1038 );
buf ( n5133 , R_1638_15815818 );
buf ( n5134 , R_9fa_123b77d8 );
buf ( n5135 , R_e82_13df3ef8 );
buf ( n5136 , R_1019_158858f8 );
buf ( n5137 , R_863_13d47318 );
buf ( n5138 , R_14a1_117ed938 );
buf ( n5139 , R_eb2_11c6d2f8 );
buf ( n5140 , R_fe9_1162ed98 );
buf ( n5141 , R_14d1_1587ae58 );
buf ( n5142 , R_9ca_1587bd58 );
buf ( n5143 , R_893_13ccf238 );
buf ( n5144 , R_1608_117f45f8 );
buf ( n5145 , R_6f3_17012cc8 );
buf ( n5146 , R_1189_13de2d78 );
buf ( n5147 , R_1950_123b8098 );
buf ( n5148 , R_d12_13cd6d58 );
buf ( n5149 , R_b6a_140afff8 );
buf ( n5150 , R_17a8_13d3cf58 );
buf ( n5151 , R_1331_148755f8 );
buf ( n5152 , R_e9f_17016288 );
buf ( n5153 , R_9dd_156ab8b8 );
buf ( n5154 , R_161b_13d3ca58 );
buf ( n5155 , R_14be_13b98478 );
buf ( n5156 , R_880_117ea2d8 );
buf ( n5157 , R_ffc_13b8acd8 );
buf ( n5158 , R_1789_13cca9b8 );
buf ( n5159 , R_196f_13bf01d8 );
buf ( n5160 , R_d31_156b13f8 );
buf ( n5161 , R_116a_13c23e58 );
buf ( n5162 , R_1350_11632498 );
buf ( n5163 , R_b4b_156ad398 );
buf ( n5164 , R_712_13b90d18 );
buf ( n5165 , R_e92_117f2ed8 );
buf ( n5166 , R_9ea_123b7e18 );
buf ( n5167 , R_1628_123b7698 );
buf ( n5168 , R_14b1_14a16e98 );
buf ( n5169 , R_873_14a14238 );
buf ( n5170 , R_1009_13b980b8 );
buf ( n5171 , R_bf2_170099e8 );
buf ( n5172 , R_12a9_1162d0d8 );
buf ( n5173 , R_1211_150e5278 );
buf ( n5174 , R_c8a_150e3798 );
buf ( n5175 , R_1830_13bf6358 );
buf ( n5176 , R_66b_150e1498 );
buf ( n5177 , R_5d3_158808f8 );
buf ( n5178 , R_18c8_13cd9f58 );
buf ( n5179 , R_a42_15888198 );
buf ( n5180 , R_81b_12fbec18 );
buf ( n5181 , R_1061_13d3c558 );
buf ( n5182 , R_1459_17016aa8 );
buf ( n5183 , R_1680_1486aab8 );
buf ( n5184 , R_e3a_123bb798 );
buf ( n5185 , R_17ef_15889958 );
buf ( n5186 , R_1909_15815e58 );
buf ( n5187 , R_6ac_12fc1918 );
buf ( n5188 , R_bb1_14874d38 );
buf ( n5189 , R_12ea_13ddf358 );
buf ( n5190 , R_11d0_170096c8 );
buf ( n5191 , R_ccb_117ec038 );
buf ( n5192 , R_592_13c23958 );
buf ( n5193 , R_fee_14b29f58 );
buf ( n5194 , R_ead_13c22378 );
buf ( n5195 , R_9cf_1162e118 );
buf ( n5196 , R_14cc_123c0b58 );
buf ( n5197 , R_160d_123bff78 );
buf ( n5198 , R_88e_123c0fb8 );
buf ( n5199 , R_8ff_156b7c58 );
buf ( n5200 , R_f1e_15880038 );
buf ( n5201 , R_153d_15811218 );
buf ( n5202 , R_159c_15815db8 );
buf ( n5203 , R_f7d_13cd0778 );
buf ( n5204 , R_95e_13b98018 );
buf ( n5205 , R_189d_13cd3518 );
buf ( n5206 , R_127e_13d4f118 );
buf ( n5207 , R_c5f_12fbfa78 );
buf ( n5208 , R_640_140b2258 );
buf ( n5209 , R_5fe_15888558 );
buf ( n5210 , R_c1d_13dfb1f8 );
buf ( n5211 , R_123c_15fee708 );
buf ( n5212 , R_185b_14b21538 );
buf ( n5213 , R_15d1_123b63d8 );
buf ( n5214 , R_fb2_15810818 );
buf ( n5215 , R_8ca_15815bd8 );
buf ( n5216 , R_993_11c6b598 );
buf ( n5217 , R_ee9_1700fca8 );
buf ( n5218 , R_1508_156b7898 );
buf ( n5219 , R_121c_158871f8 );
buf ( n5220 , R_129e_13d3cb98 );
buf ( n5221 , R_183b_13c20bb8 );
buf ( n5222 , R_c7f_13cd6ad8 );
buf ( n5223 , R_660_156ba458 );
buf ( n5224 , R_5de_123b7cd8 );
buf ( n5225 , R_18bd_140b9878 );
buf ( n5226 , R_bfd_11c6f238 );
buf ( n5227 , R_16b4_117ead78 );
buf ( n5228 , R_e06_1580ff58 );
buf ( n5229 , R_7e7_15885858 );
buf ( n5230 , R_1a44_1162c4f8 );
buf ( n5231 , R_a76_13d38638 );
buf ( n5232 , R_1095_156b0ef8 );
buf ( n5233 , R_1425_13d571d8 );
buf ( n5234 , R_8e5_150db318 );
buf ( n5235 , R_15b6_1580e838 );
buf ( n5236 , R_f04_15885038 );
buf ( n5237 , R_f97_1700c288 );
buf ( n5238 , R_1523_140b8e78 );
buf ( n5239 , R_978_156b6498 );
buf ( n5240 , R_914_13d54c58 );
buf ( n5241 , R_f33_13d59258 );
buf ( n5242 , R_1552_13ccfa58 );
buf ( n5243 , R_1587_140aacd8 );
buf ( n5244 , R_f68_140acb78 );
buf ( n5245 , R_949_14b26a38 );
buf ( n5246 , R_15c0_158147d8 );
buf ( n5247 , R_8db_1580e158 );
buf ( n5248 , R_fa1_1162ffb8 );
buf ( n5249 , R_efa_13bf5818 );
buf ( n5250 , R_982_13debcf8 );
buf ( n5251 , R_1519_15813e78 );
buf ( n5252 , R_164e_117eb138 );
buf ( n5253 , R_148b_15886118 );
buf ( n5254 , R_a10_13df0f78 );
buf ( n5255 , R_e6c_15ff0d28 );
buf ( n5256 , R_102f_123c08d8 );
buf ( n5257 , R_84d_15feee88 );
buf ( n5258 , R_1703_13c254d8 );
buf ( n5259 , R_10e4_158894f8 );
buf ( n5260 , R_ac5_15883558 );
buf ( n5261 , R_798_123beb78 );
buf ( n5262 , R_db7_14869938 );
buf ( n5263 , R_13d6_156ae8d8 );
buf ( n5264 , R_19f5_13d2c2b8 );
buf ( n5265 , R_eb7_11c6d1b8 );
buf ( n5266 , R_fe4_12fc21d8 );
buf ( n5267 , R_14d6_1008b178 );
buf ( n5268 , R_9c5_14b21d58 );
buf ( n5269 , R_898_123b5c58 );
buf ( n5270 , R_1603_14872fd8 );
buf ( n5271 , R_1714_15889638 );
buf ( n5272 , R_10f5_140b5f98 );
buf ( n5273 , R_ad6_14873258 );
buf ( n5274 , R_787_14a0e838 );
buf ( n5275 , R_da6_13ddc158 );
buf ( n5276 , R_13c5_15fee208 );
buf ( n5277 , R_19e4_13de3a98 );
buf ( n5278 , R_98b_13b8dcf8 );
buf ( n5279 , R_ef1_13b924d8 );
buf ( n5280 , R_8d2_156ad578 );
buf ( n5281 , R_faa_156b0458 );
buf ( n5282 , R_1510_13d1f0b8 );
buf ( n5283 , R_15c9_13bf0b38 );
buf ( n5284 , R_aa7_13d451f8 );
buf ( n5285 , R_7b6_14a18018 );
buf ( n5286 , R_dd5_124c5258 );
buf ( n5287 , R_10c6_1700ff28 );
buf ( n5288 , R_13f4_14a0b778 );
buf ( n5289 , R_16e5_13c07ed8 );
buf ( n5290 , R_1a13_117ef058 );
buf ( n5291 , R_839_14b28f18 );
buf ( n5292 , R_e58_158814d8 );
buf ( n5293 , R_a24_123b5938 );
buf ( n5294 , R_1043_14b26538 );
buf ( n5295 , R_1477_117f0098 );
buf ( n5296 , R_1662_13df1978 );
buf ( n5297 , R_854_15ff3e88 );
buf ( n5298 , R_e73_14b288d8 );
buf ( n5299 , R_a09_123bb158 );
buf ( n5300 , R_1028_117f4eb8 );
buf ( n5301 , R_1492_13cd4378 );
buf ( n5302 , R_1647_12fc19b8 );
buf ( n5303 , R_be8_15ffcee8 );
buf ( n5304 , R_5c9_14b27438 );
buf ( n5305 , R_675_156aec98 );
buf ( n5306 , R_c94_13b8fb98 );
buf ( n5307 , R_1207_156b81f8 );
buf ( n5308 , R_12b3_13ddf718 );
buf ( n5309 , R_1826_140b01d8 );
buf ( n5310 , R_18d2_13c290d8 );
buf ( n5311 , R_cac_123c1058 );
buf ( n5312 , R_5b1_13d28e38 );
buf ( n5313 , R_68d_1700f2a8 );
buf ( n5314 , R_bd0_13ccc538 );
buf ( n5315 , R_11ef_117f3d38 );
buf ( n5316 , R_12cb_123bfe38 );
buf ( n5317 , R_180e_1580c7b8 );
buf ( n5318 , R_18ea_14a115d8 );
buf ( n5319 , R_d75_1486bc38 );
buf ( n5320 , R_756_13b8ae18 );
buf ( n5321 , R_b07_140aaa58 );
buf ( n5322 , R_1126_156aaeb8 );
buf ( n5323 , R_1394_15814878 );
buf ( n5324 , R_1745_123b4cb8 );
buf ( n5325 , R_19b3_123bc558 );
buf ( n5326 , R_d7a_13b95ef8 );
buf ( n5327 , R_75b_15814558 );
buf ( n5328 , R_b02_14a13f18 );
buf ( n5329 , R_1121_150e9c38 );
buf ( n5330 , R_1399_158830f8 );
buf ( n5331 , R_1740_13cd6fd8 );
buf ( n5332 , R_19b8_15812c58 );
buf ( n5333 , R_c0a_14a19ff8 );
buf ( n5334 , R_5eb_15feeac8 );
buf ( n5335 , R_653_123be358 );
buf ( n5336 , R_c72_13df6fb8 );
buf ( n5337 , R_1229_156b7938 );
buf ( n5338 , R_1291_14a0d758 );
buf ( n5339 , R_1848_14a197d8 );
buf ( n5340 , R_18b0_15815a98 );
buf ( n5341 , R_a96_150e8478 );
buf ( n5342 , R_7c7_13d45c98 );
buf ( n5343 , R_de6_13c05778 );
buf ( n5344 , R_10b5_156ab6d8 );
buf ( n5345 , R_1405_14a192d8 );
buf ( n5346 , R_16d4_14868c18 );
buf ( n5347 , R_1a24_116348d8 );
buf ( n5348 , R_85f_13dd89b8 );
buf ( n5349 , R_e7e_140ad6b8 );
buf ( n5350 , R_9fe_13c02d98 );
buf ( n5351 , R_101d_123b5d98 );
buf ( n5352 , R_149d_156b8dd8 );
buf ( n5353 , R_163c_1486a6f8 );
buf ( n5354 , R_d9b_13d3dbd8 );
buf ( n5355 , R_77c_116359b8 );
buf ( n5356 , R_ae1_15fed768 );
buf ( n5357 , R_1100_10085818 );
buf ( n5358 , R_13ba_15881d98 );
buf ( n5359 , R_171f_13bf08b8 );
buf ( n5360 , R_19d9_1700c508 );
buf ( n5361 , R_889_15ff9b08 );
buf ( n5362 , R_9d4_11c6e6f8 );
buf ( n5363 , R_ea8_13d1fe78 );
buf ( n5364 , R_ff3_117efc38 );
buf ( n5365 , R_14c7_140b4918 );
buf ( n5366 , R_1612_13cd0278 );
buf ( n5367 , R_582_14869118 );
buf ( n5368 , R_cdb_14a0ae18 );
buf ( n5369 , R_ba1_13d29338 );
buf ( n5370 , R_6bc_13cd53b8 );
buf ( n5371 , R_11c0_13deef98 );
buf ( n5372 , R_12fa_11631638 );
buf ( n5373 , R_17df_13cd0e58 );
buf ( n5374 , R_1919_1587e2d8 );
buf ( n5375 , R_e24_13ddcfb8 );
buf ( n5376 , R_a58_14a18a18 );
buf ( n5377 , R_805_1580a7d8 );
buf ( n5378 , R_1077_11c6d898 );
buf ( n5379 , R_1443_13d3f9d8 );
buf ( n5380 , R_1696_156afd78 );
buf ( n5381 , R_1a62_14b1b138 );
buf ( n5382 , R_94a_156b24d8 );
buf ( n5383 , R_f32_116350f8 );
buf ( n5384 , R_913_100840f8 );
buf ( n5385 , R_f69_117f0c78 );
buf ( n5386 , R_1551_150dde38 );
buf ( n5387 , R_1588_150e7d98 );
buf ( n5388 , R_a50_13df7698 );
buf ( n5389 , R_e2c_15881e38 );
buf ( n5390 , R_80d_14a16a38 );
buf ( n5391 , R_106f_156ad938 );
buf ( n5392 , R_144b_1486ce58 );
buf ( n5393 , R_168e_123bbc98 );
buf ( n5394 , R_6fe_13bf5318 );
buf ( n5395 , R_b5f_13cd4918 );
buf ( n5396 , R_d1d_13def2b8 );
buf ( n5397 , R_117e_14a0ccb8 );
buf ( n5398 , R_133c_117f2938 );
buf ( n5399 , R_179d_10085138 );
buf ( n5400 , R_195b_14b1c8f8 );
buf ( n5401 , R_cb3_1587b358 );
buf ( n5402 , R_5aa_13dd5678 );
buf ( n5403 , R_694_11636b38 );
buf ( n5404 , R_bc9_124c3d18 );
buf ( n5405 , R_11e8_13ccd258 );
buf ( n5406 , R_12d2_123bdc78 );
buf ( n5407 , R_1807_117ee298 );
buf ( n5408 , R_18f1_156aba98 );
buf ( n5409 , R_c1c_156ba3b8 );
buf ( n5410 , R_5fd_14a10958 );
buf ( n5411 , R_641_123b90d8 );
buf ( n5412 , R_c60_158171b8 );
buf ( n5413 , R_123b_1162cd18 );
buf ( n5414 , R_127f_13b8a558 );
buf ( n5415 , R_185a_15814cd8 );
buf ( n5416 , R_189e_13bf8e78 );
buf ( n5417 , R_877_13d3e498 );
buf ( n5418 , R_9e6_14b28838 );
buf ( n5419 , R_e96_156b4a58 );
buf ( n5420 , R_1005_13c1edb8 );
buf ( n5421 , R_14b5_15882018 );
buf ( n5422 , R_1624_10086cb8 );
buf ( n5423 , R_db5_117ece98 );
buf ( n5424 , R_796_156b0138 );
buf ( n5425 , R_ac7_148725d8 );
buf ( n5426 , R_10e6_11630918 );
buf ( n5427 , R_13d4_15882bf8 );
buf ( n5428 , R_1705_10085db8 );
buf ( n5429 , R_19f3_1008c618 );
buf ( n5430 , R_96d_1162e7f8 );
buf ( n5431 , R_f0f_13d3d9f8 );
buf ( n5432 , R_8f0_13d29838 );
buf ( n5433 , R_f8c_117f2578 );
buf ( n5434 , R_152e_117f3f18 );
buf ( n5435 , R_15ab_13ccc358 );
buf ( n5436 , R_587_124c5118 );
buf ( n5437 , R_cd6_13d39178 );
buf ( n5438 , R_ba6_156ad9d8 );
buf ( n5439 , R_6b7_13c0b718 );
buf ( n5440 , R_11c5_13d39538 );
buf ( n5441 , R_12f5_158104f8 );
buf ( n5442 , R_17e4_156acf38 );
buf ( n5443 , R_1914_10084f58 );
buf ( n5444 , R_846_100885b8 );
buf ( n5445 , R_e65_15810318 );
buf ( n5446 , R_a17_13ccf878 );
buf ( n5447 , R_1036_140b5278 );
buf ( n5448 , R_1484_11c6b778 );
buf ( n5449 , R_1655_1700cdc8 );
buf ( n5450 , R_a45_17017188 );
buf ( n5451 , R_e37_10083018 );
buf ( n5452 , R_818_13b8dbb8 );
buf ( n5453 , R_1064_1700d5e8 );
buf ( n5454 , R_1456_13cd8518 );
buf ( n5455 , R_1683_1587f6d8 );
buf ( n5456 , R_57d_14b1ef18 );
buf ( n5457 , R_ce0_1580ccb8 );
buf ( n5458 , R_b9c_15884e58 );
buf ( n5459 , R_6c1_156b1538 );
buf ( n5460 , R_11bb_117ed2f8 );
buf ( n5461 , R_12ff_17012408 );
buf ( n5462 , R_17da_123bf398 );
buf ( n5463 , R_191e_140b0c78 );
buf ( n5464 , R_d58_13df39f8 );
buf ( n5465 , R_b24_15815958 );
buf ( n5466 , R_739_123c1698 );
buf ( n5467 , R_1143_13cd7078 );
buf ( n5468 , R_1377_158873d8 );
buf ( n5469 , R_1762_140aef18 );
buf ( n5470 , R_1996_156b4058 );
buf ( n5471 , R_95f_13bf9918 );
buf ( n5472 , R_f1d_15ff80c8 );
buf ( n5473 , R_8fe_13d4f898 );
buf ( n5474 , R_f7e_156b42d8 );
buf ( n5475 , R_153c_13c1d698 );
buf ( n5476 , R_159d_1162b198 );
buf ( n5477 , R_aa5_156b4238 );
buf ( n5478 , R_7b8_1162e9d8 );
buf ( n5479 , R_dd7_140b62b8 );
buf ( n5480 , R_10c4_12fc1878 );
buf ( n5481 , R_13f6_1700d728 );
buf ( n5482 , R_16e3_123b4d58 );
buf ( n5483 , R_1a15_13d3e998 );
buf ( n5484 , R_b0c_123c1878 );
buf ( n5485 , R_d70_13b96038 );
buf ( n5486 , R_751_13bf12b8 );
buf ( n5487 , R_112b_13d5c3b8 );
buf ( n5488 , R_138f_13df66f8 );
buf ( n5489 , R_174a_13d24658 );
buf ( n5490 , R_19ae_1587f818 );
buf ( n5491 , R_a8b_117f7898 );
buf ( n5492 , R_7d2_10082a78 );
buf ( n5493 , R_df1_15884778 );
buf ( n5494 , R_10aa_13c28458 );
buf ( n5495 , R_1410_13cd5a98 );
buf ( n5496 , R_16c9_13c03018 );
buf ( n5497 , R_1a2f_15886b18 );
buf ( n5498 , R_d7f_117f5ef8 );
buf ( n5499 , R_760_13cce6f8 );
buf ( n5500 , R_afd_156ae018 );
buf ( n5501 , R_111c_13c0f138 );
buf ( n5502 , R_139e_15ff9428 );
buf ( n5503 , R_173b_13d23758 );
buf ( n5504 , R_19bd_150e0c78 );
buf ( n5505 , R_70f_14b26038 );
buf ( n5506 , R_b4e_158835f8 );
buf ( n5507 , R_d2e_15ff2d08 );
buf ( n5508 , R_116d_14a0bc78 );
buf ( n5509 , R_134d_13cd26b8 );
buf ( n5510 , R_178c_13d39718 );
buf ( n5511 , R_196c_117ef418 );
buf ( n5512 , R_705_17018768 );
buf ( n5513 , R_b58_12fc00b8 );
buf ( n5514 , R_d24_13c0ca78 );
buf ( n5515 , R_1177_13d5b558 );
buf ( n5516 , R_1343_13d298d8 );
buf ( n5517 , R_1796_156ae338 );
buf ( n5518 , R_1962_13d5d218 );
buf ( n5519 , R_c9d_13c00ef8 );
buf ( n5520 , R_bdf_117f0638 );
buf ( n5521 , R_5c0_117ea0f8 );
buf ( n5522 , R_67e_14a0b8b8 );
buf ( n5523 , R_11fe_124c36d8 );
buf ( n5524 , R_12bc_13b981f8 );
buf ( n5525 , R_181d_123ba758 );
buf ( n5526 , R_18db_11c6d7f8 );
buf ( n5527 , R_ebc_1580cfd8 );
buf ( n5528 , R_89d_11c693d8 );
buf ( n5529 , R_9c0_13d46b98 );
buf ( n5530 , R_fdf_158176b8 );
buf ( n5531 , R_14db_156b5e58 );
buf ( n5532 , R_15fe_140b97d8 );
buf ( n5533 , R_ee1_13d40c98 );
buf ( n5534 , R_99b_156b3838 );
buf ( n5535 , R_8c2_15813518 );
buf ( n5536 , R_fba_140aebf8 );
buf ( n5537 , R_1500_1700e8a8 );
buf ( n5538 , R_15d9_13d53538 );
buf ( n5539 , R_eda_13d57638 );
buf ( n5540 , R_9a2_13c28bd8 );
buf ( n5541 , R_8bb_13d43498 );
buf ( n5542 , R_fc1_156b40f8 );
buf ( n5543 , R_14f9_13cd6178 );
buf ( n5544 , R_15e0_13cd0458 );
buf ( n5545 , R_d8b_150dc7b8 );
buf ( n5546 , R_76c_150e63f8 );
buf ( n5547 , R_af1_13b8c3f8 );
buf ( n5548 , R_1110_13d5cdb8 );
buf ( n5549 , R_13aa_14b1d898 );
buf ( n5550 , R_172f_11c6dbb8 );
buf ( n5551 , R_19c9_1509b4f8 );
buf ( n5552 , R_55a_158145f8 );
buf ( n5553 , R_6e4_11630a58 );
buf ( n5554 , R_b79_13ccfd78 );
buf ( n5555 , R_d03_124c2eb8 );
buf ( n5556 , R_1198_117f3b58 );
buf ( n5557 , R_1322_15ff6ea8 );
buf ( n5558 , R_17b7_15810bd8 );
buf ( n5559 , R_1941_117ed4d8 );
buf ( n5560 , R_6cf_1486c6d8 );
buf ( n5561 , R_56f_14a0b598 );
buf ( n5562 , R_cee_13cd9c38 );
buf ( n5563 , R_b8e_150e97d8 );
buf ( n5564 , R_11ad_13d569b8 );
buf ( n5565 , R_130d_124c3818 );
buf ( n5566 , R_17cc_117e9298 );
buf ( n5567 , R_192c_13b94918 );
buf ( n5568 , R_94b_100881f8 );
buf ( n5569 , R_f31_13c231d8 );
buf ( n5570 , R_912_11630f58 );
buf ( n5571 , R_f6a_117ea058 );
buf ( n5572 , R_1550_17014668 );
buf ( n5573 , R_1589_123b7198 );
buf ( n5574 , R_bd7_14a0ef18 );
buf ( n5575 , R_ca5_1007eb58 );
buf ( n5576 , R_5b8_170170e8 );
buf ( n5577 , R_686_15810f98 );
buf ( n5578 , R_11f6_14b22bb8 );
buf ( n5579 , R_12c4_15ff0008 );
buf ( n5580 , R_1815_156b1cb8 );
buf ( n5581 , R_18e3_13ccb9f8 );
buf ( n5582 , R_6e0_14a15f98 );
buf ( n5583 , R_55e_148707d8 );
buf ( n5584 , R_cff_14a0b458 );
buf ( n5585 , R_b7d_156b6df8 );
buf ( n5586 , R_119c_14872ad8 );
buf ( n5587 , R_131e_13dd6e38 );
buf ( n5588 , R_17bb_13bf1d58 );
buf ( n5589 , R_193d_11c70638 );
buf ( n5590 , R_d92_14b21358 );
buf ( n5591 , R_773_117f54f8 );
buf ( n5592 , R_aea_17012908 );
buf ( n5593 , R_1109_15ff3de8 );
buf ( n5594 , R_13b1_150dc358 );
buf ( n5595 , R_1728_13d5beb8 );
buf ( n5596 , R_19d0_14870af8 );
buf ( n5597 , R_e12_13b8cc18 );
buf ( n5598 , R_a6a_13d1d218 );
buf ( n5599 , R_7f3_148688f8 );
buf ( n5600 , R_1089_123b6838 );
buf ( n5601 , R_1431_15812ed8 );
buf ( n5602 , R_16a8_123bf118 );
buf ( n5603 , R_1a50_117ed6b8 );
buf ( n5604 , R_6f7_117e93d8 );
buf ( n5605 , R_b66_14a0f238 );
buf ( n5606 , R_d16_13c1b7f8 );
buf ( n5607 , R_1185_13d1ecf8 );
buf ( n5608 , R_1335_13bf1f38 );
buf ( n5609 , R_17a4_14b1ea18 );
buf ( n5610 , R_1954_15ff1ae8 );
buf ( n5611 , R_e17_13df86d8 );
buf ( n5612 , R_a65_14b22b18 );
buf ( n5613 , R_7f8_1700bec8 );
buf ( n5614 , R_1084_13d39038 );
buf ( n5615 , R_1436_15fef608 );
buf ( n5616 , R_16a3_15ff2768 );
buf ( n5617 , R_1a55_123b5898 );
buf ( n5618 , R_a21_1587bad8 );
buf ( n5619 , R_83c_13cd7398 );
buf ( n5620 , R_e5b_123bf898 );
buf ( n5621 , R_1040_1008ac78 );
buf ( n5622 , R_147a_13c04378 );
buf ( n5623 , R_165f_13cd97d8 );
buf ( n5624 , R_bfc_13d53cb8 );
buf ( n5625 , R_5dd_123b45d8 );
buf ( n5626 , R_661_13d3c2d8 );
buf ( n5627 , R_c80_1008ca78 );
buf ( n5628 , R_121b_14b24698 );
buf ( n5629 , R_129f_1008b7b8 );
buf ( n5630 , R_183a_156acc18 );
buf ( n5631 , R_18be_14a0de38 );
buf ( n5632 , R_c1b_123b48f8 );
buf ( n5633 , R_5fc_140b3518 );
buf ( n5634 , R_642_14a0d118 );
buf ( n5635 , R_c61_13c06718 );
buf ( n5636 , R_123a_15ffcf88 );
buf ( n5637 , R_1280_14a106d8 );
buf ( n5638 , R_1859_13d25378 );
buf ( n5639 , R_189f_14a13c98 );
buf ( n5640 , R_556_13d2a2d8 );
buf ( n5641 , R_6e8_12fbf4d8 );
buf ( n5642 , R_b75_156ae838 );
buf ( n5643 , R_d07_156abe58 );
buf ( n5644 , R_1194_1580f058 );
buf ( n5645 , R_1326_11c684d8 );
buf ( n5646 , R_17b3_13ddb4d8 );
buf ( n5647 , R_1945_14b22898 );
buf ( n5648 , R_bf1_13df18d8 );
buf ( n5649 , R_5d2_10088f18 );
buf ( n5650 , R_66c_123c06f8 );
buf ( n5651 , R_c8b_13c0e5f8 );
buf ( n5652 , R_1210_117f56d8 );
buf ( n5653 , R_12aa_140afb98 );
buf ( n5654 , R_182f_13d58998 );
buf ( n5655 , R_18c9_11c6eb58 );
buf ( n5656 , R_cc0_1580fcd8 );
buf ( n5657 , R_59d_13df9d58 );
buf ( n5658 , R_6a1_13cd9b98 );
buf ( n5659 , R_bbc_13d4e678 );
buf ( n5660 , R_11db_124c45d8 );
buf ( n5661 , R_12df_13d27178 );
buf ( n5662 , R_17fa_13beb8b8 );
buf ( n5663 , R_18fe_1587ca78 );
buf ( n5664 , R_d63_117f68f8 );
buf ( n5665 , R_b19_158882d8 );
buf ( n5666 , R_744_123bea38 );
buf ( n5667 , R_1138_14869ed8 );
buf ( n5668 , R_1382_13b8b958 );
buf ( n5669 , R_1757_13de1978 );
buf ( n5670 , R_19a1_123b3598 );
buf ( n5671 , R_db3_14869898 );
buf ( n5672 , R_794_17016788 );
buf ( n5673 , R_ac9_15811cb8 );
buf ( n5674 , R_10e8_140b1538 );
buf ( n5675 , R_13d2_13c292b8 );
buf ( n5676 , R_1707_13ddd9b8 );
buf ( n5677 , R_19f1_13cce518 );
buf ( n5678 , R_ecd_13d5b5f8 );
buf ( n5679 , R_9af_1587fdb8 );
buf ( n5680 , R_8ae_11631778 );
buf ( n5681 , R_fce_13c051d8 );
buf ( n5682 , R_14ec_156b01d8 );
buf ( n5683 , R_15ed_1008af98 );
buf ( n5684 , R_da4_13cd7438 );
buf ( n5685 , R_785_116381b8 );
buf ( n5686 , R_ad8_117f7a78 );
buf ( n5687 , R_10f7_1587f598 );
buf ( n5688 , R_13c3_13cd0b38 );
buf ( n5689 , R_1716_123b6bf8 );
buf ( n5690 , R_19e2_13d567d8 );
buf ( n5691 , R_58c_1587fe58 );
buf ( n5692 , R_cd1_1486dc18 );
buf ( n5693 , R_bab_13df0e38 );
buf ( n5694 , R_6b2_14867ef8 );
buf ( n5695 , R_11ca_123bd9f8 );
buf ( n5696 , R_12f0_158817f8 );
buf ( n5697 , R_17e9_123bb5b8 );
buf ( n5698 , R_190f_15881b18 );
buf ( n5699 , R_979_117efcd8 );
buf ( n5700 , R_f03_13c06f38 );
buf ( n5701 , R_8e4_123b2b98 );
buf ( n5702 , R_f98_13d588f8 );
buf ( n5703 , R_1522_15817d98 );
buf ( n5704 , R_15b7_11636bd8 );
buf ( n5705 , R_c09_14a18bf8 );
buf ( n5706 , R_5ea_1162b558 );
buf ( n5707 , R_654_150e54f8 );
buf ( n5708 , R_c73_15810958 );
buf ( n5709 , R_1228_150e4ff8 );
buf ( n5710 , R_1292_117e9fb8 );
buf ( n5711 , R_1847_13d54898 );
buf ( n5712 , R_18b1_1162ae78 );
buf ( n5713 , R_ec7_10083838 );
buf ( n5714 , R_8a8_140b6858 );
buf ( n5715 , R_9b5_156b6038 );
buf ( n5716 , R_fd4_13bef878 );
buf ( n5717 , R_14e6_123be178 );
buf ( n5718 , R_15f3_1580b958 );
buf ( n5719 , R_6dc_13d56738 );
buf ( n5720 , R_562_11630198 );
buf ( n5721 , R_cfb_156b77f8 );
buf ( n5722 , R_b81_14b23658 );
buf ( n5723 , R_11a0_117f1a38 );
buf ( n5724 , R_131a_13cd6678 );
buf ( n5725 , R_17bf_1162eed8 );
buf ( n5726 , R_1939_13b99198 );
buf ( n5727 , R_85b_150e9ff8 );
buf ( n5728 , R_e7a_13df06b8 );
buf ( n5729 , R_a02_13d20378 );
buf ( n5730 , R_1021_14873438 );
buf ( n5731 , R_1499_13c056d8 );
buf ( n5732 , R_1640_15816e98 );
buf ( n5733 , R_6c6_14b27a78 );
buf ( n5734 , R_578_13c06678 );
buf ( n5735 , R_ce5_117e9518 );
buf ( n5736 , R_b97_116328f8 );
buf ( n5737 , R_11b6_123b6478 );
buf ( n5738 , R_1304_150e5a98 );
buf ( n5739 , R_17d5_13cd9eb8 );
buf ( n5740 , R_1923_10086ad8 );
buf ( n5741 , R_aa3_123ba9d8 );
buf ( n5742 , R_7ba_17013308 );
buf ( n5743 , R_dd9_1587f4f8 );
buf ( n5744 , R_10c2_13de4358 );
buf ( n5745 , R_13f8_14866c38 );
buf ( n5746 , R_16e1_1587e058 );
buf ( n5747 , R_1a17_13d3a398 );
buf ( n5748 , R_ea3_117f04f8 );
buf ( n5749 , R_884_124c4358 );
buf ( n5750 , R_9d9_14a0c178 );
buf ( n5751 , R_ff8_14a15098 );
buf ( n5752 , R_14c2_13d50e78 );
buf ( n5753 , R_1617_13de3e58 );
buf ( n5754 , R_e0d_13c081f8 );
buf ( n5755 , R_a6f_140ab4f8 );
buf ( n5756 , R_7ee_117eb4f8 );
buf ( n5757 , R_108e_117ecf38 );
buf ( n5758 , R_142c_13d55f18 );
buf ( n5759 , R_16ad_15885df8 );
buf ( n5760 , R_1a4b_13d3a118 );
buf ( n5761 , R_e01_13b8ca38 );
buf ( n5762 , R_a7b_150e6f38 );
buf ( n5763 , R_7e2_116332f8 );
buf ( n5764 , R_109a_140adc58 );
buf ( n5765 , R_1420_1580acd8 );
buf ( n5766 , R_16b9_13b972f8 );
buf ( n5767 , R_1a3f_13cd8f18 );
buf ( n5768 , R_597_156aeab8 );
buf ( n5769 , R_cc6_1486fd38 );
buf ( n5770 , R_bb6_13d58fd8 );
buf ( n5771 , R_6a7_140b7938 );
buf ( n5772 , R_11d5_14871bd8 );
buf ( n5773 , R_12e5_14b28bf8 );
buf ( n5774 , R_17f4_156b4cd8 );
buf ( n5775 , R_1904_140b9058 );
buf ( n5776 , R_dfa_1486ff18 );
buf ( n5777 , R_a82_116368b8 );
buf ( n5778 , R_7db_150dd1b8 );
buf ( n5779 , R_10a1_123b8598 );
buf ( n5780 , R_1419_13df1b58 );
buf ( n5781 , R_16c0_13b994b8 );
buf ( n5782 , R_1a38_13ccab98 );
buf ( n5783 , R_911_14b22078 );
buf ( n5784 , R_94c_123bc7d8 );
buf ( n5785 , R_f30_12fbf898 );
buf ( n5786 , R_f6b_13c0a6d8 );
buf ( n5787 , R_154f_1700ea88 );
buf ( n5788 , R_158a_13c25758 );
buf ( n5789 , R_d44_13b99418 );
buf ( n5790 , R_b38_13d23618 );
buf ( n5791 , R_725_13d4f618 );
buf ( n5792 , R_1157_14a13298 );
buf ( n5793 , R_1363_124c4718 );
buf ( n5794 , R_1776_15882518 );
buf ( n5795 , R_1982_15816fd8 );
buf ( n5796 , R_983_1700b4c8 );
buf ( n5797 , R_ef9_1007e338 );
buf ( n5798 , R_8da_1587ba38 );
buf ( n5799 , R_fa2_15ffaf08 );
buf ( n5800 , R_1518_13c09ff8 );
buf ( n5801 , R_15c1_13c1e138 );
buf ( n5802 , R_d41_13bf8f18 );
buf ( n5803 , R_722_14b26fd8 );
buf ( n5804 , R_b3b_14a0f378 );
buf ( n5805 , R_115a_156af9b8 );
buf ( n5806 , R_1360_156aa5f8 );
buf ( n5807 , R_1779_13dec3d8 );
buf ( n5808 , R_197f_1700ba68 );
buf ( n5809 , R_7fd_13d29658 );
buf ( n5810 , R_e1c_156b8158 );
buf ( n5811 , R_a60_124c2738 );
buf ( n5812 , R_107f_13d55ab8 );
buf ( n5813 , R_143b_13cd5458 );
buf ( n5814 , R_169e_13d59618 );
buf ( n5815 , R_1a5a_117ecd58 );
buf ( n5816 , R_a94_158121b8 );
buf ( n5817 , R_7c9_13c1bb18 );
buf ( n5818 , R_de8_13df22d8 );
buf ( n5819 , R_10b3_17011328 );
buf ( n5820 , R_1407_140b9cd8 );
buf ( n5821 , R_16d2_150e0098 );
buf ( n5822 , R_1a26_14868678 );
buf ( n5823 , R_e9a_14a0e1f8 );
buf ( n5824 , R_87b_123b2e18 );
buf ( n5825 , R_9e2_148680d8 );
buf ( n5826 , R_1001_100877f8 );
buf ( n5827 , R_14b9_150dda78 );
buf ( n5828 , R_1620_117efff8 );
buf ( n5829 , R_bc2_1580b098 );
buf ( n5830 , R_cba_13c20118 );
buf ( n5831 , R_5a3_13b98298 );
buf ( n5832 , R_69b_13bf94b8 );
buf ( n5833 , R_11e1_1486a798 );
buf ( n5834 , R_12d9_123ba118 );
buf ( n5835 , R_1800_15888378 );
buf ( n5836 , R_18f8_156ac538 );
buf ( n5837 , R_960_13ccf418 );
buf ( n5838 , R_f1c_13df79b8 );
buf ( n5839 , R_8fd_123b6fb8 );
buf ( n5840 , R_f7f_140aa558 );
buf ( n5841 , R_153b_117f5d18 );
buf ( n5842 , R_159e_14871db8 );
buf ( n5843 , R_d47_13d27998 );
buf ( n5844 , R_b35_1587cc58 );
buf ( n5845 , R_728_140ba318 );
buf ( n5846 , R_1154_117e95b8 );
buf ( n5847 , R_1366_17015568 );
buf ( n5848 , R_1773_156ac2b8 );
buf ( n5849 , R_1985_1162c3b8 );
buf ( n5850 , R_b11_15883698 );
buf ( n5851 , R_d6b_123b8958 );
buf ( n5852 , R_74c_150e17b8 );
buf ( n5853 , R_1130_13bef0f8 );
buf ( n5854 , R_138a_13d25cd8 );
buf ( n5855 , R_174f_13df2058 );
buf ( n5856 , R_19a9_1486eed8 );
buf ( n5857 , R_6ec_13c03b58 );
buf ( n5858 , R_b71_140afd78 );
buf ( n5859 , R_d0b_1587d158 );
buf ( n5860 , R_1190_13c09198 );
buf ( n5861 , R_132a_13d44bb8 );
buf ( n5862 , R_17af_123b9d58 );
buf ( n5863 , R_1949_140b51d8 );
buf ( n5864 , R_815_158140f8 );
buf ( n5865 , R_a48_13bed6b8 );
buf ( n5866 , R_e34_13cd7e38 );
buf ( n5867 , R_1067_13b93ab8 );
buf ( n5868 , R_1453_15ff99c8 );
buf ( n5869 , R_1686_1008c258 );
buf ( n5870 , R_af8_148696b8 );
buf ( n5871 , R_d84_156b3e78 );
buf ( n5872 , R_765_13df9678 );
buf ( n5873 , R_1117_140b2398 );
buf ( n5874 , R_13a3_123bd598 );
buf ( n5875 , R_1736_117f1218 );
buf ( n5876 , R_19c2_14871098 );
buf ( n5877 , R_d3e_14870198 );
buf ( n5878 , R_71f_123b6e78 );
buf ( n5879 , R_b3e_11631138 );
buf ( n5880 , R_115d_1008bd58 );
buf ( n5881 , R_135d_13cd9d78 );
buf ( n5882 , R_177c_11629258 );
buf ( n5883 , R_197c_13bec8f8 );
buf ( n5884 , R_96e_1162bff8 );
buf ( n5885 , R_f0e_17010f68 );
buf ( n5886 , R_8ef_13dd96d8 );
buf ( n5887 , R_f8d_13cd51d8 );
buf ( n5888 , R_152d_13d1f8d8 );
buf ( n5889 , R_15ac_12fc1418 );
buf ( n5890 , R_ee8_13d55658 );
buf ( n5891 , R_994_13c086f8 );
buf ( n5892 , R_8c9_1162f838 );
buf ( n5893 , R_fb3_11c6c7b8 );
buf ( n5894 , R_1507_14b218f8 );
buf ( n5895 , R_15d2_11c6e978 );
buf ( n5896 , R_ed3_13b93018 );
buf ( n5897 , R_9a9_140ac3f8 );
buf ( n5898 , R_8b4_150e2e38 );
buf ( n5899 , R_fc8_14875238 );
buf ( n5900 , R_14f2_13cd1718 );
buf ( n5901 , R_15e7_150e0e58 );
buf ( n5902 , R_c1a_13d3c198 );
buf ( n5903 , R_5fb_156b22f8 );
buf ( n5904 , R_643_117ea698 );
buf ( n5905 , R_c62_1162c598 );
buf ( n5906 , R_1239_15817938 );
buf ( n5907 , R_1281_158887d8 );
buf ( n5908 , R_1858_13bea9b8 );
buf ( n5909 , R_18a0_123bfcf8 );
buf ( n5910 , R_98c_13c21f18 );
buf ( n5911 , R_ef0_13d51418 );
buf ( n5912 , R_8d1_12fc06f8 );
buf ( n5913 , R_fab_14a127f8 );
buf ( n5914 , R_150f_15817398 );
buf ( n5915 , R_15ca_156b71b8 );
buf ( n5916 , R_c95_123be2b8 );
buf ( n5917 , R_be7_1162d858 );
buf ( n5918 , R_5c8_15feeca8 );
buf ( n5919 , R_676_13d37e18 );
buf ( n5920 , R_1206_13ddcc98 );
buf ( n5921 , R_12b4_10087938 );
buf ( n5922 , R_1825_1486a298 );
buf ( n5923 , R_18d3_17018f88 );
buf ( n5924 , R_d5b_150e0958 );
buf ( n5925 , R_b21_14b21e98 );
buf ( n5926 , R_73c_13bec858 );
buf ( n5927 , R_1140_13b98798 );
buf ( n5928 , R_137a_13dd7018 );
buf ( n5929 , R_175f_15ff7f88 );
buf ( n5930 , R_1999_117f2118 );
buf ( n5931 , R_d4a_13df40d8 );
buf ( n5932 , R_b32_13c268d8 );
buf ( n5933 , R_72b_11632c18 );
buf ( n5934 , R_1151_11638898 );
buf ( n5935 , R_1369_117f5138 );
buf ( n5936 , R_1770_124c2a58 );
buf ( n5937 , R_1988_150dfaf8 );
buf ( n5938 , R_db1_13bf06d8 );
buf ( n5939 , R_792_13ccb638 );
buf ( n5940 , R_acb_13d2a378 );
buf ( n5941 , R_10ea_13d2b598 );
buf ( n5942 , R_13d0_1700b388 );
buf ( n5943 , R_1709_1162a298 );
buf ( n5944 , R_19ef_150de1f8 );
buf ( n5945 , R_ae3_14b24738 );
buf ( n5946 , R_d99_156abef8 );
buf ( n5947 , R_77a_13c0f3b8 );
buf ( n5948 , R_1102_11632358 );
buf ( n5949 , R_13b8_13c29c18 );
buf ( n5950 , R_1721_14870f58 );
buf ( n5951 , R_19d7_13de38b8 );
buf ( n5952 , R_6d8_1580ebf8 );
buf ( n5953 , R_566_140b4f58 );
buf ( n5954 , R_cf7_13d26778 );
buf ( n5955 , R_b85_13df3958 );
buf ( n5956 , R_11a4_140b1178 );
buf ( n5957 , R_1316_13c24718 );
buf ( n5958 , R_17c3_13df1e78 );
buf ( n5959 , R_1935_14a13798 );
buf ( n5960 , R_a0d_14a0f198 );
buf ( n5961 , R_850_1700cbe8 );
buf ( n5962 , R_e6f_117ee6f8 );
buf ( n5963 , R_102c_156ae3d8 );
buf ( n5964 , R_148e_17014208 );
buf ( n5965 , R_164b_123b8638 );
buf ( n5966 , R_f2f_13ccded8 );
buf ( n5967 , R_910_158144b8 );
buf ( n5968 , R_94d_13de1dd8 );
buf ( n5969 , R_f6c_140aca38 );
buf ( n5970 , R_154e_158131f8 );
buf ( n5971 , R_158b_123b5078 );
buf ( n5972 , R_70c_1162a338 );
buf ( n5973 , R_b51_13df4c18 );
buf ( n5974 , R_d2b_123bacf8 );
buf ( n5975 , R_1170_13ddca18 );
buf ( n5976 , R_134a_123bdb38 );
buf ( n5977 , R_178f_14a0df78 );
buf ( n5978 , R_1969_13c0e918 );
buf ( n5979 , R_ec1_13c0ddd8 );
buf ( n5980 , R_8a2_13dd9638 );
buf ( n5981 , R_9bb_14a13d38 );
buf ( n5982 , R_fda_14876098 );
buf ( n5983 , R_14e0_117ea9b8 );
buf ( n5984 , R_15f9_13d4fcf8 );
buf ( n5985 , R_d3b_150e4a58 );
buf ( n5986 , R_71c_150dba98 );
buf ( n5987 , R_b41_100844b8 );
buf ( n5988 , R_1160_14a16498 );
buf ( n5989 , R_135a_156b8838 );
buf ( n5990 , R_177f_13ccedd8 );
buf ( n5991 , R_1979_156ad7f8 );
buf ( n5992 , R_80a_11c686b8 );
buf ( n5993 , R_a53_13d54ed8 );
buf ( n5994 , R_e29_124c3138 );
buf ( n5995 , R_1072_13d5c598 );
buf ( n5996 , R_1448_156b5098 );
buf ( n5997 , R_1691_13bf8478 );
buf ( n5998 , R_1a67_13d3a898 );
buf ( n5999 , R_aa1_13ccbd18 );
buf ( n6000 , R_7bc_13ccc218 );
buf ( n6001 , R_ddb_15812618 );
buf ( n6002 , R_10c0_15816d58 );
buf ( n6003 , R_13fa_14b29a58 );
buf ( n6004 , R_16df_10084eb8 );
buf ( n6005 , R_1a19_11c70a98 );
buf ( n6006 , R_a1e_13de1338 );
buf ( n6007 , R_83f_123bc5f8 );
buf ( n6008 , R_e5e_13c25258 );
buf ( n6009 , R_103d_123b2738 );
buf ( n6010 , R_147d_13d53e98 );
buf ( n6011 , R_165c_123b57f8 );
buf ( n6012 , R_c74_14b242d8 );
buf ( n6013 , R_c08_13ded7d8 );
buf ( n6014 , R_5e9_15816178 );
buf ( n6015 , R_655_13c026b8 );
buf ( n6016 , R_1227_123b72d8 );
buf ( n6017 , R_1293_1008c6b8 );
buf ( n6018 , R_1846_13c22af8 );
buf ( n6019 , R_18b2_150dd4d8 );
buf ( n6020 , R_a14_11632038 );
buf ( n6021 , R_849_123c1af8 );
buf ( n6022 , R_e68_15887658 );
buf ( n6023 , R_1033_13bf8518 );
buf ( n6024 , R_1487_1007fc38 );
buf ( n6025 , R_1652_11635418 );
buf ( n6026 , R_68e_11630eb8 );
buf ( n6027 , R_bcf_1486c4f8 );
buf ( n6028 , R_cad_150e5c78 );
buf ( n6029 , R_5b0_13d20c38 );
buf ( n6030 , R_11ee_13df5938 );
buf ( n6031 , R_12cc_156aee78 );
buf ( n6032 , R_180d_13d29dd8 );
buf ( n6033 , R_18eb_13cd2bb8 );
buf ( n6034 , R_7e9_13b903b8 );
buf ( n6035 , R_e08_14a11498 );
buf ( n6036 , R_a74_13c02a78 );
buf ( n6037 , R_1093_123bddb8 );
buf ( n6038 , R_1427_1580dd98 );
buf ( n6039 , R_16b2_123b89f8 );
buf ( n6040 , R_1a46_150dff58 );
buf ( n6041 , R_c81_140ac718 );
buf ( n6042 , R_bfb_117e8f78 );
buf ( n6043 , R_5dc_13cd21b8 );
buf ( n6044 , R_662_11c6af58 );
buf ( n6045 , R_121a_13dd6bb8 );
buf ( n6046 , R_12a0_156af7d8 );
buf ( n6047 , R_1839_10083a18 );
buf ( n6048 , R_18bf_13cd63f8 );
buf ( n6049 , R_d4d_14b1c218 );
buf ( n6050 , R_b2f_14a168f8 );
buf ( n6051 , R_72e_15885178 );
buf ( n6052 , R_114e_14866878 );
buf ( n6053 , R_136c_13d5ce58 );
buf ( n6054 , R_176d_15883e18 );
buf ( n6055 , R_198b_123ba938 );
buf ( n6056 , R_bb0_11635198 );
buf ( n6057 , R_6ad_14b295f8 );
buf ( n6058 , R_591_123b56b8 );
buf ( n6059 , R_ccc_13c02f78 );
buf ( n6060 , R_11cf_13dedd78 );
buf ( n6061 , R_12eb_156ab598 );
buf ( n6062 , R_17ee_117f2a78 );
buf ( n6063 , R_190a_1162b238 );
buf ( n6064 , R_7d4_14a0fe18 );
buf ( n6065 , R_df3_14b1e478 );
buf ( n6066 , R_a89_13dd9278 );
buf ( n6067 , R_10a8_13d52958 );
buf ( n6068 , R_1412_11c6f198 );
buf ( n6069 , R_16c7_13d27d58 );
buf ( n6070 , R_1a31_140b9d78 );
buf ( n6071 , R_c19_1700d408 );
buf ( n6072 , R_5fa_13df88b8 );
buf ( n6073 , R_644_13d23938 );
buf ( n6074 , R_c63_1162e258 );
buf ( n6075 , R_1238_13df9a38 );
buf ( n6076 , R_1282_13c2acf8 );
buf ( n6077 , R_1857_13cd2ed8 );
buf ( n6078 , R_18a1_156aefb8 );
buf ( n6079 , R_6f0_140ae658 );
buf ( n6080 , R_b6d_123b4178 );
buf ( n6081 , R_d0f_150df0f8 );
buf ( n6082 , R_118c_14a17898 );
buf ( n6083 , R_132e_13bed758 );
buf ( n6084 , R_17ab_13cd0d18 );
buf ( n6085 , R_194d_1008c438 );
buf ( n6086 , R_802_13d3e5d8 );
buf ( n6087 , R_e21_14a0aaf8 );
buf ( n6088 , R_a5b_13bf7e38 );
buf ( n6089 , R_107a_13d1ed98 );
buf ( n6090 , R_1440_124c4d58 );
buf ( n6091 , R_1699_140b0318 );
buf ( n6092 , R_1a5f_124c5618 );
buf ( n6093 , R_8fc_13bebd18 );
buf ( n6094 , R_961_12fbe358 );
buf ( n6095 , R_f1b_13ddafd8 );
buf ( n6096 , R_f80_1486f478 );
buf ( n6097 , R_153a_116341f8 );
buf ( n6098 , R_159f_1008d338 );
buf ( n6099 , R_ada_15812f78 );
buf ( n6100 , R_da2_156b5ef8 );
buf ( n6101 , R_783_123ba898 );
buf ( n6102 , R_10f9_123b7a58 );
buf ( n6103 , R_13c1_13d3bfb8 );
buf ( n6104 , R_1718_156b8018 );
buf ( n6105 , R_19e0_13dd4ef8 );
buf ( n6106 , R_6cb_117f2258 );
buf ( n6107 , R_573_1162dfd8 );
buf ( n6108 , R_cea_13d5be18 );
buf ( n6109 , R_b92_13c01998 );
buf ( n6110 , R_11b1_1700a208 );
buf ( n6111 , R_1309_117e8898 );
buf ( n6112 , R_17d0_156b8d38 );
buf ( n6113 , R_1928_14a0f738 );
buf ( n6114 , R_eb1_156b8f18 );
buf ( n6115 , R_892_11c69018 );
buf ( n6116 , R_9cb_13bed1b8 );
buf ( n6117 , R_fea_13d2b3b8 );
buf ( n6118 , R_14d0_13ccf698 );
buf ( n6119 , R_1609_13cd30b8 );
buf ( n6120 , R_67f_13cd88d8 );
buf ( n6121 , R_c9e_1580ee78 );
buf ( n6122 , R_bde_123b3138 );
buf ( n6123 , R_5bf_117f0b38 );
buf ( n6124 , R_11fd_1162f3d8 );
buf ( n6125 , R_12bd_13bf9698 );
buf ( n6126 , R_181c_13bf7758 );
buf ( n6127 , R_18dc_15817258 );
buf ( n6128 , R_c8c_13b97258 );
buf ( n6129 , R_bf0_13c26d38 );
buf ( n6130 , R_5d1_14875af8 );
buf ( n6131 , R_66d_1700eda8 );
buf ( n6132 , R_120f_156b0a98 );
buf ( n6133 , R_12ab_1486c278 );
buf ( n6134 , R_182e_116366d8 );
buf ( n6135 , R_18ca_11c708b8 );
buf ( n6136 , R_f2e_13dddb98 );
buf ( n6137 , R_90f_13b8e3d8 );
buf ( n6138 , R_94e_117f3c98 );
buf ( n6139 , R_f6d_13bf7a78 );
buf ( n6140 , R_154d_13df8c78 );
buf ( n6141 , R_158c_13d278f8 );
buf ( n6142 , R_702_13de3598 );
buf ( n6143 , R_b5b_13d45bf8 );
buf ( n6144 , R_d21_156ac038 );
buf ( n6145 , R_117a_14b292d8 );
buf ( n6146 , R_1340_123bbab8 );
buf ( n6147 , R_1799_13df1018 );
buf ( n6148 , R_195f_13b92e38 );
buf ( n6149 , R_d38_156afaf8 );
buf ( n6150 , R_719_13d1d498 );
buf ( n6151 , R_b44_13df7238 );
buf ( n6152 , R_1163_13b91358 );
buf ( n6153 , R_1357_13d5bcd8 );
buf ( n6154 , R_1782_1486c138 );
buf ( n6155 , R_1976_14b1de38 );
buf ( n6156 , R_695_13b93b58 );
buf ( n6157 , R_bc8_13dfb3d8 );
buf ( n6158 , R_cb4_15817078 );
buf ( n6159 , R_5a9_156b6998 );
buf ( n6160 , R_11e7_13bf3298 );
buf ( n6161 , R_12d3_14b28338 );
buf ( n6162 , R_1806_123b6dd8 );
buf ( n6163 , R_18f2_13d40338 );
buf ( n6164 , R_a06_158876f8 );
buf ( n6165 , R_857_14874dd8 );
buf ( n6166 , R_e76_13bf0958 );
buf ( n6167 , R_1025_13d59438 );
buf ( n6168 , R_1495_14870238 );
buf ( n6169 , R_1644_15ff4d88 );
buf ( n6170 , R_6fb_156b9378 );
buf ( n6171 , R_b62_123bb298 );
buf ( n6172 , R_d1a_117ee1f8 );
buf ( n6173 , R_1181_148748d8 );
buf ( n6174 , R_1339_1580de38 );
buf ( n6175 , R_17a0_13dd7478 );
buf ( n6176 , R_1958_156ae5b8 );
buf ( n6177 , R_97a_117eaff8 );
buf ( n6178 , R_f02_13d538f8 );
buf ( n6179 , R_8e3_13c107b8 );
buf ( n6180 , R_f99_1580efb8 );
buf ( n6181 , R_1521_148676d8 );
buf ( n6182 , R_15b8_13b93e78 );
buf ( n6183 , R_829_13b954f8 );
buf ( n6184 , R_a34_156b03b8 );
buf ( n6185 , R_e48_15813d38 );
buf ( n6186 , R_1053_13cd3478 );
buf ( n6187 , R_1467_13b8be58 );
buf ( n6188 , R_1672_13cd1df8 );
buf ( n6189 , R_e89_13de0078 );
buf ( n6190 , R_9f3_156b0598 );
buf ( n6191 , R_86a_13b94378 );
buf ( n6192 , R_1012_123bf618 );
buf ( n6193 , R_14a8_13becdf8 );
buf ( n6194 , R_1631_1486c9f8 );
buf ( n6195 , R_acd_1008bfd8 );
buf ( n6196 , R_daf_123b59d8 );
buf ( n6197 , R_790_13d2bd18 );
buf ( n6198 , R_10ec_1700b6a8 );
buf ( n6199 , R_13ce_13df2a58 );
buf ( n6200 , R_170b_14b26178 );
buf ( n6201 , R_19ed_148709b8 );
buf ( n6202 , R_a31_13cd7d98 );
buf ( n6203 , R_82c_140b1e98 );
buf ( n6204 , R_e4b_116316d8 );
buf ( n6205 , R_1050_13d3d138 );
buf ( n6206 , R_146a_123bd318 );
buf ( n6207 , R_166f_140ad118 );
buf ( n6208 , R_eac_1007f418 );
buf ( n6209 , R_88d_13bf99b8 );
buf ( n6210 , R_9d0_17010748 );
buf ( n6211 , R_fef_1580b138 );
buf ( n6212 , R_14cb_13d44258 );
buf ( n6213 , R_160e_11632a38 );
buf ( n6214 , R_826_13c24cb8 );
buf ( n6215 , R_a37_158112b8 );
buf ( n6216 , R_e45_15fee168 );
buf ( n6217 , R_1056_15fedc68 );
buf ( n6218 , R_1464_13d3fa78 );
buf ( n6219 , R_1675_14b28dd8 );
buf ( n6220 , R_eb6_11c69518 );
buf ( n6221 , R_897_11c69338 );
buf ( n6222 , R_9c6_156ad258 );
buf ( n6223 , R_fe5_14b1f4b8 );
buf ( n6224 , R_14d5_14871a98 );
buf ( n6225 , R_1604_13beed38 );
buf ( n6226 , R_9ef_14a126b8 );
buf ( n6227 , R_e8d_13c07578 );
buf ( n6228 , R_86e_13ded738 );
buf ( n6229 , R_100e_100810d8 );
buf ( n6230 , R_14ac_13cce158 );
buf ( n6231 , R_162d_13c0adb8 );
buf ( n6232 , R_7cb_14a0acd8 );
buf ( n6233 , R_dea_123c0798 );
buf ( n6234 , R_a92_13d25238 );
buf ( n6235 , R_10b1_13d55478 );
buf ( n6236 , R_1409_1587f638 );
buf ( n6237 , R_16d0_13c02ed8 );
buf ( n6238 , R_1a28_14a12398 );
buf ( n6239 , R_ee0_13d1ffb8 );
buf ( n6240 , R_99c_14a0f418 );
buf ( n6241 , R_8c1_14b25818 );
buf ( n6242 , R_fbb_123b70f8 );
buf ( n6243 , R_14ff_1580bf98 );
buf ( n6244 , R_15da_140ba138 );
buf ( n6245 , R_687_14b23fb8 );
buf ( n6246 , R_bd6_13dd71f8 );
buf ( n6247 , R_ca6_123bd098 );
buf ( n6248 , R_5b7_117e8cf8 );
buf ( n6249 , R_11f5_15815318 );
buf ( n6250 , R_12c5_14a0f7d8 );
buf ( n6251 , R_1814_170116e8 );
buf ( n6252 , R_18e4_12fc1d78 );
buf ( n6253 , R_812_12fc0018 );
buf ( n6254 , R_a4b_13bf22f8 );
buf ( n6255 , R_e31_13bee338 );
buf ( n6256 , R_106a_13d56a58 );
buf ( n6257 , R_1450_1580a738 );
buf ( n6258 , R_1689_14a0c218 );
buf ( n6259 , R_e85_156aa878 );
buf ( n6260 , R_9f7_13d246f8 );
buf ( n6261 , R_866_15ffb868 );
buf ( n6262 , R_1016_156af698 );
buf ( n6263 , R_14a4_11c6ec98 );
buf ( n6264 , R_1635_15ff7588 );
buf ( n6265 , R_8ee_140ae338 );
buf ( n6266 , R_96f_13d3b8d8 );
buf ( n6267 , R_f0d_13d4fa78 );
buf ( n6268 , R_f8e_13d541b8 );
buf ( n6269 , R_152c_156b2258 );
buf ( n6270 , R_15ad_13d58218 );
buf ( n6271 , R_9de_124c3458 );
buf ( n6272 , R_e9e_123b9038 );
buf ( n6273 , R_87f_117f0958 );
buf ( n6274 , R_ffd_13c27f58 );
buf ( n6275 , R_14bd_13cd71b8 );
buf ( n6276 , R_161c_156b6178 );
buf ( n6277 , R_aec_14866b98 );
buf ( n6278 , R_d90_10081718 );
buf ( n6279 , R_771_1007ee78 );
buf ( n6280 , R_110b_14b24f58 );
buf ( n6281 , R_13af_158110d8 );
buf ( n6282 , R_172a_11c6feb8 );
buf ( n6283 , R_19ce_11c6fc38 );
buf ( n6284 , R_6d4_15ff47e8 );
buf ( n6285 , R_56a_17018268 );
buf ( n6286 , R_cf3_150e21b8 );
buf ( n6287 , R_b89_13cd67b8 );
buf ( n6288 , R_11a8_13c0ab38 );
buf ( n6289 , R_1312_15881758 );
buf ( n6290 , R_17c7_1580cf38 );
buf ( n6291 , R_1931_11c6b4f8 );
buf ( n6292 , R_7be_13d51918 );
buf ( n6293 , R_ddd_10083fb8 );
buf ( n6294 , R_a9f_140b7b18 );
buf ( n6295 , R_10be_1162c138 );
buf ( n6296 , R_13fc_13b967b8 );
buf ( n6297 , R_16dd_15ffb728 );
buf ( n6298 , R_1a1b_13d3ab18 );
buf ( n6299 , R_a2e_1580aeb8 );
buf ( n6300 , R_82f_14b26cb8 );
buf ( n6301 , R_e4e_13dec798 );
buf ( n6302 , R_104d_13de2af8 );
buf ( n6303 , R_146d_156b1998 );
buf ( n6304 , R_166c_117f5958 );
buf ( n6305 , R_d50_156b51d8 );
buf ( n6306 , R_b2c_12fc0478 );
buf ( n6307 , R_731_15ffaa08 );
buf ( n6308 , R_114b_13ddbed8 );
buf ( n6309 , R_136f_11c6c718 );
buf ( n6310 , R_176a_11628f38 );
buf ( n6311 , R_198e_150e3518 );
buf ( n6312 , R_ed9_15ff7948 );
buf ( n6313 , R_9a3_13c1fad8 );
buf ( n6314 , R_8ba_116386b8 );
buf ( n6315 , R_fc2_1700f7a8 );
buf ( n6316 , R_14f8_117f15d8 );
buf ( n6317 , R_15e1_150dcd58 );
buf ( n6318 , R_b16_13c1c1f8 );
buf ( n6319 , R_d66_13b8b1d8 );
buf ( n6320 , R_747_158864d8 );
buf ( n6321 , R_1135_156b68f8 );
buf ( n6322 , R_1385_1580b278 );
buf ( n6323 , R_1754_156add98 );
buf ( n6324 , R_19a4_13d4fd98 );
buf ( n6325 , R_823_11c6f2d8 );
buf ( n6326 , R_a3a_14871318 );
buf ( n6327 , R_e42_156ade38 );
buf ( n6328 , R_1059_13c0f318 );
buf ( n6329 , R_1461_14a1a138 );
buf ( n6330 , R_1678_14a0fd78 );
buf ( n6331 , R_8d9_158837d8 );
buf ( n6332 , R_984_15882d38 );
buf ( n6333 , R_ef8_15816998 );
buf ( n6334 , R_fa3_15815458 );
buf ( n6335 , R_1517_156ad898 );
buf ( n6336 , R_15c2_11630c38 );
buf ( n6337 , R_af3_13beae18 );
buf ( n6338 , R_d89_117e8938 );
buf ( n6339 , R_76a_123bceb8 );
buf ( n6340 , R_1112_13c20c58 );
buf ( n6341 , R_13a8_117f4a58 );
buf ( n6342 , R_1731_1008a818 );
buf ( n6343 , R_19c7_13d38bd8 );
buf ( n6344 , R_b04_156aed38 );
buf ( n6345 , R_d78_13cd7758 );
buf ( n6346 , R_759_11629938 );
buf ( n6347 , R_1123_15ffb908 );
buf ( n6348 , R_1397_13d37a58 );
buf ( n6349 , R_1742_13d237f8 );
buf ( n6350 , R_19b6_14b20778 );
buf ( n6351 , R_c64_13c1fdf8 );
buf ( n6352 , R_c18_12fc23b8 );
buf ( n6353 , R_5f9_13b8f238 );
buf ( n6354 , R_645_140b2118 );
buf ( n6355 , R_1237_1162dad8 );
buf ( n6356 , R_1283_14a18798 );
buf ( n6357 , R_1856_117f4878 );
buf ( n6358 , R_18a2_13d53998 );
buf ( n6359 , R_f2d_100818f8 );
buf ( n6360 , R_90e_11629898 );
buf ( n6361 , R_94f_15888738 );
buf ( n6362 , R_f6e_14a188d8 );
buf ( n6363 , R_154c_14a147d8 );
buf ( n6364 , R_158d_15ff0a08 );
buf ( n6365 , R_9eb_117ef2d8 );
buf ( n6366 , R_e91_1580e3d8 );
buf ( n6367 , R_872_13c0c7f8 );
buf ( n6368 , R_100a_117f81f8 );
buf ( n6369 , R_14b0_124c2f58 );
buf ( n6370 , R_1629_14a0b6d8 );
buf ( n6371 , R_656_15886bb8 );
buf ( n6372 , R_c75_156b0db8 );
buf ( n6373 , R_c07_124c4cb8 );
buf ( n6374 , R_5e8_1162f298 );
buf ( n6375 , R_1226_13b8e018 );
buf ( n6376 , R_1294_13b91ad8 );
buf ( n6377 , R_1845_13cd83d8 );
buf ( n6378 , R_18b3_13d1e118 );
buf ( n6379 , R_ba0_156b4698 );
buf ( n6380 , R_6bd_13c0ec38 );
buf ( n6381 , R_581_13d1d8f8 );
buf ( n6382 , R_cdc_13cd9378 );
buf ( n6383 , R_11bf_123b6c98 );
buf ( n6384 , R_12fb_150e3018 );
buf ( n6385 , R_17de_14b20458 );
buf ( n6386 , R_191a_123b2cd8 );
buf ( n6387 , R_d5e_14a10278 );
buf ( n6388 , R_b1e_13df7418 );
buf ( n6389 , R_73f_1587b998 );
buf ( n6390 , R_113d_13d58498 );
buf ( n6391 , R_137d_14a11b78 );
buf ( n6392 , R_175c_1587b218 );
buf ( n6393 , R_199c_17017408 );
buf ( n6394 , R_b09_15884f98 );
buf ( n6395 , R_d73_1580b4f8 );
buf ( n6396 , R_754_15811d58 );
buf ( n6397 , R_1128_10084d78 );
buf ( n6398 , R_1392_14a15db8 );
buf ( n6399 , R_1747_17018588 );
buf ( n6400 , R_19b1_13dd9f98 );
buf ( n6401 , R_d35_14a11858 );
buf ( n6402 , R_716_156b9c38 );
buf ( n6403 , R_b47_140af4b8 );
buf ( n6404 , R_1166_13ccdcf8 );
buf ( n6405 , R_1354_13d41738 );
buf ( n6406 , R_1785_1162d218 );
buf ( n6407 , R_1973_14a18338 );
buf ( n6408 , R_a2b_13c1e6d8 );
buf ( n6409 , R_832_13df5c58 );
buf ( n6410 , R_e51_156ab278 );
buf ( n6411 , R_104a_14a108b8 );
buf ( n6412 , R_1470_15887bf8 );
buf ( n6413 , R_1669_158828d8 );
buf ( n6414 , R_e81_1007dc58 );
buf ( n6415 , R_9fb_1486fb58 );
buf ( n6416 , R_862_156ab138 );
buf ( n6417 , R_101a_13d5a798 );
buf ( n6418 , R_14a0_13d38818 );
buf ( n6419 , R_1639_1162abf8 );
buf ( n6420 , R_ba5_140b4af8 );
buf ( n6421 , R_6b8_1580d898 );
buf ( n6422 , R_586_15ff8488 );
buf ( n6423 , R_cd7_156b7e38 );
buf ( n6424 , R_11c4_117ecad8 );
buf ( n6425 , R_12f6_17015ba8 );
buf ( n6426 , R_17e3_13c1dd78 );
buf ( n6427 , R_1915_14a17f78 );
buf ( n6428 , R_aff_140aba98 );
buf ( n6429 , R_d7d_148714f8 );
buf ( n6430 , R_75e_10084418 );
buf ( n6431 , R_111e_11635918 );
buf ( n6432 , R_139c_1580e0b8 );
buf ( n6433 , R_173d_13deffd8 );
buf ( n6434 , R_19bb_13df9df8 );
buf ( n6435 , R_7dd_13d28898 );
buf ( n6436 , R_dfc_156b9ff8 );
buf ( n6437 , R_a80_13ddc8d8 );
buf ( n6438 , R_109f_13cd2cf8 );
buf ( n6439 , R_141b_12fc10f8 );
buf ( n6440 , R_16be_13bf0098 );
buf ( n6441 , R_1a3a_156b79d8 );
buf ( n6442 , R_9d5_15ff1908 );
buf ( n6443 , R_ea7_14a124d8 );
buf ( n6444 , R_888_13deebd8 );
buf ( n6445 , R_ff4_13cd7b18 );
buf ( n6446 , R_14c6_13cd5d18 );
buf ( n6447 , R_1613_123bc198 );
buf ( n6448 , R_677_13c0c758 );
buf ( n6449 , R_c96_13c0d838 );
buf ( n6450 , R_be6_1162cf98 );
buf ( n6451 , R_5c7_1162f1f8 );
buf ( n6452 , R_1205_156b94b8 );
buf ( n6453 , R_12b5_158816b8 );
buf ( n6454 , R_1824_13c04f58 );
buf ( n6455 , R_18d4_13beb958 );
buf ( n6456 , R_f1a_124c4f38 );
buf ( n6457 , R_8fb_13c1e9f8 );
buf ( n6458 , R_962_14a15ef8 );
buf ( n6459 , R_f81_1580d438 );
buf ( n6460 , R_1539_14b267b8 );
buf ( n6461 , R_15a0_15ff32a8 );
buf ( n6462 , R_d28_156b3fb8 );
buf ( n6463 , R_709_117ea4b8 );
buf ( n6464 , R_b54_13c04c38 );
buf ( n6465 , R_1173_15810778 );
buf ( n6466 , R_1347_13dd5f38 );
buf ( n6467 , R_1792_13d39858 );
buf ( n6468 , R_1966_12fc2098 );
buf ( n6469 , R_a1b_123c17d8 );
buf ( n6470 , R_842_13bf4738 );
buf ( n6471 , R_e61_13cd0958 );
buf ( n6472 , R_103a_13ccdbb8 );
buf ( n6473 , R_1480_117f1e98 );
buf ( n6474 , R_1659_13c1fcb8 );
buf ( n6475 , R_820_17013088 );
buf ( n6476 , R_a3d_11c6bc78 );
buf ( n6477 , R_e3f_123c0e78 );
buf ( n6478 , R_105c_13dd87d8 );
buf ( n6479 , R_145e_13d5a3d8 );
buf ( n6480 , R_167b_14a19878 );
buf ( n6481 , R_ebb_13def998 );
buf ( n6482 , R_89c_1486e898 );
buf ( n6483 , R_9c1_13cd04f8 );
buf ( n6484 , R_fe0_15fee7a8 );
buf ( n6485 , R_14da_13b95818 );
buf ( n6486 , R_15ff_117f1538 );
buf ( n6487 , R_8d0_13ccd078 );
buf ( n6488 , R_98d_13cceab8 );
buf ( n6489 , R_eef_15ff2308 );
buf ( n6490 , R_fac_13df65b8 );
buf ( n6491 , R_150e_13bed398 );
buf ( n6492 , R_15cb_1580a558 );
buf ( n6493 , R_663_13c24218 );
buf ( n6494 , R_c82_11633bb8 );
buf ( n6495 , R_bfa_117f1d58 );
buf ( n6496 , R_5db_13c0d798 );
buf ( n6497 , R_1219_156b0f98 );
buf ( n6498 , R_12a1_15811e98 );
buf ( n6499 , R_1838_123c2098 );
buf ( n6500 , R_18c0_13ddb258 );
buf ( n6501 , R_bbb_13c08dd8 );
buf ( n6502 , R_6a2_14870cd8 );
buf ( n6503 , R_59c_1700ffc8 );
buf ( n6504 , R_cc1_13d5b0f8 );
buf ( n6505 , R_11da_14b1dcf8 );
buf ( n6506 , R_12e0_14b29c38 );
buf ( n6507 , R_17f9_13ddb438 );
buf ( n6508 , R_18ff_1162d538 );
buf ( n6509 , R_ecc_123bde58 );
buf ( n6510 , R_9b0_1587f458 );
buf ( n6511 , R_8ad_10082e38 );
buf ( n6512 , R_fcf_14a0e798 );
buf ( n6513 , R_14eb_140ad258 );
buf ( n6514 , R_15ee_117f3158 );
buf ( n6515 , R_d13_13c25e38 );
buf ( n6516 , R_6f4_156b4918 );
buf ( n6517 , R_b69_11c6e8d8 );
buf ( n6518 , R_1188_13cd35b8 );
buf ( n6519 , R_1332_11637d58 );
buf ( n6520 , R_17a7_117f6a38 );
buf ( n6521 , R_1951_156b6b78 );
buf ( n6522 , R_acf_13d503d8 );
buf ( n6523 , R_dad_13cd3838 );
buf ( n6524 , R_78e_13b929d8 );
buf ( n6525 , R_10ee_1587c438 );
buf ( n6526 , R_13cc_1587b3f8 );
buf ( n6527 , R_170d_12fbf9d8 );
buf ( n6528 , R_19eb_15ff53c8 );
buf ( n6529 , R_8c8_12fbe038 );
buf ( n6530 , R_ee7_13c03dd8 );
buf ( n6531 , R_995_13d50518 );
buf ( n6532 , R_fb4_156b0e58 );
buf ( n6533 , R_1506_156b9e18 );
buf ( n6534 , R_15d3_123b5ed8 );
buf ( n6535 , R_b9b_13dfa118 );
buf ( n6536 , R_6c2_14b1d618 );
buf ( n6537 , R_57c_13d464b8 );
buf ( n6538 , R_ce1_13d27358 );
buf ( n6539 , R_11ba_13cda458 );
buf ( n6540 , R_1300_13dec478 );
buf ( n6541 , R_17d9_156af918 );
buf ( n6542 , R_191f_14a0d578 );
buf ( n6543 , R_7e4_117f6c18 );
buf ( n6544 , R_e03_13b8c718 );
buf ( n6545 , R_a79_13d52db8 );
buf ( n6546 , R_1098_13cd2438 );
buf ( n6547 , R_1422_13cd7f78 );
buf ( n6548 , R_16b7_14b28518 );
buf ( n6549 , R_1a41_150e4d78 );
buf ( n6550 , R_ae5_17012048 );
buf ( n6551 , R_d97_1162ab58 );
buf ( n6552 , R_778_13d52098 );
buf ( n6553 , R_1104_13dd7a18 );
buf ( n6554 , R_13b6_14a17118 );
buf ( n6555 , R_1723_13d50018 );
buf ( n6556 , R_19d5_117edc58 );
buf ( n6557 , R_d53_13c0ae58 );
buf ( n6558 , R_b29_13b95c78 );
buf ( n6559 , R_734_14a0f558 );
buf ( n6560 , R_1148_117f6218 );
buf ( n6561 , R_1372_11c6cd58 );
buf ( n6562 , R_1767_11c691f8 );
buf ( n6563 , R_1991_13cd58b8 );
buf ( n6564 , R_f2c_15814d78 );
buf ( n6565 , R_90d_158848b8 );
buf ( n6566 , R_950_140b3798 );
buf ( n6567 , R_f6f_14a1a318 );
buf ( n6568 , R_154b_11632218 );
buf ( n6569 , R_158e_14a0b1d8 );
buf ( n6570 , R_ec6_13d37b98 );
buf ( n6571 , R_8a7_1580e6f8 );
buf ( n6572 , R_9b6_14a0cc18 );
buf ( n6573 , R_fd5_1580cc18 );
buf ( n6574 , R_14e5_13b8fd78 );
buf ( n6575 , R_15f4_170165a8 );
buf ( n6576 , R_7c0_100854f8 );
buf ( n6577 , R_ddf_13b92898 );
buf ( n6578 , R_a9d_1162c318 );
buf ( n6579 , R_10bc_140b7d98 );
buf ( n6580 , R_13fe_13cd60d8 );
buf ( n6581 , R_16db_156aaf58 );
buf ( n6582 , R_1a1d_13cd9ff8 );
buf ( n6583 , R_7f5_13b9a1d8 );
buf ( n6584 , R_e14_123bf078 );
buf ( n6585 , R_a68_150dbbd8 );
buf ( n6586 , R_1087_1587ad18 );
buf ( n6587 , R_1433_13dd7978 );
buf ( n6588 , R_16a6_13df8458 );
buf ( n6589 , R_1a52_11c70778 );
buf ( n6590 , R_646_156ad618 );
buf ( n6591 , R_c65_10086538 );
buf ( n6592 , R_c17_13ccb3b8 );
buf ( n6593 , R_5f8_1580f418 );
buf ( n6594 , R_1236_1587e558 );
buf ( n6595 , R_1284_14a1a458 );
buf ( n6596 , R_1855_10084a58 );
buf ( n6597 , R_18a3_1700b1a8 );
buf ( n6598 , R_69c_156b9058 );
buf ( n6599 , R_bc1_13bee298 );
buf ( n6600 , R_cbb_13ccbbd8 );
buf ( n6601 , R_5a2_15813658 );
buf ( n6602 , R_11e0_1587e878 );
buf ( n6603 , R_12da_14b29d78 );
buf ( n6604 , R_17ff_14a10b38 );
buf ( n6605 , R_18f9_14a16718 );
buf ( n6606 , R_adc_156ae6f8 );
buf ( n6607 , R_da0_13bf5db8 );
buf ( n6608 , R_781_13d42f98 );
buf ( n6609 , R_10fb_10085778 );
buf ( n6610 , R_13bf_123bf6b8 );
buf ( n6611 , R_171a_150deb58 );
buf ( n6612 , R_19de_117ef918 );
buf ( n6613 , R_9e7_13d54578 );
buf ( n6614 , R_e95_13d26ef8 );
buf ( n6615 , R_876_13d41698 );
buf ( n6616 , R_1006_13c08f18 );
buf ( n6617 , R_14b4_1700e268 );
buf ( n6618 , R_1625_13b96d58 );
buf ( n6619 , R_807_13cd8478 );
buf ( n6620 , R_e26_1700df48 );
buf ( n6621 , R_a56_124c4ad8 );
buf ( n6622 , R_1075_15883b98 );
buf ( n6623 , R_1445_15880218 );
buf ( n6624 , R_1694_13d218b8 );
buf ( n6625 , R_1a64_13ccac38 );
buf ( n6626 , R_a28_13cd9918 );
buf ( n6627 , R_835_140b35b8 );
buf ( n6628 , R_e54_14a179d8 );
buf ( n6629 , R_1047_14b26df8 );
buf ( n6630 , R_1473_156b60d8 );
buf ( n6631 , R_1666_14a165d8 );
buf ( n6632 , R_b0e_14a15818 );
buf ( n6633 , R_d6e_14a0c998 );
buf ( n6634 , R_74f_13c24678 );
buf ( n6635 , R_112d_1162be18 );
buf ( n6636 , R_138d_13b92258 );
buf ( n6637 , R_174c_116339d8 );
buf ( n6638 , R_19ac_14b1b4f8 );
buf ( n6639 , R_bb5_13cd29d8 );
buf ( n6640 , R_6a8_1162e618 );
buf ( n6641 , R_596_13dd6398 );
buf ( n6642 , R_cc7_123b4b78 );
buf ( n6643 , R_11d4_15ff30c8 );
buf ( n6644 , R_12e6_14a0ff58 );
buf ( n6645 , R_17f3_13ddb578 );
buf ( n6646 , R_1905_1486dfd8 );
buf ( n6647 , R_baa_14a15278 );
buf ( n6648 , R_6b3_17011288 );
buf ( n6649 , R_58b_140b1c18 );
buf ( n6650 , R_cd2_13d24dd8 );
buf ( n6651 , R_11c9_14b25278 );
buf ( n6652 , R_12f1_1587da18 );
buf ( n6653 , R_17e8_1587c078 );
buf ( n6654 , R_1910_12fc0978 );
buf ( n6655 , R_66e_17014348 );
buf ( n6656 , R_c8d_123b7ff8 );
buf ( n6657 , R_bef_14a167b8 );
buf ( n6658 , R_5d0_13c1db98 );
buf ( n6659 , R_120e_13c0d518 );
buf ( n6660 , R_12ac_13ccaf58 );
buf ( n6661 , R_182d_140b0098 );
buf ( n6662 , R_18cb_123b9e98 );
buf ( n6663 , R_8b3_13c0d298 );
buf ( n6664 , R_ed2_1580c538 );
buf ( n6665 , R_9aa_124c51b8 );
buf ( n6666 , R_fc9_13b8d118 );
buf ( n6667 , R_14f1_150e8978 );
buf ( n6668 , R_15e8_15884db8 );
buf ( n6669 , R_8e2_13bf6858 );
buf ( n6670 , R_97b_150e7a78 );
buf ( n6671 , R_f01_14a13e78 );
buf ( n6672 , R_f9a_116364f8 );
buf ( n6673 , R_1520_1162d678 );
buf ( n6674 , R_15b9_13d21a98 );
buf ( n6675 , R_7fa_123bbbf8 );
buf ( n6676 , R_e19_13d59ed8 );
buf ( n6677 , R_a63_14a16678 );
buf ( n6678 , R_1082_13c09d78 );
buf ( n6679 , R_1438_13bf2398 );
buf ( n6680 , R_16a1_14a16cb8 );
buf ( n6681 , R_1a57_13c28a98 );
buf ( n6682 , R_81d_1580d078 );
buf ( n6683 , R_a40_123bcd78 );
buf ( n6684 , R_e3c_117f2c58 );
buf ( n6685 , R_105f_13de2558 );
buf ( n6686 , R_145b_11633e38 );
buf ( n6687 , R_167e_1486d858 );
buf ( n6688 , R_7f0_13b90458 );
buf ( n6689 , R_e0f_140ab138 );
buf ( n6690 , R_a6d_117ee838 );
buf ( n6691 , R_108c_13bf90f8 );
buf ( n6692 , R_142e_11632538 );
buf ( n6693 , R_16ab_140b8d38 );
buf ( n6694 , R_1a4d_11c70bd8 );
buf ( n6695 , R_7d6_14b1e3d8 );
buf ( n6696 , R_df5_1580eab8 );
buf ( n6697 , R_a87_14a10138 );
buf ( n6698 , R_10a6_117efa58 );
buf ( n6699 , R_1414_1162b9b8 );
buf ( n6700 , R_16c5_14a10db8 );
buf ( n6701 , R_1a33_1486ebb8 );
buf ( n6702 , R_f0c_140b21b8 );
buf ( n6703 , R_8ed_11636d18 );
buf ( n6704 , R_970_13c0f818 );
buf ( n6705 , R_f8f_11632fd8 );
buf ( n6706 , R_152b_13beb778 );
buf ( n6707 , R_15ae_123b2eb8 );
buf ( n6708 , R_e6b_13b8ded8 );
buf ( n6709 , R_a11_158133d8 );
buf ( n6710 , R_84c_13bef918 );
buf ( n6711 , R_1030_140b72f8 );
buf ( n6712 , R_148a_140b0598 );
buf ( n6713 , R_164f_13d52778 );
buf ( n6714 , R_afa_123c0c98 );
buf ( n6715 , R_d82_13cd1858 );
buf ( n6716 , R_763_1580e298 );
buf ( n6717 , R_1119_1587c118 );
buf ( n6718 , R_13a1_158898b8 );
buf ( n6719 , R_1738_11c6f878 );
buf ( n6720 , R_19c0_1007ded8 );
buf ( n6721 , R_e7d_15811538 );
buf ( n6722 , R_9ff_13d245b8 );
buf ( n6723 , R_85e_13cd3018 );
buf ( n6724 , R_101e_13d5d8f8 );
buf ( n6725 , R_149c_13d5a978 );
buf ( n6726 , R_163d_13ccd438 );
buf ( n6727 , R_b8d_156aae18 );
buf ( n6728 , R_6d0_1162bb98 );
buf ( n6729 , R_56e_10086e98 );
buf ( n6730 , R_cef_14870eb8 );
buf ( n6731 , R_11ac_13c24498 );
buf ( n6732 , R_130e_14a17758 );
buf ( n6733 , R_17cb_14a0e478 );
buf ( n6734 , R_192d_123becb8 );
buf ( n6735 , R_d32_13d20558 );
buf ( n6736 , R_713_15882978 );
buf ( n6737 , R_b4a_13d22cb8 );
buf ( n6738 , R_1169_123b7c38 );
buf ( n6739 , R_1351_14a14558 );
buf ( n6740 , R_1788_13ccae18 );
buf ( n6741 , R_1970_124c43f8 );
buf ( n6742 , R_7cd_13d58df8 );
buf ( n6743 , R_dec_156ae518 );
buf ( n6744 , R_a90_13dd8058 );
buf ( n6745 , R_10af_117f0818 );
buf ( n6746 , R_140b_1580d1b8 );
buf ( n6747 , R_16ce_117ebe58 );
buf ( n6748 , R_1a2a_15810e58 );
buf ( n6749 , R_e72_13c1e8b8 );
buf ( n6750 , R_a0a_13d54438 );
buf ( n6751 , R_853_123bd778 );
buf ( n6752 , R_1029_13cd2898 );
buf ( n6753 , R_1491_117f33d8 );
buf ( n6754 , R_1648_15ff12c8 );
buf ( n6755 , R_80f_13d449d8 );
buf ( n6756 , R_a4e_13b8e798 );
buf ( n6757 , R_e2e_13dd57b8 );
buf ( n6758 , R_106d_13b8b598 );
buf ( n6759 , R_144d_13cd65d8 );
buf ( n6760 , R_168c_15ff1c28 );
buf ( R_187c_13cca558 , n17500 );
buf ( R_125d_156aaaf8 , n18225 );
buf ( R_c3e_13d2c178 , C0 );
buf ( R_61f_117eb278 , n18227 );
buf ( R_187d_117f5b38 , n19650 );
buf ( R_125e_13b8fe18 , C0 );
buf ( R_c3f_123b4358 , n19652 );
buf ( R_187b_13ccb278 , n19654 );
buf ( R_620_13dfb518 , n19656 );
buf ( R_125c_15816b78 , n19657 );
buf ( R_c3d_13c22918 , n20662 );
buf ( R_61e_14a0c538 , C0 );
buf ( R_5e7_10080958 , n20664 );
buf ( R_c06_170189e8 , C0 );
buf ( R_18b4_1162f978 , n20666 );
buf ( R_1225_13c08298 , n21799 );
buf ( R_1844_117ef378 , n21801 );
buf ( R_1295_123bcf58 , n22004 );
buf ( R_c76_15ff42e8 , C0 );
buf ( R_657_13bf5c78 , n22006 );
buf ( R_187e_140ac0d8 , C0 );
buf ( R_125f_13c0f638 , n22008 );
buf ( R_c40_1580a9b8 , n22010 );
buf ( R_621_11c70318 , n22304 );
buf ( R_187a_13ddd2d8 , C0 );
buf ( R_61d_123b84f8 , n22341 );
buf ( R_125b_1162bf58 , n22342 );
buf ( R_c3c_15ff9928 , n22344 );
buf ( R_12be_13ccf378 , C0 );
buf ( R_5be_11c6a738 , C0 );
buf ( R_bdd_17016508 , n22401 );
buf ( R_c9f_11636598 , n22403 );
buf ( R_11fc_13ddf7b8 , n22405 );
buf ( R_680_10085638 , n22407 );
buf ( R_181b_13d430d8 , n22409 );
buf ( R_18dd_13c062b8 , n22478 );
buf ( R_180c_156b4eb8 , n22480 );
buf ( R_12cd_13d535d8 , n22638 );
buf ( R_5af_1700c3c8 , n22652 );
buf ( R_cae_14a14ff8 , C0 );
buf ( R_bce_15ff4608 , C0 );
buf ( R_68f_13befcd8 , n22654 );
buf ( R_18ec_13d204b8 , n22656 );
buf ( R_11ed_116361d8 , n22713 );
buf ( R_187f_15811038 , n22715 );
buf ( R_1260_13d3b6f8 , n22717 );
buf ( R_c41_14a0bef8 , n22737 );
buf ( R_622_123b3bd8 , C0 );
buf ( R_61c_13d56378 , n22739 );
buf ( R_c3b_150e7c58 , n22741 );
buf ( R_1879_15ff5c88 , n22787 );
buf ( R_125a_13bf58b8 , C0 );
buf ( R_f82_13c1cd38 , C0 );
buf ( R_963_13c209d8 , n22789 );
buf ( R_8fa_117ec678 , C0 );
buf ( R_f19_15ff0648 , n379402 );
buf ( R_1538_13d29bf8 , n379404 );
buf ( R_15a1_150e22f8 , n379800 );
buf ( R_158f_13cd9058 , n379801 );
buf ( R_f70_17015608 , n379803 );
buf ( R_951_156b2578 , n379843 );
buf ( R_90c_13c0e0f8 , n379845 );
buf ( R_f2b_140b8838 , n379846 );
buf ( R_154a_1587f278 , C0 );
buf ( R_1880_13c22738 , n379848 );
buf ( R_1261_13ccc0d8 , n379892 );
buf ( R_c42_117eb818 , C0 );
buf ( R_623_140b3158 , n379894 );
buf ( R_61b_11c70458 , n379896 );
buf ( R_c3a_13b96218 , C0 );
buf ( R_1259_13d23578 , n379941 );
buf ( R_1878_1162da38 , n379942 );
buf ( R_ce6_14875d78 , C0 );
buf ( R_1924_13d1df38 , n379943 );
buf ( R_11b5_13d56f58 , n380201 );
buf ( R_577_1162c818 , n380202 );
buf ( R_6c7_10082438 , n380204 );
buf ( R_17d4_13cda278 , n380205 );
buf ( R_1305_10081fd8 , n380795 );
buf ( R_b96_15812b18 , C0 );
buf ( R_1881_156b0638 , n380863 );
buf ( R_1262_12fc1698 , C0 );
buf ( R_c43_140b0138 , n380864 );
buf ( R_624_13d421d8 , n380866 );
buf ( R_61a_14b2a318 , C0 );
buf ( R_c39_117eaeb8 , n380900 );
buf ( R_1258_117e8618 , n380901 );
buf ( R_1877_1162cdb8 , n380902 );
buf ( R_119b_15ffa3c8 , n380904 );
buf ( R_55d_13b8e5b8 , n380905 );
buf ( R_131f_158106d8 , n380907 );
buf ( R_6e1_13c0fb38 , n380939 );
buf ( R_17ba_15fed6c8 , C0 );
buf ( R_b7c_13b96e98 , n380941 );
buf ( R_193e_123b6018 , C0 );
buf ( R_d00_117ec358 , n380943 );
buf ( R_1323_13d5b878 , n380944 );
buf ( R_6e5_15ff5328 , n381001 );
buf ( R_559_13c024d8 , n381002 );
buf ( R_1197_13bf4918 , n381003 );
buf ( R_1942_11c6dd98 , C0 );
buf ( R_d04_14a16df8 , n381005 );
buf ( R_17b6_13dec158 , C0 );
buf ( R_b78_13c10c18 , n381007 );
buf ( R_13ca_13d2c718 , C0 );
buf ( R_19e9_13bf62b8 , n381020 );
buf ( R_170f_150defb8 , n381022 );
buf ( R_10f0_140b1ad8 , n381023 );
buf ( R_ad1_11c6ac38 , n381080 );
buf ( R_78c_13d5d3f8 , n381082 );
buf ( R_dab_140b3dd8 , n381083 );
buf ( R_883_13b936f8 , n381084 );
buf ( R_ff9_11631958 , n381489 );
buf ( R_ea2_150dd758 , C0 );
buf ( R_9da_13cd8018 , C0 );
buf ( R_1618_117f3658 , n381491 );
buf ( R_14c1_123ba4d8 , n381565 );
buf ( R_b5e_14a0f918 , C0 );
buf ( R_179c_123bb018 , n381567 );
buf ( R_133d_13cd4e18 , n381626 );
buf ( R_6ff_14a0a918 , n381627 );
buf ( R_195c_150ddf78 , n381628 );
buf ( R_117d_123b8c78 , n381706 );
buf ( R_d1e_124c2cd8 , C0 );
buf ( R_5f7_12fbf758 , n381708 );
buf ( R_c16_13df9858 , C0 );
buf ( R_1235_15880cb8 , n381836 );
buf ( R_1854_1580fd78 , n381837 );
buf ( R_18a4_13bf2d98 , n381838 );
buf ( R_1285_100890f8 , n381871 );
buf ( R_c66_13bed2f8 , C0 );
buf ( R_647_13d51af8 , n381873 );
buf ( R_1882_13d1fbf8 , C0 );
buf ( R_1263_123be498 , n381874 );
buf ( R_c44_13c229b8 , n381875 );
buf ( R_625_13c1e638 , n381885 );
buf ( R_619_156b6718 , n381932 );
buf ( R_c38_117efd78 , n381933 );
buf ( R_1257_14a0f0f8 , n381934 );
buf ( R_1876_15ffcb28 , C0 );
buf ( R_985_1587c4d8 , n382047 );
buf ( R_1516_12fc1eb8 , C0 );
buf ( R_15c3_13c02078 , n382048 );
buf ( R_8d8_13d22fd8 , n382050 );
buf ( R_fa4_13d1e898 , n382051 );
buf ( R_ef7_1162bd78 , n382053 );
buf ( R_1663_124c2698 , n382054 );
buf ( R_838_1580b8b8 , n382055 );
buf ( R_a25_13bf4ff8 , n382064 );
buf ( R_1476_1486bd78 , C0 );
buf ( R_1044_13d57818 , n382066 );
buf ( R_e57_13b8f738 , n382068 );
buf ( R_15fa_13c0bb78 , C0 );
buf ( R_ec0_13c1bf78 , n382070 );
buf ( R_fdb_15ff7308 , n382072 );
buf ( R_14df_14a0cdf8 , n382074 );
buf ( R_9bc_15812758 , n382075 );
buf ( R_8a1_13d21818 , n382535 );
buf ( R_1883_13d41058 , n382536 );
buf ( R_1264_13c02758 , n382538 );
buf ( R_c45_13d24c98 , n382555 );
buf ( R_626_123b86d8 , C0 );
buf ( R_618_1587ea58 , n382556 );
buf ( R_c37_13c0bfd8 , n382557 );
buf ( R_1256_13d54258 , C0 );
buf ( R_1875_158179d8 , n382623 );
buf ( R_1145_13b98658 , n382892 );
buf ( R_737_116313b8 , n382893 );
buf ( R_b26_1486a518 , C0 );
buf ( R_d56_117e9d38 , C0 );
buf ( R_1764_13ccf7d8 , n382894 );
buf ( R_1375_13c275f8 , n382972 );
buf ( R_1994_123bac58 , n382973 );
buf ( R_143d_13bf2258 , n383007 );
buf ( R_a5e_1587ed78 , C0 );
buf ( R_e1e_13c1bbb8 , C0 );
buf ( R_107d_15888418 , n383173 );
buf ( R_7ff_13cd45f8 , n383175 );
buf ( R_169c_15885fd8 , n383176 );
buf ( R_1a5c_13de04d8 , n383177 );
buf ( R_1a48_13c1ff38 , n383178 );
buf ( R_a72_1486d358 , C0 );
buf ( R_1429_13d23438 , n383197 );
buf ( R_1091_14a11d58 , n383344 );
buf ( R_e0a_13bfa3b8 , C0 );
buf ( R_16b0_140aae18 , n383346 );
buf ( R_7eb_123b8278 , n383347 );
buf ( R_12c6_13cd49b8 , C0 );
buf ( R_5b6_117f1f38 , C0 );
buf ( R_ca7_140b4418 , n383348 );
buf ( R_bd5_13d51698 , n383399 );
buf ( R_688_13b99af8 , n383400 );
buf ( R_11f4_13d1e6b8 , n383401 );
buf ( R_18e5_13d45658 , n383497 );
buf ( R_1813_13d29c98 , n383499 );
buf ( R_16d9_14a17cf8 , n383611 );
buf ( R_1a1f_11c70958 , n383612 );
buf ( R_1400_14b29b98 , n383614 );
buf ( R_de1_13cd0638 , n383922 );
buf ( R_7c2_15ffa508 , C0 );
buf ( R_a9b_100865d8 , n383923 );
buf ( R_10ba_15881938 , C0 );
buf ( R_1805_14b271b8 , n384048 );
buf ( R_5a8_123b8318 , n384053 );
buf ( R_cb5_170107e8 , n384198 );
buf ( R_bc7_13c2a758 , n384200 );
buf ( R_696_10082ed8 , C0 );
buf ( R_18f3_15ffc628 , n384201 );
buf ( R_11e6_14b222f8 , C0 );
buf ( R_12d4_11634d38 , n384202 );
buf ( R_119f_156b4738 , n384204 );
buf ( R_561_1162a658 , n384205 );
buf ( R_6dd_117f36f8 , n384215 );
buf ( R_131b_15ff76c8 , n384216 );
buf ( R_17be_15816538 , C0 );
buf ( R_b80_13cd8338 , n384217 );
buf ( R_cfc_1700d2c8 , n384219 );
buf ( R_193a_15885718 , C0 );
buf ( R_5da_13df70f8 , C0 );
buf ( R_18c1_11c6f738 , n384660 );
buf ( R_bf9_13d28ed8 , n384696 );
buf ( R_12a2_13bf2578 , C0 );
buf ( R_1218_13d28078 , n384697 );
buf ( R_c83_13d59f78 , n384698 );
buf ( R_1837_13deb9d8 , n384699 );
buf ( R_664_123b47b8 , n384701 );
buf ( R_e39_156b3518 , n384764 );
buf ( R_a43_14b1feb8 , n384765 );
buf ( R_81a_13cceb58 , C0 );
buf ( R_1062_117eedd8 , C0 );
buf ( R_1458_13df07f8 , n384766 );
buf ( R_1681_140b99b8 , n384940 );
buf ( R_1327_124c2b98 , n384941 );
buf ( R_6e9_156b3158 , n384993 );
buf ( R_555_13d59b18 , n384994 );
buf ( R_1193_13b97438 , n384995 );
buf ( R_1946_14a16858 , C0 );
buf ( R_d08_13d59938 , n384997 );
buf ( R_b74_123c0478 , n384998 );
buf ( R_17b2_13cd6498 , C0 );
buf ( R_113a_117eb458 , C0 );
buf ( R_742_14a129d8 , C0 );
buf ( R_b1b_11629758 , n384999 );
buf ( R_d61_11633618 , n385029 );
buf ( R_1380_15887338 , n385030 );
buf ( R_1759_14874518 , n385047 );
buf ( R_199f_13d3c9b8 , n385048 );
buf ( R_1884_13cd1c18 , n385049 );
buf ( R_1265_156b0818 , n385080 );
buf ( R_c46_1580b598 , C0 );
buf ( R_627_117efb98 , n385081 );
buf ( R_617_158807b8 , n385082 );
buf ( R_c36_156b63f8 , C0 );
buf ( R_1255_1580dbb8 , n385111 );
buf ( R_1874_13df9c18 , n385113 );
buf ( R_87a_13c286d8 , C0 );
buf ( R_1002_14a17938 , C0 );
buf ( R_e99_123ba258 , n385183 );
buf ( R_9e3_170110a8 , n385184 );
buf ( R_1621_117eacd8 , n385192 );
buf ( R_14b8_123b31d8 , n385193 );
buf ( R_edf_117f5bd8 , n385194 );
buf ( R_14fe_13d55518 , C0 );
buf ( R_15db_117f7258 , n385196 );
buf ( R_fbc_13beb9f8 , n385198 );
buf ( R_8c0_11631ef8 , n385199 );
buf ( R_99d_13cd4d78 , n385226 );
buf ( R_845_15888918 , n386562 );
buf ( R_1656_117f4af8 , C0 );
buf ( R_1483_13d53d58 , n386564 );
buf ( R_a18_12fbdef8 , n386565 );
buf ( R_e64_14875058 , n386566 );
buf ( R_1037_15815098 , n386567 );
buf ( R_d8e_11630878 , C0 );
buf ( R_172c_13d39d58 , n386568 );
buf ( R_13ad_14a12618 , n386632 );
buf ( R_19cc_13cda1d8 , n386633 );
buf ( R_110d_13dd5cb8 , n386684 );
buf ( R_aee_117e9478 , C0 );
buf ( R_76f_117f4378 , n386685 );
buf ( R_ccd_13b8c8f8 , n386743 );
buf ( R_590_13dd64d8 , n386744 );
buf ( R_17ed_156b36f8 , n386755 );
buf ( R_190b_14872038 , n386756 );
buf ( R_6ae_156ab958 , C0 );
buf ( R_baf_1700cd28 , n386757 );
buf ( R_12ec_124c3778 , n386758 );
buf ( R_11ce_11c6cad8 , C0 );
buf ( R_17a3_150e7398 , n386759 );
buf ( R_1336_148754b8 , C0 );
buf ( R_6f8_13c1c018 , n386761 );
buf ( R_1184_150e6498 , n386763 );
buf ( R_1955_14b235b8 , n30863 );
buf ( R_d17_14b27398 , n30864 );
buf ( R_b65_13dde318 , n387114 );
buf ( R_1885_1486cdb8 , n387158 );
buf ( R_1266_14a12438 , C0 );
buf ( R_c47_100803b8 , n387160 );
buf ( R_628_117eb098 , n387161 );
buf ( R_616_170152e8 , C0 );
buf ( R_c35_123b88b8 , n30990 );
buf ( R_1254_150e59f8 , n30991 );
buf ( R_1873_12fc2278 , n30993 );
buf ( R_74a_1008cb18 , C0 );
buf ( R_1132_15880e98 , C0 );
buf ( R_d69_14b23158 , n31029 );
buf ( R_b13_140b3d38 , n31031 );
buf ( R_1388_140aaf58 , n31032 );
buf ( R_19a7_140b9b98 , n31034 );
buf ( R_1751_1007feb8 , n31048 );
buf ( R_b57_13ccd6b8 , n31049 );
buf ( R_1344_117f3018 , n31050 );
buf ( R_1795_1008b678 , n31136 );
buf ( R_706_1580bd18 , C0 );
buf ( R_1963_13d1f478 , n31137 );
buf ( R_1176_17015b08 , C0 );
buf ( R_d25_15882298 , n31189 );
buf ( R_1590_150e4b98 , n31190 );
buf ( R_f71_124c4998 , n31718 );
buf ( R_952_14b26e98 , C0 );
buf ( R_90b_13d41af8 , n31720 );
buf ( R_f2a_1162a158 , C0 );
buf ( R_1549_1587ff98 , n31797 );
buf ( R_5c6_15816218 , C0 );
buf ( R_12b6_1587db58 , C0 );
buf ( R_be5_140b5818 , n31827 );
buf ( R_c97_156b09f8 , n31828 );
buf ( R_1204_13c23b38 , n31829 );
buf ( R_678_15884ef8 , n31830 );
buf ( R_1823_13d53df8 , n31831 );
buf ( R_18d5_11636098 , n31977 );
buf ( R_ed8_117e9c98 , n31978 );
buf ( R_15e2_14a140f8 , C0 );
buf ( R_14f7_13b965d8 , n31980 );
buf ( R_fc3_14b27e38 , n31981 );
buf ( R_8b9_14875e18 , n32058 );
buf ( R_9a4_117ee018 , n32059 );
buf ( R_1a04_13c22b98 , n32060 );
buf ( R_13e5_13de07f8 , n32092 );
buf ( R_16f4_123b9fd8 , n32093 );
buf ( R_dc6_14873f78 , C0 );
buf ( R_10d5_13b94a58 , n32107 );
buf ( R_7a7_116355f8 , n32108 );
buf ( R_ab6_15814e18 , C0 );
buf ( R_1886_11638c58 , C0 );
buf ( R_1267_14b23f18 , n32109 );
buf ( R_c48_13bf5e58 , n32110 );
buf ( R_629_150e7e38 , n32120 );
buf ( R_615_13c1d7d8 , n32155 );
buf ( R_c34_15ff1228 , n32156 );
buf ( R_1253_13d222b8 , n32157 );
buf ( R_1872_13ccb4f8 , C0 );
buf ( R_16f6_116389d8 , C0 );
buf ( R_10d7_156b5778 , n32158 );
buf ( R_ab8_156ac8f8 , n32159 );
buf ( R_1a02_13cd8298 , C0 );
buf ( R_13e3_14a0a7d8 , n32161 );
buf ( R_7a5_13d456f8 , n32193 );
buf ( R_dc4_11634b58 , n32194 );
buf ( R_b4d_1700f208 , n32233 );
buf ( R_710_156ac718 , n32234 );
buf ( R_178b_1580ca38 , n32235 );
buf ( R_196d_117eb8b8 , n32253 );
buf ( R_d2f_13dedf58 , n32254 );
buf ( R_116c_140b8338 , n32256 );
buf ( R_134e_13d282f8 , C0 );
buf ( R_1a06_1486e1b8 , C0 );
buf ( R_13e7_116377b8 , n32257 );
buf ( R_dc8_1162b058 , n32258 );
buf ( R_7a9_123bd458 , n32269 );
buf ( R_16f2_158857b8 , C0 );
buf ( R_ab4_12fbed58 , n32270 );
buf ( R_10d3_158899f8 , n32272 );
buf ( R_85a_156b1a38 , C0 );
buf ( R_1498_15811c18 , n32273 );
buf ( R_1641_150db8b8 , n32360 );
buf ( R_a03_123bd818 , n32361 );
buf ( R_e79_13cd8658 , n32373 );
buf ( R_1022_11c6cf38 , C0 );
buf ( R_150d_14b21678 , n32393 );
buf ( R_15cc_14a0ba98 , n32394 );
buf ( R_8cf_13ded9b8 , n32395 );
buf ( R_fad_140ac038 , n32413 );
buf ( R_eee_11632e98 , C0 );
buf ( R_98e_12fbecb8 , C0 );
buf ( R_13bd_13df6c98 , n32426 );
buf ( R_19dc_156b6858 , n32427 );
buf ( R_171c_117ecb78 , n32428 );
buf ( R_10fd_117eef18 , n32449 );
buf ( R_ade_13dd7658 , C0 );
buf ( R_77f_117f4558 , n32450 );
buf ( R_d9e_13ddc3d8 , C0 );
buf ( R_16f8_14a0e018 , n32451 );
buf ( R_10d9_123b9538 , n32469 );
buf ( R_aba_13c29678 , C0 );
buf ( R_7a3_13ccb138 , n32470 );
buf ( R_dc2_158108b8 , C0 );
buf ( R_13e1_156b8478 , n32484 );
buf ( R_1a00_123b7f58 , n32485 );
buf ( R_971_13df5618 , n32497 );
buf ( R_8ec_123bbd38 , n32498 );
buf ( R_15af_14866eb8 , n32499 );
buf ( R_f0b_13cd72f8 , n32500 );
buf ( R_f90_15812438 , n32501 );
buf ( R_152a_13df8818 , C0 );
buf ( R_c15_15fee528 , n32531 );
buf ( R_1234_15ff9e28 , n32532 );
buf ( R_1853_13dd8738 , n32533 );
buf ( R_18a5_170177c8 , n32591 );
buf ( R_1286_124c4858 , C0 );
buf ( R_c67_13ccba98 , n32592 );
buf ( R_648_15814058 , n32593 );
buf ( R_5f6_13cce018 , C0 );
buf ( R_c05_14866d78 , n32625 );
buf ( R_18b5_10087cf8 , n32671 );
buf ( R_1224_13ccff58 , n32673 );
buf ( R_1296_13dda7b8 , C0 );
buf ( R_1843_1580a878 , n32674 );
buf ( R_c77_13d523b8 , n32675 );
buf ( R_658_140ae1f8 , n32677 );
buf ( R_5e6_13d46698 , C0 );
buf ( R_1a08_14b1b958 , n32678 );
buf ( R_13e9_13d22358 , n32705 );
buf ( R_dca_14b297d8 , C0 );
buf ( R_7ab_15887ab8 , n32706 );
buf ( R_ab2_13df75f8 , C0 );
buf ( R_10d1_13d55d38 , n32716 );
buf ( R_16f0_14b1e978 , n32717 );
buf ( R_d87_123bae38 , n32718 );
buf ( R_1733_15ff79e8 , n32719 );
buf ( R_13a6_156b1718 , C0 );
buf ( R_1114_13d46ff8 , n32720 );
buf ( R_19c5_13bf6ad8 , n32728 );
buf ( R_af5_13c1b6b8 , n32832 );
buf ( R_768_158896d8 , n32833 );
buf ( R_964_123c1f58 , n32834 );
buf ( R_8f9_117ee658 , n32979 );
buf ( R_f18_14a19d78 , n32980 );
buf ( R_1537_117e9b58 , n32982 );
buf ( R_15a2_13ccce98 , C0 );
buf ( R_f83_14a0e978 , n32983 );
buf ( R_1887_17018da8 , n32984 );
buf ( R_1268_13d38278 , n32985 );
buf ( R_c49_123b36d8 , n33005 );
buf ( R_62a_13d42278 , C0 );
buf ( R_614_13c2a258 , n33006 );
buf ( R_c33_150e7bb8 , n33007 );
buf ( R_1252_116378f8 , C0 );
buf ( R_1871_13defad8 , n33076 );
buf ( R_11a3_13c1be38 , n33077 );
buf ( R_565_13ddbb18 , n33078 );
buf ( R_6d9_11636818 , n33090 );
buf ( R_1317_1580c5d8 , n33091 );
buf ( R_17c2_13c03518 , C0 );
buf ( R_b84_156b5278 , n33092 );
buf ( R_cf8_15881a78 , n33093 );
buf ( R_1936_13d2a558 , C0 );
buf ( R_13b4_156abb38 , n33094 );
buf ( R_19d3_13bf92d8 , n33095 );
buf ( R_1725_13cd9a58 , n33107 );
buf ( R_1106_14b1c718 , C0 );
buf ( R_ae7_13cd22f8 , n33108 );
buf ( R_776_14873bb8 , C0 );
buf ( R_d95_15815778 , n33140 );
buf ( R_feb_1486c818 , n33141 );
buf ( R_eb0_13d53498 , n33142 );
buf ( R_14cf_14b1bd18 , n33143 );
buf ( R_9cc_158172f8 , n33144 );
buf ( R_160a_17010ce8 , C0 );
buf ( R_891_13b8ab98 , n33163 );
buf ( R_132b_1007f7d8 , n33164 );
buf ( R_6ed_140b6538 , n33206 );
buf ( R_118f_14b1ee78 , n33207 );
buf ( R_194a_13d2ae18 , C0 );
buf ( R_d0c_13dee8b8 , n33208 );
buf ( R_b70_13d20f58 , n33209 );
buf ( R_17ae_13d29a18 , C0 );
buf ( R_1a3c_13b95278 , n33210 );
buf ( R_109d_10084878 , n33218 );
buf ( R_141d_13d441b8 , n33247 );
buf ( R_16bc_14a0bdb8 , n33248 );
buf ( R_dfe_15ff38e8 , C0 );
buf ( R_7df_1587d338 , n33249 );
buf ( R_a7e_14a0bb38 , C0 );
buf ( R_151f_12fbe998 , n33251 );
buf ( R_97c_13d528b8 , n33252 );
buf ( R_15ba_1008b0d8 , C0 );
buf ( R_8e1_15889818 , n33274 );
buf ( R_f00_17017ae8 , n33275 );
buf ( R_f9b_13b974d8 , n33276 );
buf ( R_16fa_14b299b8 , C0 );
buf ( R_10db_13cd6cb8 , n33277 );
buf ( R_abc_15882b58 , n33278 );
buf ( R_7a1_15ffcd08 , n33288 );
buf ( R_dc0_117f53b8 , n33289 );
buf ( R_13df_156b9238 , n33290 );
buf ( R_19fe_13c01fd8 , C0 );
buf ( R_5cf_124c4678 , n33291 );
buf ( R_12ad_13cca878 , n33321 );
buf ( R_bee_156ac498 , C0 );
buf ( R_c8e_156b6cb8 , C0 );
buf ( R_120d_123be218 , n33334 );
buf ( R_66f_13df8d18 , n33335 );
buf ( R_182c_13b90598 , n33336 );
buf ( R_18cc_170190c8 , n33337 );
buf ( R_1505_13d27858 , n33345 );
buf ( R_15d4_13d3a078 , n33346 );
buf ( R_fb5_13c265b8 , n33361 );
buf ( R_8c7_13ccf738 , n33362 );
buf ( R_996_13cd1498 , C0 );
buf ( R_ee6_156ae158 , C0 );
buf ( R_1a0a_140b9238 , C0 );
buf ( R_13eb_150e7438 , n33363 );
buf ( R_dcc_15815c78 , n33364 );
buf ( R_7ad_1008c078 , n33381 );
buf ( R_ab0_11629618 , n33383 );
buf ( R_10cf_1580df78 , n33384 );
buf ( R_16ee_123bf758 , C0 );
buf ( R_1660_13dd6258 , n33385 );
buf ( R_83b_117f03b8 , n33386 );
buf ( R_a22_156b92d8 , C0 );
buf ( R_1479_13ddc518 , n33448 );
buf ( R_1041_14a0db18 , n33483 );
buf ( R_e5a_11633118 , C0 );
buf ( R_1711_11c69d38 , n33595 );
buf ( R_10f2_1486ad38 , C0 );
buf ( R_ad3_13d5a5b8 , n33596 );
buf ( R_78a_13dfa2f8 , C0 );
buf ( R_da9_123bc9b8 , n33621 );
buf ( R_13c8_11628e98 , n33622 );
buf ( R_19e7_14a10098 , n33623 );
buf ( R_eb5_13cd9cd8 , n33659 );
buf ( R_fe6_13df1d38 , C0 );
buf ( R_14d4_13c27a58 , n33660 );
buf ( R_9c7_140af5f8 , n33661 );
buf ( R_896_123b6658 , C0 );
buf ( R_1605_156b1b78 , n34655 );
buf ( R_1888_1580c858 , n34656 );
buf ( R_1269_13b99c38 , n34685 );
buf ( R_c4a_14a0cb78 , C0 );
buf ( R_62b_1162a1f8 , n34686 );
buf ( R_613_124c47b8 , n34687 );
buf ( R_c32_14b23518 , C0 );
buf ( R_1251_13d3fed8 , n34698 );
buf ( R_1870_13b92bb8 , n34699 );
buf ( R_16cc_156ba318 , n34700 );
buf ( R_1a2c_156b08b8 , n34701 );
buf ( R_140d_11638258 , n34712 );
buf ( R_dee_13c0e058 , C0 );
buf ( R_7cf_123bbe78 , n34713 );
buf ( R_a8e_170160a8 , C0 );
buf ( R_10ad_10082618 , n34722 );
buf ( R_11b0_13b99f58 , n34723 );
buf ( R_572_140ab458 , n34724 );
buf ( R_6cc_117e8a78 , n34725 );
buf ( R_130a_13dda498 , C0 );
buf ( R_17cf_13d389f8 , n34726 );
buf ( R_b91_14b1f418 , n34808 );
buf ( R_ceb_13d56d78 , n34809 );
buf ( R_1929_13cd4af8 , n34851 );
buf ( R_f72_13c2a1b8 , C0 );
buf ( R_953_14b20a98 , n34852 );
buf ( R_90a_156ae658 , C0 );
buf ( R_f29_11630698 , n34883 );
buf ( R_1548_140ac538 , n34884 );
buf ( R_1591_13c25618 , n34891 );
buf ( R_16fc_156b9a58 , n34892 );
buf ( R_10dd_13d551f8 , n34914 );
buf ( R_abe_14a15958 , C0 );
buf ( R_79f_140af7d8 , n34915 );
buf ( R_dbe_13cd4c38 , C0 );
buf ( R_13dd_15884b38 , n34926 );
buf ( R_19fc_13b96fd8 , n34927 );
buf ( R_ff0_123b3b38 , n34928 );
buf ( R_eab_11634518 , n34929 );
buf ( R_9d1_13d4ed58 , n35125 );
buf ( R_14ca_11631e58 , C0 );
buf ( R_160f_170102e8 , n35126 );
buf ( R_88c_116319f8 , n35127 );
buf ( R_e36_13c05b38 , C0 );
buf ( R_a46_11637e98 , C0 );
buf ( R_817_116294d8 , n35128 );
buf ( R_1065_13c0b218 , n35143 );
buf ( R_1455_117ef238 , n35172 );
buf ( R_1684_13dd5ad8 , n35173 );
buf ( R_e2b_13d28578 , n35174 );
buf ( R_a51_11630ff8 , n35210 );
buf ( R_80c_13d2acd8 , n35211 );
buf ( R_1070_150e2d98 , n35212 );
buf ( R_1a69_11c6fe18 , n35218 );
buf ( R_168f_13d295b8 , n35219 );
buf ( R_144a_1580c678 , C0 );
buf ( R_1a0c_13ccacd8 , n35220 );
buf ( R_13ed_13cd4ff8 , n35231 );
buf ( R_dce_14871f98 , C0 );
buf ( R_7af_11633578 , n35232 );
buf ( R_aae_15814238 , C0 );
buf ( R_10cd_13d20878 , n35248 );
buf ( R_16ec_13df6a18 , n35249 );
buf ( R_1889_13bf9c38 , n35290 );
buf ( R_126a_15886a78 , C0 );
buf ( R_c4b_13cd76b8 , n35291 );
buf ( R_62c_10086038 , n35292 );
buf ( R_612_10088dd8 , C0 );
buf ( R_c31_13b90778 , n35323 );
buf ( R_1250_13d58c18 , n35324 );
buf ( R_186f_1162dcb8 , n35325 );
buf ( R_1a21_150e5598 , n35330 );
buf ( R_1402_140b1cb8 , C0 );
buf ( R_de3_140b0778 , n35331 );
buf ( R_7c4_13cd5138 , n35332 );
buf ( R_a99_13cd0a98 , n35465 );
buf ( R_10b8_13bea7d8 , n35466 );
buf ( R_16d7_15888a58 , n35467 );
buf ( R_b23_1587bc18 , n35468 );
buf ( R_d59_14868cb8 , n35503 );
buf ( R_1378_14b28158 , n35504 );
buf ( R_1761_11631f98 , n35521 );
buf ( R_1997_13d45158 , n35522 );
buf ( R_1142_117f06d8 , C0 );
buf ( R_73a_13de1158 , C0 );
buf ( R_1a35_1486d7b8 , n35528 );
buf ( R_16c3_13c01498 , n35529 );
buf ( R_1416_1162ee38 , C0 );
buf ( R_df7_117f35b8 , n35530 );
buf ( R_7d8_156abc78 , n35531 );
buf ( R_a85_17014168 , n35586 );
buf ( R_10a4_1486b0f8 , n35587 );
buf ( R_a59_14a1a1d8 , n35606 );
buf ( R_e23_13df5f78 , n35607 );
buf ( R_1078_1580f558 , n35608 );
buf ( R_804_156b6f38 , n35609 );
buf ( R_1697_13d59d98 , n35610 );
buf ( R_1a61_14a195f8 , n35612 );
buf ( R_1442_14a18c98 , C0 );
buf ( R_1096_13dd6f78 , C0 );
buf ( R_1424_13b906d8 , n35613 );
buf ( R_16b5_13c045f8 , n35621 );
buf ( R_e05_140ad938 , n35646 );
buf ( R_7e6_1486dd58 , C0 );
buf ( R_a77_100895f8 , n35647 );
buf ( R_1a43_170104c8 , n35648 );
buf ( R_15ef_15889318 , n35650 );
buf ( R_ecb_13df7198 , n35652 );
buf ( R_14ea_13cd2078 , C0 );
buf ( R_fd0_13cd59f8 , n35653 );
buf ( R_8ac_15889278 , n35654 );
buf ( R_9b1_1008a3b8 , n35662 );
buf ( R_cc2_14a11218 , C0 );
buf ( R_17f8_13c28d18 , n35663 );
buf ( R_59b_15812bb8 , n35668 );
buf ( R_1900_1486c318 , n35669 );
buf ( R_6a3_11c69658 , n35670 );
buf ( R_bba_13deb7f8 , C0 );
buf ( R_12e1_123bbf18 , n35689 );
buf ( R_11d9_14a18518 , n35727 );
buf ( R_1125_124c3e58 , n35782 );
buf ( R_d76_156b6218 , C0 );
buf ( R_b06_14b24af8 , C0 );
buf ( R_1395_13c0d978 , n35817 );
buf ( R_19b4_14a10598 , n35818 );
buf ( R_1744_11c6e3d8 , n35819 );
buf ( R_757_13d3ceb8 , n35820 );
buf ( R_16fe_123b51b8 , C0 );
buf ( R_10df_156b31f8 , n35821 );
buf ( R_ac0_123c19b8 , n35822 );
buf ( R_79d_13ddd698 , n35832 );
buf ( R_dbc_13d207d8 , n35833 );
buf ( R_13db_13d412d8 , n35834 );
buf ( R_19fa_140afeb8 , C0 );
buf ( R_188a_14a0dd98 , C0 );
buf ( R_126b_170193e8 , n35835 );
buf ( R_c4c_14874a18 , n35836 );
buf ( R_62d_123c23b8 , n35849 );
buf ( R_611_156aa558 , n35863 );
buf ( R_c30_13cd8158 , n35864 );
buf ( R_124f_13cd9418 , n35865 );
buf ( R_186e_1162cb38 , C0 );
buf ( R_1233_13d5c318 , n35866 );
buf ( R_1852_11635698 , C0 );
buf ( R_18a6_15885218 , C0 );
buf ( R_1287_13c29e98 , n35867 );
buf ( R_c68_12fc1cd8 , n35868 );
buf ( R_649_150e1f38 , n35894 );
buf ( R_5f5_13bf7398 , n35923 );
buf ( R_c14_13defe98 , n35924 );
buf ( R_18c2_13d5d998 , C0 );
buf ( R_bf8_13bf77f8 , n35925 );
buf ( R_12a3_14b20278 , n35926 );
buf ( R_1217_123bdd18 , n35927 );
buf ( R_c84_123bee98 , n35928 );
buf ( R_1836_14a16038 , C0 );
buf ( R_665_117eefb8 , n35956 );
buf ( R_5d9_15fed588 , n35981 );
buf ( R_84f_1587bdf8 , n35982 );
buf ( R_148d_156b2d98 , n36009 );
buf ( R_164c_156b65d8 , n36010 );
buf ( R_a0e_13cd5098 , C0 );
buf ( R_e6e_13c1e818 , C0 );
buf ( R_102d_14a14878 , n36018 );
buf ( R_d7b_1007dbb8 , n36019 );
buf ( R_1120_13cd3158 , n36020 );
buf ( R_139a_12fbf398 , C0 );
buf ( R_b01_1587af98 , n36068 );
buf ( R_19b9_116327b8 , n36076 );
buf ( R_75c_13d54b18 , n36077 );
buf ( R_173f_14a0d1b8 , n36078 );
buf ( R_ca0_117f3978 , n36079 );
buf ( R_bdc_14867a98 , n36080 );
buf ( R_11fb_13d26638 , n36081 );
buf ( R_681_13c02c58 , n36104 );
buf ( R_18de_1162c638 , C0 );
buf ( R_181a_15887fb8 , C0 );
buf ( R_12bf_12fbe3f8 , n36105 );
buf ( R_5bd_123b9678 , n36116 );
buf ( R_1a0e_1486b698 , C0 );
buf ( R_13ef_156ba1d8 , n36117 );
buf ( R_dd0_12fc0798 , n36118 );
buf ( R_7b1_14a13478 , n36145 );
buf ( R_aac_116311d8 , n36146 );
buf ( R_10cb_150dccb8 , n36147 );
buf ( R_16ea_140b6cb8 , C0 );
buf ( R_ffe_13ccf198 , C0 );
buf ( R_e9d_13d27038 , n36184 );
buf ( R_9df_14a17398 , n36185 );
buf ( R_161d_13b962b8 , n36191 );
buf ( R_14bc_117f0598 , n36192 );
buf ( R_87e_140b08b8 , C0 );
buf ( R_5a1_13d446b8 , n36197 );
buf ( R_cbc_12fc1b98 , n36198 );
buf ( R_bc0_13dfb338 , n36199 );
buf ( R_69d_11c69798 , n36223 );
buf ( R_18fa_140b5098 , C0 );
buf ( R_11df_15880998 , n36224 );
buf ( R_12db_156b4af8 , n36225 );
buf ( R_17fe_1580f5f8 , C0 );
buf ( R_191b_13c25f78 , n36226 );
buf ( R_580_1162b4b8 , n36227 );
buf ( R_6be_158101d8 , C0 );
buf ( R_17dd_14872358 , n36233 );
buf ( R_12fc_15813dd8 , n36234 );
buf ( R_b9f_140b49b8 , n36235 );
buf ( R_cdd_13bf42d8 , n36265 );
buf ( R_11be_150e4378 , C0 );
buf ( R_eba_13d29158 , C0 );
buf ( R_fe1_13d2bef8 , n36274 );
buf ( R_14d9_13c21338 , n36302 );
buf ( R_9c2_116297f8 , C0 );
buf ( R_89b_117ed118 , n36303 );
buf ( R_1600_117e96f8 , n36304 );
buf ( R_585_14a19b98 , n36305 );
buf ( R_1916_150e99b8 , C0 );
buf ( R_17e2_123c1d78 , C0 );
buf ( R_6b9_150dc998 , n36332 );
buf ( R_ba4_13c04d78 , n36333 );
buf ( R_12f7_117f4ff8 , n36334 );
buf ( R_11c3_117ee158 , n36335 );
buf ( R_cd8_150deab8 , n36336 );
buf ( R_15c4_13d46e18 , n36337 );
buf ( R_8d7_13de10b8 , n36338 );
buf ( R_fa5_13df4858 , n36355 );
buf ( R_ef6_13c1f358 , C0 );
buf ( R_986_11631278 , C0 );
buf ( R_1515_13ccb8b8 , n36365 );
buf ( R_11a7_123b9b78 , n36366 );
buf ( R_569_12fbfd98 , n36367 );
buf ( R_6d5_14b25958 , n36378 );
buf ( R_1313_1587dab8 , n36379 );
buf ( R_17c6_13d290b8 , C0 );
buf ( R_b88_14a0d9d8 , n36380 );
buf ( R_cf4_13bea558 , n36381 );
buf ( R_1932_13cd1538 , C0 );
buf ( R_1778_11631598 , n36382 );
buf ( R_d42_1580f918 , C0 );
buf ( R_1159_148722b8 , n36393 );
buf ( R_1361_14a18658 , n36422 );
buf ( R_b3a_11637678 , C0 );
buf ( R_1980_15883a58 , n36423 );
buf ( R_723_14a0aeb8 , n36424 );
buf ( R_ec5_123c1eb8 , n36481 );
buf ( R_fd6_15ff7448 , C0 );
buf ( R_14e4_14a121b8 , n36482 );
buf ( R_9b7_117eaaf8 , n36483 );
buf ( R_8a6_156b3018 , C0 );
buf ( R_15f5_140ade38 , n36523 );
buf ( R_d45_117f4418 , n36533 );
buf ( R_1775_140b5d18 , n36551 );
buf ( R_1364_13c1d918 , n36552 );
buf ( R_1156_15ff6fe8 , C0 );
buf ( R_1983_100863f8 , n36553 );
buf ( R_726_13d39498 , C0 );
buf ( R_b37_10089b98 , n36554 );
buf ( R_15e9_11636db8 , n36596 );
buf ( R_14f0_13b92398 , n36597 );
buf ( R_fca_156b44b8 , C0 );
buf ( R_8b2_11629078 , C0 );
buf ( R_9ab_14866698 , n36598 );
buf ( R_ed1_158870b8 , n36701 );
buf ( R_1632_117f1178 , C0 );
buf ( R_9f4_1486d2b8 , n36702 );
buf ( R_e88_124c4498 , n36703 );
buf ( R_1013_14a135b8 , n36705 );
buf ( R_14a7_15814af8 , n36706 );
buf ( R_869_14a19e18 , n36811 );
buf ( R_132f_13c0b8f8 , n36812 );
buf ( R_6f1_150df878 , n36836 );
buf ( R_118b_14b27618 , n36837 );
buf ( R_194e_14b236f8 , C0 );
buf ( R_d10_123b2d78 , n36838 );
buf ( R_b6c_123b8138 , n36839 );
buf ( R_17aa_13dfac58 , C0 );
buf ( R_188b_117e9978 , n36840 );
buf ( R_126c_1580edd8 , n36841 );
buf ( R_c4d_13d24b58 , n36853 );
buf ( R_62e_13bf7438 , C0 );
buf ( R_610_14a186f8 , n36855 );
buf ( R_c2f_14a0c038 , n36856 );
buf ( R_124e_117ee338 , C0 );
buf ( R_186d_15fee348 , n36905 );
buf ( R_e8c_1587e738 , n36906 );
buf ( R_162e_123b25f8 , C0 );
buf ( R_9f0_140abe58 , n36907 );
buf ( R_14ab_13dd50d8 , n36908 );
buf ( R_86d_14a18dd8 , n36916 );
buf ( R_100f_13d5dad8 , n36917 );
buf ( R_8f8_15ff8668 , n36918 );
buf ( R_f17_14a18e78 , n36919 );
buf ( R_1536_14a0dc58 , C0 );
buf ( R_15a3_12fc08d8 , n36920 );
buf ( R_f84_117e8d98 , n36921 );
buf ( R_965_140b2578 , n36929 );
buf ( R_d71_14b23018 , n36960 );
buf ( R_b0b_13c21e78 , n36961 );
buf ( R_1390_17016a08 , n36962 );
buf ( R_19af_11636458 , n36963 );
buf ( R_1749_117ec178 , n36969 );
buf ( R_752_15ff64a8 , C0 );
buf ( R_112a_1587e0f8 , C0 );
buf ( R_18b6_13bf3018 , C0 );
buf ( R_1223_13dd8418 , n36970 );
buf ( R_1297_13b99738 , n36971 );
buf ( R_1842_123b43f8 , C0 );
buf ( R_c78_15887018 , n36972 );
buf ( R_659_123b34f8 , n36984 );
buf ( R_5e5_13df0578 , n36995 );
buf ( R_c04_13cd6f38 , n36996 );
buf ( R_954_17014988 , n36997 );
buf ( R_909_13d3efd8 , n37005 );
buf ( R_f28_13bf6fd8 , n37006 );
buf ( R_1547_13df7b98 , n37007 );
buf ( R_1592_156b9918 , C0 );
buf ( R_f73_13d22a38 , n37008 );
buf ( R_70d_13beb098 , n37022 );
buf ( R_178e_13c1cb58 , C0 );
buf ( R_196a_156b6d58 , C0 );
buf ( R_d2c_14a0ec98 , n37023 );
buf ( R_116f_13d3e7b8 , n37024 );
buf ( R_134b_15ff6cc8 , n37025 );
buf ( R_b50_15815598 , n37026 );
buf ( R_caf_156adc58 , n37027 );
buf ( R_bcd_1162baf8 , n37062 );
buf ( R_690_13c1e098 , n37063 );
buf ( R_18ed_124c3278 , n37096 );
buf ( R_11ec_1008d0b8 , n37097 );
buf ( R_12ce_13c071b8 , C0 );
buf ( R_180b_1008abd8 , n37098 );
buf ( R_5ae_13cd7ed8 , n37103 );
buf ( R_177b_1007d6b8 , n37104 );
buf ( R_d3f_13cd10d8 , n37105 );
buf ( R_115c_150e8f18 , n37106 );
buf ( R_135e_11c696f8 , C0 );
buf ( R_b3d_13dddeb8 , n37431 );
buf ( R_720_13d395d8 , n37432 );
buf ( R_197d_14a15458 , n37440 );
buf ( R_1700_140ae8d8 , n37441 );
buf ( R_10e1_13c07758 , n37459 );
buf ( R_ac2_156ad2f8 , C0 );
buf ( R_79b_15886398 , n37460 );
buf ( R_dba_116373f8 , C0 );
buf ( R_13d9_14a14378 , n37471 );
buf ( R_19f8_117ef558 , n37472 );
buf ( R_595_13def178 , n37477 );
buf ( R_17f2_1580c998 , C0 );
buf ( R_1906_13ccad78 , C0 );
buf ( R_6a9_15ff4ba8 , n37487 );
buf ( R_bb4_117f4d78 , n37488 );
buf ( R_12e7_13cd42d8 , n37489 );
buf ( R_11d3_1162b0f8 , n37490 );
buf ( R_cc8_123b7738 , n37491 );
buf ( R_d48_13c21c98 , n37492 );
buf ( R_1772_14a16998 , C0 );
buf ( R_1367_15880858 , n37493 );
buf ( R_1153_117f1678 , n37494 );
buf ( R_1986_11c6c038 , C0 );
buf ( R_729_117f72f8 , n37518 );
buf ( R_b34_158825b8 , n37519 );
buf ( R_ff5_13c2a618 , n37534 );
buf ( R_ea6_150dd7f8 , C0 );
buf ( R_9d6_13c01f38 , C0 );
buf ( R_14c5_14a0e518 , n37548 );
buf ( R_1614_156b2b18 , n37549 );
buf ( R_887_14a18298 , n37550 );
buf ( R_848_13ddf218 , n37551 );
buf ( R_1653_14869438 , n37552 );
buf ( R_1486_156afe18 , C0 );
buf ( R_a15_1700ed08 , n37561 );
buf ( R_e67_117f4e18 , n37562 );
buf ( R_1034_156ac5d8 , n37563 );
buf ( R_8eb_150db1d8 , n37564 );
buf ( R_15b0_1580bdb8 , n37565 );
buf ( R_f0a_14a0ce98 , C0 );
buf ( R_f91_117f6f38 , n37574 );
buf ( R_1529_123bca58 , n37616 );
buf ( R_972_13ccc038 , C0 );
buf ( R_1a10_123b4718 , n37617 );
buf ( R_13f1_13d24298 , n37651 );
buf ( R_dd2_14a19198 , C0 );
buf ( R_7b3_13c07938 , n37652 );
buf ( R_aaa_13b8cfd8 , C0 );
buf ( R_10c9_15812a78 , n37657 );
buf ( R_16e8_13cd8d38 , n37658 );
buf ( R_d64_15ff5968 , n37659 );
buf ( R_b18_117f40f8 , n37660 );
buf ( R_1383_13c2a438 , n37661 );
buf ( R_19a2_117f01d8 , C0 );
buf ( R_1756_123c0f18 , C0 );
buf ( R_1137_13d20ff8 , n37662 );
buf ( R_745_13c1d5f8 , n37685 );
buf ( R_1636_14b22618 , C0 );
buf ( R_9f8_13decdd8 , n37686 );
buf ( R_e84_14875b98 , n37687 );
buf ( R_1017_13d3bbf8 , n37688 );
buf ( R_865_13d4e7b8 , n37693 );
buf ( R_14a3_11c6d078 , n37694 );
buf ( R_83e_13d43ad8 , C0 );
buf ( R_a1f_13d22d58 , n37695 );
buf ( R_147c_1580d398 , n37696 );
buf ( R_103e_13d57958 , C0 );
buf ( R_e5d_1486ddf8 , n37725 );
buf ( R_165d_13bec038 , n37806 );
buf ( R_1494_117f6718 , n37807 );
buf ( R_1645_11c6c178 , n37819 );
buf ( R_a07_14b251d8 , n37820 );
buf ( R_e75_1580a5f8 , n37884 );
buf ( R_1026_158103b8 , C0 );
buf ( R_856_13cd2a78 , C0 );
buf ( R_188c_13d39ad8 , n37885 );
buf ( R_126d_11636638 , n37915 );
buf ( R_c4e_13c0fe58 , C0 );
buf ( R_62f_116305f8 , n37916 );
buf ( R_60f_13bf44b8 , n37917 );
buf ( R_c2e_156b6c18 , C0 );
buf ( R_124d_123b5438 , n38002 );
buf ( R_186c_15817758 , n38003 );
buf ( R_57b_12fc1f58 , n38004 );
buf ( R_6c3_14a11718 , n38005 );
buf ( R_17d8_13bf24d8 , n38006 );
buf ( R_1301_13ccee78 , n38018 );
buf ( R_b9a_140b40f8 , C0 );
buf ( R_ce2_156b49b8 , C0 );
buf ( R_11b9_13d5d5d8 , n38032 );
buf ( R_1920_117ea198 , n38033 );
buf ( R_1713_14a0f878 , n38034 );
buf ( R_10f4_13de4c18 , n38035 );
buf ( R_ad5_117ed1b8 , n38044 );
buf ( R_788_117e8ed8 , n38045 );
buf ( R_da7_11635ff8 , n38046 );
buf ( R_13c6_123c10f8 , C0 );
buf ( R_19e5_1580eb58 , n38053 );
buf ( R_e90_11637038 , n38054 );
buf ( R_9ec_117eb958 , n38055 );
buf ( R_162a_117ec0d8 , C0 );
buf ( R_14af_156abdb8 , n38056 );
buf ( R_871_1587f138 , n38060 );
buf ( R_100b_11631d18 , n38061 );
buf ( R_111b_1580faf8 , n38062 );
buf ( R_139f_150df058 , n38063 );
buf ( R_afc_117f8158 , n38064 );
buf ( R_19be_13ccfff8 , C0 );
buf ( R_761_12fbf078 , n38087 );
buf ( R_173a_156b5a98 , C0 );
buf ( R_d80_13c1d418 , n38088 );
buf ( R_58a_13ddaf38 , n38089 );
buf ( R_1911_124c4038 , n38125 );
buf ( R_17e7_15883198 , n38126 );
buf ( R_6b4_15881bb8 , n38127 );
buf ( R_ba9_13d5c958 , n38162 );
buf ( R_12f2_17013c68 , C0 );
buf ( R_11c8_11634fb8 , n38163 );
buf ( R_cd3_13c06178 , n38164 );
buf ( R_6fc_13de34f8 , n38165 );
buf ( R_1180_13ddc298 , n38166 );
buf ( R_1959_14a14698 , n38188 );
buf ( R_d1b_13cd9558 , n38189 );
buf ( R_b61_13d22538 , n38224 );
buf ( R_179f_150e5818 , n38225 );
buf ( R_133a_13d57138 , C0 );
buf ( R_be4_15817bb8 , n38226 );
buf ( R_c98_13dec298 , n38227 );
buf ( R_1203_1587d978 , n38228 );
buf ( R_679_123b7918 , n38240 );
buf ( R_1822_117e9018 , C0 );
buf ( R_18d6_13c2ad98 , C0 );
buf ( R_5c5_1162b5f8 , n38255 );
buf ( R_12b7_117f83d8 , n38256 );
buf ( R_ca8_14a11038 , n38257 );
buf ( R_bd4_11637ad8 , n38258 );
buf ( R_689_158869d8 , n38268 );
buf ( R_11f3_116300f8 , n38269 );
buf ( R_18e6_156b1678 , C0 );
buf ( R_1812_11c6f558 , C0 );
buf ( R_12c7_13b97c58 , n38270 );
buf ( R_5b5_11637fd8 , n38271 );
buf ( R_177e_14b1a738 , C0 );
buf ( R_d3c_13b8b278 , n38272 );
buf ( R_115f_156ac7b8 , n38273 );
buf ( R_135b_13d38b38 , n38274 );
buf ( R_b40_158142d8 , n38275 );
buf ( R_71d_13c1ea98 , n38285 );
buf ( R_197a_13c0a318 , C0 );
buf ( R_e16_17018088 , C0 );
buf ( R_1085_13c03e78 , n38298 );
buf ( R_7f7_15888b98 , n38299 );
buf ( R_16a4_158821f8 , n38300 );
buf ( R_1a54_13de0438 , n38301 );
buf ( R_1435_10082258 , n38313 );
buf ( R_a66_15882838 , C0 );
buf ( R_703_14867bd8 , n38314 );
buf ( R_1960_1162c958 , n38315 );
buf ( R_1179_13d3c7d8 , n38358 );
buf ( R_d22_13d599d8 , C0 );
buf ( R_b5a_13bf68f8 , C0 );
buf ( R_1341_13d458d8 , n38369 );
buf ( R_1798_1700e9e8 , n38370 );
buf ( R_171e_13df60b8 , C0 );
buf ( R_10ff_13ddcab8 , n38371 );
buf ( R_ae0_14a11f38 , n38372 );
buf ( R_77d_13d27df8 , n38395 );
buf ( R_d9c_13ccd4d8 , n38396 );
buf ( R_13bb_1587d478 , n38397 );
buf ( R_19da_13dd5a38 , C0 );
buf ( R_108a_1486e938 , C0 );
buf ( R_e11_13cd8c98 , n38409 );
buf ( R_16a9_14a130b8 , n38417 );
buf ( R_7f2_156b2938 , C0 );
buf ( R_1a4f_13d3a618 , n38418 );
buf ( R_a6b_13b8e1f8 , n38419 );
buf ( R_1430_13dd84b8 , n38420 );
buf ( R_d4b_117f6178 , n38421 );
buf ( R_176f_13d447f8 , n38422 );
buf ( R_136a_13c26838 , C0 );
buf ( R_1150_15ff71c8 , n38423 );
buf ( R_1989_13ccbc78 , n38431 );
buf ( R_72c_10083c98 , n38432 );
buf ( R_b31_13d44c58 , n38449 );
buf ( R_814_13d51eb8 , n38450 );
buf ( R_1068_1580ea18 , n38451 );
buf ( R_1687_123b81d8 , n38452 );
buf ( R_1452_13df0938 , C0 );
buf ( R_e33_14a0c3f8 , n38453 );
buf ( R_a49_14a0eb58 , n38469 );
buf ( R_1851_13d5b058 , n38820 );
buf ( R_18a7_13b96858 , n38821 );
buf ( R_1288_13c1daf8 , n38822 );
buf ( R_c69_156af738 , n38847 );
buf ( R_64a_11629438 , C0 );
buf ( R_5f4_140b13f8 , n38848 );
buf ( R_c13_1162db78 , n38849 );
buf ( R_1232_156aaa58 , C0 );
buf ( R_15bb_117f3338 , n38850 );
buf ( R_8e0_14a0f698 , n38851 );
buf ( R_f9c_14a104f8 , n38852 );
buf ( R_eff_13d381d8 , n38853 );
buf ( R_151e_15883af8 , C0 );
buf ( R_97d_14a16178 , n38865 );
buf ( R_1702_13cd9198 , C0 );
buf ( R_10e3_117f2f78 , n38866 );
buf ( R_ac4_1700f028 , n38867 );
buf ( R_799_13d5a018 , n38879 );
buf ( R_db8_150e6998 , n38880 );
buf ( R_13d7_14b1d1b8 , n38881 );
buf ( R_19f6_1580aa58 , C0 );
buf ( R_14fd_156b56d8 , n38890 );
buf ( R_15dc_123bfd98 , n38891 );
buf ( R_fbd_14a0b098 , n38908 );
buf ( R_8bf_14875f58 , n38909 );
buf ( R_99e_15ff9388 , C0 );
buf ( R_ede_11634338 , C0 );
buf ( R_188d_17018e48 , n38934 );
buf ( R_126e_150e04f8 , C0 );
buf ( R_c4f_15814918 , n38935 );
buf ( R_630_13d25558 , n38936 );
buf ( R_60e_13cd3d38 , C0 );
buf ( R_c2d_1580aaf8 , n38958 );
buf ( R_124c_13d40018 , n38959 );
buf ( R_186b_13d42bd8 , n38960 );
buf ( R_1a23_13d52458 , n38961 );
buf ( R_1404_1486a8d8 , n38962 );
buf ( R_de5_11633a78 , n38972 );
buf ( R_7c6_156b9738 , C0 );
buf ( R_a97_13c05e58 , n38973 );
buf ( R_10b6_124c3638 , C0 );
buf ( R_16d5_123bc4b8 , n38987 );
buf ( R_bed_13b90db8 , n39019 );
buf ( R_c8f_117ef4b8 , n39020 );
buf ( R_120c_13ddcd38 , n39021 );
buf ( R_670_13ccfaf8 , n39022 );
buf ( R_182b_13cd80b8 , n39023 );
buf ( R_18cd_13c1ca18 , n39058 );
buf ( R_5ce_14b1ded8 , C0 );
buf ( R_12ae_13c1f178 , C0 );
buf ( R_bc6_13cd7bb8 , C0 );
buf ( R_697_13bf83d8 , n39059 );
buf ( R_18f4_15881cf8 , n39060 );
buf ( R_11e5_1162add8 , n39114 );
buf ( R_12d5_17015928 , n39125 );
buf ( R_1804_150e44b8 , n39126 );
buf ( R_5a7_12fbe178 , n39131 );
buf ( R_cb6_1162e398 , C0 );
buf ( R_110f_15887518 , n39132 );
buf ( R_19ca_156b8a18 , C0 );
buf ( R_af0_17012a48 , n39133 );
buf ( R_76d_156b1df8 , n39145 );
buf ( R_d8c_15814b98 , n39146 );
buf ( R_172e_117ed438 , C0 );
buf ( R_13ab_13b99878 , n39147 );
buf ( R_1a12_13d52ef8 , C0 );
buf ( R_13f3_156b74d8 , n39148 );
buf ( R_dd4_140ac5d8 , n39149 );
buf ( R_7b5_13c1f718 , n39165 );
buf ( R_aa8_14a0ea18 , n39166 );
buf ( R_10c7_13df2c38 , n39167 );
buf ( R_16e6_156b9eb8 , C0 );
buf ( R_15cd_13cd86f8 , n39214 );
buf ( R_8ce_13d1e2f8 , C0 );
buf ( R_fae_13bf6df8 , C0 );
buf ( R_eed_15812578 , n39224 );
buf ( R_98f_117f62b8 , n39225 );
buf ( R_150c_15ff3848 , n39226 );
buf ( R_908_123c0658 , n39227 );
buf ( R_f27_13cd08b8 , n39228 );
buf ( R_1546_14a18f18 , C0 );
buf ( R_1593_13d58e98 , n39229 );
buf ( R_f74_158805d8 , n39230 );
buf ( R_955_1580f0f8 , n39237 );
buf ( R_d5c_1580ed38 , n39238 );
buf ( R_137b_13d5cc78 , n39239 );
buf ( R_175e_15813478 , C0 );
buf ( R_199a_117e8b18 , C0 );
buf ( R_113f_123b3098 , n39240 );
buf ( R_73d_13c220f8 , n39249 );
buf ( R_b20_13c06c18 , n39250 );
buf ( R_163a_13d3ddb8 , C0 );
buf ( R_9fc_14a0b818 , n39251 );
buf ( R_e80_11633ed8 , n39252 );
buf ( R_101b_123b6518 , n39253 );
buf ( R_861_124c3bd8 , n39259 );
buf ( R_149f_123b5e38 , n39260 );
buf ( R_1080_14a149b8 , n39261 );
buf ( R_7fc_13d3f258 , n39262 );
buf ( R_169f_124c2d78 , n39263 );
buf ( R_1a59_117eded8 , n39269 );
buf ( R_143a_14a0edd8 , C0 );
buf ( R_a61_1700dd68 , n39286 );
buf ( R_e1b_13cd1178 , n39287 );
buf ( R_140f_117f1cb8 , n39288 );
buf ( R_df0_13c09cd8 , n39289 );
buf ( R_7d1_14b28978 , n39312 );
buf ( R_a8c_123c0338 , n39313 );
buf ( R_10ab_13df0398 , n39314 );
buf ( R_16ca_13d52f98 , C0 );
buf ( R_1a2e_13c22698 , C0 );
buf ( R_b10_14b21fd8 , n39315 );
buf ( R_138b_156b0318 , n39316 );
buf ( R_19aa_14a194b8 , C0 );
buf ( R_174e_15811a38 , C0 );
buf ( R_74d_117f0e58 , n39330 );
buf ( R_112f_156aac38 , n39331 );
buf ( R_d6c_156b62b8 , n39332 );
buf ( R_1781_1162d5d8 , n39379 );
buf ( R_d39_15811b78 , n39392 );
buf ( R_1162_124c2558 , C0 );
buf ( R_1358_156b8e78 , n39393 );
buf ( R_b43_13c06858 , n39394 );
buf ( R_71a_117ee798 , C0 );
buf ( R_1977_15880b78 , n39395 );
buf ( R_1108_13ccfb98 , n39396 );
buf ( R_ae9_1580cd58 , n39435 );
buf ( R_774_1700a7a8 , n39436 );
buf ( R_d93_13cce0b8 , n39437 );
buf ( R_13b2_15886898 , C0 );
buf ( R_1727_14870e18 , n39438 );
buf ( R_19d1_123b5b18 , n39446 );
buf ( R_188e_11c6a698 , C0 );
buf ( R_126f_14b23c98 , n39447 );
buf ( R_c50_13d471d8 , n39448 );
buf ( R_631_13ddd7d8 , n39458 );
buf ( R_60d_117f3a18 , n39470 );
buf ( R_c2c_13d2c498 , n39471 );
buf ( R_124b_156b97d8 , n39472 );
buf ( R_186a_13ddb118 , C0 );
buf ( R_fdc_1162ca98 , n39473 );
buf ( R_14de_13c202f8 , C0 );
buf ( R_9bd_11632cb8 , n39481 );
buf ( R_8a0_13bf81f8 , n39482 );
buf ( R_15fb_123ba078 , n39483 );
buf ( R_ebf_13b91678 , n39484 );
buf ( R_e94_148719f8 , n39485 );
buf ( R_9e8_15ff97e8 , n39486 );
buf ( R_1626_13de2918 , C0 );
buf ( R_14b3_13dde9f8 , n39487 );
buf ( R_875_156aea18 , n39488 );
buf ( R_1007_15881578 , n39489 );
buf ( R_14f6_11638938 , C0 );
buf ( R_fc4_1580d578 , n39490 );
buf ( R_8b8_123ba2f8 , n39491 );
buf ( R_9a5_117ecc18 , n39499 );
buf ( R_ed7_14a0da78 , n39500 );
buf ( R_15e3_123c0158 , n39501 );
buf ( R_e0c_1700d0e8 , n39502 );
buf ( R_16ae_123b38b8 , C0 );
buf ( R_7ed_117ef738 , n39510 );
buf ( R_1a4a_12fc1c38 , C0 );
buf ( R_a70_150dbc78 , n39511 );
buf ( R_142b_15889bd8 , n39512 );
buf ( R_108f_13de36d8 , n39513 );
buf ( R_d4e_11c6b6d8 , C0 );
buf ( R_176c_13ddfcb8 , n39514 );
buf ( R_136d_11634dd8 , n39524 );
buf ( R_114d_158861b8 , n39543 );
buf ( R_198c_13d53a38 , n39544 );
buf ( R_72f_11637498 , n39545 );
buf ( R_b2e_170098a8 , C0 );
buf ( R_8f7_13b8e298 , n39546 );
buf ( R_f16_1587d838 , C0 );
buf ( R_1535_13ded2d8 , n39581 );
buf ( R_15a4_1162bcd8 , n39582 );
buf ( R_f85_170174a8 , n39689 );
buf ( R_966_156acd58 , C0 );
buf ( R_12a4_13cd0db8 , n39690 );
buf ( R_1216_13c26518 , C0 );
buf ( R_c85_13d505b8 , n39713 );
buf ( R_1835_13b8eb58 , n39787 );
buf ( R_666_13cd8798 , C0 );
buf ( R_5d8_14a11fd8 , n39788 );
buf ( R_18c3_156b8c98 , n39789 );
buf ( R_bf7_156b4418 , n39790 );
buf ( R_15d5_117ed898 , n39828 );
buf ( R_fb6_14b24558 , C0 );
buf ( R_8c6_13d442f8 , C0 );
buf ( R_997_123bb478 , n39829 );
buf ( R_ee5_14a14af8 , n39858 );
buf ( R_1504_13d553d8 , n39859 );
buf ( R_6d1_158167b8 , n39868 );
buf ( R_130f_156ab4f8 , n39869 );
buf ( R_17ca_150df9b8 , C0 );
buf ( R_b8c_124c3ef8 , n39870 );
buf ( R_cf0_11c6a878 , n39871 );
buf ( R_192e_150e8a18 , C0 );
buf ( R_11ab_13d29d38 , n39872 );
buf ( R_56d_156b76b8 , n39873 );
buf ( R_1704_13bf4238 , n39874 );
buf ( R_10e5_14871778 , n39889 );
buf ( R_ac6_1587bcb8 , C0 );
buf ( R_797_14b1c178 , n39890 );
buf ( R_db6_13ddd058 , C0 );
buf ( R_13d5_1587c618 , n39903 );
buf ( R_19f4_150e3ab8 , n39904 );
buf ( R_1298_156b1d58 , n39905 );
buf ( R_1841_13d2c538 , n39922 );
buf ( R_c79_156b5598 , n39934 );
buf ( R_65a_14874ab8 , C0 );
buf ( R_5e4_13bf0278 , n39935 );
buf ( R_c03_14a0d2f8 , n39936 );
buf ( R_18b7_13ccd1b8 , n39937 );
buf ( R_1222_14b1acd8 , C0 );
buf ( R_1073_14b20f98 , n39938 );
buf ( R_809_13d3e678 , n39999 );
buf ( R_1a66_123b6158 , C0 );
buf ( R_1692_117f31f8 , C0 );
buf ( R_1447_13b93338 , n40000 );
buf ( R_e28_156abbd8 , n40001 );
buf ( R_a54_13cce838 , n40002 );
buf ( R_1054_13bf8ab8 , n40003 );
buf ( R_1466_13d5abf8 , C0 );
buf ( R_1673_1580e798 , n40004 );
buf ( R_e47_1587b178 , n40005 );
buf ( R_a35_117f5db8 , n40010 );
buf ( R_828_10081f38 , n40011 );
buf ( R_1469_1587ee18 , n40025 );
buf ( R_1051_11635c38 , n40074 );
buf ( R_e4a_11629118 , C0 );
buf ( R_1670_1007f238 , n40075 );
buf ( R_82b_13cd7258 , n40076 );
buf ( R_a32_1486afb8 , C0 );
buf ( R_1187_117f4198 , n40077 );
buf ( R_1952_14a0c0d8 , C0 );
buf ( R_d14_13dee778 , n40078 );
buf ( R_b68_10089d78 , n40079 );
buf ( R_17a6_15811f38 , C0 );
buf ( R_1333_117f21b8 , n40080 );
buf ( R_6f5_13d43678 , n40091 );
buf ( R_6c8_1580d758 , n40092 );
buf ( R_1306_1580d938 , C0 );
buf ( R_17d3_13d3a578 , n40093 );
buf ( R_b95_117f7618 , n40129 );
buf ( R_ce7_13d27218 , n40130 );
buf ( R_1925_15ff0328 , n40161 );
buf ( R_11b4_13b8ec98 , n40162 );
buf ( R_576_13d2bf98 , n40163 );
buf ( R_e00_13cd8bf8 , n40164 );
buf ( R_7e1_150e4058 , n40217 );
buf ( R_a7c_156b7118 , n40218 );
buf ( R_1a3e_14a0b278 , C0 );
buf ( R_109b_123bd4f8 , n40219 );
buf ( R_141f_1008c578 , n40220 );
buf ( R_16ba_156b6e98 , C0 );
buf ( R_188f_156b5458 , n40221 );
buf ( R_1270_14a103b8 , n40222 );
buf ( R_c51_11630af8 , n40233 );
buf ( R_632_13ccde38 , C0 );
buf ( R_60c_13dd9c78 , n40234 );
buf ( R_c2b_14b23478 , n40235 );
buf ( R_124a_140b7898 , C0 );
buf ( R_1869_14b29cd8 , n40289 );
buf ( R_1a14_117ebbd8 , n40290 );
buf ( R_13f5_13cd8a18 , n40302 );
buf ( R_dd6_13de0d98 , C0 );
buf ( R_7b7_15816a38 , n40303 );
buf ( R_aa6_13d28c58 , C0 );
buf ( R_10c5_11632998 , n40316 );
buf ( R_16e4_10087078 , n40317 );
buf ( R_190c_13d1d998 , n40318 );
buf ( R_6af_124c33b8 , n40319 );
buf ( R_bae_1587b5d8 , C0 );
buf ( R_12ed_14a176b8 , n40328 );
buf ( R_11cd_13cd27f8 , n40353 );
buf ( R_cce_116331b8 , C0 );
buf ( R_58f_156b9558 , n40354 );
buf ( R_17ec_13dd7fb8 , n40355 );
buf ( R_1057_123bd278 , n40356 );
buf ( R_1463_124c4b78 , n40357 );
buf ( R_1676_140ae6f8 , C0 );
buf ( R_e44_148741f8 , n40358 );
buf ( R_a38_150dc3f8 , n40359 );
buf ( R_825_123b3278 , n40400 );
buf ( R_18a8_1580c8f8 , n40401 );
buf ( R_1289_13c09738 , n40431 );
buf ( R_c6a_15811fd8 , C0 );
buf ( R_64b_1007d938 , n40432 );
buf ( R_5f3_116307d8 , n40433 );
buf ( R_c12_1162cc78 , C0 );
buf ( R_1231_13dee9f8 , n40465 );
buf ( R_1850_1587f778 , n40466 );
buf ( R_146c_14872f38 , n40467 );
buf ( R_104e_1580f7d8 , C0 );
buf ( R_e4d_14b20d18 , n40491 );
buf ( R_166d_13d20058 , n40499 );
buf ( R_82e_1580f2d8 , C0 );
buf ( R_a2f_123b3db8 , n40500 );
buf ( R_19c3_116340b8 , n40501 );
buf ( R_af7_13cd2d98 , n40502 );
buf ( R_766_13c07618 , C0 );
buf ( R_1735_13bf9f58 , n40507 );
buf ( R_d85_13dd7518 , n40517 );
buf ( R_13a4_150ea138 , n40518 );
buf ( R_1116_13c02438 , C0 );
buf ( R_df9_13dd9458 , n40531 );
buf ( R_7da_14a16fd8 , C0 );
buf ( R_a83_13b9a278 , n40532 );
buf ( R_10a2_123b3d18 , C0 );
buf ( R_1a37_1587f958 , n40533 );
buf ( R_16c1_13d3d458 , n40542 );
buf ( R_1418_13d2b1d8 , n40543 );
buf ( R_ea1_156b5c78 , n40580 );
buf ( R_9db_13c05bd8 , n40581 );
buf ( R_1619_15888d78 , n40587 );
buf ( R_14c0_17012fe8 , n40588 );
buf ( R_882_13dee458 , C0 );
buf ( R_ffa_11c68f78 , C0 );
buf ( R_1967_15ff9608 , n40589 );
buf ( R_1172_170122c8 , C0 );
buf ( R_d29_13bed898 , n40599 );
buf ( R_1348_156b1178 , n40600 );
buf ( R_b53_1162fe78 , n40601 );
buf ( R_1791_15ff73a8 , n40641 );
buf ( R_70a_13dee818 , C0 );
buf ( R_8ea_13b91c18 , C0 );
buf ( R_15b1_140b0d18 , n40673 );
buf ( R_f09_13d4f9d8 , n40679 );
buf ( R_f92_13b99238 , C0 );
buf ( R_1528_13cca918 , n40680 );
buf ( R_973_12fc1738 , n40681 );
buf ( R_907_13d1cef8 , n40682 );
buf ( R_f26_13d51378 , C0 );
buf ( R_1545_13ddab78 , n40713 );
buf ( R_1594_123b52f8 , n40714 );
buf ( R_f75_1587ec38 , n40733 );
buf ( R_956_117f3bf8 , C0 );
buf ( R_a1c_13d42098 , n40734 );
buf ( R_147f_15ffd208 , n40735 );
buf ( R_103b_12fbfbb8 , n40736 );
buf ( R_e60_13b98dd8 , n40737 );
buf ( R_165a_156b9418 , C0 );
buf ( R_841_13de1e78 , n40772 );
buf ( R_1715_13c03ab8 , n40787 );
buf ( R_10f6_1587fc78 , C0 );
buf ( R_ad7_11c6aaf8 , n40788 );
buf ( R_786_13bf7938 , C0 );
buf ( R_da5_13c24c18 , n40798 );
buf ( R_13c4_156adbb8 , n40799 );
buf ( R_19e3_13b8b4f8 , n40800 );
buf ( R_15c5_13cce478 , n40826 );
buf ( R_8d6_14a156d8 , C0 );
buf ( R_fa6_13ccd7f8 , C0 );
buf ( R_ef5_13c0f8b8 , n40896 );
buf ( R_987_148737f8 , n40897 );
buf ( R_1514_13d4ea38 , n40898 );
buf ( R_d36_13cd2938 , C0 );
buf ( R_1165_1700dae8 , n40912 );
buf ( R_1355_13c0e2d8 , n40923 );
buf ( R_b46_12fbedf8 , C0 );
buf ( R_717_13c1ebd8 , n40924 );
buf ( R_1974_13b938d8 , n40925 );
buf ( R_1784_14b1b3b8 , n40926 );
buf ( R_156d_13b91d58 , n40958 );
buf ( R_f4e_13d2bb38 , C0 );
buf ( R_156c_1486f8d8 , n40959 );
buf ( R_92f_1587e418 , n40960 );
buf ( R_f4d_158174d8 , n40990 );
buf ( R_92e_15880df8 , C0 );
buf ( R_156e_13bee0b8 , C0 );
buf ( R_f4f_13d1f298 , n40991 );
buf ( R_930_117f5818 , n40992 );
buf ( R_156b_13cd6a38 , n40993 );
buf ( R_f4c_13d4edf8 , n40994 );
buf ( R_92d_13b93838 , n41023 );
buf ( R_156f_1700c828 , n41024 );
buf ( R_f50_13d5d038 , n41025 );
buf ( R_931_1007f198 , n41049 );
buf ( R_92c_13bef238 , n41050 );
buf ( R_156a_14a0d7f8 , C0 );
buf ( R_f4b_1162df38 , n41051 );
buf ( R_682_13dd6a78 , C0 );
buf ( R_11fa_12fbfe38 , C0 );
buf ( R_18df_1162e1b8 , n41052 );
buf ( R_1819_117f44b8 , n41093 );
buf ( R_12c0_156b3478 , n41094 );
buf ( R_5bc_150db098 , n41095 );
buf ( R_ca1_15888af8 , n41105 );
buf ( R_bdb_123b9178 , n41106 );
buf ( R_1890_13c0a4f8 , n41107 );
buf ( R_1271_13cd3e78 , n41138 );
buf ( R_c52_11629cf8 , C0 );
buf ( R_633_1587c6b8 , n41139 );
buf ( R_60b_17014c08 , n41140 );
buf ( R_c2a_13c01d58 , C0 );
buf ( R_1249_150de798 , n41169 );
buf ( R_1868_13cd62b8 , n41170 );
buf ( R_105a_14a112b8 , C0 );
buf ( R_1460_158862f8 , n41171 );
buf ( R_1679_13cd44b8 , n41178 );
buf ( R_e41_14a14e18 , n41188 );
buf ( R_a3b_13cd1998 , n41189 );
buf ( R_822_117e9158 , C0 );
buf ( R_1570_13d44118 , n41190 );
buf ( R_f51_13ccb778 , n41212 );
buf ( R_932_15810d18 , C0 );
buf ( R_92b_14a180b8 , n41213 );
buf ( R_f4a_1162c8b8 , C0 );
buf ( R_1569_13bede38 , n41226 );
buf ( R_163e_12fc0338 , C0 );
buf ( R_a00_13df4df8 , n41227 );
buf ( R_e7c_13c08798 , n41228 );
buf ( R_101f_117ed9d8 , n41229 );
buf ( R_85d_117f4738 , n41235 );
buf ( R_149b_13cd1038 , n41236 );
buf ( R_146f_117f47d8 , n41237 );
buf ( R_104b_158885f8 , n41238 );
buf ( R_e50_12fbe858 , n41239 );
buf ( R_166a_1587c938 , C0 );
buf ( R_831_156b2398 , n41275 );
buf ( R_a2c_11c701d8 , n41276 );
buf ( R_801_150e6e98 , n41317 );
buf ( R_169a_13b94878 , C0 );
buf ( R_1a5e_1162d3f8 , C0 );
buf ( R_143f_13b8c218 , n41318 );
buf ( R_a5c_13b8c178 , n41319 );
buf ( R_e20_13ddd0f8 , n41320 );
buf ( R_107b_156b2118 , n41321 );
buf ( R_d51_13df3b38 , n41332 );
buf ( R_1769_14b21038 , n41349 );
buf ( R_1370_13cd2618 , n41350 );
buf ( R_114a_13c218d8 , C0 );
buf ( R_198f_13d28bb8 , n41351 );
buf ( R_732_13d55fb8 , C0 );
buf ( R_b2b_13ccd2f8 , n41352 );
buf ( R_1571_1580af58 , n41369 );
buf ( R_f52_12fc1ff8 , C0 );
buf ( R_933_14868718 , n41370 );
buf ( R_92a_13c01a38 , C0 );
buf ( R_f49_13d4f4d8 , n41393 );
buf ( R_1568_1580c218 , n41394 );
buf ( R_1706_15814eb8 , C0 );
buf ( R_10e7_14a160d8 , n41395 );
buf ( R_ac8_156afa58 , n41396 );
buf ( R_795_14a12b18 , n41407 );
buf ( R_db4_117edd98 , n41408 );
buf ( R_13d3_13b90f98 , n41409 );
buf ( R_19f2_12fbf258 , C0 );
buf ( R_17b9_156b0b38 , n41440 );
buf ( R_193f_13d3aa78 , n41441 );
buf ( R_b7b_13befeb8 , n41442 );
buf ( R_d01_140ab318 , n41467 );
buf ( R_119a_13b8a5f8 , C0 );
buf ( R_1320_14b27f78 , n41468 );
buf ( R_55c_11630e18 , n41469 );
buf ( R_6e2_158149b8 , C0 );
buf ( R_106b_117f3518 , n41470 );
buf ( R_168a_117eb598 , C0 );
buf ( R_144f_14b26718 , n41471 );
buf ( R_e30_123b3e58 , n41472 );
buf ( R_a4c_170172c8 , n41473 );
buf ( R_811_15882478 , n41509 );
buf ( R_1406_148665f8 , C0 );
buf ( R_de7_1007fcd8 , n41510 );
buf ( R_7c8_156b7f78 , n41511 );
buf ( R_a95_117f6cb8 , n41563 );
buf ( R_10b4_13d3d598 , n41564 );
buf ( R_16d3_1700be28 , n41565 );
buf ( R_1a25_13b9a318 , n41569 );
buf ( R_1572_156b67b8 , C0 );
buf ( R_f53_123c01f8 , n41570 );
buf ( R_934_156b0958 , n41571 );
buf ( R_929_13d5bf58 , n41588 );
buf ( R_f48_13c256b8 , n41589 );
buf ( R_1567_13b91e98 , n41590 );
buf ( R_1943_11c70598 , n41591 );
buf ( R_d05_13c0cd98 , n41600 );
buf ( R_b77_13d415f8 , n41601 );
buf ( R_17b5_14a12118 , n41615 );
buf ( R_1324_15887298 , n41616 );
buf ( R_6e6_13becb78 , C0 );
buf ( R_558_116299d8 , n41617 );
buf ( R_1196_13d4f398 , C0 );
buf ( R_e98_13d433f8 , n41618 );
buf ( R_9e4_13cccdf8 , n41619 );
buf ( R_1622_13c044b8 , C0 );
buf ( R_14b7_13d21318 , n41620 );
buf ( R_879_15884c78 , n41625 );
buf ( R_1003_124c39f8 , n41626 );
buf ( R_1a16_1486b418 , C0 );
buf ( R_13f7_13d24338 , n41627 );
buf ( R_dd8_1587fd18 , n41628 );
buf ( R_7b9_13c0f458 , n41638 );
buf ( R_aa4_13c1d0f8 , n41639 );
buf ( R_10c3_13ccbef8 , n41640 );
buf ( R_16e2_140b6df8 , C0 );
buf ( R_1573_14a0c498 , n41641 );
buf ( R_f54_11632858 , n41642 );
buf ( R_935_150e5318 , n41661 );
buf ( R_928_156aab98 , n41662 );
buf ( R_f47_13cd9238 , n41663 );
buf ( R_1566_123b2a58 , C0 );
buf ( R_a0b_11637858 , n41664 );
buf ( R_e71_14b21a38 , n41671 );
buf ( R_102a_11c6ccb8 , C0 );
buf ( R_852_14b1d938 , C0 );
buf ( R_1490_13bf8158 , n41672 );
buf ( R_1649_13dd4f98 , n41685 );
buf ( R_a12_1008b358 , C0 );
buf ( R_e6a_156b7a78 , C0 );
buf ( R_1031_14b25778 , n41694 );
buf ( R_84b_156ad1b8 , n41695 );
buf ( R_1650_13dd4e58 , n41696 );
buf ( R_1489_13c21978 , n41708 );
buf ( R_7e8_1486a0b8 , n41709 );
buf ( R_1a45_1162e2f8 , n41714 );
buf ( R_a75_156b0778 , n41729 );
buf ( R_1426_11637718 , C0 );
buf ( R_1094_13d28398 , n41730 );
buf ( R_16b3_117efeb8 , n41731 );
buf ( R_e07_13d453d8 , n41732 );
buf ( R_17bd_1162b918 , n41750 );
buf ( R_b7f_14a0be58 , n41751 );
buf ( R_cfd_13d1d038 , n41761 );
buf ( R_193b_13d39f38 , n41762 );
buf ( R_119e_13c1bcf8 , C0 );
buf ( R_560_12fbf118 , n41763 );
buf ( R_6de_13cd4058 , C0 );
buf ( R_131c_13c245d8 , n41764 );
buf ( R_1891_123b9858 , n41799 );
buf ( R_1272_13dd9ef8 , C0 );
buf ( R_c53_15ff5148 , n41800 );
buf ( R_634_11631818 , n41801 );
buf ( R_60a_156b2758 , C0 );
buf ( R_c29_13cd0598 , n41831 );
buf ( R_1248_12fbfcf8 , n41832 );
buf ( R_1867_14a0ded8 , n41833 );
buf ( R_9cd_13d1f518 , n41843 );
buf ( R_14ce_1008b5d8 , C0 );
buf ( R_160b_14b24cd8 , n41844 );
buf ( R_890_11628df8 , n41845 );
buf ( R_fec_13ccc5d8 , n41846 );
buf ( R_eaf_13d5baf8 , n41847 );
buf ( R_15bc_15889138 , n41848 );
buf ( R_8df_11637358 , n41849 );
buf ( R_f9d_158889b8 , n41861 );
buf ( R_efe_11632b78 , C0 );
buf ( R_97e_13c29718 , C0 );
buf ( R_151d_1700bc48 , n41870 );
buf ( R_ae2_123bdef8 , C0 );
buf ( R_77b_17011828 , n41871 );
buf ( R_d9a_13c047d8 , C0 );
buf ( R_13b9_15ffc948 , n41882 );
buf ( R_19d8_14870b98 , n41883 );
buf ( R_1720_156b9198 , n41884 );
buf ( R_1101_140b7398 , n41931 );
buf ( R_1202_15881898 , C0 );
buf ( R_67a_13de2878 , C0 );
buf ( R_1821_117f1c18 , n41974 );
buf ( R_18d7_1580f378 , n41975 );
buf ( R_5c4_14868fd8 , n41976 );
buf ( R_12b8_11631b38 , n41977 );
buf ( R_be3_13de2198 , n41978 );
buf ( R_c99_13c029d8 , n41990 );
buf ( R_fd1_13c1d058 , n42009 );
buf ( R_14e9_14868538 , n42038 );
buf ( R_9b2_1580b6d8 , C0 );
buf ( R_8ab_14a0fc38 , n42039 );
buf ( R_15f0_140ae3d8 , n42040 );
buf ( R_eca_14a11df8 , C0 );
buf ( R_1574_13cd7cf8 , n42041 );
buf ( R_f55_14b1ac38 , n42060 );
buf ( R_936_140acf38 , C0 );
buf ( R_927_124c4178 , n42061 );
buf ( R_f46_14a0af58 , C0 );
buf ( R_1565_1700e808 , n42126 );
buf ( R_14d3_1580e5b8 , n42127 );
buf ( R_9c8_15fef248 , n42128 );
buf ( R_895_13d532b8 , n42157 );
buf ( R_1606_1007ef18 , C0 );
buf ( R_eb4_117eda78 , n42158 );
buf ( R_fe7_1162ba58 , n42159 );
buf ( R_8f6_156b7b18 , C0 );
buf ( R_f15_158819d8 , n42168 );
buf ( R_15a5_158168f8 , n42185 );
buf ( R_1534_123b9c18 , n42186 );
buf ( R_f86_13c1ce78 , C0 );
buf ( R_967_11c68938 , n42187 );
buf ( R_1901_15817ed8 , n42218 );
buf ( R_6a4_1162c1d8 , n42219 );
buf ( R_bb9_156ab1d8 , n42231 );
buf ( R_12e2_11636a98 , C0 );
buf ( R_11d8_156aa738 , n42232 );
buf ( R_cc3_15887c98 , n42233 );
buf ( R_59a_117f76b8 , n42238 );
buf ( R_17f7_117e9838 , n42239 );
buf ( R_105d_123b4998 , n42252 );
buf ( R_145d_123bec18 , n42264 );
buf ( R_167c_140b6178 , n42265 );
buf ( R_e3e_150da7d8 , C0 );
buf ( R_a3e_11635cd8 , C0 );
buf ( R_81f_156b45f8 , n42266 );
buf ( R_120b_13def358 , n42267 );
buf ( R_671_140b4058 , n42276 );
buf ( R_182a_117ef698 , C0 );
buf ( R_18ce_156b4e18 , C0 );
buf ( R_5cd_14a185b8 , n42278 );
buf ( R_12af_15ff69a8 , n42279 );
buf ( R_bec_124c2878 , n42280 );
buf ( R_c90_117eb778 , n42281 );
buf ( R_1386_14a0c7b8 , C0 );
buf ( R_19a5_1008a598 , n42289 );
buf ( R_1753_13cd1218 , n42290 );
buf ( R_748_13d3b518 , n42291 );
buf ( R_1134_1580ad78 , n42292 );
buf ( R_d67_13d3caf8 , n42293 );
buf ( R_b15_156b2078 , n42303 );
buf ( R_128a_15880718 , C0 );
buf ( R_c6b_14a13518 , n42304 );
buf ( R_64c_148739d8 , n42305 );
buf ( R_5f2_13dd5538 , C0 );
buf ( R_c11_15ff5aa8 , n42334 );
buf ( R_1230_124c42b8 , n42335 );
buf ( R_184f_1587fa98 , n42336 );
buf ( R_18a9_11c6f918 , n42347 );
buf ( R_bbf_1587ddd8 , n42348 );
buf ( R_69e_123b5bb8 , C0 );
buf ( R_18fb_13df16f8 , n42349 );
buf ( R_11de_10089058 , C0 );
buf ( R_12dc_13c0bc18 , n42350 );
buf ( R_17fd_13d408d8 , n42391 );
buf ( R_5a0_11631db8 , n42396 );
buf ( R_cbd_14872df8 , n42407 );
buf ( R_691_15883378 , n42417 );
buf ( R_18ee_14a171b8 , C0 );
buf ( R_11eb_13d4f078 , n42418 );
buf ( R_12cf_158850d8 , n42419 );
buf ( R_180a_13d3fc58 , C0 );
buf ( R_5ad_14a0c2b8 , n42424 );
buf ( R_cb0_13de1658 , n42425 );
buf ( R_bcc_13df1f18 , n42426 );
buf ( R_1472_13d3c698 , C0 );
buf ( R_1048_13df8bd8 , n42427 );
buf ( R_e53_10087b18 , n42428 );
buf ( R_1667_13beaf58 , n42429 );
buf ( R_834_15888698 , n42430 );
buf ( R_a29_13de0618 , n42440 );
buf ( R_1575_13d42598 , n42466 );
buf ( R_f56_13c0c578 , C0 );
buf ( R_937_15886c58 , n42467 );
buf ( R_926_158846d8 , C0 );
buf ( R_f45_13d4f438 , n42488 );
buf ( R_1564_1587b038 , n42489 );
buf ( R_906_14a145f8 , C0 );
buf ( R_f25_13d24e78 , n42508 );
buf ( R_1544_124c4fd8 , n42509 );
buf ( R_1595_14b1f698 , n42514 );
buf ( R_f76_117f6fd8 , C0 );
buf ( R_957_15888878 , n42515 );
buf ( R_c7a_140ac998 , C0 );
buf ( R_65b_1580b778 , n42516 );
buf ( R_5e3_117eba98 , n42517 );
buf ( R_c02_123b2f58 , C0 );
buf ( R_18b8_12fc05b8 , n42518 );
buf ( R_1221_15812cf8 , n42557 );
buf ( R_1299_14b1fc38 , n42588 );
buf ( R_1840_13d549d8 , n42589 );
buf ( R_1947_156ac3f8 , n42590 );
buf ( R_d09_150dd438 , n42599 );
buf ( R_b73_117f7938 , n42600 );
buf ( R_17b1_14a0dcf8 , n42646 );
buf ( R_1328_13d2aeb8 , n42647 );
buf ( R_6ea_123bbb58 , C0 );
buf ( R_1192_1587dbf8 , C0 );
buf ( R_137e_13c27738 , C0 );
buf ( R_175b_15883ff8 , n42648 );
buf ( R_199d_1008a6d8 , n42656 );
buf ( R_113c_13d20eb8 , n42657 );
buf ( R_740_13bf6b78 , n42658 );
buf ( R_b1d_123c1918 , n42697 );
buf ( R_d5f_15888c38 , n42698 );
buf ( R_fcb_13def8f8 , n42699 );
buf ( R_8b1_170124a8 , n42726 );
buf ( R_9ac_14a190f8 , n42727 );
buf ( R_ed0_13d23d98 , n42728 );
buf ( R_15ea_1580e658 , C0 );
buf ( R_14ef_123bead8 , n42729 );
buf ( R_d33_123bd8b8 , n42730 );
buf ( R_1168_156b6fd8 , n42731 );
buf ( R_1352_13c10b78 , C0 );
buf ( R_b49_14a158b8 , n42753 );
buf ( R_714_1587c898 , n42754 );
buf ( R_1971_13ddfe98 , n42762 );
buf ( R_1787_1486e2f8 , n42763 );
buf ( R_68a_14a15b38 , C0 );
buf ( R_11f2_1162a6f8 , C0 );
buf ( R_18e7_13c08c98 , n42764 );
buf ( R_1811_117e9a18 , n42778 );
buf ( R_12c8_140aa878 , n42779 );
buf ( R_5b4_140b2a78 , n42780 );
buf ( R_ca9_15887e78 , n42789 );
buf ( R_bd3_13c0e9b8 , n42790 );
buf ( R_195d_15884818 , n42798 );
buf ( R_117c_14874838 , n42799 );
buf ( R_d1f_1007f698 , n42800 );
buf ( R_b5d_123bb8d8 , n42862 );
buf ( R_133e_13d55dd8 , C0 );
buf ( R_179b_12fbde58 , n42863 );
buf ( R_700_13cd9878 , n42864 );
buf ( R_1576_1700c6e8 , C0 );
buf ( R_f57_14a14198 , n42865 );
buf ( R_938_13bedc58 , n42866 );
buf ( R_925_13df1338 , n42877 );
buf ( R_f44_156b99b8 , n42878 );
buf ( R_1563_158841d8 , n42879 );
buf ( R_c86_14a12e38 , C0 );
buf ( R_1834_13cd3f18 , n42880 );
buf ( R_667_1486b558 , n42881 );
buf ( R_5d7_156b0c78 , n42882 );
buf ( R_18c4_11c709f8 , n42883 );
buf ( R_bf6_11c6f378 , C0 );
buf ( R_12a5_1162d718 , n42915 );
buf ( R_1215_117f51d8 , n42927 );
buf ( R_1892_13d3b1f8 , C0 );
buf ( R_1273_13dd5c18 , n42928 );
buf ( R_c54_13becd58 , n42929 );
buf ( R_635_13d2c678 , n42941 );
buf ( R_609_1580ef18 , n42952 );
buf ( R_c28_140ba098 , n42953 );
buf ( R_1247_13ccda78 , n42954 );
buf ( R_1866_13bf9eb8 , C0 );
buf ( R_9d2_13ccb958 , C0 );
buf ( R_14c9_117f80b8 , n42966 );
buf ( R_1610_1700a988 , n42967 );
buf ( R_88b_1587e5f8 , n42968 );
buf ( R_ff1_13b8bd18 , n42977 );
buf ( R_eaa_13dd6618 , C0 );
buf ( R_1708_11630558 , n42978 );
buf ( R_10e9_123c2138 , n42992 );
buf ( R_aca_14a131f8 , C0 );
buf ( R_793_12fc2138 , n42993 );
buf ( R_db2_123b68d8 , C0 );
buf ( R_13d1_156ac998 , n43007 );
buf ( R_19f0_13d47138 , n43008 );
buf ( R_7d3_13dd99f8 , n43009 );
buf ( R_a8a_150e0ef8 , C0 );
buf ( R_10a9_1486ae78 , n43013 );
buf ( R_16c8_13dfaed8 , n43014 );
buf ( R_1a30_14a19698 , n43015 );
buf ( R_1411_13dfa438 , n43026 );
buf ( R_df2_150e09f8 , C0 );
buf ( R_14e3_11634838 , n43027 );
buf ( R_9b8_13d43b78 , n43028 );
buf ( R_8a5_13bee798 , n43056 );
buf ( R_15f6_117f0458 , C0 );
buf ( R_ec4_11c68a78 , n43057 );
buf ( R_fd7_116387f8 , n43058 );
buf ( R_17c1_13d57d18 , n43070 );
buf ( R_b83_13bedd98 , n43071 );
buf ( R_cf9_1587d798 , n43083 );
buf ( R_1937_150e3c98 , n43084 );
buf ( R_11a2_13c05138 , C0 );
buf ( R_564_15815278 , n43085 );
buf ( R_6da_13c00f98 , C0 );
buf ( R_1318_1008a9f8 , n43086 );
buf ( R_faf_158866b8 , n43087 );
buf ( R_8cd_15ff2ee8 , n43122 );
buf ( R_eec_117f7078 , n43123 );
buf ( R_990_11633c58 , n43124 );
buf ( R_150b_13cd8dd8 , n43125 );
buf ( R_15ce_13df0898 , C0 );
buf ( R_1766_116318b8 , C0 );
buf ( R_1373_15810598 , n43126 );
buf ( R_1147_13b8d438 , n43127 );
buf ( R_1992_13b8d1b8 , C0 );
buf ( R_735_13cd4cd8 , n43139 );
buf ( R_b28_1162fab8 , n43140 );
buf ( R_d54_150e15d8 , n43141 );
buf ( R_1577_13d44ed8 , n43142 );
buf ( R_f58_13d3e178 , n43143 );
buf ( R_939_123b2878 , n43165 );
buf ( R_924_140b7118 , n43166 );
buf ( R_f43_140aeab8 , n43167 );
buf ( R_1562_100874d8 , C0 );
buf ( R_17ce_13d50b58 , C0 );
buf ( R_b90_14a17e38 , n43168 );
buf ( R_cec_156b8fb8 , n43169 );
buf ( R_192a_13df93f8 , C0 );
buf ( R_11af_156b2a78 , n43170 );
buf ( R_571_13b96ad8 , n43171 );
buf ( R_6cd_150dc5d8 , n43184 );
buf ( R_130b_14b1eab8 , n43185 );
buf ( R_19b7_117f7758 , n43186 );
buf ( R_75a_150de5b8 , C0 );
buf ( R_1741_100824d8 , n43202 );
buf ( R_d79_1008a638 , n43214 );
buf ( R_1122_150e9a58 , C0 );
buf ( R_1398_10083978 , n43215 );
buf ( R_b03_158129d8 , n43216 );
buf ( R_14d8_13cd4698 , n43217 );
buf ( R_9c3_13befa58 , n43218 );
buf ( R_89a_117edb18 , C0 );
buf ( R_1601_13d272b8 , n43248 );
buf ( R_eb9_11638438 , n43280 );
buf ( R_fe2_13defdf8 , C0 );
buf ( R_13f9_1580cb78 , n43291 );
buf ( R_dda_117f7118 , C0 );
buf ( R_7bb_13bf54f8 , n43292 );
buf ( R_aa2_12fc1a58 , C0 );
buf ( R_10c1_13b901d8 , n43297 );
buf ( R_16e0_158811b8 , n43298 );
buf ( R_1a18_156b8bf8 , n43299 );
buf ( R_fbe_13cd90f8 , C0 );
buf ( R_8be_13df3278 , C0 );
buf ( R_99f_123b6b58 , n43300 );
buf ( R_edd_13b99cd8 , n43307 );
buf ( R_15dd_156aef18 , n43333 );
buf ( R_14fc_140b09f8 , n43334 );
buf ( R_19b2_150e0318 , C0 );
buf ( R_1746_123b75f8 , C0 );
buf ( R_755_14a13338 , n43346 );
buf ( R_1127_13de3318 , n43347 );
buf ( R_d74_17011d28 , n43348 );
buf ( R_b08_150dce98 , n43350 );
buf ( R_1393_11c68c58 , n43351 );
buf ( R_1956_15813158 , C0 );
buf ( R_d18_156b9698 , n43352 );
buf ( R_b64_156b3a18 , n43353 );
buf ( R_17a2_117e8758 , C0 );
buf ( R_1337_13d20af8 , n43354 );
buf ( R_6f9_17012b88 , n43365 );
buf ( R_1183_1580f698 , n43366 );
buf ( R_bb3_17013d08 , n43367 );
buf ( R_12e8_14b1e158 , n43368 );
buf ( R_11d2_124c3318 , C0 );
buf ( R_cc9_11c6e018 , n43377 );
buf ( R_594_13cd9698 , n43382 );
buf ( R_17f1_13c0bdf8 , n43392 );
buf ( R_1907_13ccaa58 , n43393 );
buf ( R_6aa_13de4038 , C0 );
buf ( R_ba3_13cd5bd8 , n43394 );
buf ( R_12f8_13cd2758 , n43395 );
buf ( R_11c2_13c1fc18 , C0 );
buf ( R_cd9_14b1f878 , n43407 );
buf ( R_584_12fc0bf8 , n43408 );
buf ( R_1917_13d21f98 , n43409 );
buf ( R_17e1_13d37878 , n43419 );
buf ( R_6ba_11637b78 , C0 );
buf ( R_8e9_13cd6b78 , n43449 );
buf ( R_15b2_117f08b8 , C0 );
buf ( R_f08_156b5db8 , n43450 );
buf ( R_f93_13b92758 , n43451 );
buf ( R_1527_13ccaeb8 , n43452 );
buf ( R_974_13c0c2f8 , n43453 );
buf ( R_ad9_150e2a78 , n43464 );
buf ( R_784_13dfa4d8 , n43465 );
buf ( R_da3_14a0cd58 , n43466 );
buf ( R_13c2_13d2a4b8 , C0 );
buf ( R_19e1_1700c5a8 , n43470 );
buf ( R_1717_13df61f8 , n43471 );
buf ( R_10f8_156b7258 , n43472 );
buf ( R_1578_123bab18 , n43473 );
buf ( R_f59_13c10358 , n43495 );
buf ( R_93a_1486f978 , C0 );
buf ( R_923_11632178 , n43496 );
buf ( R_f42_14b1f9b8 , C0 );
buf ( R_1561_13bf4a58 , n43504 );
buf ( R_1060_13c0b358 , n43505 );
buf ( R_145a_14a12bb8 , C0 );
buf ( R_167f_14a19378 , n43506 );
buf ( R_e3b_13dd7f18 , n43507 );
buf ( R_a41_14a10d18 , n43520 );
buf ( R_81c_13bf79d8 , n43521 );
buf ( R_12fd_1007d9d8 , n43532 );
buf ( R_b9e_123ba618 , C0 );
buf ( R_cde_13d39218 , C0 );
buf ( R_11bd_11c6dcf8 , n43550 );
buf ( R_191c_1580c038 , n43551 );
buf ( R_57f_158160d8 , n43552 );
buf ( R_6bf_13df4e98 , n43553 );
buf ( R_17dc_15ff5508 , n43554 );
buf ( R_1893_117f0d18 , n43555 );
buf ( R_1274_156b1218 , n43556 );
buf ( R_c55_13cce338 , n43568 );
buf ( R_636_123c1238 , C0 );
buf ( R_608_13d58678 , n43569 );
buf ( R_c27_13bf2a78 , n43570 );
buf ( R_1246_14b229d8 , C0 );
buf ( R_1865_156b4d78 , n43605 );
buf ( R_772_11634a18 , C0 );
buf ( R_d91_13c0fdb8 , n43614 );
buf ( R_13b0_1486d0d8 , n43615 );
buf ( R_1729_123b6338 , n43631 );
buf ( R_19cf_11c70c78 , n43632 );
buf ( R_110a_156b12b8 , C0 );
buf ( R_aeb_11638758 , n43633 );
buf ( R_e78_117ef0f8 , n43634 );
buf ( R_1023_15ff3ac8 , n43635 );
buf ( R_859_13c0f098 , n43648 );
buf ( R_1497_116337f8 , n43649 );
buf ( R_1642_1162e578 , C0 );
buf ( R_a04_13c22e18 , n43650 );
buf ( R_76b_13ddaad8 , n43651 );
buf ( R_d8a_10085458 , C0 );
buf ( R_1730_11c6fd78 , n43652 );
buf ( R_13a9_15887978 , n43663 );
buf ( R_1111_11629c58 , n43704 );
buf ( R_19c8_123b61f8 , n43705 );
buf ( R_af2_11635558 , C0 );
buf ( R_1045_13c2abb8 , n43719 );
buf ( R_e56_13c1f0d8 , C0 );
buf ( R_1664_1700d9a8 , n43720 );
buf ( R_837_13d43c18 , n43721 );
buf ( R_a26_13c28c78 , C0 );
buf ( R_1475_123b8bd8 , n43733 );
buf ( R_e63_156b1358 , n43734 );
buf ( R_1038_10085f98 , n43735 );
buf ( R_1657_13cd2c58 , n43736 );
buf ( R_844_117f3ab8 , n43737 );
buf ( R_1482_140b29d8 , C0 );
buf ( R_a19_156ad4d8 , n43741 );
buf ( R_18f5_1587d518 , n43769 );
buf ( R_11e4_158159f8 , n43770 );
buf ( R_12d6_11c6c5d8 , C0 );
buf ( R_1803_123b54d8 , n43771 );
buf ( R_5a6_13ccf5f8 , n43776 );
buf ( R_cb7_1162c458 , n43777 );
buf ( R_bc5_14a0c5d8 , n43790 );
buf ( R_698_14a0feb8 , n43791 );
buf ( R_194b_15882658 , n43792 );
buf ( R_d0d_1580bef8 , n43802 );
buf ( R_b6f_117eb638 , n43803 );
buf ( R_17ad_156b4f58 , n43845 );
buf ( R_132c_158823d8 , n43846 );
buf ( R_6ee_14a0faf8 , C0 );
buf ( R_118e_156ab3b8 , C0 );
buf ( R_75f_14870918 , n43847 );
buf ( R_173c_123b9218 , n43848 );
buf ( R_d7e_11634018 , C0 );
buf ( R_111d_13beeb58 , n43887 );
buf ( R_139d_100868f8 , n43899 );
buf ( R_afe_15ff7ee8 , C0 );
buf ( R_19bc_17010248 , n43900 );
buf ( R_1175_11634c98 , n43941 );
buf ( R_d26_1587cf78 , C0 );
buf ( R_b56_13c236d8 , C0 );
buf ( R_1345_13cd4738 , n43952 );
buf ( R_1794_15813338 , n43953 );
buf ( R_707_13d580d8 , n43954 );
buf ( R_1964_13d42b38 , n43955 );
buf ( R_f24_13b92938 , n43956 );
buf ( R_1543_15ff0828 , n43957 );
buf ( R_1596_15ff8a28 , C0 );
buf ( R_f77_158124d8 , n43958 );
buf ( R_958_13df5bb8 , n43959 );
buf ( R_905_13d4f758 , n43967 );
buf ( R_1579_13b8d078 , n43973 );
buf ( R_f5a_15884d18 , C0 );
buf ( R_93b_1580c3f8 , n43974 );
buf ( R_922_140af198 , C0 );
buf ( R_f41_156b7cf8 , n44008 );
buf ( R_1560_14a14cd8 , n44009 );
buf ( R_c6c_14b20318 , n44010 );
buf ( R_64d_13ccebf8 , n44022 );
buf ( R_5f1_15814c38 , n44031 );
buf ( R_c10_15817898 , n44032 );
buf ( R_122f_13d22038 , n44033 );
buf ( R_184e_14b1b8b8 , C0 );
buf ( R_18aa_11638b18 , C0 );
buf ( R_128b_1587eaf8 , n44034 );
buf ( R_1695_14a12ed8 , n44050 );
buf ( R_1a63_1486ec58 , n44051 );
buf ( R_1444_15ff0788 , n44052 );
buf ( R_a57_13d5aa18 , n44053 );
buf ( R_e25_14a17078 , n44062 );
buf ( R_1076_1587b678 , C0 );
buf ( R_806_14a0bd18 , C0 );
buf ( R_fb7_15887158 , n44063 );
buf ( R_8c5_1008b2b8 , n44086 );
buf ( R_998_13d573b8 , n44087 );
buf ( R_ee4_15ff7da8 , n44088 );
buf ( R_1503_150daf58 , n44089 );
buf ( R_15d6_117ed398 , C0 );
buf ( R_7ca_150de978 , C0 );
buf ( R_a93_156af4b8 , n44090 );
buf ( R_10b2_100826b8 , C0 );
buf ( R_16d1_156b27f8 , n44103 );
buf ( R_1a27_13cd2118 , n44104 );
buf ( R_1408_1587fbd8 , n44105 );
buf ( R_de9_13cd12b8 , n44115 );
buf ( R_9e0_15ffc9e8 , n44116 );
buf ( R_161e_123b8a98 , C0 );
buf ( R_14bb_10081cb8 , n44117 );
buf ( R_87d_123b9498 , n44122 );
buf ( R_fff_12fbe5d8 , n44123 );
buf ( R_e9c_13df34f8 , n44124 );
buf ( R_ba8_123c12d8 , n44125 );
buf ( R_12f3_11634f18 , n44126 );
buf ( R_11c7_17013b28 , n44127 );
buf ( R_cd4_13c2b018 , n44128 );
buf ( R_589_14a19058 , n44129 );
buf ( R_1912_156aacd8 , C0 );
buf ( R_17e6_140b2758 , C0 );
buf ( R_6b5_1587d658 , n44143 );
buf ( R_f14_13d26458 , n44144 );
buf ( R_15a6_1162eb18 , C0 );
buf ( R_1533_14b268f8 , n44145 );
buf ( R_f87_11637998 , n44146 );
buf ( R_968_13d2b958 , n44147 );
buf ( R_8f5_13bebe58 , n44165 );
buf ( R_8d5_150e1c18 , n44194 );
buf ( R_fa7_12fbff78 , n44195 );
buf ( R_ef4_1162ea78 , n44196 );
buf ( R_988_15814198 , n44197 );
buf ( R_1513_13c06498 , n44198 );
buf ( R_15c6_12fbf2f8 , C0 );
buf ( R_8b7_15ffa468 , n44199 );
buf ( R_9a6_13d46058 , C0 );
buf ( R_ed6_13d57598 , C0 );
buf ( R_15e4_156aeb58 , n44200 );
buf ( R_14f5_13c29178 , n44208 );
buf ( R_fc5_13b8d258 , n44224 );
buf ( R_acc_13df8638 , n44225 );
buf ( R_791_13d42818 , n44234 );
buf ( R_db0_13bf9418 , n44235 );
buf ( R_13cf_123c2318 , n44236 );
buf ( R_19ee_11630cd8 , C0 );
buf ( R_170a_13d25698 , C0 );
buf ( R_10eb_13debbb8 , n44237 );
buf ( R_19ad_1587f9f8 , n44245 );
buf ( R_174b_15ff3528 , n44246 );
buf ( R_750_1008c9d8 , n44247 );
buf ( R_112c_13c015d8 , n44248 );
buf ( R_d6f_117eae18 , n44249 );
buf ( R_b0d_13d41c38 , n44286 );
buf ( R_138e_158113f8 , C0 );
buf ( R_168d_156b2f78 , n44301 );
buf ( R_144c_14a0dbb8 , n44302 );
buf ( R_e2d_1587d3d8 , n44312 );
buf ( R_a4f_15814418 , n44313 );
buf ( R_80e_156ac218 , C0 );
buf ( R_106e_14a15318 , C0 );
buf ( R_157a_156b4198 , C0 );
buf ( R_f5b_1162d7b8 , n44314 );
buf ( R_93c_13b933d8 , n44315 );
buf ( R_921_15813298 , n44326 );
buf ( R_f40_13cd1fd8 , n44327 );
buf ( R_155f_148745b8 , n44328 );
buf ( R_1275_13d26bd8 , n44358 );
buf ( R_c56_12fbf438 , C0 );
buf ( R_637_14b20db8 , n44359 );
buf ( R_607_15886258 , n44360 );
buf ( R_c26_13d3ac58 , C0 );
buf ( R_1245_13d261d8 , n44371 );
buf ( R_1864_13ddb2f8 , n44372 );
buf ( R_1894_13cd6998 , n44373 );
buf ( R_9d7_1580ac38 , n44374 );
buf ( R_1615_150e0598 , n44396 );
buf ( R_14c4_15ffa148 , n44397 );
buf ( R_886_156aa9b8 , C0 );
buf ( R_ff6_13d424f8 , C0 );
buf ( R_ea5_13d23b18 , n44430 );
buf ( R_1a51_13cda098 , n44435 );
buf ( R_a69_123b4f38 , n44447 );
buf ( R_1432_14b1d258 , C0 );
buf ( R_1088_13bec3f8 , n44448 );
buf ( R_e13_140ab1d8 , n44449 );
buf ( R_16a7_156afb98 , n44450 );
buf ( R_7f4_14b238d8 , n44451 );
buf ( R_17c5_12fc1058 , n44471 );
buf ( R_b87_140b0db8 , n44472 );
buf ( R_cf5_156ab818 , n44483 );
buf ( R_1933_11633258 , n44484 );
buf ( R_11a6_13c243f8 , C0 );
buf ( R_568_13ccd9d8 , n44485 );
buf ( R_6d6_13ccc498 , C0 );
buf ( R_1314_13b93158 , n44486 );
buf ( R_a81_11c6b098 , n44508 );
buf ( R_10a0_148694d8 , n44509 );
buf ( R_1a39_150e4cd8 , n44513 );
buf ( R_16bf_13d3e8f8 , n44514 );
buf ( R_141a_13ccc678 , C0 );
buf ( R_dfb_123b4c18 , n44515 );
buf ( R_7dc_14b22578 , n44516 );
buf ( R_116b_13ddcb58 , n44517 );
buf ( R_134f_14b1c7b8 , n44518 );
buf ( R_b4c_13d41eb8 , n44519 );
buf ( R_711_140b8798 , n44529 );
buf ( R_178a_13b96538 , C0 );
buf ( R_196e_150e3658 , C0 );
buf ( R_d30_13df5118 , n44530 );
buf ( R_b99_13df2ff8 , n44541 );
buf ( R_ce3_10088b58 , n44542 );
buf ( R_11b8_156b8798 , n44543 );
buf ( R_1921_13b91df8 , n44577 );
buf ( R_57a_13ccb818 , n44578 );
buf ( R_6c4_15887798 , n44579 );
buf ( R_17d7_11c6faf8 , n44580 );
buf ( R_1302_12fbe8f8 , C0 );
buf ( R_65c_117f0278 , n44581 );
buf ( R_5e2_117ef198 , C0 );
buf ( R_c01_13df0118 , n44614 );
buf ( R_18b9_13ded058 , n44623 );
buf ( R_1220_117f77f8 , n44624 );
buf ( R_129a_14a10ef8 , C0 );
buf ( R_183f_140b7f78 , n44625 );
buf ( R_c7b_1580c178 , n44626 );
buf ( R_7bd_12fc1558 , n44635 );
buf ( R_aa0_11c6be58 , n44636 );
buf ( R_10bf_13df54d8 , n44637 );
buf ( R_16de_13de3138 , C0 );
buf ( R_1a1a_156b8ab8 , C0 );
buf ( R_13fb_156b4b98 , n44638 );
buf ( R_ddc_11632df8 , n44639 );
buf ( R_a7a_11c6b1d8 , C0 );
buf ( R_1a40_140b6d58 , n44640 );
buf ( R_1099_116354b8 , n44651 );
buf ( R_1421_117ef7d8 , n44662 );
buf ( R_16b8_13d3ea38 , n44663 );
buf ( R_e02_15ff37a8 , C0 );
buf ( R_7e3_15812118 , n44664 );
buf ( R_1a56_13bf0818 , C0 );
buf ( R_1437_123bad98 , n44665 );
buf ( R_a64_13beb318 , n44666 );
buf ( R_e18_156afc38 , n44667 );
buf ( R_1083_123c0a18 , n44668 );
buf ( R_7f9_156b30b8 , n44697 );
buf ( R_16a2_150e9418 , C0 );
buf ( R_18e0_13c201b8 , n44698 );
buf ( R_1818_140b47d8 , n44699 );
buf ( R_12c1_123bb838 , n44725 );
buf ( R_5bb_156b5638 , n44726 );
buf ( R_ca2_13dd9d18 , C0 );
buf ( R_bda_13b985b8 , C0 );
buf ( R_683_11634478 , n44727 );
buf ( R_11f9_13ccd938 , n44766 );
buf ( R_157b_1486f0b8 , n44767 );
buf ( R_f5c_13de2378 , n44768 );
buf ( R_93d_117f0ef8 , n44795 );
buf ( R_920_13df90d8 , n44796 );
buf ( R_f3f_13bf1a38 , n44797 );
buf ( R_155e_123c0d38 , C0 );
buf ( R_8de_13d4e0d8 , C0 );
buf ( R_f9e_13b8a738 , C0 );
buf ( R_efd_123bfed8 , n44811 );
buf ( R_97f_123c21d8 , n44812 );
buf ( R_151c_13d5c4f8 , n44813 );
buf ( R_15bd_13df43f8 , n44836 );
buf ( R_1763_13d44618 , n44837 );
buf ( R_1995_17017548 , n44845 );
buf ( R_1144_17018948 , n44846 );
buf ( R_738_1700bce8 , n44847 );
buf ( R_b25_1162ad38 , n44863 );
buf ( R_d57_13c242b8 , n44864 );
buf ( R_1376_117f5098 , C0 );
buf ( R_9be_140aaaf8 , C0 );
buf ( R_89f_156b2ed8 , n44865 );
buf ( R_15fc_13c28db8 , n44866 );
buf ( R_ebe_13cd5c78 , C0 );
buf ( R_fdd_1162dd58 , n44877 );
buf ( R_14dd_123b8db8 , n44888 );
buf ( R_14aa_13c0f9f8 , C0 );
buf ( R_86c_13df77d8 , n44889 );
buf ( R_1010_15884278 , n44890 );
buf ( R_e8b_15880ad8 , n44891 );
buf ( R_162f_15ff7808 , n44892 );
buf ( R_9f1_123be718 , n44902 );
buf ( R_1457_13d54758 , n44903 );
buf ( R_1682_1587fb38 , C0 );
buf ( R_e38_150debf8 , n44904 );
buf ( R_a44_1580d618 , n44905 );
buf ( R_819_14873898 , n44941 );
buf ( R_1063_13cd8978 , n44942 );
buf ( R_1a4c_156b8b58 , n44943 );
buf ( R_a6e_117ec3f8 , C0 );
buf ( R_142d_14b1c998 , n44953 );
buf ( R_108d_14a0a878 , n44968 );
buf ( R_e0e_156b9f58 , C0 );
buf ( R_16ac_13bf1218 , n44969 );
buf ( R_7ef_1700c788 , n44970 );
buf ( R_1014_13c079d8 , n44971 );
buf ( R_868_1587de78 , n44972 );
buf ( R_14a6_10081998 , C0 );
buf ( R_1633_117e9ab8 , n44973 );
buf ( R_9f5_13d25c38 , n44983 );
buf ( R_e87_15ff9ce8 , n44984 );
buf ( R_1829_123b40d8 , n45020 );
buf ( R_18cf_13ded238 , n45021 );
buf ( R_5cc_156aa698 , n45022 );
buf ( R_12b0_14a177f8 , n45023 );
buf ( R_beb_13cca738 , n45024 );
buf ( R_c91_15ff1cc8 , n45033 );
buf ( R_120a_13cd9738 , C0 );
buf ( R_672_13c06fd8 , C0 );
buf ( R_779_13cd2258 , n45045 );
buf ( R_d98_13b958b8 , n45046 );
buf ( R_13b7_1700e308 , n45047 );
buf ( R_19d6_117ecfd8 , C0 );
buf ( R_1722_123b5a78 , C0 );
buf ( R_1103_117f7bb8 , n45048 );
buf ( R_ae4_11634ab8 , n45049 );
buf ( R_c57_15814f58 , n45050 );
buf ( R_638_14a151d8 , n45051 );
buf ( R_606_13d50838 , C0 );
buf ( R_c25_10083bf8 , n45073 );
buf ( R_1244_13ddb898 , n45074 );
buf ( R_1863_123b9f38 , n45075 );
buf ( R_1895_13df3a98 , n45105 );
buf ( R_1276_123bda98 , C0 );
buf ( R_1042_13cd6718 , C0 );
buf ( R_e59_1587dd38 , n45117 );
buf ( R_1661_13de0758 , n45148 );
buf ( R_83a_13d21598 , C0 );
buf ( R_a23_14869cf8 , n45149 );
buf ( R_1478_13cd7618 , n45150 );
buf ( R_668_11c6aff8 , n45151 );
buf ( R_5d6_13d24158 , C0 );
buf ( R_18c5_123b5f78 , n45183 );
buf ( R_bf5_123ba7f8 , n45209 );
buf ( R_12a6_148674f8 , C0 );
buf ( R_1214_15886cf8 , n45210 );
buf ( R_c87_13c21bf8 , n45211 );
buf ( R_1833_117f3838 , n45212 );
buf ( R_1820_14872a38 , n45213 );
buf ( R_18d8_13b8ef18 , n45214 );
buf ( R_5c3_10080778 , n45215 );
buf ( R_12b9_140abb38 , n45239 );
buf ( R_be2_13b98338 , C0 );
buf ( R_c9a_13cd1f38 , C0 );
buf ( R_1201_15ff65e8 , n45282 );
buf ( R_67b_13c02bb8 , n45283 );
buf ( R_1542_14a19cd8 , C0 );
buf ( R_1597_117ee478 , n45284 );
buf ( R_f78_156af198 , n45285 );
buf ( R_959_11631bd8 , n45291 );
buf ( R_904_13bebbd8 , n45292 );
buf ( R_f23_13c2b338 , n45293 );
buf ( R_157c_14a0eab8 , n45294 );
buf ( R_f5d_15817c58 , n45317 );
buf ( R_93e_13cd6858 , C0 );
buf ( R_91f_117f7d98 , n45318 );
buf ( R_f3e_1700a708 , C0 );
buf ( R_155d_1700fa28 , n45346 );
buf ( R_764_150dee78 , n45347 );
buf ( R_1737_13cd6538 , n45348 );
buf ( R_d83_150dc678 , n45349 );
buf ( R_1118_13cce3d8 , n45350 );
buf ( R_13a2_13df95d8 , C0 );
buf ( R_af9_14b1bc78 , n45391 );
buf ( R_19c1_15811358 , n45399 );
buf ( R_14ae_14b22438 , C0 );
buf ( R_870_158800d8 , n45400 );
buf ( R_100c_14b1bef8 , n45401 );
buf ( R_e8f_13c27cd8 , n45402 );
buf ( R_9ed_150e3a18 , n45411 );
buf ( R_162b_13d24478 , n45412 );
buf ( R_64e_12fbeb78 , C0 );
buf ( R_5f0_13d25738 , n45413 );
buf ( R_c0f_1587ef58 , n45414 );
buf ( R_122e_14a181f8 , C0 );
buf ( R_184d_1486ac98 , n45429 );
buf ( R_18ab_13bf9d78 , n45430 );
buf ( R_128c_11c6a378 , n45431 );
buf ( R_c6d_13d3be78 , n45441 );
buf ( R_d11_117f09f8 , n45450 );
buf ( R_b6b_13c0e878 , n45451 );
buf ( R_17a9_15ff62c8 , n45466 );
buf ( R_1330_1580d6b8 , n45467 );
buf ( R_6f2_123ba398 , C0 );
buf ( R_118a_13c1eef8 , C0 );
buf ( R_194f_13c0e738 , n45468 );
buf ( R_1758_14a14eb8 , n45469 );
buf ( R_19a0_13c204d8 , n45470 );
buf ( R_1139_117ef878 , n45481 );
buf ( R_743_13d5a478 , n45482 );
buf ( R_b1a_13c01038 , C0 );
buf ( R_d62_15811df8 , C0 );
buf ( R_1381_123b3a98 , n45494 );
buf ( R_e6d_123b7238 , n45550 );
buf ( R_102e_150ddd98 , C0 );
buf ( R_84e_15883418 , C0 );
buf ( R_164d_14a0c678 , n45564 );
buf ( R_148c_1580e8d8 , n45565 );
buf ( R_a0f_15ffbae8 , n45566 );
buf ( R_12ee_13d3d958 , C0 );
buf ( R_11cc_14a11a38 , n45567 );
buf ( R_ccf_15812258 , n45568 );
buf ( R_58e_150e4558 , n45569 );
buf ( R_17eb_150e6538 , n45570 );
buf ( R_190d_14b294b8 , n45600 );
buf ( R_6b0_14a172f8 , n45601 );
buf ( R_bad_15883c38 , n45637 );
buf ( R_1018_13d2a878 , n45638 );
buf ( R_864_13c09238 , n45639 );
buf ( R_14a2_13cd9e18 , C0 );
buf ( R_1637_1162fbf8 , n45640 );
buf ( R_9f9_156b7438 , n45652 );
buf ( R_e83_15886438 , n45653 );
buf ( R_1a5b_13df6158 , n45654 );
buf ( R_143c_15ff2a88 , n45655 );
buf ( R_a5f_13df1518 , n45656 );
buf ( R_e1d_13c288b8 , n45665 );
buf ( R_107e_13c1c298 , C0 );
buf ( R_7fe_117f30b8 , C0 );
buf ( R_169d_156abf98 , n45683 );
buf ( R_15b3_13cd6e98 , n45684 );
buf ( R_f07_13b953b8 , n45685 );
buf ( R_f94_13d25198 , n45686 );
buf ( R_1526_1486bf58 , C0 );
buf ( R_975_13d529f8 , n45693 );
buf ( R_8e8_117f0bd8 , n45694 );
buf ( R_78f_1162c9f8 , n45695 );
buf ( R_dae_11c6d578 , C0 );
buf ( R_13cd_14a162b8 , n45704 );
buf ( R_19ec_15814738 , n45705 );
buf ( R_170c_13ccdd98 , n45706 );
buf ( R_10ed_15882dd8 , n45721 );
buf ( R_ace_15885cb8 , C0 );
buf ( R_157d_13cd56d8 , n45728 );
buf ( R_f5e_140b53b8 , C0 );
buf ( R_93f_13d57778 , n45729 );
buf ( R_91e_15886f78 , C0 );
buf ( R_f3d_11634798 , n45748 );
buf ( R_155c_156adf78 , n45749 );
buf ( R_782_15ffd168 , C0 );
buf ( R_da1_14b290f8 , n45759 );
buf ( R_13c0_117f6b78 , n45760 );
buf ( R_19df_117eb318 , n45761 );
buf ( R_1719_13c1f8f8 , n45776 );
buf ( R_10fa_13decd38 , C0 );
buf ( R_adb_17014708 , n45777 );
buf ( R_a88_13cd40f8 , n45778 );
buf ( R_10a7_117eb1d8 , n45779 );
buf ( R_16c6_158880f8 , C0 );
buf ( R_1a32_15818018 , C0 );
buf ( R_1413_13d57ef8 , n45780 );
buf ( R_df4_17013f88 , n45781 );
buf ( R_7d5_15889098 , n45789 );
buf ( R_639_13df0cf8 , n45800 );
buf ( R_605_14b1c3f8 , n45810 );
buf ( R_c24_11632d58 , n45811 );
buf ( R_1243_158151d8 , n45812 );
buf ( R_1862_140b94b8 , C0 );
buf ( R_1896_13c0a598 , C0 );
buf ( R_1277_13c27378 , n45813 );
buf ( R_c58_13dddc38 , n45814 );
buf ( R_15a7_17013448 , n45815 );
buf ( R_1532_156b4ff8 , C0 );
buf ( R_f88_13d225d8 , n45816 );
buf ( R_969_13cce298 , n45822 );
buf ( R_8f4_156b9af8 , n45823 );
buf ( R_f13_13c2b478 , n45824 );
buf ( R_1750_14a13018 , n45825 );
buf ( R_74b_123b9998 , n45826 );
buf ( R_1131_13d21c78 , n45841 );
buf ( R_d6a_13c0c118 , C0 );
buf ( R_b12_1587bb78 , C0 );
buf ( R_1389_13c2a4d8 , n45852 );
buf ( R_19a8_124c5578 , n45853 );
buf ( R_a9e_13de43f8 , C0 );
buf ( R_10bd_1162e6b8 , n45862 );
buf ( R_16dc_14b1f058 , n45863 );
buf ( R_1a1c_13cda138 , n45864 );
buf ( R_13fd_14a0e0b8 , n45875 );
buf ( R_dde_15ffc448 , C0 );
buf ( R_7bf_123bb0b8 , n45876 );
buf ( R_1027_13c277d8 , n45877 );
buf ( R_855_14a117b8 , n45888 );
buf ( R_1493_13bee3d8 , n45889 );
buf ( R_1646_13ccbdb8 , C0 );
buf ( R_a08_15ffa5a8 , n45890 );
buf ( R_e74_123b4678 , n45891 );
buf ( R_12d0_14a11cb8 , n45892 );
buf ( R_1809_13d4f7f8 , n45933 );
buf ( R_5ac_11c6e838 , n45938 );
buf ( R_cb1_13d2c998 , n45947 );
buf ( R_bcb_1007e3d8 , n45948 );
buf ( R_692_1587be98 , C0 );
buf ( R_18ef_13d28758 , n45949 );
buf ( R_11ea_1580f238 , C0 );
buf ( R_991_1007ff58 , n45957 );
buf ( R_eeb_12fbe0d8 , n45958 );
buf ( R_150a_14a0b3b8 , C0 );
buf ( R_15cf_10085958 , n45959 );
buf ( R_fb0_117f5318 , n45960 );
buf ( R_8cc_13bf3338 , n45961 );
buf ( R_ce8_11c6a7d8 , n45962 );
buf ( R_1926_116372b8 , C0 );
buf ( R_11b3_13cd3fb8 , n45963 );
buf ( R_575_15817438 , n45964 );
buf ( R_6c9_13dee318 , n45973 );
buf ( R_1307_15ff2da8 , n45974 );
buf ( R_17d2_156b8978 , C0 );
buf ( R_b94_1587e198 , n45975 );
buf ( R_1810_117f12b8 , n45976 );
buf ( R_12c9_17017868 , n45996 );
buf ( R_5b3_123baa78 , n45997 );
buf ( R_caa_15fedbc8 , C0 );
buf ( R_bd2_1580d9d8 , C0 );
buf ( R_68b_13ddf038 , n45998 );
buf ( R_11f1_13c2a938 , n46032 );
buf ( R_18e8_123bd638 , n46033 );
buf ( R_157e_13dee278 , C0 );
buf ( R_f5f_1162d038 , n46034 );
buf ( R_940_1486f838 , n46035 );
buf ( R_91d_14b1cdf8 , n46047 );
buf ( R_f3c_148682b8 , n46048 );
buf ( R_155b_12fc0158 , n46049 );
buf ( R_14b2_15ff2628 , C0 );
buf ( R_874_123c0298 , n46050 );
buf ( R_1008_1587dc98 , n46051 );
buf ( R_e93_13cd4878 , n46052 );
buf ( R_9e9_123b4498 , n46060 );
buf ( R_1627_156b7578 , n46061 );
buf ( R_cf1_124c34f8 , n46071 );
buf ( R_192f_14a12cf8 , n46072 );
buf ( R_11aa_117e9bf8 , C0 );
buf ( R_56c_140ab598 , n46073 );
buf ( R_6d2_1162ec58 , C0 );
buf ( R_1310_13ddf538 , n46074 );
buf ( R_17c9_11638578 , n46094 );
buf ( R_b8b_13df36d8 , n46095 );
buf ( R_a91_13ccfeb8 , n46133 );
buf ( R_10b0_117ea418 , n46134 );
buf ( R_16cf_11c6b138 , n46135 );
buf ( R_1a29_13d384f8 , n46139 );
buf ( R_140a_140aa5f8 , C0 );
buf ( R_deb_140b71b8 , n46140 );
buf ( R_7cc_13cd94b8 , n46141 );
buf ( R_1a47_100862b8 , n46142 );
buf ( R_a73_123be538 , n46143 );
buf ( R_1428_13dde3b8 , n46144 );
buf ( R_1092_15ff41a8 , C0 );
buf ( R_e09_15887a18 , n46153 );
buf ( R_16b1_13c0c258 , n46161 );
buf ( R_7ea_11c6e518 , C0 );
buf ( R_e66_170138a8 , C0 );
buf ( R_1035_1162a478 , n46174 );
buf ( R_847_14a15a98 , n46175 );
buf ( R_1654_1580fff8 , n46176 );
buf ( R_1485_117f6358 , n46189 );
buf ( R_a16_14b25638 , C0 );
buf ( R_b60_13b97b18 , n46190 );
buf ( R_179e_156b3c98 , C0 );
buf ( R_133b_13ddde18 , n46191 );
buf ( R_6fd_156b8338 , n46200 );
buf ( R_117f_13cd7578 , n46201 );
buf ( R_195a_150e1218 , C0 );
buf ( R_d1c_13d3fd98 , n46202 );
buf ( R_134c_14a11ad8 , n46203 );
buf ( R_b4f_12fbee98 , n46204 );
buf ( R_70e_124c25f8 , C0 );
buf ( R_178d_11638a78 , n46247 );
buf ( R_196b_1580a918 , n46248 );
buf ( R_d2d_13cd54f8 , n46257 );
buf ( R_116e_117ebb38 , C0 );
buf ( R_5e1_14b286f8 , n46266 );
buf ( R_c00_150df558 , n46267 );
buf ( R_18ba_11638bb8 , C0 );
buf ( R_121f_13dfa1b8 , n46268 );
buf ( R_129b_13cd3298 , n46269 );
buf ( R_183e_1587c398 , C0 );
buf ( R_c7c_11c6a558 , n46270 );
buf ( R_65d_13cd74d8 , n46280 );
buf ( R_9b3_13df8138 , n46281 );
buf ( R_8aa_13dd9a98 , C0 );
buf ( R_15f1_156b5d18 , n46311 );
buf ( R_ec9_1587c1b8 , n46338 );
buf ( R_fd2_13c05098 , C0 );
buf ( R_14e8_1700a528 , n46339 );
buf ( R_11dd_14875918 , n46388 );
buf ( R_12dd_14a0e158 , n46399 );
buf ( R_17fc_11635eb8 , n46400 );
buf ( R_59f_14a14c38 , n46405 );
buf ( R_cbe_116357d8 , C0 );
buf ( R_bbe_15881438 , C0 );
buf ( R_18fc_17009bc8 , n46406 );
buf ( R_69f_13d56b98 , n46407 );
buf ( R_1598_13cd92d8 , n46408 );
buf ( R_f79_13bf2e38 , n46425 );
buf ( R_95a_13d37698 , C0 );
buf ( R_903_117ec7b8 , n46426 );
buf ( R_f22_14a13978 , C0 );
buf ( R_1541_15886758 , n46437 );
buf ( R_12e3_17014028 , n46438 );
buf ( R_11d7_1587d5b8 , n46439 );
buf ( R_cc4_13bead78 , n46440 );
buf ( R_599_150dcf38 , n46445 );
buf ( R_17f6_117f1498 , C0 );
buf ( R_1902_14b1af58 , C0 );
buf ( R_6a5_13df56b8 , n46454 );
buf ( R_bb8_124c3b38 , n46455 );
buf ( R_14bf_150dd938 , n46456 );
buf ( R_881_150db278 , n46461 );
buf ( R_ffb_15813ab8 , n46462 );
buf ( R_ea0_13b95778 , n46463 );
buf ( R_9dc_15ff19a8 , n46464 );
buf ( R_161a_14b23bf8 , C0 );
buf ( R_1454_123b4538 , n46465 );
buf ( R_e35_11c70098 , n46477 );
buf ( R_a47_1486f3d8 , n46478 );
buf ( R_816_13c06cb8 , C0 );
buf ( R_1066_13bee838 , C0 );
buf ( R_1685_15ff1d68 , n46492 );
buf ( R_8b0_15813c98 , n46493 );
buf ( R_9ad_13de0bb8 , n46501 );
buf ( R_ecf_13c26798 , n46502 );
buf ( R_15eb_140b6498 , n46503 );
buf ( R_14ee_13d5a298 , C0 );
buf ( R_fcc_150e33d8 , n46504 );
buf ( R_101c_11c6ce98 , n46505 );
buf ( R_860_14a17b18 , n46506 );
buf ( R_149e_11c6edd8 , C0 );
buf ( R_163b_13c04b98 , n46507 );
buf ( R_9fd_117ebf98 , n46525 );
buf ( R_e7f_117f6038 , n46526 );
buf ( R_604_15811718 , n46527 );
buf ( R_c23_123bfc58 , n46528 );
buf ( R_1242_10080c78 , C0 );
buf ( R_1861_12fbf7f8 , n46552 );
buf ( R_1897_13d3d1d8 , n46553 );
buf ( R_1278_117f4f58 , n46554 );
buf ( R_c59_116304b8 , n46556 );
buf ( R_63a_13c0a278 , C0 );
buf ( R_b59_15feff68 , n46599 );
buf ( R_1342_148716d8 , C0 );
buf ( R_1797_117f7e38 , n46600 );
buf ( R_704_123b2ff8 , n46601 );
buf ( R_1961_1162de98 , n46609 );
buf ( R_1178_13cd24d8 , n46610 );
buf ( R_d23_11c68618 , n46611 );
buf ( R_157f_13b8ce98 , n46612 );
buf ( R_f60_140af9b8 , n46613 );
buf ( R_941_13df8b38 , n46629 );
buf ( R_91c_13df6d38 , n46630 );
buf ( R_f3b_15810c78 , n46631 );
buf ( R_155a_15882338 , C0 );
buf ( R_e5c_117f6df8 , n46632 );
buf ( R_165e_117edf78 , C0 );
buf ( R_83d_13c24ad8 , n46665 );
buf ( R_a20_15883738 , n46666 );
buf ( R_147b_1700f5c8 , n46667 );
buf ( R_103f_123b9ad8 , n46668 );
buf ( R_5ef_1162a018 , n46669 );
buf ( R_c0e_158802b8 , C0 );
buf ( R_122d_150e4eb8 , n46680 );
buf ( R_184c_14a19418 , n46681 );
buf ( R_18ac_117f13f8 , n46682 );
buf ( R_128d_123b2af8 , n46712 );
buf ( R_c6e_15ff6408 , C0 );
buf ( R_64f_13bf1ad8 , n46713 );
buf ( R_9a0_13dd6078 , n46714 );
buf ( R_edc_123be678 , n46715 );
buf ( R_15de_15ff2268 , C0 );
buf ( R_14fb_13c29038 , n46716 );
buf ( R_fbf_150e4f58 , n46717 );
buf ( R_8bd_13cd5ef8 , n46740 );
buf ( R_1998_14b279d8 , n46741 );
buf ( R_1141_1580bbd8 , n46758 );
buf ( R_73b_14a15638 , n46759 );
buf ( R_b22_13cce8d8 , C0 );
buf ( R_d5a_13bf6178 , C0 );
buf ( R_1379_123bdbd8 , n46771 );
buf ( R_1760_117f7f78 , n46772 );
buf ( R_1981_1587b7b8 , n46780 );
buf ( R_b39_15ffae68 , n46794 );
buf ( R_724_117ec8f8 , n46795 );
buf ( R_1777_1587ccf8 , n46796 );
buf ( R_d43_13beedd8 , n46797 );
buf ( R_1362_150dfcd8 , C0 );
buf ( R_1158_13bf0f98 , n46798 );
buf ( R_770_15888058 , n46799 );
buf ( R_d8f_11629f78 , n46800 );
buf ( R_13ae_13bf3478 , C0 );
buf ( R_172b_156b88d8 , n46801 );
buf ( R_19cd_117ed578 , n46809 );
buf ( R_110c_15810458 , n46810 );
buf ( R_aed_14a0e298 , n46850 );
buf ( R_1449_14b26678 , n46860 );
buf ( R_e2a_13c29858 , C0 );
buf ( R_a52_140af378 , C0 );
buf ( R_80b_158154f8 , n46861 );
buf ( R_1071_123c1378 , n46875 );
buf ( R_1a68_117ed618 , n46876 );
buf ( R_1690_13c216f8 , n46877 );
buf ( R_ef3_13cd06d8 , n46878 );
buf ( R_989_13c068f8 , n46885 );
buf ( R_1512_1162e078 , C0 );
buf ( R_15c7_13d3c4b8 , n46886 );
buf ( R_8d4_123c1738 , n46887 );
buf ( R_fa8_123be858 , n46888 );
buf ( R_1984_1162e438 , n46889 );
buf ( R_727_1700aca8 , n46890 );
buf ( R_b36_123bb338 , C0 );
buf ( R_d46_13cd3338 , C0 );
buf ( R_1774_13c26c98 , n46891 );
buf ( R_1365_150db818 , n46902 );
buf ( R_1155_17012868 , n46912 );
buf ( R_b3c_13cd4eb8 , n46913 );
buf ( R_721_156b7d98 , n46922 );
buf ( R_197e_13d5c8b8 , C0 );
buf ( R_177a_123c1418 , C0 );
buf ( R_d40_11635af8 , n46923 );
buf ( R_115b_123bf2f8 , n46924 );
buf ( R_135f_11c6da78 , n46925 );
buf ( R_894_1587b2b8 , n46926 );
buf ( R_1607_123bd138 , n46927 );
buf ( R_eb3_123b5cf8 , n46928 );
buf ( R_fe8_15816678 , n46929 );
buf ( R_14d2_11636e58 , C0 );
buf ( R_9c9_13cce798 , n46937 );
buf ( R_160c_117f74d8 , n46938 );
buf ( R_88f_13c0d338 , n46939 );
buf ( R_fed_12fc1198 , n46945 );
buf ( R_eae_13cd1d58 , C0 );
buf ( R_9ce_1162c6d8 , C0 );
buf ( R_14cd_10081178 , n46955 );
buf ( R_dac_14a109f8 , n46956 );
buf ( R_13cb_13ccf0f8 , n46957 );
buf ( R_19ea_11629b18 , C0 );
buf ( R_170e_1580e338 , C0 );
buf ( R_10ef_14a199b8 , n46958 );
buf ( R_ad0_123b65b8 , n46959 );
buf ( R_78d_15817618 , n46971 );
buf ( R_999_1008a138 , n46979 );
buf ( R_ee3_158135b8 , n46980 );
buf ( R_1502_117ea238 , C0 );
buf ( R_15d7_11c6ab98 , n46981 );
buf ( R_fb8_156b7bb8 , n46982 );
buf ( R_8c4_117f8018 , n46983 );
buf ( R_efc_12fc14b8 , n46984 );
buf ( R_980_13d2b9f8 , n46985 );
buf ( R_151b_14a153b8 , n46986 );
buf ( R_15be_11629bb8 , C0 );
buf ( R_8dd_13d1dcb8 , n47008 );
buf ( R_f9f_13bf1858 , n47009 );
buf ( R_8a4_13cd4418 , n47010 );
buf ( R_15f7_117ea878 , n47011 );
buf ( R_ec3_14a15e58 , n47012 );
buf ( R_fd8_117f1718 , n47013 );
buf ( R_14e2_13ddc478 , C0 );
buf ( R_9b9_1008a458 , n47021 );
buf ( R_1580_123b3958 , n47022 );
buf ( R_f61_14867318 , n47049 );
buf ( R_942_140b3a18 , C0 );
buf ( R_91b_156b0d18 , n47050 );
buf ( R_f3a_1007f4b8 , C0 );
buf ( R_1559_13c234f8 , n47059 );
buf ( R_1441_13ded378 , n47070 );
buf ( R_a5a_13c097d8 , C0 );
buf ( R_e22_117eccb8 , C0 );
buf ( R_1079_13beb6d8 , n47080 );
buf ( R_803_140b8158 , n47081 );
buf ( R_1698_15811998 , n47082 );
buf ( R_1a60_14b1b778 , n47083 );
buf ( R_1987_140b7cf8 , n47084 );
buf ( R_72a_158127f8 , C0 );
buf ( R_b33_13d2aaf8 , n47085 );
buf ( R_d49_15811678 , n47094 );
buf ( R_1771_17009c68 , n47107 );
buf ( R_1368_1587e9b8 , n47108 );
buf ( R_1152_13c0bd58 , C0 );
buf ( R_5d5_123be038 , n47120 );
buf ( R_18c6_13d3a1b8 , C0 );
buf ( R_bf4_1587cb18 , n47121 );
buf ( R_12a7_15817cf8 , n47122 );
buf ( R_1213_140ad078 , n47123 );
buf ( R_c88_17017cc8 , n47124 );
buf ( R_1832_123bc2d8 , C0 );
buf ( R_669_116322b8 , n47134 );
buf ( R_769_150da558 , n47143 );
buf ( R_d88_117f22f8 , n47144 );
buf ( R_1732_123b2558 , C0 );
buf ( R_13a7_13c08ab8 , n47145 );
buf ( R_1113_123c1e18 , n47146 );
buf ( R_19c6_13cd18f8 , C0 );
buf ( R_af4_1580feb8 , n47147 );
buf ( R_b3f_13c22198 , n47148 );
buf ( R_71e_140aec98 , C0 );
buf ( R_197b_123c14b8 , n47149 );
buf ( R_177d_17012728 , n47163 );
buf ( R_d3d_13c053b8 , n47171 );
buf ( R_115e_15885c18 , C0 );
buf ( R_135c_13cda3b8 , n47172 );
buf ( R_12d7_13cd2578 , n47173 );
buf ( R_1802_13d3fbb8 , C0 );
buf ( R_5a5_13d375f8 , n47178 );
buf ( R_cb8_11c6c218 , n47179 );
buf ( R_bc4_14b2a138 , n47180 );
buf ( R_699_15888ff8 , n47191 );
buf ( R_18f6_124c27d8 , C0 );
buf ( R_11e3_1162fa18 , n47192 );
buf ( R_b67_13cd4f58 , n47193 );
buf ( R_17a5_116334d8 , n47234 );
buf ( R_1334_13cd5598 , n47235 );
buf ( R_6f6_117f1858 , C0 );
buf ( R_1186_11635d78 , C0 );
buf ( R_1953_117eb6d8 , n47236 );
buf ( R_d15_123b5578 , n47247 );
buf ( R_603_13ddbe38 , n47248 );
buf ( R_c22_117f71b8 , C0 );
buf ( R_1241_1162a5b8 , n47281 );
buf ( R_1860_13ccdf78 , n47282 );
buf ( R_1898_11c6bb38 , n47283 );
buf ( R_1279_15887478 , n47315 );
buf ( R_c5a_14a16538 , C0 );
buf ( R_63b_15883cd8 , n47316 );
buf ( R_10bb_1587d8d8 , n47317 );
buf ( R_16da_124c3db8 , C0 );
buf ( R_1a1e_11c6ed38 , C0 );
buf ( R_13ff_17012c28 , n47318 );
buf ( R_de0_13d3abb8 , n47319 );
buf ( R_7c1_156b3bf8 , n47329 );
buf ( R_a9c_1162e4d8 , n47330 );
buf ( R_18d0_117f1358 , n47331 );
buf ( R_5cb_12fc0d38 , n47332 );
buf ( R_12b1_124c38b8 , n47363 );
buf ( R_bea_13ccb098 , C0 );
buf ( R_c92_150e3838 , C0 );
buf ( R_1209_14a0aa58 , n47400 );
buf ( R_673_14a13fb8 , n47401 );
buf ( R_1828_1580ab98 , n47402 );
buf ( R_14b6_1587d1f8 , C0 );
buf ( R_878_13c100d8 , n47403 );
buf ( R_1004_156ab318 , n47404 );
buf ( R_e97_14866918 , n47405 );
buf ( R_9e5_1587d6f8 , n47414 );
buf ( R_1623_13b96178 , n47415 );
buf ( R_11d1_1162f6f8 , n47425 );
buf ( R_cca_117eebf8 , C0 );
buf ( R_593_117ee0b8 , n47430 );
buf ( R_17f0_100833d8 , n47431 );
buf ( R_1908_1162f5b8 , n47432 );
buf ( R_6ab_13ccbe58 , n47433 );
buf ( R_bb2_15810278 , C0 );
buf ( R_12e9_13d26818 , n47443 );
buf ( R_f89_13d51738 , n47461 );
buf ( R_96a_1587c258 , C0 );
buf ( R_8f3_10082b18 , n47462 );
buf ( R_f12_1162b2d8 , C0 );
buf ( R_15a8_14b25db8 , n47463 );
buf ( R_1531_13c0ac78 , n47471 );
buf ( R_12c2_13d4e2b8 , C0 );
buf ( R_5ba_13b94d78 , C0 );
buf ( R_ca3_13ddaa38 , n47472 );
buf ( R_bd9_13d54398 , n47502 );
buf ( R_684_117f5a98 , n47503 );
buf ( R_11f8_13bf1538 , n47504 );
buf ( R_18e1_17010388 , n47523 );
buf ( R_1817_1580f9b8 , n47524 );
buf ( R_a7f_117ebc78 , n47525 );
buf ( R_1a3b_13d275d8 , n47526 );
buf ( R_109e_14a11538 , C0 );
buf ( R_16bd_117eb9f8 , n47535 );
buf ( R_141c_123b3f98 , n47536 );
buf ( R_dfd_1700cf08 , n47547 );
buf ( R_7de_15881ed8 , C0 );
buf ( R_f95_13d51058 , n47553 );
buf ( R_1525_140b5598 , n47589 );
buf ( R_976_140b2f78 , C0 );
buf ( R_8e7_13dd8ff8 , n47590 );
buf ( R_15b4_13dee598 , n47591 );
buf ( R_f06_14b29238 , C0 );
buf ( R_899_13d5a8d8 , n47608 );
buf ( R_1602_13c28ef8 , C0 );
buf ( R_eb8_13c1c0b8 , n47609 );
buf ( R_fe3_13ccb598 , n47610 );
buf ( R_14d7_14a0fb98 , n47611 );
buf ( R_9c4_123c1a58 , n47612 );
buf ( R_1599_13bf40f8 , n47618 );
buf ( R_f7a_13d510f8 , C0 );
buf ( R_95b_15813838 , n47619 );
buf ( R_902_14a0aff8 , C0 );
buf ( R_f21_15812398 , n47641 );
buf ( R_1540_14871458 , n47642 );
buf ( R_1321_156b1038 , n47669 );
buf ( R_1199_13cd3bf8 , n47706 );
buf ( R_6e3_140b27f8 , n47707 );
buf ( R_55b_13d54f78 , n47708 );
buf ( R_1940_117ed758 , n47709 );
buf ( R_17b8_14b1ca38 , n47710 );
buf ( R_d02_14b21998 , C0 );
buf ( R_b7a_140b8298 , C0 );
buf ( R_ed5_123b27d8 , n47718 );
buf ( R_15e5_13d3e0d8 , n47741 );
buf ( R_14f4_1580cad8 , n47742 );
buf ( R_fc6_117f2078 , C0 );
buf ( R_8b6_12fbe7b8 , C0 );
buf ( R_9a7_13dd6118 , n47743 );
buf ( R_d96_13c23778 , C0 );
buf ( R_13b5_124c31d8 , n47755 );
buf ( R_19d4_123b6798 , n47756 );
buf ( R_1724_117edcf8 , n47757 );
buf ( R_1105_158130b8 , n47801 );
buf ( R_ae6_14873e38 , C0 );
buf ( R_777_17012228 , n47802 );
buf ( R_1581_10080458 , n47847 );
buf ( R_f62_13ccaff8 , C0 );
buf ( R_943_156b21b8 , n47848 );
buf ( R_91a_13d23e38 , C0 );
buf ( R_f39_117f5778 , n47867 );
buf ( R_1558_15ffb2c8 , n47868 );
buf ( R_88a_15880c18 , C0 );
buf ( R_ff2_13d42638 , C0 );
buf ( R_ea9_15810ef8 , n47900 );
buf ( R_9d3_12fc1e18 , n47901 );
buf ( R_14c8_13d50d38 , n47902 );
buf ( R_1611_13df2b98 , n47965 );
buf ( R_5c2_150db138 , C0 );
buf ( R_12ba_158138d8 , C0 );
buf ( R_be1_10082898 , n47995 );
buf ( R_c9b_13b977f8 , n47996 );
buf ( R_1200_13d3d778 , n47997 );
buf ( R_67c_13dec978 , n47998 );
buf ( R_181f_156b4558 , n47999 );
buf ( R_18d9_117f3e78 , n48012 );
buf ( R_1743_15ff3488 , n48013 );
buf ( R_758_13cd0ef8 , n48014 );
buf ( R_1124_14a17d98 , n48015 );
buf ( R_d77_14a0ca38 , n48016 );
buf ( R_1396_156ace98 , C0 );
buf ( R_b05_13d37d78 , n48025 );
buf ( R_19b5_13cd3c98 , n48033 );
buf ( R_d9f_1580b818 , n48034 );
buf ( R_13be_156af5f8 , C0 );
buf ( R_19dd_13d56238 , n48038 );
buf ( R_171b_14a0ac38 , n48039 );
buf ( R_10fc_13d52c78 , n48040 );
buf ( R_add_17015ce8 , n48050 );
buf ( R_780_13cd31f8 , n48051 );
buf ( R_198a_12fc1af8 , C0 );
buf ( R_72d_13d467d8 , n48064 );
buf ( R_b30_156ac358 , n48065 );
buf ( R_d4c_11633d98 , n48066 );
buf ( R_176e_12fbe678 , C0 );
buf ( R_136b_15810638 , n48067 );
buf ( R_114f_123ba1b8 , n48068 );
buf ( R_119d_123ba578 , n48077 );
buf ( R_55f_13cce658 , n48078 );
buf ( R_6df_13bf5ef8 , n48079 );
buf ( R_131d_14a11c18 , n48090 );
buf ( R_17bc_15886d98 , n48091 );
buf ( R_b7e_123b7eb8 , C0 );
buf ( R_cfe_123b7418 , C0 );
buf ( R_193c_123b6298 , n48092 );
buf ( R_b42_116296b8 , C0 );
buf ( R_71b_13cd8fb8 , n48093 );
buf ( R_1978_1587e698 , n48094 );
buf ( R_1780_1587b718 , n48095 );
buf ( R_d3a_117f6678 , C0 );
buf ( R_1161_13beb3b8 , n48105 );
buf ( R_1359_11c6d9d8 , n48116 );
buf ( R_1325_156ac178 , n48127 );
buf ( R_6e7_15882fb8 , n48128 );
buf ( R_557_15885f38 , n48129 );
buf ( R_1195_116363b8 , n48169 );
buf ( R_1944_124c2918 , n48170 );
buf ( R_d06_13dde818 , C0 );
buf ( R_b76_13d41b98 , C0 );
buf ( R_17b4_13d29ab8 , n48171 );
buf ( R_1020_117ed258 , n48172 );
buf ( R_85c_1580fc38 , n48173 );
buf ( R_149a_13bf0ef8 , C0 );
buf ( R_163f_13de4218 , n48174 );
buf ( R_a01_156b1498 , n48191 );
buf ( R_e7b_1486b738 , n48192 );
buf ( R_11c1_123b5618 , n48202 );
buf ( R_cda_156b9878 , C0 );
buf ( R_1918_15880f38 , n48203 );
buf ( R_583_13cccb78 , n48204 );
buf ( R_17e0_14a15d18 , n48205 );
buf ( R_6bb_117f2398 , n48206 );
buf ( R_ba2_14a0e5b8 , C0 );
buf ( R_12f9_13d5c9f8 , n48217 );
buf ( R_5ee_12fc0c98 , C0 );
buf ( R_c0d_13b93fb8 , n48244 );
buf ( R_122c_14b217b8 , n48245 );
buf ( R_18ad_13cd6358 , n48272 );
buf ( R_184b_1486d3f8 , n48273 );
buf ( R_128e_13b91a38 , C0 );
buf ( R_c6f_150e83d8 , n48274 );
buf ( R_650_116346f8 , n48275 );
buf ( R_5e0_13df04d8 , n48276 );
buf ( R_bff_123b92b8 , n48277 );
buf ( R_18bb_11c6f698 , n48278 );
buf ( R_121e_14b1d438 , C0 );
buf ( R_129c_1007ebf8 , n48279 );
buf ( R_183d_15882e78 , n48292 );
buf ( R_c7d_13c108f8 , n48303 );
buf ( R_65e_13d43998 , C0 );
buf ( R_75d_156ad118 , n48313 );
buf ( R_173e_148678b8 , C0 );
buf ( R_d7c_123be998 , n48314 );
buf ( R_111f_14a110d8 , n48315 );
buf ( R_139b_156b35b8 , n48316 );
buf ( R_b00_13ccf558 , n48317 );
buf ( R_19ba_17014d48 , C0 );
buf ( R_a78_13cd1cb8 , n48318 );
buf ( R_1a42_15817118 , C0 );
buf ( R_1097_13d240b8 , n48319 );
buf ( R_1423_13c05a98 , n48320 );
buf ( R_16b6_140aab98 , C0 );
buf ( R_e04_156b17b8 , n48321 );
buf ( R_7e5_14b1e798 , n48329 );
buf ( R_746_170166e8 , C0 );
buf ( R_1136_13d56558 , C0 );
buf ( R_d65_1008bb78 , n48339 );
buf ( R_b17_123bcc38 , n48340 );
buf ( R_1384_140b3298 , n48341 );
buf ( R_19a3_117eaa58 , n48342 );
buf ( R_1755_10087258 , n48351 );
buf ( R_c21_1700d4a8 , n48380 );
buf ( R_1240_11630238 , n48381 );
buf ( R_185f_13bf7118 , n48382 );
buf ( R_1899_156b1fd8 , n48392 );
buf ( R_127a_14b28298 , C0 );
buf ( R_c5b_13d26278 , n48393 );
buf ( R_63c_1587b538 , n48394 );
buf ( R_602_156afff8 , C0 );
buf ( R_753_116336b8 , n48395 );
buf ( R_1129_13ccc3f8 , n48434 );
buf ( R_d72_13b95e58 , C0 );
buf ( R_b0a_156ad438 , C0 );
buf ( R_1391_15886578 , n48445 );
buf ( R_19b0_17014a28 , n48446 );
buf ( R_1748_117eeab8 , n48447 );
buf ( R_e32_13c05c78 , C0 );
buf ( R_a4a_117e8bb8 , C0 );
buf ( R_813_11631318 , n48448 );
buf ( R_1069_116369f8 , n48459 );
buf ( R_1688_156b6a38 , n48460 );
buf ( R_1451_150e6b78 , n48471 );
buf ( R_cdf_150dfa58 , n48472 );
buf ( R_11bc_11c6a9b8 , n48473 );
buf ( R_191d_13c10678 , n48500 );
buf ( R_57e_1162f338 , n48501 );
buf ( R_6c0_13b98c98 , n48502 );
buf ( R_17db_117f6858 , n48503 );
buf ( R_12fe_116291b8 , C0 );
buf ( R_b9d_14872678 , n48542 );
buf ( R_1349_13d26db8 , n48552 );
buf ( R_b52_1162a978 , C0 );
buf ( R_1790_117e9798 , n48553 );
buf ( R_70b_17018808 , n48554 );
buf ( R_1968_13bf0318 , n48555 );
buf ( R_d2a_15fef568 , C0 );
buf ( R_1171_117f5278 , n48596 );
buf ( R_192b_11633cf8 , n48597 );
buf ( R_11ae_123bc238 , C0 );
buf ( R_570_117ec218 , n48598 );
buf ( R_6ce_13dee1d8 , C0 );
buf ( R_130c_15ff67c8 , n48599 );
buf ( R_17cd_13b91858 , n48614 );
buf ( R_b8f_14b25b38 , n48615 );
buf ( R_ced_14a0a558 , n48625 );
buf ( R_1582_150e7ed8 , C0 );
buf ( R_f63_13cca7d8 , n48626 );
buf ( R_944_13d1fab8 , n48627 );
buf ( R_919_123bdf98 , n48641 );
buf ( R_f38_13d26958 , n48642 );
buf ( R_1557_14a16c18 , n48643 );
buf ( R_10ae_123b9358 , C0 );
buf ( R_16cd_117eee78 , n48654 );
buf ( R_1a2b_140accb8 , n48655 );
buf ( R_140c_11c6f058 , n48656 );
buf ( R_ded_14a14738 , n48666 );
buf ( R_7ce_13d45d38 , C0 );
buf ( R_a8f_17014de8 , n48667 );
buf ( R_10a5_13d564b8 , n48673 );
buf ( R_16c4_1580f878 , n48674 );
buf ( R_1a34_14a19558 , n48675 );
buf ( R_1415_158165d8 , n48686 );
buf ( R_df6_156b2bb8 , C0 );
buf ( R_7d7_13c29998 , n48687 );
buf ( R_a86_123bc0f8 , C0 );
buf ( R_165b_13de0898 , n48688 );
buf ( R_840_156b26b8 , n48689 );
buf ( R_a1d_14a15778 , n48693 );
buf ( R_147e_11638078 , C0 );
buf ( R_103c_140b0ef8 , n48694 );
buf ( R_e5f_150e3d38 , n48695 );
buf ( R_11c6_13def038 , C0 );
buf ( R_cd5_13cd09f8 , n48706 );
buf ( R_588_13de09d8 , n48707 );
buf ( R_1913_13beef18 , n48708 );
buf ( R_17e5_150de518 , n48719 );
buf ( R_6b6_13d519b8 , C0 );
buf ( R_ba7_13d2ca38 , n48720 );
buf ( R_12f4_11c6ca38 , n48721 );
buf ( R_19e8_15888e18 , n48722 );
buf ( R_1710_13bf6718 , n48723 );
buf ( R_10f1_124c52f8 , n48734 );
buf ( R_ad2_156b8658 , C0 );
buf ( R_78b_1162ddf8 , n48735 );
buf ( R_daa_1008ced8 , C0 );
buf ( R_13c9_13de18d8 , n48747 );
buf ( R_11a1_117e91f8 , n48783 );
buf ( R_563_13d1ea78 , n48784 );
buf ( R_6db_13dd91d8 , n48785 );
buf ( R_1319_117f10d8 , n48796 );
buf ( R_17c0_15ff4888 , n48797 );
buf ( R_b82_13beff58 , C0 );
buf ( R_cfa_14b21ad8 , C0 );
buf ( R_1938_13df6ab8 , n48798 );
buf ( R_82a_14a0cfd8 , C0 );
buf ( R_a33_11c70278 , n48799 );
buf ( R_1468_158803f8 , n48800 );
buf ( R_1052_117f42d8 , C0 );
buf ( R_1671_13dd6898 , n48805 );
buf ( R_e49_15ff8f28 , n48814 );
buf ( R_1329_14a16ad8 , n48824 );
buf ( R_6eb_13d45b58 , n48825 );
buf ( R_1191_15881618 , n48839 );
buf ( R_1948_13c26a18 , n48840 );
buf ( R_d0a_158820b8 , C0 );
buf ( R_b72_13c103f8 , C0 );
buf ( R_17b0_13decf18 , n48841 );
buf ( R_a36_13b92438 , C0 );
buf ( R_827_123b8f98 , n48842 );
buf ( R_1055_11635738 , n48865 );
buf ( R_1465_14a18ab8 , n48877 );
buf ( R_1674_11636c78 , n48878 );
buf ( R_e46_15884098 , C0 );
buf ( R_851_11635238 , n48886 );
buf ( R_148f_13df4358 , n48887 );
buf ( R_164a_13c1e318 , C0 );
buf ( R_a0c_100899b8 , n48888 );
buf ( R_e70_117ec538 , n48889 );
buf ( R_102b_13d38d18 , n48890 );
buf ( R_198d_156b4378 , n48898 );
buf ( R_730_123bb518 , n48899 );
buf ( R_b2d_124c29b8 , n48915 );
buf ( R_d4f_13cd15d8 , n48916 );
buf ( R_176b_150e5bd8 , n48917 );
buf ( R_136e_15ff6b88 , C0 );
buf ( R_114c_140b06d8 , n48918 );
buf ( R_16f5_13d39b78 , n48932 );
buf ( R_1a03_14b23338 , n48933 );
buf ( R_10d6_150df4b8 , C0 );
buf ( R_13e4_13cd99b8 , n48934 );
buf ( R_ab7_1700b748 , n48935 );
buf ( R_dc5_15ff3f28 , n48959 );
buf ( R_7a6_150dad78 , C0 );
buf ( R_1a05_1162d498 , n48963 );
buf ( R_13e6_1486e578 , C0 );
buf ( R_dc7_13cd2398 , n48964 );
buf ( R_16f3_10088bf8 , n48965 );
buf ( R_7a8_13beac38 , n48966 );
buf ( R_10d4_13d1de98 , n48967 );
buf ( R_ab5_13df25f8 , n49003 );
buf ( R_82d_13c24b78 , n49039 );
buf ( R_a30_117ef9b8 , n49040 );
buf ( R_146b_150da9b8 , n49041 );
buf ( R_104f_170118c8 , n49042 );
buf ( R_e4c_13ddfd58 , n49043 );
buf ( R_166e_123be3f8 , C0 );
buf ( R_73e_15883878 , C0 );
buf ( R_b1f_11631098 , n49044 );
buf ( R_d5d_11636778 , n49054 );
buf ( R_137c_11634e78 , n49055 );
buf ( R_175d_13df13d8 , n49064 );
buf ( R_199b_150dc8f8 , n49065 );
buf ( R_113e_10081ad8 , C0 );
buf ( R_b45_13cce978 , n49072 );
buf ( R_718_123b4fd8 , n49073 );
buf ( R_1975_13deedb8 , n49081 );
buf ( R_1783_15817e38 , n49082 );
buf ( R_d37_13d26d18 , n49083 );
buf ( R_1164_13df29b8 , n49084 );
buf ( R_1356_15884958 , C0 );
buf ( R_16f7_140b9558 , n49085 );
buf ( R_10d8_13d55158 , n49086 );
buf ( R_ab9_14a16358 , n49113 );
buf ( R_1a01_14a0bf98 , n49118 );
buf ( R_7a4_13cca698 , n49119 );
buf ( R_13e2_13d50338 , C0 );
buf ( R_dc3_13d5b918 , n49120 );
buf ( R_1509_13c080b8 , n49128 );
buf ( R_15d0_13d5d7b8 , n49129 );
buf ( R_fb1_17011fa8 , n49142 );
buf ( R_8cb_1162afb8 , n49143 );
buf ( R_992_158117b8 , C0 );
buf ( R_eea_158843b8 , C0 );
buf ( R_1a07_15817f78 , n49144 );
buf ( R_13e8_13d57458 , n49145 );
buf ( R_dc9_13dedb98 , n49154 );
buf ( R_7aa_14a113f8 , C0 );
buf ( R_ab3_13ccea18 , n49155 );
buf ( R_16f1_13c2b298 , n49170 );
buf ( R_10d2_14a0f4b8 , C0 );
buf ( R_84a_1700eee8 , C0 );
buf ( R_1651_100849b8 , n49183 );
buf ( R_1488_15811858 , n49184 );
buf ( R_a13_117f7ed8 , n49185 );
buf ( R_e69_14b24ff8 , n49193 );
buf ( R_1032_15884638 , C0 );
buf ( R_1434_15884a98 , n49194 );
buf ( R_a67_1587c9d8 , n49195 );
buf ( R_e15_117f6538 , n49206 );
buf ( R_1086_158844f8 , C0 );
buf ( R_16a5_1587d018 , n49214 );
buf ( R_7f6_14a10318 , C0 );
buf ( R_1a53_11c70b38 , n49215 );
buf ( R_f7b_13c24f38 , n49216 );
buf ( R_95c_13b8ad78 , n49217 );
buf ( R_901_15ff0dc8 , n49223 );
buf ( R_f20_11633078 , n49224 );
buf ( R_153f_140abef8 , n49225 );
buf ( R_159a_13d58d58 , C0 );
buf ( R_1a20_117f5638 , n49226 );
buf ( R_1401_14a19918 , n49237 );
buf ( R_de2_123bef38 , C0 );
buf ( R_7c3_14a0f058 , n49238 );
buf ( R_a9a_15816f38 , C0 );
buf ( R_10b9_15ff6908 , n49244 );
buf ( R_16d8_14b209f8 , n49245 );
buf ( R_1583_13b8ba98 , n49246 );
buf ( R_f64_123b9718 , n49247 );
buf ( R_945_123bcaf8 , n49261 );
buf ( R_918_13c20ed8 , n49262 );
buf ( R_f37_158875b8 , n49263 );
buf ( R_1556_140b5db8 , C0 );
buf ( R_a39_17016d28 , n49276 );
buf ( R_824_140b4b98 , n49277 );
buf ( R_1058_13b8c7b8 , n49278 );
buf ( R_1462_13d228f8 , C0 );
buf ( R_1677_1008aef8 , n49279 );
buf ( R_e43_140ab8b8 , n49280 );
buf ( R_123f_12fc2458 , n49281 );
buf ( R_185e_100815d8 , C0 );
buf ( R_189a_15ff14a8 , C0 );
buf ( R_127b_13de1a18 , n49282 );
buf ( R_c5c_140b8518 , n49283 );
buf ( R_63d_13df0438 , n49293 );
buf ( R_601_14a12c58 , n49303 );
buf ( R_c20_1486b7d8 , n49304 );
buf ( R_15fd_156b4c38 , n49327 );
buf ( R_ebd_117f1ad8 , n49335 );
buf ( R_fde_13d429f8 , C0 );
buf ( R_14dc_13ddc5b8 , n49336 );
buf ( R_9bf_15ff2128 , n49337 );
buf ( R_89e_123bbdd8 , C0 );
buf ( R_16f9_13cd6218 , n49349 );
buf ( R_10da_14a0d4d8 , C0 );
buf ( R_abb_14b262b8 , n49350 );
buf ( R_7a2_13de1fb8 , C0 );
buf ( R_dc1_13c211f8 , n49360 );
buf ( R_13e0_1486e4d8 , n49361 );
buf ( R_19ff_123b42b8 , n49362 );
buf ( R_1739_15ff78a8 , n49365 );
buf ( R_d81_140ad4d8 , n49374 );
buf ( R_111a_13d42ef8 , C0 );
buf ( R_13a0_117f2bb8 , n49375 );
buf ( R_afb_13bf4af8 , n49376 );
buf ( R_19bf_117f5e58 , n49377 );
buf ( R_762_156b33d8 , C0 );
buf ( R_1a09_1162d358 , n49381 );
buf ( R_13ea_1580dc58 , C0 );
buf ( R_dcb_1162f798 , n49382 );
buf ( R_7ac_13c08838 , n49383 );
buf ( R_ab1_150e1b78 , n49396 );
buf ( R_10d0_150e7938 , n49397 );
buf ( R_16ef_14a136f8 , n49398 );
buf ( R_a6c_123b7378 , n49399 );
buf ( R_142f_117f79d8 , n49400 );
buf ( R_108b_156b83d8 , n49401 );
buf ( R_e10_14a0b4f8 , n49402 );
buf ( R_16aa_150e47d8 , C0 );
buf ( R_7f1_123bc378 , n49411 );
buf ( R_1a4e_123b60b8 , C0 );
buf ( R_5b2_1486f018 , n49412 );
buf ( R_cab_15fee028 , n49413 );
buf ( R_bd1_1587dfb8 , n49441 );
buf ( R_68c_123c1b98 , n49442 );
buf ( R_11f0_13cd3a18 , n49443 );
buf ( R_18e9_13b98a18 , n49474 );
buf ( R_180f_13c1cbf8 , n49475 );
buf ( R_12ca_14a13dd8 , C0 );
buf ( R_1000_13d4e858 , n49476 );
buf ( R_e9b_13cd5f98 , n49477 );
buf ( R_9e1_13bea878 , n49486 );
buf ( R_161f_10080098 , n49487 );
buf ( R_14ba_1580ba98 , C0 );
buf ( R_87c_13dee6d8 , n49488 );
buf ( R_830_1008cc58 , n49489 );
buf ( R_a2d_13d43f38 , n49494 );
buf ( R_146e_17010ba8 , C0 );
buf ( R_104c_13d1f658 , n49495 );
buf ( R_e4f_13ccef18 , n49496 );
buf ( R_166b_116345b8 , n49497 );
buf ( R_ff7_13c0cf78 , n49498 );
buf ( R_ea4_117ea738 , n49499 );
buf ( R_9d8_156b6ad8 , n49500 );
buf ( R_1616_17009da8 , C0 );
buf ( R_14c3_116384d8 , n49501 );
buf ( R_885_13de02f8 , n49506 );
buf ( R_11b7_11c6de38 , n49507 );
buf ( R_1922_13c26018 , C0 );
buf ( R_579_13d5d358 , n49508 );
buf ( R_6c5_13d59398 , n49517 );
buf ( R_17d6_11c6d258 , C0 );
buf ( R_1303_156b3d38 , n49518 );
buf ( R_b98_14b1aeb8 , n49519 );
buf ( R_ce4_117f17b8 , n49520 );
buf ( R_96b_15816c18 , n49521 );
buf ( R_8f2_158891d8 , C0 );
buf ( R_f11_124c3598 , n49527 );
buf ( R_15a9_1007e0b8 , n49558 );
buf ( R_1530_13c1c5b8 , n49559 );
buf ( R_f8a_1580da78 , C0 );
buf ( R_5ab_13d20b98 , n49564 );
buf ( R_cb2_15883eb8 , C0 );
buf ( R_bca_1162ecf8 , C0 );
buf ( R_693_1580e978 , n49565 );
buf ( R_18f0_14868178 , n49566 );
buf ( R_11e9_12fc0518 , n49577 );
buf ( R_12d1_15ff4388 , n49585 );
buf ( R_1808_117ec998 , n49586 );
buf ( R_112e_124c40d8 , C0 );
buf ( R_d6d_10080278 , n49596 );
buf ( R_b0f_150e1e98 , n49597 );
buf ( R_138c_14a12938 , n49598 );
buf ( R_19ab_1486d5d8 , n49599 );
buf ( R_174d_13c05318 , n49601 );
buf ( R_74e_117e9dd8 , C0 );
buf ( R_5d4_1587e918 , n49602 );
buf ( R_18c7_117ed7f8 , n49603 );
buf ( R_bf3_158826f8 , n49604 );
buf ( R_12a8_140b92d8 , n49605 );
buf ( R_1212_13debed8 , C0 );
buf ( R_c89_15886078 , n49614 );
buf ( R_1831_13b99eb8 , n49624 );
buf ( R_66a_117f7c58 , C0 );
buf ( R_16fb_13d39a38 , n49625 );
buf ( R_10dc_140acad8 , n49626 );
buf ( R_abd_12fbf938 , n49642 );
buf ( R_7a0_1162cef8 , n49643 );
buf ( R_dbf_13d1dd58 , n49644 );
buf ( R_13de_13bf51d8 , C0 );
buf ( R_19fd_13c22cd8 , n49648 );
buf ( R_a62_11630378 , C0 );
buf ( R_e1a_13d29f18 , C0 );
buf ( R_1081_156ae298 , n49658 );
buf ( R_7fb_13c27c38 , n49659 );
buf ( R_16a0_1007f9b8 , n49660 );
buf ( R_1a58_123b6a18 , n49661 );
buf ( R_1439_11637c18 , n49672 );
buf ( R_1511_1162c778 , n49679 );
buf ( R_15c8_10085a98 , n49680 );
buf ( R_8d3_15fefba8 , n49681 );
buf ( R_fa9_150dc218 , n49691 );
buf ( R_ef2_13d3af78 , C0 );
buf ( R_98a_11629578 , C0 );
buf ( R_151a_15ff8d48 , C0 );
buf ( R_15bf_15ff4f68 , n49692 );
buf ( R_8dc_13dd7b58 , n49693 );
buf ( R_fa0_1162a838 , n49694 );
buf ( R_efb_13ccc2b8 , n49695 );
buf ( R_981_156acad8 , n49703 );
buf ( R_133f_11636ef8 , n49704 );
buf ( R_179a_13ccf918 , C0 );
buf ( R_701_13dd6438 , n49713 );
buf ( R_195e_15817578 , C0 );
buf ( R_117b_156b5f98 , n49714 );
buf ( R_d20_1162aa18 , n49715 );
buf ( R_b5c_116370d8 , n49716 );
buf ( R_c0c_13d3f7f8 , n49717 );
buf ( R_122b_117ec498 , n49718 );
buf ( R_18ae_13d39998 , C0 );
buf ( R_184a_124c54d8 , C0 );
buf ( R_128f_123b97b8 , n49719 );
buf ( R_c70_15885998 , n49720 );
buf ( R_651_14a122f8 , n49729 );
buf ( R_5ed_13cccad8 , n49741 );
buf ( R_1a0b_1486ee38 , n49742 );
buf ( R_13ec_117f2758 , n49743 );
buf ( R_dcd_13d1e438 , n49753 );
buf ( R_7ae_13d3c058 , C0 );
buf ( R_aaf_140af698 , n49754 );
buf ( R_10ce_11637538 , C0 );
buf ( R_16ed_156af558 , n49767 );
buf ( R_a55_12fbef38 , n49784 );
buf ( R_e27_13d405b8 , n49785 );
buf ( R_1074_14b1a878 , n49786 );
buf ( R_808_13c22c38 , n49787 );
buf ( R_1693_13cd4558 , n49788 );
buf ( R_1a65_1587f8b8 , n49789 );
buf ( R_1446_1587eff8 , C0 );
buf ( R_a3c_150e6038 , n49790 );
buf ( R_821_117f1b78 , n49800 );
buf ( R_105b_13cd2f78 , n49801 );
buf ( R_145f_13b8d398 , n49802 );
buf ( R_167a_13df45d8 , C0 );
buf ( R_e40_13c26f18 , n49803 );
buf ( R_1584_1580b318 , n49804 );
buf ( R_f65_13d3b5b8 , n49828 );
buf ( R_946_14a10a98 , C0 );
buf ( R_917_117f5458 , n49829 );
buf ( R_f36_14a118f8 , C0 );
buf ( R_1555_15815638 , n49859 );
buf ( R_cd0_117f6d58 , n49860 );
buf ( R_58d_1587f3b8 , n49861 );
buf ( R_17ea_15ffadc8 , C0 );
buf ( R_190e_13bf3d38 , C0 );
buf ( R_6b1_15ffc808 , n49870 );
buf ( R_bac_13c0a098 , n49871 );
buf ( R_12ef_14b277f8 , n49872 );
buf ( R_11cb_15ff6f48 , n49873 );
buf ( R_977_1580b1d8 , n49874 );
buf ( R_8e6_1580c0d8 , C0 );
buf ( R_15b5_14866f58 , n49897 );
buf ( R_f05_123b8ef8 , n49902 );
buf ( R_f96_15885538 , C0 );
buf ( R_1524_1162d178 , n49903 );
buf ( R_11a5_156b5138 , n49914 );
buf ( R_567_13bf17b8 , n49915 );
buf ( R_6d7_12fc12d8 , n49916 );
buf ( R_1315_123b2698 , n49927 );
buf ( R_17c4_13ccc718 , n49928 );
buf ( R_b86_123b9a38 , C0 );
buf ( R_cf6_14b29738 , C0 );
buf ( R_1934_123bf7f8 , n49929 );
buf ( R_1338_116375d8 , n49930 );
buf ( R_6fa_13bec218 , C0 );
buf ( R_1182_13c1c658 , C0 );
buf ( R_1957_13d3ec18 , n49931 );
buf ( R_d19_13def3f8 , n49942 );
buf ( R_b63_15ffbb88 , n49943 );
buf ( R_17a1_117f24d8 , n49957 );
buf ( R_132d_1587ce38 , n49966 );
buf ( R_6ef_158893b8 , n49967 );
buf ( R_118d_124c3958 , n49980 );
buf ( R_194c_1587cbb8 , n49981 );
buf ( R_d0e_13c10998 , C0 );
buf ( R_b6e_117ef5f8 , C0 );
buf ( R_17ac_1486cb38 , n49982 );
buf ( R_12b2_156ab458 , C0 );
buf ( R_be9_14867638 , n50011 );
buf ( R_c93_14a12258 , n50012 );
buf ( R_1208_13bec358 , n50013 );
buf ( R_674_123c0018 , n50014 );
buf ( R_1827_13c01b78 , n50015 );
buf ( R_18d1_117e98d8 , n50026 );
buf ( R_5ca_13ccca38 , C0 );
buf ( R_16fd_13bf4378 , n50037 );
buf ( R_10de_140b68f8 , C0 );
buf ( R_abf_13befd78 , n50038 );
buf ( R_79e_15817b18 , C0 );
buf ( R_dbd_117f2b18 , n50048 );
buf ( R_13dc_13d1ce58 , n50049 );
buf ( R_19fb_150e3978 , n50050 );
buf ( R_858_150dae18 , n50051 );
buf ( R_1496_13b8b098 , C0 );
buf ( R_1643_1162c278 , n50052 );
buf ( R_a05_117f4cd8 , n50069 );
buf ( R_e77_1486b878 , n50070 );
buf ( R_1024_11635058 , n50071 );
buf ( R_733_10086998 , n50072 );
buf ( R_b2a_150dd2f8 , C0 );
buf ( R_d52_1580c498 , C0 );
buf ( R_1768_15813b58 , n50073 );
buf ( R_1371_156b10d8 , n50086 );
buf ( R_1149_156aff58 , n50132 );
buf ( R_1990_117f1df8 , n50133 );
buf ( R_185d_1162a0b8 , n50141 );
buf ( R_189b_123bccd8 , n50142 );
buf ( R_127c_1580f198 , n50143 );
buf ( R_c5d_13bf88d8 , n50153 );
buf ( R_63e_170163c8 , C0 );
buf ( R_600_150e8798 , n50154 );
buf ( R_c1f_117ebdb8 , n50155 );
buf ( R_123e_13ccb318 , C0 );
buf ( R_bfe_17018b28 , C0 );
buf ( R_18bc_123b9df8 , n50156 );
buf ( R_121d_11632718 , n50167 );
buf ( R_129d_117f6998 , n50197 );
buf ( R_183c_14b21498 , n50198 );
buf ( R_c7e_14a0d6b8 , C0 );
buf ( R_65f_14874978 , n50199 );
buf ( R_5df_13c24178 , n50200 );
buf ( R_833_117f3dd8 , n50201 );
buf ( R_a2a_14869bb8 , C0 );
buf ( R_1471_140adbb8 , n50214 );
buf ( R_1049_11636138 , n50227 );
buf ( R_e52_13d4e498 , C0 );
buf ( R_1668_13b909f8 , n50228 );
buf ( R_15df_14b24c38 , n50229 );
buf ( R_14fa_15ff7128 , C0 );
buf ( R_fc0_13beba98 , n50230 );
buf ( R_8bc_14a0e338 , n50231 );
buf ( R_9a1_123b5758 , n50239 );
buf ( R_edb_17017048 , n50240 );
buf ( R_1a0d_13ccaaf8 , n50244 );
buf ( R_13ee_13d23398 , C0 );
buf ( R_dcf_13cccfd8 , n50245 );
buf ( R_7b0_123bf4d8 , n50246 );
buf ( R_aad_14873a78 , n50259 );
buf ( R_10cc_13cd01d8 , n50260 );
buf ( R_16eb_150e81f8 , n50261 );
buf ( R_172d_13cda318 , n50266 );
buf ( R_13ac_116343d8 , n50267 );
buf ( R_110e_14a11998 , C0 );
buf ( R_19cb_13d3a758 , n50268 );
buf ( R_aef_13d50dd8 , n50269 );
buf ( R_76e_13bf8d38 , C0 );
buf ( R_d8d_13dd52b8 , n50279 );
buf ( R_715_13b94ff8 , n50290 );
buf ( R_1972_156aa918 , C0 );
buf ( R_1786_140b5778 , C0 );
buf ( R_d34_15ff3b68 , n50291 );
buf ( R_1167_1587c7f8 , n50292 );
buf ( R_1353_123c05b8 , n50293 );
buf ( R_b48_15814378 , n50294 );
buf ( R_17fb_11c6bd18 , n50295 );
buf ( R_59e_13cd0098 , n50300 );
buf ( R_cbf_15fed948 , n50301 );
buf ( R_bbd_13b8f418 , n50366 );
buf ( R_18fd_15882798 , n50393 );
buf ( R_6a0_117edbb8 , n50394 );
buf ( R_11dc_150db458 , n50395 );
buf ( R_12de_117e9658 , C0 );
buf ( R_19db_123b8458 , n50396 );
buf ( R_171d_13d45e78 , n50411 );
buf ( R_10fe_117ebd18 , C0 );
buf ( R_adf_13ccfcd8 , n50412 );
buf ( R_77e_123bcff8 , C0 );
buf ( R_d9d_12fc0298 , n50422 );
buf ( R_13bc_13c07cf8 , n50423 );
buf ( R_142a_14a0f2d8 , C0 );
buf ( R_1090_1486e7f8 , n50424 );
buf ( R_e0b_156b7758 , n50425 );
buf ( R_16af_1486be18 , n50426 );
buf ( R_7ec_123b4038 , n50427 );
buf ( R_1a49_13ccbb38 , n50431 );
buf ( R_a71_117f59f8 , n50475 );
buf ( R_15f2_13d4fe38 , C0 );
buf ( R_ec8_15883058 , n50476 );
buf ( R_fd3_10088798 , n50477 );
buf ( R_14e7_14b1ce98 , n50478 );
buf ( R_9b4_13bf5b38 , n50479 );
buf ( R_8a9_13c21298 , n50500 );
buf ( R_ece_11634bf8 , C0 );
buf ( R_15ec_13d3f4d8 , n50501 );
buf ( R_14ed_117f5f98 , n50507 );
buf ( R_fcd_1580d258 , n50519 );
buf ( R_8af_13ddfb78 , n50520 );
buf ( R_9ae_140b18f8 , C0 );
buf ( R_1501_117f0a98 , n50527 );
buf ( R_15d8_11c6ea18 , n50528 );
buf ( R_fb9_15ff0be8 , n50541 );
buf ( R_8c3_10081498 , n50542 );
buf ( R_99a_15ffaaa8 , C0 );
buf ( R_ee2_13cd1b78 , C0 );
buf ( R_1712_11637178 , C0 );
buf ( R_10f3_14a19238 , n50543 );
buf ( R_ad4_14a0a5f8 , n50544 );
buf ( R_789_140b2cf8 , n50553 );
buf ( R_da8_140b3838 , n50554 );
buf ( R_13c7_13df0ed8 , n50555 );
buf ( R_19e6_11636958 , C0 );
buf ( R_95d_117f8338 , n50561 );
buf ( R_900_140b74d8 , n50562 );
buf ( R_f1f_1587f1d8 , n50563 );
buf ( R_153e_13d410f8 , C0 );
buf ( R_159b_1162f658 , n50564 );
buf ( R_f7c_15ffc268 , n50565 );
buf ( R_cc5_13b8c858 , n50575 );
buf ( R_598_17015108 , n50580 );
buf ( R_17f5_13c1c798 , n50590 );
buf ( R_1903_1162d2b8 , n50591 );
buf ( R_6a6_15816df8 , C0 );
buf ( R_bb7_14a17a78 , n50592 );
buf ( R_12e4_13df4678 , n50593 );
buf ( R_11d6_13cccf38 , C0 );
buf ( R_a4d_14a159f8 , n50609 );
buf ( R_810_1007f918 , n50610 );
buf ( R_106c_13cd4238 , n50611 );
buf ( R_168b_13d20d78 , n50612 );
buf ( R_144e_17019028 , C0 );
buf ( R_e2f_123b83b8 , n50613 );
buf ( R_f66_1700e448 , C0 );
buf ( R_947_13cd36f8 , n50614 );
buf ( R_916_12fbefd8 , C0 );
buf ( R_f35_13dd5fd8 , n50636 );
buf ( R_1554_13c04918 , n50637 );
buf ( R_1585_117efe18 , n50648 );
buf ( R_16ff_13b95318 , n50649 );
buf ( R_10e0_1580e478 , n50650 );
buf ( R_ac1_13d23078 , n50662 );
buf ( R_79c_1162d8f8 , n50663 );
buf ( R_dbb_1580e018 , n50664 );
buf ( R_13da_123c03d8 , C0 );
buf ( R_19f9_13cd81f8 , n50668 );
buf ( R_a3f_13c012b8 , n50669 );
buf ( R_81e_140b4cd8 , C0 );
buf ( R_105e_156ba278 , C0 );
buf ( R_145c_13ddc0b8 , n50670 );
buf ( R_167d_124c5438 , n50675 );
buf ( R_e3d_15889778 , n50685 );
buf ( R_be0_117ea5f8 , n50686 );
buf ( R_c9c_13b8ed38 , n50687 );
buf ( R_11ff_14a17618 , n50688 );
buf ( R_67d_156b7398 , n50698 );
buf ( R_181e_13c04e18 , C0 );
buf ( R_18da_13cd38d8 , C0 );
buf ( R_5c1_13c0a818 , n50705 );
buf ( R_12bb_13b8a918 , n50706 );
buf ( R_ca4_156b1c18 , n50707 );
buf ( R_bd8_117e87f8 , n50708 );
buf ( R_685_13bf38d8 , n50717 );
buf ( R_11f7_10080b38 , n50718 );
buf ( R_18e2_13becfd8 , C0 );
buf ( R_1816_14b1ff58 , C0 );
buf ( R_12c3_10083478 , n50719 );
buf ( R_5b9_140b2bb8 , n50724 );
buf ( R_1630_123b9cb8 , n50725 );
buf ( R_e8a_14b1db18 , C0 );
buf ( R_9f2_10089418 , C0 );
buf ( R_14a9_156acb78 , n50736 );
buf ( R_1011_12fbe218 , n50752 );
buf ( R_86b_124c4e98 , n50753 );
buf ( R_1726_14869a78 , C0 );
buf ( R_19d2_13d533f8 , C0 );
buf ( R_1107_13df9038 , n50754 );
buf ( R_ae8_13bef5f8 , n50755 );
buf ( R_775_158109f8 , n50766 );
buf ( R_d94_12fbf6b8 , n50767 );
buf ( R_13b3_13d40158 , n50768 );
buf ( R_1658_13bf9ff8 , n50769 );
buf ( R_843_150e0458 , n50770 );
buf ( R_1481_117e8e38 , n50782 );
buf ( R_a1a_15fefd88 , C0 );
buf ( R_1039_13ddba78 , n50793 );
buf ( R_e62_13c23098 , C0 );
buf ( R_1a0f_13c24038 , n50794 );
buf ( R_13f0_11c6e338 , n50795 );
buf ( R_dd1_13de4a38 , n50805 );
buf ( R_7b2_13bf2898 , C0 );
buf ( R_aab_13c1cfb8 , n50806 );
buf ( R_10ca_1700ac08 , C0 );
buf ( R_16e9_15ff3668 , n50820 );
buf ( R_1793_150de018 , n50821 );
buf ( R_708_14a0d258 , n50822 );
buf ( R_1965_13ccb6d8 , n50830 );
buf ( R_1174_11c6c358 , n50831 );
buf ( R_d27_13dee138 , n50832 );
buf ( R_b55_15ffb0e8 , n50847 );
buf ( R_1346_13d3f2f8 , C0 );
buf ( R_e1f_123b6ab8 , n50848 );
buf ( R_107c_117f4058 , n50849 );
buf ( R_800_13d219f8 , n50850 );
buf ( R_169b_150e49b8 , n50851 );
buf ( R_1a5d_1486e398 , n50852 );
buf ( R_143e_14a19f58 , C0 );
buf ( R_a5d_15880498 , n50868 );
buf ( R_1a22_15810b38 , C0 );
buf ( R_1403_124c5398 , n50869 );
buf ( R_de4_117f6498 , n50870 );
buf ( R_7c5_15ffbe08 , n50879 );
buf ( R_a98_1486db78 , n50880 );
buf ( R_10b7_14a17578 , n50881 );
buf ( R_16d6_14a10458 , C0 );
buf ( R_1a2d_13b8fcd8 , n50886 );
buf ( R_140e_13def718 , C0 );
buf ( R_def_13d3eb78 , n50887 );
buf ( R_7d0_156b2e38 , n50888 );
buf ( R_a8d_11632678 , n50900 );
buf ( R_10ac_156b5958 , n50901 );
buf ( R_16cb_156b72f8 , n50902 );
buf ( R_1634_17018c68 , n50903 );
buf ( R_9f6_158867f8 , C0 );
buf ( R_e86_14a183d8 , C0 );
buf ( R_1015_14b1e6f8 , n50913 );
buf ( R_867_15881398 , n50914 );
buf ( R_14a5_11629ed8 , n50926 );
buf ( R_e8e_150da878 , C0 );
buf ( R_9ee_13d54618 , C0 );
buf ( R_162c_13b96c18 , n50927 );
buf ( R_14ad_12fbf618 , n50937 );
buf ( R_86f_15ff83e8 , n50938 );
buf ( R_100d_158136f8 , n50951 );
buf ( R_189c_14a10c78 , n50952 );
buf ( R_127d_11636318 , n50982 );
buf ( R_c5e_15882a18 , C0 );
buf ( R_63f_156b5b38 , n50983 );
buf ( R_5ff_13d40ab8 , n50984 );
buf ( R_c1e_14a0b958 , C0 );
buf ( R_123d_13ddd5f8 , n50994 );
buf ( R_185c_11630738 , n50995 );
buf ( R_141e_13b90818 , C0 );
buf ( R_16bb_123b7d78 , n50996 );
buf ( R_dff_117eeb58 , n50997 );
buf ( R_7e0_13dfacf8 , n50998 );
buf ( R_a7d_123b7af8 , n51041 );
buf ( R_1a3d_156b9cd8 , n51045 );
buf ( R_109c_13b98d38 , n51046 );
buf ( R_cb9_150db638 , n51057 );
buf ( R_bc3_156b6678 , n51058 );
buf ( R_69a_13b8b6d8 , C0 );
buf ( R_18f7_13b90bd8 , n51059 );
buf ( R_11e2_13d1e4d8 , C0 );
buf ( R_12d8_13d43718 , n51060 );
buf ( R_1801_13c013f8 , n51073 );
buf ( R_5a4_15ff7d08 , n51078 );
buf ( R_13a5_13d45338 , n51090 );
buf ( R_1115_11630b98 , n51102 );
buf ( R_19c4_17016fa8 , n51103 );
buf ( R_af6_117f49b8 , C0 );
buf ( R_767_117f2d98 , n51104 );
buf ( R_d86_15fef7e8 , C0 );
buf ( R_1734_1580c718 , n51105 );
buf ( R_836_123b33b8 , C0 );
buf ( R_a27_117ede38 , n51106 );
buf ( R_1474_13c042d8 , n51107 );
buf ( R_1046_123bc918 , C0 );
buf ( R_e55_124c3a98 , n51118 );
buf ( R_1665_156ac678 , n51127 );
buf ( R_122a_14a0b318 , C0 );
buf ( R_18af_11c6f7d8 , n51128 );
buf ( R_1849_140b6358 , n51140 );
buf ( R_1290_13dd8b98 , n51141 );
buf ( R_c71_14a11e98 , n51150 );
buf ( R_652_13d386d8 , C0 );
buf ( R_5ec_14868df8 , n51151 );
buf ( R_c0b_13b8c038 , n51152 );
buf ( R_574_13d4ec18 , n51153 );
buf ( R_6ca_156b3f18 , C0 );
buf ( R_1308_117f2438 , n51154 );
buf ( R_17d1_11c6fa58 , n51165 );
buf ( R_b93_15881078 , n51166 );
buf ( R_ce9_156b86f8 , n51175 );
buf ( R_1927_123bb6f8 , n51176 );
buf ( R_11b2_14a101d8 , C0 );
buf ( R_8f1_14a0fcd8 , n51196 );
buf ( R_f10_156ab778 , n51197 );
buf ( R_15aa_13c1f498 , C0 );
buf ( R_152f_158884b8 , n51198 );
buf ( R_f8b_13dda218 , n51199 );
buf ( R_96c_15ff4e28 , n51200 );
buf ( R_948_15ff1728 , n51201 );
buf ( R_915_158834b8 , n51211 );
buf ( R_f34_123bd958 , n51212 );
buf ( R_1553_1162fdd8 , n51213 );
buf ( R_1586_13cd7938 , C0 );
buf ( R_f67_156b54f8 , n51214 );
buf ( R_1701_117ee5b8 , n51224 );
buf ( R_10e2_13b97cf8 , C0 );
buf ( R_ac3_13d41ff8 , n51225 );
buf ( R_79a_13b8d758 , C0 );
buf ( R_db9_13d4e358 , n51239 );
buf ( R_13d8_13c10178 , n51240 );
buf ( R_19f7_123b4218 , n51241 );
buf ( R_ec2_156acdf8 , C0 );
buf ( R_fd9_13cd6038 , n51248 );
buf ( R_14e1_13d4fbb8 , n51260 );
buf ( R_9ba_13d3b018 , C0 );
buf ( R_8a3_117f3298 , n51261 );
buf ( R_15f8_150dd618 , n51262 );
buf ( R_b1c_10084238 , n51263 );
buf ( R_d60_1700c1e8 , n51264 );
buf ( R_137f_13d27fd8 , n51265 );
buf ( R_175a_15fedda8 , C0 );
buf ( R_199e_123b8d18 , C0 );
buf ( R_113b_11c703b8 , n51266 );
buf ( R_741_156b0278 , n51276 );
buf ( R_15e6_140b4238 , C0 );
buf ( R_14f3_10088a18 , n51277 );
buf ( R_fc7_117e8c58 , n51278 );
buf ( R_8b5_13ccefb8 , n51298 );
buf ( R_9a8_14a19af8 , n51299 );
buf ( R_ed4_150e1998 , n51300 );
buf ( R_d68_15885b78 , n51301 );
buf ( R_b14_11c6b8b8 , n51302 );
buf ( R_1387_117eaf58 , n51303 );
buf ( R_19a6_14a19738 , C0 );
buf ( R_1752_150e4738 , C0 );
buf ( R_749_123b2918 , n51312 );
buf ( R_1133_1587e378 , n51313 );
buf ( R_1417_15ff4428 , n51314 );
buf ( R_df8_15888eb8 , n51315 );
buf ( R_7d9_124c3098 , n51324 );
buf ( R_a84_13b8b778 , n51325 );
buf ( R_10a3_13c1e4f8 , n51326 );
buf ( R_1a36_14b1b318 , C0 );
buf ( R_16c2_156b1e98 , C0 );
buf ( R_1a11_123b7b98 , n51330 );
buf ( R_13f2_13de2738 , C0 );
buf ( R_dd3_14a19a58 , n51331 );
buf ( R_7b4_15885a38 , n51332 );
buf ( R_aa9_13cd5818 , n51354 );
buf ( R_10c8_14a14058 , n51355 );
buf ( R_16e7_117eea18 , n51356 );
buf ( R_b27_10087e38 , n51357 );
buf ( R_d55_117f0f98 , n51368 );
buf ( R_1765_12fbdf98 , n51381 );
buf ( R_1374_17015888 , n51382 );
buf ( R_1146_123bed58 , C0 );
buf ( R_1993_13d53b78 , n51383 );
buf ( R_736_15ff9108 , C0 );
buf ( R_56b_123b7558 , n51384 );
buf ( R_6d3_1007e1f8 , n51385 );
buf ( R_1311_10087a78 , n51396 );
buf ( R_17c8_13d50a18 , n51397 );
buf ( R_b8a_14b26858 , C0 );
buf ( R_cf2_14a17438 , C0 );
buf ( R_1930_13c083d8 , n51398 );
buf ( R_11a9_117f1038 , n51409 );
buf ( R_1638_15815818 , n51410 );
buf ( R_9fa_123b77d8 , C0 );
buf ( R_e82_13df3ef8 , C0 );
buf ( R_1019_158858f8 , n51418 );
buf ( R_863_13d47318 , n51419 );
buf ( R_14a1_117ed938 , n51431 );
buf ( R_eb2_11c6d2f8 , C0 );
buf ( R_fe9_1162ed98 , n51437 );
buf ( R_14d1_1587ae58 , n51449 );
buf ( R_9ca_1587bd58 , C0 );
buf ( R_893_13ccf238 , n51450 );
buf ( R_1608_117f45f8 , n51451 );
buf ( R_6f3_17012cc8 , n51452 );
buf ( R_1189_13de2d78 , n51493 );
buf ( R_1950_123b8098 , n51494 );
buf ( R_d12_13cd6d58 , C0 );
buf ( R_b6a_140afff8 , C0 );
buf ( R_17a8_13d3cf58 , n51495 );
buf ( R_1331_148755f8 , n51506 );
buf ( R_e9f_17016288 , n51507 );
buf ( R_9dd_156ab8b8 , n51517 );
buf ( R_161b_13d3ca58 , n51518 );
buf ( R_14be_13b98478 , C0 );
buf ( R_880_117ea2d8 , n51519 );
buf ( R_ffc_13b8acd8 , n51520 );
buf ( R_1789_13cca9b8 , n51530 );
buf ( R_196f_13bf01d8 , n51531 );
buf ( R_d31_156b13f8 , n51540 );
buf ( R_116a_13c23e58 , C0 );
buf ( R_1350_11632498 , n51541 );
buf ( R_b4b_156ad398 , n51542 );
buf ( R_712_13b90d18 , C0 );
buf ( R_e92_117f2ed8 , C0 );
buf ( R_9ea_123b7e18 , C0 );
buf ( R_1628_123b7698 , n51543 );
buf ( R_14b1_14a16e98 , n51555 );
buf ( R_873_14a14238 , n51556 );
buf ( R_1009_13b980b8 , n51566 );
buf ( R_bf2_170099e8 , C0 );
buf ( R_12a9_1162d0d8 , n51589 );
buf ( R_1211_150e5278 , n51600 );
buf ( R_c8a_150e3798 , C0 );
buf ( R_1830_13bf6358 , n51601 );
buf ( R_66b_150e1498 , n51602 );
buf ( R_5d3_158808f8 , n51603 );
buf ( R_18c8_13cd9f58 , n51604 );
buf ( R_a42_15888198 , C0 );
buf ( R_81b_12fbec18 , n51605 );
buf ( R_1061_13d3c558 , n51616 );
buf ( R_1459_17016aa8 , n51627 );
buf ( R_1680_1486aab8 , n51628 );
buf ( R_e3a_123bb798 , C0 );
buf ( R_17ef_15889958 , n51629 );
buf ( R_1909_15815e58 , n51659 );
buf ( R_6ac_12fc1918 , n51660 );
buf ( R_bb1_14874d38 , n51672 );
buf ( R_12ea_13ddf358 , C0 );
buf ( R_11d0_170096c8 , n51673 );
buf ( R_ccb_117ec038 , n51674 );
buf ( R_592_13c23958 , n51675 );
buf ( R_fee_14b29f58 , C0 );
buf ( R_ead_13c22378 , n51683 );
buf ( R_9cf_1162e118 , n51684 );
buf ( R_14cc_123c0b58 , n51685 );
buf ( R_160d_123bff78 , n51714 );
buf ( R_88e_123c0fb8 , C0 );
buf ( R_8ff_156b7c58 , n51715 );
buf ( R_f1e_15880038 , C0 );
buf ( R_153d_15811218 , n51747 );
buf ( R_159c_15815db8 , n51748 );
buf ( R_f7d_13cd0778 , n51770 );
buf ( R_95e_13b98018 , C0 );
buf ( R_189d_13cd3518 , n51780 );
buf ( R_127e_13d4f118 , C0 );
buf ( R_c5f_12fbfa78 , n51781 );
buf ( R_640_140b2258 , n51782 );
buf ( R_5fe_15888558 , C0 );
buf ( R_c1d_13dfb1f8 , n51806 );
buf ( R_123c_15fee708 , n51807 );
buf ( R_185b_14b21538 , n51808 );
buf ( R_15d1_123b63d8 , n51831 );
buf ( R_fb2_15810818 , C0 );
buf ( R_8ca_15815bd8 , C0 );
buf ( R_993_11c6b598 , n51832 );
buf ( R_ee9_1700fca8 , n51840 );
buf ( R_1508_156b7898 , n51841 );
buf ( R_121c_158871f8 , n51842 );
buf ( R_129e_13d3cb98 , C0 );
buf ( R_183b_13c20bb8 , n51843 );
buf ( R_c7f_13cd6ad8 , n51844 );
buf ( R_660_156ba458 , n51845 );
buf ( R_5de_123b7cd8 , C0 );
buf ( R_18bd_140b9878 , n51856 );
buf ( R_bfd_11c6f238 , n51882 );
buf ( R_16b4_117ead78 , n51883 );
buf ( R_e06_1580ff58 , C0 );
buf ( R_7e7_15885858 , n51884 );
buf ( R_1a44_1162c4f8 , n51885 );
buf ( R_a76_13d38638 , C0 );
buf ( R_1095_156b0ef8 , n51888 );
buf ( R_1425_13d571d8 , n51899 );
buf ( R_8e5_150db318 , n51923 );
buf ( R_15b6_1580e838 , C0 );
buf ( R_f04_15885038 , n51924 );
buf ( R_f97_1700c288 , n51925 );
buf ( R_1523_140b8e78 , n51926 );
buf ( R_978_156b6498 , n51927 );
buf ( R_914_13d54c58 , n51928 );
buf ( R_f33_13d59258 , n51929 );
buf ( R_1552_13ccfa58 , C0 );
buf ( R_1587_140aacd8 , n51930 );
buf ( R_f68_140acb78 , n51931 );
buf ( R_949_14b26a38 , n51945 );
buf ( R_15c0_158147d8 , n51946 );
buf ( R_8db_1580e158 , n51947 );
buf ( R_fa1_1162ffb8 , n51957 );
buf ( R_efa_13bf5818 , C0 );
buf ( R_982_13debcf8 , C0 );
buf ( R_1519_15813e78 , n51965 );
buf ( R_164e_117eb138 , C0 );
buf ( R_148b_15886118 , n51966 );
buf ( R_a10_13df0f78 , n51967 );
buf ( R_e6c_15ff0d28 , n51968 );
buf ( R_102f_123c08d8 , n51969 );
buf ( R_84d_15feee88 , n52025 );
buf ( R_1703_13c254d8 , n52026 );
buf ( R_10e4_158894f8 , n52027 );
buf ( R_ac5_15883558 , n52033 );
buf ( R_798_123beb78 , n52034 );
buf ( R_db7_14869938 , n52035 );
buf ( R_13d6_156ae8d8 , C0 );
buf ( R_19f5_13d2c2b8 , n52039 );
buf ( R_eb7_11c6d1b8 , n52040 );
buf ( R_fe4_12fc21d8 , n52041 );
buf ( R_14d6_1008b178 , C0 );
buf ( R_9c5_14b21d58 , n52049 );
buf ( R_898_123b5c58 , n52050 );
buf ( R_1603_14872fd8 , n52051 );
buf ( R_1714_15889638 , n52052 );
buf ( R_10f5_140b5f98 , n52068 );
buf ( R_ad6_14873258 , C0 );
buf ( R_787_14a0e838 , n52069 );
buf ( R_da6_13ddc158 , C0 );
buf ( R_13c5_15fee208 , n52081 );
buf ( R_19e4_13de3a98 , n52082 );
buf ( R_98b_13b8dcf8 , n52083 );
buf ( R_ef1_13b924d8 , n52089 );
buf ( R_8d2_156ad578 , C0 );
buf ( R_faa_156b0458 , C0 );
buf ( R_1510_13d1f0b8 , n52090 );
buf ( R_15c9_13bf0b38 , n52117 );
buf ( R_aa7_13d451f8 , n52118 );
buf ( R_7b6_14a18018 , C0 );
buf ( R_dd5_124c5258 , n52130 );
buf ( R_10c6_1700ff28 , C0 );
buf ( R_13f4_14a0b778 , n52131 );
buf ( R_16e5_13c07ed8 , n52139 );
buf ( R_1a13_117ef058 , n52140 );
buf ( R_839_14b28f18 , n52148 );
buf ( R_e58_158814d8 , n52149 );
buf ( R_a24_123b5938 , n52150 );
buf ( R_1043_14b26538 , n52151 );
buf ( R_1477_117f0098 , n52152 );
buf ( R_1662_13df1978 , C0 );
buf ( R_854_15ff3e88 , n52153 );
buf ( R_e73_14b288d8 , n52154 );
buf ( R_a09_123bb158 , n52157 );
buf ( R_1028_117f4eb8 , n52158 );
buf ( R_1492_13cd4378 , C0 );
buf ( R_1647_12fc19b8 , n52159 );
buf ( R_be8_15ffcee8 , n52160 );
buf ( R_5c9_14b27438 , n52170 );
buf ( R_675_156aec98 , n52182 );
buf ( R_c94_13b8fb98 , n52183 );
buf ( R_1207_156b81f8 , n52184 );
buf ( R_12b3_13ddf718 , n52185 );
buf ( R_1826_140b01d8 , C0 );
buf ( R_18d2_13c290d8 , C0 );
buf ( R_cac_123c1058 , n52186 );
buf ( R_5b1_13d28e38 , n52187 );
buf ( R_68d_1700f2a8 , n52199 );
buf ( R_bd0_13ccc538 , n52200 );
buf ( R_11ef_117f3d38 , n52201 );
buf ( R_12cb_123bfe38 , n52202 );
buf ( R_180e_1580c7b8 , C0 );
buf ( R_18ea_14a115d8 , C0 );
buf ( R_d75_1486bc38 , n52213 );
buf ( R_756_13b8ae18 , C0 );
buf ( R_b07_140aaa58 , n52214 );
buf ( R_1126_156aaeb8 , C0 );
buf ( R_1394_15814878 , n52215 );
buf ( R_1745_123b4cb8 , n52221 );
buf ( R_19b3_123bc558 , n52222 );
buf ( R_d7a_13b95ef8 , C0 );
buf ( R_75b_15814558 , n52223 );
buf ( R_b02_14a13f18 , C0 );
buf ( R_1121_150e9c38 , n52236 );
buf ( R_1399_158830f8 , n52247 );
buf ( R_1740_13cd6fd8 , n52248 );
buf ( R_19b8_15812c58 , n52249 );
buf ( R_c0a_14a19ff8 , C0 );
buf ( R_5eb_15feeac8 , n52250 );
buf ( R_653_123be358 , n52251 );
buf ( R_c72_13df6fb8 , C0 );
buf ( R_1229_156b7938 , n52261 );
buf ( R_1291_14a0d758 , n52289 );
buf ( R_1848_14a197d8 , n52290 );
buf ( R_18b0_15815a98 , n52291 );
buf ( R_a96_150e8478 , C0 );
buf ( R_7c7_13d45c98 , n52292 );
buf ( R_de6_13c05778 , C0 );
buf ( R_10b5_156ab6d8 , n52297 );
buf ( R_1405_14a192d8 , n52308 );
buf ( R_16d4_14868c18 , n52309 );
buf ( R_1a24_116348d8 , n52310 );
buf ( R_85f_13dd89b8 , n52311 );
buf ( R_e7e_140ad6b8 , C0 );
buf ( R_9fe_13c02d98 , C0 );
buf ( R_101d_123b5d98 , n52319 );
buf ( R_149d_156b8dd8 , n52331 );
buf ( R_163c_1486a6f8 , n52332 );
buf ( R_d9b_13d3dbd8 , n52333 );
buf ( R_77c_116359b8 , n52334 );
buf ( R_ae1_15fed768 , n52344 );
buf ( R_1100_10085818 , n52345 );
buf ( R_13ba_15881d98 , C0 );
buf ( R_171f_13bf08b8 , n52346 );
buf ( R_19d9_1700c508 , n52354 );
buf ( R_889_15ff9b08 , n52362 );
buf ( R_9d4_11c6e6f8 , n52363 );
buf ( R_ea8_13d1fe78 , n52364 );
buf ( R_ff3_117efc38 , n52365 );
buf ( R_14c7_140b4918 , n52366 );
buf ( R_1612_13cd0278 , C0 );
buf ( R_582_14869118 , n52367 );
buf ( R_cdb_14a0ae18 , n52368 );
buf ( R_ba1_13d29338 , n52380 );
buf ( R_6bc_13cd53b8 , n52381 );
buf ( R_11c0_13deef98 , n52382 );
buf ( R_12fa_11631638 , C0 );
buf ( R_17df_13cd0e58 , n52383 );
buf ( R_1919_1587e2d8 , n52414 );
buf ( R_e24_13ddcfb8 , n52415 );
buf ( R_a58_14a18a18 , n52416 );
buf ( R_805_1580a7d8 , n52449 );
buf ( R_1077_11c6d898 , n52450 );
buf ( R_1443_13d3f9d8 , n52451 );
buf ( R_1696_156afd78 , C0 );
buf ( R_1a62_14b1b138 , C0 );
buf ( R_94a_156b24d8 , C0 );
buf ( R_f32_116350f8 , C0 );
buf ( R_913_100840f8 , n52452 );
buf ( R_f69_117f0c78 , n52478 );
buf ( R_1551_150dde38 , n52487 );
buf ( R_1588_150e7d98 , n52488 );
buf ( R_a50_13df7698 , n52489 );
buf ( R_e2c_15881e38 , n52490 );
buf ( R_80d_14a16a38 , n52525 );
buf ( R_106f_156ad938 , n52526 );
buf ( R_144b_1486ce58 , n52527 );
buf ( R_168e_123bbc98 , C0 );
buf ( R_6fe_13bf5318 , C0 );
buf ( R_b5f_13cd4918 , n52528 );
buf ( R_d1d_13def2b8 , n52537 );
buf ( R_117e_14a0ccb8 , C0 );
buf ( R_133c_117f2938 , n52538 );
buf ( R_179d_10085138 , n52579 );
buf ( R_195b_14b1c8f8 , n52580 );
buf ( R_cb3_1587b358 , n52581 );
buf ( R_5aa_13dd5678 , n52586 );
buf ( R_694_11636b38 , n52587 );
buf ( R_bc9_124c3d18 , n52606 );
buf ( R_11e8_13ccd258 , n52607 );
buf ( R_12d2_123bdc78 , C0 );
buf ( R_1807_117ee298 , n52608 );
buf ( R_18f1_156aba98 , n52637 );
buf ( R_c1c_156ba3b8 , n52638 );
buf ( R_5fd_14a10958 , n52647 );
buf ( R_641_123b90d8 , n52656 );
buf ( R_c60_158171b8 , n52657 );
buf ( R_123b_1162cd18 , n52658 );
buf ( R_127f_13b8a558 , n52659 );
buf ( R_185a_15814cd8 , C0 );
buf ( R_189e_13bf8e78 , C0 );
buf ( R_877_13d3e498 , n52660 );
buf ( R_9e6_14b28838 , C0 );
buf ( R_e96_156b4a58 , C0 );
buf ( R_1005_13c1edb8 , n52672 );
buf ( R_14b5_15882018 , n52684 );
buf ( R_1624_10086cb8 , n52685 );
buf ( R_db5_117ece98 , n52696 );
buf ( R_796_156b0138 , C0 );
buf ( R_ac7_148725d8 , n52697 );
buf ( R_10e6_11630918 , C0 );
buf ( R_13d4_15882bf8 , n52698 );
buf ( R_1705_10085db8 , n52708 );
buf ( R_19f3_1008c618 , n52709 );
buf ( R_96d_1162e7f8 , n52716 );
buf ( R_f0f_13d3d9f8 , n52717 );
buf ( R_8f0_13d29838 , n52718 );
buf ( R_f8c_117f2578 , n52719 );
buf ( R_152e_117f3f18 , C0 );
buf ( R_15ab_13ccc358 , n52720 );
buf ( R_587_124c5118 , n52721 );
buf ( R_cd6_13d39178 , C0 );
buf ( R_ba6_156ad9d8 , C0 );
buf ( R_6b7_13c0b718 , n52722 );
buf ( R_11c5_13d39538 , n52731 );
buf ( R_12f5_158104f8 , n52742 );
buf ( R_17e4_156acf38 , n52743 );
buf ( R_1914_10084f58 , n52744 );
buf ( R_846_100885b8 , C0 );
buf ( R_e65_15810318 , n52752 );
buf ( R_a17_13ccf878 , n52753 );
buf ( R_1036_140b5278 , C0 );
buf ( R_1484_11c6b778 , n52754 );
buf ( R_1655_1700cdc8 , n52763 );
buf ( R_a45_17017188 , n52770 );
buf ( R_e37_10083018 , n52771 );
buf ( R_818_13b8dbb8 , n52772 );
buf ( R_1064_1700d5e8 , n52773 );
buf ( R_1456_13cd8518 , C0 );
buf ( R_1683_1587f6d8 , n52774 );
buf ( R_57d_14b1ef18 , n52775 );
buf ( R_ce0_1580ccb8 , n52776 );
buf ( R_b9c_15884e58 , n52777 );
buf ( R_6c1_156b1538 , n52786 );
buf ( R_11bb_117ed2f8 , n52787 );
buf ( R_12ff_17012408 , n52788 );
buf ( R_17da_123bf398 , C0 );
buf ( R_191e_140b0c78 , C0 );
buf ( R_d58_13df39f8 , n52789 );
buf ( R_b24_15815958 , n52790 );
buf ( R_739_123c1698 , n52801 );
buf ( R_1143_13cd7078 , n52802 );
buf ( R_1377_158873d8 , n52803 );
buf ( R_1762_140aef18 , C0 );
buf ( R_1996_156b4058 , C0 );
buf ( R_95f_13bf9918 , n52804 );
buf ( R_f1d_15ff80c8 , n52820 );
buf ( R_8fe_13d4f898 , C0 );
buf ( R_f7e_156b42d8 , C0 );
buf ( R_153c_13c1d698 , n52821 );
buf ( R_159d_1162b198 , n52826 );
buf ( R_aa5_156b4238 , n52840 );
buf ( R_7b8_1162e9d8 , n52841 );
buf ( R_dd7_140b62b8 , n52842 );
buf ( R_10c4_12fc1878 , n52843 );
buf ( R_13f6_1700d728 , C0 );
buf ( R_16e3_123b4d58 , n52844 );
buf ( R_1a15_13d3e998 , n52849 );
buf ( R_b0c_123c1878 , n52850 );
buf ( R_d70_13b96038 , n52851 );
buf ( R_751_13bf12b8 , n52860 );
buf ( R_112b_13d5c3b8 , n52861 );
buf ( R_138f_13df66f8 , n52862 );
buf ( R_174a_13d24658 , C0 );
buf ( R_19ae_1587f818 , C0 );
buf ( R_a8b_117f7898 , n52863 );
buf ( R_7d2_10082a78 , C0 );
buf ( R_df1_15884778 , n52873 );
buf ( R_10aa_13c28458 , C0 );
buf ( R_1410_13cd5a98 , n52874 );
buf ( R_16c9_13c03018 , n52885 );
buf ( R_1a2f_15886b18 , n52886 );
buf ( R_d7f_117f5ef8 , n52887 );
buf ( R_760_13cce6f8 , n52888 );
buf ( R_afd_156ae018 , n52901 );
buf ( R_111c_13c0f138 , n52902 );
buf ( R_139e_15ff9428 , C0 );
buf ( R_173b_13d23758 , n52903 );
buf ( R_19bd_150e0c78 , n52911 );
buf ( R_70f_14b26038 , n52912 );
buf ( R_b4e_158835f8 , C0 );
buf ( R_d2e_15ff2d08 , C0 );
buf ( R_116d_14a0bc78 , n52926 );
buf ( R_134d_13cd26b8 , n52935 );
buf ( R_178c_13d39718 , n52936 );
buf ( R_196c_117ef418 , n52937 );
buf ( R_705_17018768 , n52947 );
buf ( R_b58_12fc00b8 , n52948 );
buf ( R_d24_13c0ca78 , n52949 );
buf ( R_1177_13d5b558 , n52950 );
buf ( R_1343_13d298d8 , n52951 );
buf ( R_1796_156ae338 , C0 );
buf ( R_1962_13d5d218 , C0 );
buf ( R_c9d_13c00ef8 , n52961 );
buf ( R_bdf_117f0638 , n52962 );
buf ( R_5c0_117ea0f8 , n52963 );
buf ( R_67e_14a0b8b8 , C0 );
buf ( R_11fe_124c36d8 , C0 );
buf ( R_12bc_13b981f8 , n52964 );
buf ( R_181d_123ba758 , n52978 );
buf ( R_18db_11c6d7f8 , n52979 );
buf ( R_ebc_1580cfd8 , n52980 );
buf ( R_89d_11c693d8 , n53000 );
buf ( R_9c0_13d46b98 , n53001 );
buf ( R_fdf_158176b8 , n53002 );
buf ( R_14db_156b5e58 , n53003 );
buf ( R_15fe_140b97d8 , C0 );
buf ( R_ee1_13d40c98 , n53013 );
buf ( R_99b_156b3838 , n53014 );
buf ( R_8c2_15813518 , C0 );
buf ( R_fba_140aebf8 , C0 );
buf ( R_1500_1700e8a8 , n53015 );
buf ( R_15d9_13d53538 , n53039 );
buf ( R_eda_13d57638 , C0 );
buf ( R_9a2_13c28bd8 , C0 );
buf ( R_8bb_13d43498 , n53040 );
buf ( R_fc1_156b40f8 , n53053 );
buf ( R_14f9_13cd6178 , n53060 );
buf ( R_15e0_13cd0458 , n53061 );
buf ( R_d8b_150dc7b8 , n53062 );
buf ( R_76c_150e63f8 , n53063 );
buf ( R_af1_13b8c3f8 , n53076 );
buf ( R_1110_13d5cdb8 , n53077 );
buf ( R_13aa_14b1d898 , C0 );
buf ( R_172f_11c6dbb8 , n53078 );
buf ( R_19c9_1509b4f8 , n53086 );
buf ( R_55a_158145f8 , n53087 );
buf ( R_6e4_11630a58 , n53088 );
buf ( R_b79_13ccfd78 , n53100 );
buf ( R_d03_124c2eb8 , n53101 );
buf ( R_1198_117f3b58 , n53102 );
buf ( R_1322_15ff6ea8 , C0 );
buf ( R_17b7_15810bd8 , n53103 );
buf ( R_1941_117ed4d8 , n53129 );
buf ( R_6cf_1486c6d8 , n53130 );
buf ( R_56f_14a0b598 , n53131 );
buf ( R_cee_13cd9c38 , C0 );
buf ( R_b8e_150e97d8 , C0 );
buf ( R_11ad_13d569b8 , n53148 );
buf ( R_130d_124c3818 , n53157 );
buf ( R_17cc_117e9298 , n53158 );
buf ( R_192c_13b94918 , n53159 );
buf ( R_94b_100881f8 , n53160 );
buf ( R_f31_13c231d8 , n53178 );
buf ( R_912_11630f58 , C0 );
buf ( R_f6a_117ea058 , C0 );
buf ( R_1550_17014668 , n53179 );
buf ( R_1589_123b7198 , n53185 );
buf ( R_bd7_14a0ef18 , n53186 );
buf ( R_ca5_1007eb58 , n53195 );
buf ( R_5b8_170170e8 , n53196 );
buf ( R_686_15810f98 , C0 );
buf ( R_11f6_14b22bb8 , C0 );
buf ( R_12c4_15ff0008 , n53197 );
buf ( R_1815_156b1cb8 , n53210 );
buf ( R_18e3_13ccb9f8 , n53211 );
buf ( R_6e0_14a15f98 , n53212 );
buf ( R_55e_148707d8 , n53213 );
buf ( R_cff_14a0b458 , n53214 );
buf ( R_b7d_156b6df8 , n53225 );
buf ( R_119c_14872ad8 , n53226 );
buf ( R_131e_13dd6e38 , C0 );
buf ( R_17bb_13bf1d58 , n53227 );
buf ( R_193d_11c70638 , n53253 );
buf ( R_d92_14b21358 , C0 );
buf ( R_773_117f54f8 , n53254 );
buf ( R_aea_17012908 , C0 );
buf ( R_1109_15ff3de8 , n53268 );
buf ( R_13b1_150dc358 , n53280 );
buf ( R_1728_13d5beb8 , n53281 );
buf ( R_19d0_14870af8 , n53282 );
buf ( R_e12_13b8cc18 , C0 );
buf ( R_a6a_13d1d218 , C0 );
buf ( R_7f3_148688f8 , n53283 );
buf ( R_1089_123b6838 , n53292 );
buf ( R_1431_15812ed8 , n53303 );
buf ( R_16a8_123bf118 , n53304 );
buf ( R_1a50_117ed6b8 , n53305 );
buf ( R_6f7_117e93d8 , n53306 );
buf ( R_b66_14a0f238 , C0 );
buf ( R_d16_13c1b7f8 , C0 );
buf ( R_1185_13d1ecf8 , n53319 );
buf ( R_1335_13bf1f38 , n53330 );
buf ( R_17a4_14b1ea18 , n53331 );
buf ( R_1954_15ff1ae8 , n53332 );
buf ( R_e17_13df86d8 , n53333 );
buf ( R_a65_14b22b18 , n53373 );
buf ( R_7f8_1700bec8 , n53374 );
buf ( R_1084_13d39038 , n53375 );
buf ( R_1436_15fef608 , C0 );
buf ( R_16a3_15ff2768 , n53376 );
buf ( R_1a55_123b5898 , n53380 );
buf ( R_a21_1587bad8 , n53383 );
buf ( R_83c_13cd7398 , n53384 );
buf ( R_e5b_123bf898 , n53385 );
buf ( R_1040_1008ac78 , n53386 );
buf ( R_147a_13c04378 , C0 );
buf ( R_165f_13cd97d8 , n53387 );
buf ( R_bfc_13d53cb8 , n53388 );
buf ( R_5dd_123b45d8 , n53397 );
buf ( R_661_13d3c2d8 , n53407 );
buf ( R_c80_1008ca78 , n53408 );
buf ( R_121b_14b24698 , n53409 );
buf ( R_129f_1008b7b8 , n53410 );
buf ( R_183a_156acc18 , C0 );
buf ( R_18be_14a0de38 , C0 );
buf ( R_c1b_123b48f8 , n53411 );
buf ( R_5fc_140b3518 , n53412 );
buf ( R_642_14a0d118 , C0 );
buf ( R_c61_13c06718 , n53421 );
buf ( R_123a_15ffcf88 , C0 );
buf ( R_1280_14a106d8 , n53422 );
buf ( R_1859_13d25378 , n53433 );
buf ( R_189f_14a13c98 , n53434 );
buf ( R_556_13d2a2d8 , n53435 );
buf ( R_6e8_12fbf4d8 , n53436 );
buf ( R_b75_156ae838 , n53446 );
buf ( R_d07_156abe58 , n53447 );
buf ( R_1194_1580f058 , n53448 );
buf ( R_1326_11c684d8 , C0 );
buf ( R_17b3_13ddb4d8 , n53449 );
buf ( R_1945_14b22898 , n53474 );
buf ( R_bf1_13df18d8 , n53505 );
buf ( R_5d2_10088f18 , C0 );
buf ( R_66c_123c06f8 , n53506 );
buf ( R_c8b_13c0e5f8 , n53507 );
buf ( R_1210_117f56d8 , n53508 );
buf ( R_12aa_140afb98 , C0 );
buf ( R_182f_13d58998 , n53509 );
buf ( R_18c9_11c6eb58 , n53520 );
buf ( R_cc0_1580fcd8 , n53521 );
buf ( R_59d_13df9d58 , n53526 );
buf ( R_6a1_13cd9b98 , n53535 );
buf ( R_bbc_13d4e678 , n53536 );
buf ( R_11db_124c45d8 , n53537 );
buf ( R_12df_13d27178 , n53538 );
buf ( R_17fa_13beb8b8 , C0 );
buf ( R_18fe_1587ca78 , C0 );
buf ( R_d63_117f68f8 , n53539 );
buf ( R_b19_158882d8 , n53550 );
buf ( R_744_123bea38 , n53551 );
buf ( R_1138_14869ed8 , n53552 );
buf ( R_1382_13b8b958 , C0 );
buf ( R_1757_13de1978 , n53553 );
buf ( R_19a1_123b3598 , n53561 );
buf ( R_db3_14869898 , n53562 );
buf ( R_794_17016788 , n53563 );
buf ( R_ac9_15811cb8 , n53572 );
buf ( R_10e8_140b1538 , n53573 );
buf ( R_13d2_13c292b8 , C0 );
buf ( R_1707_13ddd9b8 , n53574 );
buf ( R_19f1_13cce518 , n53578 );
buf ( R_ecd_13d5b5f8 , n53586 );
buf ( R_9af_1587fdb8 , n53587 );
buf ( R_8ae_11631778 , C0 );
buf ( R_fce_13c051d8 , C0 );
buf ( R_14ec_156b01d8 , n53588 );
buf ( R_15ed_1008af98 , n53612 );
buf ( R_da4_13cd7438 , n53613 );
buf ( R_785_116381b8 , n53622 );
buf ( R_ad8_117f7a78 , n53623 );
buf ( R_10f7_1587f598 , n53624 );
buf ( R_13c3_13cd0b38 , n53625 );
buf ( R_1716_123b6bf8 , C0 );
buf ( R_19e2_13d567d8 , C0 );
buf ( R_58c_1587fe58 , n53626 );
buf ( R_cd1_1486dc18 , n53636 );
buf ( R_bab_13df0e38 , n53637 );
buf ( R_6b2_14867ef8 , C0 );
buf ( R_11ca_123bd9f8 , C0 );
buf ( R_12f0_158817f8 , n53638 );
buf ( R_17e9_123bb5b8 , n53648 );
buf ( R_190f_15881b18 , n53649 );
buf ( R_979_117efcd8 , n53653 );
buf ( R_f03_13c06f38 , n53654 );
buf ( R_8e4_123b2b98 , n53655 );
buf ( R_f98_13d588f8 , n53656 );
buf ( R_1522_15817d98 , C0 );
buf ( R_15b7_11636bd8 , n53657 );
buf ( R_c09_14a18bf8 , n53687 );
buf ( R_5ea_1162b558 , C0 );
buf ( R_654_150e54f8 , n53688 );
buf ( R_c73_15810958 , n53689 );
buf ( R_1228_150e4ff8 , n53690 );
buf ( R_1292_117e9fb8 , C0 );
buf ( R_1847_13d54898 , n53691 );
buf ( R_18b1_1162ae78 , n53697 );
buf ( R_ec7_10083838 , n53698 );
buf ( R_8a8_140b6858 , n53699 );
buf ( R_9b5_156b6038 , n53707 );
buf ( R_fd4_13bef878 , n53708 );
buf ( R_14e6_123be178 , C0 );
buf ( R_15f3_1580b958 , n53709 );
buf ( R_6dc_13d56738 , n53710 );
buf ( R_562_11630198 , n53711 );
buf ( R_cfb_156b77f8 , n53712 );
buf ( R_b81_14b23658 , n53724 );
buf ( R_11a0_117f1a38 , n53725 );
buf ( R_131a_13cd6678 , C0 );
buf ( R_17bf_1162eed8 , n53726 );
buf ( R_1939_13b99198 , n53754 );
buf ( R_85b_150e9ff8 , n53755 );
buf ( R_e7a_13df06b8 , C0 );
buf ( R_a02_13d20378 , C0 );
buf ( R_1021_14873438 , n53763 );
buf ( R_1499_13c056d8 , n53774 );
buf ( R_1640_15816e98 , n53775 );
buf ( R_6c6_14b27a78 , C0 );
buf ( R_578_13c06678 , n53776 );
buf ( R_ce5_117e9518 , n53786 );
buf ( R_b97_116328f8 , n53787 );
buf ( R_11b6_123b6478 , C0 );
buf ( R_1304_150e5a98 , n53788 );
buf ( R_17d5_13cd9eb8 , n53836 );
buf ( R_1923_10086ad8 , n53837 );
buf ( R_aa3_123ba9d8 , n53838 );
buf ( R_7ba_17013308 , C0 );
buf ( R_dd9_1587f4f8 , n53849 );
buf ( R_10c2_13de4358 , C0 );
buf ( R_13f8_14866c38 , n53850 );
buf ( R_16e1_1587e058 , n53867 );
buf ( R_1a17_13d3a398 , n53868 );
buf ( R_ea3_117f04f8 , n53869 );
buf ( R_884_124c4358 , n53870 );
buf ( R_9d9_14a0c178 , n53881 );
buf ( R_ff8_14a15098 , n53882 );
buf ( R_14c2_13d50e78 , C0 );
buf ( R_1617_13de3e58 , n53883 );
buf ( R_e0d_13c081f8 , n53893 );
buf ( R_a6f_140ab4f8 , n53894 );
buf ( R_7ee_117eb4f8 , C0 );
buf ( R_108e_117ecf38 , C0 );
buf ( R_142c_13d55f18 , n53895 );
buf ( R_16ad_15885df8 , n53903 );
buf ( R_1a4b_13d3a118 , n53904 );
buf ( R_e01_13b8ca38 , n53913 );
buf ( R_a7b_150e6f38 , n53914 );
buf ( R_7e2_116332f8 , C0 );
buf ( R_109a_140adc58 , C0 );
buf ( R_1420_1580acd8 , n53915 );
buf ( R_16b9_13b972f8 , n53923 );
buf ( R_1a3f_13cd8f18 , n53924 );
buf ( R_597_156aeab8 , n53929 );
buf ( R_cc6_1486fd38 , C0 );
buf ( R_bb6_13d58fd8 , C0 );
buf ( R_6a7_140b7938 , n53930 );
buf ( R_11d5_14871bd8 , n53956 );
buf ( R_12e5_14b28bf8 , n53958 );
buf ( R_17f4_156b4cd8 , n53959 );
buf ( R_1904_140b9058 , n53960 );
buf ( R_dfa_1486ff18 , C0 );
buf ( R_a82_116368b8 , C0 );
buf ( R_7db_150dd1b8 , n53961 );
buf ( R_10a1_123b8598 , n53974 );
buf ( R_1419_13df1b58 , n53985 );
buf ( R_16c0_13b994b8 , n53986 );
buf ( R_1a38_13ccab98 , n53987 );
buf ( R_911_14b22078 , n53996 );
buf ( R_94c_123bc7d8 , n53997 );
buf ( R_f30_12fbf898 , n53998 );
buf ( R_f6b_13c0a6d8 , n53999 );
buf ( R_154f_1700ea88 , n54000 );
buf ( R_158a_13c25758 , C0 );
buf ( R_d44_13b99418 , n54001 );
buf ( R_b38_13d23618 , n54002 );
buf ( R_725_13d4f618 , n54012 );
buf ( R_1157_14a13298 , n54013 );
buf ( R_1363_124c4718 , n54014 );
buf ( R_1776_15882518 , C0 );
buf ( R_1982_15816fd8 , C0 );
buf ( R_983_1700b4c8 , n54015 );
buf ( R_ef9_1007e338 , n54021 );
buf ( R_8da_1587ba38 , C0 );
buf ( R_fa2_15ffaf08 , C0 );
buf ( R_1518_13c09ff8 , n54022 );
buf ( R_15c1_13c1e138 , n54048 );
buf ( R_d41_13bf8f18 , n54058 );
buf ( R_722_14b26fd8 , C0 );
buf ( R_b3b_14a0f378 , n54059 );
buf ( R_115a_156af9b8 , C0 );
buf ( R_1360_156aa5f8 , n54060 );
buf ( R_1779_13dec3d8 , n54072 );
buf ( R_197f_1700ba68 , n54073 );
buf ( R_7fd_13d29658 , n54099 );
buf ( R_e1c_156b8158 , n54100 );
buf ( R_a60_124c2738 , n54101 );
buf ( R_107f_13d55ab8 , n54102 );
buf ( R_143b_13cd5458 , n54103 );
buf ( R_169e_13d59618 , C0 );
buf ( R_1a5a_117ecd58 , C0 );
buf ( R_a94_158121b8 , n54104 );
buf ( R_7c9_13c1bb18 , n54113 );
buf ( R_de8_13df22d8 , n54114 );
buf ( R_10b3_17011328 , n54115 );
buf ( R_1407_140b9cd8 , n54116 );
buf ( R_16d2_150e0098 , C0 );
buf ( R_1a26_14868678 , C0 );
buf ( R_e9a_14a0e1f8 , C0 );
buf ( R_87b_123b2e18 , n54117 );
buf ( R_9e2_148680d8 , C0 );
buf ( R_1001_100877f8 , n54129 );
buf ( R_14b9_150dda78 , n54140 );
buf ( R_1620_117efff8 , n54141 );
buf ( R_bc2_1580b098 , C0 );
buf ( R_cba_13c20118 , C0 );
buf ( R_5a3_13b98298 , n54146 );
buf ( R_69b_13bf94b8 , n54147 );
buf ( R_11e1_1486a798 , n54160 );
buf ( R_12d9_123ba118 , n54168 );
buf ( R_1800_15888378 , n54169 );
buf ( R_18f8_156ac538 , n54170 );
buf ( R_960_13ccf418 , n54171 );
buf ( R_f1c_13df79b8 , n54172 );
buf ( R_8fd_123b6fb8 , n54191 );
buf ( R_f7f_140aa558 , n54192 );
buf ( R_153b_117f5d18 , n54193 );
buf ( R_159e_14871db8 , C0 );
buf ( R_d47_13d27998 , n54194 );
buf ( R_b35_1587cc58 , n54206 );
buf ( R_728_140ba318 , n54207 );
buf ( R_1154_117e95b8 , n54208 );
buf ( R_1366_17015568 , C0 );
buf ( R_1773_156ac2b8 , n54209 );
buf ( R_1985_1162c3b8 , n54217 );
buf ( R_b11_15883698 , n54228 );
buf ( R_d6b_123b8958 , n54229 );
buf ( R_74c_150e17b8 , n54230 );
buf ( R_1130_13bef0f8 , n54231 );
buf ( R_138a_13d25cd8 , C0 );
buf ( R_174f_13df2058 , n54232 );
buf ( R_19a9_1486eed8 , n54240 );
buf ( R_6ec_13c03b58 , n54241 );
buf ( R_b71_140afd78 , n54252 );
buf ( R_d0b_1587d158 , n54253 );
buf ( R_1190_13c09198 , n54254 );
buf ( R_132a_13d44bb8 , C0 );
buf ( R_17af_123b9d58 , n54255 );
buf ( R_1949_140b51d8 , n54284 );
buf ( R_815_158140f8 , n54317 );
buf ( R_a48_13bed6b8 , n54318 );
buf ( R_e34_13cd7e38 , n54319 );
buf ( R_1067_13b93ab8 , n54320 );
buf ( R_1453_15ff99c8 , n54321 );
buf ( R_1686_1008c258 , C0 );
buf ( R_af8_148696b8 , n54322 );
buf ( R_d84_156b3e78 , n54323 );
buf ( R_765_13df9678 , n54332 );
buf ( R_1117_140b2398 , n54333 );
buf ( R_13a3_123bd598 , n54334 );
buf ( R_1736_117f1218 , C0 );
buf ( R_19c2_14871098 , C0 );
buf ( R_d3e_14870198 , C0 );
buf ( R_71f_123b6e78 , n54335 );
buf ( R_b3e_11631138 , C0 );
buf ( R_115d_1008bd58 , n54349 );
buf ( R_135d_13cd9d78 , n54360 );
buf ( R_177c_11629258 , n54361 );
buf ( R_197c_13bec8f8 , n54362 );
buf ( R_96e_1162bff8 , C0 );
buf ( R_f0e_17010f68 , C0 );
buf ( R_8ef_13dd96d8 , n54363 );
buf ( R_f8d_13cd51d8 , n54369 );
buf ( R_152d_13d1f8d8 , n54400 );
buf ( R_15ac_12fc1418 , n54401 );
buf ( R_ee8_13d55658 , n54402 );
buf ( R_994_13c086f8 , n54403 );
buf ( R_8c9_1162f838 , n54426 );
buf ( R_fb3_11c6c7b8 , n54427 );
buf ( R_1507_14b218f8 , n54428 );
buf ( R_15d2_11c6e978 , C0 );
buf ( R_ed3_13b93018 , n54429 );
buf ( R_9a9_140ac3f8 , n54437 );
buf ( R_8b4_150e2e38 , n54438 );
buf ( R_fc8_14875238 , n54439 );
buf ( R_14f2_13cd1718 , C0 );
buf ( R_15e7_150e0e58 , n54440 );
buf ( R_c1a_13d3c198 , C0 );
buf ( R_5fb_156b22f8 , n54441 );
buf ( R_643_117ea698 , n54442 );
buf ( R_c62_1162c598 , C0 );
buf ( R_1239_15817938 , n54452 );
buf ( R_1281_158887d8 , n54479 );
buf ( R_1858_13bea9b8 , n54480 );
buf ( R_18a0_123bfcf8 , n54481 );
buf ( R_98c_13c21f18 , n54482 );
buf ( R_ef0_13d51418 , n54483 );
buf ( R_8d1_12fc06f8 , n54501 );
buf ( R_fab_14a127f8 , n54502 );
buf ( R_150f_15817398 , n54503 );
buf ( R_15ca_156b71b8 , C0 );
buf ( R_c95_123be2b8 , n54514 );
buf ( R_be7_1162d858 , n54515 );
buf ( R_5c8_15feeca8 , n54516 );
buf ( R_676_13d37e18 , C0 );
buf ( R_1206_13ddcc98 , C0 );
buf ( R_12b4_10087938 , n54517 );
buf ( R_1825_1486a298 , n54527 );
buf ( R_18d3_17018f88 , n54528 );
buf ( R_d5b_150e0958 , n54529 );
buf ( R_b21_14b21e98 , n54544 );
buf ( R_73c_13bec858 , n54545 );
buf ( R_1140_13b98798 , n54546 );
buf ( R_137a_13dd7018 , C0 );
buf ( R_175f_15ff7f88 , n54547 );
buf ( R_1999_117f2118 , n54555 );
buf ( R_d4a_13df40d8 , C0 );
buf ( R_b32_13c268d8 , C0 );
buf ( R_72b_11632c18 , n54556 );
buf ( R_1151_11638898 , n54564 );
buf ( R_1369_117f5138 , n54575 );
buf ( R_1770_124c2a58 , n54576 );
buf ( R_1988_150dfaf8 , n54577 );
buf ( R_db1_13bf06d8 , n54587 );
buf ( R_792_13ccb638 , C0 );
buf ( R_acb_13d2a378 , n54588 );
buf ( R_10ea_13d2b598 , C0 );
buf ( R_13d0_1700b388 , n54589 );
buf ( R_1709_1162a298 , n54602 );
buf ( R_19ef_150de1f8 , n54603 );
buf ( R_ae3_14b24738 , n54604 );
buf ( R_d99_156abef8 , n54615 );
buf ( R_77a_13c0f3b8 , C0 );
buf ( R_1102_11632358 , C0 );
buf ( R_13b8_13c29c18 , n54616 );
buf ( R_1721_14870f58 , n54619 );
buf ( R_19d7_13de38b8 , n54620 );
buf ( R_6d8_1580ebf8 , n54621 );
buf ( R_566_140b4f58 , n54622 );
buf ( R_cf7_13d26778 , n54623 );
buf ( R_b85_13df3958 , n54631 );
buf ( R_11a4_140b1178 , n54632 );
buf ( R_1316_13c24718 , C0 );
buf ( R_17c3_13df1e78 , n54633 );
buf ( R_1935_14a13798 , n54652 );
buf ( R_a0d_14a0f198 , n54661 );
buf ( R_850_1700cbe8 , n54662 );
buf ( R_e6f_117ee6f8 , n54663 );
buf ( R_102c_156ae3d8 , n54664 );
buf ( R_148e_17014208 , C0 );
buf ( R_164b_123b8638 , n54665 );
buf ( R_f2f_13ccded8 , n54666 );
buf ( R_910_158144b8 , n54667 );
buf ( R_94d_13de1dd8 , n54674 );
buf ( R_f6c_140aca38 , n54675 );
buf ( R_154e_158131f8 , C0 );
buf ( R_158b_123b5078 , n54676 );
buf ( R_70c_1162a338 , n54677 );
buf ( R_b51_13df4c18 , n54724 );
buf ( R_d2b_123bacf8 , n54725 );
buf ( R_1170_13ddca18 , n54726 );
buf ( R_134a_123bdb38 , C0 );
buf ( R_178f_14a0df78 , n54727 );
buf ( R_1969_13c0e918 , n54735 );
buf ( R_ec1_13c0ddd8 , n54744 );
buf ( R_8a2_13dd9638 , C0 );
buf ( R_9bb_14a13d38 , n54745 );
buf ( R_fda_14876098 , C0 );
buf ( R_14e0_117ea9b8 , n54746 );
buf ( R_15f9_13d4fcf8 , n54771 );
buf ( R_d3b_150e4a58 , n54772 );
buf ( R_71c_150dba98 , n54773 );
buf ( R_b41_100844b8 , n54781 );
buf ( R_1160_14a16498 , n54782 );
buf ( R_135a_156b8838 , C0 );
buf ( R_177f_13ccedd8 , n54783 );
buf ( R_1979_156ad7f8 , n54791 );
buf ( R_80a_11c686b8 , C0 );
buf ( R_a53_13d54ed8 , n54792 );
buf ( R_e29_124c3138 , n54801 );
buf ( R_1072_13d5c598 , C0 );
buf ( R_1448_156b5098 , n54802 );
buf ( R_1691_13bf8478 , n54813 );
buf ( R_1a67_13d3a898 , n54814 );
buf ( R_aa1_13ccbd18 , n54823 );
buf ( R_7bc_13ccc218 , n54824 );
buf ( R_ddb_15812618 , n54825 );
buf ( R_10c0_15816d58 , n54826 );
buf ( R_13fa_14b29a58 , C0 );
buf ( R_16df_10084eb8 , n54827 );
buf ( R_1a19_11c70a98 , n54831 );
buf ( R_a1e_13de1338 , C0 );
buf ( R_83f_123bc5f8 , n54832 );
buf ( R_e5e_13c25258 , C0 );
buf ( R_103d_123b2738 , n54847 );
buf ( R_147d_13d53e98 , n54859 );
buf ( R_165c_123b57f8 , n54860 );
buf ( R_c74_14b242d8 , n54861 );
buf ( R_c08_13ded7d8 , n54862 );
buf ( R_5e9_15816178 , n54871 );
buf ( R_655_13c026b8 , n54883 );
buf ( R_1227_123b72d8 , n54884 );
buf ( R_1293_1008c6b8 , n54885 );
buf ( R_1846_13c22af8 , C0 );
buf ( R_18b2_150dd4d8 , C0 );
buf ( R_a14_11632038 , n54886 );
buf ( R_849_123c1af8 , n54894 );
buf ( R_e68_15887658 , n54895 );
buf ( R_1033_13bf8518 , n54896 );
buf ( R_1487_1007fc38 , n54897 );
buf ( R_1652_11635418 , C0 );
buf ( R_68e_11630eb8 , C0 );
buf ( R_bcf_1486c4f8 , n54898 );
buf ( R_cad_150e5c78 , n54907 );
buf ( R_5b0_13d20c38 , n54912 );
buf ( R_11ee_13df5938 , C0 );
buf ( R_12cc_156aee78 , n54913 );
buf ( R_180d_13d29dd8 , n54922 );
buf ( R_18eb_13cd2bb8 , n54923 );
buf ( R_7e9_13b903b8 , n54931 );
buf ( R_e08_14a11498 , n54932 );
buf ( R_a74_13c02a78 , n54933 );
buf ( R_1093_123bddb8 , n54934 );
buf ( R_1427_1580dd98 , n54935 );
buf ( R_16b2_123b89f8 , C0 );
buf ( R_1a46_150dff58 , C0 );
buf ( R_c81_140ac718 , n54944 );
buf ( R_bfb_117e8f78 , n54945 );
buf ( R_5dc_13cd21b8 , n54946 );
buf ( R_662_11c6af58 , C0 );
buf ( R_121a_13dd6bb8 , C0 );
buf ( R_12a0_156af7d8 , n54947 );
buf ( R_1839_10083a18 , n54956 );
buf ( R_18bf_13cd63f8 , n54957 );
buf ( R_d4d_14b1c218 , n54967 );
buf ( R_b2f_14a168f8 , n54968 );
buf ( R_72e_15885178 , C0 );
buf ( R_114e_14866878 , C0 );
buf ( R_136c_13d5ce58 , n54969 );
buf ( R_176d_15883e18 , n54982 );
buf ( R_198b_123ba938 , n54983 );
buf ( R_bb0_11635198 , n54984 );
buf ( R_6ad_14b295f8 , n54996 );
buf ( R_591_123b56b8 , n54997 );
buf ( R_ccc_13c02f78 , n54998 );
buf ( R_11cf_13dedd78 , n54999 );
buf ( R_12eb_156ab598 , n55000 );
buf ( R_17ee_117f2a78 , C0 );
buf ( R_190a_1162b238 , C0 );
buf ( R_7d4_14a0fe18 , n55001 );
buf ( R_df3_14b1e478 , n55002 );
buf ( R_a89_13dd9278 , n55042 );
buf ( R_10a8_13d52958 , n55043 );
buf ( R_1412_11c6f198 , C0 );
buf ( R_16c7_13d27d58 , n55044 );
buf ( R_1a31_140b9d78 , n55048 );
buf ( R_c19_1700d408 , n55076 );
buf ( R_5fa_13df88b8 , C0 );
buf ( R_644_13d23938 , n55077 );
buf ( R_c63_1162e258 , n55078 );
buf ( R_1238_13df9a38 , n55079 );
buf ( R_1282_13c2acf8 , C0 );
buf ( R_1857_13cd2ed8 , n55080 );
buf ( R_18a1_156aefb8 , n55090 );
buf ( R_6f0_140ae658 , n55091 );
buf ( R_b6d_123b4178 , n55102 );
buf ( R_d0f_150df0f8 , n55103 );
buf ( R_118c_14a17898 , n55104 );
buf ( R_132e_13bed758 , C0 );
buf ( R_17ab_13cd0d18 , n55105 );
buf ( R_194d_1008c438 , n55132 );
buf ( R_802_13d3e5d8 , C0 );
buf ( R_e21_14a0aaf8 , n55141 );
buf ( R_a5b_13bf7e38 , n55142 );
buf ( R_107a_13d1ed98 , C0 );
buf ( R_1440_124c4d58 , n55143 );
buf ( R_1699_140b0318 , n55154 );
buf ( R_1a5f_124c5618 , n55155 );
buf ( R_8fc_13bebd18 , n55156 );
buf ( R_961_12fbe358 , n55162 );
buf ( R_f1b_13ddafd8 , n55163 );
buf ( R_f80_1486f478 , n55164 );
buf ( R_153a_116341f8 , C0 );
buf ( R_159f_1008d338 , n55165 );
buf ( R_ada_15812f78 , C0 );
buf ( R_da2_156b5ef8 , C0 );
buf ( R_783_123ba898 , n55166 );
buf ( R_10f9_123b7a58 , n55180 );
buf ( R_13c1_13d3bfb8 , n55192 );
buf ( R_1718_156b8018 , n55193 );
buf ( R_19e0_13dd4ef8 , n55194 );
buf ( R_6cb_117f2258 , n55195 );
buf ( R_573_1162dfd8 , n55196 );
buf ( R_cea_13d5be18 , C0 );
buf ( R_b92_13c01998 , C0 );
buf ( R_11b1_1700a208 , n55206 );
buf ( R_1309_117e8898 , n55216 );
buf ( R_17d0_156b8d38 , n55217 );
buf ( R_1928_14a0f738 , n55218 );
buf ( R_eb1_156b8f18 , n55227 );
buf ( R_892_11c69018 , C0 );
buf ( R_9cb_13bed1b8 , n55228 );
buf ( R_fea_13d2b3b8 , C0 );
buf ( R_14d0_13ccf698 , n55229 );
buf ( R_1609_13cd30b8 , n55260 );
buf ( R_67f_13cd88d8 , n55261 );
buf ( R_c9e_1580ee78 , C0 );
buf ( R_bde_123b3138 , C0 );
buf ( R_5bf_117f0b38 , n55262 );
buf ( R_11fd_1162f3d8 , n55297 );
buf ( R_12bd_13bf9698 , n55321 );
buf ( R_181c_13bf7758 , n55322 );
buf ( R_18dc_15817258 , n55323 );
buf ( R_c8c_13b97258 , n55324 );
buf ( R_bf0_13c26d38 , n55325 );
buf ( R_5d1_14875af8 , n55334 );
buf ( R_66d_1700eda8 , n55346 );
buf ( R_120f_156b0a98 , n55347 );
buf ( R_12ab_1486c278 , n55348 );
buf ( R_182e_116366d8 , C0 );
buf ( R_18ca_11c708b8 , C0 );
buf ( R_f2e_13dddb98 , C0 );
buf ( R_90f_13b8e3d8 , n55349 );
buf ( R_94e_117f3c98 , C0 );
buf ( R_f6d_13bf7a78 , n55371 );
buf ( R_154d_13df8c78 , n55382 );
buf ( R_158c_13d278f8 , n55383 );
buf ( R_702_13de3598 , C0 );
buf ( R_b5b_13d45bf8 , n55384 );
buf ( R_d21_156ac038 , n55393 );
buf ( R_117a_14b292d8 , C0 );
buf ( R_1340_123bbab8 , n55394 );
buf ( R_1799_13df1018 , n55412 );
buf ( R_195f_13b92e38 , n55413 );
buf ( R_d38_156afaf8 , n55414 );
buf ( R_719_13d1d498 , n55425 );
buf ( R_b44_13df7238 , n55426 );
buf ( R_1163_13b91358 , n55427 );
buf ( R_1357_13d5bcd8 , n55428 );
buf ( R_1782_1486c138 , C0 );
buf ( R_1976_14b1de38 , C0 );
buf ( R_695_13b93b58 , n55439 );
buf ( R_bc8_13dfb3d8 , n55440 );
buf ( R_cb4_15817078 , n55441 );
buf ( R_5a9_156b6998 , n55446 );
buf ( R_11e7_13bf3298 , n55447 );
buf ( R_12d3_14b28338 , n55448 );
buf ( R_1806_123b6dd8 , C0 );
buf ( R_18f2_13d40338 , C0 );
buf ( R_a06_158876f8 , C0 );
buf ( R_857_14874dd8 , n55449 );
buf ( R_e76_13bf0958 , C0 );
buf ( R_1025_13d59438 , n55457 );
buf ( R_1495_14870238 , n55469 );
buf ( R_1644_15ff4d88 , n55470 );
buf ( R_6fb_156b9378 , n55471 );
buf ( R_b62_123bb298 , C0 );
buf ( R_d1a_117ee1f8 , C0 );
buf ( R_1181_148748d8 , n55485 );
buf ( R_1339_1580de38 , n55496 );
buf ( R_17a0_13dd7478 , n55497 );
buf ( R_1958_156ae5b8 , n55498 );
buf ( R_97a_117eaff8 , C0 );
buf ( R_f02_13d538f8 , C0 );
buf ( R_8e3_13c107b8 , n55499 );
buf ( R_f99_1580efb8 , n55503 );
buf ( R_1521_148676d8 , n55511 );
buf ( R_15b8_13b93e78 , n55512 );
buf ( R_829_13b954f8 , n55522 );
buf ( R_a34_156b03b8 , n55523 );
buf ( R_e48_15813d38 , n55524 );
buf ( R_1053_13cd3478 , n55525 );
buf ( R_1467_13b8be58 , n55526 );
buf ( R_1672_13cd1df8 , C0 );
buf ( R_e89_13de0078 , n55538 );
buf ( R_9f3_156b0598 , n55539 );
buf ( R_86a_13b94378 , C0 );
buf ( R_1012_123bf618 , C0 );
buf ( R_14a8_13becdf8 , n55540 );
buf ( R_1631_1486c9f8 , n55551 );
buf ( R_acd_1008bfd8 , n55563 );
buf ( R_daf_123b59d8 , n55564 );
buf ( R_790_13d2bd18 , n55565 );
buf ( R_10ec_1700b6a8 , n55566 );
buf ( R_13ce_13df2a58 , C0 );
buf ( R_170b_14b26178 , n55567 );
buf ( R_19ed_148709b8 , n55571 );
buf ( R_a31_13cd7d98 , n55577 );
buf ( R_82c_140b1e98 , n55578 );
buf ( R_e4b_116316d8 , n55579 );
buf ( R_1050_13d3d138 , n55580 );
buf ( R_146a_123bd318 , C0 );
buf ( R_166f_140ad118 , n55581 );
buf ( R_eac_1007f418 , n55582 );
buf ( R_88d_13bf99b8 , n55597 );
buf ( R_9d0_17010748 , n55598 );
buf ( R_fef_1580b138 , n55599 );
buf ( R_14cb_13d44258 , n55600 );
buf ( R_160e_11632a38 , C0 );
buf ( R_826_13c24cb8 , C0 );
buf ( R_a37_158112b8 , n55601 );
buf ( R_e45_15fee168 , n55611 );
buf ( R_1056_15fedc68 , C0 );
buf ( R_1464_13d3fa78 , n55612 );
buf ( R_1675_14b28dd8 , n55617 );
buf ( R_eb6_11c69518 , C0 );
buf ( R_897_11c69338 , n55618 );
buf ( R_9c6_156ad258 , C0 );
buf ( R_fe5_14b1f4b8 , n55623 );
buf ( R_14d5_14871a98 , n55635 );
buf ( R_1604_13beed38 , n55636 );
buf ( R_9ef_14a126b8 , n55637 );
buf ( R_e8d_13c07578 , n55645 );
buf ( R_86e_13ded738 , C0 );
buf ( R_100e_100810d8 , C0 );
buf ( R_14ac_13cce158 , n55646 );
buf ( R_162d_13c0adb8 , n55659 );
buf ( R_7cb_14a0acd8 , n55660 );
buf ( R_dea_123c0798 , C0 );
buf ( R_a92_13d25238 , C0 );
buf ( R_10b1_13d55478 , n55666 );
buf ( R_1409_1587f638 , n55676 );
buf ( R_16d0_13c02ed8 , n55677 );
buf ( R_1a28_14a12398 , n55678 );
buf ( R_ee0_13d1ffb8 , n55679 );
buf ( R_99c_14a0f418 , n55680 );
buf ( R_8c1_14b25818 , n55707 );
buf ( R_fbb_123b70f8 , n55708 );
buf ( R_14ff_1580bf98 , n55709 );
buf ( R_15da_140ba138 , C0 );
buf ( R_687_14b23fb8 , n55710 );
buf ( R_bd6_13dd71f8 , C0 );
buf ( R_ca6_123bd098 , C0 );
buf ( R_5b7_117e8cf8 , n55711 );
buf ( R_11f5_15815318 , n55751 );
buf ( R_12c5_14a0f7d8 , n55774 );
buf ( R_1814_170116e8 , n55775 );
buf ( R_18e4_12fc1d78 , n55776 );
buf ( R_812_12fc0018 , C0 );
buf ( R_a4b_13bf22f8 , n55777 );
buf ( R_e31_13bee338 , n55787 );
buf ( R_106a_13d56a58 , C0 );
buf ( R_1450_1580a738 , n55788 );
buf ( R_1689_14a0c218 , n55799 );
buf ( R_e85_156aa878 , n55806 );
buf ( R_9f7_13d246f8 , n55807 );
buf ( R_866_15ffb868 , C0 );
buf ( R_1016_156af698 , C0 );
buf ( R_14a4_11c6ec98 , n55808 );
buf ( R_1635_15ff7588 , n55821 );
buf ( R_8ee_140ae338 , C0 );
buf ( R_96f_13d3b8d8 , n55822 );
buf ( R_f0d_13d4fa78 , n55827 );
buf ( R_f8e_13d541b8 , C0 );
buf ( R_152c_156b2258 , n55828 );
buf ( R_15ad_13d58218 , n55852 );
buf ( R_9de_124c3458 , C0 );
buf ( R_e9e_123b9038 , C0 );
buf ( R_87f_117f0958 , n55853 );
buf ( R_ffd_13c27f58 , n55865 );
buf ( R_14bd_13cd71b8 , n55876 );
buf ( R_161c_156b6178 , n55877 );
buf ( R_aec_14866b98 , n55878 );
buf ( R_d90_10081718 , n55879 );
buf ( R_771_1007ee78 , n55888 );
buf ( R_110b_14b24f58 , n55889 );
buf ( R_13af_158110d8 , n55890 );
buf ( R_172a_11c6feb8 , C0 );
buf ( R_19ce_11c6fc38 , C0 );
buf ( R_6d4_15ff47e8 , n55891 );
buf ( R_56a_17018268 , n55892 );
buf ( R_cf3_150e21b8 , n55893 );
buf ( R_b89_13cd67b8 , n55901 );
buf ( R_11a8_13c0ab38 , n55902 );
buf ( R_1312_15881758 , C0 );
buf ( R_17c7_1580cf38 , n55903 );
buf ( R_1931_11c6b4f8 , n55928 );
buf ( R_7be_13d51918 , C0 );
buf ( R_ddd_10083fb8 , n55938 );
buf ( R_a9f_140b7b18 , n55939 );
buf ( R_10be_1162c138 , C0 );
buf ( R_13fc_13b967b8 , n55940 );
buf ( R_16dd_15ffb728 , n55951 );
buf ( R_1a1b_13d3ab18 , n55952 );
buf ( R_a2e_1580aeb8 , C0 );
buf ( R_82f_14b26cb8 , n55953 );
buf ( R_e4e_13dec798 , C0 );
buf ( R_104d_13de2af8 , n55966 );
buf ( R_146d_156b1998 , n55976 );
buf ( R_166c_117f5958 , n55977 );
buf ( R_d50_156b51d8 , n55978 );
buf ( R_b2c_12fc0478 , n55979 );
buf ( R_731_15ffaa08 , n55988 );
buf ( R_114b_13ddbed8 , n55989 );
buf ( R_136f_11c6c718 , n55990 );
buf ( R_176a_11628f38 , C0 );
buf ( R_198e_150e3518 , C0 );
buf ( R_ed9_15ff7948 , n56001 );
buf ( R_9a3_13c1fad8 , n56002 );
buf ( R_8ba_116386b8 , C0 );
buf ( R_fc2_1700f7a8 , C0 );
buf ( R_14f8_117f15d8 , n56003 );
buf ( R_15e1_150dcd58 , n56031 );
buf ( R_b16_13c1c1f8 , C0 );
buf ( R_d66_13b8b1d8 , C0 );
buf ( R_747_158864d8 , n56032 );
buf ( R_1135_156b68f8 , n56043 );
buf ( R_1385_1580b278 , n56055 );
buf ( R_1754_156add98 , n56056 );
buf ( R_19a4_13d4fd98 , n56057 );
buf ( R_823_11c6f2d8 , n56058 );
buf ( R_a3a_14871318 , C0 );
buf ( R_e42_156ade38 , C0 );
buf ( R_1059_13c0f318 , n56066 );
buf ( R_1461_14a1a138 , n56077 );
buf ( R_1678_14a0fd78 , n56078 );
buf ( R_8d9_158837d8 , n56098 );
buf ( R_984_15882d38 , n56099 );
buf ( R_ef8_15816998 , n56100 );
buf ( R_fa3_15815458 , n56101 );
buf ( R_1517_156ad898 , n56102 );
buf ( R_15c2_11630c38 , C0 );
buf ( R_af3_13beae18 , n56103 );
buf ( R_d89_117e8938 , n56112 );
buf ( R_76a_123bceb8 , C0 );
buf ( R_1112_13c20c58 , C0 );
buf ( R_13a8_117f4a58 , n56113 );
buf ( R_1731_1008a818 , n56121 );
buf ( R_19c7_13d38bd8 , n56122 );
buf ( R_b04_156aed38 , n56123 );
buf ( R_d78_13cd7758 , n56124 );
buf ( R_759_11629938 , n56135 );
buf ( R_1123_15ffb908 , n56136 );
buf ( R_1397_13d37a58 , n56137 );
buf ( R_1742_13d237f8 , C0 );
buf ( R_19b6_14b20778 , C0 );
buf ( R_c64_13c1fdf8 , n56138 );
buf ( R_c18_12fc23b8 , n56139 );
buf ( R_5f9_13b8f238 , n56150 );
buf ( R_645_140b2118 , n56159 );
buf ( R_1237_1162dad8 , n56160 );
buf ( R_1283_14a18798 , n56161 );
buf ( R_1856_117f4878 , C0 );
buf ( R_18a2_13d53998 , C0 );
buf ( R_f2d_100818f8 , n56180 );
buf ( R_90e_11629898 , C0 );
buf ( R_94f_15888738 , n56181 );
buf ( R_f6e_14a188d8 , C0 );
buf ( R_154c_14a147d8 , n56182 );
buf ( R_158d_15ff0a08 , n56183 );
buf ( R_9eb_117ef2d8 , n56184 );
buf ( R_e91_1580e3d8 , n56215 );
buf ( R_872_13c0c7f8 , C0 );
buf ( R_100a_117f81f8 , C0 );
buf ( R_14b0_124c2f58 , n56216 );
buf ( R_1629_14a0b6d8 , n56223 );
buf ( R_656_15886bb8 , C0 );
buf ( R_c75_156b0db8 , n56234 );
buf ( R_c07_124c4cb8 , n56235 );
buf ( R_5e8_1162f298 , n56236 );
buf ( R_1226_13b8e018 , C0 );
buf ( R_1294_13b91ad8 , n56237 );
buf ( R_1845_13cd83d8 , n56248 );
buf ( R_18b3_13d1e118 , n56249 );
buf ( R_ba0_156b4698 , n56250 );
buf ( R_6bd_13c0ec38 , n56260 );
buf ( R_581_13d1d8f8 , n56261 );
buf ( R_cdc_13cd9378 , n56262 );
buf ( R_11bf_123b6c98 , n56263 );
buf ( R_12fb_150e3018 , n56264 );
buf ( R_17de_14b20458 , C0 );
buf ( R_191a_123b2cd8 , C0 );
buf ( R_d5e_14a10278 , C0 );
buf ( R_b1e_13df7418 , C0 );
buf ( R_73f_1587b998 , n56265 );
buf ( R_113d_13d58498 , n56281 );
buf ( R_137d_14a11b78 , n56293 );
buf ( R_175c_1587b218 , n56294 );
buf ( R_199c_17017408 , n56295 );
buf ( R_b09_15884f98 , n56305 );
buf ( R_d73_1580b4f8 , n56306 );
buf ( R_754_15811d58 , n56307 );
buf ( R_1128_10084d78 , n56308 );
buf ( R_1392_14a15db8 , C0 );
buf ( R_1747_17018588 , n56309 );
buf ( R_19b1_13dd9f98 , n56317 );
buf ( R_d35_14a11858 , n56328 );
buf ( R_716_156b9c38 , C0 );
buf ( R_b47_140af4b8 , n56329 );
buf ( R_1166_13ccdcf8 , C0 );
buf ( R_1354_13d41738 , n56330 );
buf ( R_1785_1162d218 , n56343 );
buf ( R_1973_14a18338 , n56344 );
buf ( R_a2b_13c1e6d8 , n56345 );
buf ( R_832_13df5c58 , C0 );
buf ( R_e51_156ab278 , n56355 );
buf ( R_104a_14a108b8 , C0 );
buf ( R_1470_15887bf8 , n56356 );
buf ( R_1669_158828d8 , n56366 );
buf ( R_e81_1007dc58 , n56377 );
buf ( R_9fb_1486fb58 , n56378 );
buf ( R_862_156ab138 , C0 );
buf ( R_101a_13d5a798 , C0 );
buf ( R_14a0_13d38818 , n56379 );
buf ( R_1639_1162abf8 , n56390 );
buf ( R_ba5_140b4af8 , n56399 );
buf ( R_6b8_1580d898 , n56400 );
buf ( R_586_15ff8488 , n56401 );
buf ( R_cd7_156b7e38 , n56402 );
buf ( R_11c4_117ecad8 , n56403 );
buf ( R_12f6_17015ba8 , C0 );
buf ( R_17e3_13c1dd78 , n56404 );
buf ( R_1915_14a17f78 , n56432 );
buf ( R_aff_140aba98 , n56433 );
buf ( R_d7d_148714f8 , n56443 );
buf ( R_75e_10084418 , C0 );
buf ( R_111e_11635918 , C0 );
buf ( R_139c_1580e0b8 , n56444 );
buf ( R_173d_13deffd8 , n56446 );
buf ( R_19bb_13df9df8 , n56447 );
buf ( R_7dd_13d28898 , n56454 );
buf ( R_dfc_156b9ff8 , n56455 );
buf ( R_a80_13ddc8d8 , n56456 );
buf ( R_109f_13cd2cf8 , n56457 );
buf ( R_141b_12fc10f8 , n56458 );
buf ( R_16be_13bf0098 , C0 );
buf ( R_1a3a_156b79d8 , C0 );
buf ( R_9d5_15ff1908 , n56468 );
buf ( R_ea7_14a124d8 , n56469 );
buf ( R_888_13deebd8 , n56470 );
buf ( R_ff4_13cd7b18 , n56471 );
buf ( R_14c6_13cd5d18 , C0 );
buf ( R_1613_123bc198 , n56472 );
buf ( R_677_13c0c758 , n56473 );
buf ( R_c96_13c0d838 , C0 );
buf ( R_be6_1162cf98 , C0 );
buf ( R_5c7_1162f1f8 , n56474 );
buf ( R_1205_156b94b8 , n56485 );
buf ( R_12b5_158816b8 , n56512 );
buf ( R_1824_13c04f58 , n56513 );
buf ( R_18d4_13beb958 , n56514 );
buf ( R_f1a_124c4f38 , C0 );
buf ( R_8fb_13c1e9f8 , n56515 );
buf ( R_962_14a15ef8 , C0 );
buf ( R_f81_1580d438 , n56534 );
buf ( R_1539_14b267b8 , n56542 );
buf ( R_15a0_15ff32a8 , n56543 );
buf ( R_d28_156b3fb8 , n56544 );
buf ( R_709_117ea4b8 , n56554 );
buf ( R_b54_13c04c38 , n56555 );
buf ( R_1173_15810778 , n56556 );
buf ( R_1347_13dd5f38 , n56557 );
buf ( R_1792_13d39858 , C0 );
buf ( R_1966_12fc2098 , C0 );
buf ( R_a1b_123c17d8 , n56558 );
buf ( R_842_13bf4738 , C0 );
buf ( R_e61_13cd0958 , n56564 );
buf ( R_103a_13ccdbb8 , C0 );
buf ( R_1480_117f1e98 , n56565 );
buf ( R_1659_13c1fcb8 , n56576 );
buf ( R_820_17013088 , n56577 );
buf ( R_a3d_11c6bc78 , n56584 );
buf ( R_e3f_123c0e78 , n56585 );
buf ( R_105c_13dd87d8 , n56586 );
buf ( R_145e_13d5a3d8 , C0 );
buf ( R_167b_14a19878 , n56587 );
buf ( R_ebb_13def998 , n56588 );
buf ( R_89c_1486e898 , n56589 );
buf ( R_9c1_13cd04f8 , n56597 );
buf ( R_fe0_15fee7a8 , n56598 );
buf ( R_14da_13b95818 , C0 );
buf ( R_15ff_117f1538 , n56599 );
buf ( R_8d0_13ccd078 , n56600 );
buf ( R_98d_13cceab8 , n56608 );
buf ( R_eef_15ff2308 , n56609 );
buf ( R_fac_13df65b8 , n56610 );
buf ( R_150e_13bed398 , C0 );
buf ( R_15cb_1580a558 , n56611 );
buf ( R_663_13c24218 , n56612 );
buf ( R_c82_11633bb8 , C0 );
buf ( R_bfa_117f1d58 , C0 );
buf ( R_5db_13c0d798 , n56613 );
buf ( R_1219_156b0f98 , n56624 );
buf ( R_12a1_15811e98 , n56648 );
buf ( R_1838_123c2098 , n56649 );
buf ( R_18c0_13ddb258 , n56650 );
buf ( R_bbb_13c08dd8 , n56651 );
buf ( R_6a2_14870cd8 , C0 );
buf ( R_59c_1700ffc8 , n56656 );
buf ( R_cc1_13d5b0f8 , n56665 );
buf ( R_11da_14b1dcf8 , C0 );
buf ( R_12e0_14b29c38 , n56666 );
buf ( R_17f9_13ddb438 , n56676 );
buf ( R_18ff_1162d538 , n56677 );
buf ( R_ecc_123bde58 , n56678 );
buf ( R_9b0_1587f458 , n56679 );
buf ( R_8ad_10082e38 , n56700 );
buf ( R_fcf_14a0e798 , n56701 );
buf ( R_14eb_140ad258 , n56702 );
buf ( R_15ee_117f3158 , C0 );
buf ( R_d13_13c25e38 , n56703 );
buf ( R_6f4_156b4918 , n56704 );
buf ( R_b69_11c6e8d8 , n56738 );
buf ( R_1188_13cd35b8 , n56739 );
buf ( R_1332_11637d58 , C0 );
buf ( R_17a7_117f6a38 , n56740 );
buf ( R_1951_156b6b78 , n56764 );
buf ( R_acf_13d503d8 , n56765 );
buf ( R_dad_13cd3838 , n56775 );
buf ( R_78e_13b929d8 , C0 );
buf ( R_10ee_1587c438 , C0 );
buf ( R_13cc_1587b3f8 , n56776 );
buf ( R_170d_12fbf9d8 , n56787 );
buf ( R_19eb_15ff53c8 , n56788 );
buf ( R_8c8_12fbe038 , n56789 );
buf ( R_ee7_13c03dd8 , n56790 );
buf ( R_995_13d50518 , n56798 );
buf ( R_fb4_156b0e58 , n56799 );
buf ( R_1506_156b9e18 , C0 );
buf ( R_15d3_123b5ed8 , n56800 );
buf ( R_b9b_13dfa118 , n56801 );
buf ( R_6c2_14b1d618 , C0 );
buf ( R_57c_13d464b8 , n56802 );
buf ( R_ce1_13d27358 , n56811 );
buf ( R_11ba_13cda458 , C0 );
buf ( R_1300_13dec478 , n56812 );
buf ( R_17d9_156af918 , n56822 );
buf ( R_191f_14a0d578 , n56823 );
buf ( R_7e4_117f6c18 , n56824 );
buf ( R_e03_13b8c718 , n56825 );
buf ( R_a79_13d52db8 , n56834 );
buf ( R_1098_13cd2438 , n56835 );
buf ( R_1422_13cd7f78 , C0 );
buf ( R_16b7_14b28518 , n56836 );
buf ( R_1a41_150e4d78 , n56841 );
buf ( R_ae5_17012048 , n56854 );
buf ( R_d97_1162ab58 , n56855 );
buf ( R_778_13d52098 , n56856 );
buf ( R_1104_13dd7a18 , n56857 );
buf ( R_13b6_14a17118 , C0 );
buf ( R_1723_13d50018 , n56858 );
buf ( R_19d5_117edc58 , n56866 );
buf ( R_d53_13c0ae58 , n56867 );
buf ( R_b29_13b95c78 , n56878 );
buf ( R_734_14a0f558 , n56879 );
buf ( R_1148_117f6218 , n56880 );
buf ( R_1372_11c6cd58 , C0 );
buf ( R_1767_11c691f8 , n56881 );
buf ( R_1991_13cd58b8 , n56889 );
buf ( R_f2c_15814d78 , n56890 );
buf ( R_90d_158848b8 , n56894 );
buf ( R_950_140b3798 , n56895 );
buf ( R_f6f_14a1a318 , n56896 );
buf ( R_154b_11632218 , n56897 );
buf ( R_158e_14a0b1d8 , C0 );
buf ( R_ec6_13d37b98 , C0 );
buf ( R_8a7_1580e6f8 , n56898 );
buf ( R_9b6_14a0cc18 , C0 );
buf ( R_fd5_1580cc18 , n56913 );
buf ( R_14e5_13b8fd78 , n56925 );
buf ( R_15f4_170165a8 , n56926 );
buf ( R_7c0_100854f8 , n56927 );
buf ( R_ddf_13b92898 , n56928 );
buf ( R_a9d_1162c318 , n56941 );
buf ( R_10bc_140b7d98 , n56942 );
buf ( R_13fe_13cd60d8 , C0 );
buf ( R_16db_156aaf58 , n56943 );
buf ( R_1a1d_13cd9ff8 , n56947 );
buf ( R_7f5_13b9a1d8 , n56954 );
buf ( R_e14_123bf078 , n56955 );
buf ( R_a68_150dbbd8 , n56956 );
buf ( R_1087_1587ad18 , n56957 );
buf ( R_1433_13dd7978 , n56958 );
buf ( R_16a6_13df8458 , C0 );
buf ( R_1a52_11c70778 , C0 );
buf ( R_646_156ad618 , C0 );
buf ( R_c65_10086538 , n56967 );
buf ( R_c17_13ccb3b8 , n56968 );
buf ( R_5f8_1580f418 , n56969 );
buf ( R_1236_1587e558 , C0 );
buf ( R_1284_14a1a458 , n56970 );
buf ( R_1855_10084a58 , n56980 );
buf ( R_18a3_1700b1a8 , n56981 );
buf ( R_69c_156b9058 , n56982 );
buf ( R_bc1_13bee298 , n56993 );
buf ( R_cbb_13ccbbd8 , n56994 );
buf ( R_5a2_15813658 , n56999 );
buf ( R_11e0_1587e878 , n57000 );
buf ( R_12da_14b29d78 , C0 );
buf ( R_17ff_14a10b38 , n57001 );
buf ( R_18f9_14a16718 , n57030 );
buf ( R_adc_156ae6f8 , n57031 );
buf ( R_da0_13bf5db8 , n57032 );
buf ( R_781_13d42f98 , n57041 );
buf ( R_10fb_10085778 , n57042 );
buf ( R_13bf_123bf6b8 , n57043 );
buf ( R_171a_150deb58 , C0 );
buf ( R_19de_117ef918 , C0 );
buf ( R_9e7_13d54578 , n57044 );
buf ( R_e95_13d26ef8 , n57052 );
buf ( R_876_13d41698 , C0 );
buf ( R_1006_13c08f18 , C0 );
buf ( R_14b4_1700e268 , n57053 );
buf ( R_1625_13b96d58 , n57057 );
buf ( R_807_13cd8478 , n57058 );
buf ( R_e26_1700df48 , C0 );
buf ( R_a56_124c4ad8 , C0 );
buf ( R_1075_15883b98 , n57069 );
buf ( R_1445_15880218 , n57080 );
buf ( R_1694_13d218b8 , n57081 );
buf ( R_1a64_13ccac38 , n57082 );
buf ( R_a28_13cd9918 , n57083 );
buf ( R_835_140b35b8 , n57092 );
buf ( R_e54_14a179d8 , n57093 );
buf ( R_1047_14b26df8 , n57094 );
buf ( R_1473_156b60d8 , n57095 );
buf ( R_1666_14a165d8 , C0 );
buf ( R_b0e_14a15818 , C0 );
buf ( R_d6e_14a0c998 , C0 );
buf ( R_74f_13c24678 , n57096 );
buf ( R_112d_1162be18 , n57110 );
buf ( R_138d_13b92258 , n57119 );
buf ( R_174c_116339d8 , n57120 );
buf ( R_19ac_14b1b4f8 , n57121 );
buf ( R_bb5_13cd29d8 , n57133 );
buf ( R_6a8_1162e618 , n57134 );
buf ( R_596_13dd6398 , n57139 );
buf ( R_cc7_123b4b78 , n57140 );
buf ( R_11d4_15ff30c8 , n57141 );
buf ( R_12e6_14a0ff58 , C0 );
buf ( R_17f3_13ddb578 , n57142 );
buf ( R_1905_1486dfd8 , n57170 );
buf ( R_baa_14a15278 , C0 );
buf ( R_6b3_17011288 , n57171 );
buf ( R_58b_140b1c18 , n57172 );
buf ( R_cd2_13d24dd8 , C0 );
buf ( R_11c9_14b25278 , n57182 );
buf ( R_12f1_1587da18 , n57193 );
buf ( R_17e8_1587c078 , n57194 );
buf ( R_1910_12fc0978 , n57195 );
buf ( R_66e_17014348 , C0 );
buf ( R_c8d_123b7ff8 , n57205 );
buf ( R_bef_14a167b8 , n57206 );
buf ( R_5d0_13c1db98 , n57207 );
buf ( R_120e_13c0d518 , C0 );
buf ( R_12ac_13ccaf58 , n57208 );
buf ( R_182d_140b0098 , n57217 );
buf ( R_18cb_123b9e98 , n57218 );
buf ( R_8b3_13c0d298 , n57219 );
buf ( R_ed2_1580c538 , C0 );
buf ( R_9aa_124c51b8 , C0 );
buf ( R_fc9_13b8d118 , n57228 );
buf ( R_14f1_150e8978 , n57235 );
buf ( R_15e8_15884db8 , n57236 );
buf ( R_8e2_13bf6858 , C0 );
buf ( R_97b_150e7a78 , n57237 );
buf ( R_f01_14a13e78 , n57241 );
buf ( R_f9a_116364f8 , C0 );
buf ( R_1520_1162d678 , n57242 );
buf ( R_15b9_13d21a98 , n57260 );
buf ( R_7fa_123bbbf8 , C0 );
buf ( R_e19_13d59ed8 , n57271 );
buf ( R_a63_14a16678 , n57272 );
buf ( R_1082_13c09d78 , C0 );
buf ( R_1438_13bf2398 , n57273 );
buf ( R_16a1_14a16cb8 , n57286 );
buf ( R_1a57_13c28a98 , n57287 );
buf ( R_81d_1580d078 , n57295 );
buf ( R_a40_123bcd78 , n57296 );
buf ( R_e3c_117f2c58 , n57297 );
buf ( R_105f_13de2558 , n57298 );
buf ( R_145b_11633e38 , n57299 );
buf ( R_167e_1486d858 , C0 );
buf ( R_7f0_13b90458 , n57300 );
buf ( R_e0f_140ab138 , n57301 );
buf ( R_a6d_117ee838 , n57314 );
buf ( R_108c_13bf90f8 , n57315 );
buf ( R_142e_11632538 , C0 );
buf ( R_16ab_140b8d38 , n57316 );
buf ( R_1a4d_11c70bd8 , n57320 );
buf ( R_7d6_14b1e3d8 , C0 );
buf ( R_df5_1580eab8 , n57331 );
buf ( R_a87_14a10138 , n57332 );
buf ( R_10a6_117efa58 , C0 );
buf ( R_1414_1162b9b8 , n57333 );
buf ( R_16c5_14a10db8 , n57344 );
buf ( R_1a33_1486ebb8 , n57345 );
buf ( R_f0c_140b21b8 , n57346 );
buf ( R_8ed_11636d18 , n57371 );
buf ( R_970_13c0f818 , n57372 );
buf ( R_f8f_11632fd8 , n57373 );
buf ( R_152b_13beb778 , n57374 );
buf ( R_15ae_123b2eb8 , C0 );
buf ( R_e6b_13b8ded8 , n57375 );
buf ( R_a11_158133d8 , n57390 );
buf ( R_84c_13bef918 , n57391 );
buf ( R_1030_140b72f8 , n57392 );
buf ( R_148a_140b0598 , C0 );
buf ( R_164f_13d52778 , n57393 );
buf ( R_afa_123c0c98 , C0 );
buf ( R_d82_13cd1858 , C0 );
buf ( R_763_1580e298 , n57394 );
buf ( R_1119_1587c118 , n57407 );
buf ( R_13a1_158898b8 , n57419 );
buf ( R_1738_11c6f878 , n57420 );
buf ( R_19c0_1007ded8 , n57421 );
buf ( R_e7d_15811538 , n57428 );
buf ( R_9ff_13d245b8 , n57429 );
buf ( R_85e_13cd3018 , C0 );
buf ( R_101e_13d5d8f8 , C0 );
buf ( R_149c_13d5a978 , n57430 );
buf ( R_163d_13ccd438 , n57438 );
buf ( R_b8d_156aae18 , n57448 );
buf ( R_6d0_1162bb98 , n57449 );
buf ( R_56e_10086e98 , n57450 );
buf ( R_cef_14870eb8 , n57451 );
buf ( R_11ac_13c24498 , n57452 );
buf ( R_130e_14a17758 , C0 );
buf ( R_17cb_14a0e478 , n57453 );
buf ( R_192d_123becb8 , n57475 );
buf ( R_d32_13d20558 , C0 );
buf ( R_713_15882978 , n57476 );
buf ( R_b4a_13d22cb8 , C0 );
buf ( R_1169_123b7c38 , n57486 );
buf ( R_1351_14a14558 , n57497 );
buf ( R_1788_13ccae18 , n57498 );
buf ( R_1970_124c43f8 , n57499 );
buf ( R_7cd_13d58df8 , n57510 );
buf ( R_dec_156ae518 , n57511 );
buf ( R_a90_13dd8058 , n57512 );
buf ( R_10af_117f0818 , n57513 );
buf ( R_140b_1580d1b8 , n57514 );
buf ( R_16ce_117ebe58 , C0 );
buf ( R_1a2a_15810e58 , C0 );
buf ( R_e72_13c1e8b8 , C0 );
buf ( R_a0a_13d54438 , C0 );
buf ( R_853_123bd778 , n57515 );
buf ( R_1029_13cd2898 , n57523 );
buf ( R_1491_117f33d8 , n57534 );
buf ( R_1648_15ff12c8 , n57535 );
buf ( R_80f_13d449d8 , n57536 );
buf ( R_a4e_13b8e798 , C0 );
buf ( R_e2e_13dd57b8 , C0 );
buf ( R_106d_13b8b598 , n57547 );
buf ( R_144d_13cd65d8 , n57557 );
buf ( R_168c_15ff1c28 , n57558 );
buf ( n17499 , RI15b3e9d0_1);
buf ( n17500 , n17499 );
not ( n17501 , RI15b51198_632);
nor ( n17502 , n17501 , RI15b51210_633);
nor ( n17503 , RI15b51120_631 , RI15b51288_634);
and ( n17504 , n17502 , n17503 );
not ( n17505 , RI15b54690_745);
nand ( n17506 , n17504 , n17505 );
not ( n17507 , n17506 );
nand ( n17508 , RI15b56760_815 , RI15b567d8_816);
not ( n17509 , n17508 );
not ( n17510 , RI15b566e8_814);
and ( n17511 , n17509 , n17510 );
nand ( n17512 , n17507 , n17511 );
not ( n17513 , n17512 );
nand ( n17514 , RI15b570c0_835 , RI15b57138_836);
not ( n17515 , n17514 );
and ( n17516 , n17515 , RI15b571b0_837);
nand ( n17517 , n17516 , RI15b57228_838);
not ( n17518 , RI15b572a0_839);
nor ( n17519 , n17517 , n17518 );
nand ( n17520 , n17519 , RI15b57318_840);
not ( n17521 , RI15b57390_841);
nor ( n17522 , n17520 , n17521 );
nand ( n17523 , n17522 , RI15b57408_842);
not ( n17524 , n17523 );
nand ( n17525 , RI15b567d8_816 , RI15b56850_817);
not ( n17526 , RI15b568c8_818);
nor ( n17527 , n17525 , n17526 );
nand ( n17528 , n17527 , RI15b56940_819);
not ( n17529 , RI15b569b8_820);
nor ( n17530 , n17528 , n17529 );
and ( n17531 , n17530 , RI15b56a30_821);
nand ( n17532 , n17531 , RI15b56aa8_822);
not ( n17533 , RI15b56b20_823);
nor ( n17534 , n17532 , n17533 );
nand ( n17535 , n17534 , RI15b56b98_824);
not ( n17536 , RI15b56c10_825);
nor ( n17537 , n17535 , n17536 );
and ( n17538 , n17537 , RI15b56c88_826);
nand ( n17539 , n17538 , RI15b56d00_827);
not ( n17540 , RI15b56d78_828);
nor ( n17541 , n17539 , n17540 );
nand ( n17542 , n17541 , RI15b56df0_829);
not ( n17543 , RI15b56e68_830);
nor ( n17544 , n17542 , n17543 );
nand ( n17545 , n17544 , RI15b56ee0_831);
not ( n17546 , RI15b56f58_832);
nor ( n17547 , n17545 , n17546 );
nand ( n17548 , n17547 , RI15b56fd0_833);
not ( n17549 , RI15b57048_834);
nor ( n17550 , n17548 , n17549 );
nand ( n17551 , n17550 , RI15b56760_815);
not ( n17552 , n17551 );
buf ( n17553 , n17552 );
nand ( n17554 , n17524 , n17553 );
not ( n17555 , RI15b57480_843);
nor ( n17556 , n17554 , n17555 );
nand ( n17557 , n17556 , RI15b574f8_844);
not ( n17558 , RI15b57570_845);
and ( n17559 , n17557 , n17558 );
not ( n17560 , n17557 );
and ( n17561 , n17560 , RI15b57570_845);
nor ( n17562 , n17559 , n17561 );
not ( n17563 , n17562 );
nand ( n17564 , n17563 , n17507 );
buf ( n17565 , n17564 );
not ( n17566 , n17565 );
or ( n17567 , n17513 , n17566 );
not ( n17568 , n17508 );
not ( n17569 , RI15b56850_817);
and ( n17570 , n17568 , n17569 );
and ( n17571 , n17508 , RI15b56850_817);
nor ( n17572 , n17570 , n17571 );
not ( n17573 , n17572 );
nand ( n17574 , n17567 , n17573 );
nand ( n17575 , n17562 , n17507 );
buf ( n17576 , n17575 );
buf ( n17577 , n17576 );
not ( n17578 , n17577 );
nor ( n17579 , n17573 , n17511 );
nand ( n17580 , n17578 , n17579 );
not ( n17581 , RI15b4d340_499);
nor ( n17582 , RI15b50e50_625 , RI15b50ec8_626);
and ( n17583 , n17582 , RI15b50f40_627);
not ( n17584 , RI15b50fb8_628);
nand ( n17585 , n17583 , n17584 );
not ( n17586 , n17585 );
not ( n17587 , RI15b51030_629);
nand ( n17588 , n17586 , n17587 );
not ( n17589 , n17588 );
not ( n17590 , n17589 );
or ( n17591 , n17581 , n17590 );
nand ( n17592 , RI15b50ec8_626 , RI15b50f40_627);
buf ( n17593 , n17592 );
nor ( n17594 , n17593 , RI15b50e50_625);
not ( n17595 , RI15b50fb8_628);
and ( n17596 , n17594 , n17595 );
nand ( n17597 , n17596 , n17587 );
not ( n17598 , n17597 );
not ( n17599 , RI15b4dac0_515);
not ( n17600 , n17599 );
and ( n17601 , n17598 , n17600 );
not ( n17602 , RI15b50f40_627);
nand ( n17603 , n17602 , RI15b50ec8_626);
nor ( n17604 , n17603 , RI15b50e50_625);
not ( n17605 , n17604 );
not ( n17606 , RI15b50fb8_628);
nor ( n17607 , n17605 , n17606 );
nand ( n17608 , n17607 , n17587 );
not ( n17609 , n17608 );
and ( n17610 , n17609 , RI15b4e9c0_547);
nor ( n17611 , n17601 , n17610 );
nand ( n17612 , n17591 , n17611 );
not ( n17613 , RI15b4ed80_555);
not ( n17614 , n17603 );
nand ( n17615 , n17614 , RI15b50e50_625);
not ( n17616 , RI15b50fb8_628);
nor ( n17617 , n17615 , n17616 );
and ( n17618 , n17617 , n17587 );
not ( n17619 , n17618 );
or ( n17620 , n17613 , n17619 );
nand ( n17621 , RI15b50e50_625 , RI15b50ec8_626);
not ( n17622 , n17621 );
nand ( n17623 , n17622 , RI15b50f40_627);
not ( n17624 , RI15b50fb8_628);
nor ( n17625 , n17623 , n17624 );
nand ( n17626 , n17625 , n17587 );
not ( n17627 , n17626 );
nand ( n17628 , n17627 , RI15b4fc80_587);
nand ( n17629 , n17620 , n17628 );
nor ( n17630 , n17612 , n17629 );
not ( n17631 , RI15b50ec8_626);
nand ( n17632 , n17631 , RI15b50e50_625);
buf ( n17633 , n17632 );
not ( n17634 , n17633 );
not ( n17635 , RI15b50f40_627);
nand ( n17636 , n17634 , n17635 );
not ( n17637 , RI15b50fb8_628);
nor ( n17638 , n17636 , n17637 );
and ( n17639 , n17638 , n17587 );
nand ( n17640 , n17639 , RI15b4e600_539);
not ( n17641 , n17636 );
nor ( n17642 , RI15b50fb8_628 , RI15b51030_629);
nand ( n17643 , n17641 , n17642 );
not ( n17644 , n17643 );
not ( n17645 , RI15b4c800_475);
not ( n17646 , n17645 );
and ( n17647 , n17644 , n17646 );
not ( n17648 , RI15b50f40_627);
nor ( n17649 , n17633 , n17648 );
nor ( n17650 , RI15b50fb8_628 , RI15b51030_629);
and ( n17651 , n17649 , n17650 );
not ( n17652 , n17651 );
not ( n17653 , RI15b4d700_507);
nor ( n17654 , n17652 , n17653 );
nor ( n17655 , n17647 , n17654 );
not ( n17656 , RI15b50f40_627);
and ( n17657 , n17582 , n17656 );
nand ( n17658 , n17657 , n17650 );
not ( n17659 , n17658 );
not ( n17660 , RI15b4c440_467);
not ( n17661 , n17660 );
and ( n17662 , n17659 , n17661 );
nand ( n17663 , n17604 , n17650 );
not ( n17664 , RI15b4cbc0_483);
nor ( n17665 , n17663 , n17664 );
nor ( n17666 , n17662 , n17665 );
not ( n17667 , n17615 );
nand ( n17668 , n17667 , n17642 );
not ( n17669 , n17668 );
nand ( n17670 , n17669 , RI15b4cf80_491);
and ( n17671 , n17640 , n17655 , n17666 , n17670 );
and ( n17672 , n17583 , RI15b50fb8_628);
and ( n17673 , n17672 , n17587 );
and ( n17674 , n17673 , RI15b4f140_563);
and ( n17675 , n17594 , RI15b50fb8_628);
and ( n17676 , n17675 , n17587 );
not ( n17677 , n17676 );
not ( n17678 , RI15b4f8c0_579);
nor ( n17679 , n17677 , n17678 );
nor ( n17680 , n17674 , n17679 );
nand ( n17681 , n17657 , RI15b50fb8_628);
nor ( n17682 , n17681 , RI15b51030_629);
buf ( n17683 , n17682 );
nand ( n17684 , n17683 , RI15b4e240_531);
not ( n17685 , n17649 );
not ( n17686 , RI15b50fb8_628);
nor ( n17687 , n17685 , n17686 );
nand ( n17688 , n17687 , n17587 );
not ( n17689 , n17688 );
nand ( n17690 , n17689 , RI15b4f500_571);
nor ( n17691 , n17623 , RI15b50fb8_628);
nand ( n17692 , n17691 , n17587 );
not ( n17693 , n17692 );
nand ( n17694 , n17693 , RI15b4de80_523);
and ( n17695 , n17684 , n17690 , n17694 );
nand ( n17696 , n17630 , n17671 , n17680 , n17695 );
not ( n17697 , n17696 );
not ( n17698 , RI15b4d3b8_500);
not ( n17699 , n17589 );
or ( n17700 , n17698 , n17699 );
not ( n17701 , n17597 );
not ( n17702 , RI15b4db38_516);
not ( n17703 , n17702 );
and ( n17704 , n17701 , n17703 );
and ( n17705 , n17609 , RI15b4ea38_548);
nor ( n17706 , n17704 , n17705 );
nand ( n17707 , n17700 , n17706 );
not ( n17708 , RI15b4edf8_556);
not ( n17709 , n17618 );
or ( n17710 , n17708 , n17709 );
nand ( n17711 , n17627 , RI15b4fcf8_588);
nand ( n17712 , n17710 , n17711 );
nor ( n17713 , n17707 , n17712 );
nand ( n17714 , n17639 , RI15b4e678_540);
not ( n17715 , n17643 );
not ( n17716 , RI15b4c878_476);
not ( n17717 , n17716 );
and ( n17718 , n17715 , n17717 );
and ( n17719 , n17651 , RI15b4d778_508);
nor ( n17720 , n17718 , n17719 );
not ( n17721 , n17663 );
and ( n17722 , n17721 , RI15b4cc38_484);
not ( n17723 , RI15b4c4b8_468);
nor ( n17724 , n17658 , n17723 );
nor ( n17725 , n17722 , n17724 );
nand ( n17726 , n17669 , RI15b4cff8_492);
and ( n17727 , n17714 , n17720 , n17725 , n17726 );
and ( n17728 , n17673 , RI15b4f1b8_564);
not ( n17729 , RI15b4f938_580);
nor ( n17730 , n17677 , n17729 );
nor ( n17731 , n17728 , n17730 );
nand ( n17732 , n17683 , RI15b4e2b8_532);
nand ( n17733 , n17689 , RI15b4f578_572);
nand ( n17734 , n17693 , RI15b4def8_524);
and ( n17735 , n17732 , n17733 , n17734 );
nand ( n17736 , n17713 , n17727 , n17731 , n17735 );
not ( n17737 , RI15b4d598_504);
not ( n17738 , n17589 );
or ( n17739 , n17737 , n17738 );
not ( n17740 , n17597 );
not ( n17741 , RI15b4dd18_520);
not ( n17742 , n17741 );
and ( n17743 , n17740 , n17742 );
and ( n17744 , n17609 , RI15b4ec18_552);
nor ( n17745 , n17743 , n17744 );
nand ( n17746 , n17739 , n17745 );
not ( n17747 , RI15b4efd8_560);
not ( n17748 , n17618 );
or ( n17749 , n17747 , n17748 );
nand ( n17750 , n17627 , RI15b4fed8_592);
nand ( n17751 , n17749 , n17750 );
nor ( n17752 , n17746 , n17751 );
nand ( n17753 , n17639 , RI15b4e858_544);
not ( n17754 , n17643 );
not ( n17755 , RI15b4ca58_480);
not ( n17756 , n17755 );
and ( n17757 , n17754 , n17756 );
not ( n17758 , RI15b4d958_512);
nor ( n17759 , n17652 , n17758 );
nor ( n17760 , n17757 , n17759 );
not ( n17761 , n17663 );
not ( n17762 , RI15b4ce18_488);
not ( n17763 , n17762 );
and ( n17764 , n17761 , n17763 );
not ( n17765 , RI15b4c698_472);
nor ( n17766 , n17658 , n17765 );
nor ( n17767 , n17764 , n17766 );
nand ( n17768 , n17669 , RI15b4d1d8_496);
and ( n17769 , n17753 , n17760 , n17767 , n17768 );
not ( n17770 , n17672 );
nor ( n17771 , n17770 , RI15b51030_629);
not ( n17772 , n17771 );
not ( n17773 , n17772 );
not ( n17774 , RI15b4f398_568);
not ( n17775 , n17774 );
and ( n17776 , n17773 , n17775 );
and ( n17777 , n17676 , RI15b4fb18_584);
nor ( n17778 , n17776 , n17777 );
nand ( n17779 , n17683 , RI15b4e498_536);
not ( n17780 , n17688 );
nand ( n17781 , n17780 , RI15b4f758_576);
nand ( n17782 , n17693 , RI15b4e0d8_528);
and ( n17783 , n17779 , n17781 , n17782 );
nand ( n17784 , n17752 , n17769 , n17778 , n17783 );
and ( n17785 , n17697 , n17736 , n17784 );
not ( n17786 , RI15b4d4a8_502);
not ( n17787 , n17589 );
or ( n17788 , n17786 , n17787 );
not ( n17789 , n17597 );
not ( n17790 , RI15b4dc28_518);
not ( n17791 , n17790 );
and ( n17792 , n17789 , n17791 );
and ( n17793 , n17609 , RI15b4eb28_550);
nor ( n17794 , n17792 , n17793 );
nand ( n17795 , n17788 , n17794 );
not ( n17796 , RI15b4eee8_558);
not ( n17797 , n17618 );
or ( n17798 , n17796 , n17797 );
nand ( n17799 , n17627 , RI15b4fde8_590);
nand ( n17800 , n17798 , n17799 );
nor ( n17801 , n17795 , n17800 );
not ( n17802 , n17643 );
not ( n17803 , RI15b4c968_478);
not ( n17804 , n17803 );
and ( n17805 , n17802 , n17804 );
not ( n17806 , RI15b4d868_510);
nor ( n17807 , n17652 , n17806 );
nor ( n17808 , n17805 , n17807 );
not ( n17809 , n17663 );
not ( n17810 , RI15b4cd28_486);
not ( n17811 , n17810 );
and ( n17812 , n17809 , n17811 );
not ( n17813 , RI15b4c5a8_470);
nor ( n17814 , n17658 , n17813 );
nor ( n17815 , n17812 , n17814 );
nand ( n17816 , n17669 , RI15b4d0e8_494);
nand ( n17817 , n17808 , n17815 , n17816 );
not ( n17818 , n17639 );
not ( n17819 , RI15b4e768_542);
nor ( n17820 , n17818 , n17819 );
nor ( n17821 , n17817 , n17820 );
and ( n17822 , n17771 , RI15b4f2a8_566);
and ( n17823 , n17676 , RI15b4fa28_582);
nor ( n17824 , n17822 , n17823 );
and ( n17825 , n17683 , RI15b4e3a8_534);
not ( n17826 , RI15b4f668_574);
not ( n17827 , n17689 );
or ( n17828 , n17826 , n17827 );
nand ( n17829 , n17693 , RI15b4dfe8_526);
nand ( n17830 , n17828 , n17829 );
nor ( n17831 , n17825 , n17830 );
nand ( n17832 , n17801 , n17821 , n17824 , n17831 );
not ( n17833 , n17832 );
not ( n17834 , RI15b4d430_501);
not ( n17835 , n17589 );
or ( n17836 , n17834 , n17835 );
not ( n17837 , n17597 );
not ( n17838 , RI15b4dbb0_517);
not ( n17839 , n17838 );
and ( n17840 , n17837 , n17839 );
and ( n17841 , n17609 , RI15b4eab0_549);
nor ( n17842 , n17840 , n17841 );
nand ( n17843 , n17836 , n17842 );
not ( n17844 , RI15b4ee70_557);
not ( n17845 , n17618 );
or ( n17846 , n17844 , n17845 );
nand ( n17847 , n17627 , RI15b4fd70_589);
nand ( n17848 , n17846 , n17847 );
nor ( n17849 , n17843 , n17848 );
not ( n17850 , RI15b4c8f0_477);
not ( n17851 , n17643 );
not ( n17852 , n17851 );
or ( n17853 , n17850 , n17852 );
nand ( n17854 , n17651 , RI15b4d7f0_509);
nand ( n17855 , n17853 , n17854 );
not ( n17856 , RI15b4d070_493);
nor ( n17857 , n17668 , n17856 );
nor ( n17858 , n17855 , n17857 );
nand ( n17859 , n17639 , RI15b4e6f0_541);
not ( n17860 , RI15b4c530_469);
nor ( n17861 , n17658 , n17860 );
not ( n17862 , RI15b4ccb0_485);
nor ( n17863 , n17663 , n17862 );
nor ( n17864 , n17861 , n17863 );
and ( n17865 , n17858 , n17859 , n17864 );
and ( n17866 , n17673 , RI15b4f230_565);
not ( n17867 , RI15b4f9b0_581);
nor ( n17868 , n17677 , n17867 );
nor ( n17869 , n17866 , n17868 );
and ( n17870 , n17683 , RI15b4e330_533);
not ( n17871 , RI15b4f5f0_573);
not ( n17872 , n17689 );
or ( n17873 , n17871 , n17872 );
nand ( n17874 , n17693 , RI15b4df70_525);
nand ( n17875 , n17873 , n17874 );
nor ( n17876 , n17870 , n17875 );
nand ( n17877 , n17849 , n17865 , n17869 , n17876 );
not ( n17878 , n17877 );
not ( n17879 , RI15b4d520_503);
not ( n17880 , n17589 );
or ( n17881 , n17879 , n17880 );
not ( n17882 , n17597 );
not ( n17883 , RI15b4dca0_519);
not ( n17884 , n17883 );
and ( n17885 , n17882 , n17884 );
and ( n17886 , n17609 , RI15b4eba0_551);
nor ( n17887 , n17885 , n17886 );
nand ( n17888 , n17881 , n17887 );
not ( n17889 , RI15b4ef60_559);
not ( n17890 , n17618 );
or ( n17891 , n17889 , n17890 );
nand ( n17892 , n17627 , RI15b4fe60_591);
nand ( n17893 , n17891 , n17892 );
nor ( n17894 , n17888 , n17893 );
nand ( n17895 , n17639 , RI15b4e7e0_543);
not ( n17896 , n17643 );
not ( n17897 , RI15b4c9e0_479);
not ( n17898 , n17897 );
and ( n17899 , n17896 , n17898 );
not ( n17900 , RI15b4d8e0_511);
nor ( n17901 , n17652 , n17900 );
nor ( n17902 , n17899 , n17901 );
and ( n17903 , n17721 , RI15b4cda0_487);
not ( n17904 , RI15b4c620_471);
nor ( n17905 , n17658 , n17904 );
nor ( n17906 , n17903 , n17905 );
nand ( n17907 , n17669 , RI15b4d160_495);
and ( n17908 , n17895 , n17902 , n17906 , n17907 );
and ( n17909 , n17771 , RI15b4f320_567);
and ( n17910 , n17676 , RI15b4faa0_583);
nor ( n17911 , n17909 , n17910 );
nand ( n17912 , n17683 , RI15b4e420_535);
nand ( n17913 , n17689 , RI15b4f6e0_575);
nand ( n17914 , n17693 , RI15b4e060_527);
and ( n17915 , n17912 , n17913 , n17914 );
nand ( n17916 , n17894 , n17908 , n17911 , n17915 );
not ( n17917 , n17916 );
and ( n17918 , n17833 , n17878 , n17917 );
nand ( n17919 , n17851 , RI15b4c788_474);
nand ( n17920 , n17669 , RI15b4cf08_490);
nand ( n17921 , n17651 , RI15b4d688_506);
nand ( n17922 , n17919 , n17920 , n17921 );
not ( n17923 , RI15b4c3c8_466);
not ( n17924 , n17658 );
not ( n17925 , n17924 );
or ( n17926 , n17923 , n17925 );
nand ( n17927 , n17721 , RI15b4cb48_482);
nand ( n17928 , n17926 , n17927 );
nor ( n17929 , n17922 , n17928 );
nand ( n17930 , n17771 , RI15b4f0c8_562);
nand ( n17931 , n17639 , RI15b4e588_538);
nand ( n17932 , n17676 , RI15b4f848_578);
nand ( n17933 , n17929 , n17930 , n17931 , n17932 );
and ( n17934 , n17689 , RI15b4f488_570);
and ( n17935 , n17693 , RI15b4de08_522);
nor ( n17936 , n17934 , n17935 );
nand ( n17937 , n17683 , RI15b4e1c8_530);
nand ( n17938 , n17936 , n17937 );
nor ( n17939 , n17933 , n17938 );
and ( n17940 , n17589 , RI15b4d2c8_498);
not ( n17941 , RI15b4ed08_554);
not ( n17942 , n17618 );
or ( n17943 , n17941 , n17942 );
nand ( n17944 , n17627 , RI15b4fc08_586);
nand ( n17945 , n17943 , n17944 );
not ( n17946 , n17608 );
nand ( n17947 , n17946 , RI15b4e948_546);
not ( n17948 , n17597 );
nand ( n17949 , n17948 , RI15b4da48_514);
nand ( n17950 , n17947 , n17949 );
nor ( n17951 , n17940 , n17945 , n17950 );
nand ( n17952 , n17939 , n17951 );
not ( n17953 , RI15b4d250_497);
not ( n17954 , n17589 );
or ( n17955 , n17953 , n17954 );
not ( n17956 , n17597 );
not ( n17957 , RI15b4d9d0_513);
not ( n17958 , n17957 );
and ( n17959 , n17956 , n17958 );
and ( n17960 , n17609 , RI15b4e8d0_545);
nor ( n17961 , n17959 , n17960 );
nand ( n17962 , n17955 , n17961 );
not ( n17963 , RI15b4ec90_553);
not ( n17964 , n17618 );
or ( n17965 , n17963 , n17964 );
nand ( n17966 , n17627 , RI15b4fb90_585);
nand ( n17967 , n17965 , n17966 );
nor ( n17968 , n17962 , n17967 );
nand ( n17969 , n17639 , RI15b4e510_537);
not ( n17970 , n17643 );
not ( n17971 , RI15b4c710_473);
not ( n17972 , n17971 );
and ( n17973 , n17970 , n17972 );
not ( n17974 , RI15b4d610_505);
nor ( n17975 , n17652 , n17974 );
nor ( n17976 , n17973 , n17975 );
and ( n17977 , n17721 , RI15b4cad0_481);
not ( n17978 , RI15b4c350_465);
nor ( n17979 , n17658 , n17978 );
nor ( n17980 , n17977 , n17979 );
nand ( n17981 , n17669 , RI15b4ce90_489);
and ( n17982 , n17969 , n17976 , n17980 , n17981 );
and ( n17983 , n17673 , RI15b4f050_561);
not ( n17984 , RI15b4f7d0_577);
nor ( n17985 , n17677 , n17984 );
nor ( n17986 , n17983 , n17985 );
nand ( n17987 , n17683 , RI15b4e150_529);
nand ( n17988 , n17689 , RI15b4f410_569);
nand ( n17989 , n17693 , RI15b4dd90_521);
and ( n17990 , n17987 , n17988 , n17989 );
nand ( n17991 , n17968 , n17982 , n17986 , n17990 );
nand ( n17992 , n17952 , n17991 );
not ( n17993 , n17992 );
and ( n17994 , n17785 , n17918 , n17993 );
buf ( n17995 , n17642 );
not ( n17996 , n17995 );
not ( n17997 , n17996 );
not ( n17998 , RI15b4c1e8_462);
nand ( n17999 , n17998 , RI15b50f40_627);
not ( n18000 , n17999 );
nor ( n18001 , RI15b4c0f8_460 , RI15b4c170_461);
or ( n18002 , n18001 , RI15b50ec8_626);
not ( n18003 , n17582 );
not ( n18004 , RI15b50e50_625);
nand ( n18005 , n18004 , RI15b4c170_461);
nand ( n18006 , RI15b4c0f8_460 , RI15b4c170_461);
buf ( n18007 , n18006 );
nand ( n18008 , n18002 , n18003 , n18005 , n18007 );
not ( n18009 , n18008 );
or ( n18010 , n18000 , n18009 );
not ( n18011 , RI15b50f40_627);
nand ( n18012 , n18011 , RI15b4c1e8_462);
nand ( n18013 , n18010 , n18012 );
nand ( n18014 , n18013 , RI15b4c260_463);
not ( n18015 , n18014 );
nand ( n18016 , n18015 , RI15b50fb8_628 , RI15b51030_629);
not ( n18017 , n18016 );
nor ( n18018 , n18013 , RI15b4c260_463);
not ( n18019 , n18018 );
not ( n18020 , RI15b50fb8_628);
nand ( n18021 , n18019 , n18014 , n18020 );
not ( n18022 , n18021 );
or ( n18023 , n18017 , n18022 );
nand ( n18024 , n18023 , RI15b4c2d8_464);
nand ( n18025 , n18018 , n17587 , RI15b50fb8_628);
nand ( n18026 , n18024 , n18025 );
not ( n18027 , n18026 );
or ( n18028 , n17997 , n18027 );
not ( n18029 , RI15b50fb8_628);
not ( n18030 , n18018 );
nand ( n18031 , n18030 , n18014 );
not ( n18032 , n18031 );
or ( n18033 , n18029 , n18032 );
nand ( n18034 , n18033 , n18021 );
nor ( n18035 , RI15b4c2d8_464 , RI15b51030_629);
and ( n18036 , n18034 , n18035 );
not ( n18037 , RI15b4c2d8_464);
or ( n18038 , n18018 , RI15b50fb8_628);
nand ( n18039 , n18038 , n18014 , RI15b51030_629);
not ( n18040 , n18039 );
or ( n18041 , n18037 , n18040 );
not ( n18042 , n18018 );
not ( n18043 , n17995 );
not ( n18044 , n18043 );
and ( n18045 , n18042 , n18044 );
nor ( n18046 , n18014 , RI15b51030_629);
nor ( n18047 , n18045 , n18046 );
nand ( n18048 , n18041 , n18047 );
not ( n18049 , n18048 );
nor ( n18050 , n18036 , n18049 );
nand ( n18051 , n18028 , n18050 );
and ( n18052 , n18012 , n17999 );
and ( n18053 , n18008 , n18052 );
nor ( n18054 , n18008 , n18052 );
nor ( n18055 , n18053 , n18054 );
nand ( n18056 , n18048 , n18055 );
not ( n18057 , RI15b4c0f8_460);
and ( n18058 , n18057 , RI15b50e50_625);
not ( n18059 , n18058 );
not ( n18060 , RI15b50ec8_626);
and ( n18061 , n18060 , RI15b4c170_461);
not ( n18062 , RI15b4c170_461);
and ( n18063 , n18062 , RI15b50ec8_626);
nor ( n18064 , n18061 , n18063 );
not ( n18065 , n18064 );
or ( n18066 , n18059 , n18065 );
or ( n18067 , n18064 , n18058 );
nand ( n18068 , n18066 , n18067 );
nand ( n18069 , n18048 , n18068 );
and ( n18070 , n18056 , n18069 );
nand ( n18071 , n18051 , n18070 );
nand ( n18072 , RI15b667c8_1362 , RI15b66840_1363);
nand ( n18073 , n18072 , n17505 );
nand ( n18074 , n17994 , n18071 , n18073 );
not ( n18075 , RI15b51288_634);
and ( n18076 , n18075 , RI15b51210_633);
and ( n18077 , n18076 , n17501 , RI15b51120_631);
not ( n18078 , n18077 );
or ( n18079 , n18074 , n18078 );
nor ( n18080 , RI15b557e8_782 , RI15b55860_783);
not ( n18081 , RI15b558d8_784);
nand ( n18082 , n18080 , n18081 );
or ( n18083 , n18079 , n18082 );
not ( n18084 , RI15b56670_813);
not ( n18085 , n18084 );
not ( n18086 , n18079 );
not ( n18087 , n18086 );
or ( n18088 , n18085 , n18087 );
not ( n18089 , n17991 );
nor ( n18090 , n18089 , n17952 );
nand ( n18091 , n17785 , n17918 , n18090 );
and ( n18092 , RI15b547f8_748 , RI15b54870_749);
or ( n18093 , RI15b547f8_748 , RI15b54870_749);
not ( n18094 , RI15b54780_747);
nand ( n18095 , n18093 , n18094 );
nor ( n18096 , n18092 , n18095 );
nand ( n18097 , n18096 , n18072 );
nor ( n18098 , n18097 , RI15b54690_745);
nor ( n18099 , n18091 , n18098 );
and ( n18100 , n18071 , n18077 );
buf ( n18101 , n18100 );
nand ( n18102 , n18099 , n18101 );
nand ( n18103 , n18088 , n18102 );
not ( n18104 , n18103 );
nand ( n18105 , n18083 , n18104 );
and ( n18106 , n18105 , RI15b55950_785);
not ( n18107 , n17833 );
nand ( n18108 , n17785 , n18107 );
not ( n18109 , n18108 );
not ( n18110 , n17917 );
nor ( n18111 , n17878 , n18110 );
nand ( n18112 , n18109 , n18111 );
not ( n18113 , n17952 );
and ( n18114 , n18089 , n18113 );
nor ( n18115 , n17993 , n18114 );
nor ( n18116 , n18112 , n18115 );
not ( n18117 , n17877 );
and ( n18118 , n18117 , n17916 );
and ( n18119 , n18090 , n18118 );
nand ( n18120 , n18109 , n18119 );
not ( n18121 , n18120 );
nor ( n18122 , n18116 , n18121 );
not ( n18123 , n17736 );
and ( n18124 , n18123 , n17697 , n17833 );
buf ( n18125 , n18110 );
nand ( n18126 , n18124 , n18114 , n17784 , n18125 );
nand ( n18127 , n18122 , n18126 );
not ( n18128 , n18118 );
nor ( n18129 , n18128 , n17992 );
nand ( n18130 , n18109 , n18129 );
not ( n18131 , n18130 );
nor ( n18132 , n18127 , n18131 );
not ( n18133 , n17994 );
and ( n18134 , n18123 , n17696 , n18089 );
and ( n18135 , n17784 , n17832 );
and ( n18136 , n18134 , n18135 , n18118 );
buf ( n18137 , n17952 );
not ( n18138 , n18137 );
nand ( n18139 , n18136 , n18138 );
nand ( n18140 , n18133 , n18139 );
nand ( n18141 , n18136 , n18137 );
nand ( n18142 , n18091 , n18141 );
nor ( n18143 , n18140 , n18142 );
buf ( n18144 , n18143 );
not ( n18145 , n18144 );
buf ( n18146 , n18071 );
not ( n18147 , n18146 );
buf ( n18148 , n18147 );
not ( n18149 , n18148 );
nand ( n18150 , n18132 , n18145 , n18149 );
nand ( n18151 , n18150 , n18077 );
nor ( n18152 , RI15b51198_632 , RI15b51210_633);
not ( n18153 , n18152 );
or ( n18154 , n18153 , n18075 , RI15b51120_631);
not ( n18155 , n18154 );
and ( n18156 , n18076 , RI15b51120_631 , RI15b51198_632);
nor ( n18157 , n18155 , n18156 );
not ( n18158 , n18152 );
not ( n18159 , n18075 );
and ( n18160 , n18158 , n18159 );
and ( n18161 , n18152 , n18075 );
nor ( n18162 , n18160 , n18161 );
not ( n18163 , n18162 );
nand ( n18164 , n18163 , RI15b51120_631);
nand ( n18165 , n17502 , n18075 , RI15b51120_631);
not ( n18166 , RI15b51120_631);
nand ( n18167 , n18076 , n18166 , RI15b51198_632);
nand ( n18168 , n18165 , n18167 );
not ( n18169 , n18168 );
and ( n18170 , n18076 , n17501 , n18166 );
not ( n18171 , n18170 );
nand ( n18172 , n18157 , n18164 , n18169 , n18171 );
buf ( n18173 , n17504 );
buf ( n18174 , n18173 );
not ( n18175 , n18174 );
nor ( n18176 , n18175 , n17505 );
or ( n18177 , n18172 , n18176 );
not ( n18178 , n18177 );
nand ( n18179 , n18151 , n18178 );
and ( n18180 , n18179 , RI15b57750_849);
nand ( n18181 , n18071 , n18072 );
not ( n18182 , n18181 );
buf ( n18183 , n17994 );
nand ( n18184 , n18182 , n18183 , n17505 );
not ( n18185 , n18091 );
nand ( n18186 , n18185 , n18146 , n18098 );
nand ( n18187 , n18184 , n18186 );
and ( n18188 , n18187 , n18077 );
not ( n18189 , n18188 );
nand ( n18190 , RI15b57660_847 , RI15b576d8_848);
not ( n18191 , n18190 );
not ( n18192 , RI15b57750_849);
and ( n18193 , n18191 , n18192 );
and ( n18194 , n18190 , RI15b57750_849);
nor ( n18195 , n18193 , n18194 );
or ( n18196 , n18189 , n18195 );
or ( n18197 , n18079 , n18084 );
not ( n18198 , n18197 );
not ( n18199 , n18082 );
nor ( n18200 , n18199 , RI15b55950_785);
and ( n18201 , n18198 , n18200 );
not ( n18202 , n18101 );
not ( n18203 , n18136 );
nor ( n18204 , n18202 , n18203 );
not ( n18205 , n17592 );
nand ( n18206 , n18205 , RI15b50e50_625);
not ( n18207 , RI15b50fb8_628);
and ( n18208 , n18206 , n18207 );
not ( n18209 , n18206 );
and ( n18210 , n18209 , RI15b50fb8_628);
nor ( n18211 , n18208 , n18210 );
not ( n18212 , n18211 );
not ( n18213 , n18212 );
buf ( n18214 , n18213 );
buf ( n18215 , n18214 );
and ( n18216 , n18204 , n18215 );
nand ( n18217 , RI15b51120_631 , RI15b51288_634);
or ( n18218 , n18153 , n18217 );
not ( n18219 , n18218 );
and ( n18220 , n18219 , RI15b56850_817);
nor ( n18221 , n18201 , n18216 , n18220 );
nand ( n18222 , n18196 , n18221 );
nor ( n18223 , n18106 , n18180 , n18222 );
nand ( n18224 , n17574 , n17580 , n18223 );
buf ( n18225 , n18224 );
buf ( n18226 , RI15b3ea48_2);
buf ( n18227 , n18226 );
nand ( n18228 , RI15b5c4a8_1014 , RI15b5c520_1015);
not ( n18229 , RI15b5c598_1016);
nor ( n18230 , n18228 , n18229 );
nand ( n18231 , n18230 , RI15b5c430_1013);
not ( n18232 , RI15b5c610_1017);
nor ( n18233 , n18231 , n18232 );
nand ( n18234 , n18233 , RI15b5c688_1018);
not ( n18235 , RI15b5c700_1019);
nor ( n18236 , n18234 , n18235 );
not ( n18237 , n18236 );
not ( n18238 , RI15b5c778_1020);
not ( n18239 , n18238 );
and ( n18240 , n18237 , n18239 );
and ( n18241 , n18236 , n18238 );
nor ( n18242 , n18240 , n18241 );
not ( n18243 , n18242 );
not ( n18244 , RI15b5d2b8_1044);
nand ( n18245 , n18244 , RI15b5d330_1045);
not ( n18246 , RI15b5d330_1045);
nand ( n18247 , n18246 , RI15b5d2b8_1044);
nand ( n18248 , n18245 , n18247 );
not ( n18249 , RI15b5d2b8_1044);
and ( n18250 , n18248 , n18249 );
not ( n18251 , RI15b5d420_1047);
nand ( n18252 , RI15b5d2b8_1044 , RI15b5d330_1045);
not ( n18253 , n18252 );
nand ( n18254 , n18253 , RI15b5d3a8_1046);
not ( n18255 , n18254 );
or ( n18256 , n18251 , n18255 );
not ( n18257 , RI15b5d420_1047);
nand ( n18258 , n18257 , RI15b5d3a8_1046);
nor ( n18259 , n18252 , n18258 );
not ( n18260 , n18259 );
nand ( n18261 , n18256 , n18260 );
buf ( n18262 , n18261 );
not ( n18263 , RI15b5d3a8_1046);
nand ( n18264 , RI15b5d2b8_1044 , RI15b5d330_1045);
not ( n18265 , n18264 );
or ( n18266 , n18263 , n18265 );
not ( n18267 , n18264 );
not ( n18268 , RI15b5d3a8_1046);
nand ( n18269 , n18267 , n18268 );
nand ( n18270 , n18266 , n18269 );
not ( n18271 , n18270 );
and ( n18272 , n18250 , n18262 , n18271 );
buf ( n18273 , n18272 );
and ( n18274 , n18273 , RI15b5b440_979);
nand ( n18275 , n18248 , RI15b5d2b8_1044);
not ( n18276 , n18275 );
and ( n18277 , n18276 , n18262 , n18271 );
buf ( n18278 , n18277 );
and ( n18279 , n18278 , RI15b5b080_971);
nor ( n18280 , n18274 , n18279 );
not ( n18281 , n18248 );
nand ( n18282 , n18281 , RI15b5d2b8_1044);
not ( n18283 , n18282 );
nand ( n18284 , n18283 , n18262 , n18271 );
not ( n18285 , n18284 );
buf ( n18286 , n18285 );
and ( n18287 , n18286 , RI15b5a900_955);
not ( n18288 , n18248 );
and ( n18289 , n18288 , n18249 );
not ( n18290 , n18289 );
not ( n18291 , n18270 );
not ( n18292 , n18291 );
nor ( n18293 , n18290 , n18292 );
nand ( n18294 , n18293 , n18262 );
not ( n18295 , RI15b5acc0_963);
nor ( n18296 , n18294 , n18295 );
nor ( n18297 , n18287 , n18296 );
nand ( n18298 , n18280 , n18297 );
not ( n18299 , n18282 );
and ( n18300 , n18262 , n18299 , n18292 );
and ( n18301 , n18300 , RI15b5b800_987);
not ( n18302 , RI15b5d330_1045);
nand ( n18303 , n18302 , RI15b5d3a8_1046);
nor ( n18304 , n18303 , RI15b5d2b8_1044);
nand ( n18305 , n18262 , n18304 );
buf ( n18306 , n18305 );
not ( n18307 , n18306 );
and ( n18308 , n18307 , RI15b5bbc0_995);
nor ( n18309 , n18301 , n18308 );
not ( n18310 , n18270 );
not ( n18311 , n18310 );
and ( n18312 , n18276 , n18262 , n18311 );
buf ( n18313 , n18312 );
nand ( n18314 , n18313 , RI15b5bf80_1003);
not ( n18315 , n18291 );
and ( n18316 , n18250 , n18262 , n18315 );
buf ( n18317 , n18316 );
nand ( n18318 , n18317 , RI15b5c340_1011);
nand ( n18319 , n18309 , n18314 , n18318 );
nor ( n18320 , n18298 , n18319 );
not ( n18321 , n18282 );
not ( n18322 , n18254 );
not ( n18323 , n18322 );
not ( n18324 , RI15b5d420_1047);
not ( n18325 , n18324 );
and ( n18326 , n18323 , n18325 );
nor ( n18327 , n18326 , n18259 );
buf ( n18328 , n18327 );
and ( n18329 , n18321 , n18328 , n18315 );
buf ( n18330 , n18329 );
and ( n18331 , n18330 , RI15b59a00_923);
buf ( n18332 , n18327 );
nand ( n18333 , n18332 , n18304 );
buf ( n18334 , n18333 );
not ( n18335 , n18334 );
and ( n18336 , n18335 , RI15b59dc0_931);
nor ( n18337 , n18331 , n18336 );
not ( n18338 , n18275 );
and ( n18339 , n18338 , n18332 , n18270 );
not ( n18340 , n18339 );
not ( n18341 , n18340 );
nand ( n18342 , n18341 , RI15b5a180_939);
and ( n18343 , n18250 , n18328 , n18311 );
not ( n18344 , n18343 );
not ( n18345 , n18344 );
nand ( n18346 , n18345 , RI15b5a540_947);
nand ( n18347 , n18337 , n18342 , n18346 );
not ( n18348 , n18270 );
and ( n18349 , n18250 , n18328 , n18348 );
not ( n18350 , n18349 );
not ( n18351 , n18350 );
nand ( n18352 , n18351 , RI15b59640_915);
and ( n18353 , n18276 , n18328 , n18271 );
not ( n18354 , n18353 );
not ( n18355 , n18354 );
nand ( n18356 , n18355 , RI15b59280_907);
not ( n18357 , n18282 );
and ( n18358 , n18357 , n18332 , n18291 );
not ( n18359 , n18358 );
not ( n18360 , n18359 );
nand ( n18361 , n18360 , RI15b58b00_891);
and ( n18362 , n18332 , n18289 , n18310 );
nand ( n18363 , n18362 , RI15b58ec0_899);
nand ( n18364 , n18352 , n18356 , n18361 , n18363 );
nor ( n18365 , n18347 , n18364 );
nand ( n18366 , n18320 , n18365 );
not ( n18367 , n18366 );
and ( n18368 , n18234 , n18235 );
not ( n18369 , n18234 );
and ( n18370 , n18369 , RI15b5c700_1019);
nor ( n18371 , n18368 , n18370 );
not ( n18372 , n18371 );
nand ( n18373 , n18367 , n18372 );
not ( n18374 , n18373 );
not ( n18375 , n18338 );
not ( n18376 , n18375 );
not ( n18377 , n18292 );
nand ( n18378 , n18376 , n18262 , n18377 );
not ( n18379 , n18378 );
not ( n18380 , RI15b5b008_970);
not ( n18381 , n18380 );
and ( n18382 , n18379 , n18381 );
not ( n18383 , n18250 );
not ( n18384 , n18383 );
not ( n18385 , n18271 );
not ( n18386 , n18385 );
nand ( n18387 , n18384 , n18262 , n18386 );
not ( n18388 , RI15b5b3c8_978);
nor ( n18389 , n18387 , n18388 );
nor ( n18390 , n18382 , n18389 );
buf ( n18391 , n18343 );
and ( n18392 , n18391 , RI15b5a4c8_946);
and ( n18393 , n18341 , RI15b5a108_938);
nor ( n18394 , n18392 , n18393 );
not ( n18395 , n18286 );
not ( n18396 , n18395 );
not ( n18397 , RI15b5a888_954);
not ( n18398 , n18397 );
and ( n18399 , n18396 , n18398 );
not ( n18400 , RI15b5ac48_962);
nor ( n18401 , n18294 , n18400 );
nor ( n18402 , n18399 , n18401 );
and ( n18403 , n18330 , RI15b59988_922);
and ( n18404 , n18335 , RI15b59d48_930);
nor ( n18405 , n18403 , n18404 );
nand ( n18406 , n18390 , n18394 , n18402 , n18405 );
not ( n18407 , n18375 );
nand ( n18408 , n18407 , n18262 , n18385 );
not ( n18409 , n18408 );
not ( n18410 , RI15b5bf08_1002);
not ( n18411 , n18410 );
and ( n18412 , n18409 , n18411 );
and ( n18413 , n18317 , RI15b5c2c8_1010);
nor ( n18414 , n18412 , n18413 );
not ( n18415 , n18351 );
not ( n18416 , n18415 );
not ( n18417 , RI15b595c8_914);
not ( n18418 , n18417 );
and ( n18419 , n18416 , n18418 );
not ( n18420 , RI15b59208_906);
nor ( n18421 , n18354 , n18420 );
nor ( n18422 , n18419 , n18421 );
not ( n18423 , n18360 );
not ( n18424 , n18423 );
not ( n18425 , RI15b58a88_890);
not ( n18426 , n18425 );
and ( n18427 , n18424 , n18426 );
not ( n18428 , n18362 );
not ( n18429 , RI15b58e48_898);
nor ( n18430 , n18428 , n18429 );
nor ( n18431 , n18427 , n18430 );
and ( n18432 , n18300 , RI15b5b788_986);
and ( n18433 , n18307 , RI15b5bb48_994);
nor ( n18434 , n18432 , n18433 );
nand ( n18435 , n18414 , n18422 , n18431 , n18434 );
nor ( n18436 , n18406 , n18435 );
buf ( n18437 , n18436 );
and ( n18438 , n18233 , RI15b5c688_1018);
not ( n18439 , n18233 );
not ( n18440 , RI15b5c688_1018);
and ( n18441 , n18439 , n18440 );
nor ( n18442 , n18438 , n18441 );
not ( n18443 , n18442 );
nand ( n18444 , n18437 , n18443 );
not ( n18445 , n18444 );
not ( n18446 , RI15b5c430_1013);
nor ( n18447 , n18446 , n18228 );
and ( n18448 , n18447 , RI15b5c598_1016);
not ( n18449 , n18447 );
and ( n18450 , n18449 , n18229 );
nor ( n18451 , n18448 , n18450 );
not ( n18452 , n18451 );
not ( n18453 , RI15b5be18_1000);
nor ( n18454 , n18408 , n18453 );
not ( n18455 , n18383 );
nand ( n18456 , n18455 , n18262 , n18292 );
not ( n18457 , RI15b5c1d8_1008);
nor ( n18458 , n18456 , n18457 );
nor ( n18459 , n18454 , n18458 );
not ( n18460 , n18353 );
not ( n18461 , RI15b59118_904);
nor ( n18462 , n18460 , n18461 );
not ( n18463 , RI15b594d8_912);
nor ( n18464 , n18350 , n18463 );
nor ( n18465 , n18462 , n18464 );
not ( n18466 , n18285 );
not ( n18467 , n18466 );
not ( n18468 , RI15b5a798_952);
not ( n18469 , n18468 );
and ( n18470 , n18467 , n18469 );
not ( n18471 , RI15b5ab58_960);
nor ( n18472 , n18294 , n18471 );
nor ( n18473 , n18470 , n18472 );
and ( n18474 , n18329 , RI15b59898_920);
not ( n18475 , RI15b59c58_928);
nor ( n18476 , n18334 , n18475 );
nor ( n18477 , n18474 , n18476 );
nand ( n18478 , n18459 , n18465 , n18473 , n18477 );
not ( n18479 , n18387 );
not ( n18480 , RI15b5b2d8_976);
not ( n18481 , n18480 );
and ( n18482 , n18479 , n18481 );
not ( n18483 , RI15b5af18_968);
nor ( n18484 , n18378 , n18483 );
nor ( n18485 , n18482 , n18484 );
not ( n18486 , n18343 );
not ( n18487 , n18486 );
not ( n18488 , RI15b5a3d8_944);
not ( n18489 , n18488 );
and ( n18490 , n18487 , n18489 );
not ( n18491 , n18339 );
not ( n18492 , RI15b5a018_936);
nor ( n18493 , n18491 , n18492 );
nor ( n18494 , n18490 , n18493 );
not ( n18495 , n18359 );
not ( n18496 , RI15b58998_888);
not ( n18497 , n18496 );
and ( n18498 , n18495 , n18497 );
not ( n18499 , RI15b58d58_896);
nor ( n18500 , n18428 , n18499 );
nor ( n18501 , n18498 , n18500 );
and ( n18502 , n18321 , n18262 , n18311 );
and ( n18503 , n18502 , RI15b5b698_984);
not ( n18504 , RI15b5ba58_992);
nor ( n18505 , n18306 , n18504 );
nor ( n18506 , n18503 , n18505 );
nand ( n18507 , n18485 , n18494 , n18501 , n18506 );
nor ( n18508 , n18478 , n18507 );
buf ( n18509 , n18508 );
nand ( n18510 , n18452 , n18509 );
not ( n18511 , n18510 );
and ( n18512 , n18330 , RI15b59820_919);
not ( n18513 , RI15b59be0_927);
nor ( n18514 , n18334 , n18513 );
nor ( n18515 , n18512 , n18514 );
nand ( n18516 , n18273 , RI15b5b260_975);
nand ( n18517 , n18278 , RI15b5aea0_967);
nand ( n18518 , n18515 , n18516 , n18517 );
and ( n18519 , n18391 , RI15b5a360_943);
and ( n18520 , n18341 , RI15b59fa0_935);
nor ( n18521 , n18519 , n18520 );
and ( n18522 , n18286 , RI15b5a720_951);
not ( n18523 , RI15b5aae0_959);
nor ( n18524 , n18294 , n18523 );
nor ( n18525 , n18522 , n18524 );
nand ( n18526 , n18521 , n18525 );
nor ( n18527 , n18518 , n18526 );
and ( n18528 , n18360 , RI15b58920_887);
not ( n18529 , RI15b58ce0_895);
nor ( n18530 , n18428 , n18529 );
nor ( n18531 , n18528 , n18530 );
nand ( n18532 , n18317 , RI15b5c160_1007);
nand ( n18533 , n18313 , RI15b5bda0_999);
nand ( n18534 , n18531 , n18532 , n18533 );
and ( n18535 , n18300 , RI15b5b620_983);
not ( n18536 , n18306 );
and ( n18537 , n18536 , RI15b5b9e0_991);
nor ( n18538 , n18535 , n18537 );
nand ( n18539 , n18351 , RI15b59460_911);
nand ( n18540 , n18353 , RI15b590a0_903);
nand ( n18541 , n18538 , n18539 , n18540 );
nor ( n18542 , n18534 , n18541 );
nand ( n18543 , n18527 , n18542 );
not ( n18544 , n18543 );
nand ( n18545 , RI15b5c430_1013 , RI15b5c4a8_1014);
not ( n18546 , RI15b5c520_1015);
and ( n18547 , n18545 , n18546 );
not ( n18548 , n18545 );
and ( n18549 , n18548 , RI15b5c520_1015);
nor ( n18550 , n18547 , n18549 );
not ( n18551 , n18550 );
nand ( n18552 , n18544 , n18551 );
not ( n18553 , n18552 );
not ( n18554 , n18378 );
not ( n18555 , RI15b5ae28_966);
not ( n18556 , n18555 );
and ( n18557 , n18554 , n18556 );
not ( n18558 , RI15b5b1e8_974);
nor ( n18559 , n18387 , n18558 );
nor ( n18560 , n18557 , n18559 );
and ( n18561 , n18317 , RI15b5c0e8_1006);
and ( n18562 , n18312 , RI15b5bd28_998);
nor ( n18563 , n18561 , n18562 );
nand ( n18564 , n18560 , n18563 );
and ( n18565 , n18300 , RI15b5b5a8_982);
not ( n18566 , RI15b5b968_990);
nor ( n18567 , n18306 , n18566 );
nor ( n18568 , n18565 , n18567 );
nand ( n18569 , n18351 , RI15b593e8_910);
nand ( n18570 , n18353 , RI15b59028_902);
nand ( n18571 , n18568 , n18569 , n18570 );
nor ( n18572 , n18564 , n18571 );
nand ( n18573 , n18286 , RI15b5a6a8_950);
nand ( n18574 , n18343 , RI15b5a2e8_942);
not ( n18575 , n18340 );
nand ( n18576 , n18575 , RI15b59f28_934);
and ( n18577 , n18262 , n18289 , n18348 );
nand ( n18578 , n18577 , RI15b5aa68_958);
nand ( n18579 , n18573 , n18574 , n18576 , n18578 );
and ( n18580 , n18360 , RI15b588a8_886);
not ( n18581 , RI15b58c68_894);
nor ( n18582 , n18428 , n18581 );
nor ( n18583 , n18580 , n18582 );
and ( n18584 , n18330 , RI15b597a8_918);
not ( n18585 , RI15b59b68_926);
nor ( n18586 , n18334 , n18585 );
nor ( n18587 , n18584 , n18586 );
nand ( n18588 , n18583 , n18587 );
nor ( n18589 , n18579 , n18588 );
nand ( n18590 , n18572 , n18589 );
not ( n18591 , n18590 );
or ( n18592 , n18446 , RI15b5c4a8_1014);
not ( n18593 , RI15b5c4a8_1014);
or ( n18594 , n18593 , RI15b5c430_1013);
nand ( n18595 , n18592 , n18594 );
not ( n18596 , n18595 );
nand ( n18597 , n18591 , n18596 );
not ( n18598 , n18597 );
nand ( n18599 , n18272 , RI15b5b170_973);
nand ( n18600 , n18277 , RI15b5adb0_965);
nand ( n18601 , n18349 , RI15b59370_909);
and ( n18602 , n18276 , n18328 , n18271 );
nand ( n18603 , n18602 , RI15b58fb0_901);
nand ( n18604 , n18599 , n18600 , n18601 , n18603 );
nand ( n18605 , n18316 , RI15b5c070_1005);
nand ( n18606 , n18312 , RI15b5bcb0_997);
and ( n18607 , n18250 , n18328 , n18292 );
nand ( n18608 , n18607 , RI15b5a270_941);
nand ( n18609 , n18339 , RI15b59eb0_933);
nand ( n18610 , n18605 , n18606 , n18608 , n18609 );
nor ( n18611 , n18604 , n18610 );
nand ( n18612 , n18285 , RI15b5a630_949);
nand ( n18613 , n18358 , RI15b58830_885);
nand ( n18614 , n18362 , RI15b58bf0_893);
nand ( n18615 , n18577 , RI15b5a9f0_957);
nand ( n18616 , n18612 , n18613 , n18614 , n18615 );
nand ( n18617 , n18502 , RI15b5b530_981);
not ( n18618 , n18282 );
and ( n18619 , n18618 , n18328 , n18292 );
nand ( n18620 , n18619 , RI15b59730_917);
not ( n18621 , n18333 );
not ( n18622 , RI15b59af0_925);
not ( n18623 , n18622 );
and ( n18624 , n18621 , n18623 );
not ( n18625 , RI15b5b8f0_989);
nor ( n18626 , n18305 , n18625 );
nor ( n18627 , n18624 , n18626 );
nand ( n18628 , n18617 , n18620 , n18627 );
nor ( n18629 , n18616 , n18628 );
nand ( n18630 , n18611 , n18629 );
not ( n18631 , n18630 );
nand ( n18632 , n18631 , RI15b5c430_1013);
not ( n18633 , n18456 );
not ( n18634 , RI15b5bff8_1004);
not ( n18635 , n18634 );
and ( n18636 , n18633 , n18635 );
not ( n18637 , RI15b5bc38_996);
nor ( n18638 , n18408 , n18637 );
nor ( n18639 , n18636 , n18638 );
not ( n18640 , n18350 );
and ( n18641 , n18640 , RI15b592f8_908);
and ( n18642 , n18353 , RI15b58f38_900);
nor ( n18643 , n18641 , n18642 );
nand ( n18644 , n18639 , n18643 );
nand ( n18645 , n18272 , RI15b5b0f8_972);
nand ( n18646 , n18277 , RI15b5ad38_964);
nand ( n18647 , n18607 , RI15b5a1f8_940);
nand ( n18648 , n18339 , RI15b59e38_932);
nand ( n18649 , n18645 , n18646 , n18647 , n18648 );
nor ( n18650 , n18644 , n18649 );
nand ( n18651 , n18285 , RI15b5a5b8_948);
nand ( n18652 , n18619 , RI15b596b8_916);
nand ( n18653 , n18502 , RI15b5b4b8_980);
nand ( n18654 , n18577 , RI15b5a978_956);
nand ( n18655 , n18651 , n18652 , n18653 , n18654 );
not ( n18656 , n18359 );
nand ( n18657 , n18656 , RI15b587b8_884);
not ( n18658 , n18333 );
and ( n18659 , n18658 , RI15b59a78_924);
not ( n18660 , RI15b5b878_988);
nor ( n18661 , n18305 , n18660 );
nor ( n18662 , n18659 , n18661 );
nand ( n18663 , n18362 , RI15b58b78_892);
nand ( n18664 , n18657 , n18662 , n18663 );
nor ( n18665 , n18655 , n18664 );
nand ( n18666 , n18650 , n18665 );
and ( n18667 , n18666 , RI15b5c3b8_1012);
nand ( n18668 , n18632 , n18667 );
or ( n18669 , n18631 , RI15b5c430_1013);
nand ( n18670 , n18668 , n18669 );
not ( n18671 , n18670 );
or ( n18672 , n18598 , n18671 );
nand ( n18673 , n18590 , n18595 );
nand ( n18674 , n18672 , n18673 );
not ( n18675 , n18674 );
or ( n18676 , n18553 , n18675 );
not ( n18677 , n18544 );
nand ( n18678 , n18677 , n18550 );
nand ( n18679 , n18676 , n18678 );
not ( n18680 , n18679 );
or ( n18681 , n18511 , n18680 );
not ( n18682 , n18509 );
nand ( n18683 , n18682 , n18451 );
nand ( n18684 , n18681 , n18683 );
and ( n18685 , n18231 , n18232 );
not ( n18686 , n18231 );
and ( n18687 , n18686 , RI15b5c610_1017);
nor ( n18688 , n18685 , n18687 );
not ( n18689 , n18688 );
not ( n18690 , n18456 );
not ( n18691 , RI15b5c250_1009);
not ( n18692 , n18691 );
and ( n18693 , n18690 , n18692 );
not ( n18694 , RI15b5be90_1001);
nor ( n18695 , n18408 , n18694 );
nor ( n18696 , n18693 , n18695 );
not ( n18697 , n18387 );
not ( n18698 , RI15b5b350_977);
not ( n18699 , n18698 );
and ( n18700 , n18697 , n18699 );
not ( n18701 , RI15b5af90_969);
nor ( n18702 , n18378 , n18701 );
nor ( n18703 , n18700 , n18702 );
not ( n18704 , n18466 );
not ( n18705 , RI15b5a810_953);
not ( n18706 , n18705 );
and ( n18707 , n18704 , n18706 );
not ( n18708 , RI15b5abd0_961);
nor ( n18709 , n18294 , n18708 );
nor ( n18710 , n18707 , n18709 );
and ( n18711 , n18300 , RI15b5b710_985);
not ( n18712 , RI15b5bad0_993);
nor ( n18713 , n18306 , n18712 );
nor ( n18714 , n18711 , n18713 );
nand ( n18715 , n18696 , n18703 , n18710 , n18714 );
not ( n18716 , n18344 );
not ( n18717 , RI15b5a450_945);
not ( n18718 , n18717 );
and ( n18719 , n18716 , n18718 );
not ( n18720 , RI15b5a090_937);
nor ( n18721 , n18491 , n18720 );
nor ( n18722 , n18719 , n18721 );
not ( n18723 , n18350 );
not ( n18724 , RI15b59550_913);
not ( n18725 , n18724 );
and ( n18726 , n18723 , n18725 );
not ( n18727 , n18602 );
not ( n18728 , RI15b59190_905);
nor ( n18729 , n18727 , n18728 );
nor ( n18730 , n18726 , n18729 );
not ( n18731 , n18359 );
not ( n18732 , RI15b58a10_889);
not ( n18733 , n18732 );
and ( n18734 , n18731 , n18733 );
not ( n18735 , RI15b58dd0_897);
nor ( n18736 , n18428 , n18735 );
nor ( n18737 , n18734 , n18736 );
and ( n18738 , n18329 , RI15b59910_921);
and ( n18739 , n18658 , RI15b59cd0_929);
nor ( n18740 , n18738 , n18739 );
nand ( n18741 , n18722 , n18730 , n18737 , n18740 );
nor ( n18742 , n18715 , n18741 );
buf ( n18743 , n18742 );
buf ( n18744 , n18743 );
nand ( n18745 , n18689 , n18744 );
nand ( n18746 , n18684 , n18745 );
not ( n18747 , n18743 );
nand ( n18748 , n18747 , n18688 );
nand ( n18749 , n18746 , n18748 );
not ( n18750 , n18749 );
or ( n18751 , n18445 , n18750 );
not ( n18752 , n18437 );
nand ( n18753 , n18752 , n18442 );
nand ( n18754 , n18751 , n18753 );
not ( n18755 , n18754 );
or ( n18756 , n18374 , n18755 );
nand ( n18757 , n18366 , n18371 );
nand ( n18758 , n18756 , n18757 );
not ( n18759 , n18758 );
or ( n18760 , n18243 , n18759 );
or ( n18761 , n18758 , n18242 );
nand ( n18762 , n18760 , n18761 );
not ( n18763 , RI15b5d420_1047);
nor ( n18764 , n18763 , RI15b5d3a8_1046);
not ( n18765 , RI15b5d498_1048);
nand ( n18766 , n18764 , n18765 );
not ( n18767 , n18766 );
not ( n18768 , n18264 );
not ( n18769 , n18768 );
not ( n18770 , n18769 );
nand ( n18771 , n18767 , n18770 );
not ( n18772 , n18771 );
not ( n18773 , n18388 );
and ( n18774 , n18772 , n18773 );
nor ( n18775 , RI15b5d2b8_1044 , RI15b5d330_1045);
not ( n18776 , n18775 );
not ( n18777 , n18776 );
nand ( n18778 , n18767 , n18777 );
nor ( n18779 , n18778 , n18397 );
nor ( n18780 , n18774 , n18779 );
not ( n18781 , n18247 );
not ( n18782 , n18781 );
not ( n18783 , n18782 );
nand ( n18784 , n18767 , n18783 );
not ( n18785 , n18784 );
not ( n18786 , n18400 );
and ( n18787 , n18785 , n18786 );
not ( n18788 , n18766 );
not ( n18789 , n18245 );
nand ( n18790 , n18788 , n18789 );
nor ( n18791 , n18790 , n18380 );
nor ( n18792 , n18787 , n18791 );
not ( n18793 , n18258 );
nand ( n18794 , n18781 , n18793 );
nor ( n18795 , n18794 , RI15b5d498_1048);
buf ( n18796 , n18795 );
and ( n18797 , n18796 , RI15b59d48_930);
nand ( n18798 , RI15b5d3a8_1046 , RI15b5d420_1047);
nor ( n18799 , n18798 , n18245 );
not ( n18800 , RI15b5d498_1048);
and ( n18801 , n18799 , n18800 );
not ( n18802 , n18801 );
not ( n18803 , n18802 );
and ( n18804 , n18803 , RI15b5bf08_1002);
nor ( n18805 , n18797 , n18804 );
not ( n18806 , n18798 );
nand ( n18807 , n18781 , n18806 );
or ( n18808 , n18807 , RI15b5d498_1048);
not ( n18809 , n18808 );
nand ( n18810 , n18809 , RI15b5bb48_994);
nand ( n18811 , n18780 , n18792 , n18805 , n18810 );
nor ( n18812 , RI15b5d3a8_1046 , RI15b5d420_1047);
not ( n18813 , RI15b5d498_1048);
nand ( n18814 , n18812 , n18813 );
not ( n18815 , n18814 );
nand ( n18816 , n18815 , n18768 );
not ( n18817 , n18816 );
not ( n18818 , n18417 );
and ( n18819 , n18817 , n18818 );
not ( n18820 , n18814 );
nand ( n18821 , n18820 , n18775 );
nor ( n18822 , n18821 , n18425 );
nor ( n18823 , n18819 , n18822 );
buf ( n18824 , n18814 );
not ( n18825 , n18824 );
not ( n18826 , n18782 );
nand ( n18827 , n18825 , n18826 );
not ( n18828 , n18827 );
not ( n18829 , n18429 );
and ( n18830 , n18828 , n18829 );
not ( n18831 , n18824 );
nand ( n18832 , n18831 , n18789 );
nor ( n18833 , n18832 , n18420 );
nor ( n18834 , n18830 , n18833 );
not ( n18835 , n18260 );
not ( n18836 , RI15b5d498_1048);
nand ( n18837 , n18835 , n18836 );
not ( n18838 , n18837 );
nand ( n18839 , n18838 , RI15b5a4c8_946);
nand ( n18840 , n18823 , n18834 , n18839 );
nor ( n18841 , n18811 , n18840 );
not ( n18842 , RI15b5a108_938);
nand ( n18843 , n18789 , n18793 );
nor ( n18844 , n18843 , RI15b5d498_1048);
buf ( n18845 , n18844 );
not ( n18846 , n18845 );
or ( n18847 , n18842 , n18846 );
nor ( n18848 , RI15b5d2b8_1044 , RI15b5d330_1045);
nand ( n18849 , n18848 , n18793 );
not ( n18850 , n18849 );
not ( n18851 , RI15b5d498_1048);
nand ( n18852 , n18850 , n18851 );
not ( n18853 , n18852 );
nand ( n18854 , n18853 , RI15b59988_922);
nand ( n18855 , n18847 , n18854 );
not ( n18856 , RI15b5c2c8_1010);
nand ( n18857 , RI15b5d3a8_1046 , RI15b5d420_1047);
not ( n18858 , n18857 );
nand ( n18859 , n18768 , n18858 );
or ( n18860 , n18859 , RI15b5d498_1048);
not ( n18861 , n18860 );
not ( n18862 , n18861 );
or ( n18863 , n18856 , n18862 );
nand ( n18864 , n18848 , n18858 );
not ( n18865 , n18864 );
not ( n18866 , RI15b5d498_1048);
nand ( n18867 , n18865 , n18866 );
not ( n18868 , n18867 );
nand ( n18869 , n18868 , RI15b5b788_986);
nand ( n18870 , n18863 , n18869 );
nor ( n18871 , n18855 , n18870 );
nand ( n18872 , n18841 , n18871 );
buf ( n18873 , n18872 );
not ( n18874 , n18771 );
not ( n18875 , n18480 );
and ( n18876 , n18874 , n18875 );
nor ( n18877 , n18778 , n18468 );
nor ( n18878 , n18876 , n18877 );
not ( n18879 , n18784 );
not ( n18880 , n18471 );
and ( n18881 , n18879 , n18880 );
nand ( n18882 , n18788 , n18789 );
nor ( n18883 , n18882 , n18483 );
nor ( n18884 , n18881 , n18883 );
buf ( n18885 , n18795 );
and ( n18886 , n18885 , RI15b59c58_928);
buf ( n18887 , n18801 );
and ( n18888 , n18887 , RI15b5be18_1000);
nor ( n18889 , n18886 , n18888 );
nand ( n18890 , n18809 , RI15b5ba58_992);
nand ( n18891 , n18878 , n18884 , n18889 , n18890 );
not ( n18892 , n18891 );
not ( n18893 , n18821 );
and ( n18894 , n18893 , RI15b58998_888);
not ( n18895 , n18816 );
and ( n18896 , n18895 , RI15b594d8_912);
nor ( n18897 , n18894 , n18896 );
not ( n18898 , n18827 );
and ( n18899 , n18898 , RI15b58d58_896);
not ( n18900 , n18832 );
and ( n18901 , n18900 , RI15b59118_904);
nor ( n18902 , n18899 , n18901 );
nand ( n18903 , n18838 , RI15b5a3d8_944);
and ( n18904 , n18897 , n18902 , n18903 );
not ( n18905 , RI15b5a018_936);
not ( n18906 , n18844 );
or ( n18907 , n18905 , n18906 );
nand ( n18908 , n18853 , RI15b59898_920);
nand ( n18909 , n18907 , n18908 );
not ( n18910 , RI15b5b698_984);
not ( n18911 , n18867 );
not ( n18912 , n18911 );
or ( n18913 , n18910 , n18912 );
not ( n18914 , n18860 );
nand ( n18915 , n18914 , RI15b5c1d8_1008);
nand ( n18916 , n18913 , n18915 );
nor ( n18917 , n18909 , n18916 );
nand ( n18918 , n18892 , n18904 , n18917 );
not ( n18919 , n18918 );
nand ( n18920 , n18873 , n18919 );
not ( n18921 , n18769 );
nand ( n18922 , n18788 , n18921 );
not ( n18923 , n18922 );
not ( n18924 , RI15b5b0f8_972);
not ( n18925 , n18924 );
and ( n18926 , n18923 , n18925 );
not ( n18927 , n18776 );
nand ( n18928 , n18767 , n18927 );
not ( n18929 , RI15b5a5b8_948);
nor ( n18930 , n18928 , n18929 );
nor ( n18931 , n18926 , n18930 );
nand ( n18932 , n18788 , n18826 );
not ( n18933 , n18932 );
not ( n18934 , RI15b5a978_956);
not ( n18935 , n18934 );
and ( n18936 , n18933 , n18935 );
not ( n18937 , RI15b5ad38_964);
nor ( n18938 , n18790 , n18937 );
nor ( n18939 , n18936 , n18938 );
not ( n18940 , RI15b59a78_924);
not ( n18941 , n18795 );
or ( n18942 , n18940 , n18941 );
nand ( n18943 , n18801 , RI15b5bc38_996);
nand ( n18944 , n18942 , n18943 );
not ( n18945 , n18944 );
nand ( n18946 , n18809 , RI15b5b878_988);
nand ( n18947 , n18931 , n18939 , n18945 , n18946 );
nand ( n18948 , n18844 , RI15b59e38_932);
nand ( n18949 , n18868 , RI15b5b4b8_980);
nand ( n18950 , n18861 , RI15b5bff8_1004);
not ( n18951 , n18852 );
nand ( n18952 , n18951 , RI15b596b8_916);
nand ( n18953 , n18948 , n18949 , n18950 , n18952 );
not ( n18954 , n18821 );
not ( n18955 , RI15b587b8_884);
not ( n18956 , n18955 );
and ( n18957 , n18954 , n18956 );
not ( n18958 , RI15b592f8_908);
nor ( n18959 , n18816 , n18958 );
nor ( n18960 , n18957 , n18959 );
not ( n18961 , n18827 );
not ( n18962 , RI15b58b78_892);
not ( n18963 , n18962 );
and ( n18964 , n18961 , n18963 );
not ( n18965 , RI15b58f38_900);
nor ( n18966 , n18832 , n18965 );
nor ( n18967 , n18964 , n18966 );
nand ( n18968 , n18838 , RI15b5a1f8_940);
nand ( n18969 , n18960 , n18967 , n18968 );
nor ( n18970 , n18947 , n18953 , n18969 );
not ( n18971 , n18970 );
not ( n18972 , n18971 );
nor ( n18973 , n18920 , n18972 );
nor ( n18974 , n18922 , n18558 );
not ( n18975 , RI15b5aa68_958);
nor ( n18976 , n18932 , n18975 );
nor ( n18977 , n18974 , n18976 );
nor ( n18978 , n18790 , n18555 );
not ( n18979 , RI15b5a6a8_950);
nor ( n18980 , n18928 , n18979 );
nor ( n18981 , n18978 , n18980 );
nand ( n18982 , n18911 , RI15b5b5a8_982);
nand ( n18983 , n18977 , n18981 , n18982 );
not ( n18984 , RI15b59b68_926);
not ( n18985 , n18795 );
or ( n18986 , n18984 , n18985 );
nand ( n18987 , n18801 , RI15b5bd28_998);
nand ( n18988 , n18986 , n18987 );
not ( n18989 , n18988 );
not ( n18990 , RI15b593e8_910);
nor ( n18991 , n18816 , n18990 );
not ( n18992 , RI15b588a8_886);
nor ( n18993 , n18821 , n18992 );
nor ( n18994 , n18991 , n18993 );
not ( n18995 , n18814 );
nand ( n18996 , n18995 , n18789 );
not ( n18997 , RI15b59028_902);
nor ( n18998 , n18996 , n18997 );
not ( n18999 , n18814 );
nand ( n19000 , n18999 , n18783 );
nor ( n19001 , n19000 , n18581 );
nor ( n19002 , n18998 , n19001 );
nand ( n19003 , n18809 , RI15b5b968_990);
nand ( n19004 , n18989 , n18994 , n19002 , n19003 );
nand ( n19005 , n18844 , RI15b59f28_934);
not ( n19006 , n18860 );
nand ( n19007 , n19006 , RI15b5c0e8_1006);
not ( n19008 , n18852 );
nand ( n19009 , n19008 , RI15b597a8_918);
nand ( n19010 , n18838 , RI15b5a2e8_942);
nand ( n19011 , n19005 , n19007 , n19009 , n19010 );
nor ( n19012 , n18983 , n19004 , n19011 );
not ( n19013 , n18882 );
not ( n19014 , RI15b5b080_971);
not ( n19015 , n19014 );
and ( n19016 , n19013 , n19015 );
not ( n19017 , RI15b5a900_955);
nor ( n19018 , n18928 , n19017 );
nor ( n19019 , n19016 , n19018 );
not ( n19020 , n18922 );
not ( n19021 , RI15b5b440_979);
not ( n19022 , n19021 );
and ( n19023 , n19020 , n19022 );
nor ( n19024 , n18932 , n18295 );
nor ( n19025 , n19023 , n19024 );
nand ( n19026 , n18911 , RI15b5b800_987);
nand ( n19027 , n19019 , n19025 , n19026 );
not ( n19028 , n19027 );
not ( n19029 , RI15b59640_915);
nor ( n19030 , n18816 , n19029 );
not ( n19031 , RI15b58b00_891);
nor ( n19032 , n18821 , n19031 );
nor ( n19033 , n19030 , n19032 );
not ( n19034 , RI15b59280_907);
nor ( n19035 , n18996 , n19034 );
not ( n19036 , RI15b58ec0_899);
nor ( n19037 , n19000 , n19036 );
nor ( n19038 , n19035 , n19037 );
nand ( n19039 , n18809 , RI15b5bbc0_995);
nand ( n19040 , n19033 , n19038 , n19039 );
not ( n19041 , RI15b59dc0_931);
buf ( n19042 , n18795 );
not ( n19043 , n19042 );
or ( n19044 , n19041 , n19043 );
not ( n19045 , n18802 );
nand ( n19046 , n19045 , RI15b5bf80_1003);
nand ( n19047 , n19044 , n19046 );
nor ( n19048 , n19040 , n19047 );
not ( n19049 , RI15b5a180_939);
not ( n19050 , n18844 );
or ( n19051 , n19049 , n19050 );
nand ( n19052 , n18951 , RI15b59a00_923);
nand ( n19053 , n19051 , n19052 );
not ( n19054 , RI15b5c340_1011);
not ( n19055 , n18914 );
or ( n19056 , n19054 , n19055 );
nand ( n19057 , n18838 , RI15b5a540_947);
nand ( n19058 , n19056 , n19057 );
nor ( n19059 , n19053 , n19058 );
nand ( n19060 , n19028 , n19048 , n19059 );
nand ( n19061 , n19012 , n19060 );
not ( n19062 , n18771 );
not ( n19063 , RI15b5b260_975);
not ( n19064 , n19063 );
and ( n19065 , n19062 , n19064 );
not ( n19066 , RI15b5a720_951);
nor ( n19067 , n18778 , n19066 );
nor ( n19068 , n19065 , n19067 );
not ( n19069 , n18784 );
not ( n19070 , n18523 );
and ( n19071 , n19069 , n19070 );
not ( n19072 , RI15b5aea0_967);
nor ( n19073 , n18882 , n19072 );
nor ( n19074 , n19071 , n19073 );
and ( n19075 , n18796 , RI15b59be0_927);
and ( n19076 , n18803 , RI15b5bda0_999);
nor ( n19077 , n19075 , n19076 );
nand ( n19078 , n18809 , RI15b5b9e0_991);
nand ( n19079 , n19068 , n19074 , n19077 , n19078 );
not ( n19080 , n18816 );
not ( n19081 , RI15b59460_911);
not ( n19082 , n19081 );
and ( n19083 , n19080 , n19082 );
not ( n19084 , RI15b58920_887);
nor ( n19085 , n18821 , n19084 );
nor ( n19086 , n19083 , n19085 );
not ( n19087 , n18827 );
not ( n19088 , n18529 );
and ( n19089 , n19087 , n19088 );
not ( n19090 , RI15b590a0_903);
nor ( n19091 , n18832 , n19090 );
nor ( n19092 , n19089 , n19091 );
nand ( n19093 , n18838 , RI15b5a360_943);
nand ( n19094 , n19086 , n19092 , n19093 );
nor ( n19095 , n19079 , n19094 );
not ( n19096 , RI15b59fa0_935);
not ( n19097 , n18845 );
or ( n19098 , n19096 , n19097 );
nand ( n19099 , n18853 , RI15b59820_919);
nand ( n19100 , n19098 , n19099 );
not ( n19101 , RI15b5b620_983);
not ( n19102 , n18911 );
or ( n19103 , n19101 , n19102 );
nand ( n19104 , n18861 , RI15b5c160_1007);
nand ( n19105 , n19103 , n19104 );
nor ( n19106 , n19100 , n19105 );
nand ( n19107 , n19095 , n19106 );
nor ( n19108 , n18771 , n18698 );
nor ( n19109 , n18932 , n18708 );
nor ( n19110 , n19108 , n19109 );
nor ( n19111 , n18790 , n18701 );
nor ( n19112 , n18928 , n18705 );
nor ( n19113 , n19111 , n19112 );
nand ( n19114 , n18911 , RI15b5b710_985);
nand ( n19115 , n19110 , n19113 , n19114 );
not ( n19116 , n18802 );
not ( n19117 , n18694 );
and ( n19118 , n19116 , n19117 );
and ( n19119 , n19042 , RI15b59cd0_929);
nor ( n19120 , n19118 , n19119 );
not ( n19121 , n18816 );
not ( n19122 , n18724 );
and ( n19123 , n19121 , n19122 );
nor ( n19124 , n18821 , n18732 );
nor ( n19125 , n19123 , n19124 );
not ( n19126 , n18827 );
not ( n19127 , n18735 );
and ( n19128 , n19126 , n19127 );
nor ( n19129 , n18996 , n18728 );
nor ( n19130 , n19128 , n19129 );
nand ( n19131 , n18809 , RI15b5bad0_993);
nand ( n19132 , n19120 , n19125 , n19130 , n19131 );
nor ( n19133 , n19115 , n19132 );
not ( n19134 , RI15b5a090_937);
not ( n19135 , n18844 );
or ( n19136 , n19134 , n19135 );
nand ( n19137 , n18853 , RI15b59910_921);
nand ( n19138 , n19136 , n19137 );
not ( n19139 , RI15b5c250_1009);
not ( n19140 , n18914 );
or ( n19141 , n19139 , n19140 );
nand ( n19142 , n18838 , RI15b5a450_945);
nand ( n19143 , n19141 , n19142 );
nor ( n19144 , n19138 , n19143 );
nand ( n19145 , n19133 , n19144 );
nand ( n19146 , n19107 , n19145 );
nor ( n19147 , n19061 , n19146 );
nand ( n19148 , n18973 , n19147 );
not ( n19149 , n18816 );
not ( n19150 , RI15b59370_909);
not ( n19151 , n19150 );
and ( n19152 , n19149 , n19151 );
not ( n19153 , RI15b58830_885);
nor ( n19154 , n18821 , n19153 );
nor ( n19155 , n19152 , n19154 );
not ( n19156 , n18778 );
nand ( n19157 , n19156 , RI15b5a630_949);
not ( n19158 , n18882 );
nand ( n19159 , n19158 , RI15b5adb0_965);
and ( n19160 , n19155 , n19157 , n19159 );
not ( n19161 , n19000 );
not ( n19162 , RI15b58bf0_893);
not ( n19163 , n19162 );
and ( n19164 , n19161 , n19163 );
not ( n19165 , RI15b58fb0_901);
nor ( n19166 , n18996 , n19165 );
nor ( n19167 , n19164 , n19166 );
not ( n19168 , n18784 );
nand ( n19169 , n19168 , RI15b5a9f0_957);
not ( n19170 , n18922 );
nand ( n19171 , n19170 , RI15b5b170_973);
and ( n19172 , n19167 , n19169 , n19171 );
not ( n19173 , n18837 );
not ( n19174 , RI15b5a270_941);
not ( n19175 , n19174 );
and ( n19176 , n19173 , n19175 );
and ( n19177 , n18861 , RI15b5c070_1005);
nor ( n19178 , n19176 , n19177 );
and ( n19179 , n18885 , RI15b59af0_925);
and ( n19180 , n18887 , RI15b5bcb0_997);
nor ( n19181 , n19179 , n19180 );
nand ( n19182 , n19160 , n19172 , n19178 , n19181 );
and ( n19183 , n18845 , RI15b59eb0_933);
and ( n19184 , n18809 , RI15b5b8f0_989);
nor ( n19185 , n19183 , n19184 );
and ( n19186 , n18853 , RI15b59730_917);
and ( n19187 , n18868 , RI15b5b530_981);
nor ( n19188 , n19186 , n19187 );
nand ( n19189 , n19185 , n19188 );
nor ( n19190 , n19182 , n19189 );
not ( n19191 , n19190 );
not ( n19192 , n19191 );
buf ( n19193 , n19192 );
nor ( n19194 , n19148 , n19193 );
not ( n19195 , RI15b5d588_1050);
nor ( n19196 , n19195 , RI15b5d6f0_1053);
not ( n19197 , n19196 );
not ( n19198 , RI15b5d600_1051);
nand ( n19199 , n19198 , RI15b5d678_1052);
or ( n19200 , n19197 , n19199 );
not ( n19201 , n19200 );
nand ( n19202 , n19194 , n19201 );
not ( n19203 , RI15b58740_883);
nand ( n19204 , n19203 , RI15b5d498_1048);
not ( n19205 , n19204 );
not ( n19206 , RI15b586c8_882);
nand ( n19207 , n19206 , RI15b5d420_1047);
not ( n19208 , n19207 );
not ( n19209 , RI15b58650_881);
nand ( n19210 , n19209 , RI15b5d3a8_1046);
not ( n19211 , n19210 );
nor ( n19212 , RI15b58560_879 , RI15b585d8_880);
or ( n19213 , n19212 , RI15b5d330_1045);
not ( n19214 , RI15b5d2b8_1044);
nand ( n19215 , n19214 , RI15b585d8_880);
nand ( n19216 , RI15b58560_879 , RI15b585d8_880);
buf ( n19217 , n19216 );
nand ( n19218 , n18776 , n19213 , n19215 , n19217 );
not ( n19219 , n19218 );
or ( n19220 , n19211 , n19219 );
nand ( n19221 , n18268 , RI15b58650_881);
nand ( n19222 , n19220 , n19221 );
not ( n19223 , n19222 );
or ( n19224 , n19208 , n19223 );
not ( n19225 , RI15b5d420_1047);
nand ( n19226 , n19225 , RI15b586c8_882);
nand ( n19227 , n19224 , n19226 );
not ( n19228 , n19227 );
or ( n19229 , n19205 , n19228 );
not ( n19230 , RI15b5d498_1048);
nand ( n19231 , n19230 , RI15b58740_883);
nand ( n19232 , n19229 , n19231 );
and ( n19233 , n19218 , RI15b5d3a8_1046);
not ( n19234 , n19218 );
and ( n19235 , n19234 , n18268 );
nor ( n19236 , n19233 , n19235 );
and ( n19237 , n19236 , n19209 );
not ( n19238 , n19236 );
and ( n19239 , n19238 , RI15b58650_881);
nor ( n19240 , n19237 , n19239 );
nand ( n19241 , n19232 , n19240 );
nand ( n19242 , n19226 , n19207 , n19231 );
not ( n19243 , n19242 );
not ( n19244 , n19222 );
or ( n19245 , n19243 , n19244 );
not ( n19246 , RI15b5d420_1047);
or ( n19247 , n19246 , RI15b5d498_1048);
nand ( n19248 , n19247 , n19206 );
nor ( n19249 , n19222 , n19248 );
or ( n19250 , n19231 , n19206 );
nand ( n19251 , n19250 , n19204 );
nor ( n19252 , n19249 , n19251 );
nand ( n19253 , n19245 , n19252 );
nand ( n19254 , n19232 , n19253 );
buf ( n19255 , n19254 );
buf ( n19256 , n18777 );
not ( n19257 , n19256 );
buf ( n19258 , n19257 );
not ( n19259 , n19258 );
and ( n19260 , n19259 , RI15b585d8_880);
not ( n19261 , RI15b585d8_880);
and ( n19262 , n18789 , n19261 );
nor ( n19263 , n19260 , n19262 );
not ( n19264 , RI15b58560_879);
or ( n19265 , n19263 , n19264 );
buf ( n19266 , n18783 );
buf ( n19267 , n19266 );
buf ( n19268 , n19212 );
and ( n19269 , n19267 , n19268 );
and ( n19270 , n19264 , RI15b585d8_880);
not ( n19271 , n19270 );
not ( n19272 , n19271 );
buf ( n19273 , n19272 );
buf ( n19274 , n18770 );
buf ( n19275 , n19274 );
and ( n19276 , n19273 , n19275 );
nor ( n19277 , n19269 , n19276 );
nand ( n19278 , n19265 , n19277 );
nand ( n19279 , n19232 , n19278 );
and ( n19280 , n19241 , n19255 , n19279 );
nor ( n19281 , n19202 , n19280 );
nand ( n19282 , n19281 , n18367 );
buf ( n19283 , n19282 );
buf ( n19284 , n19283 );
buf ( n19285 , n19284 );
not ( n19286 , n19285 );
buf ( n19287 , n19286 );
and ( n19288 , n18762 , n19287 );
not ( n19289 , RI15b5c688_1018);
buf ( n19290 , n18230 );
nand ( n19291 , RI15b5c3b8_1012 , RI15b5c430_1013);
buf ( n19292 , n19291 );
not ( n19293 , n19292 );
nand ( n19294 , n19290 , n19293 );
or ( n19295 , n19294 , n18232 );
not ( n19296 , n19295 );
or ( n19297 , n19289 , n19296 );
or ( n19298 , n19295 , RI15b5c688_1018);
nand ( n19299 , n19297 , n19298 );
not ( n19300 , n19299 );
nand ( n19301 , n18437 , n19300 );
not ( n19302 , n19301 );
buf ( n19303 , n19292 );
nor ( n19304 , n19303 , n18228 );
and ( n19305 , n19304 , n18229 );
not ( n19306 , n19304 );
and ( n19307 , n19306 , RI15b5c598_1016);
nor ( n19308 , n19305 , n19307 );
nand ( n19309 , n18508 , n19308 );
and ( n19310 , n19294 , RI15b5c610_1017);
not ( n19311 , n19294 );
and ( n19312 , n19311 , n18232 );
nor ( n19313 , n19310 , n19312 );
nand ( n19314 , n18742 , n19313 );
nand ( n19315 , n19309 , n19314 );
not ( n19316 , n18543 );
nand ( n19317 , n19293 , RI15b5c4a8_1014);
and ( n19318 , n19317 , RI15b5c520_1015);
not ( n19319 , n19317 );
and ( n19320 , n19319 , n18546 );
nor ( n19321 , n19318 , n19320 );
and ( n19322 , n19316 , n19321 );
nor ( n19323 , n19315 , n19322 );
not ( n19324 , n19323 );
and ( n19325 , n19303 , RI15b5c4a8_1014);
not ( n19326 , n19303 );
and ( n19327 , n19326 , n18593 );
nor ( n19328 , n19325 , n19327 );
nand ( n19329 , n18591 , n19328 );
not ( n19330 , n19329 );
nand ( n19331 , n18446 , RI15b5c3b8_1012);
not ( n19332 , n19331 );
not ( n19333 , n18631 );
or ( n19334 , n19332 , n19333 );
nand ( n19335 , n19334 , n18666 );
not ( n19336 , RI15b5c3b8_1012);
nand ( n19337 , n19336 , RI15b5c430_1013);
nand ( n19338 , n19335 , n18669 , n19337 );
not ( n19339 , n19338 );
or ( n19340 , n19330 , n19339 );
not ( n19341 , n19328 );
nand ( n19342 , n18590 , n19341 );
nand ( n19343 , n19340 , n19342 );
not ( n19344 , n19343 );
or ( n19345 , n19324 , n19344 );
not ( n19346 , n19315 );
or ( n19347 , n18544 , n19321 );
not ( n19348 , n19347 );
and ( n19349 , n19346 , n19348 );
not ( n19350 , n18508 );
not ( n19351 , n19308 );
nand ( n19352 , n19350 , n19351 );
not ( n19353 , n19314 );
or ( n19354 , n19352 , n19353 );
not ( n19355 , n18742 );
not ( n19356 , n19313 );
nand ( n19357 , n19355 , n19356 );
nand ( n19358 , n19354 , n19357 );
nor ( n19359 , n19349 , n19358 );
nand ( n19360 , n19345 , n19359 );
not ( n19361 , n19360 );
or ( n19362 , n19302 , n19361 );
nand ( n19363 , n18752 , n19299 );
nand ( n19364 , n19362 , n19363 );
not ( n19365 , n19295 );
nand ( n19366 , n19365 , RI15b5c688_1018);
and ( n19367 , n19366 , n18235 );
not ( n19368 , n19366 );
and ( n19369 , n19368 , RI15b5c700_1019);
nor ( n19370 , n19367 , n19369 );
nor ( n19371 , n19364 , n19370 );
not ( n19372 , n19371 );
nand ( n19373 , n18236 , RI15b5c3b8_1012);
and ( n19374 , n19373 , n18238 );
not ( n19375 , n19373 );
and ( n19376 , n19375 , RI15b5c778_1020);
nor ( n19377 , n19374 , n19376 );
and ( n19378 , n19372 , n19377 );
not ( n19379 , n19370 );
nand ( n19380 , n19379 , n18367 );
nand ( n19381 , n19364 , n19380 );
and ( n19382 , n18366 , n19370 );
nor ( n19383 , n19382 , n19377 );
nand ( n19384 , n19381 , n19383 );
not ( n19385 , n19384 );
nor ( n19386 , n19378 , n19385 );
and ( n19387 , n19281 , n18366 );
not ( n19388 , n19387 );
buf ( n19389 , n19388 );
not ( n19390 , n19389 );
buf ( n19391 , n19390 );
not ( n19392 , n19391 );
or ( n19393 , n19386 , n19392 );
nand ( n19394 , n19291 , n18593 );
nand ( n19395 , n19394 , RI15b5c520_1015);
nor ( n19396 , n19395 , n18229 );
nand ( n19397 , n19396 , RI15b5c610_1017);
nor ( n19398 , n19397 , n18440 );
nand ( n19399 , n19398 , RI15b5c700_1019);
and ( n19400 , n19399 , n18238 );
not ( n19401 , n19399 );
and ( n19402 , n19401 , RI15b5c778_1020);
nor ( n19403 , n19400 , n19402 );
not ( n19404 , n19403 );
not ( n19405 , n19398 );
and ( n19406 , n19405 , n18235 );
not ( n19407 , n19405 );
and ( n19408 , n19407 , RI15b5c700_1019);
nor ( n19409 , n19406 , n19408 );
and ( n19410 , n18366 , n19409 );
not ( n19411 , n19410 );
nor ( n19412 , n18366 , n19409 );
not ( n19413 , n19412 );
not ( n19414 , n18437 );
and ( n19415 , n19397 , RI15b5c688_1018);
not ( n19416 , n19397 );
and ( n19417 , n19416 , n18440 );
nor ( n19418 , n19415 , n19417 );
not ( n19419 , n19418 );
and ( n19420 , n19414 , n19419 );
nand ( n19421 , n18591 , n19341 );
not ( n19422 , n19421 );
nand ( n19423 , n19337 , n19331 );
nand ( n19424 , n18630 , n19423 );
not ( n19425 , n18446 );
not ( n19426 , n18631 );
or ( n19427 , n19425 , n19426 );
not ( n19428 , n18666 );
nor ( n19429 , n19428 , RI15b5c3b8_1012);
nand ( n19430 , n19427 , n19429 );
nand ( n19431 , n19424 , n19430 );
not ( n19432 , n19431 );
or ( n19433 , n19422 , n19432 );
nand ( n19434 , n18590 , n19328 );
nand ( n19435 , n19433 , n19434 );
nand ( n19436 , n18436 , n19418 );
nor ( n19437 , n19292 , n18546 );
not ( n19438 , n19437 );
nand ( n19439 , n19438 , n18228 );
and ( n19440 , n19439 , n18229 );
and ( n19441 , n19395 , RI15b5c598_1016);
nor ( n19442 , n19440 , n19441 );
and ( n19443 , n18508 , n19442 );
not ( n19444 , n19443 );
and ( n19445 , RI15b5c610_1017 , n19396 );
not ( n19446 , RI15b5c610_1017);
and ( n19447 , n19437 , RI15b5c598_1016);
nor ( n19448 , n19447 , n19290 );
and ( n19449 , n19446 , n19448 );
nor ( n19450 , n19445 , n19449 );
not ( n19451 , n19450 );
nand ( n19452 , n19451 , n18742 );
and ( n19453 , n19394 , RI15b5c520_1015);
not ( n19454 , n19394 );
and ( n19455 , n19454 , n18546 );
nor ( n19456 , n19453 , n19455 );
not ( n19457 , n19456 );
nand ( n19458 , n19316 , n19457 );
and ( n19459 , n19436 , n19444 , n19452 , n19458 );
and ( n19460 , n19435 , n19459 );
nor ( n19461 , n19420 , n19460 );
not ( n19462 , n19450 );
nor ( n19463 , n18742 , n19462 );
not ( n19464 , n19463 );
nand ( n19465 , n18543 , n19456 );
nor ( n19466 , n19443 , n19465 );
not ( n19467 , n19395 );
or ( n19468 , n19467 , RI15b5c598_1016);
nand ( n19469 , n19468 , n19448 );
nor ( n19470 , n18508 , n19469 );
or ( n19471 , n19466 , n19470 );
nand ( n19472 , n19471 , n19452 );
nand ( n19473 , n19464 , n19472 );
nand ( n19474 , n19473 , n19436 );
nand ( n19475 , n19461 , n19474 );
nand ( n19476 , n19413 , n19475 );
nand ( n19477 , n19411 , n19476 );
not ( n19478 , n19477 );
not ( n19479 , n19478 );
or ( n19480 , n19404 , n19479 );
or ( n19481 , n19478 , n19403 );
nand ( n19482 , n19480 , n19481 );
nand ( n19483 , n19192 , n19201 );
nor ( n19484 , n19148 , n19483 );
and ( n19485 , n18249 , RI15b58560_879);
and ( n19486 , n19264 , RI15b5d2b8_1044);
and ( n19487 , n18302 , RI15b585d8_880);
and ( n19488 , n19261 , RI15b5d330_1045);
nor ( n19489 , n19487 , n19488 );
not ( n19490 , n19489 );
nor ( n19491 , n19485 , n19486 , n19490 );
nor ( n19492 , n19241 , n19491 );
not ( n19493 , n19492 );
nand ( n19494 , n19493 , n19255 );
buf ( n19495 , n19494 );
not ( n19496 , n19495 );
not ( n19497 , n19496 );
and ( n19498 , n19484 , n19497 );
not ( n19499 , n19498 );
not ( n19500 , n19499 );
not ( n19501 , n19500 );
not ( n19502 , n19501 );
and ( n19503 , n19482 , n19502 );
nor ( n19504 , RI15b5d600_1051 , RI15b5d678_1052);
not ( n19505 , RI15b5d6f0_1053);
nand ( n19506 , n19195 , n19505 );
and ( n19507 , n19504 , n19506 );
not ( n19508 , n19504 );
not ( n19509 , RI15b5d588_1050);
nand ( n19510 , n19509 , RI15b5d6f0_1053);
and ( n19511 , n19508 , n19510 );
or ( n19512 , n19507 , n19511 );
not ( n19513 , n19512 );
and ( n19514 , n19513 , RI15b63e10_1273);
nor ( n19515 , n19503 , n19514 );
nand ( n19516 , n19393 , n19515 );
nor ( n19517 , n19288 , n19516 );
nor ( n19518 , n18920 , n19107 );
not ( n19519 , n19012 );
buf ( n19520 , n19060 );
nor ( n19521 , n19145 , n19519 , n19520 );
nand ( n19522 , n19518 , n19521 );
not ( n19523 , n19522 );
and ( n19524 , n19190 , n18970 );
and ( n19525 , n19523 , n19524 );
nor ( n19526 , n18919 , n18873 );
nand ( n19527 , n19147 , n19526 );
not ( n19528 , n19527 );
not ( n19529 , n19524 );
nand ( n19530 , n19191 , n18971 );
nand ( n19531 , n19529 , n19530 );
nand ( n19532 , n19528 , n19531 );
not ( n19533 , n19532 );
nor ( n19534 , n19525 , n19533 , n19200 );
not ( n19535 , n19534 );
not ( n19536 , n18971 );
and ( n19537 , n19191 , n19536 );
and ( n19538 , n19520 , n19519 , n19145 );
nand ( n19539 , n19518 , n19537 , n19538 );
nor ( n19540 , n19061 , n19145 );
nor ( n19541 , n18918 , n18872 );
nand ( n19542 , n19540 , n19541 , n19107 , n18971 );
not ( n19543 , n19542 );
nand ( n19544 , n19543 , n19192 );
nand ( n19545 , n19539 , n19544 );
not ( n19546 , n18920 );
not ( n19547 , n19107 );
nand ( n19548 , n19546 , n19538 , n19524 , n19547 );
not ( n19549 , n19542 );
not ( n19550 , n19192 );
nand ( n19551 , n19549 , n19550 );
nand ( n19552 , n19548 , n19551 );
or ( n19553 , n19545 , n19552 );
not ( n19554 , n19553 );
and ( n19555 , n18873 , n19547 );
nand ( n19556 , n19540 , n19555 , n19524 );
and ( n19557 , n19556 , n19148 );
nand ( n19558 , n19554 , n19557 );
not ( n19559 , n19558 );
not ( n19560 , n19559 );
or ( n19561 , n19535 , n19560 );
nand ( n19562 , n19524 , n19201 );
not ( n19563 , n19562 );
nand ( n19564 , n19523 , n19563 );
buf ( n19565 , n19564 );
nand ( n19566 , n19561 , n19565 );
not ( n19567 , n19495 );
not ( n19568 , n19567 );
not ( n19569 , n19484 );
or ( n19570 , n19568 , n19569 );
not ( n19571 , n19202 );
nand ( n19572 , n19571 , n19280 );
nand ( n19573 , n19570 , n19572 );
not ( n19574 , RI15b5d678_1052);
nand ( n19575 , n19574 , RI15b5d600_1051);
not ( n19576 , n19575 );
nand ( n19577 , n19576 , n19196 );
nand ( n19578 , RI15b5d600_1051 , RI15b5d678_1052);
or ( n19579 , n19506 , n19578 );
nand ( n19580 , n19577 , n19579 );
not ( n19581 , n19580 );
nor ( n19582 , RI15b5d600_1051 , RI15b5d678_1052);
not ( n19583 , n19582 );
not ( n19584 , n19583 );
and ( n19585 , n19584 , n19196 );
not ( n19586 , n19584 );
nand ( n19587 , RI15b5d588_1050 , RI15b5d6f0_1053);
not ( n19588 , n19587 );
and ( n19589 , n19586 , n19588 );
nor ( n19590 , n19585 , n19589 );
nand ( n19591 , n19581 , n19590 );
not ( n19592 , n19591 );
not ( n19593 , n19578 );
nand ( n19594 , n19196 , n19593 );
or ( n19595 , n19583 , n19510 );
nand ( n19596 , n19594 , n19595 );
not ( n19597 , n19587 );
nand ( n19598 , n19597 , n19582 );
not ( n19599 , n19598 );
nor ( n19600 , n19596 , n19599 );
nand ( n19601 , n19592 , n19600 );
nor ( n19602 , n19573 , n19601 );
nand ( n19603 , n19532 , n19556 );
or ( n19604 , n19553 , n19603 );
nand ( n19605 , n19604 , n19201 );
nand ( n19606 , n19602 , n19605 );
nor ( n19607 , n19566 , n19606 );
not ( n19608 , n19607 );
and ( n19609 , n19608 , RI15b62f10_1241);
not ( n19610 , RI15b62f10_1241);
not ( n19611 , n19610 );
nand ( n19612 , RI15b62c40_1235 , RI15b62cb8_1236);
not ( n19613 , RI15b62d30_1237);
nor ( n19614 , n19612 , n19613 );
nand ( n19615 , n19614 , RI15b62da8_1238);
not ( n19616 , RI15b62e20_1239);
nor ( n19617 , n19615 , n19616 );
nand ( n19618 , n19617 , RI15b62e98_1240);
buf ( n19619 , n19618 );
not ( n19620 , RI15b62bc8_1234);
nor ( n19621 , n19619 , n19620 );
not ( n19622 , n19621 );
or ( n19623 , n19611 , n19622 );
or ( n19624 , n19621 , n19610 );
nand ( n19625 , n19623 , n19624 );
nor ( n19626 , n19506 , n19575 );
not ( n19627 , RI15b606c0_1155);
and ( n19628 , n19626 , n19627 );
nor ( n19629 , n19506 , n19199 );
or ( n19630 , n19628 , n19629 );
and ( n19631 , n19625 , n19630 );
buf ( n19632 , n19619 );
and ( n19633 , n19632 , n19610 );
not ( n19634 , n19632 );
and ( n19635 , n19634 , RI15b62f10_1241);
nor ( n19636 , n19633 , n19635 );
buf ( n19637 , n19626 );
not ( n19638 , n19637 );
nor ( n19639 , n19638 , n19627 );
buf ( n19640 , n19639 );
buf ( n19641 , n19640 );
buf ( n19642 , n19641 );
buf ( n19643 , n19642 );
buf ( n19644 , n19643 );
buf ( n19645 , n19644 );
buf ( n19646 , n19645 );
and ( n19647 , n19636 , n19646 );
nor ( n19648 , n19609 , n19631 , n19647 );
nand ( n19649 , n19517 , n19648 );
buf ( n19650 , n19649 );
buf ( n19651 , RI15b3ea48_2);
buf ( n19652 , n19651 );
buf ( n19653 , RI15b3ea48_2);
buf ( n19654 , n19653 );
buf ( n19655 , RI15b3e9d0_1);
buf ( n19656 , n19655 );
buf ( n19657 , n19655 );
nand ( n19658 , RI15b4a370_397 , RI15b4a3e8_398);
not ( n19659 , RI15b4a460_399);
nor ( n19660 , n19658 , n19659 );
nand ( n19661 , n19660 , RI15b4a4d8_400);
not ( n19662 , RI15b4a550_401);
nor ( n19663 , n19661 , n19662 );
and ( n19664 , n19663 , RI15b4a5c8_402);
nand ( n19665 , n19664 , RI15b4a640_403);
not ( n19666 , RI15b4a6b8_404);
nor ( n19667 , n19665 , n19666 );
and ( n19668 , n19667 , RI15b4a730_405);
nand ( n19669 , n19668 , RI15b4a7a8_406);
not ( n19670 , RI15b4a820_407);
nor ( n19671 , n19669 , n19670 );
nand ( n19672 , n19671 , RI15b4a898_408);
not ( n19673 , RI15b4a910_409);
nor ( n19674 , n19672 , n19673 );
nand ( n19675 , n19674 , RI15b4a988_410);
not ( n19676 , RI15b4a2f8_396);
nor ( n19677 , n19675 , n19676 );
nand ( n19678 , n19677 , RI15b4aa00_411);
not ( n19679 , n19678 );
buf ( n19680 , n19679 );
buf ( n19681 , n19680 );
not ( n19682 , n19681 );
not ( n19683 , n19682 );
buf ( n19684 , n19683 );
not ( n19685 , n19684 );
nand ( n19686 , RI15b4aa78_412 , RI15b4aaf0_413);
not ( n19687 , RI15b4ab68_414);
nor ( n19688 , n19686 , n19687 );
and ( n19689 , n19688 , RI15b4abe0_415);
and ( n19690 , n19689 , RI15b4ac58_416);
nand ( n19691 , n19690 , RI15b4acd0_417);
not ( n19692 , RI15b4ad48_418);
nor ( n19693 , n19691 , n19692 );
and ( n19694 , n19693 , RI15b4adc0_419);
nand ( n19695 , n19694 , RI15b4ae38_420);
not ( n19696 , RI15b4aeb0_421);
nor ( n19697 , n19695 , n19696 );
nand ( n19698 , n19697 , RI15b4af28_422);
not ( n19699 , RI15b4afa0_423);
or ( n19700 , n19698 , n19699 );
nor ( n19701 , n19685 , n19700 );
and ( n19702 , n19701 , RI15b4b018_424);
not ( n19703 , n19701 );
not ( n19704 , RI15b4b018_424);
and ( n19705 , n19703 , n19704 );
nor ( n19706 , n19702 , n19705 );
not ( n19707 , n19706 );
not ( n19708 , n19683 );
not ( n19709 , n19697 );
nor ( n19710 , n19708 , n19709 );
and ( n19711 , n19710 , RI15b4af28_422);
not ( n19712 , n19710 );
not ( n19713 , RI15b4af28_422);
and ( n19714 , n19712 , n19713 );
nor ( n19715 , n19711 , n19714 );
not ( n19716 , n19715 );
not ( n19717 , RI15b4aa78_412);
and ( n19718 , n19679 , n19717 );
not ( n19719 , n19679 );
and ( n19720 , n19719 , RI15b4aa78_412);
nor ( n19721 , n19718 , n19720 );
nand ( n19722 , RI15b4a2f8_396 , RI15b4a370_397);
not ( n19723 , n19722 );
not ( n19724 , RI15b4a3e8_398);
and ( n19725 , n19723 , n19724 );
and ( n19726 , n19722 , RI15b4a3e8_398);
nor ( n19727 , n19725 , n19726 );
not ( n19728 , n19722 );
not ( n19729 , RI15b4a280_395);
and ( n19730 , n19728 , n19729 );
nand ( n19731 , n19727 , n19730 );
not ( n19732 , RI15b4a460_399);
not ( n19733 , n19732 );
buf ( n19734 , n19658 );
nor ( n19735 , n19734 , n19676 );
not ( n19736 , n19735 );
or ( n19737 , n19733 , n19736 );
not ( n19738 , RI15b4a460_399);
or ( n19739 , n19735 , n19738 );
nand ( n19740 , n19737 , n19739 );
nor ( n19741 , n19731 , n19740 );
buf ( n19742 , n19660 );
nand ( n19743 , n19742 , RI15b4a2f8_396);
and ( n19744 , n19743 , RI15b4a4d8_400);
not ( n19745 , n19743 );
not ( n19746 , RI15b4a4d8_400);
and ( n19747 , n19745 , n19746 );
nor ( n19748 , n19744 , n19747 );
nand ( n19749 , n19741 , n19748 );
not ( n19750 , n19662 );
buf ( n19751 , n19661 );
nor ( n19752 , n19751 , n19676 );
not ( n19753 , n19752 );
or ( n19754 , n19750 , n19753 );
or ( n19755 , n19752 , n19662 );
nand ( n19756 , n19754 , n19755 );
nor ( n19757 , n19749 , n19756 );
buf ( n19758 , n19663 );
nand ( n19759 , n19758 , RI15b4a2f8_396);
and ( n19760 , n19759 , RI15b4a5c8_402);
not ( n19761 , n19759 );
not ( n19762 , RI15b4a5c8_402);
and ( n19763 , n19761 , n19762 );
nor ( n19764 , n19760 , n19763 );
nand ( n19765 , n19757 , n19764 );
not ( n19766 , RI15b4a640_403);
not ( n19767 , n19766 );
not ( n19768 , n19664 );
nor ( n19769 , n19768 , n19676 );
not ( n19770 , n19769 );
or ( n19771 , n19767 , n19770 );
or ( n19772 , n19769 , n19766 );
nand ( n19773 , n19771 , n19772 );
nor ( n19774 , n19765 , n19773 );
not ( n19775 , n19665 );
nand ( n19776 , n19775 , RI15b4a2f8_396);
and ( n19777 , n19776 , RI15b4a6b8_404);
not ( n19778 , n19776 );
and ( n19779 , n19778 , n19666 );
nor ( n19780 , n19777 , n19779 );
and ( n19781 , n19774 , n19780 );
buf ( n19782 , n19667 );
nand ( n19783 , n19782 , RI15b4a2f8_396);
and ( n19784 , n19783 , RI15b4a730_405);
not ( n19785 , n19783 );
not ( n19786 , RI15b4a730_405);
and ( n19787 , n19785 , n19786 );
nor ( n19788 , n19784 , n19787 );
nand ( n19789 , n19781 , n19788 );
not ( n19790 , RI15b4a7a8_406);
not ( n19791 , n19790 );
not ( n19792 , n19668 );
nor ( n19793 , n19792 , n19676 );
not ( n19794 , n19793 );
or ( n19795 , n19791 , n19794 );
or ( n19796 , n19793 , n19790 );
nand ( n19797 , n19795 , n19796 );
nor ( n19798 , n19789 , n19797 );
not ( n19799 , n19669 );
nand ( n19800 , n19799 , RI15b4a2f8_396);
and ( n19801 , n19800 , RI15b4a820_407);
not ( n19802 , n19800 );
and ( n19803 , n19802 , n19670 );
nor ( n19804 , n19801 , n19803 );
nand ( n19805 , n19798 , n19804 );
nand ( n19806 , n19671 , RI15b4a2f8_396);
xnor ( n19807 , n19806 , RI15b4a898_408);
nor ( n19808 , n19805 , n19807 );
not ( n19809 , n19672 );
nand ( n19810 , n19809 , RI15b4a2f8_396);
and ( n19811 , n19810 , RI15b4a910_409);
not ( n19812 , n19810 );
and ( n19813 , n19812 , n19673 );
nor ( n19814 , n19811 , n19813 );
and ( n19815 , n19808 , n19814 );
buf ( n19816 , n19674 );
nand ( n19817 , n19816 , RI15b4a2f8_396);
and ( n19818 , n19817 , RI15b4a988_410);
not ( n19819 , n19817 );
not ( n19820 , RI15b4a988_410);
and ( n19821 , n19819 , n19820 );
nor ( n19822 , n19818 , n19821 );
nand ( n19823 , n19815 , n19822 );
not ( n19824 , RI15b4aa00_411);
not ( n19825 , n19824 );
buf ( n19826 , n19677 );
not ( n19827 , n19826 );
or ( n19828 , n19825 , n19827 );
or ( n19829 , n19826 , n19824 );
nand ( n19830 , n19828 , n19829 );
nor ( n19831 , n19823 , n19830 );
nand ( n19832 , n19721 , n19831 );
not ( n19833 , RI15b4aaf0_413);
nand ( n19834 , n19679 , RI15b4aa78_412);
not ( n19835 , n19834 );
or ( n19836 , n19833 , n19835 );
or ( n19837 , n19834 , RI15b4aaf0_413);
nand ( n19838 , n19836 , n19837 );
nor ( n19839 , n19832 , n19838 );
buf ( n19840 , n19679 );
not ( n19841 , n19686 );
nand ( n19842 , n19840 , n19841 );
and ( n19843 , n19842 , RI15b4ab68_414);
not ( n19844 , n19842 );
and ( n19845 , n19844 , n19687 );
nor ( n19846 , n19843 , n19845 );
nand ( n19847 , n19839 , n19846 );
not ( n19848 , n19688 );
not ( n19849 , n19848 );
nand ( n19850 , n19849 , n19680 );
not ( n19851 , RI15b4abe0_415);
and ( n19852 , n19850 , n19851 );
not ( n19853 , n19850 );
and ( n19854 , n19853 , RI15b4abe0_415);
nor ( n19855 , n19852 , n19854 );
nor ( n19856 , n19847 , n19855 );
not ( n19857 , n19689 );
not ( n19858 , n19857 );
nand ( n19859 , n19858 , n19680 );
xor ( n19860 , n19859 , RI15b4ac58_416);
and ( n19861 , n19856 , n19860 );
buf ( n19862 , n19690 );
nand ( n19863 , n19681 , n19862 );
and ( n19864 , n19863 , RI15b4acd0_417);
not ( n19865 , n19863 );
not ( n19866 , RI15b4acd0_417);
and ( n19867 , n19865 , n19866 );
nor ( n19868 , n19864 , n19867 );
nand ( n19869 , n19861 , n19868 );
not ( n19870 , n19691 );
nand ( n19871 , n19870 , n19681 );
and ( n19872 , n19871 , n19692 );
not ( n19873 , n19871 );
and ( n19874 , n19873 , RI15b4ad48_418);
nor ( n19875 , n19872 , n19874 );
nor ( n19876 , n19869 , n19875 );
nand ( n19877 , n19681 , n19693 );
and ( n19878 , n19877 , RI15b4adc0_419);
not ( n19879 , n19877 );
not ( n19880 , RI15b4adc0_419);
and ( n19881 , n19879 , n19880 );
nor ( n19882 , n19878 , n19881 );
and ( n19883 , n19876 , n19882 );
not ( n19884 , n19694 );
nor ( n19885 , n19682 , n19884 );
not ( n19886 , RI15b4ae38_420);
and ( n19887 , n19885 , n19886 );
not ( n19888 , n19885 );
and ( n19889 , n19888 , RI15b4ae38_420);
nor ( n19890 , n19887 , n19889 );
nand ( n19891 , n19883 , n19890 );
not ( n19892 , n19695 );
nand ( n19893 , n19892 , n19683 );
and ( n19894 , n19893 , n19696 );
not ( n19895 , n19893 );
and ( n19896 , n19895 , RI15b4aeb0_421);
nor ( n19897 , n19894 , n19896 );
nor ( n19898 , n19891 , n19897 );
nand ( n19899 , n19716 , n19898 );
not ( n19900 , n19698 );
nand ( n19901 , n19900 , n19684 );
and ( n19902 , n19901 , n19699 );
not ( n19903 , n19901 );
and ( n19904 , n19903 , RI15b4afa0_423);
nor ( n19905 , n19902 , n19904 );
nor ( n19906 , n19899 , n19905 );
nand ( n19907 , n19707 , n19906 );
not ( n19908 , RI15b44d30_213);
nor ( n19909 , n19908 , RI15b44cb8_212);
nor ( n19910 , RI15b44da8_214 , RI15b44e20_215);
nand ( n19911 , n19909 , n19910 );
not ( n19912 , n19911 );
not ( n19913 , RI15b47df0_317);
nand ( n19914 , n19912 , n19913 );
buf ( n19915 , n19914 );
buf ( n19916 , n19915 );
buf ( n19917 , n19916 );
buf ( n19918 , n19917 );
buf ( n19919 , n19918 );
not ( n19920 , n19919 );
not ( n19921 , n19920 );
buf ( n19922 , n19921 );
nor ( n19923 , n19907 , n19922 );
or ( n19924 , n19700 , n19704 );
not ( n19925 , RI15b4b090_425);
or ( n19926 , n19924 , n19925 );
not ( n19927 , n19926 );
nand ( n19928 , n19927 , n19681 );
and ( n19929 , n19928 , RI15b4b108_426);
not ( n19930 , n19928 );
not ( n19931 , RI15b4b108_426);
and ( n19932 , n19930 , n19931 );
nor ( n19933 , n19929 , n19932 );
buf ( n19934 , n19916 );
not ( n19935 , n19934 );
nand ( n19936 , n19933 , n19935 );
not ( n19937 , n19936 );
not ( n19938 , n19937 );
not ( n19939 , n19938 );
not ( n19940 , n19939 );
not ( n19941 , n19940 );
not ( n19942 , n19941 );
not ( n19943 , n19942 );
buf ( n19944 , n19943 );
or ( n19945 , n19923 , n19944 );
not ( n19946 , n19924 );
nand ( n19947 , n19946 , n19684 );
and ( n19948 , n19947 , n19925 );
not ( n19949 , n19947 );
and ( n19950 , n19949 , RI15b4b090_425);
nor ( n19951 , n19948 , n19950 );
nand ( n19952 , n19945 , n19951 );
not ( n19953 , RI15b4a0a0_391);
nor ( n19954 , RI15b49380_363 , RI15b493f8_364);
not ( n19955 , RI15b49470_365);
and ( n19956 , n19954 , n19955 );
not ( n19957 , RI15b494e8_366);
nand ( n19958 , n19956 , n19957 );
nor ( n19959 , n19958 , RI15b49560_367);
not ( n19960 , RI15b495d8_368);
and ( n19961 , n19959 , n19960 );
not ( n19962 , RI15b49650_369);
nand ( n19963 , n19961 , n19962 );
nor ( n19964 , n19963 , RI15b496c8_370);
not ( n19965 , RI15b49740_371);
and ( n19966 , n19964 , n19965 );
not ( n19967 , RI15b497b8_372);
nand ( n19968 , n19966 , n19967 );
nor ( n19969 , n19968 , RI15b49830_373);
not ( n19970 , RI15b498a8_374);
and ( n19971 , n19969 , n19970 );
not ( n19972 , RI15b49920_375);
nand ( n19973 , n19971 , n19972 );
nor ( n19974 , n19973 , RI15b49998_376);
not ( n19975 , RI15b49a10_377);
and ( n19976 , n19974 , n19975 );
not ( n19977 , RI15b49a88_378);
nand ( n19978 , n19976 , n19977 );
nor ( n19979 , n19978 , RI15b49b00_379);
not ( n19980 , RI15b49b78_380);
nand ( n19981 , n19979 , n19980 );
nor ( n19982 , n19981 , RI15b49bf0_381);
not ( n19983 , RI15b49c68_382);
and ( n19984 , n19982 , n19983 );
not ( n19985 , RI15b49ce0_383);
nand ( n19986 , n19984 , n19985 );
nor ( n19987 , n19986 , RI15b49d58_384);
not ( n19988 , RI15b49dd0_385);
and ( n19989 , n19987 , n19988 );
not ( n19990 , RI15b49e48_386);
nand ( n19991 , n19989 , n19990 );
nor ( n19992 , n19991 , RI15b49ec0_387);
not ( n19993 , RI15b49f38_388);
and ( n19994 , n19992 , n19993 );
not ( n19995 , RI15b49fb0_389);
nand ( n19996 , n19994 , n19995 );
nor ( n19997 , n19996 , RI15b4a028_390);
nand ( n19998 , n19953 , n19997 );
nor ( n19999 , n19998 , RI15b4a118_392);
not ( n20000 , n19999 );
not ( n20001 , RI15b42918_136);
nand ( n20002 , RI15b449e8_206 , RI15b44a60_207);
not ( n20003 , n20002 );
not ( n20004 , RI15b44b50_209);
nor ( n20005 , n20004 , RI15b44ad8_208);
nand ( n20006 , n20003 , n20005 );
not ( n20007 , n20006 );
not ( n20008 , RI15b44bc8_210);
nand ( n20009 , n20007 , n20008 );
not ( n20010 , n20009 );
not ( n20011 , n20010 );
or ( n20012 , n20001 , n20011 );
not ( n20013 , RI15b44a60_207);
nand ( n20014 , n20013 , RI15b449e8_206);
not ( n20015 , n20014 );
not ( n20016 , RI15b44b50_209);
nand ( n20017 , n20016 , RI15b44ad8_208);
not ( n20018 , n20017 );
nand ( n20019 , n20015 , n20018 );
not ( n20020 , n20019 );
nand ( n20021 , n20020 , n20008 );
not ( n20022 , n20021 );
nand ( n20023 , n20022 , RI15b41298_88);
nand ( n20024 , n20012 , n20023 );
nor ( n20025 , RI15b449e8_206 , RI15b44a60_207);
nand ( n20026 , n20025 , n20018 );
not ( n20027 , n20026 );
nand ( n20028 , n20027 , n20008 );
not ( n20029 , n20028 );
nand ( n20030 , n20029 , RI15b40ed8_80);
not ( n20031 , RI15b449e8_206);
nand ( n20032 , n20031 , RI15b44a60_207);
not ( n20033 , n20032 );
not ( n20034 , n20033 );
not ( n20035 , n20018 );
nor ( n20036 , n20034 , n20035 );
nand ( n20037 , n20036 , n20008 );
not ( n20038 , n20037 );
nand ( n20039 , n20038 , RI15b41658_96);
nor ( n20040 , RI15b44ad8_208 , RI15b44b50_209);
nand ( n20041 , n20033 , n20040 );
not ( n20042 , n20041 );
nand ( n20043 , n20042 , n20008 );
not ( n20044 , n20043 );
nand ( n20045 , n20044 , RI15b40758_64);
nand ( n20046 , n20030 , n20039 , n20045 );
nor ( n20047 , n20024 , n20046 );
nand ( n20048 , n20003 , n20018 );
not ( n20049 , n20048 );
nand ( n20050 , n20049 , n20008 );
not ( n20051 , n20050 );
and ( n20052 , n20051 , RI15b41a18_104);
not ( n20053 , RI15b42198_120);
not ( n20054 , n20014 );
buf ( n20055 , n20005 );
nand ( n20056 , n20054 , n20055 );
nor ( n20057 , n20056 , RI15b44bc8_210);
not ( n20058 , n20057 );
or ( n20059 , n20053 , n20058 );
nand ( n20060 , n20033 , n20005 );
not ( n20061 , n20060 );
nand ( n20062 , n20061 , n20008 );
not ( n20063 , n20062 );
nand ( n20064 , n20063 , RI15b42558_128);
nand ( n20065 , n20059 , n20064 );
nor ( n20066 , n20052 , n20065 );
nand ( n20067 , RI15b44ad8_208 , RI15b44b50_209);
nor ( n20068 , n20067 , RI15b44bc8_210);
not ( n20069 , n20068 );
not ( n20070 , n20069 );
nor ( n20071 , RI15b449e8_206 , RI15b44a60_207);
buf ( n20072 , n20071 );
nand ( n20073 , n20070 , n20072 );
not ( n20074 , n20073 );
not ( n20075 , RI15b42cd8_144);
not ( n20076 , n20075 );
and ( n20077 , n20074 , n20076 );
not ( n20078 , n20068 );
not ( n20079 , n20078 );
not ( n20080 , n20014 );
nand ( n20081 , n20079 , n20080 );
not ( n20082 , RI15b43098_152);
nor ( n20083 , n20081 , n20082 );
nor ( n20084 , n20077 , n20083 );
not ( n20085 , n20033 );
or ( n20086 , n20069 , n20085 );
not ( n20087 , n20086 );
and ( n20088 , n20087 , RI15b43458_160);
and ( n20089 , n20068 , n20003 );
and ( n20090 , n20089 , RI15b43818_168);
nor ( n20091 , n20088 , n20090 );
nand ( n20092 , n20072 , n20005 );
nor ( n20093 , n20092 , RI15b44bc8_210);
buf ( n20094 , n20093 );
nand ( n20095 , n20094 , RI15b41dd8_112);
not ( n20096 , n20003 );
not ( n20097 , n20040 );
nor ( n20098 , n20096 , n20097 );
nand ( n20099 , n20098 , n20008 );
not ( n20100 , n20099 );
nand ( n20101 , n20100 , RI15b40b18_72);
nand ( n20102 , n20084 , n20091 , n20095 , n20101 );
not ( n20103 , n20102 );
not ( n20104 , n20097 );
nand ( n20105 , n20054 , n20104 );
nor ( n20106 , n20105 , RI15b44bc8_210);
and ( n20107 , n20106 , RI15b40398_56);
not ( n20108 , n20071 );
not ( n20109 , n20108 );
nand ( n20110 , n20109 , n20040 );
not ( n20111 , n20110 );
nand ( n20112 , n20111 , n20008 );
not ( n20113 , RI15b3ffd8_48);
nor ( n20114 , n20112 , n20113 );
nor ( n20115 , n20107 , n20114 );
nand ( n20116 , n20047 , n20066 , n20103 , n20115 );
not ( n20117 , n20116 );
not ( n20118 , n20081 );
not ( n20119 , RI15b432f0_157);
not ( n20120 , n20119 );
and ( n20121 , n20118 , n20120 );
not ( n20122 , n20073 );
and ( n20123 , n20122 , RI15b42f30_149);
nor ( n20124 , n20121 , n20123 );
not ( n20125 , n20089 );
not ( n20126 , n20125 );
not ( n20127 , RI15b43a70_173);
not ( n20128 , n20127 );
and ( n20129 , n20126 , n20128 );
not ( n20130 , n20086 );
and ( n20131 , n20130 , RI15b436b0_165);
nor ( n20132 , n20129 , n20131 );
buf ( n20133 , n20093 );
nand ( n20134 , n20133 , RI15b42030_117);
not ( n20135 , n20099 );
nand ( n20136 , n20135 , RI15b40d70_77);
nand ( n20137 , n20124 , n20132 , n20134 , n20136 );
not ( n20138 , RI15b405f0_61);
not ( n20139 , n20106 );
or ( n20140 , n20138 , n20139 );
not ( n20141 , n20112 );
nand ( n20142 , n20141 , RI15b40230_53);
nand ( n20143 , n20140 , n20142 );
nor ( n20144 , n20137 , n20143 );
not ( n20145 , RI15b42b70_141);
not ( n20146 , n20009 );
not ( n20147 , n20146 );
or ( n20148 , n20145 , n20147 );
nand ( n20149 , n20022 , RI15b414f0_93);
nand ( n20150 , n20148 , n20149 );
not ( n20151 , n20028 );
nand ( n20152 , n20151 , RI15b41130_85);
nand ( n20153 , n20038 , RI15b418b0_101);
not ( n20154 , n20043 );
nand ( n20155 , n20154 , RI15b409b0_69);
nand ( n20156 , n20152 , n20153 , n20155 );
nor ( n20157 , n20150 , n20156 );
not ( n20158 , n20050 );
and ( n20159 , n20158 , RI15b41c70_109);
not ( n20160 , RI15b423f0_125);
not ( n20161 , n20057 );
or ( n20162 , n20160 , n20161 );
not ( n20163 , n20062 );
nand ( n20164 , n20163 , RI15b427b0_133);
nand ( n20165 , n20162 , n20164 );
nor ( n20166 , n20159 , n20165 );
nand ( n20167 , n20144 , n20157 , n20166 );
not ( n20168 , n20081 );
not ( n20169 , RI15b43110_153);
not ( n20170 , n20169 );
and ( n20171 , n20168 , n20170 );
and ( n20172 , n20122 , RI15b42d50_145);
nor ( n20173 , n20171 , n20172 );
not ( n20174 , n20125 );
not ( n20175 , RI15b43890_169);
not ( n20176 , n20175 );
and ( n20177 , n20174 , n20176 );
and ( n20178 , n20130 , RI15b434d0_161);
nor ( n20179 , n20177 , n20178 );
nand ( n20180 , n20133 , RI15b41e50_113);
not ( n20181 , n20099 );
nand ( n20182 , n20181 , RI15b40b90_73);
nand ( n20183 , n20173 , n20179 , n20180 , n20182 );
not ( n20184 , RI15b40410_57);
not ( n20185 , n20106 );
or ( n20186 , n20184 , n20185 );
nand ( n20187 , n20141 , RI15b40050_49);
nand ( n20188 , n20186 , n20187 );
nor ( n20189 , n20183 , n20188 );
not ( n20190 , RI15b42990_137);
not ( n20191 , n20146 );
or ( n20192 , n20190 , n20191 );
nand ( n20193 , n20022 , RI15b41310_89);
nand ( n20194 , n20192 , n20193 );
not ( n20195 , n20028 );
nand ( n20196 , n20195 , RI15b40f50_81);
nand ( n20197 , n20038 , RI15b416d0_97);
nand ( n20198 , n20154 , RI15b407d0_65);
nand ( n20199 , n20196 , n20197 , n20198 );
nor ( n20200 , n20194 , n20199 );
and ( n20201 , n20158 , RI15b41a90_105);
not ( n20202 , RI15b42210_121);
not ( n20203 , n20057 );
or ( n20204 , n20202 , n20203 );
nand ( n20205 , n20163 , RI15b425d0_129);
nand ( n20206 , n20204 , n20205 );
nor ( n20207 , n20201 , n20206 );
nand ( n20208 , n20189 , n20200 , n20207 );
nand ( n20209 , n20117 , n20167 , n20208 );
not ( n20210 , n20209 );
not ( n20211 , RI15b42828_134);
not ( n20212 , n20146 );
or ( n20213 , n20211 , n20212 );
nand ( n20214 , n20022 , RI15b411a8_86);
nand ( n20215 , n20213 , n20214 );
nand ( n20216 , n20195 , RI15b40de8_78);
nand ( n20217 , n20038 , RI15b41568_94);
not ( n20218 , n20043 );
nand ( n20219 , n20218 , RI15b40668_62);
nand ( n20220 , n20216 , n20217 , n20219 );
nor ( n20221 , n20215 , n20220 );
and ( n20222 , n20158 , RI15b41928_102);
not ( n20223 , RI15b420a8_118);
nor ( n20224 , n20056 , RI15b44bc8_210);
not ( n20225 , n20224 );
or ( n20226 , n20223 , n20225 );
nand ( n20227 , n20163 , RI15b42468_126);
nand ( n20228 , n20226 , n20227 );
nor ( n20229 , n20222 , n20228 );
not ( n20230 , n20073 );
not ( n20231 , RI15b42be8_142);
not ( n20232 , n20231 );
and ( n20233 , n20230 , n20232 );
not ( n20234 , RI15b42fa8_150);
nor ( n20235 , n20081 , n20234 );
nor ( n20236 , n20233 , n20235 );
not ( n20237 , n20086 );
and ( n20238 , n20237 , RI15b43368_158);
not ( n20239 , n20125 );
and ( n20240 , n20239 , RI15b43728_166);
nor ( n20241 , n20238 , n20240 );
nand ( n20242 , n20133 , RI15b41ce8_110);
nand ( n20243 , n20135 , RI15b40a28_70);
nand ( n20244 , n20236 , n20241 , n20242 , n20243 );
not ( n20245 , n20244 );
nor ( n20246 , n20105 , RI15b44bc8_210);
and ( n20247 , n20246 , RI15b402a8_54);
not ( n20248 , RI15b3fee8_46);
nor ( n20249 , n20112 , n20248 );
nor ( n20250 , n20247 , n20249 );
nand ( n20251 , n20221 , n20229 , n20245 , n20250 );
not ( n20252 , n20251 );
not ( n20253 , RI15b42a08_138);
not ( n20254 , n20009 );
not ( n20255 , n20254 );
or ( n20256 , n20253 , n20255 );
nand ( n20257 , n20022 , RI15b41388_90);
nand ( n20258 , n20256 , n20257 );
nand ( n20259 , n20195 , RI15b40fc8_82);
nand ( n20260 , n20038 , RI15b41748_98);
nand ( n20261 , n20218 , RI15b40848_66);
nand ( n20262 , n20259 , n20260 , n20261 );
nor ( n20263 , n20258 , n20262 );
and ( n20264 , n20158 , RI15b41b08_106);
not ( n20265 , RI15b42288_122);
not ( n20266 , n20224 );
or ( n20267 , n20265 , n20266 );
not ( n20268 , n20062 );
nand ( n20269 , n20268 , RI15b42648_130);
nand ( n20270 , n20267 , n20269 );
nor ( n20271 , n20264 , n20270 );
not ( n20272 , n20073 );
not ( n20273 , RI15b42dc8_146);
not ( n20274 , n20273 );
and ( n20275 , n20272 , n20274 );
not ( n20276 , RI15b43188_154);
nor ( n20277 , n20081 , n20276 );
nor ( n20278 , n20275 , n20277 );
and ( n20279 , n20237 , RI15b43548_162);
not ( n20280 , n20125 );
and ( n20281 , n20280 , RI15b43908_170);
nor ( n20282 , n20279 , n20281 );
nand ( n20283 , n20133 , RI15b41ec8_114);
nand ( n20284 , n20135 , RI15b40c08_74);
and ( n20285 , n20278 , n20282 , n20283 , n20284 );
not ( n20286 , n20112 );
not ( n20287 , RI15b400c8_50);
not ( n20288 , n20287 );
and ( n20289 , n20286 , n20288 );
and ( n20290 , n20246 , RI15b40488_58);
nor ( n20291 , n20289 , n20290 );
nand ( n20292 , n20263 , n20271 , n20285 , n20291 );
nor ( n20293 , n20252 , n20292 );
nand ( n20294 , n20210 , n20293 );
not ( n20295 , RI15b428a0_135);
not ( n20296 , n20254 );
or ( n20297 , n20295 , n20296 );
nand ( n20298 , n20022 , RI15b41220_87);
nand ( n20299 , n20297 , n20298 );
nand ( n20300 , n20151 , RI15b40e60_79);
nand ( n20301 , n20038 , RI15b415e0_95);
nand ( n20302 , n20218 , RI15b406e0_63);
nand ( n20303 , n20300 , n20301 , n20302 );
nor ( n20304 , n20299 , n20303 );
not ( n20305 , n20050 );
and ( n20306 , n20305 , RI15b419a0_103);
not ( n20307 , RI15b42120_119);
not ( n20308 , n20224 );
or ( n20309 , n20307 , n20308 );
nand ( n20310 , n20268 , RI15b424e0_127);
nand ( n20311 , n20309 , n20310 );
nor ( n20312 , n20306 , n20311 );
not ( n20313 , n20073 );
not ( n20314 , RI15b42c60_143);
not ( n20315 , n20314 );
and ( n20316 , n20313 , n20315 );
not ( n20317 , RI15b43020_151);
nor ( n20318 , n20081 , n20317 );
nor ( n20319 , n20316 , n20318 );
and ( n20320 , n20237 , RI15b433e0_159);
and ( n20321 , n20280 , RI15b437a0_167);
nor ( n20322 , n20320 , n20321 );
nand ( n20323 , n20133 , RI15b41d60_111);
nand ( n20324 , n20135 , RI15b40aa0_71);
and ( n20325 , n20319 , n20322 , n20323 , n20324 );
not ( n20326 , n20112 );
not ( n20327 , RI15b3ff60_47);
not ( n20328 , n20327 );
and ( n20329 , n20326 , n20328 );
and ( n20330 , n20246 , RI15b40320_55);
nor ( n20331 , n20329 , n20330 );
nand ( n20332 , n20304 , n20312 , n20325 , n20331 );
not ( n20333 , n20073 );
not ( n20334 , RI15b42e40_147);
not ( n20335 , n20334 );
and ( n20336 , n20333 , n20335 );
not ( n20337 , RI15b43200_155);
nor ( n20338 , n20081 , n20337 );
nor ( n20339 , n20336 , n20338 );
not ( n20340 , n20125 );
not ( n20341 , RI15b43980_171);
not ( n20342 , n20341 );
and ( n20343 , n20340 , n20342 );
and ( n20344 , n20237 , RI15b435c0_163);
nor ( n20345 , n20343 , n20344 );
nand ( n20346 , n20133 , RI15b41f40_115);
nand ( n20347 , n20135 , RI15b40c80_75);
nand ( n20348 , n20339 , n20345 , n20346 , n20347 );
not ( n20349 , RI15b40500_59);
not ( n20350 , n20106 );
or ( n20351 , n20349 , n20350 );
nand ( n20352 , n20141 , RI15b40140_51);
nand ( n20353 , n20351 , n20352 );
nor ( n20354 , n20348 , n20353 );
and ( n20355 , n20305 , RI15b41b80_107);
not ( n20356 , RI15b42300_123);
not ( n20357 , n20224 );
or ( n20358 , n20356 , n20357 );
nand ( n20359 , n20163 , RI15b426c0_131);
nand ( n20360 , n20358 , n20359 );
nor ( n20361 , n20355 , n20360 );
not ( n20362 , n20021 );
not ( n20363 , RI15b41400_91);
not ( n20364 , n20363 );
and ( n20365 , n20362 , n20364 );
and ( n20366 , n20254 , RI15b42a80_139);
nor ( n20367 , n20365 , n20366 );
not ( n20368 , RI15b417c0_99);
not ( n20369 , n20038 );
or ( n20370 , n20368 , n20369 );
nand ( n20371 , n20218 , RI15b408c0_67);
nand ( n20372 , n20370 , n20371 );
and ( n20373 , n20151 , RI15b41040_83);
nor ( n20374 , n20372 , n20373 );
nand ( n20375 , n20354 , n20361 , n20367 , n20374 );
not ( n20376 , n20375 );
not ( n20377 , RI15b42af8_140);
not ( n20378 , n20146 );
or ( n20379 , n20377 , n20378 );
nand ( n20380 , n20022 , RI15b41478_92);
nand ( n20381 , n20379 , n20380 );
nand ( n20382 , n20195 , RI15b410b8_84);
nand ( n20383 , n20038 , RI15b41838_100);
nand ( n20384 , n20154 , RI15b40938_68);
nand ( n20385 , n20382 , n20383 , n20384 );
nor ( n20386 , n20381 , n20385 );
and ( n20387 , n20305 , RI15b41bf8_108);
not ( n20388 , RI15b42378_124);
not ( n20389 , n20057 );
or ( n20390 , n20388 , n20389 );
nand ( n20391 , n20268 , RI15b42738_132);
nand ( n20392 , n20390 , n20391 );
nor ( n20393 , n20387 , n20392 );
not ( n20394 , n20073 );
not ( n20395 , RI15b42eb8_148);
not ( n20396 , n20395 );
and ( n20397 , n20394 , n20396 );
not ( n20398 , RI15b43278_156);
nor ( n20399 , n20081 , n20398 );
nor ( n20400 , n20397 , n20399 );
and ( n20401 , n20130 , RI15b43638_164);
and ( n20402 , n20089 , RI15b439f8_172);
nor ( n20403 , n20401 , n20402 );
nand ( n20404 , n20133 , RI15b41fb8_116);
nand ( n20405 , n20181 , RI15b40cf8_76);
nand ( n20406 , n20400 , n20403 , n20404 , n20405 );
not ( n20407 , n20406 );
and ( n20408 , n20246 , RI15b40578_60);
not ( n20409 , RI15b401b8_52);
nor ( n20410 , n20112 , n20409 );
nor ( n20411 , n20408 , n20410 );
nand ( n20412 , n20386 , n20393 , n20407 , n20411 );
not ( n20413 , n20412 );
nand ( n20414 , n20332 , n20376 , n20413 );
nor ( n20415 , n20294 , n20414 );
buf ( n20416 , n20415 );
not ( n20417 , RI15b3fd80_43);
nand ( n20418 , n20417 , RI15b44ad8_208);
not ( n20419 , n20418 );
not ( n20420 , n20108 );
not ( n20421 , n20420 );
not ( n20422 , RI15b3fc90_41);
not ( n20423 , RI15b3fd08_42);
nand ( n20424 , n20422 , n20423 );
not ( n20425 , RI15b44a60_207);
and ( n20426 , n20424 , n20425 );
and ( n20427 , RI15b3fc90_41 , RI15b3fd08_42);
nor ( n20428 , n20426 , n20427 );
not ( n20429 , RI15b449e8_206);
nand ( n20430 , n20429 , RI15b3fd08_42);
nand ( n20431 , n20421 , n20428 , n20430 );
not ( n20432 , n20431 );
or ( n20433 , n20419 , n20432 );
not ( n20434 , RI15b44ad8_208);
nand ( n20435 , n20434 , RI15b3fd80_43);
nand ( n20436 , n20433 , n20435 );
nand ( n20437 , n20008 , RI15b3fe70_45);
not ( n20438 , RI15b44b50_209);
nand ( n20439 , n20438 , RI15b3fdf8_44);
not ( n20440 , RI15b3fdf8_44);
nand ( n20441 , n20440 , RI15b44b50_209);
nand ( n20442 , n20437 , n20439 , n20441 );
nand ( n20443 , n20436 , n20442 );
not ( n20444 , n20443 );
not ( n20445 , RI15b3fe70_45);
not ( n20446 , n20440 );
not ( n20447 , n20436 );
or ( n20448 , n20446 , n20447 );
nand ( n20449 , RI15b3fdf8_44 , RI15b44bc8_210);
nand ( n20450 , n20448 , n20449 );
not ( n20451 , n20450 );
or ( n20452 , n20445 , n20451 );
nor ( n20453 , n20436 , RI15b3fdf8_44);
or ( n20454 , n20453 , RI15b3fe70_45);
nand ( n20455 , n20454 , n20441 );
nand ( n20456 , n20455 , n20008 );
nand ( n20457 , n20452 , n20456 );
not ( n20458 , n20457 );
or ( n20459 , n20444 , n20458 );
not ( n20460 , RI15b44bc8_210);
not ( n20461 , RI15b3fe70_45);
not ( n20462 , n20461 );
or ( n20463 , n20460 , n20462 );
not ( n20464 , n20441 );
not ( n20465 , n20436 );
or ( n20466 , n20464 , n20465 );
nand ( n20467 , n20466 , n20439 );
nand ( n20468 , n20463 , n20467 );
nand ( n20469 , n20468 , n20437 );
nand ( n20470 , n20459 , n20469 );
not ( n20471 , n20431 );
not ( n20472 , n20471 );
nand ( n20473 , n20435 , n20418 );
not ( n20474 , n20473 );
and ( n20475 , n20472 , n20474 );
and ( n20476 , n20471 , n20473 );
nor ( n20477 , n20475 , n20476 );
nand ( n20478 , n20469 , n20477 );
nand ( n20479 , n20422 , RI15b449e8_206);
not ( n20480 , n20479 );
and ( n20481 , n20425 , n20423 );
and ( n20482 , RI15b3fd08_42 , RI15b44a60_207);
nor ( n20483 , n20481 , n20482 );
not ( n20484 , n20483 );
or ( n20485 , n20480 , n20484 );
or ( n20486 , n20479 , n20483 );
nand ( n20487 , n20485 , n20486 );
nand ( n20488 , n20469 , n20487 );
nand ( n20489 , n20470 , n20478 , n20488 );
not ( n20490 , n20489 );
nand ( n20491 , RI15b3fba0_39 , RI15b668b8_1364);
not ( n20492 , n20491 );
nor ( n20493 , n20492 , RI15b47df0_317);
nor ( n20494 , n20490 , n20493 );
nand ( n20495 , n20416 , n20494 );
not ( n20496 , n20495 );
not ( n20497 , RI15b44da8_214);
nor ( n20498 , n20497 , RI15b44e20_215);
not ( n20499 , RI15b44cb8_212);
nor ( n20500 , n20499 , RI15b44d30_213);
and ( n20501 , n20498 , n20500 );
nand ( n20502 , n20496 , n20501 );
nor ( n20503 , n20000 , n20502 );
nor ( n20504 , n20502 , RI15b4a208_394);
not ( n20505 , n20294 );
nor ( n20506 , n20375 , n20412 );
not ( n20507 , n20332 );
and ( n20508 , n20506 , n20507 );
nand ( n20509 , n20505 , n20508 );
not ( n20510 , n20509 );
not ( n20511 , n20490 );
buf ( n20512 , n20511 );
and ( n20513 , RI15b48390_329 , RI15b48408_330);
nor ( n20514 , RI15b48390_329 , RI15b48408_330);
nor ( n20515 , n20513 , n20514 , RI15b48318_328);
nand ( n20516 , n20515 , n20491 );
or ( n20517 , n20516 , RI15b47df0_317);
nand ( n20518 , n20510 , n20512 , n20517 );
not ( n20519 , n20501 );
nor ( n20520 , n20518 , n20519 );
or ( n20521 , n20504 , n20520 );
or ( n20522 , n20503 , n20521 );
nand ( n20523 , n20522 , RI15b4a190_393);
nor ( n20524 , n19933 , n19917 );
not ( n20525 , n20524 );
nor ( n20526 , n20525 , n19951 );
nand ( n20527 , n19907 , n20526 );
not ( n20528 , RI15b4a208_394);
or ( n20529 , n20502 , n20528 );
nor ( n20530 , n20529 , RI15b4a190_393);
and ( n20531 , n20000 , n20530 );
not ( n20532 , RI15b4b2e8_430);
nand ( n20533 , RI15b4b1f8_428 , RI15b4b270_429);
nor ( n20534 , n20532 , n20533 );
and ( n20535 , RI15b4b360_431 , RI15b4b3d8_432);
nand ( n20536 , n20534 , n20535 );
nand ( n20537 , RI15b4b450_433 , RI15b4b4c8_434);
nor ( n20538 , n20536 , n20537 );
and ( n20539 , n20538 , RI15b4b540_435);
nand ( n20540 , n20539 , RI15b4b5b8_436);
not ( n20541 , n20540 );
and ( n20542 , RI15b4b630_437 , RI15b4b6a8_438);
nand ( n20543 , n20541 , n20542 );
nand ( n20544 , RI15b4b720_439 , RI15b4b798_440);
nor ( n20545 , n20543 , n20544 );
not ( n20546 , RI15b4b888_442);
not ( n20547 , RI15b4b810_441);
nor ( n20548 , n20546 , n20547 );
nand ( n20549 , n20545 , n20548 );
nand ( n20550 , RI15b4b900_443 , RI15b4b978_444);
nor ( n20551 , n20549 , n20550 );
and ( n20552 , n20551 , RI15b4b9f0_445);
nand ( n20553 , n20552 , RI15b4ba68_446);
nand ( n20554 , RI15b4bae0_447 , RI15b4bb58_448);
nor ( n20555 , n20553 , n20554 );
and ( n20556 , n20555 , RI15b4bbd0_449 , RI15b4bc48_450);
and ( n20557 , n20556 , RI15b4bcc0_451 , RI15b4bd38_452);
and ( n20558 , n20557 , RI15b4bdb0_453 , RI15b4be28_454);
nand ( n20559 , n20558 , RI15b4bea0_455 , RI15b4bf18_456);
not ( n20560 , n20489 );
nor ( n20561 , n20560 , n20516 );
nand ( n20562 , n20561 , n20510 , n19913 );
nand ( n20563 , n20416 , n20511 , n20493 );
and ( n20564 , n20562 , n20563 );
not ( n20565 , n20564 );
and ( n20566 , n20565 , n20501 );
not ( n20567 , n20566 );
not ( n20568 , n20567 );
and ( n20569 , n20559 , n20568 );
not ( n20570 , n20416 );
not ( n20571 , n20292 );
and ( n20572 , n20375 , n20571 , n20412 );
not ( n20573 , n20208 );
and ( n20574 , n20573 , n20167 , n20116 );
nand ( n20575 , n20572 , n20574 );
not ( n20576 , n20251 );
nand ( n20577 , n20507 , n20576 );
nor ( n20578 , n20575 , n20577 );
not ( n20579 , n20578 );
nand ( n20580 , n20570 , n20579 );
buf ( n20581 , n20572 );
and ( n20582 , n20332 , n20576 );
buf ( n20583 , n20582 );
nand ( n20584 , n20581 , n20583 , n20574 );
nand ( n20585 , n20509 , n20584 );
nor ( n20586 , n20580 , n20585 );
nand ( n20587 , n20375 , n20412 );
nor ( n20588 , n20294 , n20587 );
and ( n20589 , n20588 , n20332 );
nand ( n20590 , n20376 , n20573 , n20412 );
buf ( n20591 , n20167 );
nand ( n20592 , n20117 , n20591 );
nor ( n20593 , n20590 , n20592 );
not ( n20594 , n20577 );
nand ( n20595 , n20593 , n20594 );
nand ( n20596 , n20507 , n20251 );
not ( n20597 , n20596 );
not ( n20598 , n20209 );
nand ( n20599 , n20597 , n20581 , n20598 );
nand ( n20600 , n20595 , n20599 );
nor ( n20601 , n20589 , n20600 );
not ( n20602 , n20582 );
nand ( n20603 , n20602 , n20596 );
and ( n20604 , n20375 , n20413 , n20292 );
nand ( n20605 , n20598 , n20604 );
nor ( n20606 , n20603 , n20605 );
not ( n20607 , n20606 );
and ( n20608 , n20586 , n20601 , n20607 );
not ( n20609 , n20608 );
not ( n20610 , n20512 );
nor ( n20611 , n20606 , n20610 );
nand ( n20612 , n20609 , n20601 , n20611 );
nand ( n20613 , n20612 , n20501 );
not ( n20614 , RI15b44da8_214);
nand ( n20615 , n19908 , n20614 );
not ( n20616 , n20615 );
not ( n20617 , RI15b44e20_215);
and ( n20618 , n20616 , n20617 );
and ( n20619 , n20615 , RI15b44e20_215);
nor ( n20620 , n20618 , n20619 );
or ( n20621 , n20620 , n20499 );
nand ( n20622 , n20499 , RI15b44e20_215);
or ( n20623 , n20615 , n20622 );
not ( n20624 , n20498 );
nand ( n20625 , RI15b44cb8_212 , RI15b44d30_213);
nor ( n20626 , n20624 , n20625 );
not ( n20627 , n20626 );
and ( n20628 , n20623 , n20627 );
not ( n20629 , n19909 );
or ( n20630 , n20624 , n20629 );
not ( n20631 , n20630 );
not ( n20632 , n20625 );
nand ( n20633 , n20632 , n19910 );
not ( n20634 , n20633 );
nor ( n20635 , n20624 , RI15b44cb8_212 , RI15b44d30_213);
nor ( n20636 , n20631 , n20634 , n20635 );
and ( n20637 , n19912 , RI15b47df0_317);
not ( n20638 , n20637 );
and ( n20639 , n20621 , n20628 , n20636 , n20638 );
and ( n20640 , n20613 , n20639 );
not ( n20641 , n20640 );
nor ( n20642 , n20569 , n20641 );
not ( n20643 , RI15b4bf90_457);
or ( n20644 , n20642 , n20643 );
not ( n20645 , n20559 );
buf ( n20646 , n20566 );
buf ( n20647 , n20646 );
and ( n20648 , n20645 , n20647 , n20643 );
not ( n20649 , n20615 );
nand ( n20650 , n20649 , RI15b44cb8_212 , RI15b44e20_215);
buf ( n20651 , n20650 );
not ( n20652 , n20651 );
not ( n20653 , n20652 );
not ( n20654 , n20653 );
buf ( n20655 , n20654 );
buf ( n20656 , n20655 );
and ( n20657 , n20656 , RI15b4b090_425);
nor ( n20658 , n20648 , n20657 );
nand ( n20659 , n20644 , n20658 );
nor ( n20660 , n20531 , n20659 );
nand ( n20661 , n19952 , n20523 , n20527 , n20660 );
buf ( n20662 , n20661 );
buf ( n20663 , RI15b3ea48_2);
buf ( n20664 , n20663 );
buf ( n20665 , RI15b3e9d0_1);
buf ( n20666 , n20665 );
nand ( n20667 , RI15b4ffc8_594 , RI15b50040_595);
nand ( n20668 , RI15b500b8_596 , RI15b50130_597);
nor ( n20669 , n20667 , n20668 );
and ( n20670 , RI15b501a8_598 , RI15b50220_599);
nand ( n20671 , n20669 , n20670 );
not ( n20672 , RI15b50298_600);
nor ( n20673 , n20671 , n20672 );
nand ( n20674 , n20673 , RI15b50310_601);
not ( n20675 , RI15b50388_602);
nor ( n20676 , n20674 , n20675 );
nand ( n20677 , n20676 , RI15b50400_603);
not ( n20678 , RI15b50478_604);
nor ( n20679 , n20677 , n20678 );
not ( n20680 , n20679 );
nand ( n20681 , RI15b504f0_605 , RI15b50568_606);
not ( n20682 , RI15b505e0_607);
nor ( n20683 , n20681 , n20682 );
nand ( n20684 , n20683 , RI15b50658_608);
not ( n20685 , RI15b506d0_609);
nor ( n20686 , n20684 , n20685 );
nand ( n20687 , n20686 , RI15b50748_610);
not ( n20688 , n20687 );
nand ( n20689 , n20688 , RI15b507c0_611);
nor ( n20690 , n20680 , n20689 );
and ( n20691 , n20690 , RI15b50838_612);
not ( n20692 , n20691 );
and ( n20693 , RI15b508b0_613 , n20692 );
not ( n20694 , RI15b508b0_613);
and ( n20695 , n20694 , n20691 );
nor ( n20696 , n20693 , n20695 );
not ( n20697 , n20696 );
buf ( n20698 , n20680 );
buf ( n20699 , n20698 );
and ( n20700 , n20699 , RI15b50748_610);
buf ( n20701 , n20698 );
not ( n20702 , RI15b50748_610);
nand ( n20703 , n20686 , n20702 );
or ( n20704 , n20701 , n20703 );
not ( n20705 , n20686 );
nand ( n20706 , n20705 , RI15b50748_610);
nand ( n20707 , n20704 , n20706 );
nor ( n20708 , n20700 , n20707 );
not ( n20709 , n20708 );
buf ( n20710 , n20699 );
and ( n20711 , n20710 , RI15b50658_608);
not ( n20712 , RI15b50658_608);
nand ( n20713 , n20683 , n20712 );
or ( n20714 , n20710 , n20713 );
not ( n20715 , n20683 );
nand ( n20716 , n20715 , RI15b50658_608);
nand ( n20717 , n20714 , n20716 );
nor ( n20718 , n20711 , n20717 );
not ( n20719 , n20718 );
buf ( n20720 , n18211 );
not ( n20721 , n20720 );
not ( n20722 , n17621 );
not ( n20723 , RI15b50f40_627);
and ( n20724 , n20722 , n20723 );
and ( n20725 , n17621 , RI15b50f40_627);
nor ( n20726 , n20724 , n20725 );
not ( n20727 , n20726 );
not ( n20728 , RI15b50e50_625);
nand ( n20729 , n20728 , RI15b50ec8_626);
nand ( n20730 , n20729 , n17632 );
not ( n20731 , RI15b50e50_625);
and ( n20732 , n20730 , n20731 );
nand ( n20733 , n20727 , n20732 );
not ( n20734 , n20733 );
nand ( n20735 , n20721 , n20734 );
not ( n20736 , n20735 );
not ( n20737 , RI15b4e0d8_528);
not ( n20738 , n20737 );
and ( n20739 , n20736 , n20738 );
not ( n20740 , n18213 );
nor ( n20741 , n20730 , RI15b50e50_625);
not ( n20742 , n20741 );
nor ( n20743 , n20742 , n20726 );
nand ( n20744 , n20740 , n20743 );
not ( n20745 , n20744 );
not ( n20746 , n20745 );
nor ( n20747 , n20746 , n17758 );
nor ( n20748 , n20739 , n20747 );
not ( n20749 , n20720 );
not ( n20750 , n20726 );
nand ( n20751 , n20730 , RI15b50e50_625);
not ( n20752 , n20751 );
nand ( n20753 , n20750 , n20752 );
not ( n20754 , n20753 );
nand ( n20755 , n20749 , n20754 );
not ( n20756 , n20755 );
not ( n20757 , n17741 );
and ( n20758 , n20756 , n20757 );
not ( n20759 , n20752 );
not ( n20760 , n20726 );
nor ( n20761 , n20759 , n20760 );
nand ( n20762 , n20761 , n20720 );
buf ( n20763 , n20762 );
not ( n20764 , n20763 );
and ( n20765 , n20764 , RI15b4ec18_552);
nor ( n20766 , n20758 , n20765 );
not ( n20767 , n17615 );
and ( n20768 , n18212 , n20767 );
not ( n20769 , n20768 );
not ( n20770 , n20769 );
not ( n20771 , RI15b4d598_504);
not ( n20772 , n20771 );
and ( n20773 , n20770 , n20772 );
not ( n20774 , n18212 );
not ( n20775 , n18206 );
nand ( n20776 , n20774 , n20775 );
buf ( n20777 , n20776 );
not ( n20778 , n20777 );
and ( n20779 , n20778 , RI15b4e498_536);
nor ( n20780 , n20773 , n20779 );
not ( n20781 , n18212 );
not ( n20782 , n20732 );
nor ( n20783 , n20782 , n20760 );
nand ( n20784 , n20781 , n20783 );
not ( n20785 , n20784 );
not ( n20786 , RI15b4efd8_560);
not ( n20787 , n20786 );
and ( n20788 , n20785 , n20787 );
not ( n20789 , n18212 );
and ( n20790 , n20741 , n20726 );
nand ( n20791 , n20789 , n20790 );
not ( n20792 , RI15b4e858_544);
nor ( n20793 , n20791 , n20792 );
nor ( n20794 , n20788 , n20793 );
nand ( n20795 , n20748 , n20766 , n20780 , n20794 );
not ( n20796 , n18212 );
nand ( n20797 , n20796 , n20734 );
not ( n20798 , n20797 );
not ( n20799 , RI15b4fed8_592);
not ( n20800 , n20799 );
and ( n20801 , n20798 , n20800 );
not ( n20802 , n18212 );
nand ( n20803 , n20802 , n20743 );
not ( n20804 , n20803 );
not ( n20805 , n20804 );
not ( n20806 , RI15b4f758_576);
nor ( n20807 , n20805 , n20806 );
nor ( n20808 , n20801 , n20807 );
nand ( n20809 , n20796 , n20754 );
not ( n20810 , n20809 );
not ( n20811 , RI15b4fb18_584);
not ( n20812 , n20811 );
and ( n20813 , n20810 , n20812 );
not ( n20814 , n20720 );
nor ( n20815 , n20751 , n20760 );
nand ( n20816 , n20814 , n20815 );
not ( n20817 , n20816 );
and ( n20818 , n20817 , RI15b4ce18_488);
nor ( n20819 , n20813 , n20818 );
not ( n20820 , n20720 );
nand ( n20821 , n20820 , n20775 );
buf ( n20822 , n20821 );
not ( n20823 , n20822 );
not ( n20824 , n17765 );
and ( n20825 , n20823 , n20824 );
nand ( n20826 , n20720 , n20767 );
buf ( n20827 , n20826 );
not ( n20828 , n20827 );
and ( n20829 , n20828 , RI15b4f398_568);
nor ( n20830 , n20825 , n20829 );
not ( n20831 , n20726 );
nor ( n20832 , n20782 , n20831 );
not ( n20833 , n20720 );
nand ( n20834 , n20832 , n20833 );
buf ( n20835 , n20834 );
not ( n20836 , n20835 );
not ( n20837 , RI15b4d1d8_496);
not ( n20838 , n20837 );
and ( n20839 , n20836 , n20838 );
not ( n20840 , n20720 );
nand ( n20841 , n20840 , n20790 );
buf ( n20842 , n20841 );
nor ( n20843 , n20842 , n17755 );
nor ( n20844 , n20839 , n20843 );
nand ( n20845 , n20808 , n20819 , n20830 , n20844 );
nor ( n20846 , n20795 , n20845 );
buf ( n20847 , n20846 );
buf ( n20848 , n20847 );
buf ( n20849 , n20848 );
not ( n20850 , n20849 );
not ( n20851 , n20735 );
not ( n20852 , RI15b4e060_527);
not ( n20853 , n20852 );
and ( n20854 , n20851 , n20853 );
not ( n20855 , n20744 );
not ( n20856 , n20855 );
nor ( n20857 , n20856 , n17900 );
nor ( n20858 , n20854 , n20857 );
not ( n20859 , RI15b4cda0_487);
nor ( n20860 , n20816 , n20859 );
nor ( n20861 , n20755 , n17883 );
nor ( n20862 , n20860 , n20861 );
not ( n20863 , n20835 );
not ( n20864 , RI15b4d160_495);
not ( n20865 , n20864 );
and ( n20866 , n20863 , n20865 );
nor ( n20867 , n20842 , n17897 );
nor ( n20868 , n20866 , n20867 );
not ( n20869 , n20768 );
not ( n20870 , RI15b4d520_503);
nor ( n20871 , n20869 , n20870 );
nor ( n20872 , n20822 , n17904 );
nor ( n20873 , n20871 , n20872 );
nand ( n20874 , n20858 , n20862 , n20868 , n20873 );
not ( n20875 , n20797 );
not ( n20876 , RI15b4fe60_591);
not ( n20877 , n20876 );
and ( n20878 , n20875 , n20877 );
not ( n20879 , n20803 );
not ( n20880 , n20879 );
not ( n20881 , RI15b4f6e0_575);
nor ( n20882 , n20880 , n20881 );
nor ( n20883 , n20878 , n20882 );
not ( n20884 , n20763 );
not ( n20885 , RI15b4eba0_551);
not ( n20886 , n20885 );
and ( n20887 , n20884 , n20886 );
not ( n20888 , RI15b4faa0_583);
nor ( n20889 , n20809 , n20888 );
nor ( n20890 , n20887 , n20889 );
not ( n20891 , n20827 );
not ( n20892 , RI15b4f320_567);
not ( n20893 , n20892 );
and ( n20894 , n20891 , n20893 );
not ( n20895 , RI15b4e420_535);
nor ( n20896 , n20777 , n20895 );
nor ( n20897 , n20894 , n20896 );
not ( n20898 , n20784 );
not ( n20899 , RI15b4ef60_559);
not ( n20900 , n20899 );
and ( n20901 , n20898 , n20900 );
not ( n20902 , RI15b4e7e0_543);
nor ( n20903 , n20791 , n20902 );
nor ( n20904 , n20901 , n20903 );
nand ( n20905 , n20883 , n20890 , n20897 , n20904 );
nor ( n20906 , n20874 , n20905 );
not ( n20907 , n20906 );
buf ( n20908 , n20907 );
not ( n20909 , n20908 );
buf ( n20910 , n20669 );
not ( n20911 , RI15b50220_599);
or ( n20912 , n20910 , n20911 );
buf ( n20913 , n20910 );
and ( n20914 , n20911 , RI15b501a8_598);
and ( n20915 , n20913 , n20914 );
not ( n20916 , RI15b501a8_598);
and ( n20917 , n20916 , RI15b50220_599);
nor ( n20918 , n20915 , n20917 );
nand ( n20919 , n20912 , n20918 );
not ( n20920 , n20919 );
nand ( n20921 , n20909 , n20920 );
not ( n20922 , n20921 );
and ( n20923 , n20913 , RI15b501a8_598);
not ( n20924 , n20913 );
and ( n20925 , n20924 , n20916 );
nor ( n20926 , n20923 , n20925 );
not ( n20927 , n20926 );
not ( n20928 , n20809 );
nand ( n20929 , n20928 , RI15b4fa28_582);
nand ( n20930 , n20764 , RI15b4eb28_550);
not ( n20931 , n20797 );
nand ( n20932 , n20931 , RI15b4fde8_590);
not ( n20933 , n20880 );
nand ( n20934 , n20933 , RI15b4f668_574);
nand ( n20935 , n20929 , n20930 , n20932 , n20934 );
not ( n20936 , n20784 );
nand ( n20937 , n20936 , RI15b4eee8_558);
not ( n20938 , n20791 );
nand ( n20939 , n20938 , RI15b4e768_542);
nand ( n20940 , n20778 , RI15b4e3a8_534);
nand ( n20941 , n20828 , RI15b4f2a8_566);
nand ( n20942 , n20937 , n20939 , n20940 , n20941 );
nor ( n20943 , n20935 , n20942 );
not ( n20944 , n20755 );
nand ( n20945 , n20944 , RI15b4dc28_518);
nand ( n20946 , n20817 , RI15b4cd28_486);
not ( n20947 , n20835 );
nand ( n20948 , n20947 , RI15b4d0e8_494);
not ( n20949 , n20842 );
nand ( n20950 , n20949 , RI15b4c968_478);
nand ( n20951 , n20945 , n20946 , n20948 , n20950 );
not ( n20952 , n20735 );
nand ( n20953 , n20952 , RI15b4dfe8_526);
nand ( n20954 , n20745 , RI15b4d868_510);
not ( n20955 , n20822 );
nand ( n20956 , n20955 , RI15b4c5a8_470);
not ( n20957 , n20869 );
nand ( n20958 , n20957 , RI15b4d4a8_502);
nand ( n20959 , n20953 , n20954 , n20956 , n20958 );
nor ( n20960 , n20951 , n20959 );
nand ( n20961 , n20943 , n20960 );
not ( n20962 , n20961 );
nand ( n20963 , n20927 , n20962 );
not ( n20964 , n20963 );
not ( n20965 , n20735 );
not ( n20966 , RI15b4def8_524);
not ( n20967 , n20966 );
and ( n20968 , n20965 , n20967 );
nor ( n20969 , n20842 , n17716 );
nor ( n20970 , n20968 , n20969 );
not ( n20971 , RI15b4cc38_484);
nor ( n20972 , n20816 , n20971 );
nor ( n20973 , n20755 , n17702 );
nor ( n20974 , n20972 , n20973 );
not ( n20975 , n20835 );
not ( n20976 , RI15b4cff8_492);
not ( n20977 , n20976 );
and ( n20978 , n20975 , n20977 );
not ( n20979 , RI15b4d778_508);
nor ( n20980 , n20744 , n20979 );
nor ( n20981 , n20978 , n20980 );
not ( n20982 , RI15b4d3b8_500);
nor ( n20983 , n20769 , n20982 );
not ( n20984 , n20821 );
not ( n20985 , n20984 );
nor ( n20986 , n20985 , n17723 );
nor ( n20987 , n20983 , n20986 );
nand ( n20988 , n20970 , n20974 , n20981 , n20987 );
not ( n20989 , n20784 );
not ( n20990 , RI15b4edf8_556);
not ( n20991 , n20990 );
and ( n20992 , n20989 , n20991 );
not ( n20993 , RI15b4ea38_548);
nor ( n20994 , n20763 , n20993 );
nor ( n20995 , n20992 , n20994 );
not ( n20996 , n20797 );
not ( n20997 , RI15b4fcf8_588);
not ( n20998 , n20997 );
and ( n20999 , n20996 , n20998 );
not ( n21000 , RI15b4f578_572);
nor ( n21001 , n20803 , n21000 );
nor ( n21002 , n20999 , n21001 );
not ( n21003 , n20827 );
not ( n21004 , RI15b4f1b8_564);
not ( n21005 , n21004 );
and ( n21006 , n21003 , n21005 );
not ( n21007 , RI15b4e2b8_532);
nor ( n21008 , n20777 , n21007 );
nor ( n21009 , n21006 , n21008 );
not ( n21010 , n20809 );
not ( n21011 , n17729 );
and ( n21012 , n21010 , n21011 );
not ( n21013 , RI15b4e678_540);
nor ( n21014 , n20791 , n21013 );
nor ( n21015 , n21012 , n21014 );
nand ( n21016 , n20995 , n21002 , n21009 , n21015 );
nor ( n21017 , n20988 , n21016 );
and ( n21018 , n20667 , RI15b500b8_596);
not ( n21019 , n20667 );
not ( n21020 , RI15b500b8_596);
and ( n21021 , n21019 , n21020 );
nor ( n21022 , n21018 , n21021 );
nand ( n21023 , n21017 , n21022 );
not ( n21024 , n20816 );
not ( n21025 , n17862 );
and ( n21026 , n21024 , n21025 );
and ( n21027 , n20931 , RI15b4fd70_589);
nor ( n21028 , n21026 , n21027 );
and ( n21029 , n20804 , RI15b4f5f0_573);
and ( n21030 , n20928 , RI15b4f9b0_581);
nor ( n21031 , n21029 , n21030 );
nand ( n21032 , n21028 , n21031 );
not ( n21033 , n20835 );
nand ( n21034 , n21033 , RI15b4d070_493);
not ( n21035 , n20842 );
nand ( n21036 , n21035 , RI15b4c8f0_477);
not ( n21037 , n20827 );
nand ( n21038 , n21037 , RI15b4f230_565);
nand ( n21039 , n20984 , RI15b4c530_469);
nand ( n21040 , n21034 , n21036 , n21038 , n21039 );
nor ( n21041 , n21032 , n21040 );
nand ( n21042 , n20944 , RI15b4dbb0_517);
not ( n21043 , n20763 );
nand ( n21044 , n21043 , RI15b4eab0_549);
nand ( n21045 , n20936 , RI15b4ee70_557);
nand ( n21046 , n20938 , RI15b4e6f0_541);
nand ( n21047 , n21042 , n21044 , n21045 , n21046 );
nand ( n21048 , n20952 , RI15b4df70_525);
nand ( n21049 , n20745 , RI15b4d7f0_509);
not ( n21050 , n20777 );
nand ( n21051 , n21050 , RI15b4e330_533);
nand ( n21052 , n20768 , RI15b4d430_501);
nand ( n21053 , n21048 , n21049 , n21051 , n21052 );
nor ( n21054 , n21047 , n21053 );
nand ( n21055 , n21041 , n21054 );
not ( n21056 , n21055 );
and ( n21057 , n20667 , RI15b50130_597);
nor ( n21058 , n21020 , RI15b50130_597);
not ( n21059 , n21058 );
or ( n21060 , n21059 , n20667 );
nand ( n21061 , n21020 , RI15b50130_597);
nand ( n21062 , n21060 , n21061 );
nor ( n21063 , n21057 , n21062 );
nand ( n21064 , n21056 , n21063 );
nand ( n21065 , n21023 , n21064 );
nand ( n21066 , n20952 , RI15b4de80_523);
nand ( n21067 , n20947 , RI15b4cf80_491);
not ( n21068 , n20822 );
nand ( n21069 , n21068 , RI15b4c440_467);
not ( n21070 , n20769 );
nand ( n21071 , n21070 , RI15b4d340_499);
nand ( n21072 , n21066 , n21067 , n21069 , n21071 );
nand ( n21073 , n20944 , RI15b4dac0_515);
nand ( n21074 , n20817 , RI15b4cbc0_483);
nand ( n21075 , n20855 , RI15b4d700_507);
nand ( n21076 , n20949 , RI15b4c800_475);
nand ( n21077 , n21073 , n21074 , n21075 , n21076 );
nor ( n21078 , n21072 , n21077 );
nand ( n21079 , n20928 , RI15b4f8c0_579);
nand ( n21080 , n20764 , RI15b4e9c0_547);
nand ( n21081 , n20933 , RI15b4f500_571);
nand ( n21082 , n20936 , RI15b4ed80_555);
nand ( n21083 , n21079 , n21080 , n21081 , n21082 );
nand ( n21084 , n20931 , RI15b4fc80_587);
nand ( n21085 , n20938 , RI15b4e600_539);
nand ( n21086 , n20778 , RI15b4e240_531);
nand ( n21087 , n20828 , RI15b4f140_563);
nand ( n21088 , n21084 , n21085 , n21086 , n21087 );
nor ( n21089 , n21083 , n21088 );
nand ( n21090 , n21078 , n21089 );
not ( n21091 , RI15b50040_595);
not ( n21092 , n21091 );
not ( n21093 , RI15b4ffc8_594);
not ( n21094 , n21093 );
or ( n21095 , n21092 , n21094 );
nand ( n21096 , n21095 , n20667 );
not ( n21097 , n21096 );
nor ( n21098 , n21090 , n21097 );
nor ( n21099 , n21065 , n21098 );
not ( n21100 , n21099 );
not ( n21101 , n20735 );
not ( n21102 , RI15b4de08_522);
not ( n21103 , n21102 );
and ( n21104 , n21101 , n21103 );
and ( n21105 , n20936 , RI15b4ed08_554);
nor ( n21106 , n21104 , n21105 );
not ( n21107 , n20821 );
not ( n21108 , RI15b4c3c8_466);
not ( n21109 , n21108 );
and ( n21110 , n21107 , n21109 );
not ( n21111 , RI15b4c788_474);
nor ( n21112 , n20841 , n21111 );
nor ( n21113 , n21110 , n21112 );
not ( n21114 , n20768 );
not ( n21115 , n21114 );
not ( n21116 , RI15b4d2c8_498);
not ( n21117 , n21116 );
and ( n21118 , n21115 , n21117 );
not ( n21119 , n20826 );
not ( n21120 , n21119 );
not ( n21121 , RI15b4f0c8_562);
nor ( n21122 , n21120 , n21121 );
nor ( n21123 , n21118 , n21122 );
not ( n21124 , n20791 );
not ( n21125 , RI15b4e588_538);
not ( n21126 , n21125 );
and ( n21127 , n21124 , n21126 );
not ( n21128 , n20776 );
not ( n21129 , n21128 );
not ( n21130 , RI15b4e1c8_530);
nor ( n21131 , n21129 , n21130 );
nor ( n21132 , n21127 , n21131 );
nand ( n21133 , n21106 , n21113 , n21123 , n21132 );
not ( n21134 , n20835 );
not ( n21135 , RI15b4cf08_490);
not ( n21136 , n21135 );
and ( n21137 , n21134 , n21136 );
not ( n21138 , n20763 );
and ( n21139 , n21138 , RI15b4e948_546);
nor ( n21140 , n21137 , n21139 );
not ( n21141 , n20797 );
not ( n21142 , RI15b4fc08_586);
not ( n21143 , n21142 );
and ( n21144 , n21141 , n21143 );
and ( n21145 , n20855 , RI15b4d688_506);
nor ( n21146 , n21144 , n21145 );
not ( n21147 , n20816 );
not ( n21148 , RI15b4cb48_482);
not ( n21149 , n21148 );
and ( n21150 , n21147 , n21149 );
not ( n21151 , RI15b4da48_514);
nor ( n21152 , n20755 , n21151 );
nor ( n21153 , n21150 , n21152 );
not ( n21154 , n20809 );
not ( n21155 , RI15b4f848_578);
not ( n21156 , n21155 );
and ( n21157 , n21154 , n21156 );
not ( n21158 , RI15b4f488_570);
nor ( n21159 , n20803 , n21158 );
nor ( n21160 , n21157 , n21159 );
nand ( n21161 , n21140 , n21146 , n21153 , n21160 );
nor ( n21162 , n21133 , n21161 );
not ( n21163 , n21162 );
not ( n21164 , RI15b4dd90_521);
nor ( n21165 , n20735 , n21164 );
nor ( n21166 , n20755 , n17957 );
nor ( n21167 , n21165 , n21166 );
and ( n21168 , n20817 , RI15b4cad0_481);
and ( n21169 , n20984 , RI15b4c350_465);
nor ( n21170 , n21168 , n21169 );
nand ( n21171 , n21167 , n21170 );
not ( n21172 , RI15b4ce90_489);
nor ( n21173 , n20834 , n21172 );
nor ( n21174 , n20841 , n17971 );
nor ( n21175 , n21173 , n21174 );
not ( n21176 , RI15b4fb90_585);
nor ( n21177 , n20797 , n21176 );
nor ( n21178 , n20809 , n17984 );
nor ( n21179 , n21177 , n21178 );
nand ( n21180 , n21175 , n21179 );
nor ( n21181 , n21171 , n21180 );
not ( n21182 , RI15b4e8d0_545);
nor ( n21183 , n20762 , n21182 );
not ( n21184 , RI15b4e510_537);
nor ( n21185 , n20791 , n21184 );
nor ( n21186 , n21183 , n21185 );
and ( n21187 , n20936 , RI15b4ec90_553);
and ( n21188 , n20879 , RI15b4f410_569);
nor ( n21189 , n21187 , n21188 );
nand ( n21190 , n21186 , n21189 );
not ( n21191 , n20744 );
nand ( n21192 , n21191 , RI15b4d610_505);
nand ( n21193 , n21119 , RI15b4f050_561);
nand ( n21194 , n20768 , RI15b4d250_497);
nand ( n21195 , n21128 , RI15b4e150_529);
nand ( n21196 , n21192 , n21193 , n21194 , n21195 );
nor ( n21197 , n21190 , n21196 );
nand ( n21198 , n21181 , n21197 );
nand ( n21199 , n21198 , RI15b4ff50_593);
not ( n21200 , n21199 );
or ( n21201 , n21163 , n21200 );
nand ( n21202 , n21201 , n21093 );
not ( n21203 , n21199 );
not ( n21204 , n21162 );
nand ( n21205 , n21203 , n21204 );
nand ( n21206 , n21202 , n21205 );
not ( n21207 , n21206 );
or ( n21208 , n21100 , n21207 );
not ( n21209 , n21065 );
not ( n21210 , n21090 );
nor ( n21211 , n21210 , n21096 );
and ( n21212 , n21209 , n21211 );
not ( n21213 , n21064 );
nor ( n21214 , n21017 , n21022 );
not ( n21215 , n21214 );
or ( n21216 , n21213 , n21215 );
not ( n21217 , n21055 );
not ( n21218 , n21217 );
not ( n21219 , n21063 );
nand ( n21220 , n21218 , n21219 );
nand ( n21221 , n21216 , n21220 );
nor ( n21222 , n21212 , n21221 );
nand ( n21223 , n21208 , n21222 );
not ( n21224 , n21223 );
or ( n21225 , n20964 , n21224 );
not ( n21226 , n20962 );
nand ( n21227 , n21226 , n20926 );
nand ( n21228 , n21225 , n21227 );
not ( n21229 , n21228 );
or ( n21230 , n20922 , n21229 );
nand ( n21231 , n20908 , n20919 );
nand ( n21232 , n21230 , n21231 );
not ( n21233 , n20671 );
and ( n21234 , n21233 , RI15b50298_600);
not ( n21235 , n21233 );
and ( n21236 , n21235 , n20672 );
nor ( n21237 , n21234 , n21236 );
nand ( n21238 , n21232 , n21237 );
not ( n21239 , n21238 );
or ( n21240 , n20850 , n21239 );
not ( n21241 , n21232 );
not ( n21242 , n21237 );
and ( n21243 , n21241 , n21242 );
not ( n21244 , RI15b50388_602);
not ( n21245 , n20674 );
or ( n21246 , n21244 , n21245 );
or ( n21247 , n20674 , RI15b50388_602);
nand ( n21248 , n21246 , n21247 );
not ( n21249 , n20673 );
not ( n21250 , RI15b50310_601);
and ( n21251 , n21249 , n21250 );
not ( n21252 , n21249 );
and ( n21253 , n21252 , RI15b50310_601);
nor ( n21254 , n21251 , n21253 );
nand ( n21255 , n21248 , n21254 );
nor ( n21256 , n21243 , n21255 );
nand ( n21257 , n21240 , n21256 );
and ( n21258 , n20698 , RI15b505e0_607);
nor ( n21259 , n20681 , RI15b505e0_607);
not ( n21260 , n21259 );
or ( n21261 , n20698 , n21260 );
nand ( n21262 , n20681 , RI15b505e0_607);
nand ( n21263 , n21261 , n21262 );
nor ( n21264 , n21258 , n21263 );
not ( n21265 , n21264 );
and ( n21266 , n20698 , RI15b504f0_605);
not ( n21267 , n20698 );
not ( n21268 , RI15b504f0_605);
and ( n21269 , n21267 , n21268 );
nor ( n21270 , n21266 , n21269 );
not ( n21271 , n20677 );
not ( n21272 , n21271 );
and ( n21273 , n21272 , RI15b50478_604);
not ( n21274 , n21272 );
and ( n21275 , n21274 , n20678 );
nor ( n21276 , n21273 , n21275 );
not ( n21277 , n20676 );
and ( n21278 , n21277 , RI15b50400_603);
not ( n21279 , n21277 );
not ( n21280 , RI15b50400_603);
and ( n21281 , n21279 , n21280 );
nor ( n21282 , n21278 , n21281 );
nor ( n21283 , n21270 , n21276 , n21282 );
and ( n21284 , n20701 , RI15b50568_606);
not ( n21285 , RI15b50568_606);
nand ( n21286 , n21285 , RI15b504f0_605);
or ( n21287 , n20698 , n21286 );
nand ( n21288 , n21268 , RI15b50568_606);
nand ( n21289 , n21287 , n21288 );
nor ( n21290 , n21284 , n21289 );
not ( n21291 , n21290 );
nand ( n21292 , n21265 , n21283 , n21291 );
nor ( n21293 , n21257 , n21292 );
nand ( n21294 , n20719 , n21293 );
and ( n21295 , n20710 , RI15b506d0_609);
nor ( n21296 , n20684 , RI15b506d0_609);
not ( n21297 , n21296 );
or ( n21298 , n20710 , n21297 );
nand ( n21299 , n20684 , RI15b506d0_609);
nand ( n21300 , n21298 , n21299 );
nor ( n21301 , n21295 , n21300 );
nor ( n21302 , n21294 , n21301 );
buf ( n21303 , n21302 );
nand ( n21304 , n20709 , n21303 );
and ( n21305 , n20701 , RI15b507c0_611);
nor ( n21306 , n20687 , RI15b507c0_611);
not ( n21307 , n21306 );
or ( n21308 , n20701 , n21307 );
nand ( n21309 , n20687 , RI15b507c0_611);
nand ( n21310 , n21308 , n21309 );
nor ( n21311 , n21305 , n21310 );
nor ( n21312 , n21304 , n21311 );
not ( n21313 , n20690 );
not ( n21314 , RI15b50838_612);
and ( n21315 , n21313 , n21314 );
not ( n21316 , n21313 );
and ( n21317 , n21316 , RI15b50838_612);
nor ( n21318 , n21315 , n21317 );
and ( n21319 , n21312 , n21318 );
nand ( n21320 , n20697 , n21319 );
and ( n21321 , n20692 , RI15b50928_614);
not ( n21322 , RI15b508b0_613);
nor ( n21323 , n21322 , RI15b50928_614);
not ( n21324 , n21323 );
not ( n21325 , n20691 );
or ( n21326 , n21324 , n21325 );
nand ( n21327 , n21322 , RI15b50928_614);
nand ( n21328 , n21326 , n21327 );
nor ( n21329 , n21321 , n21328 );
and ( n21330 , n21320 , n21329 );
not ( n21331 , n21320 );
not ( n21332 , n21329 );
and ( n21333 , n21331 , n21332 );
nor ( n21334 , n21330 , n21333 );
nor ( n21335 , n18130 , n18078 );
not ( n21336 , n18056 );
and ( n21337 , n18057 , RI15b4c170_461);
and ( n21338 , n21337 , n17622 );
or ( n21339 , n18003 , n18062 );
or ( n21340 , n20729 , RI15b4c170_461);
nand ( n21341 , n21339 , n21340 );
and ( n21342 , n21341 , RI15b4c0f8_460);
not ( n21343 , n17633 );
buf ( n21344 , n18001 );
and ( n21345 , n21343 , n21344 );
nor ( n21346 , n21338 , n21342 , n21345 );
nor ( n21347 , n18049 , n21346 );
nor ( n21348 , n21336 , n21347 );
and ( n21349 , n18051 , n21348 );
not ( n21350 , n21349 );
nand ( n21351 , n21335 , n21350 );
not ( n21352 , n20849 );
nor ( n21353 , n21351 , n21352 );
buf ( n21354 , n21353 );
buf ( n21355 , n21354 );
buf ( n21356 , n21355 );
buf ( n21357 , n21356 );
not ( n21358 , n21357 );
buf ( n21359 , n21358 );
not ( n21360 , n21359 );
buf ( n21361 , n21360 );
buf ( n21362 , n21361 );
and ( n21363 , n21334 , n21362 );
nand ( n21364 , RI15b4ff50_593 , RI15b4ffc8_594);
nand ( n21365 , n21364 , n21091 );
not ( n21366 , n20668 );
nand ( n21367 , n21365 , n21366 );
not ( n21368 , n20670 );
nor ( n21369 , n21367 , n21368 );
nand ( n21370 , n21369 , RI15b50298_600);
nor ( n21371 , n21370 , n21250 );
nand ( n21372 , n21371 , RI15b50388_602);
nor ( n21373 , n21372 , n21280 );
and ( n21374 , n21373 , RI15b50478_604);
not ( n21375 , n20689 );
and ( n21376 , n21374 , n21375 );
and ( n21377 , n21376 , RI15b50838_612);
not ( n21378 , n21377 );
and ( n21379 , RI15b508b0_613 , n21378 );
not ( n21380 , RI15b508b0_613);
and ( n21381 , n21380 , n21377 );
nor ( n21382 , n21379 , n21381 );
not ( n21383 , n21382 );
and ( n21384 , n21365 , n21020 );
not ( n21385 , n21365 );
and ( n21386 , n21385 , RI15b500b8_596);
nor ( n21387 , n21384 , n21386 );
not ( n21388 , n21387 );
buf ( n21389 , n21017 );
not ( n21390 , n21389 );
not ( n21391 , n21390 );
not ( n21392 , n21391 );
or ( n21393 , n21388 , n21392 );
and ( n21394 , n21364 , RI15b50040_595);
not ( n21395 , n21364 );
and ( n21396 , n21395 , n21091 );
nor ( n21397 , n21394 , n21396 );
not ( n21398 , n21397 );
nand ( n21399 , n21210 , n21398 );
not ( n21400 , n21399 );
nand ( n21401 , n21162 , n21093 );
not ( n21402 , RI15b4ff50_593);
and ( n21403 , n21198 , n21402 );
nand ( n21404 , n21401 , n21403 );
nor ( n21405 , n21093 , RI15b4ff50_593);
not ( n21406 , n21405 );
nand ( n21407 , n21093 , RI15b4ff50_593);
nand ( n21408 , n21406 , n21407 );
nand ( n21409 , n21204 , n21408 );
nand ( n21410 , n21404 , n21409 );
not ( n21411 , n21410 );
or ( n21412 , n21400 , n21411 );
not ( n21413 , n21210 );
nand ( n21414 , n21413 , n21397 );
nand ( n21415 , n21412 , n21414 );
nand ( n21416 , n21393 , n21415 );
and ( n21417 , n21369 , n20672 );
not ( n21418 , n21369 );
and ( n21419 , n21418 , RI15b50298_600);
nor ( n21420 , n21417 , n21419 );
nand ( n21421 , n20846 , n21420 );
not ( n21422 , RI15b50220_599);
not ( n21423 , n21367 );
or ( n21424 , n21422 , n21423 );
not ( n21425 , n21367 );
and ( n21426 , n21425 , n20914 );
nor ( n21427 , n21426 , n20917 );
nand ( n21428 , n21424 , n21427 );
not ( n21429 , n21428 );
nand ( n21430 , n21429 , n20906 );
and ( n21431 , n21421 , n21430 );
not ( n21432 , n21058 );
not ( n21433 , n21365 );
or ( n21434 , n21432 , n21433 );
not ( n21435 , n21365 );
and ( n21436 , n21435 , RI15b50130_597);
not ( n21437 , n21061 );
nor ( n21438 , n21436 , n21437 );
nand ( n21439 , n21434 , n21438 );
not ( n21440 , n21439 );
nand ( n21441 , n21217 , n21440 );
buf ( n21442 , n21441 );
and ( n21443 , n21367 , RI15b501a8_598);
not ( n21444 , n21367 );
and ( n21445 , n21444 , n20916 );
nor ( n21446 , n21443 , n21445 );
nand ( n21447 , n20962 , n21446 );
nand ( n21448 , n21431 , n21442 , n21447 );
or ( n21449 , n21416 , n21448 );
nor ( n21450 , n21017 , n21387 );
nand ( n21451 , n21441 , n21450 );
not ( n21452 , n21217 );
nand ( n21453 , n21452 , n21439 );
nand ( n21454 , n21451 , n21453 );
and ( n21455 , n21454 , n21431 , n21447 );
nor ( n21456 , n20962 , n21446 );
nand ( n21457 , n21456 , n21430 );
not ( n21458 , n20906 );
nand ( n21459 , n21458 , n21428 );
nand ( n21460 , n21457 , n21459 );
nand ( n21461 , n21460 , n21421 );
not ( n21462 , n20847 );
not ( n21463 , n21420 );
nand ( n21464 , n21462 , n21463 );
nand ( n21465 , n21461 , n21464 );
nor ( n21466 , n21455 , n21465 );
nand ( n21467 , n21449 , n21466 );
and ( n21468 , n21370 , n21250 );
not ( n21469 , n21370 );
and ( n21470 , n21469 , RI15b50310_601);
nor ( n21471 , n21468 , n21470 );
nand ( n21472 , n21467 , n21471 );
not ( n21473 , n21371 );
not ( n21474 , n21473 );
not ( n21475 , RI15b50388_602);
and ( n21476 , n21474 , n21475 );
and ( n21477 , n21473 , RI15b50388_602);
nor ( n21478 , n21476 , n21477 );
nor ( n21479 , n21472 , n21478 );
and ( n21480 , RI15b504f0_605 , n21374 );
not ( n21481 , RI15b504f0_605);
not ( n21482 , n21374 );
and ( n21483 , n21481 , n21482 );
nor ( n21484 , n21480 , n21483 );
not ( n21485 , RI15b50478_604);
not ( n21486 , n21373 );
not ( n21487 , n21486 );
or ( n21488 , n21485 , n21487 );
or ( n21489 , n21486 , RI15b50478_604);
nand ( n21490 , n21488 , n21489 );
and ( n21491 , n21372 , n21280 );
not ( n21492 , n21372 );
and ( n21493 , n21492 , RI15b50400_603);
nor ( n21494 , n21491 , n21493 );
nand ( n21495 , n21484 , n21490 , n21494 );
and ( n21496 , n21482 , RI15b505e0_607);
or ( n21497 , n21482 , n21260 );
nand ( n21498 , n21497 , n21262 );
nor ( n21499 , n21496 , n21498 );
and ( n21500 , n21482 , RI15b50568_606);
or ( n21501 , n21482 , n21286 );
nand ( n21502 , n21501 , n21288 );
nor ( n21503 , n21500 , n21502 );
nor ( n21504 , n21495 , n21499 , n21503 );
and ( n21505 , n21479 , n21504 );
and ( n21506 , n21482 , RI15b50658_608);
or ( n21507 , n21482 , n20713 );
nand ( n21508 , n21507 , n20716 );
nor ( n21509 , n21506 , n21508 );
not ( n21510 , n21509 );
nand ( n21511 , n21505 , n21510 );
and ( n21512 , n21482 , RI15b506d0_609);
or ( n21513 , n21482 , n21297 );
nand ( n21514 , n21513 , n21299 );
nor ( n21515 , n21512 , n21514 );
nor ( n21516 , n21511 , n21515 );
and ( n21517 , n21482 , RI15b50748_610);
or ( n21518 , n21482 , n20703 );
nand ( n21519 , n21518 , n20706 );
nor ( n21520 , n21517 , n21519 );
not ( n21521 , n21520 );
and ( n21522 , n21516 , n21521 );
buf ( n21523 , n21522 );
and ( n21524 , n21482 , RI15b507c0_611);
or ( n21525 , n21482 , n21307 );
nand ( n21526 , n21525 , n21309 );
nor ( n21527 , n21524 , n21526 );
not ( n21528 , n21527 );
and ( n21529 , n21523 , n21528 );
not ( n21530 , n21376 );
and ( n21531 , n21530 , RI15b50838_612);
not ( n21532 , n21530 );
and ( n21533 , n21532 , n21314 );
nor ( n21534 , n21531 , n21533 );
not ( n21535 , n21534 );
and ( n21536 , n21529 , n21535 );
nand ( n21537 , n21383 , n21536 );
not ( n21538 , n21377 );
not ( n21539 , n21538 );
nand ( n21540 , n21539 , n21323 );
nand ( n21541 , n21538 , RI15b50928_614);
and ( n21542 , n21540 , n21541 , n21327 );
not ( n21543 , n21542 );
and ( n21544 , n21537 , n21543 );
not ( n21545 , n21537 );
and ( n21546 , n21545 , n21542 );
nor ( n21547 , n21544 , n21546 );
nor ( n21548 , n18120 , n18078 );
not ( n21549 , n21548 );
and ( n21550 , n20731 , RI15b4c0f8_460);
nor ( n21551 , n21550 , n18058 );
nand ( n21552 , n21551 , n18064 );
nand ( n21553 , n21336 , n21552 );
nand ( n21554 , n18051 , n21553 );
not ( n21555 , n21554 );
not ( n21556 , n21555 );
not ( n21557 , n21556 );
nor ( n21558 , n21549 , n21557 );
buf ( n21559 , n21558 );
not ( n21560 , n21559 );
buf ( n21561 , n21560 );
buf ( n21562 , n21561 );
not ( n21563 , n21562 );
buf ( n21564 , n21563 );
not ( n21565 , n21564 );
or ( n21566 , n21547 , n21565 );
nor ( n21567 , n21364 , n21091 );
and ( n21568 , n21567 , n21366 );
nand ( n21569 , n21568 , n20670 );
and ( n21570 , n21569 , RI15b50298_600);
not ( n21571 , n21569 );
and ( n21572 , n21571 , n20672 );
nor ( n21573 , n21570 , n21572 );
not ( n21574 , n21573 );
not ( n21575 , n20848 );
or ( n21576 , n21574 , n21575 );
and ( n21577 , n21568 , RI15b501a8_598);
not ( n21578 , n21568 );
and ( n21579 , n21578 , n20916 );
nor ( n21580 , n21577 , n21579 );
not ( n21581 , n21580 );
nand ( n21582 , n20962 , n21581 );
or ( n21583 , n21568 , n20911 );
and ( n21584 , n21568 , n20914 );
nor ( n21585 , n21584 , n20917 );
nand ( n21586 , n21583 , n21585 );
not ( n21587 , n21586 );
nand ( n21588 , n20906 , n21587 );
nand ( n21589 , n21582 , n21588 );
not ( n21590 , n21452 );
not ( n21591 , RI15b50130_597);
not ( n21592 , n21567 );
not ( n21593 , n21592 );
or ( n21594 , n21591 , n21593 );
and ( n21595 , n21567 , n21058 );
nor ( n21596 , n21595 , n21437 );
nand ( n21597 , n21594 , n21596 );
not ( n21598 , n21597 );
and ( n21599 , n21590 , n21598 );
nor ( n21600 , n21589 , n21599 );
not ( n21601 , n21600 );
not ( n21602 , n21162 );
not ( n21603 , n21198 );
not ( n21604 , n21603 );
and ( n21605 , n21602 , n21604 );
nor ( n21606 , n21605 , n21405 );
nand ( n21607 , n21202 , n21606 );
nand ( n21608 , n21210 , n21397 );
and ( n21609 , n21607 , n21608 );
nor ( n21610 , n21210 , n21397 );
nor ( n21611 , n21609 , n21610 );
and ( n21612 , n21592 , n21020 );
not ( n21613 , n21592 );
and ( n21614 , n21613 , RI15b500b8_596);
nor ( n21615 , n21612 , n21614 );
not ( n21616 , n21615 );
and ( n21617 , n21389 , n21616 );
or ( n21618 , n21611 , n21617 );
nand ( n21619 , n21390 , n21615 );
nand ( n21620 , n21618 , n21619 );
not ( n21621 , n21620 );
or ( n21622 , n21601 , n21621 );
not ( n21623 , n21589 );
not ( n21624 , n21590 );
nand ( n21625 , n21624 , n21597 );
not ( n21626 , n21625 );
and ( n21627 , n21623 , n21626 );
not ( n21628 , n20962 );
nand ( n21629 , n21628 , n21580 );
not ( n21630 , n21588 );
or ( n21631 , n21629 , n21630 );
nand ( n21632 , n20907 , n21586 );
nand ( n21633 , n21631 , n21632 );
nor ( n21634 , n21627 , n21633 );
nand ( n21635 , n21622 , n21634 );
nand ( n21636 , n21576 , n21635 );
buf ( n21637 , n21636 );
and ( n21638 , n20679 , RI15b4ff50_593);
buf ( n21639 , n21638 );
not ( n21640 , n20703 );
and ( n21641 , n21639 , n21640 );
not ( n21642 , n20706 );
nor ( n21643 , n21641 , n21642 );
not ( n21644 , n21639 );
nand ( n21645 , n21644 , RI15b50748_610);
and ( n21646 , n21643 , n21645 );
and ( n21647 , n21639 , n21306 );
not ( n21648 , n21309 );
nor ( n21649 , n21647 , n21648 );
not ( n21650 , n21639 );
nand ( n21651 , n21650 , RI15b507c0_611);
and ( n21652 , n21649 , n21651 );
nand ( n21653 , n21646 , n21652 );
not ( n21654 , n20847 );
not ( n21655 , n21573 );
and ( n21656 , n21654 , n21655 );
not ( n21657 , n21249 );
nand ( n21658 , n21657 , RI15b4ff50_593);
and ( n21659 , n21658 , n21250 );
not ( n21660 , n21658 );
and ( n21661 , n21660 , RI15b50310_601);
nor ( n21662 , n21659 , n21661 );
nor ( n21663 , n21656 , n21662 );
not ( n21664 , n21639 );
and ( n21665 , n21664 , RI15b504f0_605);
not ( n21666 , n21664 );
and ( n21667 , n21666 , n21268 );
nor ( n21668 , n21665 , n21667 );
and ( n21669 , n21638 , n21375 );
not ( n21670 , n21669 );
and ( n21671 , n21670 , RI15b50838_612);
not ( n21672 , n21670 );
and ( n21673 , n21672 , n21314 );
nor ( n21674 , n21671 , n21673 );
nand ( n21675 , n21271 , RI15b4ff50_593);
and ( n21676 , n21675 , n20678 );
not ( n21677 , n21675 );
and ( n21678 , n21677 , RI15b50478_604);
nor ( n21679 , n21676 , n21678 );
not ( n21680 , n21277 );
nand ( n21681 , n21680 , RI15b4ff50_593);
and ( n21682 , n21681 , n21280 );
not ( n21683 , n21681 );
and ( n21684 , n21683 , RI15b50400_603);
nor ( n21685 , n21682 , n21684 );
not ( n21686 , RI15b50388_602);
or ( n21687 , n20674 , n21402 );
not ( n21688 , n21687 );
or ( n21689 , n21686 , n21688 );
or ( n21690 , n21687 , RI15b50388_602);
nand ( n21691 , n21689 , n21690 );
nor ( n21692 , n21679 , n21685 , n21691 );
nand ( n21693 , n21663 , n21668 , n21674 , n21692 );
nor ( n21694 , n21653 , n21693 );
and ( n21695 , n21639 , n21296 );
not ( n21696 , n21299 );
nor ( n21697 , n21695 , n21696 );
nand ( n21698 , n21650 , RI15b506d0_609);
and ( n21699 , n21697 , n21698 );
not ( n21700 , n20713 );
and ( n21701 , n21639 , n21700 );
not ( n21702 , n20716 );
nor ( n21703 , n21701 , n21702 );
nand ( n21704 , n21664 , RI15b50658_608);
and ( n21705 , n21703 , n21704 );
and ( n21706 , n21639 , n21259 );
not ( n21707 , n21262 );
nor ( n21708 , n21706 , n21707 );
nand ( n21709 , n21650 , RI15b505e0_607);
and ( n21710 , n21708 , n21709 );
not ( n21711 , n21286 );
and ( n21712 , n21639 , n21711 );
not ( n21713 , n21288 );
nor ( n21714 , n21712 , n21713 );
nand ( n21715 , n21664 , RI15b50568_606);
and ( n21716 , n21714 , n21715 );
and ( n21717 , n21699 , n21705 , n21710 , n21716 );
nand ( n21718 , n21669 , RI15b50838_612);
and ( n21719 , RI15b508b0_613 , n21718 );
not ( n21720 , RI15b508b0_613);
not ( n21721 , n21718 );
and ( n21722 , n21720 , n21721 );
nor ( n21723 , n21719 , n21722 );
and ( n21724 , n21694 , n21717 , n21723 );
nand ( n21725 , n21637 , n21724 );
not ( n21726 , RI15b50928_614);
buf ( n21727 , n21718 );
not ( n21728 , n21727 );
not ( n21729 , n21728 );
not ( n21730 , n21729 );
or ( n21731 , n21726 , n21730 );
and ( n21732 , n21728 , n21323 );
not ( n21733 , n21327 );
nor ( n21734 , n21732 , n21733 );
nand ( n21735 , n21731 , n21734 );
and ( n21736 , n21725 , n21735 );
nor ( n21737 , n21725 , n21735 );
nor ( n21738 , n21736 , n21737 );
not ( n21739 , n21738 );
not ( n21740 , n21351 );
not ( n21741 , n20849 );
and ( n21742 , n21740 , n21741 );
not ( n21743 , n21742 );
buf ( n21744 , n21743 );
buf ( n21745 , n21744 );
not ( n21746 , n21745 );
buf ( n21747 , n21746 );
buf ( n21748 , n21747 );
and ( n21749 , n21739 , n21748 );
or ( n21750 , n18162 , RI15b51120_631);
not ( n21751 , n21750 );
and ( n21752 , n21751 , RI15b57fc0_867);
nor ( n21753 , n21749 , n21752 );
nand ( n21754 , n21566 , n21753 );
nor ( n21755 , n21363 , n21754 );
not ( n21756 , n17551 );
not ( n21757 , n21756 );
not ( n21758 , RI15b570c0_835);
not ( n21759 , n21758 );
and ( n21760 , n21757 , n21759 );
and ( n21761 , n17552 , n21758 );
nor ( n21762 , n21760 , n21761 );
not ( n21763 , n21762 );
or ( n21764 , n17507 , n18170 );
buf ( n21765 , n21764 );
buf ( n21766 , n21765 );
buf ( n21767 , n21766 );
buf ( n21768 , n21767 );
buf ( n21769 , n21768 );
buf ( n21770 , n21769 );
buf ( n21771 , n21770 );
and ( n21772 , n21763 , n21771 );
not ( n21773 , n17550 );
buf ( n21774 , n18176 );
buf ( n21775 , n21774 );
buf ( n21776 , n21775 );
buf ( n21777 , n21776 );
nand ( n21778 , n21773 , n21777 );
not ( n21779 , n21349 );
not ( n21780 , n21335 );
or ( n21781 , n21779 , n21780 );
nand ( n21782 , n21548 , n21555 );
nand ( n21783 , n21781 , n21782 );
nor ( n21784 , n18121 , n18131 );
and ( n21785 , n21784 , n18077 );
and ( n21786 , n18157 , n18218 );
nand ( n21787 , n21786 , n18164 , n18169 );
or ( n21788 , n21783 , n21785 , n21787 );
not ( n21789 , n21788 );
and ( n21790 , n21778 , n21789 );
not ( n21791 , n21790 );
and ( n21792 , n21791 , RI15b570c0_835);
not ( n21793 , n21773 );
buf ( n21794 , n21777 );
and ( n21795 , n21793 , n21794 );
and ( n21796 , n21795 , n21758 );
nor ( n21797 , n21772 , n21792 , n21796 );
nand ( n21798 , n21755 , n21797 );
buf ( n21799 , n21798 );
buf ( n21800 , RI15b3e9d0_1);
buf ( n21801 , n21800 );
not ( n21802 , n17576 );
not ( n21803 , RI15b56a30_821);
not ( n21804 , n21803 );
nand ( n21805 , n17530 , RI15b56760_815);
not ( n21806 , n21805 );
not ( n21807 , n21806 );
or ( n21808 , n21804 , n21807 );
or ( n21809 , n21806 , n21803 );
nand ( n21810 , n21808 , n21809 );
not ( n21811 , n21810 );
nand ( n21812 , n17527 , RI15b56760_815);
xnor ( n21813 , n21812 , RI15b56940_819);
not ( n21814 , n21813 );
nand ( n21815 , n17572 , n17511 );
not ( n21816 , RI15b568c8_818);
not ( n21817 , n21816 );
buf ( n21818 , n17525 );
not ( n21819 , RI15b56760_815);
nor ( n21820 , n21818 , n21819 );
not ( n21821 , n21820 );
or ( n21822 , n21817 , n21821 );
not ( n21823 , RI15b568c8_818);
or ( n21824 , n21820 , n21823 );
nand ( n21825 , n21822 , n21824 );
nor ( n21826 , n21815 , n21825 );
nand ( n21827 , n21814 , n21826 );
not ( n21828 , n17529 );
buf ( n21829 , n17528 );
not ( n21830 , RI15b56760_815);
nor ( n21831 , n21829 , n21830 );
not ( n21832 , n21831 );
or ( n21833 , n21828 , n21832 );
or ( n21834 , n21831 , n17529 );
nand ( n21835 , n21833 , n21834 );
nor ( n21836 , n21827 , n21835 );
nand ( n21837 , n21811 , n21836 );
not ( n21838 , RI15b56aa8_822);
not ( n21839 , n21838 );
not ( n21840 , n17531 );
not ( n21841 , RI15b56760_815);
nor ( n21842 , n21840 , n21841 );
not ( n21843 , n21842 );
or ( n21844 , n21839 , n21843 );
or ( n21845 , n21842 , n21838 );
nand ( n21846 , n21844 , n21845 );
nor ( n21847 , n21837 , n21846 );
not ( n21848 , n17532 );
nand ( n21849 , n21848 , RI15b56760_815);
and ( n21850 , n21849 , RI15b56b20_823);
not ( n21851 , n21849 );
and ( n21852 , n21851 , n17533 );
nor ( n21853 , n21850 , n21852 );
and ( n21854 , n21847 , n21853 );
buf ( n21855 , n17534 );
nand ( n21856 , n21855 , RI15b56760_815);
and ( n21857 , n21856 , RI15b56b98_824);
not ( n21858 , n21856 );
not ( n21859 , RI15b56b98_824);
and ( n21860 , n21858 , n21859 );
nor ( n21861 , n21857 , n21860 );
nand ( n21862 , n21854 , n21861 );
not ( n21863 , n17536 );
buf ( n21864 , n17535 );
not ( n21865 , RI15b56760_815);
nor ( n21866 , n21864 , n21865 );
not ( n21867 , n21866 );
or ( n21868 , n21863 , n21867 );
or ( n21869 , n21866 , n17536 );
nand ( n21870 , n21868 , n21869 );
nor ( n21871 , n21862 , n21870 );
buf ( n21872 , n17537 );
nand ( n21873 , n21872 , RI15b56760_815);
and ( n21874 , n21873 , RI15b56c88_826);
not ( n21875 , n21873 );
not ( n21876 , RI15b56c88_826);
and ( n21877 , n21875 , n21876 );
nor ( n21878 , n21874 , n21877 );
nand ( n21879 , n21871 , n21878 );
nand ( n21880 , n17538 , RI15b56760_815);
not ( n21881 , RI15b56d00_827);
and ( n21882 , n21880 , n21881 );
not ( n21883 , n21880 );
and ( n21884 , n21883 , RI15b56d00_827);
nor ( n21885 , n21882 , n21884 );
nor ( n21886 , n21879 , n21885 );
not ( n21887 , n17539 );
nand ( n21888 , n21887 , RI15b56760_815);
and ( n21889 , n21888 , RI15b56d78_828);
not ( n21890 , n21888 );
and ( n21891 , n21890 , n17540 );
nor ( n21892 , n21889 , n21891 );
and ( n21893 , n21886 , n21892 );
buf ( n21894 , n17541 );
nand ( n21895 , n21894 , RI15b56760_815);
and ( n21896 , n21895 , RI15b56df0_829);
not ( n21897 , n21895 );
not ( n21898 , RI15b56df0_829);
and ( n21899 , n21897 , n21898 );
nor ( n21900 , n21896 , n21899 );
nand ( n21901 , n21893 , n21900 );
not ( n21902 , n17543 );
not ( n21903 , n17542 );
nand ( n21904 , n21903 , RI15b56760_815);
not ( n21905 , n21904 );
not ( n21906 , n21905 );
or ( n21907 , n21902 , n21906 );
or ( n21908 , n21905 , n17543 );
nand ( n21909 , n21907 , n21908 );
nor ( n21910 , n21901 , n21909 );
buf ( n21911 , n21910 );
buf ( n21912 , n17544 );
nand ( n21913 , n21912 , RI15b56760_815);
and ( n21914 , n21913 , RI15b56ee0_831);
not ( n21915 , n21913 );
not ( n21916 , RI15b56ee0_831);
and ( n21917 , n21915 , n21916 );
nor ( n21918 , n21914 , n21917 );
not ( n21919 , n21918 );
nor ( n21920 , n21911 , n21919 );
and ( n21921 , n21802 , n21920 );
not ( n21922 , n18187 );
not ( n21923 , RI15b57750_849);
nor ( n21924 , n21923 , n18190 );
nand ( n21925 , n21924 , RI15b577c8_850);
not ( n21926 , RI15b57840_851);
nor ( n21927 , n21925 , n21926 );
and ( n21928 , RI15b578b8_852 , RI15b57930_853);
nand ( n21929 , n21927 , n21928 );
not ( n21930 , RI15b579a8_854);
nor ( n21931 , n21929 , n21930 );
and ( n21932 , n21931 , RI15b57a20_855);
nand ( n21933 , n21932 , RI15b57a98_856);
not ( n21934 , RI15b57b10_857);
nor ( n21935 , n21933 , n21934 );
not ( n21936 , RI15b57b88_858);
not ( n21937 , RI15b57c00_859);
nor ( n21938 , n21936 , n21937 );
and ( n21939 , n21935 , n21938 );
not ( n21940 , RI15b57c78_860);
not ( n21941 , RI15b57cf0_861);
nor ( n21942 , n21940 , n21941 );
nand ( n21943 , n21939 , n21942 );
not ( n21944 , n21943 );
or ( n21945 , n21922 , n21944 );
not ( n21946 , n18150 );
nand ( n21947 , n21945 , n21946 );
and ( n21948 , n21947 , RI15b57de0_863);
not ( n21949 , n18074 );
not ( n21950 , n21949 );
nor ( n21951 , n18082 , RI15b55950_785);
not ( n21952 , RI15b559c8_786);
and ( n21953 , n21951 , n21952 );
not ( n21954 , RI15b55a40_787);
nand ( n21955 , n21953 , n21954 );
nor ( n21956 , n21955 , RI15b55ab8_788);
not ( n21957 , RI15b55b30_789);
and ( n21958 , n21956 , n21957 );
not ( n21959 , RI15b55ba8_790);
nand ( n21960 , n21958 , n21959 );
nor ( n21961 , n21960 , RI15b55c20_791);
not ( n21962 , RI15b55c98_792);
and ( n21963 , n21961 , n21962 );
not ( n21964 , RI15b55d10_793);
nand ( n21965 , n21963 , n21964 );
nor ( n21966 , n21965 , RI15b55d88_794);
not ( n21967 , RI15b55e00_795);
and ( n21968 , n21966 , n21967 );
not ( n21969 , RI15b55e78_796);
nand ( n21970 , n21968 , n21969 );
nor ( n21971 , n21970 , RI15b55ef0_797);
not ( n21972 , RI15b55f68_798);
and ( n21973 , n21971 , n21972 );
not ( n21974 , n21973 );
or ( n21975 , n21950 , n21974 );
nand ( n21976 , n21949 , n18084 );
not ( n21977 , n18148 );
nand ( n21978 , n18099 , n21977 );
and ( n21979 , n21976 , n21978 );
nand ( n21980 , n21975 , n21979 );
and ( n21981 , n21980 , RI15b55fe0_799);
or ( n21982 , n18074 , n18084 );
or ( n21983 , n21982 , n21973 , RI15b55fe0_799);
not ( n21984 , RI15b57de0_863);
and ( n21985 , n21944 , n21984 , RI15b57d68_862);
not ( n21986 , RI15b57d68_862);
and ( n21987 , n21986 , RI15b57de0_863);
nor ( n21988 , n21985 , n21987 );
or ( n21989 , n21922 , n21988 );
nand ( n21990 , n21983 , n21989 );
nor ( n21991 , n21948 , n21981 , n21990 );
or ( n21992 , n21991 , n18078 );
and ( n21993 , n18177 , RI15b57de0_863);
and ( n21994 , n18219 , RI15b56ee0_831);
nor ( n21995 , n21993 , n21994 , n21751 );
nand ( n21996 , n21992 , n21995 );
nor ( n21997 , n21921 , n21996 );
nand ( n21998 , n21911 , n17507 );
not ( n21999 , n21998 );
not ( n22000 , n17565 );
or ( n22001 , n21999 , n22000 );
nand ( n22002 , n22001 , n21919 );
nand ( n22003 , n21997 , n22002 );
buf ( n22004 , n22003 );
buf ( n22005 , RI15b3ea48_2);
buf ( n22006 , n22005 );
buf ( n22007 , RI15b3ea48_2);
buf ( n22008 , n22007 );
buf ( n22009 , RI15b3e9d0_1);
buf ( n22010 , n22009 );
not ( n22011 , n20637 );
not ( n22012 , RI15b66408_1354);
not ( n22013 , n22012 );
nor ( n22014 , RI15b65850_1329 , RI15b658c8_1330);
not ( n22015 , RI15b65940_1331);
and ( n22016 , n22014 , n22015 );
not ( n22017 , RI15b659b8_1332);
nand ( n22018 , n22016 , n22017 );
nor ( n22019 , n22018 , RI15b65a30_1333);
not ( n22020 , RI15b65aa8_1334);
and ( n22021 , n22019 , n22020 );
not ( n22022 , RI15b65b20_1335);
nand ( n22023 , n22021 , n22022 );
nor ( n22024 , n22023 , RI15b65b98_1336);
not ( n22025 , RI15b65c10_1337);
nand ( n22026 , n22024 , n22025 );
nor ( n22027 , n22026 , RI15b65c88_1338);
not ( n22028 , RI15b65d00_1339);
not ( n22029 , RI15b65d78_1340);
not ( n22030 , RI15b65df0_1341);
and ( n22031 , n22027 , n22028 , n22029 , n22030 );
not ( n22032 , RI15b65e68_1342);
nand ( n22033 , n22031 , n22032 );
nor ( n22034 , n22033 , RI15b65ee0_1343);
not ( n22035 , RI15b65f58_1344);
not ( n22036 , RI15b65fd0_1345);
not ( n22037 , RI15b66048_1346);
and ( n22038 , n22034 , n22035 , n22036 , n22037 );
not ( n22039 , RI15b660c0_1347);
and ( n22040 , n22038 , n22039 );
not ( n22041 , RI15b66138_1348);
nand ( n22042 , n22040 , n22041 );
nor ( n22043 , n22042 , RI15b661b0_1349);
not ( n22044 , RI15b66228_1350);
nand ( n22045 , n22043 , n22044 );
not ( n22046 , n22045 );
not ( n22047 , RI15b662a0_1351);
nand ( n22048 , n22046 , n22047 );
nor ( n22049 , n22048 , RI15b66318_1352);
not ( n22050 , RI15b66390_1353);
nand ( n22051 , n22049 , n22050 );
not ( n22052 , n22051 );
or ( n22053 , n22013 , n22052 );
not ( n22054 , RI15b66480_1355);
nand ( n22055 , n22054 , RI15b66408_1354);
nand ( n22056 , n22053 , n22055 );
not ( n22057 , n22056 );
not ( n22058 , n22048 );
not ( n22059 , RI15b66318_1352);
nand ( n22060 , n22058 , n22059 );
nand ( n22061 , n22060 , RI15b666d8_1360);
not ( n22062 , n22061 );
not ( n22063 , RI15b66390_1353);
and ( n22064 , n22062 , n22063 );
and ( n22065 , n22061 , RI15b66390_1353);
nor ( n22066 , n22064 , n22065 );
not ( n22067 , n22051 );
nand ( n22068 , n22067 , RI15b66480_1355);
nand ( n22069 , n22057 , n22066 , n22068 );
not ( n22070 , n22069 );
not ( n22071 , RI15b66408_1354);
nand ( n22072 , n22071 , n22054 );
nor ( n22073 , n22051 , n22072 );
not ( n22074 , n22073 );
not ( n22075 , RI15b664f8_1356);
and ( n22076 , n22074 , n22075 );
buf ( n22077 , n22073 );
and ( n22078 , n22077 , RI15b664f8_1356);
nor ( n22079 , n22076 , n22078 );
nand ( n22080 , n22070 , n22079 );
not ( n22081 , n22080 );
not ( n22082 , n22081 );
not ( n22083 , RI15b664f8_1356);
and ( n22084 , n22073 , n22083 );
buf ( n22085 , n22084 );
not ( n22086 , n22085 );
not ( n22087 , n22086 );
and ( n22088 , n22082 , n22087 );
not ( n22089 , n22080 );
and ( n22090 , n22089 , n22086 );
nor ( n22091 , n22088 , n22090 );
not ( n22092 , n22091 );
or ( n22093 , n22011 , n22092 );
or ( n22094 , n20638 , RI15b666d8_1360);
nand ( n22095 , n22093 , n22094 );
and ( n22096 , n22095 , RI15b66570_1357);
and ( n22097 , n20637 , RI15b666d8_1360);
not ( n22098 , RI15b66570_1357);
nand ( n22099 , n22097 , n22098 );
nor ( n22100 , n22091 , n22099 );
nor ( n22101 , n22096 , n22100 );
buf ( n22102 , n22101 );
nand ( n22103 , RI15b3fc90_41 , RI15b3fd08_42);
not ( n22104 , n22103 );
nand ( n22105 , n22104 , RI15b3fd80_43);
and ( n22106 , n22105 , n20440 );
not ( n22107 , n22105 );
and ( n22108 , n22107 , RI15b3fdf8_44);
nor ( n22109 , n22106 , n22108 );
not ( n22110 , n22109 );
not ( n22111 , RI15b3fd80_43);
not ( n22112 , n22103 );
or ( n22113 , n22111 , n22112 );
nand ( n22114 , n20427 , n20417 );
nand ( n22115 , n22113 , n22114 );
nand ( n22116 , n22110 , n22115 );
nand ( n22117 , n20422 , RI15b3fd08_42);
buf ( n22118 , n22117 );
nor ( n22119 , n22116 , n22118 );
not ( n22120 , n22117 );
not ( n22121 , n22109 );
or ( n22122 , n22120 , n22121 );
not ( n22123 , n22115 );
nand ( n22124 , n22109 , n22123 );
nand ( n22125 , n22122 , n22124 );
nor ( n22126 , n22119 , n22125 );
and ( n22127 , n22115 , n22117 );
not ( n22128 , n22127 );
not ( n22129 , n22117 );
nand ( n22130 , n22123 , n22129 );
nand ( n22131 , n22128 , n22130 );
and ( n22132 , n22126 , n22131 );
or ( n22133 , n20422 , RI15b3fd08_42);
not ( n22134 , n22133 );
nand ( n22135 , n22132 , n22134 );
not ( n22136 , n22126 );
not ( n22137 , n22134 );
and ( n22138 , n22136 , n22137 );
buf ( n22139 , n22131 );
nor ( n22140 , n22126 , n22139 );
nor ( n22141 , n22138 , n22140 );
nand ( n22142 , n22135 , n22141 );
not ( n22143 , n22142 );
and ( n22144 , n22131 , n22134 );
not ( n22145 , n22131 );
and ( n22146 , n22145 , n22133 );
nor ( n22147 , n22144 , n22146 );
not ( n22148 , n22147 );
nand ( n22149 , n22143 , n22148 );
buf ( n22150 , n22103 );
or ( n22151 , n22149 , n22150 );
or ( n22152 , n22102 , n22151 );
not ( n22153 , RI15b66138_1348);
not ( n22154 , n22040 );
nand ( n22155 , n22154 , RI15b666d8_1360);
not ( n22156 , n22155 );
or ( n22157 , n22153 , n22156 );
or ( n22158 , n22155 , RI15b66138_1348);
nand ( n22159 , n22157 , n22158 );
buf ( n22160 , n22034 );
and ( n22161 , n22160 , n22035 );
nand ( n22162 , n22161 , n22036 );
nand ( n22163 , n22162 , RI15b666d8_1360);
not ( n22164 , n22163 );
not ( n22165 , RI15b66048_1346);
and ( n22166 , n22164 , n22165 );
and ( n22167 , n22163 , RI15b66048_1346);
nor ( n22168 , n22166 , n22167 );
not ( n22169 , n22161 );
nand ( n22170 , n22169 , RI15b666d8_1360);
not ( n22171 , n22170 );
not ( n22172 , RI15b65fd0_1345);
and ( n22173 , n22171 , n22172 );
and ( n22174 , n22170 , RI15b65fd0_1345);
nor ( n22175 , n22173 , n22174 );
nand ( n22176 , n22168 , n22175 );
not ( n22177 , n22176 );
not ( n22178 , n22038 );
nand ( n22179 , n22178 , RI15b666d8_1360);
not ( n22180 , n22179 );
not ( n22181 , RI15b660c0_1347);
and ( n22182 , n22180 , n22181 );
and ( n22183 , n22179 , RI15b660c0_1347);
nor ( n22184 , n22182 , n22183 );
nand ( n22185 , n22177 , n22184 );
nor ( n22186 , n22159 , n22185 );
not ( n22187 , n22186 );
or ( n22188 , n22187 , n20638 );
nand ( n22189 , n22188 , n22094 );
buf ( n22190 , n22042 );
nand ( n22191 , n22190 , RI15b666d8_1360);
not ( n22192 , n22191 );
not ( n22193 , RI15b661b0_1349);
and ( n22194 , n22192 , n22193 );
and ( n22195 , n22191 , RI15b661b0_1349);
nor ( n22196 , n22194 , n22195 );
not ( n22197 , n22196 );
and ( n22198 , n22189 , n22197 );
not ( n22199 , n22097 );
nor ( n22200 , n22197 , n22199 );
and ( n22201 , n22200 , n22187 );
nor ( n22202 , n22198 , n22201 );
not ( n22203 , n22202 );
buf ( n22204 , n22126 );
buf ( n22205 , n22204 );
buf ( n22206 , n22139 );
not ( n22207 , n22206 );
and ( n22208 , n22205 , n22207 );
not ( n22209 , n20424 );
buf ( n22210 , n22209 );
and ( n22211 , n22208 , n22210 );
and ( n22212 , n22203 , n22211 );
not ( n22213 , n22211 );
and ( n22214 , n22151 , n22213 , n19912 );
not ( n22215 , n20635 );
and ( n22216 , n19914 , n22215 );
not ( n22217 , n22216 );
nor ( n22218 , n22214 , n22217 );
or ( n22219 , n22109 , n22115 );
nor ( n22220 , n22219 , n22133 );
or ( n22221 , n22218 , n22220 );
nand ( n22222 , n22221 , n20623 );
nor ( n22223 , RI15b3fdf8_44 , RI15b3fe70_45);
nand ( n22224 , n22223 , n20417 );
buf ( n22225 , n22118 );
buf ( n22226 , n22225 );
buf ( n22227 , n22226 );
or ( n22228 , n22224 , n22227 );
and ( n22229 , n22222 , n22228 );
nor ( n22230 , n20620 , RI15b44cb8_212);
not ( n22231 , n22230 );
nand ( n22232 , n20621 , n22231 );
nor ( n22233 , n20623 , n20008 );
nand ( n22234 , n20650 , n20630 , n20633 );
or ( n22235 , n22232 , n22233 , n20501 , n22234 );
or ( n22236 , n22235 , n20626 );
nor ( n22237 , n22229 , n22236 );
not ( n22238 , RI15b40848_66);
or ( n22239 , n22237 , n22238 );
nand ( n22240 , n22023 , RI15b666d8_1360);
not ( n22241 , RI15b65b98_1336);
and ( n22242 , n22240 , n22241 );
not ( n22243 , n22240 );
and ( n22244 , n22243 , RI15b65b98_1336);
nor ( n22245 , n22242 , n22244 );
not ( n22246 , RI15b65aa8_1334);
not ( n22247 , n22019 );
nand ( n22248 , n22247 , RI15b666d8_1360);
not ( n22249 , n22248 );
or ( n22250 , n22246 , n22249 );
or ( n22251 , n22248 , RI15b65aa8_1334);
nand ( n22252 , n22250 , n22251 );
not ( n22253 , n22252 );
not ( n22254 , RI15b666d8_1360);
nor ( n22255 , n22021 , n22254 );
and ( n22256 , n22255 , n22022 );
not ( n22257 , n22255 );
and ( n22258 , n22257 , RI15b65b20_1335);
nor ( n22259 , n22256 , n22258 );
not ( n22260 , n22014 );
not ( n22261 , RI15b65a30_1333);
nand ( n22262 , n22018 , RI15b666d8_1360);
not ( n22263 , n22262 );
or ( n22264 , n22261 , n22263 );
or ( n22265 , n22262 , RI15b65a30_1333);
nand ( n22266 , n22264 , n22265 );
and ( n22267 , RI15b65940_1331 , RI15b666d8_1360);
nand ( n22268 , RI15b65850_1329 , RI15b666d8_1360);
nand ( n22269 , RI15b658c8_1330 , RI15b666d8_1360);
nand ( n22270 , n22268 , n22269 );
nor ( n22271 , n22267 , n22270 );
or ( n22272 , n22271 , RI15b659b8_1332);
not ( n22273 , RI15b666d8_1360);
not ( n22274 , n22016 );
not ( n22275 , n22274 );
or ( n22276 , n22273 , n22275 );
nand ( n22277 , n22276 , RI15b659b8_1332);
nand ( n22278 , n22272 , n22277 );
not ( n22279 , n22270 );
or ( n22280 , n22279 , RI15b65940_1331);
or ( n22281 , n22014 , n22254 );
nand ( n22282 , n22281 , RI15b65940_1331);
nand ( n22283 , n22280 , n22282 );
nor ( n22284 , n22260 , n22266 , n22278 , n22283 );
nand ( n22285 , n22253 , n22259 , n22284 );
nor ( n22286 , n22245 , n22285 );
or ( n22287 , n22286 , n22254 );
not ( n22288 , n22287 );
not ( n22289 , RI15b65a30_1333);
not ( n22290 , n22289 );
and ( n22291 , n22288 , n22290 );
and ( n22292 , n22287 , n22266 );
nor ( n22293 , n22291 , n22292 );
not ( n22294 , n22228 );
nor ( n22295 , n22220 , n22294 );
or ( n22296 , n22218 , n22295 );
or ( n22297 , n22293 , n22296 );
or ( n22298 , n20623 , RI15b44bc8_210);
or ( n22299 , n20571 , n22298 );
or ( n22300 , n22228 , n22299 );
nand ( n22301 , n22239 , n22297 , n22300 );
nor ( n22302 , n22212 , n22301 );
nand ( n22303 , n22152 , n22302 );
buf ( n22304 , n22303 );
buf ( n22305 , n22069 );
not ( n22306 , n22305 );
buf ( n22307 , n22079 );
not ( n22308 , n22307 );
or ( n22309 , n22306 , n22308 );
or ( n22310 , n22305 , n22307 );
nand ( n22311 , n22309 , n22310 );
and ( n22312 , n22311 , n22097 );
nor ( n22313 , n22094 , n22083 );
nor ( n22314 , n22312 , n22313 );
buf ( n22315 , n22314 );
or ( n22316 , n22315 , n22151 );
not ( n22317 , n20637 );
not ( n22318 , n22185 );
not ( n22319 , n22318 );
or ( n22320 , n22317 , n22319 );
nand ( n22321 , n22320 , n22094 );
nand ( n22322 , n22321 , n22159 );
not ( n22323 , n22159 );
nand ( n22324 , n22323 , n22185 , n22097 );
and ( n22325 , n22322 , n22324 );
not ( n22326 , n22325 );
and ( n22327 , n22326 , n22211 );
not ( n22328 , RI15b407d0_65);
or ( n22329 , n22237 , n22328 );
not ( n22330 , n22287 );
not ( n22331 , n22017 );
and ( n22332 , n22330 , n22331 );
and ( n22333 , n22287 , n22278 );
nor ( n22334 , n22332 , n22333 );
or ( n22335 , n22334 , n22296 );
or ( n22336 , n20573 , n22298 );
or ( n22337 , n22228 , n22336 );
nand ( n22338 , n22329 , n22335 , n22337 );
nor ( n22339 , n22327 , n22338 );
nand ( n22340 , n22316 , n22339 );
buf ( n22341 , n22340 );
buf ( n22342 , n18226 );
buf ( n22343 , RI15b3e9d0_1);
buf ( n22344 , n22343 );
not ( n22345 , n19918 );
not ( n22346 , n22345 );
not ( n22347 , n19749 );
not ( n22348 , n22347 );
or ( n22349 , n22346 , n22348 );
not ( n22350 , n19937 );
nand ( n22351 , n22349 , n22350 );
and ( n22352 , n22351 , n19756 );
nand ( n22353 , n20565 , n20501 );
buf ( n22354 , n22353 );
buf ( n22355 , n22354 );
buf ( n22356 , n20536 );
or ( n22357 , n22355 , n22356 , RI15b4b450_433);
buf ( n22358 , n20496 );
nand ( n22359 , n22358 , RI15b4a208_394);
not ( n22360 , n22359 );
and ( n22361 , n22360 , n20501 );
not ( n22362 , n22361 );
buf ( n22363 , n19961 );
or ( n22364 , n22362 , n22363 , RI15b49650_369);
nand ( n22365 , n22357 , n22364 );
nor ( n22366 , n22352 , n22365 );
not ( n22367 , n19756 );
buf ( n22368 , n20524 );
not ( n22369 , n22347 );
nand ( n22370 , n22367 , n22368 , n22369 );
and ( n22371 , n20565 , n22356 );
buf ( n22372 , n20612 );
nor ( n22373 , n22371 , n22372 );
not ( n22374 , RI15b4b450_433);
or ( n22375 , n22373 , n22374 );
buf ( n22376 , n22358 );
buf ( n22377 , n22376 );
buf ( n22378 , n22377 );
and ( n22379 , n22378 , n22363 );
not ( n22380 , n20528 );
not ( n22381 , n22358 );
or ( n22382 , n22380 , n22381 );
nand ( n22383 , n22382 , n20518 );
nor ( n22384 , n22379 , n22383 );
or ( n22385 , n22384 , n19962 );
nand ( n22386 , n22375 , n22385 );
nand ( n22387 , n22386 , n20501 );
not ( n22388 , n20639 );
and ( n22389 , n22388 , RI15b4b450_433);
buf ( n22390 , n20653 );
not ( n22391 , n22390 );
and ( n22392 , n22391 , RI15b4a550_401);
buf ( n22393 , n22230 );
buf ( n22394 , n22393 );
buf ( n22395 , n22394 );
buf ( n22396 , n22395 );
not ( n22397 , n22396 );
not ( n22398 , n22397 );
nor ( n22399 , n22389 , n22392 , n22398 );
nand ( n22400 , n22366 , n22370 , n22387 , n22399 );
buf ( n22401 , n22400 );
buf ( n22402 , RI15b3ea48_2);
buf ( n22403 , n22402 );
buf ( n22404 , RI15b3e9d0_1);
buf ( n22405 , n22404 );
buf ( n22406 , RI15b3e9d0_1);
buf ( n22407 , n22406 );
buf ( n22408 , RI15b3ea48_2);
buf ( n22409 , n22408 );
not ( n22410 , n19486 );
not ( n22411 , n19489 );
or ( n22412 , n22410 , n22411 );
or ( n22413 , n19489 , n19486 );
nand ( n22414 , n22412 , n22413 );
nand ( n22415 , n19232 , n22414 );
nand ( n22416 , n19241 , n19254 , n22415 );
buf ( n22417 , n22416 );
buf ( n22418 , n22417 );
not ( n22419 , n22418 );
nor ( n22420 , n19554 , n22419 );
not ( n22421 , n22420 );
nand ( n22422 , n22421 , n19201 );
or ( n22423 , n19591 , n19639 , n19596 , n19629 );
not ( n22424 , n22423 );
and ( n22425 , n22422 , n22424 );
not ( n22426 , n22425 );
nand ( n22427 , RI15b3fb28_38 , RI15b66750_1361);
not ( n22428 , n22427 );
nor ( n22429 , n22428 , RI15b606c0_1155);
not ( n22430 , n22429 );
not ( n22431 , n19551 );
not ( n22432 , n22431 );
or ( n22433 , n22430 , n22432 );
not ( n22434 , n19544 );
not ( n22435 , RI15b60be8_1166);
nand ( n22436 , n22435 , RI15b60c60_1167);
not ( n22437 , n22436 );
buf ( n22438 , n22437 );
not ( n22439 , RI15b60cd8_1168);
and ( n22440 , n22438 , n22439 );
not ( n22441 , n22440 );
nor ( n22442 , RI15b60be8_1166 , RI15b60c60_1167);
nand ( n22443 , n22442 , RI15b60cd8_1168);
nand ( n22444 , n22441 , n22443 );
nand ( n22445 , n22444 , n22429 );
not ( n22446 , n22445 );
nand ( n22447 , n22434 , n22446 );
nand ( n22448 , n22433 , n22447 );
and ( n22449 , n22448 , n22418 );
and ( n22450 , n22449 , n19201 );
or ( n22451 , n22426 , n22450 );
nand ( n22452 , n22451 , RI15b63a50_1265);
not ( n22453 , n22417 );
nor ( n22454 , n22453 , n22429 );
and ( n22455 , n22431 , n22454 );
nand ( n22456 , n22455 , n19201 );
not ( n22457 , n22456 );
buf ( n22458 , n22457 );
not ( n22459 , n22458 );
not ( n22460 , n19544 );
nand ( n22461 , n22416 , n19201 );
not ( n22462 , n22461 );
and ( n22463 , n22460 , n22462 );
buf ( n22464 , n22463 );
buf ( n22465 , n22464 );
nand ( n22466 , n22465 , n22445 );
nand ( n22467 , n22459 , n22466 );
and ( n22468 , n22467 , RI15b61c50_1201);
buf ( n22469 , n19548 );
and ( n22470 , n22469 , n19539 );
nor ( n22471 , n22470 , n22461 );
and ( n22472 , n22471 , n18249 );
not ( n22473 , n19628 );
nand ( n22474 , n22473 , n19598 );
and ( n22475 , n22474 , RI15b62b50_1233);
nor ( n22476 , n22468 , n22472 , n22475 );
nand ( n22477 , n22452 , n22476 );
buf ( n22478 , n22477 );
buf ( n22479 , RI15b3e9d0_1);
buf ( n22480 , n22479 );
not ( n22481 , RI15b56fd0_833);
not ( n22482 , n22481 );
nand ( n22483 , n17547 , RI15b56760_815);
not ( n22484 , n22483 );
not ( n22485 , n22484 );
or ( n22486 , n22482 , n22485 );
or ( n22487 , n22484 , n22481 );
nand ( n22488 , n22486 , n22487 );
not ( n22489 , n22488 );
nand ( n22490 , n21910 , n21918 );
not ( n22491 , n17546 );
buf ( n22492 , n17545 );
not ( n22493 , RI15b56760_815);
nor ( n22494 , n22492 , n22493 );
not ( n22495 , n22494 );
or ( n22496 , n22491 , n22495 );
or ( n22497 , n22494 , n17546 );
nand ( n22498 , n22496 , n22497 );
nor ( n22499 , n22490 , n22498 );
nand ( n22500 , n22489 , n22499 );
not ( n22501 , n17549 );
not ( n22502 , RI15b56760_815);
nor ( n22503 , n17548 , n22502 );
not ( n22504 , n22503 );
or ( n22505 , n22501 , n22504 );
or ( n22506 , n22503 , n17549 );
nand ( n22507 , n22505 , n22506 );
nor ( n22508 , n22500 , n22507 );
nand ( n22509 , n22508 , n21762 );
nand ( n22510 , n21756 , RI15b570c0_835);
not ( n22511 , RI15b57138_836);
and ( n22512 , n22510 , n22511 );
not ( n22513 , n22510 );
and ( n22514 , n22513 , RI15b57138_836);
nor ( n22515 , n22512 , n22514 );
nor ( n22516 , n22509 , n22515 );
nand ( n22517 , n17552 , n17515 );
and ( n22518 , n22517 , RI15b571b0_837);
not ( n22519 , n22517 );
not ( n22520 , RI15b571b0_837);
and ( n22521 , n22519 , n22520 );
nor ( n22522 , n22518 , n22521 );
nand ( n22523 , n22516 , n22522 );
nand ( n22524 , n17552 , n17516 );
not ( n22525 , RI15b57228_838);
and ( n22526 , n22524 , n22525 );
not ( n22527 , n22524 );
and ( n22528 , n22527 , RI15b57228_838);
nor ( n22529 , n22526 , n22528 );
nor ( n22530 , n22523 , n22529 );
buf ( n22531 , n17552 );
not ( n22532 , n17517 );
nand ( n22533 , n22531 , n22532 );
and ( n22534 , n22533 , RI15b572a0_839);
not ( n22535 , n22533 );
and ( n22536 , n22535 , n17518 );
nor ( n22537 , n22534 , n22536 );
nand ( n22538 , n22530 , n22537 );
nand ( n22539 , n22531 , n17519 );
not ( n22540 , RI15b57318_840);
and ( n22541 , n22539 , n22540 );
not ( n22542 , n22539 );
and ( n22543 , n22542 , RI15b57318_840);
nor ( n22544 , n22541 , n22543 );
nor ( n22545 , n22538 , n22544 );
not ( n22546 , n17520 );
nand ( n22547 , n22546 , n22531 );
and ( n22548 , n22547 , RI15b57390_841);
not ( n22549 , n22547 );
and ( n22550 , n22549 , n17521 );
nor ( n22551 , n22548 , n22550 );
and ( n22552 , n22545 , n22551 );
nand ( n22553 , n22531 , n17522 );
and ( n22554 , n22553 , RI15b57408_842);
not ( n22555 , n22553 );
not ( n22556 , RI15b57408_842);
and ( n22557 , n22555 , n22556 );
nor ( n22558 , n22554 , n22557 );
nand ( n22559 , n22552 , n22558 );
not ( n22560 , n17554 );
and ( n22561 , n22560 , RI15b57480_843);
not ( n22562 , n22560 );
and ( n22563 , n22562 , n17555 );
nor ( n22564 , n22561 , n22563 );
nor ( n22565 , n22559 , n22564 );
not ( n22566 , n22565 );
not ( n22567 , n17576 );
not ( n22568 , n17556 );
and ( n22569 , n22568 , RI15b574f8_844);
not ( n22570 , n22568 );
not ( n22571 , RI15b574f8_844);
and ( n22572 , n22570 , n22571 );
nor ( n22573 , n22569 , n22572 );
and ( n22574 , n22567 , n22573 );
not ( n22575 , n22574 );
or ( n22576 , n22566 , n22575 );
not ( n22577 , RI15b55fe0_799);
nand ( n22578 , n21973 , n22577 );
nor ( n22579 , n22578 , RI15b56058_800);
not ( n22580 , RI15b560d0_801);
and ( n22581 , n22579 , n22580 );
not ( n22582 , RI15b56148_802);
nand ( n22583 , n22581 , n22582 );
nor ( n22584 , n22583 , RI15b561c0_803);
not ( n22585 , RI15b56238_804);
and ( n22586 , n22584 , n22585 );
not ( n22587 , RI15b562b0_805);
nand ( n22588 , n22586 , n22587 );
nor ( n22589 , n22588 , RI15b56328_806);
not ( n22590 , RI15b563a0_807);
and ( n22591 , n22589 , n22590 );
not ( n22592 , RI15b56418_808);
nand ( n22593 , n22591 , n22592 );
nor ( n22594 , n22593 , RI15b56490_809);
not ( n22595 , RI15b56508_810);
nand ( n22596 , n22594 , n22595 );
not ( n22597 , n22596 );
not ( n22598 , RI15b56580_811);
nand ( n22599 , n22597 , n22598 );
not ( n22600 , n22599 );
or ( n22601 , n21982 , n18078 );
nor ( n22602 , n22601 , RI15b565f8_812);
and ( n22603 , n22600 , n22602 );
not ( n22604 , n18179 );
not ( n22605 , RI15b58470_877);
or ( n22606 , n22604 , n22605 );
not ( n22607 , n22605 );
nand ( n22608 , RI15b57d68_862 , RI15b57de0_863);
nor ( n22609 , n21943 , n22608 );
not ( n22610 , RI15b57e58_864);
not ( n22611 , RI15b57ed0_865);
nor ( n22612 , n22610 , n22611 );
and ( n22613 , n22609 , n22612 );
not ( n22614 , RI15b57f48_866);
not ( n22615 , RI15b57fc0_867);
nor ( n22616 , n22614 , n22615 );
nand ( n22617 , n22613 , n22616 );
nand ( n22618 , RI15b58038_868 , RI15b580b0_869);
nor ( n22619 , n22617 , n22618 );
and ( n22620 , n22619 , RI15b58128_870 , RI15b581a0_871);
nand ( n22621 , n22620 , RI15b58218_872 , RI15b58290_873);
not ( n22622 , RI15b58308_874);
not ( n22623 , RI15b58380_875);
nor ( n22624 , n22621 , n22622 , n22623 );
and ( n22625 , RI15b583f8_876 , n22624 );
not ( n22626 , n22625 );
or ( n22627 , n22607 , n22626 );
or ( n22628 , n22625 , n22605 );
nand ( n22629 , n22627 , n22628 );
and ( n22630 , n22629 , n18188 );
not ( n22631 , n18102 );
and ( n22632 , n22631 , RI15b56670_813);
and ( n22633 , n18219 , RI15b57570_845);
nor ( n22634 , n22630 , n22632 , n22633 );
nand ( n22635 , n22606 , n22634 );
nor ( n22636 , n22603 , n22635 );
nand ( n22637 , n22576 , n22636 );
buf ( n22638 , n22637 );
not ( n22639 , RI15b60648_1154);
and ( n22640 , n22639 , RI15b605d0_1153);
not ( n22641 , RI15b47d78_316);
and ( n22642 , n22641 , RI15b47d00_315);
nor ( n22643 , n22640 , n22642 );
not ( n22644 , RI15b541e0_735);
nand ( n22645 , n22644 , RI15b54168_734);
and ( n22646 , n22643 , n22645 );
and ( n22647 , n22646 , RI15b450f0_221);
not ( n22648 , n22646 );
and ( n22649 , n22648 , RI15b51558_640);
nor ( n22650 , n22647 , n22649 );
not ( n22651 , n22650 );
buf ( n22652 , n22651 );
buf ( n22653 , RI15b3ea48_2);
buf ( n22654 , n22653 );
buf ( n22655 , RI15b3e9d0_1);
buf ( n22656 , n22655 );
not ( n22657 , n21447 );
buf ( n22658 , n21416 );
not ( n22659 , n21450 );
nand ( n22660 , n22658 , n22659 );
buf ( n22661 , n21442 );
nand ( n22662 , n22660 , n22661 );
nand ( n22663 , n22662 , n21453 );
not ( n22664 , n22663 );
or ( n22665 , n22657 , n22664 );
not ( n22666 , n21456 );
nand ( n22667 , n22665 , n22666 );
not ( n22668 , n22667 );
and ( n22669 , n22668 , n21459 );
not ( n22670 , n21430 );
nor ( n22671 , n22669 , n22670 );
and ( n22672 , n21463 , n22671 );
not ( n22673 , n21463 );
and ( n22674 , n22667 , n21430 );
not ( n22675 , n21459 );
nor ( n22676 , n22674 , n22675 );
and ( n22677 , n22673 , n22676 );
nor ( n22678 , n22672 , n22677 );
buf ( n22679 , n21741 );
and ( n22680 , n22678 , n22679 );
not ( n22681 , n22678 );
not ( n22682 , n22679 );
and ( n22683 , n22681 , n22682 );
nor ( n22684 , n22680 , n22683 );
not ( n22685 , n21561 );
buf ( n22686 , n22685 );
not ( n22687 , n22686 );
not ( n22688 , n22687 );
and ( n22689 , n22684 , n22688 );
not ( n22690 , n21635 );
xor ( n22691 , n21573 , n22690 );
or ( n22692 , n22691 , n21745 );
and ( n22693 , n21241 , n21242 );
not ( n22694 , n21241 );
and ( n22695 , n22694 , n21237 );
nor ( n22696 , n22693 , n22695 );
and ( n22697 , n22696 , n21356 );
and ( n22698 , n21751 , RI15b57930_853);
nor ( n22699 , n22697 , n22698 );
nand ( n22700 , n22692 , n22699 );
nor ( n22701 , n22689 , n22700 );
and ( n22702 , n21788 , RI15b56a30_821);
and ( n22703 , n21810 , n21768 );
buf ( n22704 , n21794 );
not ( n22705 , n17530 );
and ( n22706 , n22705 , n21803 );
not ( n22707 , n22705 );
and ( n22708 , n22707 , RI15b56a30_821);
nor ( n22709 , n22706 , n22708 );
and ( n22710 , n22704 , n22709 );
nor ( n22711 , n22702 , n22703 , n22710 );
nand ( n22712 , n22701 , n22711 );
buf ( n22713 , n22712 );
buf ( n22714 , RI15b3ea48_2);
buf ( n22715 , n22714 );
buf ( n22716 , RI15b3e9d0_1);
buf ( n22717 , n22716 );
not ( n22718 , n20526 );
or ( n22719 , n19907 , n22718 );
nor ( n22720 , n22362 , RI15b4a190_393);
and ( n22721 , n19999 , n22720 );
not ( n22722 , RI15b4c008_458);
or ( n22723 , n20642 , n22722 );
not ( n22724 , RI15b4c008_458);
nand ( n22725 , n22724 , RI15b4bf90_457);
or ( n22726 , n20559 , n22725 );
not ( n22727 , RI15b4c008_458);
or ( n22728 , n22727 , RI15b4bf90_457);
nand ( n22729 , n22726 , n22728 );
and ( n22730 , n22729 , n20646 );
and ( n22731 , n20520 , RI15b4a208_394);
and ( n22732 , n20655 , RI15b4b108_426);
nor ( n22733 , n22730 , n22731 , n22732 );
nand ( n22734 , n22723 , n22733 );
nor ( n22735 , n22721 , n22734 );
nand ( n22736 , n22719 , n22735 );
buf ( n22737 , n22736 );
buf ( n22738 , RI15b3e9d0_1);
buf ( n22739 , n22738 );
buf ( n22740 , RI15b3ea48_2);
buf ( n22741 , n22740 );
not ( n22742 , n18372 );
not ( n22743 , n18754 );
or ( n22744 , n22742 , n22743 );
or ( n22745 , n18754 , n18372 );
nand ( n22746 , n22744 , n22745 );
and ( n22747 , n22746 , n19287 );
and ( n22748 , n19364 , n19370 );
nor ( n22749 , n22748 , n19371 );
not ( n22750 , n19390 );
or ( n22751 , n22749 , n22750 );
and ( n22752 , n18367 , n19409 );
nor ( n22753 , n18367 , n19409 );
nor ( n22754 , n22752 , n22753 );
not ( n22755 , n22754 );
not ( n22756 , n19475 );
or ( n22757 , n22755 , n22756 );
or ( n22758 , n19475 , n22754 );
nand ( n22759 , n22757 , n22758 );
not ( n22760 , n19498 );
not ( n22761 , n22760 );
and ( n22762 , n22759 , n22761 );
and ( n22763 , n19513 , RI15b63d98_1272);
nor ( n22764 , n22762 , n22763 );
nand ( n22765 , n22751 , n22764 );
nor ( n22766 , n22747 , n22765 );
and ( n22767 , n19608 , RI15b62e98_1240);
buf ( n22768 , n19617 );
nand ( n22769 , n22768 , RI15b62bc8_1234);
and ( n22770 , n22769 , RI15b62e98_1240);
not ( n22771 , n22769 );
not ( n22772 , RI15b62e98_1240);
and ( n22773 , n22771 , n22772 );
nor ( n22774 , n22770 , n22773 );
not ( n22775 , n19630 );
or ( n22776 , n22774 , n22775 );
not ( n22777 , n22768 );
and ( n22778 , n22777 , RI15b62e98_1240);
not ( n22779 , n22777 );
and ( n22780 , n22779 , n22772 );
nor ( n22781 , n22778 , n22780 );
not ( n22782 , n19645 );
or ( n22783 , n22781 , n22782 );
nand ( n22784 , n22776 , n22783 );
nor ( n22785 , n22767 , n22784 );
nand ( n22786 , n22766 , n22785 );
buf ( n22787 , n22786 );
buf ( n22788 , RI15b3ea48_2);
buf ( n22789 , n22788 );
nor ( n22790 , RI15b575e8_846 , RI15b57660_847);
not ( n22791 , RI15b576d8_848);
nand ( n22792 , n22790 , n22791 );
nand ( n22793 , n22792 , RI15b58470_877);
not ( n22794 , n22793 );
not ( n22795 , RI15b57750_849);
and ( n22796 , n22794 , n22795 );
and ( n22797 , n22793 , RI15b57750_849);
nor ( n22798 , n22796 , n22797 );
not ( n22799 , n22798 );
nor ( n22800 , RI15b575e8_846 , RI15b57660_847);
not ( n22801 , n22800 );
nand ( n22802 , n22801 , RI15b58470_877);
not ( n22803 , n22802 );
not ( n22804 , RI15b576d8_848);
and ( n22805 , n22803 , n22804 );
and ( n22806 , n22802 , RI15b576d8_848);
nor ( n22807 , n22805 , n22806 );
or ( n22808 , n22799 , n22807 );
nand ( n22809 , n22799 , n22807 );
nand ( n22810 , n22808 , n22809 );
not ( n22811 , n22810 );
nor ( n22812 , RI15b57b10_857 , RI15b57930_853 , RI15b579a8_854);
nor ( n22813 , RI15b57a20_855 , RI15b57a98_856);
nor ( n22814 , RI15b57b88_858 , RI15b57c00_859);
nand ( n22815 , n22812 , n22813 , n22814 );
nor ( n22816 , RI15b578b8_852 , RI15b57c78_860 , RI15b57cf0_861);
nor ( n22817 , RI15b57660_847 , RI15b576d8_848);
buf ( n22818 , n22817 );
nor ( n22819 , RI15b57750_849 , RI15b577c8_850);
not ( n22820 , n22819 );
not ( n22821 , n22820 );
nor ( n22822 , RI15b575e8_846 , RI15b57840_851);
nand ( n22823 , n22816 , n22818 , n22821 , n22822 );
nor ( n22824 , n22815 , n22823 );
nor ( n22825 , RI15b57d68_862 , RI15b57de0_863);
nand ( n22826 , n22824 , n22825 );
not ( n22827 , n22826 );
nor ( n22828 , RI15b57e58_864 , RI15b57ed0_865);
nand ( n22829 , n22827 , n22828 );
not ( n22830 , n22829 );
nand ( n22831 , n22614 , n22615 );
nor ( n22832 , n22831 , RI15b58038_868);
nand ( n22833 , n22830 , n22832 );
not ( n22834 , n22833 );
not ( n22835 , RI15b580b0_869);
not ( n22836 , RI15b58128_870);
and ( n22837 , n22835 , n22836 );
not ( n22838 , RI15b581a0_871);
not ( n22839 , RI15b58218_872);
nand ( n22840 , n22837 , n22838 , n22839 );
nor ( n22841 , n22840 , RI15b58290_873);
and ( n22842 , n22841 , n22622 );
nand ( n22843 , n22834 , n22842 , n22623 );
nand ( n379040 , n22843 , RI15b58470_877);
and ( n379041 , n379040 , RI15b583f8_876);
not ( n379042 , n379040 );
not ( n379043 , RI15b583f8_876);
and ( n379044 , n379042 , n379043 );
nor ( n379045 , n379041 , n379044 );
buf ( n379046 , n22843 );
nand ( n379047 , n379045 , n379046 );
not ( n379048 , n379047 );
not ( n379049 , n379048 );
nand ( n379050 , n22819 , n22817 , n22822 );
not ( n379051 , n379050 );
buf ( n379052 , n379051 );
nor ( n379053 , RI15b578b8_852 , RI15b57930_853);
nand ( n379054 , n379052 , n379053 );
not ( n379055 , n379054 );
buf ( n379056 , n22813 );
buf ( n379057 , n379056 );
and ( n379058 , n379057 , RI15b57b10_857);
nand ( n379059 , n379055 , n379058 , n21930 );
or ( n379060 , n22605 , n379057 );
nand ( n379061 , n379050 , RI15b58470_877);
buf ( n379062 , n379061 );
not ( n379063 , n21930 );
not ( n379064 , n379053 );
or ( n379065 , n379063 , n379064 );
nand ( n379066 , n379065 , RI15b58470_877);
nand ( n379067 , n379060 , n379062 , n379066 );
nand ( n379068 , n379067 , n21934 );
or ( n379069 , n21934 , RI15b58470_877);
nand ( n379070 , n379059 , n379068 , n379069 );
not ( n379071 , n379070 );
nand ( n379072 , n22798 , n22807 );
nor ( n379073 , RI15b575e8_846 , RI15b57750_849);
not ( n379074 , n379073 );
not ( n379075 , n22817 );
or ( n379076 , n379074 , n379075 );
nand ( n379077 , n379076 , RI15b58470_877);
not ( n379078 , RI15b577c8_850);
and ( n379079 , n379077 , n379078 );
not ( n379080 , n379077 );
and ( n379081 , n379080 , RI15b577c8_850);
nor ( n379082 , n379079 , n379081 );
nor ( n379083 , n379072 , n379082 );
not ( n379084 , n379061 );
not ( n379085 , RI15b578b8_852);
and ( n379086 , n379084 , n379085 );
not ( n379087 , RI15b578b8_852);
not ( n379088 , n379051 );
or ( n379089 , n379087 , n379088 );
not ( n379090 , RI15b58470_877);
nand ( n379091 , n379090 , RI15b578b8_852);
nand ( n379092 , n379089 , n379091 );
nor ( n379093 , n379086 , n379092 );
not ( n379094 , RI15b57840_851);
nor ( n379095 , n22792 , n22820 );
not ( n379096 , n379095 );
or ( n379097 , n379094 , n379096 );
not ( n379098 , RI15b58470_877);
nand ( n379099 , n379098 , RI15b57840_851);
nand ( n379100 , n379097 , n379099 );
not ( n379101 , n22792 );
and ( n379102 , n379101 , n22821 );
not ( n379103 , RI15b57840_851);
nand ( n379104 , n379103 , RI15b58470_877);
nor ( n379105 , n379102 , n379104 );
nor ( n379106 , n379100 , n379105 );
nand ( n379107 , n379093 , n379106 );
not ( n379108 , RI15b578b8_852);
nand ( n379109 , n379051 , n379108 );
not ( n379110 , RI15b57930_853);
nor ( n379111 , n379109 , n379110 );
not ( n379112 , n379111 );
not ( n379113 , RI15b58470_877);
nor ( n379114 , n379113 , RI15b57930_853);
nand ( n379115 , n379109 , n379114 );
not ( n379116 , RI15b58470_877);
nand ( n379117 , n379116 , RI15b57930_853);
nand ( n379118 , n379112 , n379115 , n379117 );
nor ( n379119 , n379107 , n379118 );
nand ( n379120 , n379083 , n379119 );
nand ( n379121 , n379055 , RI15b579a8_854);
nor ( n379122 , n22605 , RI15b579a8_854);
nand ( n379123 , n379054 , n379122 );
or ( n379124 , n21930 , RI15b58470_877);
nand ( n379125 , n379121 , n379123 , n379124 );
nor ( n379126 , n379120 , n379125 );
nor ( n379127 , n379054 , RI15b579a8_854);
not ( n379128 , n379127 );
nand ( n379129 , n379128 , RI15b58470_877);
and ( n379130 , RI15b57a20_855 , n379129 );
not ( n379131 , RI15b57a20_855);
nand ( n379132 , n379062 , n379066 );
and ( n379133 , n379131 , n379132 );
nor ( n379134 , n379130 , n379133 );
nand ( n379135 , n379126 , n379134 );
not ( n379136 , RI15b57a20_855);
not ( n379137 , n379136 );
not ( n379138 , n379127 );
or ( n379139 , n379137 , n379138 );
nand ( n379140 , n379139 , RI15b58470_877);
not ( n379141 , RI15b57a98_856);
and ( n379142 , n379140 , n379141 );
not ( n379143 , n379140 );
and ( n379144 , n379143 , RI15b57a98_856);
nor ( n379145 , n379142 , n379144 );
nor ( n379146 , n379135 , n379145 );
nand ( n379147 , n379071 , n379146 );
not ( n379148 , n21936 );
buf ( n379149 , n379109 );
buf ( n379150 , n22812 );
nand ( n379151 , n379150 , n379056 );
nor ( n379152 , n379149 , n379151 );
nor ( n379153 , n379152 , n22605 );
not ( n379154 , n379153 );
or ( n379155 , n379148 , n379154 );
not ( n379156 , n379153 );
nand ( n379157 , n379156 , RI15b57b88_858);
nand ( n379158 , n379155 , n379157 );
nor ( n379159 , n379147 , n379158 );
not ( n379160 , n21936 );
not ( n379161 , n379152 );
or ( n379162 , n379160 , n379161 );
nand ( n379163 , n379162 , RI15b58470_877);
and ( n379164 , n379163 , n21937 );
not ( n379165 , n379163 );
and ( n379166 , n379165 , RI15b57c00_859);
nor ( n379167 , n379164 , n379166 );
not ( n379168 , n379167 );
nand ( n379169 , n379159 , n379168 );
not ( n379170 , n379169 );
buf ( n379171 , n22814 );
nand ( n379172 , n379152 , n379171 );
nand ( n379173 , n379172 , RI15b58470_877);
not ( n379174 , n379173 );
not ( n379175 , RI15b57c78_860);
and ( n379176 , n379174 , n379175 );
and ( n379177 , n379173 , RI15b57c78_860);
nor ( n379178 , n379176 , n379177 );
nand ( n379179 , n379170 , n379178 );
or ( n379180 , n379172 , RI15b57c78_860);
nand ( n379181 , n379180 , RI15b58470_877);
and ( n379182 , RI15b57cf0_861 , n379181 );
not ( n379183 , RI15b57cf0_861);
not ( n379184 , RI15b58470_877);
nand ( n379185 , n379171 , n21940 );
not ( n379186 , n379185 );
or ( n379187 , n379184 , n379186 );
not ( n379188 , n379153 );
nand ( n379189 , n379187 , n379188 );
and ( n379190 , n379183 , n379189 );
nor ( n379191 , n379182 , n379190 );
not ( n379192 , n379191 );
nor ( n379193 , n379179 , n379192 );
not ( n379194 , n22824 );
nand ( n379195 , n379194 , RI15b58470_877);
and ( n379196 , n379195 , n21986 );
not ( n379197 , n379195 );
and ( n379198 , n379197 , RI15b57d68_862);
nor ( n379199 , n379196 , n379198 );
not ( n379200 , n379199 );
nand ( n379201 , n379193 , n379200 );
and ( n379202 , n22826 , RI15b58470_877);
and ( n379203 , n379202 , n22610 );
not ( n379204 , n379202 );
and ( n379205 , n379204 , RI15b57e58_864);
nor ( n379206 , n379203 , n379205 );
not ( n379207 , n21986 );
not ( n379208 , n22824 );
or ( n379209 , n379207 , n379208 );
nand ( n379210 , n379209 , RI15b58470_877);
and ( n379211 , RI15b57de0_863 , n379210 );
not ( n379212 , RI15b57de0_863);
not ( n379213 , RI15b58470_877);
not ( n379214 , RI15b57d68_862);
or ( n379215 , n379213 , n379214 );
nand ( n379216 , n379215 , n379195 );
and ( n379217 , n379212 , n379216 );
nor ( n379218 , n379211 , n379217 );
nand ( n379219 , n379206 , n379218 );
and ( n379220 , n21984 , n22610 );
nor ( n379221 , n379220 , n22605 );
nor ( n379222 , n379216 , n379221 );
or ( n379223 , n379222 , RI15b57ed0_865);
not ( n379224 , n22610 );
not ( n379225 , n22827 );
or ( n379226 , n379224 , n379225 );
nand ( n379227 , n379226 , RI15b58470_877);
nand ( n379228 , n379227 , RI15b57ed0_865);
nand ( n379229 , n379223 , n379228 );
nor ( n379230 , n379219 , n379229 );
buf ( n379231 , n22829 );
nand ( n379232 , n379231 , RI15b58470_877);
not ( n379233 , n379232 );
and ( n379234 , n379233 , n22614 );
not ( n379235 , n379233 );
and ( n379236 , n379235 , RI15b57f48_866);
nor ( n379237 , n379234 , n379236 );
nand ( n379238 , n379230 , n379237 );
not ( n379239 , RI15b57fc0_867);
not ( n379240 , n22614 );
not ( n379241 , n379231 );
not ( n379242 , n379241 );
or ( n379243 , n379240 , n379242 );
nand ( n379244 , n379243 , RI15b58470_877);
not ( n379245 , n379244 );
or ( n379246 , n379239 , n379245 );
or ( n379247 , n379244 , RI15b57fc0_867);
nand ( n379248 , n379246 , n379247 );
nor ( n379249 , n379238 , n379248 );
not ( n379250 , n22831 );
not ( n379251 , n379250 );
not ( n379252 , n379241 );
or ( n379253 , n379251 , n379252 );
nand ( n379254 , n379253 , RI15b58470_877);
and ( n379255 , RI15b58038_868 , n379254 );
not ( n379256 , RI15b58038_868);
not ( n379257 , RI15b58470_877);
not ( n379258 , n22831 );
or ( n379259 , n379257 , n379258 );
nand ( n379260 , n379259 , n379232 );
and ( n379261 , n379256 , n379260 );
nor ( n379262 , n379255 , n379261 );
nand ( n379263 , n379249 , n379262 );
nor ( n379264 , n379201 , n379263 );
nand ( n379265 , n22833 , RI15b58470_877);
buf ( n379266 , n379265 );
not ( n379267 , n379266 );
not ( n379268 , RI15b580b0_869);
and ( n379269 , n379267 , n379268 );
and ( n379270 , n379266 , RI15b580b0_869);
nor ( n379271 , n379269 , n379270 );
buf ( n379272 , n379271 );
nand ( n379273 , n379264 , n379272 );
not ( n379274 , n22833 );
nand ( n379275 , n379274 , n22837 );
nor ( n379276 , n22605 , RI15b581a0_871);
and ( n379277 , n379275 , n379276 );
not ( n379278 , n379275 );
and ( n379279 , n379278 , RI15b581a0_871);
nor ( n379280 , n379277 , n379279 );
nand ( n379281 , n22834 , n22835 );
and ( n379282 , n22836 , RI15b58470_877);
and ( n379283 , n379281 , n379282 );
not ( n379284 , n379281 );
and ( n379285 , n379284 , RI15b58128_870);
nor ( n379286 , n379283 , n379285 );
nand ( n379287 , n379280 , n379286 );
not ( n379288 , n379287 );
not ( n379289 , n379288 );
nor ( n379290 , n379273 , n379289 );
buf ( n379291 , n379290 );
not ( n379292 , n379275 );
nand ( n379293 , n379292 , n22838 );
nor ( n379294 , n22605 , RI15b58218_872);
and ( n379295 , n379293 , n379294 );
not ( n379296 , n379293 );
and ( n379297 , n379296 , RI15b58218_872);
nor ( n379298 , n379295 , n379297 );
buf ( n379299 , n379298 );
buf ( n379300 , n379299 );
buf ( n379301 , n379300 );
nand ( n379302 , n379291 , n379301 );
nor ( n379303 , n379293 , RI15b58218_872);
and ( n379304 , n379303 , RI15b58290_873);
nand ( n379305 , n22840 , RI15b58470_877);
not ( n379306 , n379305 );
not ( n379307 , n379265 );
or ( n379308 , n379306 , n379307 );
not ( n379309 , RI15b58290_873);
nand ( n379310 , n379308 , n379309 );
not ( n379311 , n379310 );
nor ( n379312 , n379304 , n379311 );
nand ( n379313 , n22834 , n22842 );
nand ( n379314 , n379313 , RI15b58470_877);
not ( n379315 , n379314 );
not ( n379316 , RI15b58380_875);
and ( n379317 , n379315 , n379316 );
and ( n379318 , n379314 , RI15b58380_875);
nor ( n379319 , n379317 , n379318 );
nand ( n379320 , n379312 , n379319 );
nor ( n379321 , n22622 , RI15b58290_873);
nand ( n379322 , n379303 , n379321 );
not ( n379323 , n22841 );
not ( n379324 , n379265 );
or ( n379325 , n379323 , n379324 );
nand ( n379326 , n379325 , n22622 );
nand ( n379327 , n22605 , RI15b58308_874);
nand ( n379328 , n379326 , n379327 );
not ( n379329 , n379328 );
nand ( n379330 , n379322 , n379329 );
nor ( n379331 , n379320 , n379330 );
buf ( n379332 , n379331 );
not ( n379333 , n379332 );
nor ( n379334 , n379302 , n379333 );
not ( n379335 , n379334 );
or ( n379336 , n379049 , n379335 );
nand ( n379337 , n379336 , RI15b58470_877);
buf ( n379338 , n379337 );
not ( n379339 , RI15b54870_749);
nand ( n379340 , n379339 , RI15b547f8_748);
or ( n379341 , n379340 , RI15b54780_747);
nor ( n379342 , n379338 , n379341 );
buf ( n379343 , n379342 );
not ( n379344 , n379343 );
or ( n379345 , n22811 , n379344 );
not ( n379346 , n22807 );
not ( n379347 , n379346 );
buf ( n379348 , n379093 );
buf ( n379349 , n379348 );
not ( n379350 , n379349 );
nor ( n379351 , n379070 , n379199 , n379350 );
nand ( n379352 , n379288 , n379298 , n379271 , n379351 );
nor ( n379353 , n379047 , n379352 );
not ( n379354 , n379134 );
not ( n379355 , n379125 );
not ( n379356 , n379118 );
buf ( n379357 , n379106 );
not ( n379358 , n379357 );
nor ( n379359 , n379358 , n22799 );
nand ( n379360 , RI15b575e8_846 , RI15b58470_877);
and ( n379361 , n379360 , RI15b57660_847);
not ( n379362 , n379360 );
not ( n379363 , RI15b57660_847);
and ( n379364 , n379362 , n379363 );
or ( n379365 , n379361 , n379364 );
not ( n379366 , n379365 );
nand ( n379367 , n379366 , n22807 );
not ( n379368 , n379082 );
not ( n379369 , n379368 );
nor ( n379370 , n379367 , n379369 );
nand ( n379371 , n379355 , n379356 , n379359 , n379370 );
nor ( n379372 , n379354 , n379371 );
nand ( n379373 , n379262 , n379372 );
not ( n379374 , n379145 );
nor ( n379375 , n379158 , n379167 );
nand ( n379376 , n379191 , n379374 , n379375 , n379178 );
nor ( n379377 , n379373 , n379376 );
and ( n379378 , n379249 , n379377 );
nand ( n379379 , n379331 , n379353 , n379378 );
and ( n379380 , n379379 , RI15b58470_877);
buf ( n379381 , n379380 );
buf ( n379382 , n379381 );
buf ( n379383 , n379382 );
nand ( n379384 , n379383 , n379365 );
not ( n379385 , n379384 );
or ( n379386 , n379347 , n379385 );
or ( n379387 , n379384 , n379346 );
nand ( n379388 , n379386 , n379387 );
nand ( n379389 , n18094 , RI15b547f8_748);
not ( n379390 , n379389 );
and ( n379391 , n379390 , RI15b54870_749);
and ( n379392 , n379388 , n379391 );
not ( n379393 , n379341 );
and ( n379394 , n379393 , n22605 );
and ( n379395 , n379394 , RI15b57750_849);
buf ( n379396 , n379390 );
not ( n379397 , n379396 );
buf ( n379398 , n379397 );
and ( n379399 , n379398 , RI15b51558_640);
nor ( n379400 , n379392 , n379395 , n379399 );
nand ( n379401 , n379345 , n379400 );
buf ( n379402 , n379401 );
buf ( n379403 , RI15b3e9d0_1);
buf ( n379404 , n379403 );
nor ( n379405 , RI15b63a50_1265 , RI15b63ac8_1266);
not ( n379406 , n379405 );
nand ( n379407 , n379406 , RI15b648d8_1296);
not ( n379408 , n379407 );
not ( n379409 , RI15b63b40_1267);
and ( n379410 , n379408 , n379409 );
and ( n379411 , n379407 , RI15b63b40_1267);
nor ( n379412 , n379410 , n379411 );
not ( n379413 , n379412 );
not ( n379414 , n379413 );
not ( n379415 , RI15b64860_1295);
nor ( n379416 , RI15b63a50_1265 , RI15b63ac8_1266);
nor ( n379417 , RI15b63c30_1269 , RI15b63ca8_1270);
nor ( n379418 , RI15b63b40_1267 , RI15b63bb8_1268);
nand ( n379419 , n379416 , n379417 , n379418 );
not ( n379420 , n379419 );
nor ( n379421 , RI15b63e10_1273 , RI15b63e88_1274);
not ( n379422 , RI15b63f00_1275);
and ( n379423 , n379421 , n379422 );
nor ( n379424 , RI15b63d20_1271 , RI15b63d98_1272);
nor ( n379425 , RI15b63f78_1276 , RI15b63ff0_1277);
not ( n379426 , RI15b64068_1278);
nand ( n379427 , n379424 , n379425 , n379426 );
not ( n379428 , n379427 );
nand ( n379429 , n379420 , n379423 , n379428 );
nor ( n379430 , n379429 , RI15b640e0_1279);
not ( n379431 , RI15b64158_1280);
and ( n379432 , n379430 , n379431 );
nor ( n379433 , RI15b641d0_1281 , RI15b64248_1282);
nand ( n379434 , n379432 , n379433 );
not ( n379435 , n379434 );
not ( n379436 , RI15b642c0_1283);
not ( n379437 , RI15b64338_1284);
and ( n379438 , n379436 , n379437 );
not ( n379439 , RI15b643b0_1285);
not ( n379440 , RI15b64428_1286);
and ( n379441 , n379439 , n379440 );
nor ( n379442 , RI15b644a0_1287 , RI15b64518_1288);
nand ( n379443 , n379435 , n379438 , n379441 , n379442 );
not ( n379444 , n379443 );
not ( n379445 , RI15b64590_1289);
not ( n379446 , RI15b64608_1290);
and ( n379447 , n379445 , n379446 );
not ( n379448 , RI15b64680_1291);
and ( n379449 , n379447 , n379448 );
nor ( n379450 , RI15b646f8_1292 , RI15b64770_1293);
not ( n379451 , RI15b647e8_1294);
and ( n379452 , n379444 , n379449 , n379450 , n379451 );
not ( n379453 , n379452 );
or ( n379454 , n379415 , n379453 );
or ( n379455 , n379452 , RI15b64860_1295);
nand ( n379456 , n379454 , n379455 );
nand ( n379457 , n379444 , n379449 , n379450 );
nand ( n379458 , n379457 , RI15b648d8_1296);
and ( n379459 , n379458 , n379451 );
not ( n379460 , n379458 );
and ( n379461 , n379460 , RI15b647e8_1294);
nor ( n379462 , n379459 , n379461 );
nor ( n379463 , n379456 , n379462 );
nor ( n379464 , RI15b63ac8_1266 , RI15b63b40_1267);
nor ( n379465 , RI15b63a50_1265 , RI15b63bb8_1268);
nand ( n379466 , n379464 , n379465 );
not ( n379467 , n379466 );
nand ( n379468 , n379417 , n379424 );
not ( n379469 , n379468 );
nand ( n379470 , n379467 , n379469 );
not ( n379471 , n379470 );
buf ( n379472 , n379421 );
nand ( n379473 , n379471 , n379472 );
not ( n379474 , RI15b63f00_1275);
and ( n379475 , n379474 , RI15b648d8_1296);
nand ( n379476 , n379473 , n379475 );
nand ( n379477 , n379466 , RI15b648d8_1296);
not ( n379478 , n379477 );
not ( n379479 , RI15b63c30_1269);
and ( n379480 , n379478 , n379479 );
not ( n379481 , n379478 );
and ( n379482 , n379481 , RI15b63c30_1269);
nor ( n379483 , n379480 , n379482 );
not ( n379484 , RI15b63d20_1271);
not ( n379485 , n379466 );
not ( n379486 , n379485 );
buf ( n379487 , n379417 );
not ( n379488 , n379487 );
nor ( n379489 , n379486 , n379488 );
not ( n379490 , n379489 );
or ( n379491 , n379484 , n379490 );
not ( n379492 , RI15b63d20_1271);
or ( n379493 , n379492 , RI15b648d8_1296);
nand ( n379494 , n379491 , n379493 );
nand ( n379495 , n379419 , RI15b648d8_1296);
nor ( n379496 , n379495 , RI15b63d20_1271);
nor ( n379497 , n379494 , n379496 );
not ( n379498 , RI15b63b40_1267);
not ( n379499 , n379498 );
not ( n379500 , n379405 );
or ( n379501 , n379499 , n379500 );
nand ( n379502 , n379501 , RI15b648d8_1296);
not ( n379503 , n379502 );
not ( n379504 , RI15b63bb8_1268);
and ( n379505 , n379503 , n379504 );
and ( n379506 , n379502 , RI15b63bb8_1268);
nor ( n379507 , n379505 , n379506 );
and ( n379508 , n379476 , n379483 , n379497 , n379507 );
not ( n379509 , RI15b63f00_1275);
nor ( n379510 , n379473 , n379509 );
not ( n379511 , RI15b63f00_1275);
nor ( n379512 , n379511 , RI15b648d8_1296);
nor ( n379513 , n379510 , n379512 );
nand ( n379514 , n379470 , RI15b648d8_1296);
not ( n379515 , n379514 );
not ( n379516 , RI15b63e10_1273);
and ( n379517 , n379515 , n379516 );
not ( n379518 , RI15b63e10_1273);
not ( n379519 , n379470 );
not ( n379520 , n379519 );
or ( n379521 , n379518 , n379520 );
not ( n379522 , RI15b648d8_1296);
nand ( n379523 , n379522 , RI15b63e10_1273);
nand ( n379524 , n379521 , n379523 );
nor ( n379525 , n379517 , n379524 );
nand ( n379526 , RI15b63d20_1271 , RI15b648d8_1296);
not ( n379527 , n379526 );
not ( n379528 , n379495 );
or ( n379529 , n379527 , n379528 );
not ( n379530 , RI15b63d98_1272);
nand ( n379531 , n379529 , n379530 );
nor ( n379532 , n379530 , RI15b63d20_1271);
nand ( n379533 , n379485 , n379487 , n379532 );
not ( n379534 , RI15b648d8_1296);
nand ( n379535 , n379534 , RI15b63d98_1272);
nand ( n379536 , n379531 , n379533 , n379535 );
not ( n379537 , n379536 );
nand ( n379538 , RI15b63c30_1269 , RI15b648d8_1296);
not ( n379539 , n379538 );
not ( n379540 , n379477 );
or ( n379541 , n379539 , n379540 );
not ( n379542 , RI15b63ca8_1270);
nand ( n379543 , n379541 , n379542 );
not ( n379544 , RI15b63ca8_1270);
nor ( n379545 , n379544 , RI15b63c30_1269);
and ( n379546 , n379485 , n379545 );
not ( n379547 , RI15b63ca8_1270);
nor ( n379548 , n379547 , RI15b648d8_1296);
nor ( n379549 , n379546 , n379548 );
nand ( n379550 , n379543 , n379549 );
not ( n379551 , n379550 );
and ( n379552 , n379513 , n379525 , n379537 , n379551 );
not ( n379553 , n379470 );
not ( n379554 , RI15b63e10_1273);
nand ( n379555 , n379553 , n379554 );
not ( n379556 , RI15b63e88_1274);
or ( n379557 , n379555 , n379556 );
or ( n379558 , n379556 , RI15b648d8_1296);
nand ( n379559 , n379557 , n379558 );
buf ( n379560 , n379553 );
and ( n379561 , n379560 , n379554 );
nand ( n379562 , n379556 , RI15b648d8_1296);
nor ( n379563 , n379561 , n379562 );
nor ( n379564 , n379559 , n379563 );
nand ( n379565 , n379508 , n379552 , n379564 );
nor ( n379566 , n379565 , n379413 );
not ( n379567 , RI15b648d8_1296);
not ( n379568 , n379423 );
not ( n379569 , n379568 );
or ( n379570 , n379567 , n379569 );
buf ( n379571 , n379514 );
nand ( n379572 , n379570 , n379571 );
not ( n379573 , RI15b63f78_1276);
and ( n379574 , n379572 , n379573 );
nor ( n379575 , n379573 , RI15b63f00_1275);
not ( n379576 , n379575 );
buf ( n379577 , n379472 );
nand ( n379578 , n379553 , n379577 );
not ( n379579 , n379578 );
not ( n379580 , n379579 );
or ( n379581 , n379576 , n379580 );
or ( n379582 , n379573 , RI15b648d8_1296);
nand ( n379583 , n379581 , n379582 );
nor ( n379584 , n379574 , n379583 );
nand ( n379585 , n379566 , n379584 );
not ( n379586 , RI15b63f00_1275);
nand ( n379587 , n379586 , n379573 );
nor ( n379588 , n379578 , n379587 );
not ( n379589 , RI15b648d8_1296);
nor ( n379590 , n379588 , n379589 );
not ( n379591 , RI15b63ff0_1277);
and ( n379592 , n379590 , n379591 );
not ( n379593 , n379590 );
and ( n379594 , n379593 , RI15b63ff0_1277);
nor ( n379595 , n379592 , n379594 );
not ( n379596 , n379595 );
nor ( n379597 , n379585 , n379596 );
buf ( n379598 , n379579 );
not ( n379599 , n379587 );
nand ( n379600 , n379598 , n379599 , n379591 , RI15b64068_1278);
not ( n379601 , n379591 );
not ( n379602 , n379588 );
or ( n379603 , n379601 , n379602 );
not ( n379604 , RI15b64068_1278);
and ( n379605 , n379604 , RI15b648d8_1296);
nand ( n379606 , n379603 , n379605 );
not ( n379607 , RI15b64068_1278);
or ( n379608 , n379607 , RI15b648d8_1296);
nand ( n379609 , n379600 , n379606 , n379608 );
not ( n379610 , n379429 );
and ( n379611 , n379610 , RI15b640e0_1279);
not ( n379612 , RI15b640e0_1279);
nor ( n379613 , n379612 , RI15b648d8_1296);
nor ( n379614 , n379611 , n379613 );
nand ( n379615 , n379429 , n379612 , RI15b648d8_1296);
nand ( n379616 , n379614 , n379615 );
nor ( n379617 , n379609 , n379616 );
buf ( n379618 , n379617 );
and ( n379619 , n379597 , n379618 );
not ( n379620 , RI15b64158_1280);
buf ( n379621 , n379430 );
not ( n379622 , n379621 );
or ( n379623 , n379620 , n379622 );
or ( n379624 , n379431 , RI15b648d8_1296);
nand ( n379625 , n379623 , n379624 );
nor ( n379626 , n379621 , n379589 , RI15b64158_1280);
nor ( n379627 , n379625 , n379626 );
nand ( n379628 , n379619 , n379627 );
not ( n379629 , n379432 );
nand ( n379630 , n379629 , RI15b648d8_1296);
not ( n379631 , n379630 );
not ( n379632 , RI15b641d0_1281);
and ( n379633 , n379631 , n379632 );
not ( n379634 , n379631 );
and ( n379635 , n379634 , RI15b641d0_1281);
nor ( n379636 , n379633 , n379635 );
not ( n379637 , n379636 );
nor ( n379638 , n379628 , n379637 );
not ( n379639 , n379434 );
nand ( n379640 , n379639 , n379438 , n379441 );
nand ( n379641 , n379640 , RI15b648d8_1296);
and ( n379642 , RI15b644a0_1287 , n379641 );
not ( n379643 , RI15b644a0_1287);
not ( n379644 , RI15b648d8_1296);
not ( n379645 , n379441 );
not ( n379646 , n379645 );
or ( n379647 , n379644 , n379646 );
not ( n379648 , n379438 );
not ( n379649 , n379639 );
or ( n379650 , n379648 , n379649 );
nand ( n379651 , n379650 , RI15b648d8_1296);
nand ( n379652 , n379647 , n379651 );
and ( n379653 , n379643 , n379652 );
nor ( n379654 , n379642 , n379653 );
nor ( n379655 , n379589 , RI15b64248_1282);
not ( n379656 , n379655 );
not ( n379657 , n379629 );
nand ( n379658 , n379657 , n379632 );
not ( n379659 , n379658 );
or ( n379660 , n379656 , n379659 );
and ( n379661 , n379657 , n379632 , RI15b64248_1282);
not ( n379662 , RI15b64248_1282);
nor ( n379663 , n379662 , RI15b648d8_1296);
nor ( n379664 , n379661 , n379663 );
nand ( n379665 , n379660 , n379664 );
not ( n379666 , n379665 );
nand ( n379667 , n379654 , n379666 );
nor ( n379668 , n379651 , RI15b643b0_1285);
nand ( n379669 , n379436 , RI15b648d8_1296);
or ( n379670 , n379639 , n379669 );
nand ( n379671 , n379639 , RI15b642c0_1283);
or ( n379672 , n379436 , RI15b648d8_1296);
nand ( n379673 , n379670 , n379671 , n379672 );
nor ( n379674 , n379668 , n379673 );
not ( n379675 , n379439 );
not ( n379676 , n379438 );
nor ( n379677 , n379434 , n379676 );
not ( n379678 , n379677 );
or ( n379679 , n379675 , n379678 );
nand ( n379680 , n379679 , RI15b648d8_1296);
and ( n379681 , n379680 , RI15b64428_1286);
not ( n379682 , n379680 );
and ( n379683 , n379682 , n379440 );
nor ( n379684 , n379681 , n379683 );
nand ( n379685 , n379651 , RI15b643b0_1285);
not ( n379686 , n379436 );
not ( n379687 , n379433 );
or ( n379688 , n379686 , n379687 );
nand ( n379689 , n379688 , RI15b648d8_1296);
nand ( n379690 , n379630 , n379689 );
and ( n379691 , n379690 , n379437 );
nor ( n379692 , n379437 , RI15b642c0_1283);
not ( n379693 , n379692 );
not ( n379694 , n379639 );
or ( n379695 , n379693 , n379694 );
or ( n379696 , n379437 , RI15b648d8_1296);
nand ( n379697 , n379695 , n379696 );
nor ( n379698 , n379691 , n379697 );
nand ( n379699 , n379674 , n379684 , n379685 , n379698 );
nor ( n379700 , n379667 , n379699 );
nand ( n379701 , n379638 , n379700 );
nor ( n379702 , n379444 , n379589 );
and ( n379703 , n379702 , RI15b64590_1289);
not ( n379704 , n379702 );
and ( n379705 , n379704 , n379445 );
nor ( n379706 , n379703 , n379705 );
not ( n379707 , n379706 );
not ( n379708 , RI15b644a0_1287);
nor ( n379709 , n379589 , n379708 );
or ( n379710 , n379652 , n379709 );
not ( n379711 , RI15b64518_1288);
nand ( n379712 , n379710 , n379711 );
nor ( n379713 , n379640 , RI15b644a0_1287);
or ( n379714 , n379713 , n379589 );
nand ( n379715 , n379714 , RI15b64518_1288);
nand ( n379716 , n379712 , n379715 );
not ( n379717 , n379716 );
nand ( n379718 , n379707 , n379717 );
nor ( n379719 , n379701 , n379718 );
not ( n379720 , RI15b646f8_1292);
not ( n379721 , n379720 );
not ( n379722 , n379449 );
nor ( n379723 , n379443 , n379722 );
not ( n379724 , n379723 );
or ( n379725 , n379721 , n379724 );
nand ( n379726 , n379725 , RI15b648d8_1296);
not ( n379727 , n379726 );
not ( n379728 , RI15b64770_1293);
and ( n379729 , n379727 , n379728 );
and ( n379730 , n379726 , RI15b64770_1293);
nor ( n379731 , n379729 , n379730 );
not ( n379732 , n379449 );
not ( n379733 , n379444 );
or ( n379734 , n379732 , n379733 );
nand ( n379735 , n379734 , RI15b648d8_1296);
and ( n379736 , n379735 , RI15b646f8_1292);
not ( n379737 , n379735 );
and ( n379738 , n379737 , n379720 );
nor ( n379739 , n379736 , n379738 );
nand ( n379740 , n379731 , n379739 );
not ( n379741 , RI15b648d8_1296);
not ( n379742 , n379447 );
not ( n379743 , n379742 );
or ( n379744 , n379741 , n379743 );
nand ( n379745 , n379443 , RI15b648d8_1296);
nand ( n379746 , n379744 , n379745 );
and ( n379747 , n379746 , n379448 );
not ( n379748 , n379447 );
not ( n379749 , n379444 );
or ( n379750 , n379748 , n379749 );
nand ( n379751 , n379750 , RI15b648d8_1296);
nand ( n379752 , n379751 , RI15b64680_1291);
not ( n379753 , n379752 );
nor ( n379754 , n379747 , n379753 );
not ( n379755 , RI15b648d8_1296);
not ( n379756 , RI15b64590_1289);
or ( n379757 , n379755 , n379756 );
nand ( n379758 , n379757 , n379745 );
and ( n379759 , n379758 , n379446 );
not ( n379760 , n379445 );
not ( n379761 , n379444 );
or ( n379762 , n379760 , n379761 );
nand ( n379763 , n379762 , RI15b648d8_1296);
nand ( n379764 , n379763 , RI15b64608_1290);
not ( n379765 , n379764 );
nor ( n379766 , n379759 , n379765 );
nand ( n379767 , n379754 , n379766 );
nor ( n379768 , n379740 , n379767 );
nand ( n379769 , n379463 , n379719 , n379768 );
buf ( n379770 , n379452 );
not ( n379771 , RI15b64860_1295);
nand ( n379772 , n379770 , n379771 );
not ( n379773 , n379772 );
and ( n379774 , n379769 , n379773 );
not ( n379775 , n379769 );
and ( n379776 , n379775 , n379772 );
nor ( n379777 , n379774 , n379776 );
nand ( n379778 , n379777 , RI15b648d8_1296);
not ( n379779 , n379778 );
and ( n379780 , n379779 , n22440 );
not ( n379781 , n379780 );
or ( n379782 , n379414 , n379781 );
and ( n379783 , n22440 , n379589 );
and ( n379784 , n379783 , RI15b63b40_1267);
and ( n379785 , n22437 , RI15b60cd8_1168);
nand ( n379786 , RI15b63a50_1265 , RI15b648d8_1296);
not ( n379787 , RI15b63ac8_1266);
and ( n379788 , n379786 , n379787 );
not ( n379789 , n379786 );
and ( n379790 , n379789 , RI15b63ac8_1266);
or ( n379791 , n379788 , n379790 );
not ( n379792 , n379791 );
and ( n379793 , n379785 , n379792 );
buf ( n379794 , n22438 );
not ( n379795 , n379794 );
buf ( n379796 , n379795 );
and ( n379797 , n379796 , RI15b5d948_1058);
nor ( n379798 , n379784 , n379793 , n379797 );
nand ( n379799 , n379782 , n379798 );
buf ( n379800 , n379799 );
buf ( n379801 , n18226 );
buf ( n379802 , RI15b3e9d0_1);
buf ( n379803 , n379802 );
not ( n379804 , n22160 );
not ( n379805 , n379804 );
not ( n379806 , n379805 );
nand ( n379807 , n379804 , RI15b666d8_1360);
not ( n379808 , n379807 );
not ( n379809 , RI15b65f58_1344);
and ( n379810 , n379808 , n379809 );
and ( n379811 , n379807 , RI15b65f58_1344);
nor ( n379812 , n379810 , n379811 );
not ( n379813 , n379812 );
or ( n379814 , n379806 , n379813 );
nand ( n379815 , n379814 , RI15b666d8_1360);
not ( n379816 , n379815 );
and ( n379817 , n20415 , n20501 );
and ( n379818 , n20489 , n20491 );
nand ( n379819 , n379817 , n379818 );
not ( n379820 , n379819 );
nand ( n379821 , n379816 , n379820 );
not ( n379822 , n379821 );
and ( n379823 , n379822 , RI15b658c8_1330);
nor ( n379824 , n20560 , n20519 );
and ( n379825 , n20510 , n379824 );
and ( n379826 , n379825 , RI15b484f8_332);
nor ( n379827 , n379823 , n379826 );
not ( n379828 , n379818 );
and ( n379829 , n379817 , n379828 );
nand ( n379830 , n20584 , n20579 );
nor ( n379831 , n379829 , n379830 , n20519 );
nand ( n379832 , n20613 , n379831 );
nand ( n379833 , n379832 , RI15b467e8_270);
nand ( n379834 , n379815 , n379820 );
not ( n379835 , n379834 );
not ( n379836 , RI15b658c8_1330);
and ( n379837 , n22268 , n379836 );
not ( n379838 , n22268 );
and ( n379839 , n379838 , RI15b658c8_1330);
nor ( n379840 , n379837 , n379839 );
nand ( n379841 , n379835 , n379840 );
nand ( n379842 , n379827 , n379833 , n379841 );
buf ( n379843 , n379842 );
buf ( n379844 , RI15b3e9d0_1);
buf ( n379845 , n379844 );
buf ( n379846 , n22402 );
buf ( n379847 , RI15b3e9d0_1);
buf ( n379848 , n379847 );
not ( n379849 , n21815 );
not ( n379850 , n379849 );
not ( n379851 , n17507 );
or ( n379852 , n379850 , n379851 );
nand ( n379853 , n379852 , n17565 );
nand ( n379854 , n379853 , n21825 );
not ( n379855 , n17576 );
nor ( n379856 , n379849 , n21825 );
nand ( n379857 , n379855 , n379856 );
buf ( n379858 , n21951 );
and ( n379859 , n21949 , n379858 );
not ( n379860 , n21979 );
nor ( n379861 , n379859 , n379860 );
or ( n379862 , n379861 , n21952 );
or ( n379863 , n379078 , n21946 );
and ( n379864 , n21924 , RI15b577c8_850);
not ( n379865 , n21924 );
and ( n379866 , n379865 , n379078 );
nor ( n379867 , n379864 , n379866 );
and ( n379868 , n18187 , n379867 );
nor ( n379869 , n21982 , n379858 , RI15b559c8_786);
buf ( n379870 , n21977 );
not ( n379871 , n379870 );
buf ( n379872 , n17625 );
buf ( n379873 , n379872 );
buf ( n379874 , n379873 );
buf ( n379875 , n379874 );
buf ( n379876 , n379875 );
buf ( n379877 , n379876 );
buf ( n379878 , n379877 );
buf ( n379879 , n379878 );
buf ( n379880 , n379879 );
not ( n379881 , n379880 );
nor ( n379882 , n379871 , n18203 , n379881 );
nor ( n379883 , n379868 , n379869 , n379882 );
nand ( n379884 , n379862 , n379863 , n379883 );
and ( n379885 , n379884 , n18077 );
and ( n379886 , n18177 , RI15b577c8_850);
not ( n379887 , RI15b568c8_818);
or ( n379888 , n18218 , n379887 );
nand ( n379889 , n379888 , n21750 );
nor ( n379890 , n379885 , n379886 , n379889 );
nand ( n379891 , n379854 , n379857 , n379890 );
buf ( n379892 , n379891 );
buf ( n379893 , RI15b3ea48_2);
buf ( n379894 , n379893 );
buf ( n379895 , RI15b3ea48_2);
buf ( n379896 , n379895 );
not ( n379897 , n17576 );
not ( n379898 , n379897 );
and ( n379899 , n17509 , RI15b566e8_814);
not ( n379900 , RI15b56760_815);
not ( n379901 , RI15b567d8_816);
and ( n379902 , n379900 , n379901 );
nor ( n379903 , n379899 , n379902 );
or ( n379904 , n379898 , n379903 );
nor ( n379905 , n17562 , n17506 );
or ( n379906 , n379901 , RI15b56760_815);
nand ( n379907 , n379901 , RI15b56760_815);
nand ( n379908 , n379906 , n379907 );
nand ( n379909 , n379905 , n379908 );
buf ( n379910 , n18080 );
not ( n379911 , n379910 );
not ( n379912 , n18086 );
or ( n379913 , n379911 , n379912 );
nand ( n379914 , n379913 , n18104 );
and ( n379915 , n379914 , RI15b558d8_784);
not ( n379916 , n18151 );
and ( n379917 , n379916 , RI15b576d8_848);
and ( n379918 , n22791 , RI15b57660_847);
and ( n379919 , n379363 , RI15b576d8_848);
nor ( n379920 , n379918 , n379919 );
or ( n379921 , n18189 , n379920 );
not ( n379922 , n379910 );
and ( n379923 , n18198 , n379922 , n18081 );
not ( n379924 , n18204 );
buf ( n379925 , n20831 );
not ( n379926 , n379925 );
not ( n379927 , n379926 );
not ( n379928 , n379927 );
or ( n379929 , n379924 , n379928 );
and ( n379930 , n18177 , RI15b576d8_848);
nor ( n379931 , n17506 , RI15b566e8_814);
not ( n379932 , n379907 );
and ( n379933 , n379931 , n379932 );
and ( n379934 , n18219 , RI15b567d8_816);
nor ( n379935 , n379930 , n379933 , n379934 );
nand ( n379936 , n379929 , n379935 );
nor ( n379937 , n379923 , n379936 );
nand ( n379938 , n379921 , n379937 );
nor ( n379939 , n379915 , n379917 , n379938 );
nand ( n379940 , n379904 , n379909 , n379939 );
buf ( n379941 , n379940 );
buf ( n379942 , n379847 );
buf ( n379943 , n19655 );
not ( n379944 , n17784 );
nand ( n379945 , n18124 , n18118 , n379944 );
not ( n379946 , n379945 );
and ( n379947 , n17993 , n18077 );
nand ( n379948 , n379946 , n379947 );
not ( n379949 , n379948 );
not ( n379950 , n379949 );
nand ( n379951 , RI15b557e8_782 , RI15b55860_783);
nor ( n379952 , n379951 , n18081 );
nand ( n379953 , n379952 , RI15b55950_785);
nor ( n379954 , n379953 , n21952 );
nand ( n379955 , n379954 , RI15b55a40_787);
not ( n379956 , RI15b55ab8_788);
nor ( n379957 , n379955 , n379956 );
and ( n379958 , n379957 , RI15b55b30_789);
nand ( n379959 , n379958 , RI15b55ba8_790);
not ( n379960 , RI15b55c20_791);
nor ( n379961 , n379959 , n379960 );
nand ( n379962 , n379961 , RI15b55c98_792);
not ( n379963 , n379962 );
and ( n379964 , n379963 , RI15b55d10_793);
nand ( n379965 , n379964 , RI15b55d88_794);
nor ( n379966 , n379965 , n21967 );
nand ( n379967 , n379966 , RI15b55e78_796);
not ( n379968 , n379967 );
and ( n379969 , n379968 , RI15b55ef0_797);
nand ( n379970 , n379969 , RI15b55f68_798);
not ( n379971 , n379970 );
nand ( n379972 , n379971 , RI15b55fe0_799);
not ( n379973 , RI15b56058_800);
nor ( n379974 , n379972 , n379973 );
nand ( n379975 , n379974 , RI15b560d0_801 , RI15b56148_802);
not ( n379976 , RI15b561c0_803);
nor ( n379977 , n379975 , n379976 );
nand ( n379978 , n379977 , RI15b56238_804);
nor ( n379979 , n379978 , n22587 );
nand ( n379980 , n379979 , RI15b56328_806);
not ( n379981 , n379980 );
or ( n379982 , n379950 , n379981 );
or ( n379983 , n379945 , n18115 );
not ( n379984 , n18140 );
nand ( n379985 , n379983 , n18122 , n379984 );
nand ( n379986 , n379985 , n21549 );
not ( n379987 , n18112 );
and ( n379988 , n379987 , n379947 );
not ( n379989 , n379988 );
not ( n379990 , n21555 );
buf ( n379991 , n379990 );
or ( n379992 , n379989 , n379991 );
nand ( n379993 , n18140 , n18077 );
nand ( n379994 , n18114 , n18077 );
not ( n379995 , n379994 );
and ( n379996 , n379987 , n379995 );
nor ( n379997 , n379945 , n379994 );
nor ( n379998 , n379996 , n379997 , n18078 );
nand ( n379999 , n379992 , n379993 , n379998 );
or ( n380000 , n379986 , n379999 );
not ( n380001 , n380000 );
nand ( n380002 , n379982 , n380001 );
not ( n380003 , n380002 );
or ( n380004 , n380003 , n22590 );
not ( n380005 , n379980 );
and ( n380006 , n380005 , n379949 , n22590 );
buf ( n380007 , n21556 );
and ( n380008 , n379988 , n380007 );
buf ( n380009 , n380008 );
buf ( n380010 , n380009 );
buf ( n380011 , n380010 );
buf ( n380012 , n380011 );
not ( n380013 , n17657 );
nor ( n380014 , n380013 , RI15b50fb8_628);
buf ( n380015 , n380014 );
buf ( n380016 , n380015 );
buf ( n380017 , n380016 );
and ( n380018 , n380017 , RI15b4d340_499);
buf ( n380019 , n17585 );
not ( n380020 , n380019 );
buf ( n380021 , n380020 );
buf ( n380022 , n380021 );
and ( n380023 , n380022 , RI15b4e240_531);
nor ( n380024 , n380018 , n380023 );
not ( n380025 , RI15b50fb8_628);
nand ( n380026 , n20767 , n380025 );
not ( n380027 , n380026 );
buf ( n380028 , n380027 );
buf ( n380029 , n380028 );
and ( n380030 , n380029 , RI15b4de80_523);
not ( n380031 , n17641 );
nor ( n380032 , n380031 , RI15b50fb8_628);
buf ( n380033 , n380032 );
buf ( n380034 , n380033 );
and ( n380035 , n380034 , RI15b4d700_507);
nor ( n380036 , n17685 , RI15b50fb8_628);
buf ( n380037 , n380036 );
buf ( n380038 , n380037 );
and ( n380039 , n380038 , RI15b4e600_539);
nor ( n380040 , n380030 , n380035 , n380039 );
buf ( n380041 , n17596 );
buf ( n380042 , n380041 );
buf ( n380043 , n380042 );
and ( n380044 , n380043 , RI15b4e9c0_547);
buf ( n380045 , n17687 );
buf ( n380046 , n380045 );
buf ( n380047 , n380046 );
and ( n380048 , n380047 , RI15b4c800_475);
nor ( n380049 , n380044 , n380048 );
buf ( n380050 , n17691 );
buf ( n380051 , n380050 );
buf ( n380052 , n380051 );
and ( n380053 , n380052 , RI15b4ed80_555);
and ( n380054 , n379874 , RI15b4cf80_491);
nor ( n380055 , n380053 , n380054 );
and ( n380056 , n380024 , n380040 , n380049 , n380055 );
buf ( n380057 , n17675 );
buf ( n380058 , n380057 );
buf ( n380059 , n380058 );
and ( n380060 , n380059 , RI15b4cbc0_483);
not ( n380061 , n17681 );
and ( n380062 , n380061 , RI15b4f140_563);
buf ( n380063 , n17672 );
buf ( n380064 , n380063 );
buf ( n380065 , n380064 );
and ( n380066 , n380065 , RI15b4c440_467);
nor ( n380067 , n380060 , n380062 , n380066 );
nor ( n380068 , n17605 , RI15b50fb8_628);
buf ( n380069 , n380068 );
buf ( n380070 , n380069 );
buf ( n380071 , n380070 );
and ( n380072 , n380071 , RI15b4dac0_515);
buf ( n380073 , n17617 );
buf ( n380074 , n380073 );
buf ( n380075 , n380074 );
and ( n380076 , n380075 , RI15b4fc80_587);
nor ( n380077 , n380072 , n380076 );
buf ( n380078 , n17607 );
buf ( n380079 , n380078 );
buf ( n380080 , n380079 );
and ( n380081 , n380080 , RI15b4f8c0_579);
buf ( n380082 , n17638 );
buf ( n380083 , n380082 );
buf ( n380084 , n380083 );
and ( n380085 , n380084 , RI15b4f500_571);
nor ( n380086 , n380081 , n380085 );
nand ( n380087 , n380056 , n380067 , n380077 , n380086 );
not ( n380088 , n380087 );
not ( n380089 , RI15b50fb8_628);
or ( n380090 , n20731 , RI15b50f40_627);
not ( n380091 , n17614 );
nand ( n380092 , n380090 , n380091 );
not ( n380093 , n380092 );
or ( n380094 , n380089 , n380093 );
not ( n380095 , n17672 );
nand ( n380096 , n380094 , n380095 );
buf ( n380097 , n20752 );
buf ( n380098 , n380097 );
and ( n380099 , n380096 , n380098 );
and ( n380100 , n380099 , RI15b4f398_568);
not ( n380101 , RI15b50fb8_628);
nand ( n380102 , n380097 , n380101 , RI15b50f40_627);
not ( n380103 , RI15b4e498_536);
or ( n380104 , n380102 , n380103 );
and ( n380105 , n380041 , RI15b4e858_544);
and ( n380106 , n380057 , RI15b4ca58_480);
nor ( n380107 , n380105 , n380106 );
and ( n380108 , n380050 , RI15b4ec18_552);
and ( n380109 , n17625 , RI15b4ce18_488);
nor ( n380110 , n380108 , n380109 );
nand ( n380111 , n380104 , n380107 , n380110 );
not ( n380112 , RI15b4c698_472);
and ( n380113 , RI15b50f40_627 , RI15b50fb8_628);
nand ( n380114 , n380097 , n380113 );
not ( n380115 , n380114 );
not ( n380116 , n380115 );
or ( n380117 , n380112 , n380116 );
and ( n380118 , n380061 , RI15b4efd8_560);
and ( n380119 , n380020 , RI15b4e0d8_528);
nor ( n380120 , n380118 , n380119 );
nand ( n380121 , n380117 , n380120 );
nor ( n380122 , n380100 , n380111 , n380121 );
and ( n380123 , n380096 , n20732 );
and ( n380124 , n380123 , RI15b4f758_576);
and ( n380125 , n380096 , n17622 );
and ( n380126 , n380125 , RI15b4fb18_584);
nor ( n380127 , n380124 , n380126 );
and ( n380128 , n380096 , n20741 );
and ( n380129 , n380128 , RI15b4fed8_592);
not ( n380130 , RI15b50fb8_628);
not ( n380131 , RI15b50f40_627);
nand ( n380132 , n380097 , n380130 , n380131 );
or ( n380133 , n380132 , n20771 );
and ( n380134 , n380068 , RI15b4d958_512);
and ( n380135 , n380027 , RI15b4dd18_520);
and ( n380136 , n380014 , RI15b4d1d8_496);
nor ( n380137 , n380134 , n380135 , n380136 );
nand ( n380138 , n380133 , n380137 );
nor ( n380139 , n380129 , n380138 );
nand ( n380140 , n380122 , n380127 , n380139 );
and ( n380141 , n380015 , RI15b4d250_497);
not ( n380142 , n380019 );
and ( n380143 , n380142 , RI15b4e150_529);
nor ( n380144 , n380141 , n380143 );
and ( n380145 , n380027 , RI15b4dd90_521);
and ( n380146 , n380032 , RI15b4d610_505);
and ( n380147 , n380036 , RI15b4e510_537);
nor ( n380148 , n380145 , n380146 , n380147 );
and ( n380149 , n380050 , RI15b4ec90_553);
and ( n380150 , n379872 , RI15b4ce90_489);
nor ( n380151 , n380149 , n380150 );
and ( n380152 , n380041 , RI15b4e8d0_545);
and ( n380153 , n380045 , RI15b4c710_473);
nor ( n380154 , n380152 , n380153 );
and ( n380155 , n380144 , n380148 , n380151 , n380154 );
and ( n380156 , n380061 , RI15b4f050_561);
and ( n380157 , n380063 , RI15b4c350_465);
and ( n380158 , n380057 , RI15b4cad0_481);
nor ( n380159 , n380156 , n380157 , n380158 );
and ( n380160 , n380069 , RI15b4d9d0_513);
and ( n380161 , n380073 , RI15b4fb90_585);
nor ( n380162 , n380160 , n380161 );
and ( n380163 , n380078 , RI15b4f7d0_577);
and ( n380164 , n380082 , RI15b4f410_569);
nor ( n380165 , n380163 , n380164 );
nand ( n380166 , n380155 , n380159 , n380162 , n380165 );
and ( n380167 , n380140 , n380166 );
and ( n380168 , n380016 , RI15b4d2c8_498);
and ( n380169 , n380021 , RI15b4e1c8_530);
nor ( n380170 , n380168 , n380169 );
and ( n380171 , n380028 , RI15b4de08_522);
and ( n380172 , n380033 , RI15b4d688_506);
and ( n380173 , n380037 , RI15b4e588_538);
nor ( n380174 , n380171 , n380172 , n380173 );
and ( n380175 , n380042 , RI15b4e948_546);
and ( n380176 , n380046 , RI15b4c788_474);
nor ( n380177 , n380175 , n380176 );
and ( n380178 , n380051 , RI15b4ed08_554);
and ( n380179 , n379873 , RI15b4cf08_490);
nor ( n380180 , n380178 , n380179 );
and ( n380181 , n380170 , n380174 , n380177 , n380180 );
and ( n380182 , n380058 , RI15b4cb48_482);
and ( n380183 , n380061 , RI15b4f0c8_562);
and ( n380184 , n380064 , RI15b4c3c8_466);
nor ( n380185 , n380182 , n380183 , n380184 );
and ( n380186 , n380070 , RI15b4da48_514);
and ( n380187 , n380074 , RI15b4fc08_586);
nor ( n380188 , n380186 , n380187 );
and ( n380189 , n380079 , RI15b4f848_578);
and ( n380190 , n380083 , RI15b4f488_570);
nor ( n380191 , n380189 , n380190 );
nand ( n380192 , n380181 , n380185 , n380188 , n380191 );
nand ( n380193 , n380167 , n380192 );
not ( n380194 , n380193 );
or ( n380195 , n380088 , n380194 );
or ( n380196 , n380193 , n380087 );
nand ( n380197 , n380195 , n380196 );
and ( n380198 , n380012 , n380197 );
nor ( n380199 , n380006 , n380198 );
nand ( n380200 , n380004 , n380199 );
buf ( n380201 , n380200 );
buf ( n380202 , RI15b5e5f0_1085);
buf ( n380203 , RI15b3ea48_2);
buf ( n380204 , n380203 );
buf ( n380205 , n379844 );
not ( n380206 , n19216 );
nand ( n380207 , n380206 , RI15b58650_881);
and ( n380208 , n380207 , n19206 );
not ( n380209 , n380207 );
and ( n380210 , n380209 , RI15b586c8_882);
nor ( n380211 , n380208 , n380210 );
not ( n380212 , n380211 );
not ( n380213 , RI15b58650_881);
not ( n380214 , n19217 );
or ( n380215 , n380213 , n380214 );
or ( n380216 , n19217 , RI15b58650_881);
nand ( n380217 , n380215 , n380216 );
and ( n380218 , n380212 , n380217 );
nand ( n380219 , n380218 , n19272 );
not ( n380220 , n19271 );
not ( n380221 , n380211 );
or ( n380222 , n380220 , n380221 );
not ( n380223 , n380217 );
nand ( n380224 , n380223 , n380211 );
nand ( n380225 , n380222 , n380224 );
not ( n380226 , n380225 );
nand ( n380227 , n380219 , n380226 );
buf ( n380228 , n380227 );
not ( n380229 , n380228 );
buf ( n380230 , n380229 );
not ( n380231 , n380217 );
buf ( n380232 , n19273 );
not ( n380233 , n380232 );
nor ( n380234 , n380231 , n380233 );
and ( n380235 , n380230 , n380234 );
not ( n380236 , n380235 );
buf ( n380237 , n19645 );
buf ( n380238 , n380237 );
not ( n380239 , n380238 );
nor ( n380240 , RI15b5ddf8_1068 , RI15b5de70_1069);
nor ( n380241 , RI15b5dee8_1070 , RI15b5df60_1071);
nor ( n380242 , RI15b5dfd8_1072 , RI15b5e050_1073);
nor ( n380243 , RI15b5e0c8_1074 , RI15b5e140_1075);
nand ( n380244 , n380240 , n380241 , n380242 , n380243 );
nor ( n380245 , RI15b5da38_1060 , RI15b5dab0_1061);
nor ( n380246 , RI15b5db28_1062 , RI15b5dba0_1063);
nor ( n380247 , RI15b5e398_1080 , RI15b5e410_1081);
nor ( n380248 , RI15b5e488_1082 , RI15b5e500_1083);
nand ( n380249 , n380245 , n380246 , n380247 , n380248 );
nor ( n380250 , n380244 , n380249 );
nor ( n380251 , RI15b5dc18_1064 , RI15b5dc90_1065);
nor ( n380252 , RI15b5dd08_1066 , RI15b5dd80_1067);
nor ( n380253 , RI15b5e1b8_1076 , RI15b5e230_1077);
nor ( n380254 , RI15b5e2a8_1078 , RI15b5e320_1079);
nand ( n380255 , n380251 , n380252 , n380253 , n380254 );
nor ( n380256 , RI15b5e578_1084 , RI15b5e5f0_1085);
nor ( n380257 , RI15b5d948_1058 , RI15b5d9c0_1059);
not ( n380258 , RI15b5e668_1086);
nand ( n380259 , n380256 , n380257 , n380258 );
nor ( n380260 , n380255 , n380259 );
nand ( n380261 , n380250 , n380260 );
nand ( n380262 , n380261 , RI15b5e6e0_1087);
buf ( n380263 , n380262 );
buf ( n380264 , n380263 );
buf ( n380265 , n380264 );
not ( n380266 , n380265 );
not ( n380267 , RI15b657d8_1328);
not ( n380268 , n380267 );
and ( n380269 , n380266 , n380268 );
buf ( n380270 , n380262 );
not ( n380271 , n380270 );
not ( n380272 , n380271 );
not ( n380273 , n380272 );
not ( n380274 , n380273 );
and ( n380275 , n380274 , RI15b3eac0_3);
nor ( n380276 , n380269 , n380275 );
not ( n380277 , n380276 );
not ( n380278 , n380277 );
not ( n380279 , n380278 );
buf ( n380280 , n380279 );
not ( n380281 , n380280 );
not ( n380282 , n380281 );
not ( n380283 , n380282 );
not ( n380284 , n380283 );
not ( n380285 , n380284 );
not ( n380286 , n380270 );
and ( n380287 , n380286 , RI15b64ab8_1300);
not ( n380288 , n380270 );
not ( n380289 , RI15b3f7e0_31);
nor ( n380290 , n380288 , n380289 );
nor ( n380291 , n380287 , n380290 );
and ( n380292 , n380271 , RI15b64b30_1301);
not ( n380293 , n380263 );
not ( n380294 , RI15b3f768_30);
nor ( n380295 , n380293 , n380294 );
nor ( n380296 , n380292 , n380295 );
buf ( n380297 , n380270 );
or ( n380298 , n380297 , RI15b64ba8_1302);
not ( n380299 , RI15b3f6f0_29);
nand ( n380300 , n380299 , n380263 );
nand ( n380301 , n380298 , n380300 );
and ( n380302 , n380291 , n380296 , n380301 );
not ( n380303 , n380263 );
and ( n380304 , n380303 , RI15b649c8_1298);
not ( n380305 , n380263 );
not ( n380306 , RI15b3f8d0_33);
nor ( n380307 , n380305 , n380306 );
nor ( n380308 , n380304 , n380307 );
not ( n380309 , n380263 );
not ( n380310 , RI15b64950_1297);
not ( n380311 , n380310 );
and ( n380312 , n380309 , n380311 );
buf ( n380313 , n380270 );
and ( n380314 , n380313 , RI15b3f948_34);
nor ( n380315 , n380312 , n380314 );
not ( n380316 , n380263 );
not ( n380317 , RI15b64a40_1299);
not ( n380318 , n380317 );
and ( n380319 , n380316 , n380318 );
and ( n380320 , n380313 , RI15b3f858_32);
nor ( n380321 , n380319 , n380320 );
and ( n380322 , n380308 , n380315 , n380321 );
not ( n380323 , n380264 );
not ( n380324 , RI15b64c20_1303);
not ( n380325 , n380324 );
and ( n380326 , n380323 , n380325 );
and ( n380327 , n380265 , RI15b3f678_28);
nor ( n380328 , n380326 , n380327 );
nand ( n380329 , n380302 , n380322 , n380328 );
not ( n380330 , n380313 );
not ( n380331 , RI15b64c98_1304);
not ( n380332 , n380331 );
and ( n380333 , n380330 , n380332 );
buf ( n380334 , n380263 );
and ( n380335 , n380334 , RI15b3f600_27);
nor ( n380336 , n380333 , n380335 );
buf ( n380337 , n380336 );
not ( n380338 , n380337 );
nor ( n380339 , n380329 , n380338 );
not ( n380340 , n380271 );
not ( n380341 , n380340 );
not ( n380342 , RI15b64d10_1305);
not ( n380343 , n380342 );
and ( n380344 , n380341 , n380343 );
and ( n380345 , n380272 , RI15b3f588_26);
nor ( n380346 , n380344 , n380345 );
not ( n380347 , n380297 );
not ( n380348 , RI15b64d88_1306);
not ( n380349 , n380348 );
and ( n380350 , n380347 , n380349 );
and ( n380351 , n380334 , RI15b3f510_25);
nor ( n380352 , n380350 , n380351 );
not ( n380353 , n380263 );
not ( n380354 , RI15b64e00_1307);
not ( n380355 , n380354 );
and ( n380356 , n380353 , n380355 );
and ( n380357 , n380297 , RI15b3f498_24);
nor ( n380358 , n380356 , n380357 );
not ( n380359 , n380263 );
not ( n380360 , RI15b64e78_1308);
not ( n380361 , n380360 );
and ( n380362 , n380359 , n380361 );
and ( n380363 , n380297 , RI15b3f420_23);
nor ( n380364 , n380362 , n380363 );
nand ( n380365 , n380346 , n380352 , n380358 , n380364 );
not ( n380366 , n380365 );
and ( n380367 , n380339 , n380366 );
buf ( n380368 , n380263 );
not ( n380369 , n380368 );
not ( n380370 , RI15b64ef0_1309);
not ( n380371 , n380370 );
and ( n380372 , n380369 , n380371 );
and ( n380373 , n380264 , RI15b3f3a8_22);
nor ( n380374 , n380372 , n380373 );
buf ( n380375 , n380374 );
not ( n380376 , n380288 );
not ( n380377 , n380376 );
not ( n380378 , RI15b64f68_1310);
not ( n380379 , n380378 );
and ( n380380 , n380377 , n380379 );
not ( n380381 , n380286 );
and ( n380382 , n380381 , RI15b3f330_21);
nor ( n380383 , n380380 , n380382 );
buf ( n380384 , n380383 );
not ( n380385 , n380297 );
not ( n380386 , RI15b64fe0_1311);
not ( n380387 , n380386 );
and ( n380388 , n380385 , n380387 );
not ( n380389 , n380286 );
and ( n380390 , n380389 , RI15b3f2b8_20);
nor ( n380391 , n380388 , n380390 );
buf ( n380392 , n380391 );
nand ( n380393 , n380367 , n380375 , n380384 , n380392 );
not ( n380394 , n380393 );
not ( n380395 , n380368 );
not ( n380396 , RI15b65058_1312);
not ( n380397 , n380396 );
and ( n380398 , n380395 , n380397 );
and ( n380399 , n380264 , RI15b3f240_19);
nor ( n380400 , n380398 , n380399 );
buf ( n380401 , n380400 );
nand ( n380402 , n380394 , n380401 );
nand ( n380403 , n380402 , n380280 );
not ( n380404 , n380403 );
not ( n380405 , n380286 );
not ( n380406 , n380405 );
not ( n380407 , RI15b650d0_1313);
not ( n380408 , n380407 );
and ( n380409 , n380406 , n380408 );
and ( n380410 , n380272 , RI15b3f1c8_18);
nor ( n380411 , n380409 , n380410 );
buf ( n380412 , n380411 );
not ( n380413 , n380412 );
not ( n380414 , n380413 );
and ( n380415 , n380404 , n380414 );
not ( n380416 , n380412 );
and ( n380417 , n380403 , n380416 );
nor ( n380418 , n380415 , n380417 );
not ( n380419 , n380297 );
not ( n380420 , RI15b65148_1314);
not ( n380421 , n380420 );
and ( n380422 , n380419 , n380421 );
and ( n380423 , n380334 , RI15b3f150_17);
nor ( n380424 , n380422 , n380423 );
not ( n380425 , n380313 );
not ( n380426 , RI15b65328_1318);
not ( n380427 , n380426 );
and ( n380428 , n380425 , n380427 );
and ( n380429 , n380334 , RI15b3ef70_13);
nor ( n380430 , n380428 , n380429 );
and ( n380431 , n380400 , n380411 , n380424 , n380430 );
not ( n380432 , n380297 );
not ( n380433 , RI15b65238_1316);
not ( n380434 , n380433 );
and ( n380435 , n380432 , n380434 );
and ( n380436 , n380272 , RI15b3f060_15);
nor ( n380437 , n380435 , n380436 );
nand ( n380438 , n380391 , n380437 );
not ( n380439 , n380376 );
not ( n380440 , RI15b652b0_1317);
not ( n380441 , n380440 );
and ( n380442 , n380439 , n380441 );
and ( n380443 , n380381 , RI15b3efe8_14);
nor ( n380444 , n380442 , n380443 );
nand ( n380445 , n380383 , n380444 );
nor ( n380446 , n380438 , n380445 );
not ( n380447 , n380297 );
not ( n380448 , RI15b651c0_1315);
not ( n380449 , n380448 );
and ( n380450 , n380447 , n380449 );
and ( n380451 , n380389 , RI15b3f0d8_16);
nor ( n380452 , n380450 , n380451 );
nand ( n380453 , n380374 , n380452 , n380336 );
not ( n380454 , n380453 );
nand ( n380455 , n380366 , n380431 , n380446 , n380454 );
nor ( n380456 , n380455 , n380329 );
buf ( n380457 , n380456 );
and ( n380458 , n380273 , RI15b65490_1321);
not ( n380459 , n380273 );
and ( n380460 , n380459 , RI15b3ee08_10);
nor ( n380461 , n380458 , n380460 );
not ( n380462 , n380265 );
not ( n380463 , RI15b65508_1322);
not ( n380464 , n380463 );
and ( n380465 , n380462 , n380464 );
not ( n380466 , n380273 );
and ( n380467 , n380466 , RI15b3ed90_9);
nor ( n380468 , n380465 , n380467 );
and ( n380469 , n380461 , n380468 );
not ( n380470 , n380273 );
and ( n380471 , n380470 , RI15b3eef8_12);
not ( n380472 , RI15b653a0_1319);
nor ( n380473 , n380265 , n380472 );
nor ( n380474 , n380471 , n380473 );
not ( n380475 , n380265 );
not ( n380476 , RI15b65418_1320);
not ( n380477 , n380476 );
and ( n380478 , n380475 , n380477 );
and ( n380479 , n380274 , RI15b3ee80_11);
nor ( n380480 , n380478 , n380479 );
nand ( n380481 , n380457 , n380469 , n380474 , n380480 );
not ( n380482 , n380481 );
not ( n380483 , n380470 );
buf ( n380484 , n380483 );
not ( n380485 , n380484 );
or ( n380486 , n380485 , RI15b65580_1323 , RI15b655f8_1324);
or ( n380487 , n380484 , RI15b3eca0_7 , RI15b3ed18_8);
nand ( n380488 , n380486 , n380487 );
nand ( n380489 , n380482 , n380488 );
and ( n380490 , n380485 , RI15b3ec28_6);
not ( n380491 , n380485 );
and ( n380492 , n380491 , RI15b65670_1325);
nor ( n380493 , n380490 , n380492 );
nor ( n380494 , n380489 , n380493 );
and ( n380495 , n380456 , n380474 , n380480 );
not ( n380496 , RI15b3ee08_10);
not ( n380497 , RI15b3ed90_9);
nand ( n380498 , n380495 , n380496 , n380497 );
nand ( n380499 , n380495 , n380496 );
nor ( n380500 , n380278 , n380497 );
nand ( n380501 , n380499 , n380500 );
not ( n380502 , n380485 );
buf ( n380503 , n380502 );
buf ( n380504 , n380503 );
not ( n380505 , n380504 );
nand ( n380506 , n380498 , n380501 , n380505 );
nor ( n380507 , n380495 , n380278 );
and ( n380508 , n380507 , n380461 );
not ( n380509 , n380507 );
not ( n380510 , n380461 );
and ( n380511 , n380509 , n380510 );
nor ( n380512 , n380508 , n380511 );
nand ( n380513 , n380506 , n380512 );
nor ( n380514 , n380494 , n380513 );
not ( n380515 , n380493 );
nor ( n380516 , n380489 , n380515 );
nor ( n380517 , n380457 , n380278 );
not ( n380518 , n380517 );
not ( n380519 , n380474 );
and ( n380520 , n380518 , n380519 );
and ( n380521 , n380517 , n380474 );
nor ( n380522 , n380520 , n380521 );
nand ( n380523 , n380457 , n380474 );
and ( n380524 , n380523 , n380480 );
not ( n380525 , n380523 );
not ( n380526 , n380480 );
and ( n380527 , n380525 , n380526 );
nor ( n380528 , n380524 , n380527 );
nand ( n380529 , n380522 , n380528 );
nor ( n380530 , n380516 , n380529 );
nand ( n380531 , n380418 , n380514 , n380530 );
not ( n380532 , n380531 );
or ( n380533 , n380285 , n380532 );
buf ( n380534 , n380485 );
not ( n380535 , n380534 );
and ( n380536 , n380535 , RI15b656e8_1326);
not ( n380537 , n380535 );
and ( n380538 , n380537 , RI15b3ebb0_5);
nor ( n380539 , n380536 , n380538 );
nand ( n380540 , n380282 , n380539 );
nand ( n380541 , n380533 , n380540 );
not ( n380542 , n380541 );
not ( n380543 , n380452 );
buf ( n380544 , n380543 );
not ( n380545 , n380544 );
not ( n380546 , n380393 );
buf ( n380547 , n380401 );
buf ( n380548 , n380424 );
and ( n380549 , n380546 , n380547 , n380412 , n380548 );
not ( n380550 , n380549 );
or ( n380551 , n380545 , n380550 );
not ( n380552 , n380430 );
buf ( n380553 , n380437 );
and ( n380554 , n380552 , n380553 );
buf ( n380555 , n380444 );
not ( n380556 , n380555 );
or ( n380557 , n380556 , n380553 );
or ( n380558 , n380555 , n380543 );
nand ( n380559 , n380557 , n380558 );
and ( n380560 , n380502 , RI15b65760_1327);
and ( n380561 , n380485 , RI15b3eb38_4);
nor ( n380562 , n380560 , n380561 );
nor ( n380563 , n380554 , n380559 , n380562 );
nand ( n380564 , n380551 , n380563 );
nand ( n380565 , n380546 , n380547 , n380412 );
and ( n380566 , n380565 , n380548 );
not ( n380567 , n380565 );
not ( n380568 , n380548 );
and ( n380569 , n380567 , n380568 );
nor ( n380570 , n380566 , n380569 );
not ( n380571 , n380481 );
and ( n380572 , n380483 , RI15b655f8_1324);
buf ( n380573 , n380466 );
and ( n380574 , n380573 , RI15b3eca0_7);
nor ( n380575 , n380572 , n380574 );
nor ( n380576 , n380571 , n380575 );
not ( n380577 , n380576 );
and ( n380578 , n380503 , RI15b65580_1323 , RI15b655f8_1324);
and ( n380579 , n380534 , RI15b3eca0_7 , RI15b3ed18_8);
nor ( n380580 , n380578 , n380579 );
nand ( n380581 , n380577 , n380489 , n380580 );
not ( n380582 , n380581 );
not ( n380583 , RI15b65490_1321);
nand ( n380584 , n380495 , n380583 );
nand ( n380585 , n380584 , n380463 );
not ( n380586 , n380585 );
not ( n380587 , n380279 );
not ( n380588 , n380584 );
or ( n380589 , n380587 , n380588 );
nand ( n380590 , n380589 , RI15b65508_1322);
not ( n380591 , n380590 );
or ( n380592 , n380586 , n380591 );
nand ( n380593 , n380592 , n380504 );
not ( n380594 , n380482 );
and ( n380595 , n380483 , RI15b65580_1323);
and ( n380596 , n380573 , RI15b3ed18_8);
nor ( n380597 , n380595 , n380596 );
not ( n380598 , n380597 );
not ( n380599 , n380598 );
and ( n380600 , n380594 , n380599 );
and ( n380601 , n380482 , n380598 );
nor ( n380602 , n380600 , n380601 );
and ( n380603 , n380597 , n380575 );
not ( n380604 , n380603 );
not ( n380605 , n380482 );
or ( n380606 , n380604 , n380605 );
nand ( n380607 , n380606 , n380493 );
nand ( n380608 , n380593 , n380602 , n380607 );
nor ( n380609 , n380582 , n380608 );
nand ( n380610 , n380570 , n380609 );
or ( n380611 , n380564 , n380610 );
not ( n380612 , n380283 );
nand ( n380613 , n380611 , n380612 );
not ( n380614 , n380549 );
buf ( n380615 , n380552 );
not ( n380616 , n380615 );
nand ( n380617 , n380614 , n380612 , n380616 );
nand ( n380618 , n380542 , n380613 , n380617 );
not ( n380619 , n380618 );
not ( n380620 , n380619 );
buf ( n380621 , n380544 );
not ( n380622 , n380621 );
and ( n380623 , n380614 , n380622 );
nand ( n380624 , n380620 , n380623 );
not ( n380625 , n380544 );
and ( n380626 , n380549 , n380625 );
buf ( n380627 , n380553 );
nand ( n380628 , n380626 , n380627 );
not ( n380629 , n380628 );
buf ( n380630 , n380555 );
nand ( n380631 , n380629 , n380630 );
buf ( n380632 , n380615 );
not ( n380633 , n380632 );
nand ( n380634 , n380618 , n380631 , n380633 );
buf ( n380635 , n380284 );
not ( n380636 , n380635 );
not ( n380637 , n380636 );
not ( n380638 , n380637 );
not ( n380639 , n380631 );
or ( n380640 , n380638 , n380639 );
not ( n380641 , n380633 );
nand ( n380642 , n380640 , n380641 );
buf ( n380643 , n380612 );
nand ( n380644 , n380614 , n380643 );
and ( n380645 , n380644 , n380621 );
buf ( n380646 , n380570 );
buf ( n380647 , n380418 );
nand ( n380648 , n380646 , n380647 );
nor ( n380649 , n380645 , n380648 );
and ( n380650 , n380624 , n380634 , n380642 , n380649 );
not ( n380651 , n380618 );
not ( n380652 , n380651 );
not ( n380653 , n380628 );
not ( n380654 , n380626 );
nand ( n380655 , n380654 , n380643 );
buf ( n380656 , n380627 );
nor ( n380657 , n380655 , n380656 );
nor ( n380658 , n380653 , n380657 );
not ( n380659 , n380658 );
and ( n380660 , n380652 , n380659 );
not ( n380661 , n380655 );
buf ( n380662 , n380656 );
nor ( n380663 , n380661 , n380662 );
and ( n380664 , n380651 , n380663 );
nor ( n380665 , n380660 , n380664 );
and ( n380666 , n380628 , n380630 );
not ( n380667 , n380666 );
not ( n380668 , n380618 );
or ( n380669 , n380667 , n380668 );
not ( n380670 , n380637 );
not ( n380671 , n380628 );
or ( n380672 , n380670 , n380671 );
not ( n380673 , n380630 );
nand ( n380674 , n380672 , n380673 );
nand ( n380675 , n380669 , n380674 );
nor ( n380676 , n380665 , n380675 );
nand ( n380677 , n380650 , n380676 );
not ( n380678 , n380522 );
nor ( n380679 , n380677 , n380678 );
not ( n380680 , n380679 );
or ( n380681 , n380239 , n380680 );
not ( n380682 , n380618 );
not ( n380683 , n380682 );
not ( n380684 , n380683 );
nand ( n380685 , n380684 , n19645 );
buf ( n380686 , n380685 );
nand ( n380687 , n380681 , n380686 );
not ( n380688 , n380528 );
not ( n380689 , n380688 );
not ( n380690 , n380683 );
or ( n380691 , n380689 , n380690 );
buf ( n380692 , n380637 );
not ( n380693 , n380692 );
nand ( n380694 , n380693 , n380526 );
nand ( n380695 , n380691 , n380694 );
and ( n380696 , n380687 , n380695 );
not ( n380697 , n380682 );
and ( n380698 , n380697 , n19645 );
not ( n380699 , n380695 );
nand ( n380700 , n380698 , n380699 );
nor ( n380701 , n380679 , n380700 );
nor ( n380702 , n380696 , n380701 );
not ( n380703 , n380702 );
not ( n380704 , n380703 );
or ( n380705 , n380236 , n380704 );
buf ( n380706 , n380609 );
buf ( n380707 , n380514 );
nand ( n380708 , n380706 , n380707 );
not ( n380709 , n380708 );
not ( n380710 , n380516 );
nand ( n380711 , n380709 , n380710 );
or ( n380712 , n380711 , n380562 );
buf ( n380713 , n380692 );
nand ( n380714 , n380712 , n380713 );
nand ( n380715 , n380714 , n380540 );
not ( n380716 , n380238 );
not ( n380717 , n380716 );
nand ( n380718 , n380715 , n380717 );
not ( n380719 , n380718 );
not ( n380720 , n380227 );
not ( n380721 , n19271 );
buf ( n380722 , n380217 );
not ( n380723 , n380722 );
or ( n380724 , n380721 , n380723 );
nand ( n380725 , n380231 , n19270 );
nand ( n380726 , n380724 , n380725 );
nand ( n380727 , n380720 , n380726 );
or ( n380728 , n19264 , RI15b585d8_880);
nor ( n380729 , n380727 , n380728 );
not ( n380730 , n380728 );
not ( n380731 , n380227 );
or ( n380732 , n380730 , n380731 );
not ( n380733 , n380726 );
nand ( n380734 , n380227 , n380733 );
nand ( n380735 , n380732 , n380734 );
nor ( n380736 , n380729 , n380735 );
not ( n380737 , n380728 );
and ( n380738 , n380726 , n380737 );
not ( n380739 , n380726 );
and ( n380740 , n380739 , n380728 );
nor ( n380741 , n380738 , n380740 );
not ( n380742 , n380741 );
nand ( n380743 , n380736 , n380742 );
or ( n380744 , n380743 , n380728 );
not ( n380745 , n380744 );
and ( n380746 , n380719 , n380745 );
not ( n380747 , n380235 );
not ( n380748 , n19637 );
buf ( n380749 , n380748 );
buf ( n380750 , n380749 );
not ( n380751 , n380750 );
and ( n380752 , n380744 , n380747 , n380751 );
nor ( n380753 , n380752 , n19630 );
buf ( n380754 , n380722 );
or ( n380755 , n380211 , n380754 );
buf ( n380756 , n19217 );
not ( n380757 , n380756 );
not ( n380758 , n380757 );
buf ( n380759 , n380758 );
nor ( n380760 , n380755 , n380759 );
or ( n380761 , n380753 , n380760 );
nand ( n380762 , n380761 , n19595 );
nor ( n380763 , RI15b586c8_882 , RI15b58740_883);
nand ( n380764 , n380763 , n19209 );
buf ( n380765 , n19268 );
buf ( n380766 , n380765 );
not ( n380767 , n380766 );
or ( n380768 , n380764 , n380767 );
nand ( n380769 , n380762 , n380768 );
not ( n380770 , n19595 );
and ( n380771 , n380770 , RI15b5d498_1048);
nor ( n380772 , n380771 , n19599 );
and ( n380773 , n19590 , n19512 );
and ( n380774 , n380772 , n380773 , n19200 , n19581 );
and ( n380775 , n380774 , n19594 );
and ( n380776 , n380769 , n380775 );
or ( n380777 , n380776 , n19031 );
buf ( n380778 , n380337 );
not ( n380779 , n380778 );
buf ( n380780 , n380779 );
buf ( n380781 , n380780 );
not ( n380782 , n380781 );
not ( n380783 , n380768 );
nor ( n380784 , n380760 , n380783 );
or ( n380785 , n380753 , n380784 );
or ( n380786 , n380782 , n380785 );
buf ( n380787 , n19520 );
or ( n380788 , n19595 , RI15b5d498_1048);
not ( n380789 , n380788 );
nand ( n380790 , n380787 , n380789 );
or ( n380791 , n380768 , n380790 );
nand ( n380792 , n380777 , n380786 , n380791 );
nor ( n380793 , n380746 , n380792 );
nand ( n380794 , n380705 , n380793 );
buf ( n380795 , n380794 );
not ( n380796 , n18242 );
nand ( n380797 , n18758 , n380796 );
nand ( n380798 , n18236 , RI15b5c778_1020);
buf ( n380799 , n380798 );
buf ( n380800 , n380799 );
and ( n380801 , n380800 , RI15b5c7f0_1021);
not ( n380802 , n380800 );
not ( n380803 , RI15b5c7f0_1021);
and ( n380804 , n380802 , n380803 );
nor ( n380805 , n380801 , n380804 );
and ( n380806 , n380797 , n380805 );
not ( n380807 , n380797 );
not ( n380808 , n380805 );
and ( n380809 , n380807 , n380808 );
nor ( n380810 , n380806 , n380809 );
not ( n380811 , n19285 );
not ( n380812 , n380811 );
not ( n380813 , n380812 );
nand ( n380814 , n380810 , n380813 );
not ( n380815 , n380803 );
nor ( n380816 , n380799 , n19336 );
not ( n380817 , n380816 );
or ( n380818 , n380815 , n380817 );
or ( n380819 , n380816 , n380803 );
nand ( n380820 , n380818 , n380819 );
nor ( n380821 , n19384 , n380820 );
not ( n380822 , n380821 );
nand ( n380823 , n19384 , n380820 );
nand ( n380824 , n380822 , n380823 );
and ( n380825 , n380824 , n19391 );
nor ( n380826 , n19399 , n18238 );
not ( n380827 , n380826 );
and ( n380828 , n380827 , n380803 );
not ( n380829 , n380827 );
and ( n380830 , n380829 , RI15b5c7f0_1021);
nor ( n380831 , n380828 , n380830 );
not ( n380832 , n380831 );
nand ( n380833 , n19477 , n19403 );
not ( n380834 , n380833 );
or ( n380835 , n380832 , n380834 );
or ( n380836 , n380833 , n380831 );
nand ( n380837 , n380835 , n380836 );
buf ( n380838 , n22761 );
and ( n380839 , n380837 , n380838 );
and ( n380840 , n19513 , RI15b63e88_1274);
nor ( n380841 , n380825 , n380839 , n380840 );
nand ( n380842 , n380814 , n380841 );
not ( n380843 , n380842 );
and ( n380844 , n19608 , RI15b62f88_1242);
nor ( n380845 , n19618 , n19610 );
buf ( n380846 , n380845 );
nand ( n380847 , n380846 , RI15b62bc8_1234);
and ( n380848 , n380847 , RI15b62f88_1242);
not ( n380849 , n380847 );
not ( n380850 , RI15b62f88_1242);
and ( n380851 , n380849 , n380850 );
nor ( n380852 , n380848 , n380851 );
not ( n380853 , n380852 );
and ( n380854 , n380853 , n19630 );
not ( n380855 , n380846 );
and ( n380856 , n380855 , n380850 );
not ( n380857 , n380855 );
and ( n380858 , n380857 , RI15b62f88_1242);
nor ( n380859 , n380856 , n380858 );
and ( n380860 , n380859 , n380238 );
nor ( n380861 , n380844 , n380854 , n380860 );
nand ( n380862 , n380843 , n380861 );
buf ( n380863 , n380862 );
buf ( n380864 , n22740 );
buf ( n380865 , RI15b3e9d0_1);
buf ( n380866 , n380865 );
not ( n380867 , n19906 );
not ( n380868 , n20524 );
buf ( n380869 , n380868 );
not ( n380870 , n380869 );
not ( n380871 , n380870 );
nor ( n380872 , n380871 , n19706 );
and ( n380873 , n380867 , n380872 );
or ( n380874 , n19998 , n20502 );
not ( n380875 , n20521 );
nand ( n380876 , n380874 , n380875 );
and ( n380877 , n380876 , RI15b4a118_392);
nor ( n380878 , n20529 , RI15b4a118_392);
not ( n380879 , n380878 );
not ( n380880 , n19998 );
or ( n380881 , n380879 , n380880 );
buf ( n380882 , n22353 );
or ( n380883 , n20558 , n380882 );
nand ( n380884 , n380883 , n20640 );
and ( n380885 , n380884 , RI15b4bf18_456);
not ( n380886 , RI15b4bf18_456);
and ( n380887 , n20558 , n380886 , RI15b4bea0_455);
nor ( n380888 , n380886 , RI15b4bea0_455);
nor ( n380889 , n380887 , n380888 );
not ( n380890 , n380889 );
and ( n380891 , n380890 , n20646 );
and ( n380892 , n20655 , RI15b4b018_424);
nor ( n380893 , n380885 , n380891 , n380892 );
nand ( n380894 , n380881 , n380893 );
nor ( n380895 , n380873 , n380877 , n380894 );
nor ( n380896 , n380867 , n19922 );
or ( n380897 , n380896 , n19943 );
nand ( n380898 , n380897 , n19706 );
nand ( n380899 , n380895 , n380898 );
buf ( n380900 , n380899 );
buf ( n380901 , n380865 );
buf ( n380902 , n22714 );
buf ( n380903 , RI15b3ea48_2);
buf ( n380904 , n380903 );
buf ( n380905 , RI15b479b8_308);
buf ( n380906 , RI15b3ea48_2);
buf ( n380907 , n380906 );
nand ( n380908 , n22142 , n22148 );
or ( n380909 , n380908 , n22133 );
or ( n380910 , n22102 , n380909 );
not ( n380911 , n22205 );
nor ( n380912 , n22123 , n22225 );
and ( n380913 , n380911 , n380912 );
and ( n380914 , n22203 , n380913 );
not ( n380915 , n380913 );
and ( n380916 , n380909 , n380915 , n19912 );
nor ( n380917 , n380916 , n22217 );
buf ( n380918 , n22124 );
buf ( n380919 , n22150 );
nor ( n380920 , n380918 , n380919 );
or ( n380921 , n380917 , n380920 );
nand ( n380922 , n380921 , n20623 );
nand ( n380923 , n20461 , RI15b3fdf8_44);
or ( n380924 , n380923 , RI15b3fd80_43);
not ( n380925 , n22210 );
or ( n380926 , n380924 , n380925 );
and ( n380927 , n380922 , n380926 );
nor ( n380928 , n380927 , n22236 );
not ( n380929 , RI15b41ec8_114);
or ( n380930 , n380928 , n380929 );
not ( n380931 , n380926 );
nor ( n380932 , n380920 , n380931 );
or ( n380933 , n380917 , n380932 );
or ( n380934 , n22293 , n380933 );
or ( n380935 , n380926 , n22299 );
nand ( n380936 , n380930 , n380934 , n380935 );
nor ( n380937 , n380914 , n380936 );
nand ( n380938 , n380910 , n380937 );
buf ( n380939 , n380938 );
buf ( n380940 , RI15b3e9d0_1);
buf ( n380941 , n380940 );
buf ( n380942 , RI15b3e9d0_1);
buf ( n380943 , n380942 );
buf ( n380944 , n380906 );
not ( n380945 , RI15b66570_1357);
not ( n380946 , n22084 );
or ( n380947 , n380945 , n380946 );
or ( n380948 , n22085 , RI15b66570_1357);
nand ( n380949 , n380947 , n380948 );
nor ( n380950 , n22080 , n380949 );
not ( n380951 , n380950 );
and ( n380952 , n22084 , n22098 );
not ( n380953 , n380952 );
not ( n380954 , RI15b665e8_1358);
and ( n380955 , n380953 , n380954 );
and ( n380956 , n380952 , RI15b665e8_1358);
nor ( n380957 , n380955 , n380956 );
not ( n380958 , n380957 );
not ( n380959 , n380958 );
or ( n380960 , n380951 , n380959 );
not ( n380961 , n380957 );
or ( n380962 , n380961 , n380950 );
nand ( n380963 , n380960 , n380962 );
and ( n380964 , n380963 , n22097 );
not ( n380965 , RI15b665e8_1358);
nor ( n380966 , n22094 , n380965 );
nor ( n380967 , n380964 , n380966 );
buf ( n380968 , n380967 );
or ( n380969 , n380968 , n380909 );
nand ( n380970 , n22196 , n22186 );
buf ( n380971 , n380970 );
or ( n380972 , n380971 , n20638 );
nand ( n380973 , n380972 , n22094 );
not ( n380974 , n22043 );
nand ( n380975 , n380974 , RI15b666d8_1360);
not ( n380976 , n380975 );
not ( n380977 , RI15b66228_1350);
and ( n380978 , n380976 , n380977 );
and ( n380979 , n380975 , RI15b66228_1350);
nor ( n380980 , n380978 , n380979 );
not ( n380981 , n380980 );
and ( n380982 , n380973 , n380981 );
nor ( n380983 , n380981 , n22199 );
and ( n380984 , n380983 , n380971 );
nor ( n380985 , n380982 , n380984 );
not ( n380986 , n380985 );
and ( n380987 , n380986 , n380913 );
not ( n380988 , RI15b41f40_115);
or ( n380989 , n380928 , n380988 );
not ( n380990 , n22287 );
not ( n380991 , n22020 );
and ( n380992 , n380990 , n380991 );
and ( n380993 , n22287 , n22252 );
nor ( n380994 , n380992 , n380993 );
or ( n380995 , n380994 , n380933 );
or ( n380996 , n20376 , n22298 );
or ( n380997 , n380926 , n380996 );
nand ( n380998 , n380989 , n380995 , n380997 );
nor ( n380999 , n380987 , n380998 );
nand ( n381000 , n380969 , n380999 );
buf ( n381001 , n381000 );
buf ( n381002 , RI15b47b98_312);
buf ( n381003 , n380903 );
buf ( n381004 , RI15b3e9d0_1);
buf ( n381005 , n381004 );
buf ( n381006 , RI15b3e9d0_1);
buf ( n381007 , n381006 );
not ( n381008 , RI15b523e0_671);
or ( n381009 , RI15b51300_635 , RI15b51378_636 , RI15b513f0_637 , RI15b51468_638);
not ( n381010 , RI15b52368_670);
nand ( n381011 , n381010 , RI15b522f0_669);
nor ( n381012 , n381008 , n381009 , n381011 , RI15b52458_672);
not ( n381013 , RI15b52278_668);
and ( n381014 , n381012 , n381013 );
buf ( n381015 , n381014 );
or ( n381016 , n381015 , n22017 );
buf ( n381017 , n381014 );
nand ( n381018 , n381017 , RI15b534c0_707);
nand ( n381019 , n381016 , n381018 );
buf ( n381020 , n381019 );
buf ( n381021 , RI15b3ea48_2);
buf ( n381022 , n381021 );
buf ( n381023 , n22479 );
not ( n381024 , n20589 );
not ( n381025 , n20590 );
nor ( n381026 , n20116 , n20292 , n20591 );
and ( n381027 , n381025 , n381026 );
not ( n381028 , n20603 );
and ( n381029 , n381027 , n381028 );
nor ( n381030 , n381029 , n20519 );
nand ( n381031 , n381024 , n381030 , n20607 );
nor ( n381032 , n20577 , n20519 );
not ( n381033 , n20605 );
nand ( n381034 , n381032 , n381033 );
not ( n381035 , n381034 );
not ( n381036 , n381035 );
nand ( n381037 , n381031 , n381036 , n20501 );
nand ( n381038 , n20332 , n20251 , n20501 );
or ( n381039 , n20605 , n381038 );
not ( n381040 , n20478 );
not ( n381041 , n20483 );
nand ( n381042 , n20429 , RI15b3fc90_41);
nand ( n381043 , n381041 , n20479 , n381042 );
nand ( n381044 , n381040 , n381043 );
nand ( n381045 , n20470 , n381044 );
buf ( n381046 , n381045 );
not ( n381047 , n381046 );
not ( n381048 , n381047 );
or ( n381049 , n381039 , n381048 );
nand ( n381050 , n20589 , n20501 );
not ( n381051 , n381032 );
not ( n381052 , n381051 );
nand ( n381053 , n381052 , n381027 );
nand ( n381054 , n381049 , n381050 , n381053 );
or ( n381055 , n381037 , n381054 );
not ( n381056 , n381055 );
or ( n381057 , n381056 , n19957 );
not ( n381058 , RI15b40050_49);
not ( n381059 , n381039 );
not ( n381060 , n381046 );
not ( n381061 , n381060 );
nand ( n381062 , n381059 , n381061 );
or ( n381063 , n381058 , n381062 );
nand ( n381064 , RI15b49380_363 , RI15b493f8_364);
not ( n381065 , RI15b49470_365);
nor ( n381066 , n381064 , n381065 );
not ( n381067 , n381066 );
and ( n381068 , n381067 , RI15b494e8_366);
not ( n381069 , n381067 );
and ( n381070 , n381069 , n19957 );
nor ( n381071 , n381068 , n381070 );
not ( n381072 , n381027 );
nor ( n381073 , n381072 , n381038 );
buf ( n381074 , n381073 );
buf ( n381075 , n381074 );
buf ( n381076 , n381075 );
not ( n381077 , n381076 );
or ( n381078 , n381071 , n381077 );
nand ( n381079 , n381057 , n381063 , n381078 );
buf ( n381080 , n381079 );
buf ( n381081 , RI15b3e9d0_1);
buf ( n381082 , n381081 );
buf ( n381083 , n20663 );
buf ( n381084 , n380903 );
nor ( n381085 , RI15b515d0_641 , RI15b51648_642);
nor ( n381086 , RI15b516c0_643 , RI15b51738_644);
nor ( n381087 , RI15b517b0_645 , RI15b51828_646);
nor ( n381088 , RI15b518a0_647 , RI15b51918_648);
nand ( n381089 , n381085 , n381086 , n381087 , n381088 );
nor ( n381090 , RI15b52110_665 , RI15b52188_666);
nor ( n381091 , RI15b514e0_639 , RI15b51558_640);
not ( n381092 , RI15b52200_667);
nand ( n381093 , n381090 , n381091 , n381092 );
nor ( n381094 , n381089 , n381093 );
not ( n381095 , n381094 );
nor ( n381096 , RI15b51990_649 , RI15b51a08_650);
nor ( n381097 , RI15b51a80_651 , RI15b51af8_652);
nor ( n381098 , RI15b51b70_653 , RI15b51be8_654);
nor ( n381099 , RI15b51c60_655 , RI15b51cd8_656);
nand ( n381100 , n381096 , n381097 , n381098 , n381099 );
nor ( n381101 , RI15b51d50_657 , RI15b51dc8_658);
nor ( n381102 , RI15b51e40_659 , RI15b51eb8_660);
nor ( n381103 , RI15b51f30_661 , RI15b51fa8_662);
nor ( n381104 , RI15b52020_663 , RI15b52098_664);
nand ( n381105 , n381101 , n381102 , n381103 , n381104 );
nor ( n381106 , n381100 , n381105 );
not ( n381107 , n381106 );
or ( n381108 , n381095 , n381107 );
nand ( n381109 , n381108 , RI15b52278_668);
buf ( n381110 , n381109 );
not ( n381111 , n381110 );
not ( n381112 , n380396 );
and ( n381113 , n381111 , n381112 );
buf ( n381114 , n381109 );
and ( n381115 , n381114 , RI15b65f58_1344);
nor ( n381116 , n381113 , n381115 );
buf ( n381117 , n381116 );
buf ( n381118 , n381117 );
nand ( n381119 , n381106 , n381094 );
nand ( n381120 , n381119 , RI15b52278_668);
buf ( n381121 , n381120 );
not ( n381122 , n381121 );
not ( n381123 , n380378 );
and ( n381124 , n381122 , n381123 );
buf ( n381125 , n381109 );
and ( n381126 , n381125 , RI15b65e68_1342);
nor ( n381127 , n381124 , n381126 );
not ( n381128 , n381121 );
not ( n381129 , n380386 );
and ( n381130 , n381128 , n381129 );
and ( n381131 , n381125 , RI15b65ee0_1343);
nor ( n381132 , n381130 , n381131 );
nand ( n381133 , n381127 , n381132 );
not ( n381134 , n381133 );
not ( n381135 , RI15b666d8_1360);
not ( n381136 , n381110 );
or ( n381137 , n381135 , n381136 );
buf ( n381138 , n381110 );
or ( n381139 , n381138 , n380267 );
nand ( n381140 , n381137 , n381139 );
not ( n381141 , n381140 );
not ( n381142 , n381141 );
not ( n381143 , n381142 );
not ( n381144 , n381143 );
not ( n381145 , n381144 );
not ( n381146 , n381145 );
not ( n381147 , n381146 );
not ( n381148 , n381147 );
not ( n381149 , n381148 );
or ( n381150 , n381134 , n381149 );
not ( n381151 , n381121 );
not ( n381152 , n380360 );
and ( n381153 , n381151 , n381152 );
and ( n381154 , n381114 , RI15b65d78_1340);
nor ( n381155 , n381153 , n381154 );
not ( n381156 , n381121 );
not ( n381157 , n380342 );
and ( n381158 , n381156 , n381157 );
and ( n381159 , n381125 , RI15b65c10_1337);
nor ( n381160 , n381158 , n381159 );
not ( n381161 , n381121 );
not ( n381162 , n380370 );
and ( n381163 , n381161 , n381162 );
and ( n381164 , n381125 , RI15b65df0_1341);
nor ( n381165 , n381163 , n381164 );
nand ( n381166 , n381155 , n381160 , n381165 );
not ( n381167 , n381121 );
not ( n381168 , n380317 );
and ( n381169 , n381167 , n381168 );
and ( n381170 , n381114 , RI15b65940_1331);
nor ( n381171 , n381169 , n381170 );
not ( n381172 , n381121 );
not ( n381173 , RI15b64ba8_1302);
not ( n381174 , n381173 );
and ( n381175 , n381172 , n381174 );
and ( n381176 , n381114 , RI15b65aa8_1334);
nor ( n381177 , n381175 , n381176 );
nand ( n381178 , n381171 , n381177 );
nor ( n381179 , n381166 , n381178 );
not ( n381180 , n381121 );
not ( n381181 , RI15b649c8_1298);
not ( n381182 , n381181 );
and ( n381183 , n381180 , n381182 );
and ( n381184 , n381125 , RI15b658c8_1330);
nor ( n381185 , n381183 , n381184 );
not ( n381186 , n381121 );
not ( n381187 , n380310 );
and ( n381188 , n381186 , n381187 );
and ( n381189 , n381125 , RI15b65850_1329);
nor ( n381190 , n381188 , n381189 );
nand ( n381191 , n381185 , n381190 );
not ( n381192 , n381121 );
not ( n381193 , n380324 );
and ( n381194 , n381192 , n381193 );
and ( n381195 , n381114 , RI15b65b20_1335);
nor ( n381196 , n381194 , n381195 );
buf ( n381197 , n381196 );
nor ( n381198 , n381121 , n380331 );
not ( n381199 , n381198 );
nand ( n381200 , n381121 , RI15b65b98_1336);
nand ( n381201 , n381199 , n381200 );
not ( n381202 , n381201 );
nand ( n381203 , n381197 , n381202 );
nor ( n381204 , n381191 , n381203 );
not ( n381205 , n381121 );
not ( n381206 , RI15b64ab8_1300);
not ( n381207 , n381206 );
and ( n381208 , n381205 , n381207 );
and ( n381209 , n381125 , RI15b659b8_1332);
nor ( n381210 , n381208 , n381209 );
not ( n381211 , n381121 );
not ( n381212 , RI15b64b30_1301);
not ( n381213 , n381212 );
and ( n381214 , n381211 , n381213 );
and ( n381215 , n381125 , RI15b65a30_1333);
nor ( n381216 , n381214 , n381215 );
nand ( n381217 , n381210 , n381216 );
or ( n381218 , n381114 , RI15b64e00_1307);
nand ( n381219 , n381121 , n22028 );
nand ( n381220 , n381218 , n381219 );
buf ( n381221 , n381119 );
and ( n381222 , RI15b52278_668 , RI15b64d88_1306);
and ( n381223 , n381221 , n381222 );
and ( n381224 , n381121 , RI15b65c88_1338);
nor ( n381225 , n381223 , n381224 );
nand ( n381226 , n381220 , n381225 );
nor ( n381227 , n381217 , n381226 );
nand ( n381228 , n381179 , n381204 , n381227 );
not ( n381229 , n381228 );
nor ( n381230 , n381229 , n381143 );
not ( n381231 , n381230 );
nand ( n381232 , n381150 , n381231 );
and ( n381233 , n381118 , n381232 );
not ( n381234 , n381118 );
or ( n381235 , n381228 , n381133 );
nand ( n381236 , n381235 , n381148 );
and ( n381237 , n381234 , n381236 );
nor ( n381238 , n381233 , n381237 );
not ( n381239 , n381238 );
buf ( n381240 , n381165 );
buf ( n381241 , n381155 );
not ( n381242 , n381241 );
not ( n381243 , n381242 );
buf ( n381244 , n381146 );
not ( n381245 , n381244 );
or ( n381246 , n381243 , n381245 );
buf ( n381247 , n381226 );
not ( n381248 , n381247 );
not ( n381249 , n381146 );
or ( n381250 , n381248 , n381249 );
buf ( n381251 , n381171 );
not ( n381252 , n381251 );
nor ( n381253 , n381191 , n381252 );
not ( n381254 , n381217 );
nand ( n381255 , n381253 , n381254 );
not ( n381256 , n381255 );
buf ( n381257 , n381177 );
nand ( n381258 , n381256 , n381257 );
buf ( n381259 , n381203 );
nor ( n381260 , n381258 , n381259 );
buf ( n381261 , n381160 );
nand ( n381262 , n381260 , n381261 );
not ( n381263 , n381144 );
not ( n381264 , n381263 );
nand ( n381265 , n381262 , n381264 );
nand ( n381266 , n381250 , n381265 );
not ( n381267 , n381266 );
nand ( n381268 , n381246 , n381267 );
and ( n381269 , n381240 , n381268 );
not ( n381270 , n381240 );
not ( n381271 , n381241 );
or ( n381272 , n381262 , n381247 , n381271 );
nand ( n381273 , n381272 , n381148 );
and ( n381274 , n381270 , n381273 );
nor ( n381275 , n381269 , n381274 );
buf ( n381276 , n381220 );
not ( n381277 , n381276 );
buf ( n381278 , n381225 );
not ( n381279 , n381278 );
not ( n381280 , n381279 );
not ( n381281 , n381146 );
or ( n381282 , n381280 , n381281 );
nand ( n381283 , n381282 , n381265 );
not ( n381284 , n381283 );
or ( n381285 , n381277 , n381284 );
not ( n381286 , n381262 );
and ( n381287 , n381286 , n381278 );
nor ( n381288 , n381287 , n381147 );
or ( n381289 , n381288 , n381276 );
nand ( n381290 , n381285 , n381289 );
not ( n381291 , n381278 );
not ( n381292 , n381291 );
and ( n381293 , n381265 , n381292 );
not ( n381294 , n381265 );
and ( n381295 , n381294 , n381291 );
nor ( n381296 , n381293 , n381295 );
not ( n381297 , n381261 );
not ( n381298 , n381297 );
not ( n381299 , n381298 );
not ( n381300 , n381259 );
not ( n381301 , n381144 );
or ( n381302 , n381300 , n381301 );
not ( n381303 , n381143 );
nand ( n381304 , n381258 , n381303 );
nand ( n381305 , n381302 , n381304 );
not ( n381306 , n381305 );
or ( n381307 , n381299 , n381306 );
or ( n381308 , n381260 , n381263 );
nand ( n381309 , n381308 , n381297 );
nand ( n381310 , n381307 , n381309 );
not ( n381311 , n381230 );
buf ( n381312 , n381127 );
buf ( n381313 , n381312 );
not ( n381314 , n381313 );
and ( n381315 , n381311 , n381314 );
and ( n381316 , n381230 , n381313 );
nor ( n381317 , n381315 , n381316 );
nor ( n381318 , n381141 , n381312 );
or ( n381319 , n381230 , n381318 );
buf ( n381320 , n381132 );
nand ( n381321 , n381319 , n381320 );
nand ( n381322 , n381317 , n381321 );
nor ( n381323 , n381310 , n381322 );
buf ( n381324 , n381197 );
not ( n381325 , n381324 );
not ( n381326 , n381325 );
not ( n381327 , n381304 );
or ( n381328 , n381326 , n381327 );
buf ( n381329 , n381325 );
or ( n381330 , n381304 , n381329 );
nand ( n381331 , n381328 , n381330 );
nor ( n381332 , n381230 , n381318 , n381320 );
not ( n381333 , n381257 );
not ( n381334 , n381333 );
buf ( n381335 , n381140 );
nand ( n381336 , n381255 , n381335 );
not ( n381337 , n381336 );
or ( n381338 , n381334 , n381337 );
not ( n381339 , n381257 );
or ( n381340 , n381336 , n381339 );
nand ( n381341 , n381338 , n381340 );
nor ( n381342 , n381332 , n381341 );
buf ( n381343 , n381216 );
not ( n381344 , n381343 );
not ( n381345 , n381344 );
buf ( n381346 , n381210 );
not ( n381347 , n381346 );
not ( n381348 , n381253 );
or ( n381349 , n381347 , n381348 );
nand ( n381350 , n381349 , n381335 );
not ( n381351 , n381350 );
or ( n381352 , n381345 , n381351 );
not ( n381353 , n381343 );
or ( n381354 , n381350 , n381353 );
nand ( n381355 , n381352 , n381354 );
nor ( n381356 , n381253 , n381141 );
buf ( n381357 , n381346 );
not ( n381358 , n381357 );
and ( n381359 , n381356 , n381358 );
not ( n381360 , n381356 );
and ( n381361 , n381360 , n381357 );
nor ( n381362 , n381359 , n381361 );
nand ( n381363 , n381140 , n381191 );
buf ( n381364 , n381251 );
and ( n381365 , n381363 , n381364 );
not ( n381366 , n381363 );
not ( n381367 , n381364 );
and ( n381368 , n381366 , n381367 );
nor ( n381369 , n381365 , n381368 );
nor ( n381370 , n381355 , n381362 , n381369 , n381191 );
nand ( n381371 , n381342 , n381370 );
nor ( n381372 , n381331 , n381371 );
not ( n381373 , n381324 );
not ( n381374 , n381373 );
not ( n381375 , n381144 );
or ( n381376 , n381374 , n381375 );
nand ( n381377 , n381376 , n381304 );
buf ( n381378 , n381202 );
and ( n381379 , n381377 , n381378 );
or ( n381380 , n381258 , n381373 );
nand ( n381381 , n381380 , n381144 );
not ( n381382 , n381378 );
and ( n381383 , n381381 , n381382 );
nor ( n381384 , n381379 , n381383 );
nand ( n381385 , n381323 , n381372 , n381384 );
nor ( n381386 , n381290 , n381296 , n381385 );
not ( n381387 , n381242 );
and ( n381388 , n381266 , n381387 );
or ( n381389 , n381262 , n381247 );
nand ( n381390 , n381389 , n381244 );
and ( n381391 , n381390 , n381242 );
nor ( n381392 , n381388 , n381391 );
nand ( n381393 , n381275 , n381386 , n381392 );
buf ( n381394 , n381148 );
buf ( n381395 , n381394 );
nand ( n381396 , n381393 , n381395 );
not ( n381397 , n381396 );
or ( n381398 , n381239 , n381397 );
nand ( n381399 , n17994 , n18077 );
or ( n381400 , n18181 , n381399 );
not ( n381401 , n381400 );
nand ( n381402 , n381398 , n381401 );
buf ( n381403 , n381395 );
not ( n381404 , n381403 );
nor ( n381405 , n381402 , n381404 );
buf ( n381406 , n381405 );
not ( n381407 , n381406 );
buf ( n381408 , n381298 );
buf ( n381409 , n381408 );
or ( n381410 , n381407 , n381409 );
not ( n381411 , n381238 );
not ( n381412 , n381393 );
not ( n381413 , n381412 );
or ( n381414 , n381411 , n381413 );
nand ( n381415 , n381414 , n381403 );
nand ( n381416 , n381415 , n381401 );
not ( n381417 , n381416 );
nand ( n381418 , n381417 , n381310 );
nand ( n381419 , n18100 , n18185 );
not ( n381420 , n381419 );
buf ( n381421 , n381420 );
buf ( n381422 , n381421 );
not ( n381423 , n381422 );
buf ( n381424 , n381423 );
nor ( n381425 , RI15b548e8_750 , RI15b54b40_755);
not ( n381426 , RI15b54bb8_756);
nand ( n381427 , n381425 , n381426 );
nor ( n381428 , RI15b54960_751 , RI15b549d8_752);
nor ( n381429 , RI15b54a50_753 , RI15b54ac8_754);
nand ( n381430 , n381428 , n381429 );
nor ( n381431 , n381427 , n381430 );
and ( n381432 , n381431 , RI15b55770_781);
nand ( n381433 , n381425 , RI15b55770_781);
nor ( n381434 , n381433 , n381430 );
not ( n381435 , RI15b54bb8_756);
nor ( n381436 , n381434 , n381435 );
nor ( n381437 , n381432 , n381436 );
not ( n381438 , n381434 );
nor ( n381439 , n381437 , n381438 );
not ( n381440 , RI15b55770_781);
nor ( n381441 , n381431 , n381440 );
not ( n381442 , RI15b54c30_757);
and ( n381443 , n381441 , n381442 );
not ( n381444 , n381441 );
and ( n381445 , n381444 , RI15b54c30_757);
nor ( n381446 , n381443 , n381445 );
nand ( n381447 , n381439 , n381446 );
or ( n381448 , n381424 , n381447 );
nor ( n381449 , n381419 , RI15b55770_781);
not ( n381450 , n381449 );
nand ( n381451 , n381448 , n381450 );
not ( n381452 , RI15b54ca8_758);
nand ( n381453 , n381431 , n381442 );
nand ( n381454 , n381453 , RI15b55770_781);
not ( n381455 , n381454 );
or ( n381456 , n381452 , n381455 );
or ( n381457 , n381454 , RI15b54ca8_758);
nand ( n381458 , n381456 , n381457 );
and ( n381459 , n381451 , n381458 );
nand ( n381460 , n381420 , RI15b55770_781);
not ( n381461 , n381460 );
not ( n381462 , n381447 );
nor ( n381463 , n381462 , n381458 );
and ( n381464 , n381461 , n381463 );
nor ( n381465 , n381459 , n381464 );
and ( n381466 , n381418 , n381465 );
nand ( n381467 , n18132 , n18144 );
nor ( n381468 , n381467 , n18078 );
not ( n381469 , n18077 );
not ( n381470 , n18127 );
or ( n381471 , n381469 , n381470 );
not ( n381472 , n21335 );
nand ( n381473 , n381471 , n381472 );
nor ( n381474 , n381468 , n381473 );
buf ( n381475 , n381474 );
buf ( n381476 , n18183 );
buf ( n381477 , n381476 );
and ( n381478 , n18181 , n381477 );
nand ( n381479 , n18147 , n18077 );
or ( n381480 , n381479 , n18091 );
or ( n381481 , n18203 , n18078 );
nand ( n381482 , n381480 , n381481 , n18077 );
nor ( n381483 , n381478 , n381482 );
nand ( n381484 , n381475 , n381483 );
buf ( n381485 , n381484 );
buf ( n381486 , n381485 );
nand ( n381487 , n381486 , RI15b52f98_696);
nand ( n381488 , n381410 , n381466 , n381487 );
buf ( n381489 , n381488 );
buf ( n381490 , RI15b3e9d0_1);
buf ( n381491 , n381490 );
and ( n381492 , n380228 , n380726 );
buf ( n381493 , n380766 );
and ( n381494 , n381492 , n381493 );
not ( n381495 , n381494 );
buf ( n381496 , n19645 );
buf ( n381497 , n381496 );
not ( n381498 , n381497 );
not ( n381499 , n380677 );
not ( n381500 , n381499 );
or ( n381501 , n381498 , n381500 );
nand ( n381502 , n381501 , n380686 );
and ( n381503 , n381502 , n380678 );
nand ( n381504 , n380698 , n380522 );
nor ( n381505 , n381499 , n381504 );
nor ( n381506 , n381503 , n381505 );
not ( n381507 , n381506 );
not ( n381508 , n381507 );
or ( n381509 , n381495 , n381508 );
not ( n381510 , n380539 );
and ( n381511 , n380708 , n381510 );
and ( n381512 , n380710 , n380539 );
nor ( n381513 , n381511 , n381512 );
not ( n381514 , n380710 );
not ( n381515 , n380708 );
nand ( n381516 , n381514 , n381515 );
and ( n381517 , n381513 , n381516 );
not ( n381518 , n19645 );
nor ( n381519 , n381517 , n380562 , n381518 );
not ( n381520 , n380711 );
not ( n381521 , n380283 );
and ( n381522 , n381521 , n19641 );
and ( n381523 , n381520 , n381522 , n381510 , n380562 );
or ( n381524 , n381519 , n381523 );
not ( n381525 , n380736 );
and ( n381526 , n381525 , n380741 );
nand ( n381527 , n381526 , n380757 );
not ( n381528 , n381527 );
and ( n381529 , n381524 , n381528 );
not ( n381530 , n381494 );
not ( n381531 , n380750 );
and ( n381532 , n381527 , n381530 , n381531 );
nor ( n381533 , n381532 , n19630 );
nand ( n381534 , n380211 , n380754 );
nor ( n381535 , n381534 , n380728 );
or ( n381536 , n381533 , n381535 );
nand ( n381537 , n381536 , n19595 );
nand ( n381538 , n19203 , RI15b586c8_882);
or ( n381539 , n381538 , n19209 );
not ( n381540 , n380232 );
buf ( n381541 , n381540 );
or ( n381542 , n381539 , n381541 );
nand ( n381543 , n381537 , n381542 );
and ( n381544 , n381543 , n380775 );
or ( n381545 , n381544 , n18410 );
buf ( n381546 , n380328 );
not ( n381547 , n381546 );
buf ( n381548 , n381547 );
buf ( n381549 , n381548 );
buf ( n381550 , n381549 );
not ( n381551 , n381550 );
not ( n381552 , n381535 );
not ( n381553 , n381542 );
not ( n381554 , n381553 );
and ( n381555 , n381552 , n381554 );
nor ( n381556 , n381555 , n381533 );
not ( n381557 , n381556 );
or ( n381558 , n381551 , n381557 );
not ( n381559 , n18873 );
or ( n381560 , n381559 , n380788 );
or ( n381561 , n381542 , n381560 );
nand ( n381562 , n381545 , n381558 , n381561 );
nor ( n381563 , n381529 , n381562 );
nand ( n381564 , n381509 , n381563 );
buf ( n381565 , n381564 );
buf ( n381566 , RI15b3e9d0_1);
buf ( n381567 , n381566 );
and ( n381568 , n380229 , n380733 );
nand ( n381569 , n381568 , n381493 );
not ( n381570 , n381569 );
not ( n381571 , n381570 );
buf ( n381572 , n380237 );
not ( n381573 , n381572 );
nand ( n381574 , n380624 , n380649 );
not ( n381575 , n381574 );
not ( n381576 , n380665 );
nand ( n381577 , n381575 , n381576 );
buf ( n381578 , n380675 );
nor ( n381579 , n381577 , n381578 );
not ( n381580 , n381579 );
or ( n381581 , n381573 , n381580 );
nand ( n381582 , n381581 , n380686 );
and ( n381583 , n380634 , n380642 );
not ( n381584 , n381583 );
and ( n381585 , n381582 , n381584 );
nand ( n381586 , n381583 , n380698 );
nor ( n381587 , n381579 , n381586 );
nor ( n381588 , n381585 , n381587 );
not ( n381589 , n381588 );
not ( n381590 , n381589 );
or ( n381591 , n381571 , n381590 );
and ( n381592 , n381520 , n380540 );
not ( n381593 , n19646 );
nor ( n381594 , n381592 , n381593 );
nand ( n381595 , n380711 , n380539 );
and ( n381596 , n381594 , n381595 );
not ( n381597 , n380757 );
or ( n381598 , n380743 , n381597 );
not ( n381599 , n381598 );
and ( n381600 , n381596 , n381599 );
not ( n381601 , n380750 );
and ( n381602 , n381598 , n381569 , n381601 );
nor ( n381603 , n381602 , n19630 );
nor ( n381604 , n380755 , n380728 );
or ( n381605 , n381603 , n381604 );
nand ( n381606 , n381605 , n19595 );
or ( n381607 , n380764 , n381540 );
nand ( n381608 , n381606 , n381607 );
and ( n381609 , n381608 , n380775 );
or ( n381610 , n381609 , n18728 );
buf ( n381611 , n380301 );
not ( n381612 , n381611 );
buf ( n381613 , n381612 );
buf ( n381614 , n381613 );
not ( n381615 , n381614 );
buf ( n381616 , n381615 );
not ( n381617 , n381607 );
nor ( n381618 , n381604 , n381617 );
or ( n381619 , n381603 , n381618 );
or ( n381620 , n381616 , n381619 );
nand ( n381621 , n19145 , n380789 );
or ( n381622 , n381607 , n381621 );
nand ( n381623 , n381610 , n381620 , n381622 );
nor ( n381624 , n381600 , n381623 );
nand ( n381625 , n381591 , n381624 );
buf ( n381626 , n381625 );
buf ( n381627 , n379895 );
buf ( n381628 , n22406 );
not ( n381629 , RI15b55d10_793);
not ( n381630 , n380000 );
or ( n381631 , n381629 , n381630 );
buf ( n381632 , n17593 );
xor ( n381633 , RI15b50fb8_628 , n381632 );
nor ( n381634 , n21555 , n381633 );
not ( n381635 , n380013 );
and ( n381636 , n381634 , n381635 );
and ( n381637 , n381636 , RI15b4ea38_548);
not ( n381638 , n17623 );
and ( n381639 , n381634 , n381638 );
and ( n381640 , n381639 , RI15b4e678_540);
nor ( n381641 , n381637 , n381640 );
not ( n381642 , n380031 );
and ( n381643 , n381634 , n381642 );
and ( n381644 , n381643 , RI15b4edf8_556);
not ( n381645 , n380007 );
not ( n381646 , n381645 );
buf ( n381647 , n380022 );
buf ( n381648 , n381647 );
not ( n381649 , n381648 );
not ( n381650 , n381649 );
buf ( n381651 , n381650 );
and ( n381652 , n381651 , RI15b4db38_516);
buf ( n381653 , n380047 );
buf ( n381654 , n381653 );
buf ( n381655 , n381654 );
not ( n381656 , n381655 );
not ( n381657 , n381656 );
and ( n381658 , n381657 , RI15b4fcf8_588);
nor ( n381659 , n381652 , n381658 );
not ( n381660 , n17583 );
nor ( n381661 , n381660 , n381633 );
and ( n381662 , n381661 , RI15b4f938_580);
nor ( n381663 , n381633 , n17605 );
and ( n381664 , n381663 , RI15b4f1b8_564);
nor ( n381665 , n381662 , n381664 );
not ( n381666 , n381633 );
nor ( n381667 , n381666 , n17605 );
and ( n381668 , n381667 , RI15b4d3b8_500);
and ( n381669 , n20767 , n381633 );
and ( n381670 , n381669 , RI15b4d778_508);
nor ( n381671 , n381668 , n381670 );
nor ( n381672 , n381666 , n17685 );
and ( n381673 , n381672 , RI15b4def8_524);
nor ( n381674 , n17615 , n381633 );
and ( n381675 , n381674 , RI15b4f578_572);
nor ( n381676 , n381673 , n381675 );
nand ( n381677 , n381659 , n381665 , n381671 , n381676 );
and ( n381678 , n381646 , n381677 );
and ( n381679 , n21554 , n381633 );
and ( n381680 , n381679 , n381638 );
and ( n381681 , n381680 , RI15b4c878_476);
nor ( n381682 , n381644 , n381678 , n381681 );
buf ( n381683 , n17594 );
and ( n381684 , n381679 , n381683 );
and ( n381685 , n381684 , RI15b4c4b8_468);
and ( n381686 , n381634 , n381683 );
and ( n381687 , n381686 , RI15b4e2b8_532);
nor ( n381688 , n381685 , n381687 );
and ( n381689 , n381679 , n381635 );
and ( n381690 , n381689 , RI15b4cc38_484);
and ( n381691 , n381679 , n381642 );
and ( n381692 , n381691 , RI15b4cff8_492);
nor ( n381693 , n381690 , n381692 );
nand ( n381694 , n381641 , n381682 , n381688 , n381693 );
buf ( n381695 , n379989 );
not ( n381696 , n381695 );
and ( n381697 , n381694 , n381696 );
not ( n381698 , RI15b55d10_793);
not ( n381699 , n379962 );
or ( n381700 , n381698 , n381699 );
or ( n381701 , n379962 , RI15b55d10_793);
nand ( n381702 , n381700 , n381701 );
and ( n381703 , n379949 , n381702 );
nor ( n381704 , n381697 , n381703 );
nand ( n381705 , n381631 , n381704 );
buf ( n381706 , n381705 );
buf ( n381707 , RI15b3ea48_2);
buf ( n381708 , n381707 );
nand ( n381709 , RI15b508b0_613 , RI15b50928_614);
not ( n381710 , RI15b509a0_615);
nor ( n381711 , n381709 , n381710 );
nand ( n381712 , n381711 , RI15b50a18_616);
not ( n381713 , n381712 );
and ( n381714 , n381713 , RI15b50a90_617);
not ( n381715 , RI15b50b08_618);
nand ( n381716 , n381714 , n381715 );
not ( n381717 , n381716 );
buf ( n381718 , n21539 );
not ( n381719 , n381718 );
not ( n381720 , n381719 );
nand ( n381721 , n381717 , n381720 );
not ( n381722 , n381718 );
nand ( n381723 , n381722 , RI15b50b08_618);
not ( n381724 , n381714 );
nand ( n381725 , n381724 , RI15b50b08_618);
and ( n381726 , n381721 , n381723 , n381725 );
not ( n381727 , n381726 );
nor ( n381728 , n21382 , n21527 , n21534 );
and ( n381729 , n21538 , RI15b50a18_616);
not ( n381730 , RI15b50a18_616);
nand ( n381731 , n381711 , n381730 );
or ( n381732 , n21378 , n381731 );
not ( n381733 , n381711 );
nand ( n381734 , n381733 , RI15b50a18_616);
nand ( n381735 , n381732 , n381734 );
nor ( n381736 , n381729 , n381735 );
not ( n381737 , n381736 );
nor ( n381738 , n381709 , RI15b509a0_615);
nand ( n381739 , n21539 , n381738 );
nand ( n381740 , n21538 , RI15b509a0_615);
nand ( n381741 , n381709 , RI15b509a0_615);
and ( n381742 , n381739 , n381740 , n381741 );
not ( n381743 , n381742 );
and ( n381744 , n381728 , n381737 , n21543 , n381743 );
nand ( n381745 , n21522 , n381744 );
nand ( n381746 , n381719 , RI15b50a90_617);
buf ( n381747 , n381718 );
or ( n381748 , n381712 , RI15b50a90_617);
not ( n381749 , n381748 );
nand ( n381750 , n381747 , n381749 );
nand ( n381751 , n381712 , RI15b50a90_617);
and ( n381752 , n381746 , n381750 , n381751 );
nor ( n381753 , n381745 , n381752 );
buf ( n381754 , n381753 );
not ( n381755 , n381754 );
or ( n381756 , n381727 , n381755 );
or ( n381757 , n381754 , n381726 );
nand ( n381758 , n381756 , n381757 );
and ( n381759 , n381758 , n21563 );
nor ( n381760 , n21750 , n22838 );
nor ( n381761 , n381759 , n381760 );
not ( n381762 , n20696 );
not ( n381763 , n20708 );
not ( n381764 , n21311 );
nand ( n381765 , n381762 , n381763 , n381764 , n21318 );
and ( n381766 , n20692 , RI15b50a18_616);
or ( n381767 , n20692 , n381731 );
nand ( n381768 , n381767 , n381734 );
nor ( n381769 , n381766 , n381768 );
nand ( n381770 , n20692 , RI15b509a0_615);
nand ( n381771 , n20691 , n381738 );
nand ( n381772 , n381770 , n381771 , n381741 );
not ( n381773 , n381772 );
nor ( n381774 , n381765 , n381769 , n381773 , n21329 );
and ( n381775 , n21302 , n381774 );
or ( n381776 , n20692 , n381748 );
nand ( n381777 , n20692 , RI15b50a90_617);
nand ( n381778 , n381776 , n381777 , n381751 );
nand ( n381779 , n381775 , n381778 );
buf ( n381780 , n381779 );
and ( n381781 , n20692 , RI15b50b08_618);
or ( n381782 , n20692 , n381716 );
nand ( n381783 , n381782 , n381725 );
nor ( n381784 , n381781 , n381783 );
and ( n381785 , n381780 , n381784 );
not ( n381786 , n381780 );
not ( n381787 , n381784 );
and ( n381788 , n381786 , n381787 );
nor ( n381789 , n381785 , n381788 );
buf ( n381790 , n21357 );
nand ( n381791 , n381789 , n381790 );
not ( n381792 , n21728 );
and ( n381793 , n381792 , RI15b509a0_615);
buf ( n381794 , n21727 );
not ( n381795 , n381738 );
or ( n381796 , n381794 , n381795 );
nand ( n381797 , n381796 , n381741 );
nor ( n381798 , n381793 , n381797 );
nand ( n381799 , n21737 , n381798 );
and ( n381800 , n381794 , RI15b50a18_616);
or ( n381801 , n21729 , n381731 );
nand ( n381802 , n381801 , n381734 );
nor ( n381803 , n381800 , n381802 );
not ( n381804 , n381803 );
nor ( n381805 , n381799 , n381804 );
buf ( n381806 , n381794 );
and ( n381807 , n381806 , RI15b50a90_617);
or ( n381808 , n381792 , n381748 );
nand ( n381809 , n381808 , n381751 );
nor ( n381810 , n381807 , n381809 );
nand ( n381811 , n381805 , n381810 );
not ( n381812 , n381811 );
and ( n381813 , n381806 , RI15b50b08_618);
or ( n381814 , n381792 , n381716 );
nand ( n381815 , n381814 , n381725 );
nor ( n381816 , n381813 , n381815 );
nor ( n381817 , n381812 , n381816 );
not ( n381818 , n381817 );
not ( n381819 , n381816 );
nor ( n381820 , n381811 , n381819 );
buf ( n381821 , n381820 );
not ( n381822 , n381821 );
nand ( n381823 , n381818 , n381822 );
nand ( n381824 , n381823 , n21747 );
and ( n381825 , n381761 , n381791 , n381824 );
not ( n381826 , n22537 );
and ( n381827 , n381826 , n21770 );
not ( n381828 , n21795 );
or ( n381829 , n381828 , n17517 , RI15b572a0_839);
and ( n381830 , n22704 , n17517 );
nor ( n381831 , n381830 , n21791 );
or ( n381832 , n381831 , n17518 );
nand ( n381833 , n381829 , n381832 );
nor ( n381834 , n381827 , n381833 );
nand ( n381835 , n381825 , n381834 );
buf ( n381836 , n381835 );
buf ( n381837 , n19655 );
buf ( n381838 , n22009 );
not ( n381839 , n21879 );
nor ( n381840 , n381839 , n21885 );
and ( n381841 , n21802 , n381840 );
buf ( n381842 , n21935 );
or ( n381843 , n21922 , n381842 );
nand ( n381844 , n381843 , n21946 );
and ( n381845 , n381844 , RI15b57c00_859);
buf ( n381846 , n21966 );
not ( n381847 , n381846 );
not ( n381848 , n21949 );
or ( n381849 , n381847 , n381848 );
nand ( n381850 , n381849 , n21979 );
and ( n381851 , n381850 , RI15b55e00_795);
or ( n381852 , n21982 , n381846 , RI15b55e00_795);
and ( n381853 , n381842 , n21937 , RI15b57b88_858);
and ( n381854 , n21936 , RI15b57c00_859);
nor ( n381855 , n381853 , n381854 );
or ( n381856 , n21922 , n381855 );
nand ( n381857 , n381852 , n381856 );
nor ( n381858 , n381845 , n381851 , n381857 );
or ( n381859 , n381858 , n18078 );
and ( n381860 , n18177 , RI15b57c00_859);
and ( n381861 , n18219 , RI15b56d00_827);
nor ( n381862 , n381860 , n381861 , n21751 );
nand ( n381863 , n381859 , n381862 );
nor ( n381864 , n381841 , n381863 );
nand ( n381865 , n381839 , n17507 );
not ( n381866 , n381865 );
not ( n381867 , n17565 );
or ( n381868 , n381866 , n381867 );
nand ( n381869 , n381868 , n21885 );
nand ( n381870 , n381864 , n381869 );
buf ( n381871 , n381870 );
buf ( n381872 , RI15b3ea48_2);
buf ( n381873 , n381872 );
buf ( n381874 , n381707 );
buf ( n381875 , n22343 );
or ( n381876 , n380968 , n22151 );
and ( n381877 , n380986 , n22211 );
not ( n381878 , RI15b408c0_67);
or ( n381879 , n22237 , n381878 );
or ( n381880 , n380994 , n22296 );
or ( n381881 , n22228 , n380996 );
nand ( n381882 , n381879 , n381880 , n381881 );
nor ( n381883 , n381877 , n381882 );
nand ( n381884 , n381876 , n381883 );
buf ( n381885 , n381884 );
not ( n381886 , RI15b66480_1355);
buf ( n381887 , n22066 );
not ( n381888 , n381887 );
not ( n381889 , n22067 );
and ( n381890 , n381888 , n381889 );
not ( n381891 , RI15b66408_1354);
nor ( n381892 , n381889 , n381891 );
nor ( n381893 , n381890 , n381892 );
not ( n381894 , RI15b66408_1354);
nand ( n381895 , n381887 , n381894 );
nand ( n381896 , n381893 , n381895 );
not ( n381897 , n381896 );
or ( n381898 , n381886 , n381897 );
not ( n381899 , n381888 );
not ( n381900 , n381889 );
nor ( n381901 , n381900 , n22055 );
nand ( n381902 , n381899 , n381901 );
nand ( n381903 , n381898 , n381902 );
and ( n381904 , n381903 , n22097 );
nor ( n381905 , n22094 , n22054 );
nor ( n381906 , n381904 , n381905 );
buf ( n381907 , n381906 );
or ( n381908 , n381907 , n22151 );
not ( n381909 , n22237 );
and ( n381910 , n381909 , RI15b40758_64);
buf ( n381911 , n22176 );
or ( n381912 , n381911 , n20638 );
nand ( n381913 , n381912 , n22094 );
not ( n381914 , n22184 );
nand ( n381915 , n381913 , n381914 );
nand ( n381916 , n22184 , n381911 , n22097 );
and ( n381917 , n381915 , n381916 );
or ( n381918 , n381917 , n22213 );
not ( n381919 , n22296 );
and ( n381920 , n22287 , n22283 );
not ( n381921 , n22287 );
and ( n381922 , n381921 , RI15b65940_1331);
or ( n381923 , n381920 , n381922 );
and ( n381924 , n381919 , n381923 );
not ( n381925 , n22298 );
and ( n381926 , n20116 , n381925 );
and ( n381927 , n381926 , n22294 );
nor ( n381928 , n381924 , n381927 );
nand ( n381929 , n381918 , n381928 );
nor ( n381930 , n381910 , n381929 );
nand ( n381931 , n381908 , n381930 );
buf ( n381932 , n381931 );
buf ( n381933 , n379802 );
buf ( n381934 , n379893 );
not ( n381935 , RI15b46e00_283);
not ( n381936 , n379832 );
or ( n381937 , n381935 , n381936 );
nor ( n381938 , RI15b48480_331 , RI15b486d8_336);
nor ( n381939 , RI15b48570_333 , RI15b48750_337);
nand ( n381940 , n381938 , n381939 );
nor ( n381941 , RI15b488b8_340 , RI15b48a20_343);
nor ( n381942 , RI15b48930_341 , RI15b48a98_344);
nand ( n381943 , n381941 , n381942 );
nor ( n381944 , n381940 , n381943 );
nor ( n381945 , RI15b484f8_332 , RI15b48660_335);
nor ( n381946 , RI15b485e8_334 , RI15b48840_339);
nand ( n381947 , n381945 , n381946 );
not ( n381948 , RI15b487c8_338);
not ( n381949 , RI15b489a8_342);
not ( n381950 , RI15b48b10_345);
nand ( n381951 , n381948 , n381949 , n381950 );
nor ( n381952 , n381947 , n381951 );
nand ( n381953 , n381944 , n381952 );
not ( n381954 , RI15b49308_362);
nor ( n381955 , n381953 , n381954 );
not ( n381956 , n381947 );
nor ( n381957 , RI15b487c8_338 , RI15b489a8_342);
nand ( n381958 , n381944 , n381956 , n381957 , RI15b49308_362);
or ( n381959 , n381955 , n381958 );
or ( n381960 , n381955 , RI15b48b10_345);
nand ( n381961 , n381960 , n381958 );
nand ( n381962 , n381959 , n381961 );
and ( n381963 , n379825 , n381962 );
not ( n381964 , n22031 );
and ( n381965 , n381964 , RI15b65e68_1342);
buf ( n381966 , n22033 );
not ( n381967 , n381966 );
nor ( n381968 , n381965 , n381967 );
not ( n381969 , n381968 );
not ( n381970 , n22027 );
nand ( n381971 , n381970 , RI15b666d8_1360);
and ( n381972 , n381971 , n22028 );
not ( n381973 , n381971 );
and ( n381974 , n381973 , RI15b65d00_1339);
nor ( n381975 , n381972 , n381974 );
and ( n381976 , RI15b666d8_1360 , n381975 );
not ( n381977 , RI15b666d8_1360);
not ( n381978 , n381975 );
and ( n381979 , n381977 , n381978 );
nor ( n381980 , n381976 , n381979 );
not ( n381981 , n381980 );
buf ( n381982 , n22026 );
nand ( n381983 , n381982 , RI15b666d8_1360);
not ( n381984 , n381983 );
not ( n381985 , RI15b65c88_1338);
and ( n381986 , n381984 , n381985 );
and ( n381987 , n381983 , RI15b65c88_1338);
nor ( n381988 , n381986 , n381987 );
not ( n381989 , n381988 );
not ( n381990 , RI15b666d8_1360);
and ( n381991 , n381989 , n381990 );
and ( n381992 , n381988 , RI15b666d8_1360);
nor ( n381993 , n381991 , n381992 );
not ( n381994 , n381993 );
not ( n381995 , n22024 );
nand ( n381996 , n381995 , RI15b666d8_1360);
and ( n381997 , n381996 , n22025 );
not ( n381998 , n381996 );
and ( n381999 , n381998 , RI15b65c10_1337);
or ( n382000 , n381997 , n381999 );
and ( n382001 , n382000 , n22286 , RI15b666d8_1360);
nand ( n382002 , n381994 , n382001 );
nor ( n382003 , n381981 , n382002 );
not ( n382004 , RI15b666d8_1360);
nor ( n382005 , n381970 , RI15b65d00_1339);
not ( n382006 , n382005 );
nand ( n382007 , n382006 , RI15b666d8_1360);
not ( n382008 , n382007 );
not ( n382009 , RI15b65d78_1340);
and ( n382010 , n382008 , n382009 );
and ( n382011 , n382007 , RI15b65d78_1340);
nor ( n382012 , n382010 , n382011 );
not ( n382013 , n382012 );
or ( n382014 , n382004 , n382013 );
or ( n382015 , n382012 , RI15b666d8_1360);
nand ( n382016 , n382014 , n382015 );
nand ( n382017 , n382003 , n382016 );
not ( n382018 , n382017 );
nand ( n382019 , n382005 , n22029 );
nand ( n382020 , n382019 , RI15b666d8_1360);
not ( n382021 , n382020 );
not ( n382022 , RI15b65df0_1341);
and ( n382023 , n382021 , n382022 );
and ( n382024 , n382020 , RI15b65df0_1341);
nor ( n382025 , n382023 , n382024 );
not ( n382026 , n382025 );
and ( n382027 , RI15b666d8_1360 , n382026 );
not ( n382028 , RI15b666d8_1360);
and ( n382029 , n382028 , n382025 );
nor ( n382030 , n382027 , n382029 );
and ( n382031 , n382018 , n382030 );
nand ( n382032 , n381969 , n382031 );
nand ( n382033 , n379816 , n382032 );
not ( n382034 , n382033 );
not ( n382035 , RI15b65ee0_1343);
nand ( n382036 , n381966 , RI15b666d8_1360);
not ( n382037 , n382036 );
or ( n382038 , n382035 , n382037 );
or ( n382039 , n382036 , RI15b65ee0_1343);
nand ( n382040 , n382038 , n382039 );
or ( n382041 , n382034 , n382040 );
nand ( n382042 , n382041 , n379820 );
and ( n382043 , n382034 , n382040 );
nor ( n382044 , n382042 , n382043 );
nor ( n382045 , n381963 , n382044 );
nand ( n382046 , n381937 , n382045 );
buf ( n382047 , n382046 );
buf ( n382048 , n381872 );
buf ( n382049 , RI15b3e9d0_1);
buf ( n382050 , n382049 );
buf ( n382051 , n381006 );
buf ( n382052 , RI15b3ea48_2);
buf ( n382053 , n382052 );
buf ( n382054 , n20663 );
buf ( n382055 , n382049 );
not ( n382056 , RI15b48228_326);
nor ( n382057 , RI15b47df0_317 , RI15b482a0_327);
nand ( n382058 , n382056 , n382057 );
or ( n382059 , n382058 , RI15b4b180_427);
and ( n382060 , RI15b47df0_317 , RI15b48228_326);
nor ( n382061 , n382060 , RI15b482a0_327);
nand ( n382062 , n382061 , RI15b4b1f8_428);
nand ( n382063 , n382059 , n382062 );
buf ( n382064 , n382063 );
buf ( n382065 , RI15b3e9d0_1);
buf ( n382066 , n382065 );
buf ( n382067 , RI15b3ea48_2);
buf ( n382068 , n382067 );
buf ( n382069 , RI15b3e9d0_1);
buf ( n382070 , n382069 );
buf ( n382071 , RI15b3ea48_2);
buf ( n382072 , n382071 );
buf ( n382073 , RI15b3ea48_2);
buf ( n382074 , n382073 );
buf ( n382075 , n19655 );
not ( n382076 , RI15b48318_328);
nand ( n382077 , n382076 , RI15b48390_329);
not ( n382078 , RI15b48408_330);
or ( n382079 , n382077 , n382078 );
not ( n382080 , n382079 );
not ( n382081 , n382080 );
nor ( n382082 , RI15b4b180_427 , RI15b4b1f8_428);
not ( n382083 , RI15b4b270_429);
and ( n382084 , n382082 , n382083 );
buf ( n382085 , n382084 );
not ( n382086 , RI15b4b2e8_430);
nand ( n382087 , n382085 , n382086 );
not ( n382088 , n382087 );
and ( n382089 , RI15b4b360_431 , n382088 );
not ( n382090 , n382089 );
nand ( n382091 , n382087 , RI15b4c008_458);
nor ( n382092 , n382091 , RI15b4b360_431);
not ( n382093 , n382092 );
nand ( n382094 , n382090 , n382093 );
not ( n382095 , n382094 );
nor ( n382096 , RI15b4b2e8_430 , RI15b4b360_431);
and ( n382097 , n382084 , n382096 );
nor ( n382098 , RI15b4b3d8_432 , RI15b4b450_433);
not ( n382099 , RI15b4b4c8_434);
and ( n382100 , n382098 , n382099 );
not ( n382101 , RI15b4b540_435);
nand ( n382102 , n382100 , n382101 );
nor ( n382103 , n382102 , RI15b4b5b8_436);
nand ( n382104 , n382097 , n382103 );
not ( n382105 , RI15b4b630_437);
not ( n382106 , RI15b4b6a8_438);
nand ( n382107 , n382105 , n382106 );
nor ( n382108 , n382104 , n382107 );
not ( n382109 , RI15b4b720_439);
not ( n382110 , RI15b4b798_440);
and ( n382111 , n382109 , n20547 , n382110 );
nand ( n382112 , n382108 , n382111 );
nor ( n382113 , n382112 , RI15b4b888_442);
not ( n382114 , RI15b4b900_443);
not ( n382115 , RI15b4b978_444);
and ( n382116 , n382114 , n382115 );
not ( n382117 , RI15b4b9f0_445);
nand ( n382118 , n382113 , n382116 , n382117 );
not ( n382119 , RI15b4ba68_446);
not ( n382120 , RI15b4bae0_447);
and ( n382121 , n382119 , n382120 );
not ( n382122 , RI15b4bb58_448);
nand ( n382123 , n382121 , n382122 );
nor ( n382124 , n382118 , n382123 );
not ( n382125 , RI15b4bbd0_449);
not ( n382126 , RI15b4bc48_450);
nand ( n382127 , n382125 , n382126 );
nor ( n382128 , n382127 , RI15b4bcc0_451);
and ( n382129 , n382124 , n382128 );
not ( n382130 , RI15b4bd38_452);
nand ( n382131 , n382129 , n382130 );
nand ( n382132 , n382131 , RI15b4c008_458);
not ( n382133 , n382132 );
not ( n382134 , n382133 );
not ( n382135 , RI15b4bdb0_453);
not ( n382136 , n382135 );
and ( n382137 , n382134 , n382136 );
not ( n382138 , n382132 );
and ( n382139 , n382138 , n382135 );
nor ( n382140 , n382137 , n382139 );
not ( n382141 , n382131 );
not ( n382142 , n382141 );
not ( n382143 , RI15b4be28_454);
nand ( n382144 , n382135 , n382143 );
nor ( n382145 , n382142 , n382144 );
nand ( n382146 , n382145 , n380888 );
not ( n382147 , n382131 );
nand ( n382148 , n382147 , n382135 );
not ( n382149 , RI15b4c008_458);
nor ( n382150 , n382149 , RI15b4be28_454);
and ( n382151 , n382148 , n382150 );
not ( n382152 , n382148 );
and ( n382153 , n382152 , RI15b4be28_454);
nor ( n382154 , n382151 , n382153 );
nand ( n382155 , RI15b4b180_427 , RI15b4c008_458);
and ( n382156 , n382155 , RI15b4b1f8_428);
not ( n382157 , n382155 );
not ( n382158 , RI15b4b1f8_428);
and ( n382159 , n382157 , n382158 );
nor ( n382160 , n382156 , n382159 );
and ( n382161 , n382140 , n382146 , n382154 , n382160 );
not ( n382162 , RI15b4bea0_455);
not ( n382163 , n382145 );
or ( n382164 , n382162 , n382163 );
or ( n382165 , n382145 , RI15b4bea0_455);
nand ( n382166 , n382164 , n382165 );
nor ( n382167 , n382144 , RI15b4bea0_455);
not ( n382168 , n382167 );
not ( n382169 , n382132 );
or ( n382170 , n382168 , n382169 );
nand ( n382171 , n382170 , n380886 );
not ( n382172 , n382129 );
nand ( n382173 , n382130 , RI15b4c008_458);
not ( n382174 , n382173 );
and ( n382175 , n382172 , n382174 );
and ( n382176 , n382129 , RI15b4bd38_452);
nor ( n382177 , n382175 , n382176 );
not ( n382178 , n382127 );
not ( n382179 , n382178 );
not ( n382180 , n382124 );
not ( n382181 , n382180 );
not ( n382182 , n382181 );
or ( n382183 , n382179 , n382182 );
nand ( n382184 , n382183 , RI15b4c008_458);
and ( n382185 , RI15b4bcc0_451 , n382184 );
not ( n382186 , RI15b4bcc0_451);
not ( n382187 , RI15b4c008_458);
not ( n382188 , n382127 );
or ( n382189 , n382187 , n382188 );
nand ( n382190 , n382180 , RI15b4c008_458);
nand ( n382191 , n382189 , n382190 );
and ( n382192 , n382186 , n382191 );
nor ( n382193 , n382185 , n382192 );
not ( n382194 , RI15b4c008_458);
nand ( n382195 , n382194 , RI15b4bd38_452);
nand ( n382196 , n382177 , n382193 , n382195 );
nor ( n382197 , n382196 , n20643 );
nand ( n382198 , n382171 , n382197 );
nor ( n382199 , n382166 , n382198 );
not ( n382200 , RI15b4c008_458);
not ( n382201 , n382144 );
nand ( n382202 , n382141 , n382201 );
not ( n382203 , n382202 );
or ( n382204 , n382200 , n382203 );
nor ( n382205 , RI15b4bea0_455 , RI15b4bf18_456);
nand ( n382206 , n382204 , n382205 );
and ( n382207 , n382206 , n20643 );
nand ( n382208 , n382205 , RI15b4bf90_457);
nor ( n382209 , n382202 , n382208 );
nor ( n382210 , n382207 , n382209 );
buf ( n382211 , n382100 );
not ( n382212 , n382211 );
and ( n382213 , n382084 , n382096 );
not ( n382214 , n382213 );
or ( n382215 , n382212 , n382214 );
nand ( n382216 , n382215 , RI15b4c008_458);
and ( n382217 , RI15b4b540_435 , n382216 );
not ( n382218 , RI15b4b540_435);
not ( n382219 , RI15b4c008_458);
not ( n382220 , n382211 );
not ( n382221 , n382220 );
or ( n382222 , n382219 , n382221 );
not ( n382223 , n382097 );
nand ( n382224 , n382223 , RI15b4c008_458);
nand ( n382225 , n382222 , n382224 );
and ( n382226 , n382218 , n382225 );
nor ( n382227 , n382217 , n382226 );
not ( n382228 , n382102 );
not ( n382229 , n382228 );
not ( n382230 , n382213 );
or ( n382231 , n382229 , n382230 );
nand ( n382232 , n382231 , RI15b4c008_458);
and ( n382233 , RI15b4b5b8_436 , n382232 );
not ( n382234 , RI15b4b5b8_436);
not ( n382235 , RI15b4c008_458);
not ( n382236 , n382102 );
or ( n382237 , n382235 , n382236 );
nand ( n382238 , n382237 , n382224 );
and ( n382239 , n382234 , n382238 );
nor ( n382240 , n382233 , n382239 );
nand ( n382241 , n382227 , n382240 );
not ( n382242 , n382241 );
not ( n382243 , n382213 );
not ( n382244 , n382098 );
or ( n382245 , n382243 , n382244 );
nand ( n382246 , n382245 , RI15b4c008_458);
and ( n382247 , RI15b4b4c8_434 , n382246 );
not ( n382248 , RI15b4b4c8_434);
nor ( n382249 , n382244 , RI15b4b360_431);
nand ( n382250 , n382091 , n382249 );
and ( n382251 , n382248 , n382250 );
nor ( n382252 , n382247 , n382251 );
not ( n382253 , RI15b4b3d8_432);
not ( n382254 , n382253 );
not ( n382255 , n382097 );
or ( n382256 , n382254 , n382255 );
nand ( n382257 , n382256 , RI15b4c008_458);
and ( n382258 , n382257 , RI15b4b450_433);
not ( n382259 , n382257 );
and ( n382260 , n382259 , n22374 );
nor ( n382261 , n382258 , n382260 );
nand ( n382262 , n382252 , n382261 );
not ( n382263 , n382092 );
not ( n382264 , n382213 );
nand ( n382265 , n382253 , RI15b4c008_458);
not ( n382266 , n382265 );
and ( n382267 , n382264 , n382266 );
and ( n382268 , n382213 , RI15b4b3d8_432);
nor ( n382269 , n382267 , n382268 );
not ( n382270 , n382085 );
or ( n382271 , n382270 , n382086 );
or ( n382272 , n382086 , RI15b4c008_458);
nand ( n382273 , n382271 , n382272 );
nand ( n382274 , n382086 , RI15b4c008_458);
nor ( n382275 , n382085 , n382274 );
nor ( n382276 , n382273 , n382275 );
buf ( n382277 , n382082 );
not ( n382278 , RI15b4c008_458);
nor ( n382279 , n382277 , n382278 );
not ( n382280 , RI15b4b270_429);
and ( n382281 , n382279 , n382280 );
not ( n382282 , n382279 );
and ( n382283 , n382282 , RI15b4b270_429);
nor ( n382284 , n382281 , n382283 );
and ( n382285 , n382276 , n382284 );
nand ( n382286 , n382091 , RI15b4b360_431);
nand ( n382287 , n382263 , n382269 , n382285 , n382286 );
nor ( n382288 , n382262 , n382287 );
nand ( n382289 , n382242 , n382288 );
nand ( n382290 , n382104 , RI15b4c008_458);
not ( n382291 , n382290 );
not ( n382292 , RI15b4b630_437);
and ( n382293 , n382291 , n382292 );
and ( n382294 , n382290 , RI15b4b630_437);
nor ( n382295 , n382293 , n382294 );
not ( n382296 , n382104 );
not ( n382297 , RI15b4b630_437);
nand ( n382298 , n382296 , n382297 );
and ( n382299 , n382106 , RI15b4c008_458);
and ( n382300 , n382298 , n382299 );
not ( n382301 , n382298 );
and ( n382302 , n382301 , RI15b4b6a8_438);
nor ( n382303 , n382300 , n382302 );
nand ( n382304 , n382295 , n382303 );
nor ( n382305 , n382289 , n382304 );
not ( n382306 , RI15b4c008_458);
nor ( n382307 , n382107 , RI15b4b720_439);
nand ( n382308 , n382307 , n382110 );
not ( n382309 , n382308 );
or ( n382310 , n382306 , n382309 );
nand ( n382311 , n382310 , n382290 );
not ( n382312 , n382311 );
not ( n382313 , n20547 );
and ( n382314 , n382312 , n382313 );
and ( n382315 , n382311 , n20547 );
nor ( n382316 , n382314 , n382315 );
not ( n382317 , n382108 );
and ( n382318 , n382109 , RI15b4c008_458);
and ( n382319 , n382317 , n382318 );
not ( n382320 , n382317 );
and ( n382321 , n382320 , RI15b4b720_439);
nor ( n382322 , n382319 , n382321 );
nand ( n382323 , n382316 , n382322 );
not ( n382324 , RI15b4b798_440);
not ( n382325 , n382109 );
not ( n382326 , n382108 );
or ( n382327 , n382325 , n382326 );
nand ( n382328 , n382327 , RI15b4c008_458);
not ( n382329 , n382328 );
or ( n382330 , n382324 , n382329 );
not ( n382331 , n382307 );
not ( n382332 , n382290 );
or ( n382333 , n382331 , n382332 );
nand ( n382334 , n382333 , n382110 );
nand ( n382335 , n382330 , n382334 );
nor ( n382336 , n382323 , n382335 );
and ( n382337 , n382305 , n382336 );
buf ( n382338 , n382112 );
and ( n382339 , n20546 , RI15b4c008_458);
and ( n382340 , n382338 , n382339 );
not ( n382341 , n382338 );
and ( n382342 , n382341 , RI15b4b888_442);
nor ( n382343 , n382340 , n382342 );
not ( n382344 , RI15b4c008_458);
nand ( n382345 , n382344 , RI15b4b888_442);
and ( n382346 , n382343 , n382345 );
nand ( n382347 , n382337 , n382346 );
buf ( n382348 , n382113 );
nand ( n382349 , n382348 , n382116 );
nand ( n382350 , n382349 , RI15b4c008_458);
and ( n382351 , RI15b4b9f0_445 , n382350 );
not ( n382352 , RI15b4b9f0_445);
not ( n382353 , RI15b4c008_458);
not ( n382354 , n382116 );
not ( n382355 , n382354 );
or ( n382356 , n382353 , n382355 );
not ( n382357 , n382113 );
nand ( n382358 , n382357 , RI15b4c008_458);
nand ( n382359 , n382356 , n382358 );
and ( n382360 , n382352 , n382359 );
nor ( n382361 , n382351 , n382360 );
not ( n382362 , RI15b4b900_443);
not ( n382363 , n382358 );
or ( n382364 , n382362 , n382363 );
or ( n382365 , n382358 , RI15b4b900_443);
nand ( n382366 , n382364 , n382365 );
not ( n382367 , RI15b4b978_444);
not ( n382368 , n382114 );
not ( n382369 , n382113 );
or ( n382370 , n382368 , n382369 );
nand ( n382371 , n382370 , RI15b4c008_458);
not ( n382372 , n382371 );
or ( n382373 , n382367 , n382372 );
or ( n382374 , n382371 , RI15b4b978_444);
nand ( n382375 , n382373 , n382374 );
nor ( n382376 , n382366 , n382375 );
nand ( n382377 , n382361 , n382376 );
nor ( n382378 , n382347 , n382377 );
not ( n382379 , n382118 );
not ( n382380 , n382379 );
nand ( n382381 , n382380 , RI15b4c008_458);
and ( n382382 , RI15b4ba68_446 , n382381 );
not ( n382383 , RI15b4ba68_446);
not ( n382384 , RI15b4c008_458);
nor ( n382385 , n382384 , n382117 );
nor ( n382386 , n382359 , n382385 );
not ( n382387 , n382386 );
and ( n382388 , n382383 , n382387 );
nor ( n382389 , n382382 , n382388 );
and ( n382390 , n382378 , n382389 );
not ( n382391 , n382121 );
not ( n382392 , n382379 );
or ( n382393 , n382391 , n382392 );
nand ( n382394 , n382393 , RI15b4c008_458);
and ( n382395 , RI15b4bb58_448 , n382394 );
not ( n382396 , RI15b4bb58_448);
not ( n382397 , RI15b4c008_458);
not ( n382398 , n382121 );
not ( n382399 , n382398 );
or ( n382400 , n382397 , n382399 );
nand ( n382401 , n382400 , n382386 );
and ( n382402 , n382396 , n382401 );
nor ( n382403 , n382395 , n382402 );
not ( n382404 , n382119 );
not ( n382405 , n382379 );
or ( n382406 , n382404 , n382405 );
nand ( n382407 , n382406 , RI15b4c008_458);
not ( n382408 , n382407 );
not ( n382409 , RI15b4bae0_447);
and ( n382410 , n382408 , n382409 );
and ( n382411 , n382407 , RI15b4bae0_447);
nor ( n382412 , n382410 , n382411 );
and ( n382413 , n382403 , n382412 );
nand ( n382414 , n382390 , n382413 );
not ( n382415 , RI15b4bbd0_449);
buf ( n382416 , n382190 );
not ( n382417 , n382416 );
or ( n382418 , n382415 , n382417 );
or ( n382419 , n382416 , RI15b4bbd0_449);
nand ( n382420 , n382418 , n382419 );
nor ( n382421 , n382414 , n382420 );
not ( n382422 , n382125 );
not ( n382423 , n382181 );
or ( n382424 , n382422 , n382423 );
nand ( n382425 , n382424 , RI15b4c008_458);
not ( n382426 , n382425 );
not ( n382427 , RI15b4bc48_450);
and ( n382428 , n382426 , n382427 );
and ( n382429 , n382425 , RI15b4bc48_450);
nor ( n382430 , n382428 , n382429 );
and ( n382431 , n382421 , n382430 );
nand ( n382432 , n382161 , n382199 , n382210 , n382431 );
nand ( n382433 , n382432 , RI15b4c008_458);
not ( n382434 , n382433 );
not ( n382435 , n382434 );
or ( n382436 , n382095 , n382435 );
not ( n382437 , RI15b4c008_458);
nand ( n382438 , n382437 , RI15b4b360_431);
nand ( n382439 , n382436 , n382438 );
buf ( n382440 , n382432 );
buf ( n382441 , n382276 );
not ( n382442 , RI15b4c008_458);
nor ( n382443 , n382441 , n382442 );
and ( n382444 , n382440 , n382443 );
not ( n382445 , n382272 );
nor ( n382446 , n382444 , n382445 );
and ( n382447 , n382284 , n382160 );
nand ( n382448 , n382446 , n382447 );
nor ( n382449 , n382439 , n382448 );
not ( n382450 , n382269 );
not ( n382451 , n382450 );
not ( n382452 , n382434 );
or ( n382453 , n382451 , n382452 );
not ( n382454 , RI15b4c008_458);
nand ( n382455 , n382454 , RI15b4b3d8_432);
nand ( n382456 , n382453 , n382455 );
not ( n382457 , n382456 );
nand ( n382458 , n382449 , n382457 );
not ( n382459 , n382434 );
not ( n382460 , n382459 );
not ( n382461 , n382261 );
and ( n382462 , n382460 , n382461 );
not ( n382463 , RI15b4c008_458);
and ( n382464 , n382463 , RI15b4b450_433);
nor ( n382465 , n382462 , n382464 );
not ( n382466 , n382465 );
nor ( n382467 , n382458 , n382466 );
buf ( n382468 , n382467 );
not ( n382469 , n382468 );
or ( n382470 , n382081 , n382469 );
buf ( n382471 , n382434 );
not ( n382472 , n382471 );
buf ( n382473 , n382472 );
nand ( n382474 , n382473 , n382080 );
not ( n382475 , n382474 );
not ( n382476 , n382475 );
nand ( n382477 , n382470 , n382476 );
not ( n382478 , n382252 );
not ( n382479 , n382478 );
not ( n382480 , n382434 );
or ( n382481 , n382479 , n382480 );
not ( n382482 , RI15b4c008_458);
nand ( n382483 , n382482 , RI15b4b4c8_434);
nand ( n382484 , n382481 , n382483 );
nand ( n382485 , n382477 , n382484 );
not ( n382486 , n382473 );
nand ( n382487 , n382486 , n382080 );
not ( n382488 , n382487 );
not ( n382489 , n382484 );
nand ( n382490 , n382488 , n382489 );
nor ( n382491 , n382468 , n382490 );
buf ( n382492 , n382210 );
and ( n382493 , n382492 , RI15b4bf90_457);
not ( n382494 , n382493 );
not ( n382495 , n382431 );
buf ( n382496 , n382196 );
nor ( n382497 , n382495 , n382496 );
buf ( n382498 , n382140 );
nand ( n382499 , n382497 , n382498 );
buf ( n382500 , n382154 );
not ( n382501 , n382500 );
nor ( n382502 , n382499 , n382501 );
not ( n382503 , n382166 );
and ( n382504 , n382502 , n382503 );
and ( n382505 , n382171 , n382146 );
and ( n382506 , n382504 , n382505 );
not ( n382507 , n382506 );
or ( n382508 , n382494 , n382507 );
and ( n382509 , n382078 , RI15b48390_329);
and ( n382510 , n382509 , n382076 );
and ( n382511 , n382510 , RI15b4c008_458);
nand ( n382512 , n382508 , n382511 );
buf ( n382513 , n382512 );
not ( n382514 , n382288 );
not ( n382515 , n382227 );
buf ( n382516 , n382515 );
not ( n382517 , n382516 );
and ( n382518 , n382514 , n382517 );
nor ( n382519 , n382514 , n382517 );
nor ( n382520 , n382518 , n382519 );
or ( n382521 , n382513 , n382520 );
not ( n382522 , RI15b4c008_458);
and ( n382523 , n382510 , n382522 );
and ( n382524 , n382523 , RI15b4b540_435);
buf ( n382525 , n382077 );
buf ( n382526 , n382525 );
buf ( n382527 , n382526 );
buf ( n382528 , n382527 );
buf ( n382529 , n382528 );
and ( n382530 , n382529 , RI15b45348_226);
nor ( n382531 , n382524 , n382530 );
nand ( n382532 , n382521 , n382531 );
nor ( n382533 , n382491 , n382532 );
nand ( n382534 , n382485 , n382533 );
buf ( n382535 , n382534 );
buf ( n382536 , n19653 );
buf ( n382537 , RI15b3e9d0_1);
buf ( n382538 , n382537 );
or ( n382539 , n18130 , n21349 );
buf ( n382540 , n21555 );
not ( n382541 , n382540 );
buf ( n382542 , n382541 );
not ( n382543 , n382542 );
or ( n382544 , n18120 , n382543 );
or ( n382545 , n18143 , n18072 );
not ( n382546 , n18096 );
nand ( n382547 , n18142 , n382546 );
nand ( n382548 , n382545 , n382547 );
nand ( n382549 , n382548 , n21977 , RI15b4c080_459);
nand ( n382550 , n382539 , n382544 , n382549 );
and ( n382551 , n382550 , n18077 );
and ( n382552 , n18078 , RI15b4c080_459);
nor ( n382553 , n382551 , n382552 );
not ( n382554 , n382553 );
buf ( n382555 , n382554 );
buf ( n382556 , n19655 );
buf ( n382557 , n382073 );
not ( n382558 , n18749 );
and ( n382559 , n18442 , n382558 );
not ( n382560 , n18442 );
not ( n382561 , n18684 );
and ( n382562 , n382561 , n18748 );
not ( n382563 , n18745 );
nor ( n382564 , n382562 , n382563 );
and ( n382565 , n382560 , n382564 );
nor ( n382566 , n382559 , n382565 );
or ( n382567 , n382566 , n19284 );
xnor ( n382568 , n19360 , n19299 );
or ( n382569 , n382568 , n19389 );
not ( n382570 , n19500 );
not ( n382571 , n19444 );
not ( n382572 , n19458 );
not ( n382573 , n19435 );
or ( n382574 , n382572 , n382573 );
nand ( n382575 , n382574 , n19465 );
not ( n382576 , n382575 );
or ( n382577 , n382571 , n382576 );
not ( n382578 , n19470 );
nand ( n382579 , n382577 , n382578 );
and ( n382580 , n382579 , n19452 );
nor ( n382581 , n382580 , n19463 );
not ( n382582 , n19418 );
and ( n382583 , n382581 , n382582 );
not ( n382584 , n382581 );
and ( n382585 , n382584 , n19418 );
nor ( n382586 , n382583 , n382585 );
or ( n382587 , n382570 , n382586 );
nand ( n382588 , n382567 , n382569 , n382587 );
buf ( n382589 , n18752 );
not ( n382590 , n382589 );
and ( n382591 , n382588 , n382590 );
and ( n382592 , n19513 , RI15b63d20_1271);
nor ( n382593 , n382591 , n382592 );
not ( n382594 , n382566 );
or ( n382595 , n382594 , n19285 );
and ( n382596 , n382568 , n19390 );
and ( n382597 , n382586 , n19500 );
nor ( n382598 , n382596 , n382597 );
nand ( n382599 , n382595 , n382598 );
not ( n382600 , n382590 );
nand ( n382601 , n382599 , n382600 );
and ( n382602 , n382593 , n382601 );
and ( n382603 , n19608 , RI15b62e20_1239);
not ( n382604 , RI15b62e20_1239);
not ( n382605 , n382604 );
buf ( n382606 , n19615 );
nor ( n382607 , n382606 , n19620 );
not ( n382608 , n382607 );
or ( n382609 , n382605 , n382608 );
not ( n382610 , RI15b62e20_1239);
or ( n382611 , n382607 , n382610 );
nand ( n382612 , n382609 , n382611 );
and ( n382613 , n19630 , n382612 );
buf ( n382614 , n382606 );
not ( n382615 , RI15b62e20_1239);
and ( n382616 , n382614 , n382615 );
not ( n382617 , n382614 );
and ( n382618 , n382617 , RI15b62e20_1239);
nor ( n382619 , n382616 , n382618 );
and ( n382620 , n380237 , n382619 );
nor ( n382621 , n382603 , n382613 , n382620 );
nand ( n382622 , n382602 , n382621 );
buf ( n382623 , n382622 );
buf ( n382624 , n379997 );
not ( n382625 , n382624 );
not ( n382626 , n382625 );
buf ( n382627 , n382626 );
not ( n382628 , n382627 );
buf ( n382629 , n382628 );
not ( n382630 , n382629 );
not ( n382631 , n382630 );
nand ( n382632 , RI15b548e8_750 , RI15b54960_751);
not ( n382633 , RI15b549d8_752);
nor ( n382634 , n382632 , n382633 );
and ( n382635 , RI15b54a50_753 , RI15b54ac8_754);
nand ( n382636 , n382634 , n382635 );
not ( n382637 , RI15b54b40_755);
nor ( n382638 , n382636 , n382637 );
nand ( n382639 , n382638 , RI15b54bb8_756);
not ( n382640 , n382639 );
and ( n382641 , RI15b54c30_757 , RI15b54ca8_758);
nand ( n382642 , n382640 , n382641 );
not ( n382643 , RI15b54d20_759);
nor ( n382644 , n382642 , n382643 );
nand ( n382645 , n382644 , RI15b54d98_760);
not ( n382646 , RI15b54e10_761);
nor ( n382647 , n382645 , n382646 );
and ( n382648 , n382647 , RI15b54e88_762);
and ( n382649 , n382648 , RI15b54f00_763);
nand ( n382650 , n382649 , RI15b54f78_764);
not ( n382651 , RI15b54ff0_765);
nor ( n382652 , n382650 , n382651 );
nand ( n382653 , n382652 , RI15b55068_766);
not ( n382654 , RI15b550e0_767);
nor ( n382655 , n382653 , n382654 );
nand ( n382656 , n382655 , RI15b55158_768);
not ( n382657 , RI15b551d0_769);
nor ( n382658 , n382656 , n382657 );
nand ( n382659 , n382658 , RI15b55248_770);
not ( n382660 , n382659 );
nand ( n382661 , n382660 , RI15b552c0_771);
not ( n382662 , RI15b55338_772);
nor ( n382663 , n382661 , n382662 );
and ( n382664 , n382663 , RI15b553b0_773);
not ( n382665 , RI15b554a0_775);
not ( n382666 , RI15b55428_774);
nor ( n382667 , n382665 , n382666 );
nand ( n382668 , n382664 , n382667 );
not ( n382669 , RI15b55518_776);
nor ( n382670 , n382668 , n382669 );
nand ( n382671 , n382670 , RI15b55590_777);
not ( n382672 , n382671 );
or ( n382673 , n382631 , n382672 );
nand ( n382674 , n379996 , n21557 );
nand ( n382675 , n382674 , n379989 , n379948 , n18077 );
nor ( n382676 , n379986 , n382675 );
not ( n382677 , n379993 );
nand ( n382678 , n382677 , n18181 );
and ( n382679 , n382676 , n382678 );
nand ( n382680 , n382673 , n382679 );
nor ( n382681 , n382628 , RI15b55608_778);
nor ( n382682 , n382680 , n382681 );
not ( n382683 , RI15b55680_779);
or ( n382684 , n382682 , n382683 );
not ( n382685 , n382671 );
not ( n382686 , RI15b55608_778);
nor ( n382687 , n382629 , n382686 );
and ( n382688 , n382685 , n382687 );
nand ( n382689 , n382688 , n382683 );
buf ( n382690 , n18137 );
or ( n382691 , n18181 , n381481 , n382690 );
not ( n382692 , n382691 );
buf ( n382693 , n381138 );
buf ( n382694 , n382693 );
not ( n382695 , n382694 );
not ( n382696 , n382695 );
not ( n382697 , n380965 );
and ( n382698 , n382696 , n382697 );
buf ( n382699 , n382693 );
not ( n382700 , n382699 );
and ( n382701 , n382700 , RI15b656e8_1326);
nor ( n382702 , n382698 , n382701 );
not ( n382703 , n382702 );
and ( n382704 , n382692 , n382703 );
not ( n382705 , n380193 );
nand ( n382706 , n382705 , n380087 );
not ( n382707 , n382706 );
buf ( n382708 , n380017 );
and ( n382709 , n382708 , RI15b4d3b8_500);
and ( n382710 , n381647 , RI15b4e2b8_532);
nor ( n382711 , n382709 , n382710 );
buf ( n382712 , n380029 );
and ( n382713 , n382712 , RI15b4def8_524);
buf ( n382714 , n380034 );
and ( n382715 , n382714 , RI15b4d778_508);
buf ( n382716 , n380038 );
and ( n382717 , n382716 , RI15b4e678_540);
nor ( n382718 , n382713 , n382715 , n382717 );
buf ( n382719 , n380043 );
and ( n382720 , n382719 , RI15b4ea38_548);
and ( n382721 , n381653 , RI15b4c878_476);
nor ( n382722 , n382720 , n382721 );
buf ( n382723 , n380052 );
and ( n382724 , n382723 , RI15b4edf8_556);
and ( n382725 , n379875 , RI15b4cff8_492);
nor ( n382726 , n382724 , n382725 );
and ( n382727 , n382711 , n382718 , n382722 , n382726 );
buf ( n382728 , n380059 );
and ( n382729 , n382728 , RI15b4cc38_484);
and ( n382730 , n380061 , RI15b4f1b8_564);
buf ( n382731 , n380065 );
and ( n382732 , n382731 , RI15b4c4b8_468);
nor ( n382733 , n382729 , n382730 , n382732 );
buf ( n382734 , n380071 );
and ( n382735 , n382734 , RI15b4db38_516);
buf ( n382736 , n380075 );
and ( n382737 , n382736 , RI15b4fcf8_588);
nor ( n382738 , n382735 , n382737 );
buf ( n382739 , n380080 );
and ( n382740 , n382739 , RI15b4f938_580);
buf ( n382741 , n380084 );
and ( n382742 , n382741 , RI15b4f578_572);
nor ( n382743 , n382740 , n382742 );
nand ( n382744 , n382727 , n382733 , n382738 , n382743 );
nand ( n382745 , n382707 , n382744 );
not ( n382746 , n382745 );
buf ( n382747 , n382708 );
and ( n382748 , n382747 , RI15b4d430_501);
and ( n382749 , n381648 , RI15b4e330_533);
nor ( n382750 , n382748 , n382749 );
buf ( n382751 , n382712 );
and ( n382752 , n382751 , RI15b4df70_525);
buf ( n382753 , n382714 );
and ( n382754 , n382753 , RI15b4d7f0_509);
buf ( n382755 , n382716 );
and ( n382756 , n382755 , RI15b4e6f0_541);
nor ( n382757 , n382752 , n382754 , n382756 );
buf ( n382758 , n382723 );
and ( n382759 , n382758 , RI15b4ee70_557);
and ( n382760 , n379876 , RI15b4d070_493);
nor ( n382761 , n382759 , n382760 );
buf ( n382762 , n382719 );
and ( n382763 , n382762 , RI15b4eab0_549);
and ( n382764 , n381654 , RI15b4c8f0_477);
nor ( n382765 , n382763 , n382764 );
nand ( n382766 , n382750 , n382757 , n382761 , n382765 );
not ( n382767 , n382766 );
buf ( n382768 , n382728 );
and ( n382769 , n382768 , RI15b4ccb0_485);
and ( n382770 , n380061 , RI15b4f230_565);
buf ( n382771 , n382731 );
and ( n382772 , n382771 , RI15b4c530_469);
nor ( n382773 , n382769 , n382770 , n382772 );
buf ( n382774 , n382739 );
and ( n382775 , n382774 , RI15b4f9b0_581);
buf ( n382776 , n382741 );
and ( n382777 , n382776 , RI15b4f5f0_573);
nor ( n382778 , n382775 , n382777 );
not ( n382779 , n382734 );
not ( n382780 , n382779 );
and ( n382781 , n382780 , RI15b4dbb0_517);
buf ( n382782 , n382736 );
and ( n382783 , n382782 , RI15b4fd70_589);
nor ( n382784 , n382781 , n382783 );
nand ( n382785 , n382767 , n382773 , n382778 , n382784 );
nand ( n382786 , n382746 , n382785 );
not ( n382787 , n382786 );
buf ( n382788 , n382747 );
and ( n382789 , n382788 , RI15b4d4a8_502);
and ( n382790 , n381650 , RI15b4e3a8_534);
nor ( n382791 , n382789 , n382790 );
not ( n382792 , n382751 );
not ( n382793 , n382792 );
and ( n382794 , n382793 , RI15b4dfe8_526);
buf ( n382795 , n382753 );
and ( n382796 , n382795 , RI15b4d868_510);
buf ( n382797 , n382755 );
and ( n382798 , n382797 , RI15b4e768_542);
nor ( n382799 , n382794 , n382796 , n382798 );
not ( n382800 , n382762 );
not ( n382801 , n382800 );
and ( n382802 , n382801 , RI15b4eb28_550);
buf ( n382803 , n381655 );
and ( n382804 , n382803 , RI15b4c968_478);
nor ( n382805 , n382802 , n382804 );
buf ( n382806 , n382758 );
and ( n382807 , n382806 , RI15b4eee8_558);
and ( n382808 , n379877 , RI15b4d0e8_494);
nor ( n382809 , n382807 , n382808 );
nand ( n382810 , n382791 , n382799 , n382805 , n382809 );
not ( n382811 , n382810 );
not ( n382812 , n382768 );
not ( n382813 , n382812 );
and ( n382814 , n382813 , RI15b4cd28_486);
and ( n382815 , n380061 , RI15b4f2a8_566);
buf ( n382816 , n382771 );
and ( n382817 , n382816 , RI15b4c5a8_470);
nor ( n382818 , n382814 , n382815 , n382817 );
buf ( n382819 , n382774 );
and ( n382820 , n382819 , RI15b4fa28_582);
buf ( n382821 , n382776 );
and ( n382822 , n382821 , RI15b4f668_574);
nor ( n382823 , n382820 , n382822 );
not ( n382824 , n382779 );
buf ( n382825 , n382824 );
buf ( n382826 , n382825 );
and ( n382827 , n382826 , RI15b4dc28_518);
buf ( n382828 , n382782 );
and ( n382829 , n382828 , RI15b4fde8_590);
nor ( n382830 , n382827 , n382829 );
nand ( n382831 , n382811 , n382818 , n382823 , n382830 );
nand ( n382832 , n382787 , n382831 );
not ( n382833 , n382832 );
buf ( n382834 , n382788 );
and ( n382835 , n382834 , RI15b4d520_503);
not ( n382836 , n381649 );
buf ( n382837 , n382836 );
buf ( n382838 , n382837 );
and ( n382839 , n382838 , RI15b4e420_535);
nor ( n382840 , n382835 , n382839 );
buf ( n382841 , n382793 );
buf ( n382842 , n382841 );
and ( n382843 , n382842 , RI15b4e060_527);
buf ( n382844 , n382795 );
and ( n382845 , n382844 , RI15b4d8e0_511);
buf ( n382846 , n382797 );
and ( n382847 , n382846 , RI15b4e7e0_543);
nor ( n382848 , n382843 , n382845 , n382847 );
buf ( n382849 , n382801 );
buf ( n382850 , n382849 );
and ( n382851 , n382850 , RI15b4eba0_551);
not ( n382852 , n381656 );
buf ( n382853 , n382852 );
and ( n382854 , n382853 , RI15b4c9e0_479);
nor ( n382855 , n382851 , n382854 );
buf ( n382856 , n382806 );
buf ( n382857 , n382856 );
and ( n382858 , n382857 , RI15b4ef60_559);
and ( n382859 , n379879 , RI15b4d160_495);
nor ( n382860 , n382858 , n382859 );
nand ( n382861 , n382840 , n382848 , n382855 , n382860 );
not ( n382862 , n382861 );
not ( n382863 , n382813 );
not ( n382864 , n382863 );
and ( n382865 , n382864 , RI15b4cda0_487);
and ( n382866 , n380061 , RI15b4f320_567);
buf ( n382867 , n382816 );
and ( n382868 , n382867 , RI15b4c620_471);
nor ( n382869 , n382865 , n382866 , n382868 );
buf ( n382870 , n382819 );
and ( n382871 , n382870 , RI15b4faa0_583);
buf ( n382872 , n382821 );
and ( n382873 , n382872 , RI15b4f6e0_575);
nor ( n382874 , n382871 , n382873 );
buf ( n382875 , n382826 );
and ( n382876 , n382875 , RI15b4dca0_519);
buf ( n382877 , n382828 );
and ( n382878 , n382877 , RI15b4fe60_591);
nor ( n382879 , n382876 , n382878 );
nand ( n382880 , n382862 , n382869 , n382874 , n382879 );
not ( n382881 , n382880 );
and ( n382882 , n382833 , n382881 );
and ( n382883 , n382832 , n382880 );
nor ( n382884 , n382882 , n382883 );
and ( n382885 , n379996 , n21556 );
not ( n382886 , n382885 );
nor ( n382887 , n382884 , n382886 );
buf ( n382888 , n381313 );
nor ( n382889 , n381400 , n382888 );
nor ( n382890 , n382704 , n382887 , n382889 );
nand ( n382891 , n382684 , n382689 , n382890 );
buf ( n382892 , n382891 );
buf ( n382893 , n380903 );
buf ( n382894 , n22343 );
not ( n382895 , n380229 );
not ( n382896 , n382895 );
not ( n382897 , n380725 );
and ( n382898 , n382896 , n382897 );
not ( n382899 , n382898 );
not ( n382900 , n381496 );
buf ( n382901 , n381574 );
not ( n382902 , n382901 );
or ( n382903 , n382900 , n382902 );
buf ( n382904 , n380685 );
nand ( n382905 , n382903 , n382904 );
not ( n382906 , n381576 );
not ( n382907 , n382906 );
and ( n382908 , n382905 , n382907 );
nand ( n382909 , n380698 , n382906 );
nor ( n382910 , n382909 , n382901 );
nor ( n382911 , n382908 , n382910 );
not ( n382912 , n382911 );
not ( n382913 , n382912 );
or ( n382914 , n382899 , n382913 );
buf ( n382915 , n380593 );
buf ( n382916 , n380506 );
nand ( n382917 , n382915 , n382916 );
not ( n382918 , n380512 );
nor ( n382919 , n382917 , n382918 );
buf ( n382920 , n380602 );
nand ( n382921 , n382919 , n382920 );
buf ( n382922 , n380581 );
not ( n382923 , n382922 );
nand ( n382924 , n382923 , n19644 );
or ( n382925 , n382921 , n382924 );
nand ( n382926 , n380636 , n19643 );
or ( n382927 , n382926 , n380575 );
nand ( n382928 , n382925 , n382927 );
not ( n382929 , n382923 );
and ( n382930 , n382921 , n382929 , n381522 );
or ( n382931 , n382928 , n382930 );
and ( n382932 , n380736 , n380741 );
nand ( n382933 , n382932 , n380737 );
not ( n382934 , n382933 );
and ( n382935 , n382931 , n382934 );
not ( n382936 , n382898 );
not ( n382937 , n380750 );
and ( n382938 , n382933 , n382936 , n382937 );
nor ( n382939 , n382938 , n19630 );
not ( n382940 , n380218 );
buf ( n382941 , n380759 );
nor ( n382942 , n382940 , n382941 );
or ( n382943 , n382939 , n382942 );
nand ( n382944 , n382943 , n19595 );
nand ( n382945 , n380763 , RI15b58650_881);
not ( n382946 , n381493 );
or ( n382947 , n382945 , n382946 );
nand ( n382948 , n382944 , n382947 );
and ( n382949 , n382948 , n380775 );
not ( n382950 , RI15b59820_919);
or ( n382951 , n382949 , n382950 );
buf ( n382952 , n380291 );
buf ( n382953 , n382952 );
buf ( n382954 , n382953 );
not ( n382955 , n382954 );
buf ( n382956 , n382955 );
buf ( n382957 , n382956 );
buf ( n382958 , n382957 );
not ( n382959 , n382958 );
not ( n382960 , n382942 );
not ( n382961 , n382947 );
not ( n382962 , n382961 );
and ( n382963 , n382960 , n382962 );
nor ( n382964 , n382963 , n382939 );
not ( n382965 , n382964 );
or ( n382966 , n382959 , n382965 );
or ( n382967 , n19547 , n380788 );
or ( n382968 , n382947 , n382967 );
nand ( n382969 , n382951 , n382966 , n382968 );
nor ( n382970 , n382935 , n382969 );
nand ( n382971 , n382914 , n382970 );
buf ( n382972 , n382971 );
buf ( n382973 , n379403 );
not ( n382974 , n380734 );
nand ( n382975 , n382974 , n381493 );
not ( n382976 , n382975 );
not ( n382977 , n382976 );
not ( n382978 , n381589 );
or ( n382979 , n382977 , n382978 );
not ( n382980 , n380736 );
and ( n382981 , n382980 , n380742 );
nand ( n382982 , n382981 , n380757 );
not ( n382983 , n382982 );
and ( n382984 , n381596 , n382983 );
not ( n382985 , n380750 );
and ( n382986 , n382982 , n382975 , n382985 );
nor ( n382987 , n382986 , n19630 );
buf ( n382988 , n380224 );
nor ( n382989 , n382988 , n380728 );
or ( n382990 , n382987 , n382989 );
nand ( n382991 , n382990 , n19595 );
or ( n382992 , n381538 , RI15b58650_881);
or ( n382993 , n382992 , n381540 );
nand ( n382994 , n382991 , n382993 );
and ( n382995 , n382994 , n380775 );
or ( n382996 , n382995 , n18701 );
buf ( n382997 , n381614 );
not ( n382998 , n382997 );
not ( n382999 , n382993 );
nor ( n383000 , n382989 , n382999 );
or ( n383001 , n382987 , n383000 );
or ( n383002 , n382998 , n383001 );
or ( n383003 , n382993 , n381621 );
nand ( n383004 , n382996 , n383002 , n383003 );
nor ( n383005 , n382984 , n383004 );
nand ( n383006 , n382979 , n383005 );
buf ( n383007 , n383006 );
not ( n383008 , n381453 );
not ( n383009 , RI15b54ca8_758);
not ( n383010 , RI15b54d98_760);
and ( n383011 , n383008 , n383009 , n382643 , n383010 );
not ( n383012 , RI15b54e88_762);
not ( n383013 , RI15b54f00_763);
and ( n383014 , n383011 , n382646 , n383012 , n383013 );
not ( n383015 , RI15b54f78_764);
not ( n383016 , RI15b55068_766);
and ( n383017 , n383014 , n383015 , n382651 , n383016 );
not ( n383018 , RI15b55158_768);
nand ( n383019 , n383017 , n382654 , n383018 , n382657 );
not ( n383020 , n383019 );
not ( n383021 , RI15b55248_770);
not ( n383022 , RI15b552c0_771);
nand ( n383023 , n383020 , n382662 , n383021 , n383022 );
not ( n383024 , n383023 );
not ( n383025 , RI15b553b0_773);
nand ( n383026 , n383024 , n383025 , n382666 );
nor ( n383027 , n383026 , RI15b554a0_775);
not ( n383028 , n383027 );
nand ( n383029 , n383026 , RI15b554a0_775);
nand ( n383030 , n383028 , n383029 );
nand ( n383031 , n383023 , RI15b55770_781);
not ( n383032 , n383031 );
not ( n383033 , RI15b553b0_773);
and ( n383034 , n383032 , n383033 );
and ( n383035 , n383031 , RI15b553b0_773);
nor ( n383036 , n383034 , n383035 );
buf ( n383037 , n383017 );
not ( n383038 , n383037 );
nand ( n383039 , RI15b550e0_767 , RI15b55158_768 , RI15b55248_770 , RI15b55338_772);
nor ( n383040 , n383039 , n383022 , n382657 );
nand ( n383041 , n383038 , n383040 );
not ( n383042 , n383041 );
not ( n383043 , n383023 );
or ( n383044 , n383042 , n383043 );
buf ( n383045 , n383014 );
nand ( n383046 , n383045 , n383015 , n382651 );
nand ( n383047 , n383046 , RI15b55770_781);
not ( n383048 , n383047 );
not ( n383049 , RI15b55068_766);
and ( n383050 , n383048 , n383049 );
and ( n383051 , n383047 , RI15b55068_766);
nor ( n383052 , n383050 , n383051 );
nand ( n383053 , n383044 , n383052 );
not ( n383054 , n383053 );
nand ( n383055 , n383036 , n383054 );
buf ( n383056 , n383055 );
and ( n383057 , n383030 , n383056 );
not ( n383058 , n383030 );
not ( n383059 , n383055 );
and ( n383060 , n383058 , n383059 );
nor ( n383061 , n383057 , n383060 );
not ( n383062 , n383061 );
not ( n383063 , n383056 );
not ( n383064 , n383063 );
not ( n383065 , n383064 );
and ( n383066 , n383062 , n383065 );
not ( n383067 , n383063 );
and ( n383068 , n383061 , n383067 );
nor ( n383069 , n383066 , n383068 );
and ( n383070 , RI15b55770_781 , n383069 );
not ( n383071 , RI15b55770_781);
and ( n383072 , n383071 , n382665 );
nor ( n383073 , n383070 , n383072 );
buf ( n383074 , n383073 );
not ( n383075 , n383074 );
buf ( n383076 , n383026 );
buf ( n383077 , n383076 );
not ( n383078 , RI15b55428_774);
not ( n383079 , n383023 );
nand ( n383080 , n383079 , n383025 );
not ( n383081 , n383080 );
or ( n383082 , n383078 , n383081 );
nand ( n383083 , n383082 , RI15b55770_781);
not ( n383084 , n383083 );
and ( n383085 , n383077 , n383084 );
nor ( n383086 , n382666 , RI15b55770_781);
nor ( n383087 , n383085 , n383086 );
not ( n383088 , n383038 );
nand ( n383089 , n383088 , n382654 , n383018 );
nand ( n383090 , n383089 , RI15b55770_781);
not ( n383091 , n383090 );
not ( n383092 , RI15b551d0_769);
and ( n383093 , n383091 , n383092 );
and ( n383094 , n383090 , RI15b551d0_769);
nor ( n383095 , n383093 , n383094 );
not ( n383096 , RI15b55158_768);
nand ( n383097 , n383037 , n382654 );
nand ( n383098 , n383097 , RI15b55770_781);
not ( n383099 , n383098 );
or ( n383100 , n383096 , n383099 );
or ( n383101 , n383098 , RI15b55158_768);
nand ( n383102 , n383100 , n383101 );
not ( n383103 , n383037 );
nand ( n383104 , n383103 , RI15b55770_781);
not ( n383105 , n383104 );
not ( n383106 , RI15b550e0_767);
and ( n383107 , n383105 , n383106 );
and ( n383108 , n383104 , RI15b550e0_767);
nor ( n383109 , n383107 , n383108 );
nand ( n383110 , n383109 , n383052 );
nor ( n383111 , n383102 , n383110 );
and ( n383112 , n383095 , n383111 );
buf ( n383113 , n383020 );
not ( n383114 , n383113 );
nand ( n383115 , n383114 , RI15b55770_781);
not ( n383116 , n383115 );
not ( n383117 , RI15b55248_770);
and ( n383118 , n383116 , n383117 );
and ( n383119 , n383115 , RI15b55248_770);
nor ( n383120 , n383118 , n383119 );
nand ( n383121 , n383112 , n383120 );
not ( n383122 , RI15b552c0_771);
nand ( n383123 , n383113 , n383021 );
nand ( n383124 , n383123 , RI15b55770_781);
not ( n383125 , n383124 );
or ( n383126 , n383122 , n383125 );
or ( n383127 , n383124 , RI15b552c0_771);
nand ( n383128 , n383126 , n383127 );
nor ( n383129 , n383121 , n383128 );
not ( n383130 , n383123 );
nand ( n383131 , n383130 , n383022 );
nand ( n383132 , n383131 , RI15b55770_781);
not ( n383133 , n383132 );
not ( n383134 , RI15b55338_772);
and ( n383135 , n383133 , n383134 );
and ( n383136 , n383132 , RI15b55338_772);
nor ( n383137 , n383135 , n383136 );
nand ( n383138 , n383129 , n383137 );
not ( n383139 , n383036 );
nor ( n383140 , n383138 , n383139 );
nand ( n383141 , n383087 , n383140 );
not ( n383142 , n383141 );
and ( n383143 , n381461 , n18096 );
not ( n383144 , n383143 );
nor ( n383145 , n383142 , n383144 );
and ( n383146 , n383075 , n383145 );
not ( n383147 , n18167 );
and ( n383148 , n383147 , RI15b52908_682);
nor ( n383149 , n383146 , n383148 );
not ( n383150 , n383075 );
not ( n383151 , n381421 );
or ( n383152 , n383151 , n382546 );
not ( n383153 , n383152 );
not ( n383154 , n383153 );
not ( n383155 , n383142 );
or ( n383156 , n383154 , n383155 );
or ( n383157 , n381450 , n382546 );
nand ( n383158 , n383156 , n383157 );
nand ( n383159 , n383150 , n383158 );
nand ( n383160 , n381474 , n381479 );
not ( n383161 , n382547 );
and ( n383162 , n383161 , n18077 );
nor ( n383163 , n18173 , n18170 );
nand ( n383164 , n21786 , n383163 );
and ( n383165 , n18164 , n21750 );
nand ( n383166 , n383165 , n18165 );
nor ( n383167 , n383162 , n383164 , n383166 );
nand ( n383168 , n383167 , n379993 );
nor ( n383169 , n383160 , n383168 );
not ( n383170 , n383169 );
nand ( n383171 , n383170 , RI15b53f10_729);
nand ( n383172 , n383149 , n383159 , n383171 );
buf ( n383173 , n383172 );
buf ( n383174 , RI15b3ea48_2);
buf ( n383175 , n383174 );
buf ( n383176 , n17499 );
buf ( n383177 , n22406 );
buf ( n383178 , n22404 );
not ( n383179 , n380647 );
nand ( n383180 , n383179 , n19644 );
or ( n383181 , n383180 , n382975 );
not ( n383182 , n382995 );
and ( n383183 , n383182 , RI15b5ad38_964);
nand ( n383184 , n382918 , n19642 );
or ( n383185 , n383184 , n382982 );
buf ( n383186 , n380315 );
not ( n383187 , n383186 );
buf ( n383188 , n383187 );
not ( n383189 , n383188 );
or ( n383190 , n383189 , n383001 );
buf ( n383191 , n18972 );
or ( n383192 , n383191 , n380788 );
or ( n383193 , n382993 , n383192 );
nand ( n383194 , n383185 , n383190 , n383193 );
nor ( n383195 , n383183 , n383194 );
nand ( n383196 , n383181 , n383195 );
buf ( n383197 , n383196 );
not ( n383198 , RI15b556f8_780);
not ( n383199 , n382683 );
not ( n383200 , n383076 );
nor ( n383201 , RI15b554a0_775 , RI15b55518_776);
nand ( n383202 , n383200 , n383201 );
not ( n383203 , RI15b55590_777);
nand ( n383204 , n383203 , n382686 );
nor ( n383205 , n383202 , n383204 );
buf ( n383206 , n383205 );
not ( n383207 , n383206 );
or ( n383208 , n383199 , n383207 );
nand ( n383209 , n383208 , RI15b55770_781);
not ( n383210 , n383209 );
or ( n383211 , n383198 , n383210 );
or ( n383212 , n383209 , RI15b556f8_780);
nand ( n383213 , n383211 , n383212 );
not ( n383214 , n383213 );
not ( n383215 , n383153 );
not ( n383216 , RI15b55770_781);
and ( n383217 , n383216 , n382686 );
not ( n383218 , n383216 );
nand ( n383219 , n383061 , n383063 );
not ( n383220 , n383219 );
not ( n383221 , n382669 );
nand ( n383222 , n383036 , n383054 );
buf ( n383223 , n383029 );
nor ( n383224 , n383222 , n383223 );
not ( n383225 , n383224 );
or ( n383226 , n383221 , n383225 );
not ( n383227 , n382665 );
not ( n383228 , n383222 );
not ( n383229 , n383228 );
or ( n383230 , n383227 , n383229 );
not ( n383231 , n383076 );
nand ( n383232 , n383231 , RI15b554a0_775);
nand ( n383233 , n383230 , n383232 );
and ( n383234 , n383222 , n383076 );
or ( n383235 , n383233 , n383234 );
nand ( n383236 , n383235 , RI15b55518_776);
nand ( n383237 , n383226 , n383236 );
not ( n383238 , n383237 );
nand ( n383239 , n383220 , n383238 );
not ( n383240 , n383239 );
not ( n383241 , RI15b55590_777);
not ( n383242 , n382665 );
not ( n383243 , RI15b55518_776);
and ( n383244 , n383242 , n383243 );
not ( n383245 , n383076 );
and ( n383246 , n383245 , RI15b55518_776);
nor ( n383247 , n383244 , n383246 );
not ( n383248 , n383222 );
nand ( n383249 , n383076 , n382665 );
nand ( n383250 , n383247 , n383248 , n383249 );
not ( n383251 , n383250 );
nand ( n383252 , n383251 , n383202 );
not ( n383253 , n383252 );
or ( n383254 , n383241 , n383253 );
not ( n383255 , n383223 );
not ( n383256 , n383056 );
nand ( n383257 , n383255 , n383256 );
not ( n383258 , n383257 );
nand ( n383259 , n383203 , RI15b55518_776);
not ( n383260 , n383259 );
and ( n383261 , n383258 , n383260 );
not ( n383262 , n383059 );
not ( n383263 , n383262 );
nand ( n383264 , n383263 , n383247 , n383249 );
not ( n383265 , n383202 );
and ( n383266 , n383264 , n383265 );
nor ( n383267 , n383261 , n383266 );
nand ( n383268 , n383254 , n383267 );
not ( n383269 , n383268 );
nand ( n383270 , n383240 , n383269 );
not ( n383271 , n383270 );
not ( n383272 , RI15b55590_777);
not ( n383273 , n383252 );
not ( n383274 , n383273 );
or ( n383275 , n383272 , n383274 );
nand ( n383276 , n383275 , RI15b55608_778);
not ( n383277 , n383257 );
nand ( n383278 , n382686 , RI15b55590_777 , RI15b55518_776);
not ( n383279 , n383278 );
and ( n383280 , n383277 , n383279 );
buf ( n383281 , n383264 );
and ( n383282 , n383281 , n383205 );
nor ( n383283 , n383280 , n383282 );
nand ( n383284 , n383276 , n383283 );
not ( n383285 , n383284 );
not ( n383286 , n383285 );
and ( n383287 , n383271 , n383286 );
not ( n383288 , n383268 );
nand ( n383289 , n383240 , n383288 );
not ( n383290 , n383284 );
and ( n383291 , n383289 , n383290 );
nor ( n383292 , n383287 , n383291 );
and ( n383293 , n383218 , n383292 );
nor ( n383294 , n383217 , n383293 );
not ( n383295 , RI15b55770_781);
and ( n383296 , n383295 , RI15b55590_777);
not ( n383297 , n383295 );
not ( n383298 , n383268 );
not ( n383299 , n383298 );
nand ( n383300 , n383220 , n383238 );
not ( n383301 , n383300 );
or ( n383302 , n383299 , n383301 );
or ( n383303 , n383300 , n383288 );
nand ( n383304 , n383302 , n383303 );
and ( n383305 , n383297 , n383304 );
nor ( n383306 , n383296 , n383305 );
not ( n383307 , n383237 );
not ( n383308 , n383219 );
not ( n383309 , n383308 );
or ( n383310 , n383307 , n383309 );
not ( n383311 , n383219 );
or ( n383312 , n383311 , n383237 );
nand ( n383313 , n383310 , n383312 );
and ( n383314 , n383313 , RI15b55770_781);
nor ( n383315 , n382669 , RI15b55770_781);
nor ( n383316 , n383314 , n383315 );
nor ( n383317 , n383073 , n383141 );
and ( n383318 , n383316 , n383317 );
nand ( n383319 , n383306 , n383318 );
nor ( n383320 , n383294 , n383319 );
not ( n383321 , n383206 );
nand ( n383322 , n383321 , RI15b55770_781);
and ( n383323 , n383322 , RI15b55680_779);
not ( n383324 , n383322 );
and ( n383325 , n383324 , n382683 );
nor ( n383326 , n383323 , n383325 );
and ( n383327 , n383320 , n383326 );
not ( n383328 , n383327 );
or ( n383329 , n383215 , n383328 );
nand ( n383330 , n383329 , n383157 );
not ( n383331 , n383330 );
or ( n383332 , n383214 , n383331 );
nor ( n383333 , n383213 , n383144 );
not ( n383334 , n383333 );
not ( n383335 , n383327 );
not ( n383336 , n383335 );
or ( n383337 , n383334 , n383336 );
and ( n383338 , n383170 , RI15b54168_734);
and ( n383339 , n383147 , RI15b52b60_687);
nor ( n383340 , n383338 , n383339 );
nand ( n383341 , n383337 , n383340 );
not ( n383342 , n383341 );
nand ( n383343 , n383332 , n383342 );
buf ( n383344 , n383343 );
buf ( n383345 , RI15b3e9d0_1);
buf ( n383346 , n383345 );
buf ( n383347 , n22005 );
buf ( n383348 , n381872 );
or ( n383349 , n19919 , n19731 );
nand ( n383350 , n383349 , n19938 );
nand ( n383351 , n383350 , n19740 );
not ( n383352 , n19740 );
buf ( n383353 , n20524 );
nand ( n383354 , n383352 , n383353 , n19731 );
not ( n383355 , n20534 );
and ( n383356 , n20565 , n383355 );
nor ( n383357 , n383356 , n22372 );
not ( n383358 , RI15b4b360_431);
or ( n383359 , n383357 , n383358 );
not ( n383360 , n19958 );
not ( n383361 , n383360 );
not ( n383362 , n22376 );
or ( n383363 , n383361 , n383362 );
not ( n383364 , n22383 );
nand ( n383365 , n383363 , n383364 );
and ( n383366 , n383365 , RI15b49560_367);
or ( n383367 , n20564 , n383355 , RI15b4b360_431);
not ( n383368 , n379830 );
buf ( n383369 , n20610 );
not ( n383370 , n383369 );
not ( n383371 , n383370 );
buf ( n383372 , n20003 );
not ( n383373 , n383372 );
buf ( n383374 , n20067 );
nor ( n383375 , n383373 , n383374 );
buf ( n383376 , n383375 );
buf ( n383377 , n383376 );
buf ( n383378 , n383377 );
buf ( n383379 , n383378 );
buf ( n383380 , n383379 );
not ( n383381 , n383380 );
buf ( n383382 , n383381 );
buf ( n383383 , n383382 );
not ( n383384 , n383383 );
and ( n383385 , n383384 , n20008 );
and ( n383386 , n383383 , RI15b44bc8_210);
nor ( n383387 , n383385 , n383386 );
or ( n383388 , n383368 , n383371 , n383387 );
nand ( n383389 , n383367 , n383388 );
nor ( n383390 , n22359 , n383360 , RI15b49560_367);
nor ( n383391 , n383366 , n383389 , n383390 );
nand ( n383392 , n383359 , n383391 );
nand ( n383393 , n383392 , n20501 );
and ( n383394 , n22388 , RI15b4b360_431);
and ( n383395 , n22391 , RI15b4a460_399);
not ( n383396 , n22397 );
nor ( n383397 , n383394 , n383395 , n383396 );
nand ( n383398 , n383351 , n383354 , n383393 , n383397 );
buf ( n383399 , n383398 );
buf ( n383400 , n380865 );
buf ( n383401 , n21800 );
buf ( n383402 , n22458 );
nor ( n383403 , RI15b61c50_1201 , RI15b61cc8_1202);
buf ( n383404 , n383403 );
and ( n383405 , n383402 , n383404 );
not ( n383406 , RI15b62ad8_1232);
nand ( n383407 , n22457 , n383406 );
and ( n383408 , n383407 , n22466 );
not ( n383409 , n383408 );
nor ( n383410 , n383405 , n383409 );
not ( n383411 , RI15b61d40_1203);
or ( n383412 , n383410 , n383411 );
not ( n383413 , n22422 );
and ( n383414 , n383413 , RI15b63b40_1267);
or ( n383415 , n379787 , RI15b63b40_1267);
or ( n383416 , n379498 , RI15b63ac8_1266);
nand ( n383417 , n383415 , n383416 );
and ( n383418 , n22450 , n383417 );
nand ( n383419 , RI15b63528_1254 , RI15b635a0_1255);
not ( n383420 , RI15b63618_1256);
nor ( n383421 , n383419 , n383420 );
nand ( n383422 , n383421 , RI15b63690_1257);
not ( n383423 , RI15b63708_1258);
nor ( n383424 , n383422 , n383423 );
nand ( n383425 , n383424 , RI15b63780_1259);
not ( n383426 , RI15b637f8_1260);
nor ( n383427 , n383425 , n383426 );
nand ( n383428 , n383427 , RI15b63870_1261);
not ( n383429 , RI15b638e8_1262);
or ( n383430 , n383428 , n383429 );
not ( n383431 , RI15b63960_1263);
or ( n383432 , n383430 , n383431 );
not ( n383433 , n383432 );
nand ( n383434 , RI15b63168_1246 , RI15b631e0_1247);
not ( n383435 , n383434 );
and ( n383436 , n383435 , RI15b63258_1248);
and ( n383437 , n383436 , RI15b632d0_1249);
nand ( n383438 , n383437 , RI15b63348_1250);
not ( n383439 , RI15b633c0_1251);
or ( n383440 , n383438 , n383439 );
not ( n383441 , RI15b63438_1252);
or ( n383442 , n383440 , n383441 );
not ( n383443 , n383442 );
and ( n383444 , n380845 , RI15b62f88_1242);
nand ( n383445 , n383444 , RI15b63000_1243);
not ( n383446 , RI15b63078_1244);
nor ( n383447 , n383445 , n383446 );
and ( n383448 , n383447 , RI15b62bc8_1234);
nand ( n383449 , n383448 , RI15b630f0_1245);
buf ( n383450 , n383449 );
buf ( n383451 , n383450 );
not ( n383452 , n383451 );
nand ( n383453 , n383443 , n383452 );
not ( n383454 , RI15b634b0_1253);
nor ( n383455 , n383453 , n383454 );
buf ( n383456 , n383455 );
nand ( n383457 , n383433 , n383456 );
not ( n383458 , n383457 );
not ( n383459 , RI15b639d8_1264);
and ( n383460 , n383458 , n383459 );
and ( n383461 , n383457 , RI15b639d8_1264);
nor ( n383462 , n383460 , n383461 );
not ( n383463 , n383462 );
nand ( n383464 , n383463 , n19628 );
not ( n383465 , n383464 );
nand ( n383466 , RI15b62bc8_1234 , RI15b62c40_1235);
not ( n383467 , RI15b62b50_1233);
or ( n383468 , n383466 , n383467 );
or ( n383469 , RI15b62bc8_1234 , RI15b62c40_1235);
nand ( n383470 , n383468 , n383469 );
and ( n383471 , n383465 , n383470 );
nor ( n383472 , n383414 , n383418 , n383471 );
nand ( n383473 , n383462 , n19628 );
buf ( n383474 , n383473 );
not ( n383475 , n383474 );
not ( n383476 , RI15b62c40_1235);
or ( n383477 , n383476 , RI15b62bc8_1234);
nor ( n383478 , n19620 , RI15b62c40_1235);
not ( n383479 , n383478 );
nand ( n383480 , n383477 , n383479 );
and ( n383481 , n383475 , n383480 );
or ( n383482 , n22456 , n383406 );
nor ( n383483 , n383482 , n383404 , RI15b61d40_1203);
not ( n383484 , n18386 );
buf ( n383485 , n383484 );
not ( n383486 , n383485 );
not ( n383487 , n22471 );
or ( n383488 , n383486 , n383487 );
and ( n383489 , n22423 , RI15b63b40_1267);
nor ( n383490 , n22473 , RI15b62b50_1233);
and ( n383491 , n383490 , n383478 );
and ( n383492 , n19599 , RI15b62c40_1235);
nor ( n383493 , n383489 , n383491 , n383492 );
nand ( n383494 , n383488 , n383493 );
nor ( n383495 , n383481 , n383483 , n383494 );
nand ( n383496 , n383412 , n383472 , n383495 );
buf ( n383497 , n383496 );
buf ( n383498 , RI15b3ea48_2);
buf ( n383499 , n383498 );
nand ( n383500 , n22463 , n22444 );
not ( n383501 , n19539 );
nand ( n383502 , n383501 , n22462 , n22444 );
nand ( n383503 , n383500 , n383502 );
buf ( n383504 , n383503 );
buf ( n383505 , n383504 );
nor ( n383506 , RI15b60d50_1169 , RI15b60fa8_1174);
not ( n383507 , RI15b61020_1175);
nand ( n383508 , n383506 , n383507 );
nor ( n383509 , RI15b60dc8_1170 , RI15b60e40_1171);
nor ( n383510 , RI15b60eb8_1172 , RI15b60f30_1173);
nand ( n383511 , n383509 , n383510 );
nor ( n383512 , n383508 , n383511 );
buf ( n383513 , n383512 );
and ( n383514 , n383513 , RI15b61bd8_1200);
buf ( n383515 , n383506 );
nand ( n383516 , n383515 , RI15b61bd8_1200);
nor ( n383517 , n383516 , n383511 );
not ( n383518 , RI15b61020_1175);
nor ( n383519 , n383517 , n383518 );
nor ( n383520 , n383514 , n383519 );
not ( n383521 , n383517 );
nor ( n383522 , n383520 , n383521 );
not ( n383523 , RI15b61bd8_1200);
nor ( n383524 , n383512 , n383523 );
not ( n383525 , RI15b61098_1176);
and ( n383526 , n383524 , n383525 );
not ( n383527 , n383524 );
and ( n383528 , n383527 , RI15b61098_1176);
nor ( n383529 , n383526 , n383528 );
and ( n383530 , n383522 , n383529 );
and ( n383531 , n383512 , n383525 );
buf ( n383532 , n383531 );
nor ( n383533 , n383532 , n383523 );
not ( n383534 , RI15b61110_1177);
and ( n383535 , n383533 , n383534 );
not ( n383536 , n383533 );
and ( n383537 , n383536 , RI15b61110_1177);
nor ( n383538 , n383535 , n383537 );
and ( n383539 , n383530 , n383538 );
nand ( n383540 , n383531 , n383534 );
nand ( n383541 , n383540 , RI15b61bd8_1200);
not ( n383542 , n383541 );
not ( n383543 , RI15b61188_1178);
and ( n383544 , n383542 , n383543 );
and ( n383545 , n383541 , RI15b61188_1178);
nor ( n383546 , n383544 , n383545 );
nand ( n383547 , n383539 , n383546 );
not ( n383548 , RI15b61200_1179);
nor ( n383549 , n383540 , RI15b61188_1178);
not ( n383550 , n383549 );
nand ( n383551 , n383550 , RI15b61bd8_1200);
not ( n383552 , n383551 );
or ( n383553 , n383548 , n383552 );
or ( n383554 , n383551 , RI15b61200_1179);
nand ( n383555 , n383553 , n383554 );
nor ( n383556 , n383547 , n383555 );
not ( n383557 , RI15b61200_1179);
nand ( n383558 , n383549 , n383557 );
buf ( n383559 , n383558 );
nand ( n383560 , n383559 , RI15b61bd8_1200);
and ( n383561 , n383560 , RI15b61278_1180);
not ( n383562 , n383560 );
not ( n383563 , RI15b61278_1180);
and ( n383564 , n383562 , n383563 );
nor ( n383565 , n383561 , n383564 );
nand ( n383566 , n383556 , n383565 );
nor ( n383567 , n383558 , RI15b61278_1180);
not ( n383568 , n383567 );
nand ( n383569 , n383568 , RI15b61bd8_1200);
not ( n383570 , RI15b612f0_1181);
and ( n383571 , n383569 , n383570 );
not ( n383572 , n383569 );
and ( n383573 , n383572 , RI15b612f0_1181);
nor ( n383574 , n383571 , n383573 );
nor ( n383575 , n383566 , n383574 );
and ( n383576 , n383505 , n383575 );
and ( n383577 , n383504 , n383523 );
nor ( n383578 , n383576 , n383577 );
and ( n383579 , n383567 , n383570 );
not ( n383580 , n383579 );
nand ( n383581 , n383580 , RI15b61bd8_1200);
and ( n383582 , n383581 , RI15b61368_1182);
not ( n383583 , n383581 );
not ( n383584 , RI15b61368_1182);
and ( n383585 , n383583 , n383584 );
nor ( n383586 , n383582 , n383585 );
or ( n383587 , n383578 , n383586 );
buf ( n383588 , n19552 );
not ( n383589 , n22444 );
nor ( n383590 , n383588 , n383589 );
not ( n383591 , n383590 );
not ( n383592 , n22420 );
or ( n383593 , n383591 , n383592 );
nand ( n383594 , n383593 , n19201 );
nand ( n383595 , n380773 , n19577 );
not ( n383596 , n19600 );
not ( n383597 , n19629 );
nand ( n383598 , n383597 , n380748 );
nor ( n383599 , n383595 , n383596 , n383598 );
and ( n383600 , n383594 , n383599 );
not ( n383601 , n383600 );
and ( n383602 , n383601 , RI15b5fdd8_1136);
and ( n383603 , n383503 , RI15b61bd8_1200);
not ( n383604 , n383586 );
nor ( n383605 , n383604 , n383575 );
and ( n383606 , n383603 , n383605 );
not ( n383607 , n19579 );
and ( n383608 , n383607 , RI15b5f658_1120);
nor ( n383609 , n383602 , n383606 , n383608 );
nand ( n383610 , n383587 , n383609 );
buf ( n383611 , n383610 );
buf ( n383612 , n22005 );
buf ( n383613 , RI15b3e9d0_1);
buf ( n383614 , n383613 );
not ( n383615 , n381121 );
not ( n383616 , n380407 );
and ( n383617 , n383615 , n383616 );
and ( n383618 , n381114 , RI15b65fd0_1345);
nor ( n383619 , n383617 , n383618 );
nand ( n383620 , n381196 , n383619 , n381185 );
nor ( n383621 , n383620 , n381217 );
nand ( n383622 , n381116 , n381190 );
nor ( n383623 , n381226 , n383622 );
nor ( n383624 , n381133 , n381201 );
and ( n383625 , n381179 , n383621 , n383623 , n383624 );
not ( n383626 , n381114 );
not ( n383627 , n380420 );
and ( n383628 , n383626 , n383627 );
buf ( n383629 , n381110 );
and ( n383630 , n383629 , RI15b66048_1346);
nor ( n383631 , n383628 , n383630 );
nand ( n383632 , n383625 , n383631 );
nand ( n383633 , n381110 , RI15b66138_1348);
not ( n383634 , n383633 );
buf ( n383635 , n381110 );
nor ( n383636 , n383635 , n380433 );
nor ( n383637 , n383634 , n383636 );
not ( n383638 , n381110 );
nand ( n383639 , n383638 , RI15b651c0_1315);
nand ( n383640 , n381138 , RI15b660c0_1347);
and ( n383641 , n383639 , n383640 );
and ( n383642 , n381138 , RI15b661b0_1349);
not ( n383643 , n381138 );
and ( n383644 , n383643 , RI15b652b0_1317);
nor ( n383645 , n383642 , n383644 );
nand ( n383646 , n383637 , n383641 , n383645 );
nor ( n383647 , n383632 , n383646 );
not ( n383648 , n383629 );
and ( n383649 , n383648 , RI15b65328_1318);
and ( n383650 , n381138 , RI15b66228_1350);
nor ( n383651 , n383649 , n383650 );
not ( n383652 , n381114 );
not ( n383653 , n380472 );
and ( n383654 , n383652 , n383653 );
not ( n383655 , n383638 );
and ( n383656 , n383655 , RI15b662a0_1351);
nor ( n383657 , n383654 , n383656 );
and ( n383658 , n383647 , n383651 , n383657 );
not ( n383659 , n383658 );
not ( n383660 , n383659 );
and ( n383661 , n381138 , RI15b66318_1352);
not ( n383662 , n381138 );
and ( n383663 , n383662 , RI15b65418_1320);
nor ( n383664 , n383661 , n383663 );
not ( n383665 , n381114 );
not ( n383666 , n380583 );
and ( n383667 , n383665 , n383666 );
and ( n383668 , n383629 , RI15b66390_1353);
nor ( n383669 , n383667 , n383668 );
and ( n383670 , n383664 , n383669 );
not ( n383671 , n382693 );
not ( n383672 , n380463 );
and ( n383673 , n383671 , n383672 );
and ( n383674 , n382693 , RI15b66408_1354);
nor ( n383675 , n383673 , n383674 );
and ( n383676 , n383670 , n383675 );
not ( n383677 , n382693 );
and ( n383678 , n383677 , RI15b65580_1323);
and ( n383679 , n382693 , RI15b66480_1355);
nor ( n383680 , n383678 , n383679 );
and ( n383681 , n383676 , n383680 );
and ( n383682 , n383660 , n383681 );
not ( n383683 , n382694 );
and ( n383684 , n383683 , RI15b655f8_1324);
and ( n383685 , n382699 , RI15b664f8_1356);
nor ( n383686 , n383684 , n383685 );
nand ( n383687 , n383682 , n383686 );
not ( n383688 , n383664 );
not ( n383689 , n383688 );
not ( n383690 , n383660 );
or ( n383691 , n383689 , n383690 );
not ( n383692 , n383659 );
or ( n383693 , n383692 , n383688 );
nand ( n383694 , n383691 , n383693 );
not ( n383695 , n381133 );
nand ( n383696 , n383695 , n381117 );
nor ( n383697 , n381228 , n383696 );
not ( n383698 , n381142 );
nor ( n383699 , n383697 , n383698 );
buf ( n383700 , n383619 );
and ( n383701 , n383699 , n383700 );
not ( n383702 , n383699 );
not ( n383703 , n383700 );
and ( n383704 , n383702 , n383703 );
nor ( n383705 , n383701 , n383704 );
buf ( n383706 , n383632 );
and ( n383707 , n383706 , n383641 );
not ( n383708 , n383706 );
not ( n383709 , n383641 );
and ( n383710 , n383708 , n383709 );
nor ( n383711 , n383707 , n383710 );
and ( n383712 , n383705 , n383711 );
not ( n383713 , n383645 );
not ( n383714 , n383713 );
not ( n383715 , n383625 );
nor ( n383716 , n383715 , n383709 );
not ( n383717 , n383716 );
or ( n383718 , n383714 , n383717 );
not ( n383719 , n383637 );
or ( n383720 , n383716 , n383719 );
nand ( n383721 , n383718 , n383720 );
or ( n383722 , n383715 , n383631 );
nand ( n383723 , n383715 , n383631 );
and ( n383724 , n383719 , n383645 );
not ( n383725 , n383657 );
and ( n383726 , n383725 , n383651 );
and ( n383727 , n383629 , RI15b66660_1359);
not ( n383728 , n383629 );
and ( n383729 , n383728 , RI15b65760_1327);
nor ( n383730 , n383727 , n383729 );
nor ( n383731 , n383724 , n383726 , n383730 );
nand ( n383732 , n383722 , n383723 , n383731 );
nor ( n383733 , n383721 , n383732 );
buf ( n383734 , n383647 );
not ( n383735 , n383651 );
and ( n383736 , n383734 , n383735 );
not ( n383737 , n383734 );
and ( n383738 , n383737 , n383657 );
nor ( n383739 , n383736 , n383738 );
not ( n383740 , n382695 );
and ( n383741 , n383740 , RI15b66570_1357);
not ( n383742 , n383740 );
and ( n383743 , n383742 , RI15b65670_1325);
nor ( n383744 , n383741 , n383743 );
nor ( n383745 , n382702 , n383744 );
nand ( n383746 , n383712 , n383733 , n383739 , n383745 );
nor ( n383747 , n383694 , n383746 );
nand ( n383748 , n383687 , n383747 );
not ( n383749 , n383686 );
not ( n383750 , n383749 );
not ( n383751 , n383682 );
or ( n383752 , n383750 , n383751 );
or ( n383753 , n383682 , n383749 );
nand ( n383754 , n383752 , n383753 );
nor ( n383755 , n383748 , n383754 );
not ( n383756 , n383755 );
not ( n383757 , n381145 );
not ( n383758 , n383757 );
not ( n383759 , n383659 );
or ( n383760 , n383758 , n383759 );
nand ( n383761 , n383760 , n383670 );
and ( n383762 , n383761 , n383675 );
not ( n383763 , n383659 );
not ( n383764 , n383670 );
nor ( n383765 , n383764 , n383675 );
and ( n383766 , n383763 , n383765 );
nor ( n383767 , n383762 , n383766 );
not ( n383768 , n383664 );
not ( n383769 , n383658 );
or ( n383770 , n383768 , n383769 );
nand ( n383771 , n383770 , n383757 );
not ( n383772 , n383771 );
not ( n383773 , n383669 );
not ( n383774 , n383773 );
and ( n383775 , n383772 , n383774 );
and ( n383776 , n383771 , n383773 );
nor ( n383777 , n383775 , n383776 );
nand ( n383778 , n383767 , n383777 );
not ( n383779 , n383676 );
nand ( n383780 , n383659 , n381146 );
not ( n383781 , n383780 );
or ( n383782 , n383779 , n383781 );
nand ( n383783 , n383782 , n383680 );
not ( n383784 , n383680 );
and ( n383785 , n383676 , n383784 );
nand ( n383786 , n383763 , n383785 );
nand ( n383787 , n383783 , n383786 );
nor ( n383788 , n383778 , n383787 );
not ( n383789 , n383788 );
or ( n383790 , n383756 , n383789 );
nand ( n383791 , n383790 , n381395 );
not ( n383792 , n383791 );
not ( n383793 , n383723 );
and ( n383794 , n383792 , n383793 );
nand ( n383795 , n383715 , n381395 );
not ( n383796 , n383631 );
and ( n383797 , n383795 , n383796 );
nor ( n383798 , n383794 , n383797 );
not ( n383799 , n383798 );
not ( n383800 , n383791 );
not ( n383801 , n21775 );
or ( n383802 , n383705 , n383801 );
not ( n383803 , n383802 );
nand ( n383804 , n383800 , n383803 );
nor ( n383805 , n383799 , n383804 );
not ( n383806 , n383805 );
nand ( n383807 , n383705 , n21794 );
not ( n383808 , n383807 );
nand ( n383809 , n383791 , n22704 );
not ( n383810 , n383809 );
or ( n383811 , n383808 , n383810 );
nand ( n383812 , n383811 , n383799 );
nand ( n383813 , n383806 , n383812 );
not ( n383814 , n383813 );
not ( n383815 , RI15b4c260_463);
not ( n383816 , n383815 );
not ( n383817 , n18006 );
nand ( n383818 , n383817 , RI15b4c1e8_462);
not ( n383819 , n383818 );
not ( n383820 , n383819 );
or ( n383821 , n383816 , n383820 );
nand ( n383822 , n383818 , RI15b4c260_463);
nand ( n383823 , n383821 , n383822 );
not ( n383824 , n383823 );
and ( n383825 , n17998 , n18007 );
not ( n383826 , n17998 );
not ( n383827 , n18007 );
and ( n383828 , n383826 , n383827 );
or ( n383829 , n383825 , n383828 );
not ( n383830 , n383829 );
nand ( n383831 , n383824 , n383830 );
not ( n383832 , n21337 );
nor ( n383833 , n383831 , n383832 );
not ( n383834 , n383832 );
not ( n383835 , n383823 );
or ( n383836 , n383834 , n383835 );
nand ( n383837 , n383823 , n383829 );
nand ( n383838 , n383836 , n383837 );
nor ( n383839 , n383833 , n383838 );
buf ( n383840 , n383839 );
buf ( n383841 , n383840 );
nand ( n383842 , n383829 , n21337 );
not ( n383843 , n383842 );
not ( n383844 , n383843 );
or ( n383845 , n383841 , n383844 );
or ( n383846 , n383814 , n383845 );
not ( n383847 , n383767 );
and ( n383848 , n383777 , n383847 );
nor ( n383849 , n383777 , n383847 );
nor ( n383850 , n383848 , n383849 );
nand ( n383851 , n381394 , n21776 );
nor ( n383852 , n383850 , n383851 );
not ( n383853 , n381395 );
buf ( n383854 , n21776 );
nand ( n383855 , n383853 , n383854 );
nor ( n383856 , n383855 , n383675 );
or ( n383857 , n383852 , n383856 );
not ( n383858 , n383839 );
not ( n383859 , n383832 );
not ( n383860 , n383830 );
or ( n383861 , n383859 , n383860 );
nand ( n383862 , n383861 , n383842 );
not ( n383863 , n383862 );
nor ( n383864 , n383858 , n383863 );
or ( n383865 , n18057 , RI15b4c170_461);
not ( n383866 , n383865 );
nand ( n383867 , n383864 , n383866 );
nor ( n383868 , n383839 , n383862 );
nor ( n383869 , n383839 , n383866 );
nor ( n383870 , n383868 , n383869 );
nand ( n383871 , n383867 , n383870 );
and ( n383872 , n383862 , n383866 );
not ( n383873 , n383862 );
and ( n383874 , n383873 , n383865 );
nor ( n383875 , n383872 , n383874 );
and ( n383876 , n383871 , n383875 );
nand ( n383877 , n383876 , n383866 );
not ( n383878 , n383877 );
and ( n383879 , n383857 , n383878 );
buf ( n383880 , n18174 );
not ( n383881 , n383880 );
not ( n383882 , n383881 );
and ( n383883 , n383877 , n383845 , n383882 );
nor ( n383884 , n383883 , n21764 );
nand ( n383885 , n383823 , n383830 );
buf ( n383886 , n18007 );
not ( n383887 , n383886 );
not ( n383888 , n383887 );
nor ( n383889 , n383885 , n383888 );
or ( n383890 , n383884 , n383889 );
nand ( n383891 , n383890 , n18154 );
nor ( n383892 , n383815 , RI15b4c2d8_464);
nand ( n383893 , n383892 , RI15b4c1e8_462);
nand ( n383894 , n18057 , n18062 );
or ( n383895 , n383893 , n383894 );
and ( n383896 , n383891 , n383895 );
or ( n383897 , n18154 , n17587 );
nand ( n383898 , n383897 , n18218 );
nor ( n383899 , n383898 , n18077 , n18168 );
nand ( n383900 , n383165 , n383899 );
nor ( n383901 , n383900 , n18156 );
not ( n383902 , n383901 );
nor ( n383903 , n383896 , n383902 );
or ( n383904 , n383903 , n21121 );
not ( n383905 , n381185 );
buf ( n383906 , n383905 );
buf ( n383907 , n383906 );
not ( n383908 , n383907 );
not ( n383909 , n383895 );
nor ( n383910 , n383889 , n383909 );
or ( n383911 , n383884 , n383910 );
or ( n383912 , n383908 , n383911 );
buf ( n383913 , n382690 );
not ( n383914 , n383913 );
and ( n383915 , n18155 , n17587 );
not ( n383916 , n383915 );
or ( n383917 , n383914 , n383916 );
or ( n383918 , n383895 , n383917 );
nand ( n383919 , n383904 , n383912 , n383918 );
nor ( n383920 , n383879 , n383919 );
nand ( n383921 , n383846 , n383920 );
buf ( n383922 , n383921 );
buf ( n383923 , n382067 );
nor ( n383924 , n19530 , n19200 );
not ( n383925 , n383924 );
nor ( n383926 , n19527 , n383925 );
not ( n383927 , n383926 );
buf ( n383928 , n383927 );
buf ( n383929 , n383928 );
not ( n383930 , n383929 );
not ( n383931 , n383930 );
not ( n383932 , n18258 );
not ( n383933 , n18302 );
and ( n383934 , n383932 , n383933 );
not ( n383935 , RI15b5d420_1047);
or ( n383936 , n383935 , RI15b5d330_1045);
buf ( n383937 , n18764 );
buf ( n383938 , n383937 );
not ( n383939 , n383938 );
nand ( n383940 , n383936 , n383939 );
nor ( n383941 , n383934 , n383940 );
nand ( n383942 , n18268 , RI15b5d330_1045);
and ( n383943 , n18303 , n383942 );
and ( n383944 , n19494 , n383941 , n383943 );
and ( n383945 , n383944 , n18789 );
and ( n383946 , n383945 , RI15b588a8_886);
not ( n383947 , n383941 );
and ( n383948 , n19494 , n383947 , n383943 );
and ( n383949 , n383948 , n18789 );
and ( n383950 , n383949 , RI15b5a6a8_950);
nor ( n383951 , n383946 , n383950 );
buf ( n383952 , n19258 );
not ( n383953 , n383952 );
buf ( n383954 , n383953 );
and ( n383955 , n383948 , n383954 );
and ( n383956 , n383955 , RI15b5ae28_966);
buf ( n383957 , n19275 );
buf ( n383958 , n383957 );
buf ( n383959 , n383958 );
and ( n383960 , n383948 , n383959 );
and ( n383961 , n383960 , RI15b5aa68_958);
nor ( n383962 , n383956 , n383961 );
buf ( n383963 , n19267 );
buf ( n383964 , n383963 );
and ( n383965 , n383948 , n383964 );
and ( n383966 , n383965 , RI15b5b1e8_974);
buf ( n383967 , n19495 );
buf ( n383968 , n383967 );
nor ( n383969 , n383947 , n383943 );
and ( n383970 , n383969 , n383953 );
and ( n383971 , n383970 , RI15b59f28_934);
and ( n383972 , n383969 , n383963 );
and ( n383973 , n383972 , RI15b5a2e8_942);
nor ( n383974 , n383971 , n383973 );
and ( n383975 , n383969 , n18789 );
and ( n383976 , n383975 , RI15b597a8_918);
and ( n383977 , n383969 , n383957 );
and ( n383978 , n383977 , RI15b59b68_926);
nor ( n383979 , n383976 , n383978 );
nor ( n383980 , n383941 , n383943 );
not ( n383981 , n383952 );
and ( n383982 , n383980 , n383981 );
and ( n383983 , n383982 , RI15b5bd28_998);
and ( n383984 , n383980 , n383957 );
and ( n383985 , n383984 , RI15b5b968_990);
nor ( n383986 , n383983 , n383985 );
and ( n383987 , n383980 , n383963 );
and ( n383988 , n383987 , RI15b5c0e8_1006);
and ( n383989 , n383980 , n18789 );
and ( n383990 , n383989 , RI15b5b5a8_982);
nor ( n383991 , n383988 , n383990 );
nand ( n383992 , n383974 , n383979 , n383986 , n383991 );
and ( n383993 , n383968 , n383992 );
and ( n383994 , n383944 , n383958 );
and ( n383995 , n383994 , RI15b58c68_894);
nor ( n383996 , n383966 , n383993 , n383995 );
and ( n383997 , n383944 , n383954 );
and ( n383998 , n383997 , RI15b59028_902);
and ( n383999 , n383944 , n383964 );
and ( n384000 , n383999 , RI15b593e8_910);
nor ( n384001 , n383998 , n384000 );
nand ( n384002 , n383951 , n383962 , n383996 , n384001 );
not ( n384003 , n384002 );
or ( n384004 , n383931 , n384003 );
not ( n384005 , n383927 );
not ( n384006 , n19495 );
and ( n384007 , n384005 , n384006 );
not ( n384008 , n19192 );
or ( n384009 , n384008 , n383191 );
not ( n384010 , n19537 );
nand ( n384011 , n384009 , n384010 );
nor ( n384012 , n19522 , n384011 );
or ( n384013 , n384012 , n19533 );
nand ( n384014 , n384013 , n19201 );
nor ( n384015 , n384007 , n384014 );
not ( n384016 , n19564 );
nor ( n384017 , n19527 , n19562 );
not ( n384018 , n384017 );
not ( n384019 , n384018 );
nor ( n384020 , n384016 , n384019 );
and ( n384021 , n384015 , n384020 );
not ( n384022 , n384021 );
and ( n384023 , n384022 , RI15b62100_1211);
nand ( n384024 , n19523 , n383924 );
not ( n384025 , n384024 );
not ( n384026 , RI15b62100_1211);
nand ( n384027 , RI15b61c50_1201 , RI15b61cc8_1202);
not ( n384028 , RI15b61d40_1203);
nor ( n384029 , n384027 , n384028 );
nand ( n384030 , n384029 , RI15b61db8_1204);
not ( n384031 , RI15b61e30_1205);
nor ( n384032 , n384030 , n384031 );
and ( n384033 , n384032 , RI15b61ea8_1206);
nand ( n384034 , n384033 , RI15b61f20_1207);
not ( n384035 , RI15b61f98_1208);
nor ( n384036 , n384034 , n384035 );
nand ( n384037 , n384036 , RI15b62010_1209);
not ( n384038 , RI15b62088_1210);
nor ( n384039 , n384037 , n384038 );
not ( n384040 , n384039 );
not ( n384041 , n384040 );
or ( n384042 , n384026 , n384041 );
or ( n384043 , n384040 , RI15b62100_1211);
nand ( n384044 , n384042 , n384043 );
and ( n384045 , n384025 , n384044 );
nor ( n384046 , n384023 , n384045 );
nand ( n384047 , n384004 , n384046 );
buf ( n384048 , n384047 );
and ( n384049 , n22646 , RI15b45438_228);
and ( n384050 , n22648 , RI15b518a0_647);
nor ( n384051 , n384049 , n384050 );
not ( n384052 , n384051 );
buf ( n384053 , n384052 );
and ( n384054 , n383840 , n383863 );
buf ( n384055 , n21344 );
buf ( n384056 , n384055 );
nand ( n384057 , n384054 , n384056 );
not ( n384058 , n384057 );
not ( n384059 , n384058 );
buf ( n384060 , n383734 );
nand ( n384061 , n384060 , n383651 );
and ( n384062 , n384061 , n383657 );
and ( n384063 , n383800 , n384062 );
and ( n384064 , n384061 , n381395 );
nor ( n384065 , n384064 , n383657 );
nor ( n384066 , n384063 , n384065 );
buf ( n384067 , n384066 );
not ( n384068 , n383791 );
not ( n384069 , n384060 );
nand ( n384070 , n384069 , n383651 );
not ( n384071 , n384070 );
and ( n384072 , n384068 , n384071 );
and ( n384073 , n384069 , n381395 );
nor ( n384074 , n384073 , n383651 );
nor ( n384075 , n384072 , n384074 );
not ( n384076 , n384075 );
not ( n384077 , n384076 );
and ( n384078 , n383800 , n22704 );
not ( n384079 , n384078 );
or ( n384080 , n384077 , n384079 );
nand ( n384081 , n383798 , n383705 );
not ( n384082 , n383791 );
nand ( n384083 , n383716 , n383631 );
nand ( n384084 , n384083 , n383637 );
not ( n384085 , n384084 );
and ( n384086 , n384082 , n384085 );
nand ( n384087 , n384083 , n381395 );
and ( n384088 , n384087 , n383719 );
nor ( n384089 , n384086 , n384088 );
not ( n384090 , n384083 );
nand ( n384091 , n384090 , n383637 );
and ( n384092 , n384091 , n381394 , n383645 );
not ( n384093 , n384092 );
buf ( n384094 , n383788 );
nand ( n384095 , n384094 , n383755 );
not ( n384096 , n384095 );
or ( n384097 , n384093 , n384096 );
not ( n384098 , n381394 );
not ( n384099 , n384091 );
or ( n384100 , n384098 , n384099 );
nand ( n384101 , n384100 , n383713 );
nand ( n384102 , n384097 , n384101 );
not ( n384103 , n383711 );
nor ( n384104 , n384102 , n384103 );
nand ( n384105 , n384089 , n384104 );
nor ( n384106 , n384081 , n384105 );
not ( n384107 , n384106 );
nand ( n384108 , n384107 , n384078 );
nand ( n384109 , n384080 , n384108 );
and ( n384110 , n384067 , n384109 );
not ( n384111 , n384067 );
buf ( n384112 , n21794 );
buf ( n384113 , n384112 );
nand ( n384114 , n384106 , n384113 );
not ( n384115 , n384114 );
nand ( n384116 , n384115 , n384075 );
not ( n384117 , n383809 );
not ( n384118 , n384117 );
nand ( n384119 , n384116 , n384118 );
and ( n384120 , n384111 , n384119 );
nor ( n384121 , n384110 , n384120 );
not ( n384122 , n384121 );
not ( n384123 , n384122 );
or ( n384124 , n384059 , n384123 );
not ( n384125 , n383730 );
not ( n384126 , n384125 );
buf ( n384127 , n22704 );
not ( n384128 , n384127 );
not ( n384129 , n384094 );
buf ( n384130 , n383754 );
nor ( n384131 , n384129 , n384130 );
and ( n384132 , n383687 , n383744 );
not ( n384133 , n383687 );
not ( n384134 , n383744 );
and ( n384135 , n384133 , n384134 );
nor ( n384136 , n384132 , n384135 );
nand ( n384137 , n384131 , n384136 );
nor ( n384138 , n383687 , n384134 );
and ( n384139 , n384137 , n384138 );
not ( n384140 , n384137 );
and ( n384141 , n384140 , n382703 );
nor ( n384142 , n384139 , n384141 );
not ( n384143 , n384142 );
or ( n384144 , n384128 , n384143 );
not ( n384145 , n21777 );
nor ( n384146 , n382702 , n384145 );
and ( n384147 , n384138 , n384146 );
not ( n384148 , n383855 );
nor ( n384149 , n384147 , n384148 );
nand ( n384150 , n384144 , n384149 );
not ( n384151 , n384150 );
or ( n384152 , n384126 , n384151 );
not ( n384153 , n384137 );
not ( n384154 , n384138 );
and ( n384155 , n384153 , n384154 );
not ( n384156 , n384155 );
not ( n384157 , n383851 );
nand ( n384158 , n384157 , n382703 , n383730 );
nor ( n384159 , n384156 , n384158 );
nand ( n384160 , n384138 , n383730 );
nor ( n384161 , n384153 , n384160 );
nor ( n384162 , n384159 , n384161 );
nand ( n384163 , n384152 , n384162 );
buf ( n384164 , n384163 );
not ( n384165 , n383871 );
not ( n384166 , n383875 );
and ( n384167 , n384165 , n384166 );
nand ( n384168 , n384167 , n383887 );
not ( n384169 , n384168 );
and ( n384170 , n384164 , n384169 );
and ( n384171 , n384168 , n384057 , n383882 );
nor ( n384172 , n384171 , n21764 );
or ( n384173 , n383823 , n383830 );
nor ( n384174 , n384173 , n383865 );
or ( n384175 , n384172 , n384174 );
nand ( n384176 , n384175 , n18154 );
not ( n384177 , RI15b4c2d8_464);
and ( n384178 , n383815 , n384177 );
nand ( n384179 , n384178 , n17998 );
or ( n384180 , n383832 , n384179 );
nand ( n384181 , n384176 , n384180 );
and ( n384182 , n384181 , n383901 );
or ( n384183 , n384182 , n20859 );
buf ( n384184 , n381329 );
buf ( n384185 , n384184 );
buf ( n384186 , n384185 );
not ( n384187 , n384186 );
not ( n384188 , n384180 );
nor ( n384189 , n384174 , n384188 );
or ( n384190 , n384172 , n384189 );
or ( n384191 , n384187 , n384190 );
not ( n384192 , n18125 );
or ( n384193 , n384192 , n383916 );
or ( n384194 , n384180 , n384193 );
nand ( n384195 , n384183 , n384191 , n384194 );
nor ( n384196 , n384170 , n384195 );
nand ( n384197 , n384124 , n384196 );
buf ( n384198 , n384197 );
buf ( n384199 , RI15b3ea48_2);
buf ( n384200 , n384199 );
buf ( n384201 , n22740 );
buf ( n384202 , n379847 );
buf ( n384203 , RI15b3ea48_2);
buf ( n384204 , n384203 );
buf ( n384205 , RI15b477d8_304);
or ( n384206 , n22315 , n380909 );
and ( n384207 , n22326 , n380913 );
not ( n384208 , RI15b41e50_113);
or ( n384209 , n380928 , n384208 );
or ( n384210 , n22334 , n380933 );
or ( n384211 , n380926 , n22336 );
nand ( n384212 , n384209 , n384210 , n384211 );
nor ( n384213 , n384207 , n384212 );
nand ( n384214 , n384206 , n384213 );
buf ( n384215 , n384214 );
buf ( n384216 , n382071 );
buf ( n384217 , n381006 );
buf ( n384218 , RI15b3e9d0_1);
buf ( n384219 , n384218 );
not ( n384220 , n380798 );
nand ( n384221 , n384220 , RI15b5c7f0_1021);
nand ( n384222 , RI15b5c868_1022 , RI15b5c8e0_1023);
not ( n384223 , RI15b5c958_1024);
nor ( n384224 , n384222 , n384223 );
nand ( n384225 , n384224 , RI15b5c9d0_1025);
not ( n384226 , RI15b5ca48_1026);
or ( n384227 , n384225 , n384226 );
nor ( n384228 , n384221 , n384227 );
and ( n384229 , n384228 , RI15b5cac0_1027);
nand ( n384230 , n384229 , RI15b5c3b8_1012);
not ( n384231 , n384230 );
buf ( n384232 , n384231 );
nand ( n384233 , RI15b5cb38_1028 , RI15b5cbb0_1029);
not ( n384234 , RI15b5cc28_1030);
nor ( n384235 , n384233 , n384234 );
nand ( n384236 , n384235 , RI15b5cca0_1031);
not ( n384237 , RI15b5cd18_1032);
nor ( n384238 , n384236 , n384237 );
nand ( n384239 , n384238 , RI15b5cd90_1033);
not ( n384240 , RI15b5ce08_1034);
nor ( n384241 , n384239 , n384240 );
nand ( n384242 , n384232 , n384241 );
not ( n384243 , n384242 );
and ( n384244 , n384243 , RI15b5ce80_1035);
nand ( n384245 , n384244 , RI15b5cef8_1036);
not ( n384246 , RI15b5cf70_1037);
and ( n384247 , n384245 , n384246 );
not ( n384248 , n384245 );
and ( n384249 , n384248 , RI15b5cf70_1037);
nor ( n384250 , n384247 , n384249 );
not ( n384251 , n384250 );
buf ( n384252 , n384232 );
not ( n384253 , n384252 );
not ( n384254 , n384253 );
or ( n384255 , n384254 , n384240 );
nor ( n384256 , n384239 , RI15b5ce08_1034);
nand ( n384257 , n384254 , n384256 );
nand ( n384258 , n384239 , RI15b5ce08_1034);
nand ( n384259 , n384255 , n384257 , n384258 );
not ( n384260 , n384259 );
not ( n384261 , n384230 );
nand ( n384262 , n384261 , RI15b5cb38_1028);
and ( n384263 , n384262 , RI15b5cbb0_1029);
not ( n384264 , n384262 );
not ( n384265 , RI15b5cbb0_1029);
and ( n384266 , n384264 , n384265 );
nor ( n384267 , n384263 , n384266 );
not ( n384268 , n384267 );
not ( n384269 , n384231 );
not ( n384270 , n384269 );
not ( n384271 , RI15b5cb38_1028);
and ( n384272 , n384270 , n384271 );
and ( n384273 , n384230 , RI15b5cb38_1028);
nor ( n384274 , n384272 , n384273 );
not ( n384275 , n384227 );
not ( n384276 , n384221 );
and ( n384277 , n384276 , RI15b5c3b8_1012);
nand ( n384278 , n384275 , n384277 );
not ( n384279 , RI15b5cac0_1027);
and ( n384280 , n384278 , n384279 );
not ( n384281 , n384278 );
and ( n384282 , n384281 , RI15b5cac0_1027);
or ( n384283 , n384280 , n384282 );
nand ( n384284 , n384274 , n384283 );
nor ( n384285 , n384268 , n384284 );
not ( n384286 , n384277 );
and ( n384287 , n384286 , RI15b5c8e0_1023);
not ( n384288 , RI15b5c868_1022);
nor ( n384289 , n384288 , RI15b5c8e0_1023);
not ( n384290 , n384289 );
not ( n384291 , n384277 );
or ( n384292 , n384290 , n384291 );
nand ( n384293 , n384288 , RI15b5c8e0_1023);
nand ( n384294 , n384292 , n384293 );
nor ( n384295 , n384287 , n384294 );
and ( n384296 , n384286 , RI15b5c958_1024);
nor ( n384297 , n384222 , RI15b5c958_1024);
not ( n384298 , n384297 );
not ( n384299 , n384277 );
or ( n384300 , n384298 , n384299 );
nand ( n384301 , n384222 , RI15b5c958_1024);
nand ( n384302 , n384300 , n384301 );
nor ( n384303 , n384296 , n384302 );
nand ( n384304 , n384295 , n384303 );
not ( n384305 , n380820 );
not ( n384306 , n384286 );
not ( n384307 , RI15b5c868_1022);
and ( n384308 , n384306 , n384307 );
and ( n384309 , n384286 , RI15b5c868_1022);
nor ( n384310 , n384308 , n384309 );
nand ( n384311 , n384305 , n384310 );
nor ( n384312 , n384304 , n384311 );
and ( n384313 , n384286 , RI15b5ca48_1026);
nor ( n384314 , n384225 , RI15b5ca48_1026);
nand ( n384315 , n384277 , n384314 );
nand ( n384316 , n384225 , RI15b5ca48_1026);
nand ( n384317 , n384315 , n384316 );
nor ( n384318 , n384313 , n384317 );
and ( n384319 , n384286 , RI15b5c9d0_1025);
not ( n384320 , n384224 );
nor ( n384321 , n384320 , RI15b5c9d0_1025);
not ( n384322 , n384321 );
not ( n384323 , n384277 );
or ( n384324 , n384322 , n384323 );
nand ( n384325 , n384320 , RI15b5c9d0_1025);
nand ( n384326 , n384324 , n384325 );
nor ( n384327 , n384319 , n384326 );
and ( n384328 , n384318 , n384327 );
nand ( n384329 , n384312 , n384328 , n19383 );
not ( n384330 , RI15b5cd18_1032);
not ( n384331 , n384230 );
or ( n384332 , n384330 , n384331 );
not ( n384333 , n384230 );
nor ( n384334 , n384236 , RI15b5cd18_1032);
and ( n384335 , n384333 , n384334 );
and ( n384336 , n384236 , RI15b5cd18_1032);
nor ( n384337 , n384335 , n384336 );
nand ( n384338 , n384332 , n384337 );
nor ( n384339 , n384329 , n384338 );
not ( n384340 , n384231 );
and ( n384341 , n384340 , RI15b5cc28_1030);
nor ( n384342 , n384233 , RI15b5cc28_1030);
not ( n384343 , n384342 );
not ( n384344 , n384231 );
or ( n384345 , n384343 , n384344 );
nand ( n384346 , n384233 , RI15b5cc28_1030);
nand ( n384347 , n384345 , n384346 );
nor ( n384348 , n384341 , n384347 );
not ( n384349 , n384333 );
and ( n384350 , n384349 , RI15b5cca0_1031);
not ( n384351 , RI15b5cca0_1031);
nand ( n384352 , n384235 , n384351 );
or ( n384353 , n384230 , n384352 );
not ( n384354 , n384235 );
nand ( n384355 , n384354 , RI15b5cca0_1031);
nand ( n384356 , n384353 , n384355 );
nor ( n384357 , n384350 , n384356 );
and ( n384358 , n384348 , n384357 );
and ( n384359 , n384285 , n384339 , n384358 );
nand ( n384360 , n19381 , n384359 );
not ( n384361 , RI15b5cd90_1033);
not ( n384362 , n384253 );
or ( n384363 , n384361 , n384362 );
not ( n384364 , n384238 );
nor ( n384365 , n384364 , RI15b5cd90_1033);
and ( n384366 , n384252 , n384365 );
not ( n384367 , RI15b5cd90_1033);
nor ( n384368 , n384238 , n384367 );
nor ( n384369 , n384366 , n384368 );
nand ( n384370 , n384363 , n384369 );
nor ( n384371 , n384360 , n384370 );
nand ( n384372 , n384260 , n384371 );
not ( n384373 , RI15b5ce80_1035);
and ( n384374 , n384242 , n384373 );
not ( n384375 , n384242 );
and ( n384376 , n384375 , RI15b5ce80_1035);
nor ( n384377 , n384374 , n384376 );
nor ( n384378 , n384372 , n384377 );
not ( n384379 , n384244 );
and ( n384380 , RI15b5cef8_1036 , n384379 );
not ( n384381 , RI15b5cef8_1036);
and ( n384382 , n384381 , n384244 );
nor ( n384383 , n384380 , n384382 );
nand ( n384384 , n384378 , n384383 );
buf ( n384385 , n384384 );
not ( n384386 , n384385 );
or ( n384387 , n384251 , n384386 );
nor ( n384388 , n384384 , n384250 );
not ( n384389 , n384388 );
nand ( n384390 , n384387 , n384389 );
buf ( n384391 , n19391 );
buf ( n384392 , n384391 );
nand ( n384393 , n384390 , n384392 );
nand ( n384394 , n380826 , RI15b5c7f0_1021);
buf ( n384395 , n384394 );
nor ( n384396 , n384395 , n384227 );
nand ( n384397 , n384396 , RI15b5cac0_1027);
not ( n384398 , n384397 );
nand ( n384399 , n384398 , n384241 );
nor ( n384400 , n384399 , n384373 );
or ( n384401 , n384400 , RI15b5cef8_1036);
nand ( n384402 , n384400 , RI15b5cef8_1036);
nand ( n384403 , n384401 , n384402 );
not ( n384404 , n384403 );
not ( n384405 , n384396 );
and ( n384406 , n384405 , RI15b5cac0_1027);
not ( n384407 , n384405 );
and ( n384408 , n384407 , n384279 );
nor ( n384409 , n384406 , n384408 );
not ( n384410 , n384409 );
or ( n384411 , n19475 , n19410 );
not ( n384412 , n384394 );
not ( n384413 , RI15b5c8e0_1023);
or ( n384414 , n384412 , n384413 );
nand ( n384415 , n384412 , n384289 );
nand ( n384416 , n384414 , n384415 , n384293 );
not ( n384417 , n384288 );
not ( n384418 , n384412 );
or ( n384419 , n384417 , n384418 );
nand ( n384420 , n384395 , RI15b5c868_1022);
nand ( n384421 , n384419 , n384420 );
nand ( n384422 , n384416 , n384421 , n380831 , n19403 );
buf ( n384423 , n384395 );
and ( n384424 , n384423 , RI15b5c9d0_1025);
not ( n384425 , n384321 );
not ( n384426 , n384412 );
or ( n384427 , n384425 , n384426 );
nand ( n384428 , n384427 , n384325 );
nor ( n384429 , n384424 , n384428 );
and ( n384430 , n384412 , n384297 );
and ( n384431 , n384395 , RI15b5c958_1024);
not ( n384432 , n384301 );
nor ( n384433 , n384430 , n384431 , n384432 );
nor ( n384434 , n384422 , n19412 , n384429 , n384433 );
nand ( n384435 , n384411 , n384434 );
and ( n384436 , n384423 , RI15b5ca48_1026);
not ( n384437 , n384314 );
not ( n384438 , n384412 );
or ( n384439 , n384437 , n384438 );
nand ( n384440 , n384439 , n384316 );
nor ( n384441 , n384436 , n384440 );
nor ( n384442 , n384435 , n384441 );
nand ( n384443 , n384410 , n384442 );
or ( n384444 , n384398 , RI15b5cb38_1028);
nand ( n384445 , n384398 , RI15b5cb38_1028);
nand ( n384446 , n384444 , n384445 );
nor ( n384447 , n384443 , n384446 );
buf ( n384448 , n384397 );
nand ( n384449 , n384448 , RI15b5ce08_1034);
nand ( n384450 , n384398 , n384256 );
nand ( n384451 , n384449 , n384450 , n384258 );
nand ( n384452 , n384448 , RI15b5cd18_1032);
nand ( n384453 , n384398 , n384334 );
not ( n384454 , n384336 );
nand ( n384455 , n384452 , n384453 , n384454 );
not ( n384456 , RI15b5cd90_1033);
not ( n384457 , n384448 );
or ( n384458 , n384456 , n384457 );
and ( n384459 , n384398 , n384365 );
nor ( n384460 , n384459 , n384368 );
nand ( n384461 , n384458 , n384460 );
or ( n384462 , n384398 , n384351 );
not ( n384463 , n384352 );
nand ( n384464 , n384398 , n384463 );
nand ( n384465 , n384462 , n384464 , n384355 );
and ( n384466 , n384451 , n384455 , n384461 , n384465 );
and ( n384467 , n384445 , n384265 );
not ( n384468 , n384445 );
and ( n384469 , n384468 , RI15b5cbb0_1029);
nor ( n384470 , n384467 , n384469 );
or ( n384471 , n384398 , n384234 );
nand ( n384472 , n384398 , n384342 );
nand ( n384473 , n384471 , n384472 , n384346 );
and ( n384474 , n384466 , n384470 , n384473 );
nand ( n384475 , n384447 , n384474 );
and ( n384476 , n384399 , RI15b5ce80_1035);
not ( n384477 , n384399 );
and ( n384478 , n384477 , n384373 );
nor ( n384479 , n384476 , n384478 );
nor ( n384480 , n384475 , n384479 );
nand ( n384481 , n384404 , n384480 );
buf ( n384482 , n384481 );
and ( n384483 , n384402 , RI15b5cf70_1037);
not ( n384484 , n384402 );
and ( n384485 , n384484 , n384246 );
nor ( n384486 , n384483 , n384485 );
and ( n384487 , n384482 , n384486 );
not ( n384488 , n384482 );
not ( n384489 , n384486 );
and ( n384490 , n384488 , n384489 );
nor ( n384491 , n384487 , n384490 );
not ( n384492 , n19501 );
buf ( n384493 , n384492 );
not ( n384494 , n384493 );
not ( n384495 , n384494 );
nand ( n384496 , n384491 , n384495 );
buf ( n384497 , n384229 );
nand ( n384498 , n384497 , n384241 );
and ( n384499 , n384498 , RI15b5ce80_1035);
not ( n384500 , n384498 );
and ( n384501 , n384500 , n384373 );
nor ( n384502 , n384499 , n384501 );
not ( n384503 , n384502 );
and ( n384504 , n18748 , n18757 , n18753 );
not ( n384505 , n384504 );
not ( n384506 , n18746 );
or ( n384507 , n384505 , n384506 );
not ( n384508 , n18444 );
nand ( n384509 , n384508 , n18757 );
buf ( n384510 , n384221 );
buf ( n384511 , n384510 );
and ( n384512 , n384511 , RI15b5c8e0_1023);
not ( n384513 , n384289 );
not ( n384514 , n384510 );
not ( n384515 , n384514 );
or ( n384516 , n384513 , n384515 );
nand ( n384517 , n384516 , n384293 );
nor ( n384518 , n384512 , n384517 );
not ( n384519 , n384510 );
buf ( n384520 , n384519 );
and ( n384521 , n384520 , n384288 );
and ( n384522 , n384510 , RI15b5c868_1022);
nor ( n384523 , n384521 , n384522 );
nor ( n384524 , n384518 , n384523 , n380805 , n18242 );
and ( n384525 , n384509 , n18373 , n384524 );
nand ( n384526 , n384507 , n384525 );
not ( n384527 , n384497 );
nand ( n384528 , n384527 , RI15b5ce08_1034);
nand ( n384529 , n384497 , n384256 );
nand ( n384530 , n384528 , n384529 , n384258 );
not ( n384531 , RI15b5cd90_1033);
not ( n384532 , n384497 );
not ( n384533 , n384532 );
or ( n384534 , n384531 , n384533 );
and ( n384535 , n384497 , n384365 );
nor ( n384536 , n384535 , n384368 );
nand ( n384537 , n384534 , n384536 );
not ( n384538 , RI15b5cd18_1032);
not ( n384539 , n384532 );
or ( n384540 , n384538 , n384539 );
and ( n384541 , n384497 , n384334 );
nor ( n384542 , n384541 , n384336 );
nand ( n384543 , n384540 , n384542 );
not ( n384544 , RI15b5c9d0_1025);
not ( n384545 , n384511 );
or ( n384546 , n384544 , n384545 );
and ( n384547 , n384519 , n384321 );
not ( n384548 , n384325 );
nor ( n384549 , n384547 , n384548 );
nand ( n384550 , n384546 , n384549 );
not ( n384551 , n384550 );
not ( n384552 , n384520 );
and ( n384553 , n384552 , RI15b5c958_1024);
not ( n384554 , n384297 );
not ( n384555 , n384514 );
or ( n384556 , n384554 , n384555 );
nand ( n384557 , n384556 , n384301 );
nor ( n384558 , n384553 , n384557 );
and ( n384559 , n384511 , RI15b5ca48_1026);
not ( n384560 , n384314 );
not ( n384561 , n384510 );
not ( n384562 , n384561 );
or ( n384563 , n384560 , n384562 );
nand ( n384564 , n384563 , n384316 );
nor ( n384565 , n384559 , n384564 );
not ( n384566 , n384228 );
and ( n384567 , n384566 , RI15b5cac0_1027);
not ( n384568 , n384566 );
and ( n384569 , n384568 , n384279 );
nor ( n384570 , n384567 , n384569 );
nor ( n384571 , n384551 , n384558 , n384565 , n384570 );
and ( n384572 , n384530 , n384537 , n384543 , n384571 );
nand ( n384573 , n384497 , RI15b5cb38_1028);
and ( n384574 , n384573 , n384265 );
not ( n384575 , n384573 );
and ( n384576 , n384575 , RI15b5cbb0_1029);
nor ( n384577 , n384574 , n384576 );
not ( n384578 , n384527 );
and ( n384579 , RI15b5cb38_1028 , n384578 );
not ( n384580 , RI15b5cb38_1028);
and ( n384581 , n384580 , n384532 );
nor ( n384582 , n384579 , n384581 );
and ( n384583 , n384577 , n384582 );
not ( n384584 , RI15b5cca0_1031);
buf ( n384585 , n384497 );
not ( n384586 , n384585 );
not ( n384587 , n384586 );
or ( n384588 , n384584 , n384587 );
and ( n384589 , n384585 , n384463 );
not ( n384590 , n384355 );
nor ( n384591 , n384589 , n384590 );
nand ( n384592 , n384588 , n384591 );
or ( n384593 , n384585 , n384234 );
nand ( n384594 , n384585 , n384342 );
nand ( n384595 , n384593 , n384594 , n384346 );
nand ( n384596 , n384572 , n384583 , n384592 , n384595 );
nor ( n384597 , n384526 , n384596 );
nand ( n384598 , n384503 , n384597 );
not ( n384599 , n384498 );
and ( n384600 , n384599 , RI15b5ce80_1035);
not ( n384601 , n384600 );
and ( n384602 , RI15b5cef8_1036 , n384601 );
not ( n384603 , RI15b5cef8_1036);
and ( n384604 , n384603 , n384600 );
nor ( n384605 , n384602 , n384604 );
nor ( n384606 , n384598 , n384605 );
not ( n384607 , n384606 );
nand ( n384608 , n384600 , RI15b5cef8_1036);
and ( n384609 , n384608 , n384246 );
not ( n384610 , n384608 );
and ( n384611 , n384610 , RI15b5cf70_1037);
nor ( n384612 , n384609 , n384611 );
not ( n384613 , n384612 );
and ( n384614 , n384607 , n384613 );
not ( n384615 , n384607 );
and ( n384616 , n384615 , n384612 );
nor ( n384617 , n384614 , n384616 );
and ( n384618 , n384617 , n380813 );
nor ( n384619 , n19512 , n379446 );
nor ( n384620 , n384618 , n384619 );
and ( n384621 , n384393 , n384496 , n384620 );
not ( n384622 , n383422 );
buf ( n384623 , n22782 );
not ( n384624 , n384623 );
not ( n384625 , n384624 );
or ( n384626 , n384622 , n384625 );
not ( n384627 , n19644 );
not ( n384628 , n383442 );
or ( n384629 , n384627 , n384628 );
buf ( n384630 , n383447 );
buf ( n384631 , n384630 );
not ( n384632 , n384631 );
nand ( n384633 , n384632 , n19642 );
nand ( n384634 , n19607 , n384633 );
not ( n384635 , n19642 );
nor ( n384636 , n384635 , RI15b630f0_1245);
nor ( n384637 , n384634 , n384636 );
nand ( n384638 , n384629 , n384637 );
not ( n384639 , n384638 );
nand ( n384640 , n19645 , n383454 );
nand ( n384641 , n384639 , n384640 );
not ( n384642 , n384641 );
nand ( n384643 , n384626 , n384642 );
nand ( n384644 , n384643 , RI15b63708_1258);
not ( n384645 , n383456 );
nor ( n384646 , n384645 , n383422 );
and ( n384647 , n384646 , RI15b63708_1258);
not ( n384648 , n384646 );
and ( n384649 , n384648 , n383423 );
nor ( n384650 , n384647 , n384649 );
and ( n384651 , n384650 , n19630 );
nand ( n384652 , n384630 , n19641 , RI15b630f0_1245);
not ( n384653 , n384652 );
not ( n384654 , n383442 );
and ( n384655 , n384653 , n384654 , RI15b634b0_1253);
nor ( n384656 , n383422 , RI15b63708_1258);
and ( n384657 , n384655 , n384656 );
nor ( n384658 , n384651 , n384657 );
nand ( n384659 , n384621 , n384644 , n384658 );
buf ( n384660 , n384659 );
and ( n384661 , n20565 , n20543 );
nor ( n384662 , n384661 , n22372 );
not ( n384663 , n384662 );
and ( n384664 , n384663 , RI15b4b798_440);
not ( n384665 , n19973 );
not ( n384666 , n384665 );
not ( n384667 , n22377 );
or ( n384668 , n384666 , n384667 );
nand ( n384669 , n384668 , n383364 );
and ( n384670 , n384669 , RI15b49998_376);
or ( n384671 , n22359 , n384665 , RI15b49998_376);
and ( n384672 , n382109 , RI15b4b798_440);
nor ( n384673 , n20543 , n382109 , RI15b4b798_440);
nor ( n384674 , n384672 , n384673 );
or ( n384675 , n20564 , n384674 );
nand ( n384676 , n384671 , n384675 );
nor ( n384677 , n384664 , n384670 , n384676 );
or ( n384678 , n384677 , n20519 );
not ( n384679 , n19807 );
buf ( n384680 , n19805 );
not ( n384681 , n384680 );
not ( n384682 , n19918 );
and ( n384683 , n384681 , n384682 );
not ( n384684 , n22350 );
nor ( n384685 , n384683 , n384684 );
or ( n384686 , n384679 , n384685 );
not ( n384687 , n20525 );
and ( n384688 , n384687 , n384680 , n384679 );
or ( n384689 , n20639 , n382110 );
not ( n384690 , RI15b4a898_408);
or ( n384691 , n384690 , n22390 );
not ( n384692 , n22395 );
nand ( n384693 , n384689 , n384691 , n384692 );
nor ( n384694 , n384688 , n384693 );
nand ( n384695 , n384678 , n384686 , n384694 );
buf ( n384696 , n384695 );
buf ( n384697 , n382049 );
buf ( n384698 , n381021 );
buf ( n384699 , n384203 );
buf ( n384700 , RI15b3e9d0_1);
buf ( n384701 , n384700 );
not ( n384702 , n383840 );
nand ( n384703 , n384702 , n383862 );
or ( n384704 , n384703 , n383894 );
not ( n384705 , n384704 );
not ( n384706 , n384705 );
not ( n384707 , n383694 );
not ( n384708 , n383800 );
or ( n384709 , n384707 , n384708 );
buf ( n384710 , n381403 );
not ( n384711 , n384710 );
nand ( n384712 , n384711 , n383688 );
nand ( n384713 , n384709 , n384712 );
nand ( n384714 , n384066 , n384075 );
not ( n384715 , n384714 );
nand ( n384716 , n384115 , n384715 );
nand ( n384717 , n384716 , n384118 );
and ( n384718 , n384713 , n384717 );
not ( n384719 , n384713 );
not ( n384720 , n384078 );
not ( n384721 , n384714 );
or ( n384722 , n384720 , n384721 );
nand ( n384723 , n384722 , n384108 );
and ( n384724 , n384719 , n384723 );
nor ( n384725 , n384718 , n384724 );
not ( n384726 , n384725 );
not ( n384727 , n384726 );
or ( n384728 , n384706 , n384727 );
nor ( n384729 , n382702 , n383730 );
not ( n384730 , n384729 );
not ( n384731 , n384156 );
not ( n384732 , n384731 );
or ( n384733 , n384730 , n384732 );
and ( n384734 , n384161 , n382702 );
nor ( n384735 , n384734 , n383851 );
nand ( n384736 , n384733 , n384735 );
not ( n384737 , n384736 );
nand ( n384738 , n383876 , n383887 );
not ( n384739 , n384738 );
and ( n384740 , n384737 , n384739 );
not ( n384741 , n383881 );
and ( n384742 , n384738 , n384704 , n384741 );
nor ( n384743 , n384742 , n21764 );
nor ( n384744 , n383885 , n383865 );
or ( n384745 , n384743 , n384744 );
nand ( n384746 , n384745 , n18154 );
or ( n384747 , n383893 , n383832 );
and ( n384748 , n384746 , n384747 );
nor ( n384749 , n384748 , n383902 );
or ( n384750 , n384749 , n20811 );
buf ( n384751 , n381378 );
buf ( n384752 , n384751 );
not ( n384753 , n384752 );
not ( n384754 , n384753 );
not ( n384755 , n384747 );
nor ( n384756 , n384744 , n384755 );
or ( n384757 , n384743 , n384756 );
or ( n384758 , n384754 , n384757 );
or ( n384759 , n379944 , n383916 );
or ( n384760 , n384747 , n384759 );
nand ( n384761 , n384750 , n384758 , n384760 );
nor ( n384762 , n384740 , n384761 );
nand ( n384763 , n384728 , n384762 );
buf ( n384764 , n384763 );
buf ( n384765 , n381707 );
buf ( n384766 , n22655 );
not ( n384767 , n380546 );
nand ( n384768 , n384767 , n380282 );
buf ( n384769 , n380547 );
and ( n384770 , n384768 , n384769 );
not ( n384771 , n384768 );
not ( n384772 , n384769 );
and ( n384773 , n384771 , n384772 );
nor ( n384774 , n384770 , n384773 );
nand ( n384775 , n384774 , n380637 );
buf ( n384776 , n380367 );
buf ( n384777 , n380375 );
nand ( n384778 , n384776 , n384777 );
buf ( n384779 , n380279 );
nand ( n384780 , n384778 , n384779 );
buf ( n384781 , n380384 );
not ( n384782 , n384781 );
and ( n384783 , n384780 , n384782 );
not ( n384784 , n384780 );
and ( n384785 , n384784 , n384781 );
nor ( n384786 , n384783 , n384785 );
buf ( n384787 , n380339 );
buf ( n384788 , n380346 );
buf ( n384789 , n380352 );
nand ( n384790 , n384787 , n384788 , n384789 );
nand ( n384791 , n384790 , n384779 );
buf ( n384792 , n380358 );
buf ( n384793 , n384792 );
not ( n384794 , n384793 );
and ( n384795 , n384791 , n384794 );
not ( n384796 , n384791 );
and ( n384797 , n384796 , n384793 );
nor ( n384798 , n384795 , n384797 );
nand ( n384799 , n384786 , n384798 );
buf ( n384800 , n380278 );
nor ( n384801 , n384776 , n384800 );
buf ( n384802 , n384777 );
and ( n384803 , n384801 , n384802 );
not ( n384804 , n384801 );
not ( n384805 , n384802 );
and ( n384806 , n384804 , n384805 );
nor ( n384807 , n384803 , n384806 );
nand ( n384808 , n384787 , n384788 );
and ( n384809 , n384808 , n380279 );
buf ( n384810 , n384789 );
and ( n384811 , n384809 , n384810 );
not ( n384812 , n384809 );
not ( n384813 , n384810 );
and ( n384814 , n384812 , n384813 );
nor ( n384815 , n384811 , n384814 );
not ( n384816 , n384788 );
not ( n384817 , n384816 );
not ( n384818 , n384787 );
not ( n384819 , n380278 );
nand ( n384820 , n384818 , n384819 );
not ( n384821 , n384820 );
or ( n384822 , n384817 , n384821 );
buf ( n384823 , n384816 );
or ( n384824 , n384820 , n384823 );
nand ( n384825 , n384822 , n384824 );
not ( n384826 , n380276 );
not ( n384827 , n380322 );
nand ( n384828 , n384826 , n384827 );
and ( n384829 , n384828 , n382955 );
not ( n384830 , n384828 );
and ( n384831 , n384830 , n382954 );
nor ( n384832 , n384829 , n384831 );
not ( n384833 , n384827 );
buf ( n384834 , n384833 );
nand ( n384835 , n384832 , n384834 );
not ( n384836 , n380296 );
not ( n384837 , n382952 );
nor ( n384838 , n384836 , n384837 );
not ( n384839 , n384838 );
not ( n384840 , n384827 );
not ( n384841 , n384840 );
or ( n384842 , n384839 , n384841 );
not ( n384843 , n380276 );
nand ( n384844 , n384842 , n384843 );
and ( n384845 , n384844 , n381611 );
not ( n384846 , n384844 );
and ( n384847 , n384846 , n381612 );
nor ( n384848 , n384845 , n384847 );
nor ( n384849 , n384835 , n384848 );
buf ( n384850 , n384836 );
not ( n384851 , n384850 );
not ( n384852 , n382953 );
not ( n384853 , n384840 );
or ( n384854 , n384852 , n384853 );
nand ( n384855 , n384854 , n384843 );
not ( n384856 , n384855 );
or ( n384857 , n384851 , n384856 );
buf ( n384858 , n384850 );
or ( n384859 , n384855 , n384858 );
nand ( n384860 , n384857 , n384859 );
not ( n384861 , n381546 );
not ( n384862 , n384861 );
not ( n384863 , n380302 );
not ( n384864 , n384833 );
or ( n384865 , n384863 , n384864 );
nand ( n384866 , n384865 , n380277 );
not ( n384867 , n384866 );
or ( n384868 , n384862 , n384867 );
or ( n384869 , n384866 , n381547 );
nand ( n384870 , n384868 , n384869 );
nor ( n384871 , n384860 , n384870 );
and ( n384872 , n380329 , n380277 );
and ( n384873 , n384872 , n380778 );
not ( n384874 , n384872 );
not ( n384875 , n380778 );
and ( n384876 , n384874 , n384875 );
nor ( n384877 , n384873 , n384876 );
nand ( n384878 , n384849 , n384871 , n384877 );
nor ( n384879 , n384825 , n384878 );
nand ( n384880 , n384807 , n384815 , n384879 );
nor ( n384881 , n384799 , n384880 );
not ( n384882 , n384781 );
nor ( n384883 , n384778 , n384882 );
nor ( n384884 , n384883 , n380281 );
buf ( n384885 , n380392 );
and ( n384886 , n384884 , n384885 );
not ( n384887 , n384884 );
not ( n384888 , n384885 );
and ( n384889 , n384887 , n384888 );
nor ( n384890 , n384886 , n384889 );
not ( n384891 , n384792 );
not ( n384892 , n384790 );
not ( n384893 , n384892 );
or ( n384894 , n384891 , n384893 );
nand ( n384895 , n384894 , n384779 );
not ( n384896 , n384895 );
not ( n384897 , n380364 );
not ( n384898 , n384897 );
and ( n384899 , n384896 , n384898 );
and ( n384900 , n384895 , n384897 );
nor ( n384901 , n384899 , n384900 );
nand ( n384902 , n384881 , n384890 , n384901 );
nand ( n384903 , n384902 , n380635 );
nand ( n384904 , n22462 , n22427 );
not ( n384905 , n384904 );
and ( n384906 , n22431 , n384905 );
and ( n384907 , n384775 , n384903 , n384906 );
not ( n384908 , n384877 );
nand ( n384909 , n384907 , n384908 );
not ( n384910 , n384774 );
nand ( n384911 , n384910 , n384903 );
nand ( n384912 , n384911 , n384906 );
buf ( n384913 , n384912 );
not ( n384914 , n384913 );
nand ( n384915 , n384914 , n380781 );
or ( n384916 , n19551 , n22427 );
nand ( n384917 , n384916 , n22470 , n19201 );
or ( n384918 , n22421 , n384917 );
nand ( n384919 , n384918 , RI15b5f388_1114);
buf ( n384920 , n22465 );
not ( n384921 , n384920 );
not ( n384922 , n384921 );
and ( n384923 , n384922 , n383522 );
nand ( n384924 , n22464 , n383523 );
buf ( n384925 , n384924 );
buf ( n384926 , n384925 );
not ( n384927 , n384926 );
nor ( n384928 , n384923 , n384927 );
not ( n384929 , n384928 );
not ( n384930 , n383529 );
and ( n384931 , n384929 , n384930 );
not ( n384932 , n22463 );
or ( n384933 , n384932 , n383523 );
not ( n384934 , n384933 );
not ( n384935 , n383529 );
nor ( n384936 , n384935 , n383522 );
and ( n384937 , n384934 , n384936 );
nor ( n384938 , n384931 , n384937 );
nand ( n384939 , n384909 , n384915 , n384919 , n384938 );
buf ( n384940 , n384939 );
buf ( n384941 , n381021 );
not ( n384942 , n22097 );
nand ( n384943 , n380957 , n380950 );
nand ( n384944 , n380952 , n380965 );
not ( n384945 , RI15b66660_1359);
and ( n384946 , n384944 , n384945 );
not ( n384947 , n384944 );
and ( n384948 , n384947 , RI15b66660_1359);
nor ( n384949 , n384946 , n384948 );
not ( n384950 , n384949 );
and ( n384951 , n384943 , n384950 );
not ( n384952 , n384943 );
and ( n384953 , n384952 , n384949 );
nor ( n384954 , n384951 , n384953 );
not ( n384955 , n384954 );
or ( n384956 , n384942 , n384955 );
not ( n384957 , n22094 );
nand ( n384958 , n384957 , RI15b66660_1359);
nand ( n384959 , n384956 , n384958 );
buf ( n384960 , n384959 );
not ( n384961 , n384960 );
or ( n384962 , n384961 , n380909 );
buf ( n384963 , n22045 );
nand ( n384964 , n384963 , RI15b666d8_1360);
and ( n384965 , n384964 , n22047 );
not ( n384966 , n384964 );
and ( n384967 , n384966 , RI15b662a0_1351);
nor ( n384968 , n384965 , n384967 );
not ( n384969 , n384968 );
not ( n384970 , n20637 );
not ( n384971 , n380970 );
nand ( n384972 , n384971 , n380980 );
not ( n384973 , n384972 );
not ( n384974 , n384973 );
or ( n384975 , n384970 , n384974 );
nand ( n384976 , n384975 , n22094 );
not ( n384977 , n384976 );
or ( n384978 , n384969 , n384977 );
not ( n384979 , n384968 );
not ( n384980 , n384973 );
nand ( n384981 , n384979 , n384980 , n22097 );
nand ( n384982 , n384978 , n384981 );
buf ( n384983 , n384982 );
and ( n384984 , n384983 , n380913 );
not ( n384985 , RI15b41fb8_116);
or ( n384986 , n380928 , n384985 );
or ( n384987 , n22022 , n380933 );
or ( n384988 , n20413 , n22298 );
or ( n384989 , n380926 , n384988 );
nand ( n384990 , n384986 , n384987 , n384989 );
nor ( n384991 , n384984 , n384990 );
nand ( n384992 , n384962 , n384991 );
buf ( n384993 , n384992 );
buf ( n384994 , RI15b47d78_316);
buf ( n384995 , n383174 );
buf ( n384996 , RI15b3e9d0_1);
buf ( n384997 , n384996 );
buf ( n384998 , n17499 );
buf ( n384999 , n382067 );
buf ( n385000 , n383840 );
nand ( n385001 , n383830 , n21337 );
or ( n385002 , n385000 , n385001 );
or ( n385003 , n383814 , n385002 );
and ( n385004 , n383871 , n384166 );
nand ( n385005 , n385004 , n383866 );
not ( n385006 , n385005 );
and ( n385007 , n383857 , n385006 );
not ( n385008 , n383880 );
not ( n385009 , n385008 );
and ( n385010 , n385005 , n385002 , n385009 );
nor ( n385011 , n385010 , n21764 );
buf ( n385012 , n383837 );
nor ( n385013 , n385012 , n383888 );
or ( n385014 , n385011 , n385013 );
nand ( n385015 , n385014 , n18154 );
nand ( n385016 , n383892 , n17998 );
or ( n385017 , n385016 , n383894 );
nand ( n385018 , n385015 , n385017 );
and ( n385019 , n385018 , n383901 );
or ( n385020 , n385019 , n21130 );
not ( n385021 , n385017 );
nor ( n385022 , n385013 , n385021 );
or ( n385023 , n385011 , n385022 );
or ( n385024 , n383908 , n385023 );
or ( n385025 , n385017 , n383917 );
nand ( n385026 , n385020 , n385024 , n385025 );
nor ( n385027 , n385007 , n385026 );
nand ( n385028 , n385003 , n385027 );
buf ( n385029 , n385028 );
buf ( n385030 , n381566 );
and ( n385031 , RI15b60c60_1167 , RI15b60cd8_1168);
not ( n385032 , RI15b3f9c0_35);
not ( n385033 , RI15b60738_1156);
and ( n385034 , n385032 , n385033 );
nand ( n385035 , RI15b60be8_1166 , RI15b60c60_1167);
nor ( n385036 , n385034 , n385035 , RI15b3fa38_36);
nor ( n385037 , n385031 , n385036 );
or ( n385038 , n385037 , n22427 );
not ( n385039 , n379785 );
nor ( n385040 , n22435 , RI15b60738_1156 , RI15b60c60_1167);
and ( n385041 , n385040 , RI15b3f9c0_35);
nor ( n385042 , n22443 , RI15b3fa38_36);
nand ( n385043 , RI15b3f9c0_35 , RI15b60cd8_1168);
nor ( n385044 , n22442 , n385043 );
nor ( n385045 , n385041 , n385042 , n385044 );
nand ( n385046 , n385038 , n385039 , n385045 );
buf ( n385047 , n385046 );
buf ( n385048 , n22402 );
buf ( n385049 , n17499 );
nand ( n385050 , n21826 , n17507 );
not ( n385051 , n385050 );
not ( n385052 , n17565 );
or ( n385053 , n385051 , n385052 );
nand ( n385054 , n385053 , n21813 );
not ( n385055 , n17576 );
buf ( n385056 , n385055 );
nor ( n385057 , n21826 , n21813 );
nand ( n385058 , n385056 , n385057 );
and ( n385059 , n18177 , RI15b57840_851);
not ( n385060 , n21953 );
or ( n385061 , n18074 , n385060 );
nand ( n385062 , n385061 , n21979 );
and ( n385063 , n385062 , RI15b55a40_787);
and ( n385064 , n18150 , RI15b57840_851);
or ( n385065 , n21982 , n21953 , RI15b55a40_787);
not ( n385066 , n21925 );
not ( n385067 , RI15b57840_851);
and ( n385068 , n385066 , n385067 );
and ( n385069 , n21925 , RI15b57840_851);
nor ( n385070 , n385068 , n385069 );
or ( n385071 , n21922 , n385070 );
nand ( n385072 , n385065 , n385071 );
nor ( n385073 , n385063 , n385064 , n385072 );
nor ( n385074 , n385073 , n18078 );
not ( n385075 , RI15b56940_819);
or ( n385076 , n18218 , n385075 );
nand ( n385077 , n385076 , n21750 );
nor ( n385078 , n385059 , n385074 , n385077 );
nand ( n385079 , n385054 , n385058 , n385078 );
buf ( n385080 , n385079 );
buf ( n385081 , n381707 );
buf ( n385082 , n18226 );
not ( n385083 , RI15b566e8_814);
not ( n385084 , n385055 );
or ( n385085 , n385083 , n385084 );
nand ( n385086 , n385085 , n18218 );
nand ( n385087 , n385086 , RI15b56760_815);
not ( n385088 , n379931 );
not ( n385089 , n385088 );
not ( n385090 , n17565 );
or ( n385091 , n385089 , n385090 );
not ( n385092 , RI15b56760_815);
nand ( n385093 , n385091 , n385092 );
and ( n385094 , n18179 , RI15b57660_847);
not ( n385095 , RI15b55860_783);
and ( n385096 , n385095 , RI15b557e8_782);
not ( n385097 , RI15b557e8_782);
and ( n385098 , n385097 , RI15b55860_783);
nor ( n385099 , n385096 , n385098 );
or ( n385100 , n18197 , n385099 );
buf ( n385101 , n20730 );
buf ( n385102 , n385101 );
not ( n385103 , n385102 );
or ( n385104 , n385103 , n379924 );
and ( n385105 , n18103 , RI15b55860_783);
and ( n385106 , n18188 , n379363 );
nor ( n385107 , n385105 , n385106 );
nand ( n385108 , n385100 , n385104 , n385107 );
nor ( n385109 , n385094 , n385108 );
nand ( n385110 , n385087 , n385093 , n385109 );
buf ( n385111 , n385110 );
buf ( n385112 , RI15b3e9d0_1);
buf ( n385113 , n385112 );
nand ( n385114 , n21636 , n21663 );
nor ( n385115 , n385114 , n21691 );
not ( n385116 , n21685 );
and ( n385117 , n385115 , n385116 );
not ( n385118 , n21679 );
nand ( n385119 , n385117 , n385118 );
not ( n385120 , n21668 );
nor ( n385121 , n385119 , n385120 );
nand ( n385122 , n385121 , n21716 );
not ( n385123 , n21710 );
nor ( n385124 , n385122 , n385123 );
buf ( n385125 , n385124 );
buf ( n385126 , n385125 );
nor ( n385127 , n385126 , n21705 );
not ( n385128 , n385127 );
nand ( n385129 , n385124 , n21705 );
buf ( n385130 , n385129 );
buf ( n385131 , n385130 );
nand ( n385132 , n385128 , n385131 );
not ( n385133 , n21745 );
buf ( n385134 , n385133 );
buf ( n385135 , n385134 );
nand ( n385136 , n385132 , n385135 );
not ( n385137 , n20718 );
not ( n385138 , n21293 );
or ( n385139 , n385137 , n385138 );
or ( n385140 , n21293 , n20718 );
nand ( n385141 , n385139 , n385140 );
and ( n385142 , n385141 , n21357 );
not ( n385143 , n21505 );
not ( n385144 , n21509 );
and ( n385145 , n385143 , n385144 );
and ( n385146 , n21505 , n21509 );
nor ( n385147 , n385145 , n385146 );
buf ( n385148 , n21561 );
or ( n385149 , n385147 , n385148 );
or ( n385150 , n21750 , n21941 );
nand ( n385151 , n385149 , n385150 );
nor ( n385152 , n385142 , n385151 );
nand ( n385153 , n385136 , n385152 );
not ( n385154 , n385153 );
or ( n385155 , n18143 , n18182 );
nand ( n385156 , n385155 , n382547 );
nand ( n385157 , n385156 , n18077 );
or ( n385158 , n379996 , n379988 );
nand ( n385159 , n385158 , n382540 );
not ( n385160 , n21783 );
nor ( n385161 , n383164 , n18168 );
and ( n385162 , n385159 , n385160 , n385161 , n18164 );
and ( n385163 , n385157 , n385162 );
not ( n385164 , n385163 );
and ( n385165 , n385164 , RI15b50658_608);
nand ( n385166 , n18142 , n18096 );
or ( n385167 , n385166 , n18181 );
nand ( n385168 , n385167 , n18126 );
nand ( n385169 , n385168 , n18077 );
and ( n385170 , n385169 , n381400 , n382691 );
or ( n385171 , n20718 , n385170 );
buf ( n385172 , n381468 );
buf ( n385173 , n385172 );
buf ( n385174 , n385173 );
not ( n385175 , n385174 );
or ( n385176 , n385175 , n21705 );
or ( n385177 , n382885 , n380008 );
not ( n385178 , n385177 );
or ( n385179 , n21509 , n385178 );
nand ( n385180 , n385171 , n385176 , n385179 );
nor ( n385181 , n385165 , n385180 );
nand ( n385182 , n385154 , n385181 );
buf ( n385183 , n385182 );
buf ( n385184 , n379895 );
not ( n385185 , RI15b5e848_1090);
not ( n385186 , n379795 );
or ( n385187 , n385185 , n385186 );
and ( n385188 , n385039 , n22441 );
not ( n385189 , RI15b60828_1158);
or ( n385190 , n385188 , n385189 );
nand ( n385191 , n385187 , n385190 );
buf ( n385192 , n385191 );
buf ( n385193 , n379802 );
buf ( n385194 , n382067 );
buf ( n385195 , RI15b3ea48_2);
buf ( n385196 , n385195 );
buf ( n385197 , RI15b3e9d0_1);
buf ( n385198 , n385197 );
buf ( n385199 , n380865 );
not ( n385200 , RI15b470d0_289);
buf ( n385201 , n20580 );
nand ( n385202 , n385201 , n20501 );
nand ( n385203 , n20613 , n385202 );
buf ( n385204 , n20585 );
not ( n385205 , n385204 );
nor ( n385206 , n385205 , n20519 , n20515 );
or ( n385207 , n22232 , n20634 );
nand ( n385208 , n20628 , n20651 );
nor ( n385209 , n19912 , n20635 );
not ( n385210 , n385209 );
or ( n385211 , n385206 , n385207 , n385208 , n385210 );
nor ( n385212 , n385203 , n385211 );
not ( n385213 , n385212 );
not ( n385214 , n385213 );
or ( n385215 , n385200 , n385214 );
not ( n385216 , n385205 );
not ( n385217 , n382510 );
nor ( n385218 , RI15b48318_328 , RI15b48390_329);
nand ( n385219 , n385218 , RI15b48408_330);
nand ( n385220 , n385217 , n385219 );
and ( n385221 , n385216 , n379824 , n385220 );
and ( n385222 , n385221 , RI15b48660_335);
and ( n385223 , n20631 , RI15b46950_273);
nor ( n385224 , n385222 , n385223 );
nand ( n385225 , n385215 , n385224 );
buf ( n385226 , n385225 );
nand ( n385227 , RI15b43bd8_176 , RI15b43c50_177);
not ( n385228 , RI15b43cc8_178);
nor ( n385229 , n385227 , n385228 );
nand ( n385230 , n385229 , RI15b43b60_175);
not ( n385231 , RI15b43d40_179);
nor ( n385232 , n385230 , n385231 );
nand ( n385233 , n385232 , RI15b43db8_180);
not ( n385234 , RI15b43e30_181);
nor ( n385235 , n385233 , n385234 );
nand ( n385236 , n385235 , RI15b43ea8_182);
not ( n385237 , RI15b43f20_183);
nor ( n385238 , n385236 , n385237 );
nand ( n385239 , n385238 , RI15b43f98_184);
not ( n385240 , RI15b44010_185);
nor ( n385241 , n385239 , n385240 );
buf ( n385242 , n385241 );
not ( n385243 , n385242 );
not ( n385244 , n385243 );
not ( n385245 , n385244 );
buf ( n385246 , n385245 );
buf ( n385247 , n385246 );
nand ( n385248 , n385247 , RI15b44268_190);
not ( n385249 , n385247 );
nand ( n385250 , RI15b44088_186 , RI15b44100_187);
not ( n385251 , RI15b44178_188);
nor ( n385252 , n385250 , n385251 );
nand ( n385253 , n385252 , RI15b441f0_189);
nor ( n385254 , n385253 , RI15b44268_190);
nand ( n385255 , n385249 , n385254 );
nand ( n385256 , n385253 , RI15b44268_190);
and ( n385257 , n385248 , n385255 , n385256 );
not ( n385258 , n385257 );
not ( n385259 , RI15b44a60_207);
nand ( n385260 , n385259 , RI15b449e8_206);
nand ( n385261 , n20032 , n385260 );
nand ( n385262 , n385261 , n20429 );
not ( n385263 , n385262 );
not ( n385264 , n385263 );
nand ( n385265 , RI15b449e8_206 , RI15b44a60_207);
not ( n385266 , n385265 );
and ( n385267 , n385266 , RI15b44ad8_208);
not ( n385268 , n385266 );
not ( n385269 , RI15b44ad8_208);
and ( n385270 , n385268 , n385269 );
nor ( n385271 , n385267 , n385270 );
buf ( n385272 , n385271 );
nand ( n385273 , RI15b449e8_206 , RI15b44a60_207 , RI15b44ad8_208);
and ( n385274 , n385273 , RI15b44b50_209);
not ( n385275 , n385273 );
not ( n385276 , RI15b44b50_209);
and ( n385277 , n385275 , n385276 );
nor ( n385278 , n385274 , n385277 );
nand ( n385279 , n385272 , n385278 );
nor ( n385280 , n385264 , n385279 );
buf ( n385281 , n385280 );
and ( n385282 , n385281 , RI15b41c70_109);
nand ( n385283 , n385272 , n385278 , n383372 );
not ( n385284 , n385283 );
and ( n385285 , n385284 , RI15b41130_85);
nor ( n385286 , n385282 , n385285 );
not ( n385287 , n385271 );
and ( n385288 , n385287 , n385278 , n20420 );
buf ( n385289 , n385288 );
not ( n385290 , n385289 );
not ( n385291 , n385290 );
not ( n385292 , RI15b405f0_61);
not ( n385293 , n385292 );
and ( n385294 , n385291 , n385293 );
not ( n385295 , n385273 );
and ( n385296 , n385295 , RI15b44b50_209);
not ( n385297 , n385295 );
not ( n385298 , RI15b44b50_209);
and ( n385299 , n385297 , n385298 );
nor ( n385300 , n385296 , n385299 );
nand ( n385301 , n385272 , n385300 );
not ( n385302 , n385263 );
nor ( n385303 , n385301 , n385302 );
and ( n385304 , n385303 , RI15b43a70_173);
nor ( n385305 , n385294 , n385304 );
and ( n385306 , n385287 , n385278 , n20054 );
buf ( n385307 , n385306 );
nand ( n385308 , n385307 , RI15b409b0_69);
nand ( n385309 , n385272 , n385278 , n20054 );
not ( n385310 , n385309 );
not ( n385311 , RI15b418b0_101);
not ( n385312 , n385311 );
and ( n385313 , n385310 , n385312 );
and ( n385314 , n383375 , RI15b40230_53);
nor ( n385315 , n385313 , n385314 );
nand ( n385316 , n385271 , n385278 , n20420 );
not ( n385317 , n385316 );
nand ( n385318 , n385317 , RI15b414f0_93);
and ( n385319 , n385315 , n385318 );
nand ( n385320 , n385286 , n385305 , n385308 , n385319 );
and ( n385321 , n385272 , n385300 , n20420 );
buf ( n385322 , n385321 );
and ( n385323 , n385322 , RI15b432f0_157);
not ( n385324 , n20014 );
and ( n385325 , n385272 , n385300 , n385324 );
buf ( n385326 , n385325 );
and ( n385327 , n385326 , RI15b436b0_165);
nor ( n385328 , n385323 , n385327 );
not ( n385329 , n385262 );
not ( n385330 , n20002 );
not ( n385331 , RI15b44ad8_208);
nand ( n385332 , n385331 , RI15b44b50_209);
nor ( n385333 , n385330 , n385332 );
buf ( n385334 , n385333 );
and ( n385335 , n385329 , n385334 );
and ( n385336 , n385335 , RI15b42b70_141);
buf ( n385337 , n20006 );
not ( n385338 , n385337 );
not ( n385339 , n385338 );
not ( n385340 , n385339 );
not ( n385341 , RI15b42f30_149);
not ( n385342 , n385341 );
and ( n385343 , n385340 , n385342 );
not ( n385344 , n20049 );
not ( n385345 , RI15b42030_117);
nor ( n385346 , n385344 , n385345 );
nor ( n385347 , n385343 , n385346 );
and ( n385348 , n385333 , n20025 );
and ( n385349 , n385348 , RI15b423f0_125);
not ( n385350 , n385260 );
nand ( n385351 , n385333 , n385350 );
not ( n385352 , n385351 );
and ( n385353 , n385352 , RI15b427b0_133);
nor ( n385354 , n385349 , n385353 );
nand ( n385355 , n385347 , n385354 );
nor ( n385356 , n385336 , n385355 );
nor ( n385357 , n385271 , n385300 );
and ( n385358 , n385357 , n385329 );
nand ( n385359 , n385358 , RI15b40d70_77);
nand ( n385360 , n385328 , n385356 , n385359 );
nor ( n385361 , n385320 , n385360 );
buf ( n385362 , n385361 );
buf ( n385363 , n385362 );
not ( n385364 , n385363 );
and ( n385365 , n385233 , n385234 );
not ( n385366 , n385233 );
and ( n385367 , n385366 , RI15b43e30_181);
nor ( n385368 , n385365 , n385367 );
and ( n385369 , n385364 , n385368 );
not ( n385370 , n385263 );
nor ( n385371 , n385370 , n385279 );
not ( n385372 , n385371 );
not ( n385373 , n385372 );
not ( n385374 , RI15b41bf8_108);
not ( n385375 , n385374 );
and ( n385376 , n385373 , n385375 );
and ( n385377 , n385317 , RI15b41478_92);
nor ( n385378 , n385376 , n385377 );
not ( n385379 , n385358 );
not ( n385380 , n385379 );
not ( n385381 , RI15b40cf8_76);
not ( n385382 , n385381 );
and ( n385383 , n385380 , n385382 );
and ( n385384 , n385321 , RI15b43278_156);
nor ( n385385 , n385383 , n385384 );
not ( n385386 , RI15b410b8_84);
not ( n385387 , n385284 );
or ( n385388 , n385386 , n385387 );
not ( n385389 , n20014 );
nand ( n385390 , n385389 , n385272 , n385278 );
not ( n385391 , n385390 );
not ( n385392 , RI15b41838_100);
not ( n385393 , n385392 );
and ( n385394 , n385391 , n385393 );
and ( n385395 , n385338 , RI15b42eb8_148);
nor ( n385396 , n385394 , n385395 );
nand ( n385397 , n385388 , n385396 );
not ( n385398 , n385397 );
not ( n385399 , n385325 );
not ( n385400 , n385399 );
nand ( n385401 , n385400 , RI15b43638_164);
nand ( n385402 , n385378 , n385385 , n385398 , n385401 );
not ( n385403 , n385303 );
not ( n385404 , n385403 );
not ( n385405 , RI15b439f8_172);
not ( n385406 , n385405 );
and ( n385407 , n385404 , n385406 );
and ( n385408 , n385289 , RI15b40578_60);
nor ( n385409 , n385407 , n385408 );
not ( n385410 , n385335 );
not ( n385411 , n385410 );
not ( n385412 , RI15b42af8_140);
not ( n385413 , n385412 );
and ( n385414 , n385411 , n385413 );
nand ( n385415 , n385348 , RI15b42378_124);
nand ( n385416 , n385352 , RI15b42738_132);
nor ( n385417 , n20096 , n383374 );
nand ( n385418 , n385417 , RI15b401b8_52);
nand ( n385419 , n20049 , RI15b41fb8_116);
nand ( n385420 , n385415 , n385416 , n385418 , n385419 );
nor ( n385421 , n385414 , n385420 );
nand ( n385422 , n385307 , RI15b40938_68);
nand ( n385423 , n385409 , n385421 , n385422 );
nor ( n385424 , n385402 , n385423 );
not ( n385425 , n385424 );
buf ( n385426 , n385425 );
buf ( n385427 , n385426 );
and ( n385428 , n385232 , RI15b43db8_180);
not ( n385429 , n385232 );
not ( n385430 , RI15b43db8_180);
and ( n385431 , n385429 , n385430 );
nor ( n385432 , n385428 , n385431 );
nand ( n385433 , n385427 , n385432 );
not ( n385434 , n385433 );
nor ( n385435 , n385369 , n385434 );
not ( n385436 , n385435 );
and ( n385437 , n385230 , n385231 );
not ( n385438 , n385230 );
and ( n385439 , n385438 , RI15b43d40_179);
nor ( n385440 , n385437 , n385439 );
buf ( n385441 , n385288 );
nand ( n385442 , n385441 , RI15b40500_59);
nand ( n385443 , n385307 , RI15b408c0_67);
and ( n385444 , n385442 , n385443 );
not ( n385445 , n385379 );
not ( n385446 , RI15b40c80_75);
not ( n385447 , n385446 );
and ( n385448 , n385445 , n385447 );
not ( n385449 , RI15b41040_83);
not ( n385450 , n385284 );
or ( n385451 , n385449 , n385450 );
not ( n385452 , RI15b417c0_99);
or ( n385453 , n385390 , n385452 );
nand ( n385454 , n385451 , n385453 );
nor ( n385455 , n385448 , n385454 );
not ( n385456 , n385372 );
not ( n385457 , RI15b41b80_107);
not ( n385458 , n385457 );
and ( n385459 , n385456 , n385458 );
not ( n385460 , RI15b40140_51);
not ( n385461 , n383375 );
or ( n385462 , n385460 , n385461 );
not ( n385463 , n385317 );
or ( n385464 , n385463 , n20363 );
nand ( n385465 , n385462 , n385464 );
nor ( n385466 , n385459 , n385465 );
nand ( n385467 , n385444 , n385455 , n385466 );
not ( n385468 , RI15b435c0_163);
nor ( n385469 , n385399 , n385468 );
not ( n385470 , n385301 );
buf ( n385471 , n20420 );
nand ( n385472 , n385470 , n385471 );
nor ( n385473 , n385472 , n20337 );
nor ( n385474 , n385469 , n385473 );
not ( n385475 , RI15b42a80_139);
nor ( n385476 , n385410 , n385475 );
nand ( n385477 , n385348 , RI15b42300_123);
nand ( n385478 , n385352 , RI15b426c0_131);
and ( n385479 , n385477 , n385478 );
not ( n385480 , n385337 );
not ( n385481 , n20334 );
and ( n385482 , n385480 , n385481 );
not ( n385483 , n20049 );
nor ( n385484 , n385483 , n380988 );
nor ( n385485 , n385482 , n385484 );
nand ( n385486 , n385479 , n385485 );
nor ( n385487 , n385476 , n385486 );
nand ( n385488 , n385303 , RI15b43980_171);
nand ( n385489 , n385474 , n385487 , n385488 );
nor ( n385490 , n385467 , n385489 );
not ( n385491 , n385490 );
buf ( n385492 , n385491 );
buf ( n385493 , n385492 );
xor ( n385494 , n385440 , n385493 );
nand ( n385495 , n385441 , RI15b40488_58);
nand ( n385496 , n385307 , RI15b40848_66);
and ( n385497 , n385495 , n385496 );
not ( n385498 , n385379 );
not ( n385499 , RI15b40c08_74);
not ( n385500 , n385499 );
and ( n385501 , n385498 , n385500 );
not ( n385502 , RI15b40fc8_82);
not ( n385503 , n385284 );
or ( n385504 , n385502 , n385503 );
not ( n385505 , RI15b41748_98);
or ( n385506 , n385309 , n385505 );
nand ( n385507 , n385504 , n385506 );
nor ( n385508 , n385501 , n385507 );
not ( n385509 , n385280 );
not ( n385510 , n385509 );
not ( n385511 , RI15b41b08_106);
not ( n385512 , n385511 );
and ( n385513 , n385510 , n385512 );
not ( n385514 , RI15b400c8_50);
not ( n385515 , n383375 );
or ( n385516 , n385514 , n385515 );
not ( n385517 , RI15b41388_90);
or ( n385518 , n385463 , n385517 );
nand ( n385519 , n385516 , n385518 );
nor ( n385520 , n385513 , n385519 );
nand ( n385521 , n385497 , n385508 , n385520 );
nand ( n385522 , n385303 , RI15b43908_170);
nand ( n385523 , n385335 , RI15b42a08_138);
not ( n385524 , n385348 );
not ( n385525 , RI15b42288_122);
or ( n385526 , n385524 , n385525 );
not ( n385527 , RI15b42648_130);
or ( n385528 , n385351 , n385527 );
nand ( n385529 , n385526 , n385528 );
not ( n385530 , RI15b42dc8_146);
not ( n385531 , n20007 );
or ( n385532 , n385530 , n385531 );
nand ( n385533 , n20049 , RI15b41ec8_114);
nand ( n385534 , n385532 , n385533 );
nor ( n385535 , n385529 , n385534 );
and ( n385536 , n385522 , n385523 , n385535 );
nand ( n385537 , n385326 , RI15b43548_162);
nand ( n385538 , n385321 , RI15b43188_154);
and ( n385539 , n385537 , n385538 );
nand ( n385540 , n385536 , n385539 );
nor ( n385541 , n385521 , n385540 );
not ( n385542 , n385541 );
buf ( n385543 , n385542 );
not ( n385544 , n385543 );
not ( n385545 , RI15b43b60_175);
nor ( n385546 , n385545 , n385227 );
and ( n385547 , n385546 , n385228 );
not ( n385548 , n385546 );
and ( n385549 , n385548 , RI15b43cc8_178);
nor ( n385550 , n385547 , n385549 );
nand ( n385551 , n385544 , n385550 );
not ( n385552 , n385551 );
nand ( n385553 , RI15b43b60_175 , RI15b43bd8_176);
not ( n385554 , RI15b43c50_177);
and ( n385555 , n385553 , n385554 );
not ( n385556 , n385553 );
and ( n385557 , n385556 , RI15b43c50_177);
nor ( n385558 , n385555 , n385557 );
not ( n385559 , n385558 );
nand ( n385560 , n385358 , RI15b40b90_73);
nand ( n385561 , n385307 , RI15b407d0_65);
and ( n385562 , n385560 , n385561 );
and ( n385563 , n385280 , RI15b41a90_105);
and ( n385564 , n385284 , RI15b40f50_81);
nor ( n385565 , n385563 , n385564 );
not ( n385566 , n385290 );
nand ( n385567 , n385566 , RI15b40410_57);
nand ( n385568 , n385317 , RI15b41310_89);
not ( n385569 , n385309 );
nand ( n385570 , n385569 , RI15b416d0_97);
nand ( n385571 , n383375 , RI15b40050_49);
and ( n385572 , n385568 , n385570 , n385571 );
nand ( n385573 , n385562 , n385565 , n385567 , n385572 );
not ( n385574 , RI15b42990_137);
or ( n385575 , n385410 , n385574 );
nand ( n385576 , n385348 , RI15b42210_121);
nand ( n385577 , n385352 , RI15b425d0_129);
and ( n385578 , n385576 , n385577 );
not ( n385579 , n385337 );
nand ( n385580 , n385579 , RI15b42d50_145);
nand ( n385581 , n20049 , RI15b41e50_113);
and ( n385582 , n385580 , n385581 );
nand ( n385583 , n385575 , n385578 , n385582 );
nor ( n385584 , n385472 , n20169 );
nor ( n385585 , n385583 , n385584 );
nand ( n385586 , n385303 , RI15b43890_169);
nand ( n385587 , n385326 , RI15b434d0_161);
and ( n385588 , n385586 , n385587 );
nand ( n385589 , n385585 , n385588 );
nor ( n385590 , n385573 , n385589 );
not ( n385591 , n385590 );
not ( n385592 , n385591 );
nand ( n385593 , n385559 , n385592 );
not ( n385594 , n385593 );
not ( n385595 , RI15b40398_56);
not ( n385596 , n385441 );
or ( n385597 , n385595 , n385596 );
not ( n385598 , n385263 );
nor ( n385599 , n385301 , n385598 );
nand ( n385600 , n385599 , RI15b43818_168);
nand ( n385601 , n385597 , n385600 );
not ( n385602 , RI15b40ed8_80);
not ( n385603 , n385284 );
or ( n385604 , n385602 , n385603 );
not ( n385605 , n385309 );
not ( n385606 , RI15b41658_96);
not ( n385607 , n385606 );
and ( n385608 , n385605 , n385607 );
and ( n385609 , n383375 , RI15b3ffd8_48);
nor ( n385610 , n385608 , n385609 );
nand ( n385611 , n385604 , n385610 );
nor ( n385612 , n385601 , n385611 );
not ( n385613 , RI15b41a18_104);
not ( n385614 , n385280 );
or ( n385615 , n385613 , n385614 );
nand ( n385616 , n385317 , RI15b41298_88);
nand ( n385617 , n385615 , n385616 );
not ( n385618 , n385306 );
not ( n385619 , RI15b40758_64);
nor ( n385620 , n385618 , n385619 );
nor ( n385621 , n385617 , n385620 );
not ( n385622 , RI15b40b18_72);
nor ( n385623 , n385379 , n385622 );
not ( n385624 , RI15b42918_136);
not ( n385625 , n385335 );
or ( n385626 , n385624 , n385625 );
not ( n385627 , RI15b42198_120);
not ( n385628 , n385348 );
or ( n385629 , n385627 , n385628 );
nand ( n385630 , n385352 , RI15b42558_128);
nand ( n385631 , n385629 , n385630 );
not ( n385632 , RI15b41dd8_112);
or ( n385633 , n385483 , n385632 );
not ( n385634 , n20007 );
or ( n385635 , n385634 , n20075 );
nand ( n385636 , n385633 , n385635 );
nor ( n385637 , n385631 , n385636 );
nand ( n385638 , n385626 , n385637 );
nor ( n385639 , n385623 , n385638 );
and ( n385640 , n385322 , RI15b43098_152);
and ( n385641 , n385400 , RI15b43458_160);
nor ( n385642 , n385640 , n385641 );
and ( n385643 , n385612 , n385621 , n385639 , n385642 );
or ( n385644 , RI15b43b60_175 , RI15b43bd8_176);
nand ( n385645 , n385644 , n385553 );
nand ( n385646 , n385643 , n385645 );
not ( n385647 , n385646 );
not ( n385648 , RI15b406e0_63);
not ( n385649 , n385306 );
or ( n385650 , n385648 , n385649 );
nand ( n385651 , n385358 , RI15b40aa0_71);
nand ( n385652 , n385650 , n385651 );
not ( n385653 , RI15b40320_55);
not ( n385654 , n385288 );
or ( n385655 , n385653 , n385654 );
nand ( n385656 , n385417 , RI15b3ff60_47);
nand ( n385657 , n385655 , n385656 );
nor ( n385658 , n385652 , n385657 );
not ( n385659 , RI15b433e0_159);
not ( n385660 , n385325 );
or ( n385661 , n385659 , n385660 );
nand ( n385662 , n385599 , RI15b437a0_167);
nand ( n385663 , n385661 , n385662 );
not ( n385664 , RI15b419a0_103);
not ( n385665 , n385371 );
or ( n385666 , n385664 , n385665 );
not ( n385667 , n385283 );
nand ( n385668 , n385667 , RI15b40e60_79);
nand ( n385669 , n385666 , n385668 );
nor ( n385670 , n385663 , n385669 );
not ( n385671 , RI15b43020_151);
not ( n385672 , n385321 );
or ( n385673 , n385671 , n385672 );
nand ( n385674 , n385348 , RI15b42120_119);
nand ( n385675 , n385352 , RI15b424e0_127);
not ( n385676 , n20006 );
not ( n385677 , n20314 );
and ( n385678 , n385676 , n385677 );
not ( n385679 , RI15b41d60_111);
nor ( n385680 , n20048 , n385679 );
nor ( n385681 , n385678 , n385680 );
nand ( n385682 , n385674 , n385675 , n385681 );
not ( n385683 , RI15b41220_87);
nor ( n385684 , n385316 , n385683 );
nor ( n385685 , n385682 , n385684 );
nand ( n385686 , n385673 , n385685 );
not ( n385687 , RI15b428a0_135);
not ( n385688 , n385335 );
or ( n385689 , n385687 , n385688 );
not ( n385690 , n385390 );
nand ( n385691 , n385690 , RI15b415e0_95);
nand ( n385692 , n385689 , n385691 );
nor ( n385693 , n385686 , n385692 );
nand ( n385694 , n385658 , n385670 , n385693 );
not ( n385695 , n385694 );
not ( n385696 , n385695 );
not ( n385697 , n385696 );
not ( n385698 , RI15b43368_158);
not ( n385699 , n385325 );
or ( n385700 , n385698 , n385699 );
nand ( n385701 , n385599 , RI15b43728_166);
nand ( n385702 , n385700 , n385701 );
or ( n385703 , n385472 , n20234 );
nand ( n385704 , n385338 , RI15b42be8_142);
nand ( n385705 , n385703 , n385704 );
nor ( n385706 , n385702 , n385705 );
not ( n385707 , RI15b41928_102);
not ( n385708 , n385371 );
or ( n385709 , n385707 , n385708 );
and ( n385710 , n385317 , RI15b411a8_86);
not ( n385711 , RI15b41568_94);
nor ( n385712 , n385390 , n385711 );
nor ( n385713 , n385710 , n385712 );
nand ( n385714 , n385709 , n385713 );
not ( n385715 , RI15b42828_134);
not ( n385716 , n385335 );
or ( n385717 , n385715 , n385716 );
not ( n385718 , RI15b420a8_118);
not ( n385719 , n385348 );
or ( n385720 , n385718 , n385719 );
nand ( n385721 , n385352 , RI15b42468_126);
nand ( n385722 , n385720 , n385721 );
not ( n385723 , RI15b3fee8_46);
not ( n385724 , n385417 );
or ( n385725 , n385723 , n385724 );
not ( n385726 , n20048 );
nand ( n385727 , n385726 , RI15b41ce8_110);
nand ( n385728 , n385725 , n385727 );
nor ( n385729 , n385722 , n385728 );
nand ( n385730 , n385717 , n385729 );
nor ( n385731 , n385714 , n385730 );
and ( n385732 , n385358 , RI15b40a28_70);
and ( n385733 , n385307 , RI15b40668_62);
nor ( n385734 , n385732 , n385733 );
and ( n385735 , n385441 , RI15b402a8_54);
and ( n385736 , n385284 , RI15b40de8_78);
nor ( n385737 , n385735 , n385736 );
nand ( n385738 , n385706 , n385731 , n385734 , n385737 );
nand ( n385739 , n385738 , RI15b43ae8_174);
not ( n385740 , n385739 );
not ( n385741 , n385740 );
or ( n385742 , n385697 , n385741 );
not ( n385743 , n385695 );
not ( n385744 , n385739 );
or ( n385745 , n385743 , n385744 );
nand ( n385746 , n385745 , n385545 );
nand ( n385747 , n385742 , n385746 );
not ( n385748 , n385747 );
or ( n385749 , n385647 , n385748 );
not ( n385750 , n385643 );
not ( n385751 , n385645 );
nand ( n385752 , n385750 , n385751 );
nand ( n385753 , n385749 , n385752 );
not ( n385754 , n385753 );
or ( n385755 , n385594 , n385754 );
not ( n385756 , n385592 );
nand ( n385757 , n385756 , n385558 );
nand ( n385758 , n385755 , n385757 );
not ( n385759 , n385758 );
or ( n385760 , n385552 , n385759 );
not ( n385761 , n385550 );
nand ( n385762 , n385543 , n385761 );
nand ( n385763 , n385760 , n385762 );
and ( n385764 , n385494 , n385763 );
and ( n385765 , n385440 , n385493 );
or ( n385766 , n385764 , n385765 );
not ( n385767 , n385432 );
not ( n385768 , n385427 );
nand ( n385769 , n385767 , n385768 );
nand ( n385770 , n385766 , n385769 );
not ( n385771 , n385770 );
or ( n385772 , n385436 , n385771 );
or ( n385773 , n385250 , RI15b44178_188);
or ( n385774 , n385243 , n385773 );
not ( n385775 , n385243 );
not ( n385776 , n385775 );
nand ( n385777 , n385776 , RI15b44178_188);
nand ( n385778 , n385250 , RI15b44178_188);
nand ( n385779 , n385774 , n385777 , n385778 );
not ( n385780 , RI15b44100_187);
not ( n385781 , n385245 );
or ( n385782 , n385780 , n385781 );
not ( n385783 , RI15b44100_187);
nand ( n385784 , n385783 , RI15b44088_186);
not ( n385785 , n385784 );
and ( n385786 , n385244 , n385785 );
not ( n385787 , RI15b44088_186);
nand ( n385788 , n385787 , RI15b44100_187);
not ( n385789 , n385788 );
nor ( n385790 , n385786 , n385789 );
nand ( n385791 , n385782 , n385790 );
and ( n385792 , n385775 , RI15b44088_186);
not ( n385793 , n385775 );
and ( n385794 , n385793 , n385787 );
nor ( n385795 , n385792 , n385794 );
not ( n385796 , n385368 );
and ( n385797 , n385363 , n385796 );
and ( n385798 , n385236 , n385237 );
not ( n385799 , n385236 );
and ( n385800 , n385799 , RI15b43f20_183);
nor ( n385801 , n385798 , n385800 );
not ( n385802 , n385235 );
not ( n385803 , RI15b43ea8_182);
and ( n385804 , n385802 , n385803 );
not ( n385805 , n385802 );
and ( n385806 , n385805 , RI15b43ea8_182);
nor ( n385807 , n385804 , n385806 );
nand ( n385808 , n385801 , n385807 );
not ( n385809 , n385808 );
not ( n385810 , n385239 );
not ( n385811 , n385810 );
and ( n385812 , n385811 , n385240 );
not ( n385813 , n385811 );
and ( n385814 , n385813 , RI15b44010_185);
nor ( n385815 , n385812 , n385814 );
buf ( n385816 , n385238 );
not ( n385817 , n385816 );
not ( n385818 , RI15b43f98_184);
and ( n385819 , n385817 , n385818 );
not ( n385820 , n385817 );
and ( n385821 , n385820 , RI15b43f98_184);
nor ( n385822 , n385819 , n385821 );
nand ( n385823 , n385809 , n385815 , n385822 );
nor ( n385824 , n385797 , n385823 );
and ( n385825 , n385779 , n385791 , n385795 , n385824 );
nand ( n385826 , n385772 , n385825 );
and ( n385827 , n385246 , RI15b441f0_189);
not ( n385828 , RI15b441f0_189);
nand ( n385829 , n385252 , n385828 );
or ( n385830 , n385246 , n385829 );
not ( n385831 , n385252 );
nand ( n385832 , n385831 , RI15b441f0_189);
nand ( n385833 , n385830 , n385832 );
nor ( n385834 , n385827 , n385833 );
nor ( n385835 , n385826 , n385834 );
nand ( n385836 , n385258 , n385835 );
not ( n385837 , RI15b44268_190);
nor ( n385838 , n385253 , n385837 );
nand ( n385839 , n385838 , RI15b442e0_191);
not ( n385840 , n385839 );
and ( n385841 , n385840 , RI15b44358_192);
nand ( n385842 , n385242 , n385841 );
not ( n385843 , RI15b443d0_193);
nor ( n385844 , n385842 , n385843 );
buf ( n385845 , n385844 );
not ( n385846 , n385845 );
and ( n385847 , n385846 , RI15b445b0_197);
nand ( n385848 , RI15b44448_194 , RI15b444c0_195);
not ( n385849 , RI15b44538_196);
nor ( n385850 , n385848 , n385849 );
not ( n385851 , n385850 );
nor ( n385852 , n385851 , RI15b445b0_197);
not ( n385853 , n385852 );
not ( n385854 , n385844 );
or ( n385855 , n385853 , n385854 );
nand ( n385856 , n385851 , RI15b445b0_197);
nand ( n385857 , n385855 , n385856 );
nor ( n385858 , n385847 , n385857 );
not ( n385859 , n385844 );
not ( n385860 , RI15b444c0_195);
not ( n385861 , n385860 );
and ( n385862 , n385859 , n385861 );
not ( n385863 , RI15b44448_194);
nor ( n385864 , n385863 , RI15b444c0_195);
not ( n385865 , n385864 );
not ( n385866 , n385844 );
or ( n385867 , n385865 , n385866 );
nand ( n385868 , n385863 , RI15b444c0_195);
nand ( n385869 , n385867 , n385868 );
nor ( n385870 , n385862 , n385869 );
nor ( n385871 , n385858 , n385870 );
not ( n385872 , n385844 );
not ( n385873 , n385863 );
and ( n385874 , n385872 , n385873 );
buf ( n385875 , n385844 );
and ( n385876 , n385875 , n385863 );
nor ( n385877 , n385874 , n385876 );
not ( n385878 , n385776 );
not ( n385879 , n385878 );
not ( n385880 , RI15b442e0_191);
not ( n385881 , n385880 );
and ( n385882 , n385879 , n385881 );
nand ( n385883 , n385838 , n385880 );
not ( n385884 , n385883 );
not ( n385885 , n385884 );
not ( n385886 , n385244 );
or ( n385887 , n385885 , n385886 );
not ( n385888 , n385838 );
nand ( n385889 , n385888 , RI15b442e0_191);
nand ( n385890 , n385887 , n385889 );
nor ( n385891 , n385882 , n385890 );
not ( n385892 , n385878 );
not ( n385893 , RI15b44358_192);
not ( n385894 , n385893 );
and ( n385895 , n385892 , n385894 );
nor ( n385896 , n385839 , RI15b44358_192);
not ( n385897 , n385896 );
not ( n385898 , n385244 );
or ( n385899 , n385897 , n385898 );
nand ( n385900 , n385839 , RI15b44358_192);
nand ( n385901 , n385899 , n385900 );
nor ( n385902 , n385895 , n385901 );
and ( n385903 , n385842 , RI15b443d0_193);
not ( n385904 , n385842 );
and ( n385905 , n385904 , n385843 );
nor ( n385906 , n385903 , n385905 );
nor ( n385907 , n385877 , n385891 , n385902 , n385906 );
or ( n385908 , n385875 , n385849 );
nor ( n385909 , n385848 , RI15b44538_196);
nand ( n385910 , n385875 , n385909 );
nand ( n385911 , n385848 , RI15b44538_196);
nand ( n385912 , n385908 , n385910 , n385911 );
nand ( n385913 , n385871 , n385907 , n385912 );
nor ( n385914 , n385836 , n385913 );
buf ( n385915 , n385845 );
nand ( n385916 , n385850 , RI15b445b0_197);
nor ( n385917 , n385916 , RI15b44628_198);
nand ( n385918 , n385915 , n385917 );
not ( n385919 , n385915 );
nand ( n385920 , n385919 , RI15b44628_198);
nand ( n385921 , n385916 , RI15b44628_198);
and ( n385922 , n385918 , n385920 , n385921 );
not ( n385923 , n385922 );
and ( n385924 , n385914 , n385923 );
and ( n385925 , n385919 , RI15b446a0_199);
not ( n385926 , RI15b44628_198);
nor ( n385927 , n385916 , n385926 );
not ( n385928 , n385927 );
nor ( n385929 , n385928 , RI15b446a0_199);
not ( n385930 , n385929 );
not ( n385931 , n385845 );
or ( n385932 , n385930 , n385931 );
nand ( n385933 , n385928 , RI15b446a0_199);
nand ( n385934 , n385932 , n385933 );
nor ( n385935 , n385925 , n385934 );
not ( n385936 , n385935 );
nand ( n385937 , n385924 , n385936 );
buf ( n385938 , n385915 );
buf ( n385939 , n385938 );
nand ( n385940 , n385927 , RI15b446a0_199);
nor ( n385941 , n385940 , RI15b44718_200);
nand ( n385942 , n385939 , n385941 );
not ( n385943 , n385938 );
nand ( n385944 , n385943 , RI15b44718_200);
nand ( n385945 , n385940 , RI15b44718_200);
and ( n385946 , n385942 , n385944 , n385945 );
nor ( n385947 , n385937 , n385946 );
not ( n385948 , n385915 );
and ( n385949 , n385948 , RI15b44790_201);
not ( n385950 , RI15b44718_200);
nor ( n385951 , n385940 , n385950 );
not ( n385952 , n385951 );
nor ( n385953 , n385952 , RI15b44790_201);
not ( n385954 , n385953 );
not ( n385955 , n385915 );
or ( n385956 , n385954 , n385955 );
nand ( n385957 , n385952 , RI15b44790_201);
nand ( n385958 , n385956 , n385957 );
nor ( n385959 , n385949 , n385958 );
not ( n385960 , n385959 );
nand ( n385961 , n385947 , n385960 );
and ( n385962 , n385948 , RI15b44808_202);
nand ( n385963 , n385951 , RI15b44790_201);
nor ( n385964 , n385963 , RI15b44808_202);
not ( n385965 , n385964 );
not ( n385966 , n385915 );
or ( n385967 , n385965 , n385966 );
nand ( n385968 , n385963 , RI15b44808_202);
nand ( n385969 , n385967 , n385968 );
nor ( n385970 , n385962 , n385969 );
nor ( n385971 , n385961 , n385970 );
not ( n385972 , n385971 );
and ( n385973 , n385943 , RI15b44880_203);
not ( n385974 , RI15b44808_202);
nor ( n385975 , n385963 , n385974 );
not ( n385976 , n385975 );
nor ( n385977 , n385976 , RI15b44880_203);
and ( n385978 , n385938 , n385977 );
not ( n385979 , RI15b44880_203);
nor ( n385980 , n385975 , n385979 );
nor ( n385981 , n385978 , n385980 );
not ( n385982 , n385981 );
nor ( n385983 , n385973 , n385982 );
and ( n385984 , n385972 , n385983 );
not ( n385985 , n385972 );
not ( n385986 , n385983 );
and ( n385987 , n385985 , n385986 );
nor ( n385988 , n385984 , n385987 );
buf ( n385989 , n20054 );
buf ( n385990 , n385989 );
and ( n385991 , n385990 , n20422 );
buf ( n385992 , n20085 );
buf ( n385993 , n385992 );
not ( n385994 , n385993 );
and ( n385995 , n385994 , RI15b3fc90_41);
nor ( n385996 , n385991 , n385995 );
or ( n385997 , n385996 , RI15b3fd08_42);
not ( n385998 , n385471 );
buf ( n385999 , n385998 );
not ( n386000 , n385999 );
and ( n386001 , n386000 , RI15b3fc90_41);
not ( n386002 , n383373 );
buf ( n386003 , n386002 );
and ( n386004 , n386003 , n20422 );
nor ( n386005 , n386001 , n386004 );
or ( n386006 , n386005 , n20423 );
nand ( n386007 , n385997 , n386006 );
and ( n386008 , n20469 , n386007 );
nor ( n386009 , n386008 , n381040 );
and ( n386010 , n386009 , n20470 );
nor ( n386011 , n381050 , n386010 );
not ( n386012 , n385364 );
nand ( n386013 , n386011 , n386012 );
not ( n386014 , n386013 );
buf ( n386015 , n386014 );
buf ( n386016 , n386015 );
buf ( n386017 , n386016 );
buf ( n386018 , n386017 );
buf ( n386019 , n386018 );
buf ( n386020 , n386019 );
and ( n386021 , n385988 , n386020 );
nand ( n386022 , RI15b43ae8_174 , RI15b43b60_175);
not ( n386023 , RI15b43bd8_176);
nand ( n386024 , n386022 , n386023 );
nand ( n386025 , n386024 , RI15b43c50_177);
nor ( n386026 , n386025 , n385228 );
nand ( n386027 , n386026 , RI15b43d40_179);
nor ( n386028 , n386027 , n385430 );
nand ( n386029 , n386028 , RI15b43e30_181);
nor ( n386030 , n386029 , n385803 );
nand ( n386031 , n386030 , RI15b43f20_183);
nor ( n386032 , n386031 , n385818 );
nand ( n386033 , n386032 , RI15b44010_185);
not ( n386034 , n386033 );
nand ( n386035 , n386034 , n385841 );
not ( n386036 , n386035 );
nand ( n386037 , n386036 , RI15b443d0_193);
not ( n386038 , n386037 );
buf ( n386039 , n386038 );
buf ( n386040 , n386039 );
nand ( n386041 , n386040 , n385953 );
not ( n386042 , n386039 );
buf ( n386043 , n386042 );
nand ( n386044 , n386043 , RI15b44790_201);
and ( n386045 , n386041 , n386044 , n385957 );
not ( n386046 , n386045 );
nand ( n386047 , n386039 , n385929 );
nand ( n386048 , n386042 , RI15b446a0_199);
and ( n386049 , n386047 , n386048 , n385933 );
not ( n386050 , n386049 );
not ( n386051 , n386029 );
not ( n386052 , RI15b43ea8_182);
and ( n386053 , n386051 , n386052 );
and ( n386054 , n386029 , RI15b43ea8_182);
nor ( n386055 , n386053 , n386054 );
not ( n386056 , n386055 );
not ( n386057 , n386028 );
and ( n386058 , n386057 , n385234 );
not ( n386059 , n386057 );
and ( n386060 , n386059 , RI15b43e30_181);
nor ( n386061 , n386058 , n386060 );
not ( n386062 , n386061 );
nand ( n386063 , n385363 , n386062 );
not ( n386064 , n386063 );
not ( n386065 , n385492 );
not ( n386066 , n386022 );
nand ( n386067 , n386066 , RI15b43c50_177);
or ( n386068 , n386067 , n385228 );
not ( n386069 , n385229 );
nand ( n386070 , n386068 , n386069 );
and ( n386071 , n386070 , n385231 );
not ( n386072 , n386026 );
and ( n386073 , n386072 , RI15b43d40_179);
nor ( n386074 , n386071 , n386073 );
nand ( n386075 , n386065 , n386074 );
not ( n386076 , n385426 );
and ( n386077 , n386027 , RI15b43db8_180);
not ( n386078 , n386027 );
and ( n386079 , n386078 , n385430 );
nor ( n386080 , n386077 , n386079 );
nand ( n386081 , n386076 , n386080 );
and ( n386082 , n386075 , n386081 );
not ( n386083 , n386082 );
and ( n386084 , n386025 , RI15b43cc8_178);
and ( n386085 , n386067 , n385227 );
nor ( n386086 , n386085 , RI15b43cc8_178);
nor ( n386087 , n386084 , n386086 );
nand ( n386088 , n385544 , n386087 );
not ( n386089 , n386088 );
not ( n386090 , n386024 );
and ( n386091 , n386090 , n385554 );
not ( n386092 , n386090 );
and ( n386093 , n386092 , RI15b43c50_177);
nor ( n386094 , n386091 , n386093 );
xor ( n386095 , n386094 , n385591 );
and ( n386096 , n386022 , RI15b43bd8_176);
not ( n386097 , n386022 );
and ( n386098 , n386097 , n386023 );
nor ( n386099 , n386096 , n386098 );
not ( n386100 , n386099 );
nand ( n386101 , n385643 , n386100 );
not ( n386102 , n386101 );
not ( n386103 , n385738 );
nor ( n386104 , n386103 , RI15b43ae8_174);
not ( n386105 , n386104 );
nand ( n386106 , n385695 , n385545 );
not ( n386107 , n386106 );
or ( n386108 , n386105 , n386107 );
nor ( n386109 , n385545 , RI15b43ae8_174);
and ( n386110 , n385545 , RI15b43ae8_174);
or ( n386111 , n386109 , n386110 );
nand ( n386112 , n385696 , n386111 );
nand ( n386113 , n386108 , n386112 );
not ( n386114 , n386113 );
or ( n386115 , n386102 , n386114 );
nand ( n386116 , n385750 , n386099 );
nand ( n386117 , n386115 , n386116 );
and ( n386118 , n386095 , n386117 );
and ( n386119 , n386094 , n385591 );
or ( n386120 , n386118 , n386119 );
not ( n386121 , n386120 );
or ( n386122 , n386089 , n386121 );
not ( n386123 , n386087 );
nand ( n386124 , n386123 , n385543 );
nand ( n386125 , n386122 , n386124 );
not ( n386126 , n386125 );
or ( n386127 , n386083 , n386126 );
not ( n386128 , n386074 );
and ( n386129 , n385492 , n386128 );
and ( n386130 , n386129 , n386081 );
not ( n386131 , n386080 );
and ( n386132 , n385427 , n386131 );
nor ( n386133 , n386130 , n386132 );
nand ( n386134 , n386127 , n386133 );
not ( n386135 , n386134 );
or ( n386136 , n386064 , n386135 );
not ( n386137 , n385363 );
nand ( n386138 , n386137 , n386061 );
nand ( n386139 , n386136 , n386138 );
nand ( n386140 , n386056 , n386139 );
not ( n386141 , n386030 );
not ( n386142 , n386141 );
not ( n386143 , RI15b43f20_183);
and ( n386144 , n386142 , n386143 );
and ( n386145 , n386141 , RI15b43f20_183);
nor ( n386146 , n386144 , n386145 );
nor ( n386147 , n386140 , n386146 );
buf ( n386148 , n386034 );
not ( n386149 , n386148 );
and ( n386150 , RI15b44088_186 , n386149 );
not ( n386151 , RI15b44088_186);
and ( n386152 , n386151 , n386148 );
nor ( n386153 , n386150 , n386152 );
not ( n386154 , n386032 );
and ( n386155 , n386154 , RI15b44010_185);
not ( n386156 , n386154 );
and ( n386157 , n386156 , n385240 );
nor ( n386158 , n386155 , n386157 );
and ( n386159 , n386031 , RI15b43f98_184);
not ( n386160 , n386031 );
and ( n386161 , n386160 , n385818 );
nor ( n386162 , n386159 , n386161 );
nor ( n386163 , n386153 , n386158 , n386162 );
or ( n386164 , n386148 , n385251 );
not ( n386165 , n385773 );
nand ( n386166 , n386148 , n386165 );
nand ( n386167 , n386164 , n386166 , n385778 );
not ( n386168 , n386149 );
or ( n386169 , n386168 , n385783 );
buf ( n386170 , n386148 );
nand ( n386171 , n386170 , n385785 );
nand ( n386172 , n386169 , n386171 , n385788 );
and ( n386173 , n386163 , n386167 , n386172 );
and ( n386174 , n386147 , n386173 );
not ( n386175 , n386037 );
and ( n386176 , n385863 , n386175 );
not ( n386177 , n385863 );
and ( n386178 , n386177 , n386037 );
or ( n386179 , n386176 , n386178 );
not ( n386180 , n386170 );
and ( n386181 , n386180 , RI15b44358_192);
not ( n386182 , n385896 );
not ( n386183 , n386034 );
or ( n386184 , n386182 , n386183 );
nand ( n386185 , n386184 , n385900 );
nor ( n386186 , n386181 , n386185 );
not ( n386187 , n386148 );
not ( n386188 , n385880 );
and ( n386189 , n386187 , n386188 );
not ( n386190 , n385884 );
not ( n386191 , n386034 );
or ( n386192 , n386190 , n386191 );
nand ( n386193 , n386192 , n385889 );
nor ( n386194 , n386189 , n386193 );
and ( n386195 , n386035 , RI15b443d0_193);
not ( n386196 , n386035 );
and ( n386197 , n386196 , n385843 );
nor ( n386198 , n386195 , n386197 );
nor ( n386199 , n386186 , n386194 , n386198 );
or ( n386200 , n386148 , n385837 );
nand ( n386201 , n386148 , n385254 );
nand ( n386202 , n386200 , n386201 , n385256 );
not ( n386203 , RI15b441f0_189);
not ( n386204 , n386149 );
or ( n386205 , n386203 , n386204 );
not ( n386206 , n385829 );
and ( n386207 , n386148 , n386206 );
not ( n386208 , n385832 );
nor ( n386209 , n386207 , n386208 );
nand ( n386210 , n386205 , n386209 );
and ( n386211 , n386179 , n386199 , n386202 , n386210 );
nand ( n386212 , n386037 , RI15b445b0_197);
not ( n386213 , n386037 );
nand ( n386214 , n386213 , n385852 );
nand ( n386215 , n386212 , n386214 , n385856 );
or ( n386216 , n386038 , n385849 );
not ( n386217 , n386037 );
nand ( n386218 , n386217 , n385909 );
nand ( n386219 , n386216 , n386218 , n385911 );
nand ( n386220 , n386217 , n385864 );
nand ( n386221 , n386037 , RI15b444c0_195);
nand ( n386222 , n386220 , n386221 , n385868 );
and ( n386223 , n386211 , n386215 , n386219 , n386222 );
nand ( n386224 , n386174 , n386223 );
nand ( n386225 , n386039 , n385917 );
not ( n386226 , n386039 );
nand ( n386227 , n386226 , RI15b44628_198);
and ( n386228 , n386225 , n386227 , n385921 );
nor ( n386229 , n386224 , n386228 );
nand ( n386230 , n386050 , n386229 );
not ( n386231 , n386043 );
nand ( n386232 , n386231 , n385941 );
nand ( n386233 , n386043 , RI15b44718_200);
and ( n386234 , n386232 , n386233 , n385945 );
nor ( n386235 , n386230 , n386234 );
nand ( n386236 , n386046 , n386235 );
nand ( n386237 , n386040 , n385964 );
not ( n386238 , n386040 );
nand ( n386239 , n386238 , RI15b44808_202);
and ( n386240 , n386237 , n386239 , n385968 );
nor ( n386241 , n386236 , n386240 );
not ( n386242 , n386241 );
not ( n386243 , n386040 );
not ( n386244 , n386243 );
or ( n386245 , n386244 , n385979 );
and ( n386246 , n386244 , n385977 );
nor ( n386247 , n386246 , n385980 );
nand ( n386248 , n386245 , n386247 );
not ( n386249 , n386248 );
not ( n386250 , n386249 );
and ( n386251 , n386242 , n386250 );
and ( n386252 , n386241 , n386249 );
nor ( n386253 , n386251 , n386252 );
buf ( n386254 , n20588 );
not ( n386255 , n386254 );
not ( n386256 , n381046 );
nor ( n386257 , n386255 , n386256 , n20332 );
and ( n386258 , n386257 , n20501 );
not ( n386259 , n386258 );
buf ( n386260 , n386259 );
buf ( n386261 , n386260 );
not ( n386262 , n386261 );
not ( n386263 , n386262 );
not ( n386264 , n386263 );
not ( n386265 , n386264 );
or ( n386266 , n386253 , n386265 );
not ( n386267 , RI15b44880_203);
nand ( n386268 , n385241 , RI15b43ae8_174);
not ( n386269 , n386268 );
nand ( n386270 , n386269 , n385841 );
not ( n386271 , n386270 );
nand ( n386272 , n386271 , RI15b443d0_193);
not ( n386273 , n386272 );
not ( n386274 , n386273 );
buf ( n386275 , n386274 );
buf ( n386276 , n386275 );
not ( n386277 , n386276 );
buf ( n386278 , n386277 );
not ( n386279 , n386278 );
not ( n386280 , n386279 );
or ( n386281 , n386267 , n386280 );
and ( n386282 , n386278 , n385977 );
nor ( n386283 , n386282 , n385980 );
nand ( n386284 , n386281 , n386283 );
not ( n386285 , n386284 );
not ( n386286 , n386276 );
not ( n386287 , RI15b44790_201);
or ( n386288 , n386286 , n386287 );
nand ( n386289 , n386286 , n385953 );
nand ( n386290 , n386288 , n386289 , n385957 );
not ( n386291 , n386290 );
not ( n386292 , RI15b44628_198);
not ( n386293 , n386275 );
or ( n386294 , n386292 , n386293 );
buf ( n386295 , n386274 );
not ( n386296 , n386295 );
and ( n386297 , n386296 , n385917 );
not ( n386298 , n385921 );
nor ( n386299 , n386297 , n386298 );
nand ( n386300 , n386294 , n386299 );
not ( n386301 , n386300 );
buf ( n386302 , n385738 );
not ( n386303 , n385695 );
and ( n386304 , n386302 , n386303 );
nor ( n386305 , n386304 , n386109 );
nand ( n386306 , n385746 , n386305 );
nand ( n386307 , n385643 , n386099 );
nand ( n386308 , n386306 , n386307 );
nor ( n386309 , n386022 , n385227 );
and ( n386310 , n386309 , n385228 );
not ( n386311 , n386309 );
and ( n386312 , n386311 , RI15b43cc8_178);
nor ( n386313 , n386310 , n386312 );
nand ( n386314 , n385541 , n386313 );
nand ( n386315 , n385229 , n386066 );
and ( n386316 , n386315 , RI15b43d40_179);
not ( n386317 , n386315 );
and ( n386318 , n386317 , n385231 );
nor ( n386319 , n386316 , n386318 );
nand ( n386320 , n385490 , n386319 );
or ( n386321 , n386315 , n385231 );
and ( n386322 , n386321 , RI15b43db8_180);
not ( n386323 , n386321 );
and ( n386324 , n386323 , n385430 );
nor ( n386325 , n386322 , n386324 );
nand ( n386326 , n385424 , n386325 );
nand ( n386327 , n386314 , n386320 , n386326 );
not ( n386328 , n386327 );
nand ( n386329 , n386066 , RI15b43bd8_176);
and ( n386330 , n386329 , RI15b43c50_177);
not ( n386331 , n386329 );
and ( n386332 , n386331 , n385554 );
nor ( n386333 , n386330 , n386332 );
nand ( n386334 , n385590 , n386333 );
buf ( n386335 , n386334 );
nand ( n386336 , n386328 , n386335 );
or ( n386337 , n386308 , n386336 );
not ( n386338 , n386327 );
nor ( n386339 , n385643 , n386099 );
nand ( n386340 , n386334 , n386339 );
not ( n386341 , n386340 );
and ( n386342 , n386338 , n386341 );
not ( n386343 , n386326 );
not ( n386344 , n386319 );
nand ( n386345 , n385491 , n386344 );
or ( n386346 , n386343 , n386345 );
not ( n386347 , n386325 );
nand ( n386348 , n385425 , n386347 );
nand ( n386349 , n386346 , n386348 );
nor ( n386350 , n386342 , n386349 );
not ( n386351 , n386327 );
or ( n386352 , n385590 , n386333 );
not ( n386353 , n386352 );
and ( n386354 , n386351 , n386353 );
not ( n386355 , n386313 );
nand ( n386356 , n385542 , n386355 );
nor ( n386357 , n386356 , n386343 );
buf ( n386358 , n386320 );
and ( n386359 , n386357 , n386358 );
nor ( n386360 , n386354 , n386359 );
nand ( n386361 , n386337 , n386350 , n386360 );
buf ( n386362 , n386361 );
not ( n386363 , n386321 );
nand ( n386364 , n386363 , RI15b43db8_180);
and ( n386365 , n386364 , RI15b43e30_181);
not ( n386366 , n386364 );
and ( n386367 , n386366 , n385234 );
nor ( n386368 , n386365 , n386367 );
nand ( n386369 , n385362 , n386368 );
nand ( n386370 , n386362 , n386369 );
not ( n386371 , n386268 );
not ( n386372 , n386371 );
and ( n386373 , n386372 , RI15b44178_188);
or ( n386374 , n386268 , n385773 );
nand ( n386375 , n386374 , n385778 );
nor ( n386376 , n386373 , n386375 );
not ( n386377 , n386371 );
and ( n386378 , n386377 , RI15b44268_190);
not ( n386379 , n386269 );
not ( n386380 , n385254 );
or ( n386381 , n386379 , n386380 );
nand ( n386382 , n386381 , n385256 );
nor ( n386383 , n386378 , n386382 );
not ( n386384 , n386371 );
and ( n386385 , n386384 , RI15b44100_187);
or ( n386386 , n386379 , n385784 );
nand ( n386387 , n386386 , n385788 );
nor ( n386388 , n386385 , n386387 );
and ( n386389 , n386384 , RI15b44358_192);
not ( n386390 , n385896 );
or ( n386391 , n386379 , n386390 );
nand ( n386392 , n386391 , n385900 );
nor ( n386393 , n386389 , n386392 );
nand ( n386394 , n386376 , n386383 , n386388 , n386393 );
and ( n386395 , n386372 , RI15b441f0_189);
or ( n386396 , n386379 , n385829 );
nand ( n386397 , n386396 , n385832 );
nor ( n386398 , n386395 , n386397 );
not ( n386399 , n386371 );
not ( n386400 , n385880 );
and ( n386401 , n386399 , n386400 );
or ( n386402 , n386268 , n385883 );
nand ( n386403 , n386402 , n385889 );
nor ( n386404 , n386401 , n386403 );
not ( n386405 , n386268 );
not ( n386406 , RI15b44088_186);
and ( n386407 , n386405 , n386406 );
and ( n386408 , n386377 , RI15b44088_186);
nor ( n386409 , n386407 , n386408 );
nand ( n386410 , n385810 , RI15b43ae8_174);
and ( n386411 , n386410 , RI15b44010_185);
not ( n386412 , n386410 );
and ( n386413 , n386412 , n385240 );
nor ( n386414 , n386411 , n386413 );
nand ( n386415 , n385816 , RI15b43ae8_174);
and ( n386416 , n386415 , RI15b43f98_184);
not ( n386417 , n386415 );
and ( n386418 , n386417 , n385818 );
nor ( n386419 , n386416 , n386418 );
not ( n386420 , n385236 );
nand ( n386421 , n386420 , RI15b43ae8_174);
and ( n386422 , n386421 , RI15b43f20_183);
not ( n386423 , n386421 );
and ( n386424 , n386423 , n385237 );
nor ( n386425 , n386422 , n386424 );
not ( n386426 , n385802 );
nand ( n386427 , n386426 , RI15b43ae8_174);
and ( n386428 , n386427 , RI15b43ea8_182);
not ( n386429 , n386427 );
and ( n386430 , n386429 , n385803 );
nor ( n386431 , n386428 , n386430 );
and ( n386432 , n386419 , n386425 , n386431 );
or ( n386433 , n385361 , n386368 );
and ( n386434 , n386414 , n386432 , n386433 );
nand ( n386435 , n386398 , n386404 , n386409 , n386434 );
nor ( n386436 , n386394 , n386435 );
not ( n386437 , n386273 );
not ( n386438 , n385863 );
and ( n386439 , n386437 , n386438 );
and ( n386440 , n386273 , n385863 );
nor ( n386441 , n386439 , n386440 );
buf ( n386442 , n386270 );
and ( n386443 , n386442 , RI15b443d0_193);
not ( n386444 , n386442 );
and ( n386445 , n386444 , n385843 );
nor ( n386446 , n386443 , n386445 );
nand ( n386447 , n386370 , n386436 , n386441 , n386446 );
not ( n386448 , RI15b444c0_195);
not ( n386449 , n386274 );
or ( n386450 , n386448 , n386449 );
not ( n386451 , n385864 );
not ( n386452 , n386273 );
or ( n386453 , n386451 , n386452 );
nand ( n386454 , n386453 , n385868 );
not ( n386455 , n386454 );
nand ( n386456 , n386450 , n386455 );
nor ( n386457 , n386447 , n386456 );
not ( n386458 , n385909 );
not ( n386459 , n386274 );
not ( n386460 , n386459 );
or ( n386461 , n386458 , n386460 );
nand ( n386462 , n386461 , n385911 );
not ( n386463 , n386274 );
nor ( n386464 , n386463 , n385849 );
nor ( n386465 , n386462 , n386464 );
nand ( n386466 , n386457 , n386465 );
not ( n386467 , RI15b445b0_197);
not ( n386468 , n386295 );
or ( n386469 , n386467 , n386468 );
and ( n386470 , n386463 , n385852 );
not ( n386471 , n385856 );
nor ( n386472 , n386470 , n386471 );
nand ( n386473 , n386469 , n386472 );
nor ( n386474 , n386466 , n386473 );
nand ( n386475 , n386301 , n386474 );
nand ( n386476 , n386275 , RI15b446a0_199);
nand ( n386477 , n386296 , n385929 );
nand ( n386478 , n386476 , n386477 , n385933 );
nor ( n386479 , n386475 , n386478 );
and ( n386480 , n386276 , RI15b44718_200);
not ( n386481 , n385941 );
not ( n386482 , n386275 );
not ( n386483 , n386482 );
or ( n386484 , n386481 , n386483 );
nand ( n386485 , n386484 , n385945 );
nor ( n386486 , n386480 , n386485 );
and ( n386487 , n386479 , n386486 );
nand ( n386488 , n386291 , n386487 );
or ( n386489 , n386286 , n385974 );
nand ( n386490 , n386277 , n385964 );
nand ( n386491 , n386489 , n386490 , n385968 );
nor ( n386492 , n386488 , n386491 );
not ( n386493 , n386492 );
not ( n386494 , n386493 );
or ( n386495 , n386285 , n386494 );
not ( n386496 , n386284 );
nand ( n386497 , n386496 , n386492 );
nand ( n386498 , n386495 , n386497 );
nand ( n386499 , n386011 , n385364 );
not ( n386500 , n386499 );
and ( n386501 , n386498 , n386500 );
not ( n386502 , n22398 );
nor ( n386503 , n386502 , n380886 );
nor ( n386504 , n386501 , n386503 );
nand ( n386505 , n386266 , n386504 );
nor ( n386506 , n386021 , n386505 );
not ( n386507 , n381030 );
not ( n386508 , n20608 );
or ( n386509 , n386507 , n386508 );
not ( n386510 , n381053 );
nor ( n386511 , n381074 , n386510 );
nand ( n386512 , n386509 , n386511 );
buf ( n386513 , n386512 );
buf ( n386514 , n386513 );
not ( n386515 , n386514 );
buf ( n386516 , n386515 );
not ( n386517 , n386516 );
and ( n386518 , n386517 , n386284 );
not ( n386519 , n20501 );
nand ( n386520 , n20589 , n386010 );
nand ( n386521 , n386254 , n381060 , n20507 );
nand ( n386522 , n386520 , n386521 );
not ( n386523 , n386522 );
or ( n386524 , n386519 , n386523 );
nand ( n386525 , n386524 , n20621 );
not ( n386526 , n20561 );
and ( n386527 , n20585 , n386526 );
nand ( n386528 , n386527 , n20501 );
nand ( n386529 , n381039 , n381034 );
not ( n386530 , n381046 );
and ( n386531 , n386529 , n386530 );
not ( n386532 , n20628 );
or ( n386533 , n22234 , n386532 );
or ( n386534 , n386533 , n385210 );
nor ( n386535 , n386531 , n386534 );
and ( n386536 , n20578 , n20501 );
or ( n386537 , n379817 , n386536 );
nand ( n386538 , n386537 , n379828 );
nand ( n386539 , n386528 , n386535 , n386538 );
or ( n386540 , n386525 , n386539 );
not ( n386541 , n386540 );
or ( n386542 , n386541 , n385979 );
and ( n386543 , n20585 , n20561 );
not ( n386544 , n20595 );
nor ( n386545 , n386543 , n386544 );
nor ( n386546 , n386545 , n20519 );
nand ( n386547 , n386536 , n379818 );
nand ( n386548 , n379819 , n386547 );
or ( n386549 , n386546 , n386548 );
not ( n386550 , n386549 );
or ( n386551 , n385983 , n386550 );
not ( n386552 , n381046 );
not ( n386553 , n386552 );
and ( n386554 , n381035 , n386553 );
not ( n386555 , n381062 );
or ( n386556 , n386554 , n386555 );
not ( n386557 , n386556 );
or ( n386558 , n386557 , n386249 );
nand ( n386559 , n386542 , n386551 , n386558 );
nor ( n386560 , n386518 , n386559 );
nand ( n386561 , n386506 , n386560 );
buf ( n386562 , n386561 );
buf ( n386563 , RI15b3ea48_2);
buf ( n386564 , n386563 );
buf ( n386565 , n381081 );
buf ( n386566 , n22343 );
buf ( n386567 , n380906 );
buf ( n386568 , n22406 );
buf ( n386569 , n380646 );
buf ( n386570 , n383179 );
or ( n386571 , n386569 , n386570 );
not ( n386572 , n380636 );
buf ( n386573 , n380548 );
nor ( n386574 , n386572 , n386573 );
not ( n386575 , n386574 );
nand ( n386576 , n386575 , n386569 , n386570 );
nand ( n386577 , n386571 , n386576 );
not ( n386578 , n386577 );
not ( n386579 , n380698 );
or ( n386580 , n386578 , n386579 );
not ( n386581 , n386570 );
nand ( n386582 , n386581 , n19645 );
not ( n386583 , n386582 );
not ( n386584 , n380685 );
or ( n386585 , n386583 , n386584 );
nand ( n386586 , n386585 , n386574 );
nand ( n386587 , n386580 , n386586 );
not ( n386588 , n386587 );
not ( n386589 , n380727 );
and ( n386590 , n386589 , n381493 );
not ( n386591 , n386590 );
or ( n386592 , n386588 , n386591 );
not ( n386593 , n382917 );
nand ( n386594 , n380512 , n381522 );
nor ( n386595 , n386593 , n386594 );
nand ( n386596 , n382918 , n381522 );
or ( n386597 , n382917 , n386596 );
or ( n386598 , n382926 , n380468 );
nand ( n386599 , n386597 , n386598 );
or ( n386600 , n386595 , n386599 );
not ( n386601 , n382932 );
or ( n386602 , n386601 , n380758 );
not ( n386603 , n386602 );
and ( n386604 , n386600 , n386603 );
and ( n386605 , n386602 , n386591 , n381531 );
nor ( n386606 , n386605 , n19630 );
nor ( n386607 , n382940 , n380728 );
or ( n386608 , n386606 , n386607 );
nand ( n386609 , n386608 , n19595 );
or ( n386610 , n382945 , n381541 );
nand ( n386611 , n386609 , n386610 );
and ( n386612 , n386611 , n380775 );
not ( n386613 , RI15b59eb0_933);
or ( n386614 , n386612 , n386613 );
not ( n386615 , n380308 );
not ( n386616 , n386615 );
buf ( n386617 , n386616 );
buf ( n386618 , n386617 );
not ( n386619 , n386607 );
not ( n386620 , n386610 );
not ( n386621 , n386620 );
and ( n386622 , n386619 , n386621 );
nor ( n386623 , n386622 , n386606 );
not ( n386624 , n386623 );
or ( n386625 , n386618 , n386624 );
buf ( n386626 , n19193 );
or ( n386627 , n386626 , n380788 );
or ( n386628 , n386610 , n386627 );
nand ( n386629 , n386614 , n386625 , n386628 );
nor ( n386630 , n386604 , n386629 );
nand ( n386631 , n386592 , n386630 );
buf ( n386632 , n386631 );
buf ( n386633 , n19655 );
or ( n386634 , n381396 , n381238 );
not ( n386635 , n381402 );
nand ( n386636 , n386634 , n386635 );
not ( n386637 , n382679 );
and ( n386638 , n386637 , RI15b54ff0_765);
and ( n386639 , n381636 , RI15b4ec18_552);
and ( n386640 , n381639 , RI15b4e858_544);
nor ( n386641 , n386639 , n386640 );
and ( n386642 , n381643 , RI15b4efd8_560);
not ( n386643 , n381645 );
and ( n386644 , n382837 , RI15b4dd18_520);
and ( n386645 , n382852 , RI15b4fed8_592);
nor ( n386646 , n386644 , n386645 );
and ( n386647 , n381661 , RI15b4fb18_584);
and ( n386648 , n381663 , RI15b4f398_568);
nor ( n386649 , n386647 , n386648 );
and ( n386650 , n381667 , RI15b4d598_504);
and ( n386651 , n381669 , RI15b4d958_512);
nor ( n386652 , n386650 , n386651 );
and ( n386653 , n381672 , RI15b4e0d8_528);
and ( n386654 , n381674 , RI15b4f758_576);
nor ( n386655 , n386653 , n386654 );
nand ( n386656 , n386646 , n386649 , n386652 , n386655 );
and ( n386657 , n386643 , n386656 );
and ( n386658 , n381680 , RI15b4ca58_480);
nor ( n386659 , n386642 , n386657 , n386658 );
and ( n386660 , n381684 , RI15b4c698_472);
and ( n386661 , n381686 , RI15b4e498_536);
nor ( n386662 , n386660 , n386661 );
and ( n386663 , n381689 , RI15b4ce18_488);
and ( n386664 , n381691 , RI15b4d1d8_496);
nor ( n386665 , n386663 , n386664 );
nand ( n386666 , n386641 , n386659 , n386662 , n386665 );
buf ( n386667 , n379996 );
not ( n386668 , n386667 );
not ( n386669 , n386668 );
not ( n386670 , n386669 );
not ( n386671 , n386670 );
and ( n386672 , n386666 , n386671 );
or ( n386673 , n382691 , n381118 );
not ( n386674 , n382626 );
not ( n386675 , n382650 );
not ( n386676 , RI15b54ff0_765);
and ( n386677 , n386675 , n386676 );
and ( n386678 , n382650 , RI15b54ff0_765);
nor ( n386679 , n386677 , n386678 );
or ( n386680 , n386674 , n386679 );
nand ( n386681 , n386673 , n386680 );
nor ( n386682 , n386638 , n386672 , n386681 );
nand ( n386683 , n386636 , n386682 );
buf ( n386684 , n386683 );
buf ( n386685 , n383498 );
not ( n386686 , n384078 );
nor ( n386687 , n386686 , n384102 );
not ( n386688 , n386687 );
nand ( n386689 , n383798 , n383711 );
not ( n386690 , n383705 );
nor ( n386691 , n386689 , n386690 );
nand ( n386692 , n386691 , n384089 );
not ( n386693 , n386692 );
or ( n386694 , n386688 , n386693 );
buf ( n386695 , n383809 );
not ( n386696 , n386695 );
not ( n386697 , n386689 );
not ( n386698 , n384089 );
nor ( n386699 , n386698 , n383807 );
nand ( n386700 , n386697 , n386699 );
not ( n386701 , n386700 );
or ( n386702 , n386696 , n386701 );
nand ( n386703 , n386702 , n384102 );
nand ( n386704 , n386694 , n386703 );
not ( n386705 , n386704 );
nand ( n386706 , n384054 , n383866 );
or ( n386707 , n386705 , n386706 );
not ( n386708 , n384131 );
not ( n386709 , n384136 );
and ( n386710 , n386708 , n386709 );
not ( n386711 , n386708 );
and ( n386712 , n386711 , n384136 );
nor ( n386713 , n386710 , n386712 );
nand ( n386714 , n386713 , n384157 );
nand ( n386715 , n384148 , n384134 );
nand ( n386716 , n386714 , n386715 );
nand ( n386717 , n384167 , n384056 );
not ( n386718 , n386717 );
and ( n386719 , n386716 , n386718 );
and ( n386720 , n386717 , n386706 , n385009 );
nor ( n386721 , n386720 , n21764 );
nor ( n386722 , n384173 , n383832 );
or ( n386723 , n386721 , n386722 );
nand ( n386724 , n386723 , n18154 );
or ( n386725 , n384179 , n383886 );
nand ( n386726 , n386724 , n386725 );
and ( n386727 , n386726 , n383901 );
or ( n386728 , n386727 , n17856 );
buf ( n386729 , n381353 );
buf ( n386730 , n386729 );
buf ( n386731 , n386730 );
not ( n386732 , n386731 );
not ( n386733 , n386725 );
nor ( n386734 , n386722 , n386733 );
or ( n386735 , n386721 , n386734 );
or ( n386736 , n386732 , n386735 );
buf ( n386737 , n17878 );
or ( n386738 , n386737 , n383916 );
or ( n386739 , n386725 , n386738 );
nand ( n386740 , n386728 , n386736 , n386739 );
nor ( n386741 , n386719 , n386740 );
nand ( n386742 , n386707 , n386741 );
buf ( n386743 , n386742 );
buf ( n386744 , RI15b5da38_1060);
or ( n386745 , n384021 , n384031 );
and ( n386746 , n383926 , n19495 );
not ( n386747 , n386746 );
or ( n386748 , n18496 , n386747 );
and ( n386749 , n384030 , RI15b61e30_1205);
not ( n386750 , n384030 );
and ( n386751 , n386750 , n384031 );
nor ( n386752 , n386749 , n386751 );
or ( n386753 , n386752 , n384024 );
nand ( n386754 , n386745 , n386748 , n386753 );
buf ( n386755 , n386754 );
buf ( n386756 , n384199 );
buf ( n386757 , n384199 );
buf ( n386758 , n379847 );
buf ( n386759 , n382071 );
buf ( n386760 , RI15b3e9d0_1);
buf ( n386761 , n386760 );
buf ( n386762 , RI15b3e9d0_1);
buf ( n386763 , n386762 );
not ( n386764 , n19628 );
buf ( n386765 , n383456 );
nand ( n386766 , n386765 , n383424 );
not ( n386767 , RI15b63780_1259);
and ( n386768 , n386766 , n386767 );
not ( n386769 , n386766 );
and ( n386770 , n386769 , RI15b63780_1259);
nor ( n386771 , n386768 , n386770 );
not ( n386772 , n386771 );
nand ( n386773 , n383456 , n383421 );
not ( n386774 , RI15b63690_1257);
and ( n386775 , n386773 , n386774 );
not ( n386776 , n386773 );
and ( n386777 , n386776 , RI15b63690_1257);
nor ( n386778 , n386775 , n386777 );
not ( n386779 , n386778 );
nand ( n386780 , n383455 , RI15b63528_1254);
not ( n386781 , RI15b635a0_1255);
and ( n386782 , n386780 , n386781 );
not ( n386783 , n386780 );
and ( n386784 , n386783 , RI15b635a0_1255);
nor ( n386785 , n386782 , n386784 );
not ( n386786 , n386785 );
nand ( n386787 , RI15b62bc8_1234 , RI15b62c40_1235);
not ( n386788 , n386787 );
not ( n386789 , RI15b62cb8_1236);
and ( n386790 , n386788 , n386789 );
and ( n386791 , n386787 , RI15b62cb8_1236);
nor ( n386792 , n386790 , n386791 );
nor ( n386793 , n383466 , RI15b62b50_1233);
nand ( n386794 , n386792 , n386793 );
not ( n386795 , RI15b62d30_1237);
not ( n386796 , n386795 );
buf ( n386797 , n19612 );
nor ( n386798 , n386797 , n19620 );
not ( n386799 , n386798 );
or ( n386800 , n386796 , n386799 );
not ( n386801 , RI15b62d30_1237);
or ( n386802 , n386798 , n386801 );
nand ( n386803 , n386800 , n386802 );
nor ( n386804 , n386794 , n386803 );
buf ( n386805 , n19614 );
nand ( n386806 , n386805 , RI15b62bc8_1234);
and ( n386807 , n386806 , RI15b62da8_1238);
not ( n386808 , n386806 );
not ( n386809 , RI15b62da8_1238);
and ( n386810 , n386808 , n386809 );
nor ( n386811 , n386807 , n386810 );
nand ( n386812 , n386804 , n386811 );
nor ( n386813 , n386812 , n382612 );
nand ( n386814 , n386813 , n22774 );
nor ( n386815 , n386814 , n19625 );
nand ( n386816 , n386815 , n380852 );
not ( n386817 , RI15b63000_1243);
not ( n386818 , n386817 );
nand ( n386819 , n383444 , RI15b62bc8_1234);
not ( n386820 , n386819 );
not ( n386821 , n386820 );
or ( n386822 , n386818 , n386821 );
or ( n386823 , n386820 , n386817 );
nand ( n386824 , n386822 , n386823 );
nor ( n386825 , n386816 , n386824 );
not ( n386826 , n383445 );
nand ( n386827 , n386826 , RI15b62bc8_1234);
and ( n386828 , n386827 , RI15b63078_1244);
not ( n386829 , n386827 );
and ( n386830 , n386829 , n383446 );
nor ( n386831 , n386828 , n386830 );
nand ( n386832 , n386825 , n386831 );
not ( n386833 , RI15b630f0_1245);
not ( n386834 , n386833 );
not ( n386835 , n383448 );
or ( n386836 , n386834 , n386835 );
or ( n386837 , n383448 , n386833 );
nand ( n386838 , n386836 , n386837 );
nor ( n386839 , n386832 , n386838 );
and ( n386840 , n383449 , RI15b63168_1246);
not ( n386841 , n383449 );
not ( n386842 , RI15b63168_1246);
and ( n386843 , n386841 , n386842 );
nor ( n386844 , n386840 , n386843 );
and ( n386845 , n386839 , n386844 );
not ( n386846 , n383449 );
nand ( n386847 , n386846 , RI15b63168_1246);
and ( n386848 , n386847 , RI15b631e0_1247);
not ( n386849 , n386847 );
not ( n386850 , RI15b631e0_1247);
and ( n386851 , n386849 , n386850 );
nor ( n386852 , n386848 , n386851 );
nand ( n386853 , n386845 , n386852 );
not ( n386854 , RI15b63258_1248);
not ( n386855 , n386854 );
nor ( n386856 , n383450 , n383434 );
not ( n386857 , n386856 );
or ( n386858 , n386855 , n386857 );
not ( n386859 , n383450 );
and ( n386860 , n386859 , n383435 );
or ( n386861 , n386860 , n386854 );
nand ( n386862 , n386858 , n386861 );
nor ( n386863 , n386853 , n386862 );
not ( n386864 , n383450 );
nand ( n386865 , n386864 , n383436 );
and ( n386866 , n386865 , RI15b632d0_1249);
not ( n386867 , n386865 );
not ( n386868 , RI15b632d0_1249);
and ( n386869 , n386867 , n386868 );
nor ( n386870 , n386866 , n386869 );
and ( n386871 , n386863 , n386870 );
not ( n386872 , n383451 );
nand ( n386873 , n386872 , n383437 );
and ( n386874 , n386873 , RI15b63348_1250);
not ( n386875 , n386873 );
not ( n386876 , RI15b63348_1250);
and ( n386877 , n386875 , n386876 );
nor ( n386878 , n386874 , n386877 );
nand ( n386879 , n386871 , n386878 );
not ( n386880 , n383439 );
nor ( n386881 , n383451 , n383438 );
not ( n386882 , n386881 );
or ( n386883 , n386880 , n386882 );
or ( n386884 , n386881 , n383439 );
nand ( n386885 , n386883 , n386884 );
nor ( n386886 , n386879 , n386885 );
not ( n386887 , n383452 );
nor ( n386888 , n386887 , n383440 );
and ( n386889 , n386888 , n383441 );
not ( n386890 , n386888 );
and ( n386891 , n386890 , RI15b63438_1252);
nor ( n386892 , n386889 , n386891 );
and ( n386893 , n386886 , n386892 );
and ( n386894 , n383453 , RI15b634b0_1253);
not ( n386895 , n383453 );
and ( n386896 , n386895 , n383454 );
nor ( n386897 , n386894 , n386896 );
nand ( n386898 , n386893 , n386897 );
not ( n386899 , n383455 );
and ( n386900 , n386899 , RI15b63528_1254);
not ( n386901 , n386899 );
not ( n386902 , RI15b63528_1254);
and ( n386903 , n386901 , n386902 );
nor ( n386904 , n386900 , n386903 );
not ( n386905 , n386904 );
nor ( n386906 , n386898 , n386905 );
nand ( n386907 , n386786 , n386906 );
nor ( n386908 , n386899 , n383419 );
and ( n386909 , n386908 , RI15b63618_1256);
not ( n386910 , n386908 );
and ( n386911 , n386910 , n383420 );
nor ( n386912 , n386909 , n386911 );
nor ( n386913 , n386907 , n386912 );
nand ( n386914 , n386779 , n386913 );
nor ( n386915 , n386914 , n384650 );
nand ( n386916 , n386772 , n386915 );
not ( n386917 , n386765 );
nor ( n386918 , n386917 , n383425 );
and ( n386919 , n386918 , RI15b637f8_1260);
not ( n386920 , n386918 );
and ( n386921 , n386920 , n383426 );
nor ( n386922 , n386919 , n386921 );
nor ( n386923 , n386916 , n386922 );
buf ( n386924 , n386765 );
nand ( n386925 , n386924 , n383427 );
not ( n386926 , RI15b63870_1261);
and ( n386927 , n386925 , n386926 );
not ( n386928 , n386925 );
and ( n386929 , n386928 , RI15b63870_1261);
nor ( n386930 , n386927 , n386929 );
not ( n386931 , n386930 );
nand ( n386932 , n386923 , n386931 );
not ( n386933 , n386924 );
nor ( n386934 , n386933 , n383428 );
and ( n386935 , n386934 , RI15b638e8_1262);
not ( n386936 , n386934 );
and ( n386937 , n386936 , n383429 );
nor ( n386938 , n386935 , n386937 );
nor ( n386939 , n386932 , n386938 );
not ( n386940 , n386939 );
or ( n386941 , n386764 , n386940 );
buf ( n386942 , n383473 );
not ( n386943 , n386942 );
buf ( n386944 , n386943 );
buf ( n386945 , n386944 );
buf ( n386946 , n386945 );
not ( n386947 , n386946 );
nand ( n386948 , n386941 , n386947 );
not ( n386949 , n383430 );
nand ( n386950 , n386949 , n386924 );
and ( n386951 , n386950 , n383431 );
not ( n386952 , n386950 );
and ( n386953 , n386952 , RI15b63960_1263);
nor ( n386954 , n386951 , n386953 );
nand ( n386955 , n386948 , n386954 );
not ( n386956 , RI15b61d40_1203);
and ( n386957 , n383403 , n386956 );
not ( n386958 , RI15b61db8_1204);
nand ( n386959 , n386957 , n386958 );
nor ( n386960 , n386959 , RI15b61e30_1205);
not ( n386961 , RI15b61ea8_1206);
and ( n386962 , n386960 , n386961 );
not ( n386963 , RI15b61f20_1207);
nand ( n386964 , n386962 , n386963 );
nor ( n386965 , n386964 , RI15b61f98_1208);
not ( n386966 , RI15b62010_1209);
and ( n386967 , n386965 , n386966 );
nand ( n386968 , n386967 , n384038 );
nor ( n386969 , n386968 , RI15b62100_1211);
not ( n386970 , RI15b62178_1212);
and ( n386971 , n386969 , n386970 );
not ( n386972 , RI15b621f0_1213);
nand ( n386973 , n386971 , n386972 );
nor ( n386974 , n386973 , RI15b62268_1214);
not ( n386975 , RI15b622e0_1215);
and ( n386976 , n386974 , n386975 );
not ( n386977 , RI15b62358_1216);
nand ( n386978 , n386976 , n386977 );
nor ( n386979 , n386978 , RI15b623d0_1217);
not ( n386980 , RI15b62448_1218);
nand ( n386981 , n386979 , n386980 );
nor ( n386982 , n386981 , RI15b624c0_1219);
not ( n386983 , RI15b62538_1220);
and ( n386984 , n386982 , n386983 );
not ( n386985 , RI15b625b0_1221);
nand ( n386986 , n386984 , n386985 );
nor ( n386987 , n386986 , RI15b62628_1222);
not ( n386988 , RI15b626a0_1223);
and ( n386989 , n386987 , n386988 );
not ( n386990 , RI15b62718_1224);
nand ( n386991 , n386989 , n386990 );
nor ( n386992 , n386991 , RI15b62790_1225);
not ( n386993 , RI15b62808_1226);
and ( n386994 , n386992 , n386993 );
not ( n386995 , RI15b62880_1227);
nand ( n386996 , n386994 , n386995 );
nor ( n386997 , n386996 , RI15b628f8_1228);
not ( n386998 , RI15b62970_1229);
nand ( n386999 , n386997 , n386998 );
not ( n387000 , n386999 );
not ( n387001 , RI15b629e8_1230);
nand ( n387002 , n387000 , n387001 );
not ( n387003 , n383402 );
buf ( n387004 , n387003 );
not ( n387005 , n387004 );
not ( n387006 , n387005 );
nor ( n387007 , n387002 , n387006 );
or ( n387008 , n387007 , n383409 );
nand ( n387009 , n387008 , RI15b62a60_1231);
not ( n387010 , n386939 );
not ( n387011 , n383464 );
buf ( n387012 , n387011 );
not ( n387013 , n387012 );
nor ( n387014 , n387013 , n386954 );
nand ( n387015 , n387010 , n387014 );
nor ( n387016 , n383482 , RI15b62a60_1231);
and ( n387017 , n387002 , n387016 );
not ( n387018 , n379771 );
not ( n387019 , RI15b63bb8_1268);
nand ( n387020 , RI15b63ac8_1266 , RI15b63b40_1267);
nor ( n387021 , n387019 , n387020 );
and ( n387022 , RI15b63c30_1269 , RI15b63ca8_1270);
nand ( n387023 , n387021 , n387022 );
not ( n387024 , n387023 );
and ( n387025 , n387024 , RI15b63d20_1271);
nand ( n387026 , n387025 , RI15b63d98_1272);
nor ( n387027 , n387026 , n379554 );
nand ( n387028 , n387027 , RI15b63e88_1274);
not ( n387029 , n387028 );
nand ( n387030 , n387029 , RI15b63f00_1275);
nor ( n387031 , n387030 , n379573 );
and ( n387032 , n387031 , RI15b63ff0_1277);
nand ( n387033 , n387032 , RI15b64068_1278);
nor ( n387034 , n387033 , n379612 );
and ( n387035 , n387034 , RI15b64158_1280);
nand ( n387036 , n387035 , RI15b641d0_1281 , RI15b64248_1282);
nor ( n387037 , n387036 , n379436 );
nand ( n30842 , n387037 , RI15b64338_1284);
nand ( n30843 , RI15b643b0_1285 , RI15b64428_1286);
nor ( n30844 , n30842 , n30843 );
nor ( n30845 , n379708 , n379711 );
nand ( n30846 , n30844 , n30845 );
nand ( n30847 , RI15b64590_1289 , RI15b64608_1290);
nor ( n30848 , n30846 , n30847 );
nor ( n30849 , n379720 , n379448 );
nand ( n30850 , n30848 , n30849 );
not ( n30851 , n30850 );
and ( n30852 , n30851 , RI15b64770_1293 , RI15b647e8_1294);
not ( n30853 , n30852 );
or ( n30854 , n387018 , n30853 );
or ( n30855 , n30852 , n379771 );
nand ( n30856 , n30854 , n30855 );
nand ( n30857 , n30856 , n22450 );
nand ( n30858 , n22426 , RI15b64860_1295);
nand ( n30859 , n19599 , RI15b63960_1263);
nand ( n30860 , n30857 , n30858 , n30859 );
nor ( n30861 , n387017 , n30860 );
nand ( n30862 , n386955 , n387009 , n387015 , n30861 );
buf ( n30863 , n30862 );
buf ( n30864 , n386563 );
not ( n30865 , n385807 );
buf ( n30866 , n385770 );
nand ( n30867 , n30866 , n385433 );
nand ( n30868 , n30867 , n385368 );
not ( n30869 , n30868 );
or ( n30870 , n30865 , n30869 );
or ( n30871 , n30868 , n385807 );
nand ( n30872 , n30870 , n30871 );
buf ( n30873 , n386016 );
and ( n30874 , n30872 , n30873 );
not ( n30875 , n386139 );
not ( n30876 , n386055 );
and ( n30877 , n30875 , n30876 );
and ( n30878 , n386139 , n386055 );
nor ( n30879 , n30877 , n30878 );
or ( n30880 , n30879 , n386260 );
not ( n30881 , n386369 );
not ( n30882 , n386361 );
or ( n30883 , n30881 , n30882 );
nand ( n30884 , n30883 , n386433 );
not ( n30885 , n30884 );
not ( n30886 , n30885 );
not ( n30887 , n386431 );
and ( n30888 , n30886 , n30887 );
not ( n30889 , n386431 );
nor ( n30890 , n30884 , n30889 );
buf ( n30891 , n30890 );
nor ( n30892 , n30888 , n30891 );
or ( n30893 , n386499 , n30892 );
not ( n30894 , n22396 );
or ( n30895 , n382101 , n30894 );
nand ( n30896 , n30880 , n30893 , n30895 );
nor ( n30897 , n30874 , n30896 );
not ( n30898 , n381051 );
not ( n30899 , n20593 );
not ( n30900 , n30899 );
and ( n30901 , n30898 , n30900 );
nor ( n30902 , n30901 , n386525 );
nand ( n30903 , n20586 , n20607 );
and ( n30904 , n30903 , n20501 );
nor ( n30905 , n30904 , n386533 );
nand ( n30906 , n30902 , n30905 );
nor ( n30907 , n386512 , n30906 );
not ( n30908 , n30907 );
and ( n30909 , n30908 , RI15b4a640_403);
and ( n30910 , n19773 , n22217 );
and ( n30911 , n19768 , n19766 );
not ( n30912 , n19768 );
and ( n30913 , n30912 , RI15b4a640_403);
nor ( n387110 , n30911 , n30913 );
and ( n387111 , n387110 , n20637 );
nor ( n387112 , n30909 , n30910 , n387111 );
nand ( n387113 , n30897 , n387112 );
buf ( n387114 , n387113 );
not ( n387115 , n384523 );
nor ( n387116 , n380797 , n380805 );
not ( n387117 , n387116 );
or ( n387118 , n387115 , n387117 );
or ( n387119 , n387116 , n384523 );
nand ( n387120 , n387118 , n387119 );
buf ( n387121 , n380811 );
not ( n387122 , n387121 );
not ( n387123 , n387122 );
and ( n387124 , n387120 , n387123 );
not ( n387125 , n380821 );
not ( n387126 , n384310 );
and ( n387127 , n387125 , n387126 );
not ( n387128 , n387126 );
nand ( n387129 , n387128 , n380821 );
not ( n387130 , n387129 );
nor ( n387131 , n387127 , n387130 );
buf ( n387132 , n19391 );
not ( n387133 , n387132 );
or ( n387134 , n387131 , n387133 );
not ( n387135 , n384421 );
not ( n387136 , n387135 );
not ( n387137 , n380831 );
nor ( n387138 , n380833 , n387137 );
not ( n387139 , n387138 );
or ( n387140 , n387136 , n387139 );
or ( n387141 , n387138 , n387135 );
nand ( n387142 , n387140 , n387141 );
and ( n387143 , n387142 , n384493 );
and ( n387144 , n19513 , RI15b63f00_1275);
nor ( n387145 , n387143 , n387144 );
nand ( n387146 , n387134 , n387145 );
nor ( n387147 , n387124 , n387146 );
and ( n387148 , n19608 , RI15b63000_1243);
and ( n387149 , n386824 , n19630 );
not ( n387150 , n383444 );
and ( n387151 , n387150 , n386817 );
not ( n387152 , n387150 );
and ( n387153 , n387152 , RI15b63000_1243);
nor ( n387154 , n387151 , n387153 );
and ( n387155 , n387154 , n381497 );
nor ( n387156 , n387148 , n387149 , n387155 );
nand ( n387157 , n387147 , n387156 );
buf ( n387158 , n387157 );
buf ( n387159 , RI15b3ea48_2);
buf ( n387160 , n387159 );
buf ( n387161 , n382537 );
nor ( n387162 , n19899 , n19921 );
or ( n387163 , n387162 , n19941 );
nand ( n387164 , n387163 , n19905 );
not ( n387165 , n19997 );
nor ( n387166 , n387165 , n20502 );
or ( n387167 , n387166 , n20521 );
nand ( n387168 , n387167 , RI15b4a0a0_391);
buf ( n387169 , n19899 );
not ( n387170 , n22368 );
nor ( n387171 , n387170 , n19905 );
nand ( n387172 , n387169 , n387171 );
nor ( n387173 , n20529 , RI15b4a0a0_391);
and ( n387174 , n387165 , n387173 );
not ( n387175 , RI15b4bea0_455);
not ( n387176 , n380884 );
or ( n387177 , n387175 , n387176 );
not ( n387178 , RI15b4bea0_455);
and ( n387179 , n20568 , n20558 , n387178 );
not ( n387180 , n22390 );
and ( n387181 , n387180 , RI15b4afa0_423);
nor ( n387182 , n387179 , n387181 );
nand ( n30987 , n387177 , n387182 );
nor ( n30988 , n387174 , n30987 );
nand ( n30989 , n387164 , n387168 , n387172 , n30988 );
buf ( n30990 , n30989 );
buf ( n30991 , n382537 );
buf ( n30992 , RI15b3ea48_2);
buf ( n30993 , n30992 );
not ( n30994 , n386698 );
not ( n30995 , n383807 );
not ( n30996 , n30995 );
not ( n30997 , n386697 );
or ( n30998 , n30996 , n30997 );
nand ( n30999 , n30998 , n386695 );
not ( n31000 , n30999 );
or ( n31001 , n30994 , n31000 );
not ( n31002 , n386691 );
nor ( n31003 , n386686 , n386698 );
nand ( n31004 , n31002 , n31003 );
nand ( n31005 , n31001 , n31004 );
not ( n31006 , n31005 );
or ( n31007 , n31006 , n385002 );
not ( n31008 , n384129 );
and ( n31009 , n384130 , n31008 );
not ( n31010 , n384130 );
not ( n31011 , n31008 );
and ( n31012 , n31010 , n31011 );
nor ( n31013 , n31009 , n31012 );
nor ( n31014 , n31013 , n383851 );
nor ( n31015 , n383855 , n383686 );
or ( n31016 , n31014 , n31015 );
and ( n31017 , n31016 , n385006 );
or ( n31018 , n385019 , n21007 );
buf ( n31019 , n381357 );
buf ( n31020 , n31019 );
not ( n31021 , n31020 );
not ( n31022 , n31021 );
or ( n31023 , n31022 , n385023 );
or ( n31024 , n18123 , n383916 );
or ( n31025 , n385017 , n31024 );
nand ( n31026 , n31018 , n31023 , n31025 );
nor ( n31027 , n31017 , n31026 );
nand ( n31028 , n31007 , n31027 );
buf ( n31029 , n31028 );
buf ( n31030 , RI15b3ea48_2);
buf ( n31031 , n31030 );
buf ( n31032 , n383613 );
buf ( n31033 , RI15b3ea48_2);
buf ( n31034 , n31033 );
or ( n31035 , n379794 , RI15b60738_1156);
not ( n31036 , RI15b60c60_1167);
nor ( n31037 , n31036 , RI15b60cd8_1168);
nand ( n31038 , n31037 , RI15b60be8_1166);
not ( n31039 , n31038 );
and ( n31040 , n31039 , n22428 );
and ( n31041 , n22442 , RI15b3fa38_36);
or ( n31042 , n385043 , RI15b60c60_1167);
or ( n31043 , n385035 , n385032 );
nand ( n31044 , n22442 , n22439 );
nand ( n31045 , n31042 , n31043 , n31044 );
nor ( n31046 , n31040 , n31041 , n31045 );
nand ( n31047 , n31035 , n31046 , n22441 );
buf ( n31048 , n31047 );
buf ( n31049 , n382073 );
buf ( n31050 , n22009 );
nor ( n31051 , n22469 , n384904 );
not ( n31052 , n31051 );
and ( n31053 , n384912 , n31052 );
buf ( n31054 , n384885 );
not ( n31055 , n31054 );
not ( n31056 , n31055 );
or ( n31057 , n31053 , n31056 );
not ( n31058 , n384890 );
nand ( n31059 , n384907 , n31058 );
nand ( n31060 , RI15b60d50_1169 , RI15b60dc8_1170);
not ( n31061 , RI15b60e40_1171);
nor ( n31062 , n31060 , n31061 );
and ( n31063 , RI15b60eb8_1172 , RI15b60f30_1173);
nand ( n31064 , n31062 , n31063 );
not ( n31065 , RI15b60fa8_1174);
nor ( n31066 , n31064 , n31065 );
nand ( n31067 , n31066 , RI15b61020_1175);
not ( n31068 , n31067 );
nand ( n31069 , n31068 , RI15b61098_1176);
nor ( n31070 , n31069 , n383534 );
nand ( n31071 , n31070 , RI15b61188_1178);
not ( n31072 , n31071 );
nand ( n31073 , n31072 , RI15b61200_1179);
nand ( n31074 , RI15b61278_1180 , RI15b612f0_1181);
nor ( n31075 , n31073 , n31074 );
not ( n31076 , n31075 );
not ( n31077 , n31076 );
not ( n31078 , n19565 );
not ( n31079 , n31078 );
not ( n31080 , n31079 );
not ( n31081 , n31080 );
not ( n31082 , n31081 );
not ( n31083 , n31082 );
or ( n31084 , n31077 , n31083 );
nand ( n31085 , n19554 , n19534 );
nand ( n31086 , n22417 , n22427 );
and ( n31087 , n383588 , n31086 );
or ( n31088 , n384018 , n19495 );
nand ( n31089 , n31088 , n383927 , n19201 );
nor ( n31090 , n31087 , n19545 , n31089 );
and ( n31091 , n31085 , n31090 );
nand ( n31092 , n31084 , n31091 );
and ( n31093 , n31092 , RI15b613e0_1183);
and ( n31094 , n383945 , RI15b58a88_890);
and ( n31095 , n383949 , RI15b5a888_954);
nor ( n31096 , n31094 , n31095 );
and ( n31097 , n383955 , RI15b5b008_970);
and ( n31098 , n383960 , RI15b5ac48_962);
nor ( n31099 , n31097 , n31098 );
and ( n31100 , n383965 , RI15b5b3c8_978);
and ( n31101 , n383970 , RI15b5a108_938);
and ( n31102 , n383972 , RI15b5a4c8_946);
nor ( n31103 , n31101 , n31102 );
and ( n31104 , n383975 , RI15b59988_922);
and ( n31105 , n383977 , RI15b59d48_930);
nor ( n31106 , n31104 , n31105 );
and ( n31107 , n383982 , RI15b5bf08_1002);
and ( n31108 , n383984 , RI15b5bb48_994);
nor ( n31109 , n31107 , n31108 );
and ( n31110 , n383987 , RI15b5c2c8_1010);
and ( n31111 , n383989 , RI15b5b788_986);
nor ( n31112 , n31110 , n31111 );
nand ( n31113 , n31103 , n31106 , n31109 , n31112 );
and ( n31114 , n383968 , n31113 );
and ( n31115 , n383994 , RI15b58e48_898);
nor ( n31116 , n31100 , n31114 , n31115 );
and ( n31117 , n383997 , RI15b59208_906);
and ( n31118 , n383999 , RI15b595c8_914);
nor ( n31119 , n31117 , n31118 );
nand ( n31120 , n31096 , n31099 , n31116 , n31119 );
buf ( n31121 , n384019 );
not ( n31122 , n31121 );
not ( n31123 , n31122 );
not ( n31124 , n31123 );
not ( n31125 , n31124 );
and ( n31126 , n31120 , n31125 );
buf ( n31127 , n31078 );
buf ( n31128 , n31127 );
or ( n31129 , n31076 , n383584 , RI15b613e0_1183);
not ( n31130 , RI15b613e0_1183);
or ( n31131 , n31130 , RI15b61368_1182);
nand ( n31132 , n31129 , n31131 );
and ( n31133 , n31128 , n31132 );
nor ( n31134 , n31093 , n31126 , n31133 );
nand ( n31135 , n31057 , n31059 , n31134 );
buf ( n31136 , n31135 );
buf ( n31137 , n379895 );
not ( n31138 , n384078 );
not ( n31139 , n384081 );
and ( n31140 , n31139 , n383711 );
not ( n31141 , n31139 );
and ( n31142 , n31141 , n384103 );
nor ( n31143 , n31140 , n31142 );
not ( n31144 , n31143 );
or ( n31145 , n31138 , n31144 );
nor ( n31146 , n384710 , n383641 );
nand ( n31147 , n384117 , n31146 );
nand ( n31148 , n31145 , n31147 );
not ( n31149 , n31148 );
not ( n31150 , n383864 );
or ( n31151 , n31150 , n383894 );
or ( n31152 , n31149 , n31151 );
not ( n31153 , n383778 );
not ( n31154 , n31153 );
not ( n31155 , n383787 );
and ( n31156 , n31154 , n31155 );
and ( n31157 , n31153 , n383787 );
nor ( n31158 , n31156 , n31157 );
nor ( n31159 , n31158 , n383851 );
nor ( n31160 , n383855 , n383680 );
or ( n31161 , n31159 , n31160 );
and ( n31162 , n384165 , n383875 );
nand ( n31163 , n31162 , n383887 );
not ( n31164 , n31163 );
and ( n31165 , n31161 , n31164 );
and ( n31166 , n31163 , n31151 , n384741 );
nor ( n31167 , n31166 , n21764 );
buf ( n31168 , n383831 );
nor ( n31169 , n31168 , n383865 );
or ( n31170 , n31167 , n31169 );
nand ( n31171 , n31170 , n18154 );
nand ( n31172 , n384178 , RI15b4c1e8_462);
or ( n31173 , n383832 , n31172 );
and ( n31174 , n31171 , n31173 );
nor ( n31175 , n31174 , n383902 );
or ( n31176 , n31175 , n17599 );
not ( n31177 , n381364 );
buf ( n31178 , n31177 );
not ( n31179 , n31178 );
not ( n31180 , n31173 );
nor ( n31181 , n31169 , n31180 );
or ( n31182 , n31167 , n31181 );
or ( n31183 , n31179 , n31182 );
or ( n31184 , n17697 , n383916 );
or ( n31185 , n31173 , n31184 );
nand ( n31186 , n31176 , n31183 , n31185 );
nor ( n31187 , n31165 , n31186 );
nand ( n31188 , n31152 , n31187 );
buf ( n31189 , n31188 );
buf ( n31190 , n19655 );
not ( n31191 , n379193 );
and ( n31192 , n31191 , n379199 );
not ( n31193 , n31191 );
and ( n31194 , n31193 , n379200 );
nor ( n31195 , n31192 , n31194 );
nand ( n31196 , n31195 , RI15b58470_877);
nand ( n31197 , n22605 , RI15b57d68_862);
nand ( n31198 , n31196 , n31197 );
not ( n31199 , n31198 );
not ( n31200 , n379170 );
not ( n31201 , n379178 );
and ( n31202 , n31200 , n31201 );
not ( n31203 , n31200 );
and ( n31204 , n31203 , n379178 );
nor ( n31205 , n31202 , n31204 );
nand ( n31206 , n31205 , RI15b58470_877);
nand ( n31207 , n22605 , RI15b57c78_860);
nand ( n31208 , n31206 , n31207 );
not ( n31209 , n31208 );
not ( n31210 , n379356 );
nand ( n31211 , n22798 , n22807 );
buf ( n31212 , n31211 );
not ( n31213 , n31212 );
nand ( n31214 , n31213 , n379348 , n379357 , n379368 );
not ( n31215 , n31214 );
or ( n31216 , n31210 , n31215 );
or ( n31217 , n31214 , n379356 );
nand ( n31218 , n31216 , n31217 );
and ( n31219 , n31218 , RI15b58470_877);
not ( n31220 , n379117 );
nor ( n31221 , n31219 , n31220 );
not ( n31222 , RI15b58470_877);
not ( n31223 , n379348 );
nand ( n31224 , n379083 , n379357 );
not ( n31225 , n31224 );
or ( n31226 , n31223 , n31225 );
or ( n31227 , n31224 , n379349 );
nand ( n31228 , n31226 , n31227 );
not ( n31229 , n31228 );
or ( n31230 , n31222 , n31229 );
buf ( n31231 , n379091 );
nand ( n31232 , n31230 , n31231 );
not ( n31233 , n379357 );
nor ( n31234 , n31211 , n379082 );
not ( n31235 , n31234 );
not ( n31236 , n31235 );
or ( n31237 , n31233 , n31236 );
or ( n31238 , n31235 , n379357 );
nand ( n31239 , n31237 , n31238 );
and ( n31240 , n31239 , RI15b58470_877);
not ( n31241 , n379099 );
nor ( n31242 , n31240 , n31241 );
not ( n31243 , n379072 );
not ( n31244 , n379082 );
not ( n31245 , n31244 );
and ( n31246 , n31243 , n31245 );
and ( n31247 , n31212 , n379368 );
nor ( n31248 , n31246 , n31247 );
or ( n31249 , n31248 , n22605 );
or ( n31250 , n379078 , RI15b58470_877);
nand ( n31251 , n31249 , n31250 );
buf ( n31252 , n31212 );
nor ( n31253 , n31251 , n31252 );
nand ( n31254 , n31242 , n31253 );
nor ( n31255 , n31232 , n31254 );
nand ( n31256 , n31221 , n31255 );
not ( n31257 , n379355 );
buf ( n31258 , n379120 );
not ( n31259 , n31258 );
or ( n31260 , n31257 , n31259 );
or ( n31261 , n31258 , n379355 );
nand ( n31262 , n31260 , n31261 );
nand ( n31263 , n31262 , RI15b58470_877);
nand ( n31264 , n31263 , n379124 );
nor ( n31265 , n31256 , n31264 );
not ( n31266 , n379134 );
not ( n31267 , n31266 );
buf ( n31268 , n379126 );
not ( n31269 , n31268 );
or ( n31270 , n31267 , n31269 );
or ( n31271 , n31268 , n379354 );
nand ( n31272 , n31270 , n31271 );
and ( n31273 , n31272 , RI15b58470_877);
nor ( n31274 , n379136 , RI15b58470_877);
nor ( n31275 , n31273 , n31274 );
nand ( n31276 , n31265 , n31275 );
buf ( n31277 , n379135 );
and ( n31278 , n31277 , n379145 );
not ( n31279 , n31277 );
and ( n31280 , n31279 , n379374 );
nor ( n31281 , n31278 , n31280 );
nand ( n31282 , n31281 , RI15b58470_877);
nand ( n31283 , n22605 , RI15b57a98_856);
nand ( n31284 , n31282 , n31283 );
nor ( n31285 , n31276 , n31284 );
not ( n31286 , n379070 );
not ( n31287 , n31286 );
not ( n31288 , n31287 );
buf ( n31289 , n379146 );
not ( n31290 , n31289 );
or ( n31291 , n31288 , n31290 );
not ( n31292 , n31286 );
or ( n31293 , n31289 , n31292 );
nand ( n31294 , n31291 , n31293 );
and ( n31295 , n31294 , RI15b58470_877);
not ( n31296 , n379069 );
nor ( n31297 , n31295 , n31296 );
nand ( n31298 , n31285 , n31297 );
not ( n31299 , n31298 );
and ( n31300 , n22605 , RI15b57b88_858);
not ( n31301 , n22605 );
and ( n31302 , n379147 , n379158 );
not ( n31303 , n379147 );
not ( n31304 , n379158 );
and ( n31305 , n31303 , n31304 );
nor ( n31306 , n31302 , n31305 );
and ( n31307 , n31301 , n31306 );
nor ( n31308 , n31300 , n31307 );
nand ( n31309 , n31299 , n31308 );
not ( n31310 , n379159 );
and ( n31311 , n31310 , n379167 );
not ( n31312 , n31310 );
and ( n31313 , n31312 , n379168 );
nor ( n31314 , n31311 , n31313 );
nand ( n31315 , n31314 , RI15b58470_877);
nand ( n31316 , n22605 , RI15b57c00_859);
nand ( n31317 , n31315 , n31316 );
nor ( n31318 , n31309 , n31317 );
nand ( n31319 , n31209 , n31318 );
buf ( n31320 , n379179 );
and ( n31321 , n31320 , n379192 );
not ( n31322 , n31320 );
and ( n31323 , n31322 , n379191 );
nor ( n31324 , n31321 , n31323 );
nand ( n31325 , n31324 , RI15b58470_877);
nand ( n31326 , n22605 , RI15b57cf0_861);
nand ( n31327 , n31325 , n31326 );
nor ( n31328 , n31319 , n31327 );
nand ( n31329 , n31199 , n31328 );
not ( n31330 , n379218 );
not ( n31331 , n31330 );
nor ( n31332 , n379201 , n22605 );
not ( n31333 , n31332 );
or ( n31334 , n31331 , n31333 );
nand ( n31335 , n379201 , RI15b58470_877);
not ( n31336 , n31335 );
not ( n31337 , n31330 );
and ( n31338 , n31336 , n31337 );
and ( n31339 , n22605 , RI15b57de0_863);
nor ( n31340 , n31338 , n31339 );
nand ( n31341 , n31334 , n31340 );
nor ( n31342 , n31329 , n31341 );
not ( n31343 , RI15b58470_877);
not ( n31344 , n31330 );
or ( n31345 , n31343 , n31344 );
nand ( n31346 , n31345 , n31335 );
and ( n31347 , n31346 , n379206 );
nor ( n31348 , n379206 , n31330 );
not ( n31349 , n31348 );
not ( n31350 , n31332 );
or ( n31351 , n31349 , n31350 );
nand ( n31352 , n22605 , RI15b57e58_864);
nand ( n31353 , n31351 , n31352 );
nor ( n31354 , n31347 , n31353 );
nand ( n31355 , n31342 , n31354 );
buf ( n31356 , n31332 );
buf ( n31357 , n379219 );
not ( n31358 , n379229 );
nor ( n31359 , n31357 , n31358 );
and ( n31360 , n31356 , n31359 );
and ( n31361 , n22605 , RI15b57ed0_865);
nor ( n31362 , n31360 , n31361 );
nand ( n31363 , n31357 , RI15b58470_877);
not ( n31364 , n31363 );
not ( n31365 , n31335 );
or ( n31366 , n31364 , n31365 );
nand ( n31367 , n31366 , n31358 );
nand ( n31368 , n31362 , n31367 );
nor ( n31369 , n31355 , n31368 );
buf ( n31370 , n31335 );
nand ( n31371 , n31370 , n379230 );
and ( n31372 , n31371 , n379237 );
not ( n31373 , n379230 );
nor ( n31374 , n31373 , n379237 );
not ( n31375 , n31374 );
not ( n31376 , n31356 );
not ( n31377 , n31376 );
not ( n31378 , n31377 );
or ( n31379 , n31375 , n31378 );
nand ( n31380 , n22605 , RI15b57f48_866);
nand ( n31381 , n31379 , n31380 );
nor ( n31382 , n31372 , n31381 );
nand ( n31383 , n31369 , n31382 );
buf ( n31384 , n31383 );
not ( n31385 , n31384 );
not ( n31386 , n31376 );
not ( n31387 , n379238 );
and ( n31388 , n31387 , n379248 );
and ( n31389 , n31386 , n31388 );
and ( n31390 , n22605 , RI15b57fc0_867);
nor ( n31391 , n31389 , n31390 );
not ( n31392 , n31387 );
not ( n31393 , n31370 );
or ( n31394 , n31392 , n31393 );
not ( n31395 , n379248 );
nand ( n31396 , n31394 , n31395 );
nand ( n31397 , n31391 , n31396 );
not ( n31398 , n31397 );
nand ( n31399 , n31370 , n379249 );
and ( n31400 , n31399 , n379262 );
not ( n31401 , RI15b58038_868);
not ( n31402 , n22605 );
or ( n31403 , n31401 , n31402 );
not ( n31404 , n379262 );
nand ( n31405 , n31386 , n379249 , n31404 );
nand ( n31406 , n31403 , n31405 );
nor ( n31407 , n31400 , n31406 );
buf ( n31408 , n379264 );
buf ( n31409 , n379272 );
buf ( n31410 , n31409 );
not ( n31411 , n31410 );
and ( n31412 , n31408 , n31411 );
not ( n31413 , n31408 );
and ( n31414 , n31413 , n31410 );
nor ( n31415 , n31412 , n31414 );
and ( n31416 , n31385 , n31398 , n31407 , n31415 );
buf ( n31417 , n379273 );
not ( n31418 , n31417 );
not ( n31419 , n31418 );
not ( n31420 , n379286 );
not ( n31421 , n31420 );
and ( n31422 , n31419 , n31421 );
and ( n31423 , n31418 , n31420 );
nor ( n31424 , n31422 , n31423 );
nand ( n31425 , n31416 , n31424 );
not ( n31426 , n31425 );
not ( n31427 , n31426 );
nand ( n31428 , n31418 , n379286 );
xor ( n31429 , n31428 , n379280 );
not ( n31430 , n31429 );
not ( n31431 , n31430 );
and ( n31432 , n31427 , n31431 );
and ( n31433 , n31426 , n31430 );
nor ( n31434 , n31432 , n31433 );
buf ( n31435 , n31434 );
not ( n31436 , n31435 );
not ( n31437 , n31383 );
not ( n31438 , n31397 );
nand ( n31439 , n31437 , n31438 );
not ( n31440 , n31439 );
nand ( n31441 , n31440 , n31407 );
nor ( n31442 , n31441 , n31415 );
not ( n31443 , n31442 );
or ( n31444 , n31408 , n31410 );
nand ( n31445 , n31444 , n31417 );
nand ( n31446 , n31441 , n31445 );
not ( n31447 , n31439 );
not ( n31448 , n31447 );
not ( n31449 , n31407 );
not ( n31450 , n31449 );
and ( n31451 , n31448 , n31450 );
and ( n31452 , n31447 , n31449 );
nor ( n31453 , n31451 , n31452 );
not ( n31454 , n31384 );
not ( n31455 , n31438 );
and ( n31456 , n31454 , n31455 );
and ( n31457 , n31384 , n31398 );
nor ( n31458 , n31456 , n31457 );
and ( n31459 , n379332 , n379048 , n379299 );
not ( n31460 , n31459 );
not ( n31461 , n379290 );
or ( n31462 , n31460 , n31461 );
not ( n31463 , n31317 );
and ( n31464 , n31309 , n31463 );
not ( n31465 , n31309 );
and ( n31466 , n31465 , n31317 );
nor ( n31467 , n31464 , n31466 );
not ( n31468 , n31308 );
not ( n31469 , n31468 );
not ( n31470 , n31299 );
or ( n31471 , n31469 , n31470 );
buf ( n31472 , n31299 );
or ( n31473 , n31472 , n31468 );
nand ( n31474 , n31471 , n31473 );
not ( n31475 , n31284 );
and ( n31476 , n31276 , n31475 );
not ( n31477 , n31276 );
and ( n31478 , n31477 , n31284 );
nor ( n31479 , n31476 , n31478 );
buf ( n31480 , n31265 );
nor ( n31481 , n31480 , n31275 );
not ( n31482 , n31481 );
nand ( n31483 , n31482 , n31276 );
not ( n31484 , n31221 );
xnor ( n31485 , n31484 , n31255 );
not ( n31486 , n31485 );
buf ( n31487 , n31256 );
not ( n31488 , n31264 );
and ( n31489 , n31487 , n31488 );
not ( n31490 , n31487 );
not ( n31491 , n31488 );
and ( n31492 , n31490 , n31491 );
nor ( n31493 , n31489 , n31492 );
nand ( n31494 , n31486 , n31493 );
buf ( n31495 , n31232 );
not ( n31496 , n31495 );
not ( n31497 , n31254 );
not ( n31498 , n31497 );
and ( n31499 , n31496 , n31498 );
and ( n31500 , n31495 , n31497 );
nor ( n31501 , n31499 , n31500 );
buf ( n31502 , n31253 );
not ( n31503 , n31502 );
not ( n31504 , n31242 );
not ( n31505 , n31504 );
or ( n31506 , n31503 , n31505 );
buf ( n31507 , n31502 );
or ( n31508 , n31504 , n31507 );
nand ( n31509 , n31506 , n31508 );
nand ( n31510 , n31507 , RI15b58470_877);
nor ( n31511 , n31509 , n31510 );
nand ( n31512 , n31501 , n31511 );
nor ( n31513 , n31494 , n31512 );
nand ( n31514 , n31479 , n31483 , n31513 );
not ( n31515 , n31514 );
not ( n31516 , n31285 );
not ( n31517 , n31516 );
buf ( n31518 , n31297 );
not ( n31519 , n31518 );
and ( n31520 , n31517 , n31519 );
and ( n31521 , n31516 , n31518 );
nor ( n31522 , n31520 , n31521 );
nand ( n31523 , n31515 , n31522 );
nor ( n31524 , n31474 , n31523 );
and ( n31525 , n31467 , n31524 );
nand ( n31526 , n31462 , n31525 );
buf ( n31527 , n31208 );
not ( n31528 , n31527 );
buf ( n31529 , n31318 );
not ( n31530 , n31529 );
or ( n31531 , n31528 , n31530 );
buf ( n31532 , n31527 );
or ( n31533 , n31529 , n31532 );
nand ( n31534 , n31531 , n31533 );
nor ( n31535 , n31526 , n31534 );
buf ( n31536 , n31319 );
buf ( n31537 , n31327 );
not ( n31538 , n31537 );
and ( n31539 , n31536 , n31538 );
not ( n31540 , n31536 );
and ( n31541 , n31540 , n31537 );
nor ( n31542 , n31539 , n31541 );
nand ( n31543 , n31535 , n31542 );
buf ( n31544 , n31328 );
buf ( n31545 , n31198 );
buf ( n31546 , n31545 );
or ( n31547 , n31544 , n31546 );
nand ( n31548 , n31544 , n31545 );
nand ( n31549 , n31547 , n31548 );
nor ( n31550 , n31543 , n31549 );
buf ( n31551 , n31329 );
buf ( n31552 , n31341 );
not ( n31553 , n31552 );
and ( n31554 , n31551 , n31553 );
not ( n31555 , n31551 );
and ( n31556 , n31555 , n31552 );
nor ( n31557 , n31554 , n31556 );
nand ( n31558 , n31550 , n31557 );
not ( n31559 , n31354 );
not ( n31560 , n31559 );
buf ( n31561 , n31342 );
not ( n31562 , n31561 );
or ( n31563 , n31560 , n31562 );
or ( n31564 , n31561 , n31559 );
nand ( n31565 , n31563 , n31564 );
nor ( n31566 , n31558 , n31565 );
buf ( n31567 , n31355 );
not ( n31568 , n31368 );
and ( n31569 , n31567 , n31568 );
not ( n31570 , n31567 );
and ( n31571 , n31570 , n31368 );
nor ( n31572 , n31569 , n31571 );
and ( n31573 , n31566 , n31572 );
not ( n31574 , n31369 );
buf ( n31575 , n31382 );
and ( n31576 , n31574 , n31575 );
not ( n31577 , n31574 );
not ( n31578 , n31575 );
and ( n31579 , n31577 , n31578 );
nor ( n31580 , n31576 , n31579 );
nand ( n31581 , n31458 , n31573 , n31580 );
not ( n31582 , n31581 );
nand ( n31583 , n31443 , n31446 , n31453 , n31582 );
not ( n31584 , n31583 );
and ( n31585 , n31385 , n31398 , n31407 , n31415 );
not ( n31586 , n31585 );
not ( n31587 , n31424 );
not ( n31588 , n31587 );
and ( n31589 , n31586 , n31588 );
and ( n31590 , n31585 , n31587 );
nor ( n31591 , n31589 , n31590 );
nand ( n31592 , n31584 , n31591 );
buf ( n31593 , n31592 );
not ( n31594 , n31593 );
and ( n31595 , n31436 , n31594 );
not ( n31596 , n31436 );
and ( n31597 , n31596 , n31593 );
nor ( n31598 , n31595 , n31597 );
buf ( n31599 , n379342 );
not ( n31600 , n31599 );
not ( n31601 , n31600 );
buf ( n31602 , n31601 );
not ( n31603 , n31602 );
or ( n31604 , n31598 , n31603 );
not ( n31605 , n379356 );
not ( n31606 , n379380 );
or ( n31607 , n31605 , n31606 );
nand ( n31608 , n31607 , n379117 );
not ( n31609 , n31608 );
not ( n31610 , n31609 );
nor ( n31611 , n22799 , n22605 );
not ( n31612 , n31611 );
not ( n31613 , n379379 );
or ( n31614 , n31612 , n31613 );
nand ( n31615 , n22605 , RI15b57750_849);
nand ( n31616 , n31614 , n31615 );
nand ( n31617 , n379380 , n31616 , n379370 );
not ( n31618 , n31617 );
not ( n31619 , n379358 );
not ( n31620 , n31619 );
not ( n31621 , n379380 );
or ( n31622 , n31620 , n31621 );
nand ( n31623 , n31622 , n379099 );
nand ( n31624 , n31618 , n31623 );
not ( n31625 , n379350 );
not ( n31626 , n379380 );
or ( n31627 , n31625 , n31626 );
buf ( n31628 , n31231 );
nand ( n31629 , n31627 , n31628 );
nor ( n31630 , n31624 , n31629 );
nand ( n31631 , n31610 , n31630 );
not ( n31632 , n379355 );
not ( n31633 , n379381 );
or ( n31634 , n31632 , n31633 );
nand ( n31635 , n31634 , n379124 );
not ( n31636 , n31635 );
nor ( n31637 , n31631 , n31636 );
buf ( n31638 , n379354 );
not ( n31639 , n31638 );
and ( n31640 , n31637 , n31639 );
not ( n31641 , n31292 );
not ( n31642 , n379381 );
or ( n31643 , n31641 , n31642 );
nand ( n31644 , n31643 , n379069 );
not ( n31645 , n379199 );
not ( n31646 , n379381 );
or ( n31647 , n31645 , n31646 );
nand ( n31648 , n31647 , n31197 );
nor ( n31649 , n31644 , n31648 );
not ( n31650 , n379376 );
and ( n31651 , n31649 , n31650 );
nand ( n31652 , n31640 , n31651 );
not ( n31653 , n379382 );
or ( n31654 , n31653 , n379237 );
nand ( n31655 , n31654 , n31380 );
nor ( n31656 , n31655 , n31373 );
nor ( n31657 , n31404 , n379248 );
nand ( n31658 , n31656 , n31657 );
nor ( n31659 , n31652 , n31658 );
not ( n31660 , n379382 );
or ( n31661 , n31660 , n31409 );
or ( n31662 , n22835 , RI15b58470_877);
nand ( n31663 , n31661 , n31662 );
not ( n31664 , n31663 );
and ( n31665 , n31659 , n31664 );
not ( n31666 , n31665 );
not ( n31667 , n379391 );
or ( n31668 , n31666 , n31667 );
not ( n31669 , n379330 );
not ( n31670 , n379382 );
or ( n31671 , n31669 , n31670 );
nand ( n31672 , n31671 , n379327 );
not ( n31673 , RI15b581a0_871);
not ( n31674 , n22605 );
or ( n31675 , n31673 , n31674 );
nand ( n31676 , n31675 , n379280 );
not ( n31677 , n31676 );
nand ( n31678 , n22605 , RI15b58128_870);
and ( n31679 , n379286 , n31678 );
nand ( n31680 , n31677 , n379319 , n31395 , n31679 );
not ( n31681 , n31680 );
not ( n31682 , RI15b58290_873);
not ( n31683 , n22605 );
or ( n31684 , n31682 , n31683 );
buf ( n31685 , n379312 );
nand ( n31686 , n31684 , n31685 );
not ( n31687 , n31686 );
nand ( n31688 , n31681 , n31687 , n379377 , n379045 );
nor ( n31689 , n31663 , n31672 , n31688 );
not ( n31690 , n379300 );
not ( n31691 , n31690 );
not ( n31692 , n379382 );
or ( n31693 , n31691 , n31692 );
nand ( n31694 , n22605 , RI15b58218_872);
nand ( n31695 , n31693 , n31694 );
nor ( n31696 , n31695 , n31629 );
nand ( n31697 , n31689 , n31656 , n31649 , n31696 );
nand ( n31698 , n31697 , n379383 );
and ( n31699 , n31698 , n379391 );
not ( n31700 , n31699 );
nand ( n31701 , n31668 , n31700 );
not ( n31702 , n31679 );
and ( n31703 , n31701 , n31702 );
not ( n31704 , n31698 );
nand ( n31705 , n31704 , n379391 );
not ( n31706 , n31705 );
not ( n31707 , n31706 );
not ( n31708 , n31707 );
not ( n31709 , n31708 );
or ( n31710 , n31665 , n31709 , n31702 );
and ( n31711 , n379394 , RI15b581a0_871);
buf ( n31712 , n379398 );
and ( n31713 , n31712 , RI15b51fa8_662);
nor ( n31714 , n31711 , n31713 );
nand ( n31715 , n31710 , n31714 );
nor ( n31716 , n31703 , n31715 );
nand ( n31717 , n31604 , n31716 );
buf ( n31718 , n31717 );
buf ( n31719 , RI15b3ea48_2);
buf ( n31720 , n31719 );
not ( n31721 , n384403 );
buf ( n31722 , n384480 );
not ( n31723 , n31722 );
or ( n31724 , n31721 , n31723 );
or ( n31725 , n31722 , n384403 );
nand ( n31726 , n31724 , n31725 );
buf ( n31727 , n384493 );
nand ( n31728 , n31726 , n31727 );
nor ( n31729 , n384378 , n384383 );
not ( n31730 , n31729 );
nand ( n31731 , n31730 , n384385 );
nand ( n31732 , n31731 , n387132 );
not ( n31733 , n19512 );
not ( n31734 , n379445 );
and ( n31735 , n31733 , n31734 );
not ( n31736 , n384605 );
not ( n31737 , n31736 );
not ( n31738 , n384598 );
or ( n31739 , n31737 , n31738 );
or ( n31740 , n384598 , n31736 );
nand ( n31741 , n31739 , n31740 );
and ( n31742 , n31741 , n380811 );
nor ( n31743 , n31735 , n31742 );
and ( n31744 , n31728 , n31732 , n31743 );
buf ( n31745 , n384400 );
not ( n31746 , n31745 );
not ( n31747 , n31746 );
buf ( n31748 , n31747 );
not ( n31749 , n31748 );
not ( n31750 , n31749 );
nor ( n31751 , n384017 , n383926 );
or ( n31752 , n31750 , n31751 );
not ( n31753 , n22418 );
nand ( n31754 , n19553 , n31753 );
not ( n31755 , n31754 );
and ( n31756 , n383588 , n22428 );
nand ( n31757 , n22444 , n22427 );
and ( n31758 , n19545 , n31757 );
nor ( n31759 , n31756 , n31758 );
not ( n31760 , n31759 );
or ( n31761 , n31755 , n31760 );
nand ( n31762 , n31761 , n19201 );
not ( n31763 , n19484 );
nand ( n31764 , n31763 , n31751 );
nand ( n31765 , n31764 , n19496 );
nor ( n31766 , n383598 , n19580 );
nand ( n31767 , n31765 , n31766 , n19600 , n19590 );
not ( n31768 , n19572 );
nor ( n31769 , n31767 , n31768 );
nand ( n31770 , n31762 , n31769 );
not ( n31771 , n31770 );
nand ( n31772 , n31752 , n31771 );
and ( n31773 , n31772 , RI15b5cef8_1036);
not ( n31774 , n31747 );
buf ( n31775 , n31774 );
not ( n31776 , n384018 );
and ( n31777 , n31776 , n19495 );
or ( n31778 , n31777 , n386746 );
not ( n31779 , n31778 );
or ( n31780 , n31775 , n31779 , RI15b5cef8_1036);
buf ( n31781 , n19566 );
not ( n31782 , n31781 );
buf ( n31783 , n31782 );
buf ( n31784 , n31783 );
or ( n31785 , n31784 , n384383 );
nand ( n31786 , n31780 , n31785 );
not ( n31787 , n383503 );
nor ( n31788 , n31787 , n22428 );
or ( n31789 , n19556 , n19200 );
nor ( n31790 , n31051 , n384906 );
nand ( n31791 , n31789 , n31790 );
or ( n31792 , n31788 , n31791 );
not ( n31793 , n31792 );
nor ( n31794 , n31793 , n384605 );
nor ( n31795 , n31773 , n31786 , n31794 );
nand ( n31796 , n31744 , n31795 );
buf ( n31797 , n31796 );
buf ( n31798 , n19765 );
not ( n31799 , n22345 );
or ( n31800 , n31798 , n31799 );
nand ( n31801 , n31800 , n19938 );
nand ( n31802 , n31801 , n19773 );
not ( n31803 , n19773 );
nand ( n31804 , n31803 , n383353 , n31798 );
and ( n31805 , n20641 , RI15b4b540_435);
not ( n31806 , n20502 );
buf ( n31807 , n19964 );
and ( n31808 , n31806 , n31807 );
and ( n31809 , n22383 , n20501 );
nor ( n31810 , n31808 , n31809 );
or ( n31811 , n31810 , n19965 );
not ( n31812 , n20538 );
and ( n31813 , n31812 , RI15b4b540_435);
not ( n31814 , n31812 );
and ( n31815 , n31814 , n382101 );
nor ( n31816 , n31813 , n31815 );
or ( n31817 , n31816 , n22354 );
not ( n31818 , n31807 );
and ( n31819 , n22361 , n31818 , n19965 );
or ( n31820 , n20653 , n19766 );
not ( n31821 , n22394 );
nand ( n31822 , n31820 , n31821 );
nor ( n31823 , n31819 , n31822 );
nand ( n31824 , n31811 , n31817 , n31823 );
nor ( n31825 , n31805 , n31824 );
nand ( n31826 , n31802 , n31804 , n31825 );
buf ( n31827 , n31826 );
buf ( n31828 , n22402 );
buf ( n31829 , n384700 );
buf ( n31830 , n386760 );
buf ( n31831 , n22788 );
nor ( n31832 , n384481 , n384486 );
not ( n31833 , n31745 );
not ( n31834 , n31833 );
not ( n31835 , RI15b5cfe8_1038);
or ( n31836 , n31834 , n31835 );
nand ( n31837 , RI15b5cef8_1036 , RI15b5cf70_1037);
nor ( n31838 , n31837 , RI15b5cfe8_1038);
nand ( n31839 , n31834 , n31838 );
nand ( n31840 , n31837 , RI15b5cfe8_1038);
nand ( n31841 , n31836 , n31839 , n31840 );
nand ( n31842 , n31832 , n31841 );
nor ( n31843 , n31837 , n31835 );
not ( n31844 , n31843 );
nor ( n31845 , n31844 , RI15b5d060_1039);
nand ( n31846 , n31747 , n31845 );
nand ( n31847 , n31746 , RI15b5d060_1039);
nand ( n31848 , n31844 , RI15b5d060_1039);
and ( n31849 , n31846 , n31847 , n31848 );
nor ( n31850 , n31842 , n31849 );
and ( n31851 , n31746 , RI15b5d0d8_1040);
nand ( n31852 , n31843 , RI15b5d060_1039);
or ( n31853 , n31852 , RI15b5d0d8_1040);
or ( n31854 , n31833 , n31853 );
nand ( n31855 , n31852 , RI15b5d0d8_1040);
nand ( n31856 , n31854 , n31855 );
nor ( n31857 , n31851 , n31856 );
not ( n31858 , n31857 );
and ( n31859 , n31850 , n31858 );
nand ( n31860 , n31749 , RI15b5d150_1041);
not ( n31861 , n31852 );
nand ( n31862 , n31861 , RI15b5d0d8_1040);
nor ( n31863 , n31862 , RI15b5d150_1041);
nand ( n31864 , n31748 , n31863 );
nand ( n31865 , n31862 , RI15b5d150_1041);
and ( n31866 , n31860 , n31864 , n31865 );
not ( n31867 , n31866 );
nand ( n31868 , n31859 , n31867 );
and ( n31869 , n31774 , RI15b5d1c8_1042);
not ( n31870 , n31862 );
nand ( n31871 , n31870 , RI15b5d150_1041);
or ( n31872 , n31871 , RI15b5d1c8_1042);
or ( n31873 , n31746 , n31872 );
nand ( n31874 , n31871 , RI15b5d1c8_1042);
nand ( n31875 , n31873 , n31874 );
nor ( n31876 , n31869 , n31875 );
and ( n31877 , n31868 , n31876 );
not ( n31878 , n31868 );
not ( n31879 , n31876 );
and ( n31880 , n31878 , n31879 );
nor ( n31881 , n31877 , n31880 );
not ( n31882 , n384494 );
not ( n31883 , n31882 );
not ( n31884 , n31883 );
nand ( n31885 , n31881 , n31884 );
and ( n31886 , n384379 , RI15b5cfe8_1038);
not ( n31887 , n31838 );
not ( n31888 , n384244 );
or ( n31889 , n31887 , n31888 );
nand ( n31890 , n31889 , n31840 );
nor ( n31891 , n31886 , n31890 );
and ( n31892 , n384388 , n31891 );
and ( n31893 , n384379 , RI15b5d060_1039);
not ( n31894 , n31845 );
not ( n31895 , n384244 );
or ( n31896 , n31894 , n31895 );
nand ( n31897 , n31896 , n31848 );
nor ( n31898 , n31893 , n31897 );
nand ( n31899 , n31892 , n31898 );
nand ( n31900 , n384379 , RI15b5d0d8_1040);
not ( n31901 , n31853 );
nand ( n31902 , n31901 , n384244 );
nand ( n31903 , n31900 , n31902 , n31855 );
nor ( n31904 , n31899 , n31903 );
and ( n31905 , n384379 , RI15b5d150_1041);
not ( n31906 , n31863 );
not ( n31907 , n384244 );
or ( n31908 , n31906 , n31907 );
nand ( n31909 , n31908 , n31865 );
nor ( n31910 , n31905 , n31909 );
nand ( n31911 , n31904 , n31910 );
not ( n31912 , n31911 );
and ( n31913 , n384379 , RI15b5d1c8_1042);
or ( n31914 , n384379 , n31872 );
nand ( n31915 , n31914 , n31874 );
nor ( n31916 , n31913 , n31915 );
nor ( n31917 , n31912 , n31916 );
not ( n31918 , n31917 );
nand ( n31919 , n31912 , n31916 );
nand ( n31920 , n31918 , n31919 );
buf ( n31921 , n387132 );
not ( n31922 , n31921 );
not ( n31923 , n31922 );
nand ( n31924 , n31920 , n31923 );
not ( n31925 , RI15b5d1c8_1042);
or ( n31926 , n384600 , n31925 );
or ( n31927 , n384601 , n31872 );
nand ( n31928 , n31926 , n31927 , n31874 );
not ( n31929 , n31928 );
and ( n31930 , n384606 , n384612 );
or ( n31931 , n384600 , n31835 );
nand ( n31932 , n384600 , n31838 );
nand ( n31933 , n31931 , n31932 , n31840 );
nand ( n31934 , n31930 , n31933 );
and ( n31935 , n384601 , RI15b5d060_1039);
not ( n31936 , n31845 );
not ( n31937 , n384600 );
or ( n31938 , n31936 , n31937 );
nand ( n31939 , n31938 , n31848 );
nor ( n31940 , n31935 , n31939 );
nor ( n31941 , n31934 , n31940 );
or ( n31942 , n384601 , n31853 );
nand ( n31943 , n384601 , RI15b5d0d8_1040);
nand ( n31944 , n31942 , n31943 , n31855 );
and ( n31945 , n31941 , n31944 );
and ( n31946 , n384601 , RI15b5d150_1041);
not ( n31947 , n31863 );
not ( n31948 , n384600 );
or ( n31949 , n31947 , n31948 );
nand ( n31950 , n31949 , n31865 );
nor ( n31951 , n31946 , n31950 );
not ( n31952 , n31951 );
nand ( n31953 , n31945 , n31952 );
not ( n31954 , n31953 );
or ( n31955 , n31929 , n31954 );
or ( n31956 , n31953 , n31928 );
nand ( n31957 , n31955 , n31956 );
buf ( n31958 , n380812 );
not ( n31959 , n31958 );
buf ( n31960 , n31959 );
nand ( n31961 , n31957 , n31960 );
nand ( n31962 , n19513 , RI15b64860_1295);
and ( n31963 , n31885 , n31924 , n31961 , n31962 );
buf ( n31964 , n384624 );
buf ( n31965 , n31964 );
not ( n31966 , n31965 );
not ( n31967 , n383430 );
or ( n31968 , n31966 , n31967 );
nand ( n31969 , n31968 , n384642 );
and ( n31970 , n31969 , RI15b63960_1263);
not ( n31971 , n384655 );
or ( n31972 , n31971 , n383430 , RI15b63960_1263);
nand ( n31973 , n386954 , n19630 );
nand ( n31974 , n31972 , n31973 );
nor ( n31975 , n31970 , n31974 );
nand ( n31976 , n31963 , n31975 );
buf ( n31977 , n31976 );
buf ( n31978 , n384996 );
buf ( n31979 , RI15b3ea48_2);
buf ( n31980 , n31979 );
buf ( n31981 , n382067 );
and ( n31982 , n382467 , n382489 );
not ( n31983 , n382515 );
not ( n31984 , n382434 );
or ( n31985 , n31983 , n31984 );
not ( n31986 , RI15b4c008_458);
nand ( n31987 , n31986 , RI15b4b540_435);
nand ( n31988 , n31985 , n31987 );
not ( n31989 , n31988 );
nand ( n31990 , n31982 , n31989 );
not ( n31991 , n382434 );
buf ( n31992 , n382240 );
or ( n31993 , n31991 , n31992 );
not ( n31994 , RI15b4c008_458);
nand ( n31995 , n31994 , RI15b4b5b8_436);
nand ( n31996 , n31993 , n31995 );
buf ( n31997 , n382303 );
or ( n31998 , n31991 , n31997 );
not ( n31999 , RI15b4c008_458);
nand ( n32000 , n31999 , RI15b4b6a8_438);
nand ( n32001 , n31998 , n32000 );
nor ( n32002 , n31996 , n32001 );
not ( n32003 , n382433 );
not ( n32004 , n32003 );
buf ( n32005 , n382295 );
or ( n32006 , n32004 , n32005 );
not ( n32007 , RI15b4c008_458);
nand ( n32008 , n32007 , RI15b4b630_437);
nand ( n32009 , n32006 , n32008 );
not ( n32010 , n382322 );
not ( n32011 , n32010 );
not ( n32012 , n32003 );
or ( n32013 , n32011 , n32012 );
not ( n32014 , RI15b4c008_458);
nand ( n32015 , n32014 , RI15b4b720_439);
nand ( n32016 , n32013 , n32015 );
nor ( n32017 , n32009 , n32016 );
nand ( n32018 , n32002 , n32017 );
buf ( n32019 , n32018 );
nor ( n32020 , n31990 , n32019 );
not ( n32021 , n32020 );
nor ( n32022 , n32021 , n382079 );
buf ( n32023 , n382474 );
not ( n32024 , n32023 );
or ( n32025 , n32022 , n32024 );
not ( n32026 , n382335 );
not ( n32027 , n32003 );
or ( n32028 , n32026 , n32027 );
not ( n32029 , RI15b4c008_458);
nand ( n32030 , n32029 , RI15b4b798_440);
nand ( n32031 , n32028 , n32030 );
nand ( n32032 , n32025 , n32031 );
not ( n32033 , n382473 );
nand ( n32034 , n32033 , n382080 );
buf ( n32035 , n32034 );
not ( n32036 , n32035 );
not ( n32037 , n32031 );
and ( n32038 , n32021 , n32036 , n32037 );
buf ( n32039 , n382305 );
not ( n32040 , n32039 );
nor ( n32041 , n32040 , n32010 );
not ( n32042 , n32041 );
nor ( n32043 , n32042 , n382335 );
not ( n32044 , n32043 );
not ( n32045 , n382316 );
not ( n32046 , n32045 );
and ( n32047 , n32044 , n32046 );
and ( n32048 , n32043 , n32045 );
nor ( n32049 , n32047 , n32048 );
or ( n32050 , n382513 , n32049 );
and ( n32051 , n382523 , RI15b4b810_441);
buf ( n32052 , n382528 );
and ( n32053 , n32052 , RI15b45618_232);
nor ( n32054 , n32051 , n32053 );
nand ( n32055 , n32050 , n32054 );
nor ( n32056 , n32038 , n32055 );
nand ( n32057 , n32032 , n32056 );
buf ( n32058 , n32057 );
buf ( n32059 , n22479 );
buf ( n32060 , n380940 );
not ( n32061 , n380729 );
buf ( n32062 , n32061 );
buf ( n32063 , n32062 );
not ( n32064 , n32063 );
not ( n32065 , n32064 );
not ( n32066 , n380703 );
or ( n32067 , n32065 , n32066 );
nand ( n32068 , n380741 , n380765 );
or ( n32069 , n382980 , n32068 );
not ( n32070 , n32069 );
and ( n32071 , n380719 , n32070 );
not ( n32072 , n380749 );
and ( n32073 , n32069 , n32061 , n32072 );
nor ( n32074 , n32073 , n19630 );
not ( n32075 , n380219 );
or ( n32076 , n32074 , n32075 );
nand ( n32077 , n32076 , n19595 );
not ( n32078 , n380763 );
or ( n32079 , n380207 , n32078 );
nand ( n32080 , n32077 , n32079 );
and ( n32081 , n32080 , n380775 );
not ( n32082 , RI15b5a540_947);
or ( n32083 , n32081 , n32082 );
not ( n32084 , n32079 );
nor ( n32085 , n32075 , n32084 );
or ( n32086 , n32074 , n32085 );
or ( n32087 , n380782 , n32086 );
or ( n32088 , n32079 , n380790 );
nand ( n32089 , n32083 , n32087 , n32088 );
nor ( n32090 , n32071 , n32089 );
nand ( n32091 , n32067 , n32090 );
buf ( n32092 , n32091 );
buf ( n32093 , n379403 );
not ( n32094 , RI15b54960_751);
or ( n32095 , n382679 , n32094 );
buf ( n32096 , n21204 );
not ( n32097 , n32096 );
or ( n32098 , n32097 , n382886 );
and ( n32099 , n382677 , n18182 , n383906 );
not ( n32100 , RI15b548e8_750);
or ( n32101 , n32100 , RI15b54960_751);
or ( n32102 , n32094 , RI15b548e8_750);
nand ( n32103 , n32101 , n32102 );
and ( n32104 , n382626 , n32103 );
nor ( n32105 , n32099 , n32104 );
nand ( n32106 , n32095 , n32098 , n32105 );
buf ( n32107 , n32106 );
buf ( n32108 , n22408 );
buf ( n32109 , n20663 );
buf ( n32110 , n381566 );
or ( n32111 , n384961 , n22151 );
and ( n32112 , n384983 , n22211 );
not ( n32113 , RI15b40938_68);
or ( n32114 , n22237 , n32113 );
or ( n32115 , n22022 , n22296 );
or ( n32116 , n22228 , n384988 );
nand ( n32117 , n32114 , n32115 , n32116 );
nor ( n32118 , n32112 , n32117 );
nand ( n32119 , n32111 , n32118 );
buf ( n32120 , n32119 );
not ( n32121 , n22151 );
not ( n32122 , n32121 );
xor ( n32123 , RI15b66408_1354 , n381889 );
xnor ( n32124 , n32123 , n381887 );
and ( n32125 , n32124 , n22097 );
not ( n32126 , RI15b66408_1354);
nor ( n32127 , n22094 , n32126 );
nor ( n32128 , n32125 , n32127 );
not ( n32129 , n32128 );
not ( n32130 , n32129 );
or ( n32131 , n32122 , n32130 );
and ( n32132 , n381909 , RI15b406e0_63);
nor ( n32133 , n22175 , n22199 );
and ( n32134 , n22168 , n32133 );
not ( n32135 , n22168 );
not ( n32136 , n20637 );
not ( n32137 , n22175 );
or ( n32138 , n32136 , n32137 );
nand ( n32139 , n32138 , n22094 );
and ( n32140 , n32135 , n32139 );
nor ( n32141 , n32134 , n32140 );
or ( n32142 , n32141 , n22213 );
not ( n32143 , n22287 );
nor ( n32144 , n32143 , n22268 );
and ( n32145 , n32144 , RI15b658c8_1330);
not ( n32146 , n32144 );
and ( n32147 , n32146 , n379836 );
or ( n32148 , n32145 , n32147 );
or ( n32149 , n32148 , n22296 );
or ( n32150 , n20507 , n22298 );
or ( n32151 , n22228 , n32150 );
nand ( n32152 , n32142 , n32149 , n32151 );
nor ( n32153 , n32132 , n32152 );
nand ( n32154 , n32131 , n32153 );
buf ( n32155 , n32154 );
buf ( n32156 , n382069 );
buf ( n32157 , n381707 );
buf ( n32158 , n380203 );
buf ( n32159 , n385197 );
buf ( n32160 , RI15b3ea48_2);
buf ( n32161 , n32160 );
and ( n32162 , n22142 , n22147 );
buf ( n32163 , n20427 );
buf ( n32164 , n32163 );
nand ( n32165 , n32162 , n32164 );
or ( n32166 , n380968 , n32165 );
not ( n32167 , n22206 );
nor ( n32168 , n22204 , n32167 );
buf ( n32169 , n22210 );
and ( n32170 , n32168 , n32169 );
and ( n32171 , n380986 , n32170 );
not ( n32172 , n32170 );
and ( n32173 , n32165 , n32172 , n19912 );
nor ( n32174 , n32173 , n22217 );
nand ( n32175 , n22109 , n22115 );
nor ( n32176 , n32175 , n22133 );
or ( n32177 , n32174 , n32176 );
nand ( n32178 , n32177 , n20623 );
or ( n32179 , n380923 , n20417 );
buf ( n32180 , n22226 );
or ( n32181 , n32179 , n32180 );
and ( n32182 , n32178 , n32181 );
nor ( n32183 , n32182 , n22236 );
or ( n32184 , n32183 , n385468 );
not ( n32185 , n32181 );
nor ( n32186 , n32176 , n32185 );
or ( n32187 , n32174 , n32186 );
or ( n32188 , n380994 , n32187 );
or ( n32189 , n32181 , n380996 );
nand ( n32190 , n32184 , n32188 , n32189 );
nor ( n32191 , n32171 , n32190 );
nand ( n32192 , n32166 , n32191 );
buf ( n32193 , n32192 );
buf ( n32194 , n22655 );
not ( n32195 , RI15b4a370_397);
or ( n32196 , n30907 , n32195 );
and ( n32197 , n20637 , n32195 );
or ( n32198 , n32195 , RI15b4a2f8_396);
nor ( n32199 , n19676 , RI15b4a370_397);
not ( n32200 , n32199 );
nand ( n32201 , n32198 , n32200 );
and ( n32202 , n22217 , n32201 );
not ( n32203 , n386306 );
not ( n32204 , n32203 );
nand ( n32205 , n386101 , n386116 );
not ( n32206 , n32205 );
and ( n32207 , n32204 , n32206 );
and ( n32208 , n32203 , n32205 );
nor ( n32209 , n32207 , n32208 );
or ( n32210 , n386499 , n32209 );
and ( n32211 , n385747 , n385645 );
not ( n32212 , n385747 );
and ( n32213 , n32212 , n385751 );
nor ( n32214 , n32211 , n32213 );
buf ( n32215 , n385750 );
and ( n32216 , n32214 , n32215 );
nor ( n32217 , n32214 , n32215 );
nor ( n32218 , n32216 , n32217 );
or ( n32219 , n386013 , n32218 );
not ( n32220 , n386259 );
not ( n32221 , n32205 );
buf ( n32222 , n386113 );
not ( n32223 , n32222 );
or ( n32224 , n32221 , n32223 );
or ( n32225 , n32222 , n32205 );
nand ( n32226 , n32224 , n32225 );
and ( n32227 , n32220 , n32226 );
and ( n32228 , n22394 , RI15b4b270_429);
nor ( n32229 , n32227 , n32228 );
nand ( n32230 , n32210 , n32219 , n32229 );
nor ( n32231 , n32197 , n32202 , n32230 );
nand ( n32232 , n32196 , n32231 );
buf ( n32233 , n32232 );
buf ( n32234 , n384700 );
buf ( n32235 , n382052 );
not ( n32236 , RI15b53538_708);
nand ( n32237 , n383683 , n381012 );
not ( n32238 , n32237 );
nor ( n32239 , RI15b5d768_1054 , RI15b5d7e0_1055 , RI15b5d858_1056 , RI15b5d8d0_1057);
not ( n32240 , RI15b5e758_1088);
not ( n32241 , RI15b5e848_1090);
nor ( n32242 , n32240 , n32241 , RI15b5e7d0_1089 , RI15b5e8c0_1091);
nand ( n32243 , n380484 , n32239 , n32242 );
and ( n32244 , n32238 , n32243 );
not ( n32245 , n32244 );
or ( n32246 , n32236 , n32245 );
and ( n32247 , n32237 , n32243 );
and ( n32248 , n32247 , RI15b64b30_1301);
not ( n32249 , n32243 );
and ( n32250 , n32249 , RI15b5f9a0_1127);
nor ( n32251 , n32248 , n32250 );
nand ( n32252 , n32246 , n32251 );
buf ( n32253 , n32252 );
buf ( n32254 , n380906 );
buf ( n32255 , RI15b3e9d0_1);
buf ( n32256 , n32255 );
buf ( n32257 , n382052 );
buf ( n32258 , n22655 );
not ( n32259 , n384960 );
or ( n32260 , n32259 , n32165 );
and ( n32261 , n384983 , n32170 );
not ( n32262 , RI15b43638_164);
or ( n32263 , n32183 , n32262 );
or ( n32264 , n22022 , n32187 );
or ( n32265 , n32181 , n384988 );
nand ( n32266 , n32263 , n32264 , n32265 );
nor ( n32267 , n32261 , n32266 );
nand ( n32268 , n32260 , n32267 );
buf ( n32269 , n32268 );
buf ( n32270 , n385197 );
buf ( n32271 , RI15b3ea48_2);
buf ( n32272 , n32271 );
buf ( n32273 , n22406 );
not ( n32274 , n384921 );
buf ( n32275 , n32274 );
not ( n32276 , n32275 );
not ( n32277 , RI15b615c0_1187);
nand ( n32278 , n383579 , n383584 );
nor ( n32279 , n32278 , RI15b613e0_1183);
not ( n32280 , RI15b61458_1184);
not ( n32281 , RI15b614d0_1185);
not ( n32282 , RI15b61548_1186);
and ( n32283 , n32279 , n32280 , n32281 , n32282 );
not ( n32284 , n32283 );
nand ( n32285 , n32284 , RI15b61bd8_1200);
not ( n32286 , n32285 );
or ( n32287 , n32277 , n32286 );
or ( n32288 , n32285 , RI15b615c0_1187);
nand ( n32289 , n32287 , n32288 );
not ( n32290 , n32281 );
buf ( n32291 , n32279 );
nand ( n32292 , n32291 , n32280 );
not ( n32293 , n32292 );
not ( n32294 , n32293 );
or ( n32295 , n32290 , n32294 );
nand ( n32296 , n32295 , RI15b61bd8_1200);
not ( n32297 , n32296 );
not ( n32298 , RI15b61548_1186);
and ( n32299 , n32297 , n32298 );
and ( n32300 , n32296 , RI15b61548_1186);
nor ( n32301 , n32299 , n32300 );
nand ( n32302 , n32292 , RI15b61bd8_1200);
and ( n32303 , n32302 , RI15b614d0_1185);
not ( n32304 , n32302 );
and ( n32305 , n32304 , n32281 );
nor ( n32306 , n32303 , n32305 );
nand ( n32307 , n32301 , n32306 );
nor ( n32308 , n32289 , n32307 );
not ( n32309 , RI15b615c0_1187);
and ( n32310 , n32283 , n32309 );
not ( n32311 , n32310 );
nand ( n32312 , n32311 , RI15b61bd8_1200);
not ( n32313 , n32312 );
not ( n32314 , RI15b61638_1188);
and ( n32315 , n32313 , n32314 );
and ( n32316 , n32312 , RI15b61638_1188);
nor ( n32317 , n32315 , n32316 );
nand ( n32318 , n32308 , n32317 );
not ( n32319 , RI15b616b0_1189);
not ( n32320 , RI15b61638_1188);
and ( n32321 , n32310 , n32320 );
not ( n32322 , n32321 );
nand ( n32323 , n32322 , RI15b61bd8_1200);
not ( n32324 , n32323 );
or ( n32325 , n32319 , n32324 );
or ( n32326 , n32323 , RI15b616b0_1189);
nand ( n32327 , n32325 , n32326 );
nor ( n32328 , n32318 , n32327 );
not ( n32329 , RI15b616b0_1189);
nand ( n32330 , n32321 , n32329 );
buf ( n32331 , n32330 );
nand ( n32332 , n32331 , RI15b61bd8_1200);
not ( n32333 , n32332 );
not ( n32334 , RI15b61728_1190);
and ( n32335 , n32333 , n32334 );
and ( n32336 , n32332 , RI15b61728_1190);
nor ( n32337 , n32335 , n32336 );
and ( n32338 , n32328 , n32337 );
buf ( n32339 , n32338 );
not ( n32340 , n32339 );
or ( n32341 , n32276 , n32340 );
not ( n32342 , n384926 );
not ( n32343 , n32342 );
nand ( n32344 , n32341 , n32343 );
nor ( n32345 , n32330 , RI15b61728_1190);
not ( n32346 , n32345 );
nand ( n32347 , n32346 , RI15b61bd8_1200);
not ( n32348 , n32347 );
not ( n32349 , RI15b617a0_1191);
and ( n32350 , n32348 , n32349 );
and ( n32351 , n32347 , RI15b617a0_1191);
nor ( n32352 , n32350 , n32351 );
not ( n32353 , n32352 );
nand ( n32354 , n32344 , n32353 );
nor ( n32355 , n32339 , n32353 );
nand ( n32356 , n32355 , n384934 );
nand ( n32357 , n384918 , RI15b5ec08_1098);
nand ( n32358 , n384906 , n381548 );
nand ( n32359 , n32354 , n32356 , n32357 , n32358 );
buf ( n32360 , n32359 );
buf ( n32361 , n22005 );
or ( n32362 , n385163 , n20672 );
not ( n32363 , n21573 );
and ( n32364 , n385174 , n32363 );
nor ( n32365 , n379984 , n18181 );
nor ( n32366 , n385168 , n32365 );
buf ( n32367 , n32366 );
nor ( n32368 , n32367 , n18078 );
and ( n32369 , n32368 , n21237 );
and ( n32370 , n385177 , n21463 );
nor ( n32371 , n32364 , n32369 , n32370 );
nand ( n32372 , n32362 , n22701 , n32371 );
buf ( n32373 , n32372 );
not ( n32374 , RI15b5c7f0_1021);
not ( n32375 , n31770 );
or ( n32376 , n32374 , n32375 );
not ( n32377 , n31781 );
buf ( n32378 , n32377 );
not ( n32379 , n32378 );
and ( n32380 , n32379 , n380820 );
not ( n32381 , n31757 );
nand ( n32382 , n32381 , n19545 , n22418 );
not ( n32383 , n31086 );
nand ( n32384 , n32383 , n383588 );
and ( n32385 , n32382 , n32384 , n19556 );
nor ( n32386 , n32385 , n19200 );
and ( n32387 , n32386 , n380808 );
and ( n32388 , n31778 , n380831 );
nor ( n32389 , n32380 , n32387 , n32388 );
nand ( n32390 , n32376 , n32389 );
nor ( n32391 , n380842 , n32390 );
not ( n32392 , n32391 );
buf ( n32393 , n32392 );
buf ( n32394 , n22404 );
buf ( n32395 , n380903 );
not ( n32396 , RI15b526b0_677);
buf ( n32397 , n381484 );
not ( n32398 , n32397 );
or ( n32399 , n32396 , n32398 );
not ( n32400 , n383112 );
not ( n32401 , n381422 );
or ( n32402 , n32400 , n32401 );
nand ( n32403 , n32402 , n381450 );
not ( n32404 , n383120 );
and ( n32405 , n32403 , n32404 );
not ( n32406 , n32400 );
nor ( n32407 , n32406 , n32404 );
and ( n32408 , n32407 , n381461 );
not ( n32409 , n386729 );
nor ( n32410 , n381400 , n32409 );
nor ( n32411 , n32405 , n32408 , n32410 );
nand ( n32412 , n32399 , n32411 );
buf ( n32413 , n32412 );
not ( n32414 , n386590 );
not ( n32415 , n381589 );
or ( n32416 , n32414 , n32415 );
and ( n32417 , n381596 , n386603 );
or ( n32418 , n386612 , n18720 );
buf ( n32419 , n381614 );
not ( n32420 , n32419 );
or ( n32421 , n32420 , n386624 );
or ( n32422 , n386610 , n381621 );
nand ( n32423 , n32418 , n32421 , n32422 );
nor ( n32424 , n32417 , n32423 );
nand ( n32425 , n32416 , n32424 );
buf ( n32426 , n32425 );
buf ( n32427 , n386762 );
buf ( n32428 , n380942 );
or ( n32429 , n381405 , n382692 );
not ( n32430 , n32429 );
buf ( n32431 , n381387 );
buf ( n32432 , n32431 );
or ( n32433 , n32430 , n32432 );
not ( n32434 , n381392 );
nand ( n32435 , n381417 , n32434 );
and ( n32436 , n386637 , RI15b54e10_761);
not ( n32437 , n386670 );
and ( n32438 , n381694 , n32437 );
buf ( n32439 , n382626 );
not ( n32440 , RI15b54e10_761);
not ( n32441 , n382645 );
or ( n32442 , n32440 , n32441 );
or ( n32443 , n382645 , RI15b54e10_761);
nand ( n32444 , n32442 , n32443 );
and ( n32445 , n32439 , n32444 );
nor ( n32446 , n32436 , n32438 , n32445 );
and ( n32447 , n32435 , n32446 );
nand ( n32448 , n32433 , n32447 );
buf ( n32449 , n32448 );
buf ( n32450 , n383498 );
buf ( n32451 , n384218 );
not ( n32452 , n31178 );
or ( n32453 , n32430 , n32452 );
nand ( n32454 , n381417 , n381369 );
and ( n32455 , n386637 , RI15b549d8_752);
buf ( n32456 , n21413 );
and ( n32457 , n382885 , n32456 );
buf ( n32458 , n382625 );
not ( n32459 , n32458 );
not ( n32460 , RI15b549d8_752);
not ( n32461 , n382632 );
or ( n32462 , n32460 , n32461 );
or ( n32463 , n382632 , RI15b549d8_752);
nand ( n32464 , n32462 , n32463 );
and ( n32465 , n32459 , n32464 );
nor ( n32466 , n32455 , n32457 , n32465 );
and ( n32467 , n32454 , n32466 );
nand ( n32468 , n32453 , n32467 );
buf ( n32469 , n32468 );
buf ( n32470 , n32271 );
not ( n32471 , n32064 );
not ( n32472 , n381507 );
or ( n32473 , n32471 , n32472 );
and ( n32474 , n381524 , n32070 );
not ( n32475 , RI15b5a4c8_946);
or ( n32476 , n32081 , n32475 );
buf ( n32477 , n381549 );
not ( n32478 , n32477 );
or ( n32479 , n32478 , n32086 );
or ( n32480 , n32079 , n381560 );
nand ( n32481 , n32476 , n32479 , n32480 );
nor ( n32482 , n32474 , n32481 );
nand ( n32483 , n32473 , n32482 );
buf ( n32484 , n32483 );
buf ( n32485 , n381566 );
not ( n32486 , n382001 );
not ( n32487 , n381993 );
or ( n32488 , n32486 , n32487 );
or ( n32489 , n381993 , n382001 );
nand ( n32490 , n32488 , n32489 );
and ( n32491 , n379822 , n32490 );
nor ( n32492 , n379834 , n381988 );
nor ( n32493 , n32491 , n32492 );
nand ( n32494 , n379832 , RI15b46ba8_278);
nand ( n32495 , n379825 , RI15b488b8_340);
nand ( n32496 , n32493 , n32494 , n32495 );
buf ( n32497 , n32496 );
buf ( n32498 , n382049 );
buf ( n32499 , n18226 );
buf ( n32500 , n386563 );
buf ( n32501 , n380940 );
not ( n32502 , n20525 );
buf ( n32503 , n19847 );
not ( n32504 , n19855 );
and ( n32505 , n32502 , n32503 , n32504 );
buf ( n32506 , n19984 );
and ( n32507 , n32506 , n31806 );
nor ( n32508 , n32507 , n20521 );
or ( n32509 , n32508 , n19985 );
not ( n32510 , n32506 );
not ( n32511 , n20529 );
and ( n32512 , n32510 , n32511 , n19985 );
or ( n32513 , n22353 , n20553 , RI15b4bae0_447);
or ( n32514 , n20653 , n19851 );
nand ( n32515 , n32513 , n32514 );
nor ( n32516 , n32512 , n32515 );
nand ( n32517 , n32509 , n32516 );
nor ( n32518 , n32505 , n32517 );
or ( n32519 , n32503 , n19918 );
nand ( n32520 , n32519 , n19938 );
nand ( n32521 , n32520 , n19855 );
not ( n32522 , n20639 );
not ( n32523 , n20567 );
and ( n32524 , n32523 , n20553 );
not ( n32525 , n20613 );
nor ( n32526 , n32524 , n32525 );
not ( n32527 , n32526 );
or ( n32528 , n32522 , n32527 );
nand ( n32529 , n32528 , RI15b4bae0_447);
nand ( n32530 , n32518 , n32521 , n32529 );
buf ( n32531 , n32530 );
buf ( n32532 , n22738 );
buf ( n32533 , n18226 );
not ( n32534 , n384348 );
not ( n32535 , n32534 );
not ( n32536 , n384295 );
nor ( n32537 , n387129 , n32536 );
buf ( n32538 , n384303 );
and ( n32539 , n32537 , n32538 );
nand ( n32540 , n32539 , n384328 );
nor ( n32541 , n32540 , n384284 );
nand ( n32542 , n32541 , n384267 );
buf ( n32543 , n32542 );
not ( n32544 , n32543 );
or ( n32545 , n32535 , n32544 );
nor ( n32546 , n32542 , n32534 );
not ( n32547 , n32546 );
nand ( n32548 , n32545 , n32547 );
buf ( n32549 , n31921 );
and ( n32550 , n32548 , n32549 );
not ( n32551 , n384570 );
nor ( n32552 , n384526 , n384558 );
nand ( n32553 , n32552 , n384550 );
nor ( n32554 , n32553 , n384565 );
nand ( n32555 , n32551 , n32554 );
not ( n32556 , n384583 );
nor ( n32557 , n32555 , n32556 );
buf ( n32558 , n32557 );
not ( n32559 , n32558 );
not ( n32560 , n384595 );
not ( n32561 , n32560 );
and ( n32562 , n32559 , n32561 );
and ( n32563 , n32558 , n32560 );
nor ( n32564 , n32562 , n32563 );
or ( n32565 , n32564 , n31958 );
not ( n32566 , n384473 );
buf ( n32567 , n384447 );
nand ( n32568 , n32567 , n384470 );
not ( n32569 , n32568 );
or ( n32570 , n32566 , n32569 );
or ( n32571 , n32568 , n384473 );
nand ( n32572 , n32570 , n32571 );
and ( n32573 , n32572 , n384493 );
and ( n32574 , n19513 , RI15b642c0_1283);
nor ( n32575 , n32573 , n32574 );
nand ( n32576 , n32565 , n32575 );
nor ( n32577 , n32550 , n32576 );
not ( n32578 , n383438 );
not ( n32579 , n381572 );
or ( n32580 , n32578 , n32579 );
buf ( n32581 , n384637 );
buf ( n32582 , n32581 );
nand ( n32583 , n32580 , n32582 );
and ( n32584 , n32583 , RI15b633c0_1251);
or ( n32585 , n384652 , n383438 , RI15b633c0_1251);
not ( n32586 , n386885 );
or ( n32587 , n32586 , n22775 );
nand ( n32588 , n32585 , n32587 );
nor ( n32589 , n32584 , n32588 );
nand ( n32590 , n32577 , n32589 );
buf ( n32591 , n32590 );
buf ( n32592 , n32160 );
buf ( n32593 , n382065 );
not ( n32594 , n19918 );
not ( n32595 , n32594 );
not ( n32596 , n19823 );
not ( n32597 , n32596 );
or ( n32598 , n32595 , n32597 );
nand ( n32599 , n32598 , n19938 );
and ( n32600 , n32599 , n19830 );
or ( n32601 , n22355 , n20549 , RI15b4b900_443);
not ( n32602 , n19978 );
or ( n32603 , n22362 , n32602 , RI15b49b00_379);
nand ( n32604 , n32601 , n32603 );
nor ( n32605 , n32600 , n32604 );
not ( n32606 , n19830 );
not ( n32607 , n32596 );
nand ( n32608 , n32606 , n383353 , n32607 );
and ( n32609 , n20565 , n20549 );
nor ( n32610 , n32609 , n22372 );
or ( n32611 , n32610 , n382114 );
and ( n32612 , n32602 , n22377 );
nor ( n32613 , n32612 , n22383 );
not ( n32614 , RI15b49b00_379);
or ( n32615 , n32613 , n32614 );
nand ( n32616 , n32611 , n32615 );
nand ( n32617 , n32616 , n20501 );
and ( n32618 , n22388 , RI15b4b900_443);
buf ( n32619 , n20653 );
not ( n32620 , n32619 );
buf ( n32621 , n32620 );
and ( n32622 , n32621 , RI15b4aa00_411);
nor ( n32623 , n32618 , n32622 , n22398 );
nand ( n32624 , n32605 , n32608 , n32617 , n32623 );
buf ( n32625 , n32624 );
and ( n32626 , n32557 , n384595 );
nand ( n32627 , n32626 , n384592 );
not ( n32628 , n384543 );
nor ( n32629 , n32627 , n32628 );
nand ( n32630 , n32629 , n384537 );
and ( n32631 , n32630 , n384530 );
not ( n32632 , n32630 );
not ( n32633 , n384530 );
and ( n32634 , n32632 , n32633 );
nor ( n32635 , n32631 , n32634 );
not ( n32636 , n31960 );
nor ( n32637 , n32635 , n32636 );
not ( n32638 , n384465 );
not ( n32639 , n32638 );
not ( n32640 , n384473 );
nor ( n32641 , n32568 , n32640 );
nand ( n32642 , n32639 , n32641 );
not ( n32643 , n384455 );
nor ( n32644 , n32642 , n32643 );
nand ( n32645 , n32644 , n384461 );
and ( n32646 , n32645 , n384451 );
not ( n32647 , n32645 );
not ( n32648 , n384451 );
and ( n32649 , n32647 , n32648 );
nor ( n32650 , n32646 , n32649 );
not ( n32651 , n31884 );
nor ( n32652 , n32650 , n32651 );
not ( n32653 , n384371 );
and ( n32654 , n32653 , n384259 );
not ( n32655 , n384372 );
nor ( n32656 , n32654 , n32655 );
or ( n32657 , n32656 , n31922 );
or ( n32658 , n19512 , n379708 );
nand ( n32659 , n32657 , n32658 );
nor ( n32660 , n32637 , n32652 , n32659 );
not ( n32661 , n31965 );
or ( n32662 , n32661 , RI15b63528_1254);
nand ( n32663 , n32662 , n384642 );
and ( n32664 , n32663 , RI15b635a0_1255);
and ( n32665 , n384655 , n386781 , RI15b63528_1254);
and ( n32666 , n386785 , n19630 );
nor ( n32667 , n32665 , n32666 );
not ( n32668 , n32667 );
nor ( n32669 , n32664 , n32668 );
nand ( n32670 , n32660 , n32669 );
buf ( n32671 , n32670 );
buf ( n32672 , RI15b3e9d0_1);
buf ( n32673 , n32672 );
buf ( n32674 , n385195 );
buf ( n32675 , n381021 );
buf ( n32676 , RI15b3e9d0_1);
buf ( n32677 , n32676 );
buf ( n32678 , n379403 );
not ( n32679 , n380230 );
and ( n32680 , n32679 , n380234 );
not ( n32681 , n32680 );
or ( n32682 , n383180 , n32681 );
nand ( n32683 , n382981 , n380737 );
not ( n32684 , n380750 );
and ( n32685 , n32683 , n32681 , n32684 );
nor ( n32686 , n32685 , n19630 );
nor ( n32687 , n382988 , n380759 );
or ( n32688 , n32686 , n32687 );
nand ( n32689 , n32688 , n19595 );
or ( n32690 , n382992 , n380767 );
nand ( n32691 , n32689 , n32690 );
and ( n32692 , n32691 , n380775 );
not ( n32693 , n32692 );
and ( n32694 , n32693 , RI15b5a5b8_948);
or ( n32695 , n383184 , n32683 );
not ( n32696 , n383188 );
not ( n32697 , n32690 );
nor ( n32698 , n32687 , n32697 );
or ( n32699 , n32686 , n32698 );
or ( n32700 , n32696 , n32699 );
or ( n32701 , n32690 , n383192 );
nand ( n32702 , n32695 , n32700 , n32701 );
nor ( n32703 , n32694 , n32702 );
nand ( n32704 , n32682 , n32703 );
buf ( n32705 , n32704 );
buf ( n32706 , n385195 );
or ( n32707 , n382679 , n32100 );
or ( n32708 , n21603 , n382886 );
buf ( n32709 , n381190 );
buf ( n32710 , n32709 );
not ( n32711 , n32710 );
and ( n32712 , n382677 , n18182 , n32711 );
and ( n32713 , n382626 , n32100 );
nor ( n32714 , n32712 , n32713 );
nand ( n32715 , n32707 , n32708 , n32714 );
buf ( n32716 , n32715 );
buf ( n32717 , n379403 );
buf ( n32718 , n19651 );
buf ( n32719 , n22740 );
buf ( n32720 , n386760 );
not ( n32721 , RI15b53f88_730);
not ( n32722 , n32244 );
or ( n32723 , n32721 , n32722 );
and ( n32724 , n32247 , RI15b65580_1323);
and ( n32725 , n32249 , RI15b603f0_1149);
nor ( n32726 , n32724 , n32725 );
nand ( n32727 , n32723 , n32726 );
buf ( n32728 , n32727 );
buf ( n32729 , n20035 );
not ( n32730 , n32729 );
and ( n32731 , n32730 , RI15b44a60_207);
not ( n32732 , RI15b44b50_209);
or ( n32733 , n32732 , RI15b44a60_207);
nand ( n32734 , n32733 , n385332 );
nor ( n32735 , n32731 , n32734 );
not ( n32736 , n32735 );
not ( n32737 , RI15b44ad8_208);
and ( n32738 , RI15b44a60_207 , n32737 );
not ( n32739 , RI15b44a60_207);
and ( n32740 , n32739 , RI15b44ad8_208);
nor ( n32741 , n32738 , n32740 );
and ( n32742 , n381046 , n32736 , n32741 );
not ( n32743 , n32742 );
buf ( n32744 , n385990 );
buf ( n32745 , n32744 );
not ( n32746 , n32745 );
nor ( n32747 , n32743 , n32746 );
and ( n32748 , n32747 , RI15b42a08_138);
not ( n32749 , n381048 );
not ( n32750 , n32749 );
nor ( n32751 , n32736 , n32741 );
buf ( n32752 , n386000 );
and ( n32753 , n32751 , n32752 );
and ( n32754 , n32753 , RI15b41748_98);
and ( n32755 , n32751 , n32744 );
and ( n32756 , n32755 , RI15b41b08_106);
nor ( n32757 , n32754 , n32756 );
not ( n32758 , n385993 );
and ( n32759 , n32751 , n32758 );
and ( n32760 , n32759 , RI15b40fc8_82);
buf ( n32761 , n386003 );
and ( n32762 , n32751 , n32761 );
and ( n32763 , n32762 , RI15b41388_90);
nor ( n32764 , n32760 , n32763 );
nor ( n32765 , n32735 , n32741 );
and ( n32766 , n32765 , n32752 );
and ( n32767 , n32766 , RI15b43548_162);
and ( n32768 , n32765 , n32761 );
and ( n32769 , n32768 , RI15b43188_154);
nor ( n32770 , n32767 , n32769 );
and ( n32771 , n32765 , n32744 );
and ( n32772 , n32771 , RI15b43908_170);
and ( n32773 , n32765 , n32758 );
and ( n32774 , n32773 , RI15b42dc8_146);
nor ( n32775 , n32772 , n32774 );
nand ( n32776 , n32757 , n32764 , n32770 , n32775 );
and ( n32777 , n32750 , n32776 );
nand ( n32778 , n381046 , n32735 , n32741 );
buf ( n32779 , n32761 );
not ( n32780 , n32779 );
nor ( n32781 , n32778 , n32780 );
and ( n32782 , n32781 , RI15b40488_58);
nor ( n32783 , n32748 , n32777 , n32782 );
buf ( n32784 , n32752 );
and ( n32785 , n32742 , n32784 );
and ( n32786 , n32785 , RI15b42648_130);
and ( n32787 , n32742 , n32779 );
and ( n32788 , n32787 , RI15b42288_122);
nor ( n32789 , n32786 , n32788 );
not ( n32790 , n32778 );
buf ( n32791 , n32758 );
and ( n32792 , n32790 , n32791 );
and ( n32793 , n32792 , RI15b400c8_50);
and ( n32794 , n32742 , n32791 );
and ( n32795 , n32794 , RI15b41ec8_114);
nor ( n32796 , n32793 , n32795 );
and ( n32797 , n32790 , n32784 );
and ( n32798 , n32797 , RI15b40848_66);
not ( n32799 , n32746 );
and ( n32800 , n32790 , n32799 );
and ( n32801 , n32800 , RI15b40c08_74);
nor ( n32802 , n32798 , n32801 );
nand ( n32803 , n32783 , n32789 , n32796 , n32802 );
not ( n32804 , n32803 );
buf ( n32805 , n381039 );
not ( n32806 , n32805 );
not ( n32807 , n32806 );
or ( n32808 , n32804 , n32807 );
and ( n32809 , n381055 , RI15b49920_375);
not ( n32810 , RI15b49920_375);
nand ( n32811 , n381066 , RI15b494e8_366);
not ( n32812 , RI15b49560_367);
nor ( n32813 , n32811 , n32812 );
and ( n32814 , n32813 , RI15b495d8_368);
nand ( n32815 , n32814 , RI15b49650_369);
not ( n32816 , RI15b496c8_370);
nor ( n32817 , n32815 , n32816 );
nand ( n32818 , n32817 , RI15b49740_371);
not ( n32819 , n32818 );
nand ( n32820 , n32819 , RI15b497b8_372);
not ( n32821 , RI15b49830_373);
nor ( n32822 , n32820 , n32821 );
and ( n32823 , n32822 , RI15b498a8_374);
not ( n32824 , n32823 );
not ( n32825 , n32824 );
or ( n32826 , n32810 , n32825 );
or ( n32827 , n32824 , RI15b49920_375);
nand ( n32828 , n32826 , n32827 );
and ( n32829 , n381076 , n32828 );
nor ( n32830 , n32809 , n32829 );
nand ( n32831 , n32808 , n32830 );
buf ( n32832 , n32831 );
buf ( n32833 , n32676 );
buf ( n32834 , n22404 );
not ( n32835 , n382439 );
nand ( n32836 , n382489 , n382457 , n382465 , n32835 );
nor ( n32837 , n32018 , n32836 );
buf ( n32838 , n32837 );
buf ( n32839 , n32003 );
not ( n32840 , n32839 );
not ( n32841 , n382375 );
or ( n32842 , n32840 , n32841 );
not ( n32843 , RI15b4c008_458);
nand ( n32844 , n32843 , RI15b4b978_444);
nand ( n32845 , n32842 , n32844 );
not ( n32846 , n32839 );
not ( n32847 , n382366 );
or ( n32848 , n32846 , n32847 );
not ( n32849 , RI15b4c008_458);
nand ( n32850 , n32849 , RI15b4b900_443);
nand ( n32851 , n32848 , n32850 );
nor ( n32852 , n32845 , n32851 );
not ( n32853 , n382471 );
or ( n32854 , n32853 , n382343 );
nand ( n32855 , n32854 , n382345 );
not ( n32856 , n382446 );
nor ( n32857 , n32855 , n32856 );
nand ( n32858 , n32852 , n32857 );
buf ( n32859 , n382412 );
or ( n32860 , n382472 , n32859 );
not ( n32861 , RI15b4c008_458);
nand ( n32862 , n32861 , RI15b4bae0_447);
nand ( n32863 , n32860 , n32862 );
buf ( n32864 , n382403 );
or ( n32865 , n32840 , n32864 );
not ( n32866 , RI15b4c008_458);
nand ( n32867 , n32866 , RI15b4bb58_448);
nand ( n32868 , n32865 , n32867 );
nor ( n32869 , n32863 , n32868 );
not ( n32870 , n382420 );
or ( n32871 , n32853 , n32870 );
not ( n32872 , RI15b4c008_458);
nand ( n32873 , n32872 , RI15b4bbd0_449);
nand ( n32874 , n32871 , n32873 );
nor ( n32875 , n32874 , n32031 );
nand ( n32876 , n32869 , n32875 );
nor ( n32877 , n32858 , n32876 );
not ( n32878 , n382361 );
not ( n32879 , n32878 );
not ( n32880 , n382471 );
or ( n32881 , n32879 , n32880 );
not ( n32882 , RI15b4c008_458);
nand ( n32883 , n32882 , RI15b4b9f0_445);
nand ( n32884 , n32881 , n32883 );
not ( n32885 , n382389 );
not ( n32886 , n32885 );
not ( n32887 , n382471 );
or ( n32888 , n32886 , n32887 );
not ( n32889 , RI15b4c008_458);
nand ( n32890 , n32889 , RI15b4ba68_446);
nand ( n32891 , n32888 , n32890 );
nor ( n32892 , n32884 , n32891 );
not ( n32893 , n32045 );
not ( n32894 , n32003 );
or ( n32895 , n32893 , n32894 );
not ( n32896 , RI15b4c008_458);
nand ( n32897 , n32896 , RI15b4b810_441);
nand ( n32898 , n32895 , n32897 );
nor ( n32899 , n32898 , n31988 );
and ( n32900 , n32892 , n32899 , n382447 );
nand ( n32901 , n32838 , n32877 , n32900 );
not ( n32902 , n32901 );
not ( n32903 , n382473 );
buf ( n32904 , n382193 );
not ( n32905 , n32904 );
and ( n32906 , n32903 , n32905 );
not ( n32907 , RI15b4c008_458);
and ( n32908 , n32907 , RI15b4bcc0_451);
nor ( n32909 , n32906 , n32908 );
nor ( n32910 , n382473 , n382430 );
nor ( n32911 , n382126 , RI15b4c008_458);
nor ( n32912 , n32910 , n32911 );
nand ( n32913 , n32909 , n32912 );
not ( n32914 , n382473 );
buf ( n32915 , n382177 );
not ( n32916 , n32915 );
and ( n32917 , n32914 , n32916 );
not ( n32918 , n382195 );
nor ( n32919 , n32917 , n32918 );
buf ( n32920 , n382498 );
nand ( n32921 , n32919 , n32920 );
nor ( n32922 , n32913 , n32921 );
nand ( n32923 , n32902 , n32922 );
buf ( n32924 , n32035 );
not ( n32925 , n32924 );
nand ( n32926 , n32923 , n32925 );
not ( n32927 , n32926 );
not ( n32928 , n32036 );
not ( n32929 , n32928 );
not ( n32930 , n32929 );
not ( n32931 , n382473 );
buf ( n32932 , n382503 );
not ( n32933 , n32932 );
and ( n32934 , n32931 , n32933 );
not ( n32935 , RI15b4c008_458);
and ( n32936 , n32935 , RI15b4bea0_455);
nor ( n32937 , n32934 , n32936 );
not ( n32938 , n32937 );
not ( n32939 , n32938 );
or ( n32940 , n32930 , n32939 );
not ( n32941 , n32035 );
or ( n32942 , n382143 , RI15b4c008_458);
buf ( n32943 , n382500 );
nand ( n32944 , n32942 , n32943 );
nand ( n32945 , n32941 , n32944 );
nand ( n32946 , n32940 , n32945 );
nor ( n32947 , n32927 , n32946 );
or ( n32948 , n382473 , n382505 );
or ( n32949 , n380886 , RI15b4c008_458);
nand ( n32950 , n32948 , n32949 );
or ( n32951 , n32947 , n32950 );
not ( n32952 , n32937 );
not ( n32953 , n32944 );
nand ( n32954 , n32953 , n382080 );
nor ( n32955 , n32923 , n32954 );
not ( n32956 , n32955 );
or ( n32957 , n32952 , n32956 );
buf ( n32958 , n32024 );
not ( n32959 , n32958 );
nand ( n32960 , n32957 , n32959 );
nand ( n32961 , n32960 , n32950 );
not ( n32962 , n382512 );
buf ( n32963 , n32962 );
not ( n32964 , n32963 );
not ( n32965 , n32964 );
not ( n32966 , n382506 );
buf ( n32967 , n382492 );
not ( n32968 , n32967 );
and ( n32969 , n32966 , n32968 );
and ( n32970 , n382506 , n32967 );
nor ( n32971 , n32969 , n32970 );
and ( n32972 , n32965 , n32971 );
and ( n32973 , n382523 , RI15b4bf90_457);
buf ( n32974 , n382529 );
buf ( n32975 , n32974 );
and ( n32976 , n32975 , RI15b45d98_248);
nor ( n32977 , n32972 , n32973 , n32976 );
nand ( n32978 , n32951 , n32961 , n32977 );
buf ( n32979 , n32978 );
buf ( n32980 , n22009 );
buf ( n32981 , RI15b3ea48_2);
buf ( n32982 , n32981 );
buf ( n32983 , n381021 );
buf ( n32984 , n382073 );
buf ( n32985 , n380940 );
and ( n32986 , n18156 , RI15b4c080_459);
not ( n32987 , n32986 );
not ( n32988 , n17996 );
not ( n32989 , RI15b50f40_627);
not ( n32990 , n18003 );
or ( n32991 , n32989 , n32990 );
nand ( n32992 , n32991 , n17587 );
not ( n32993 , n32992 );
or ( n32994 , n32988 , n32993 );
nand ( n32995 , n32994 , n18156 );
nand ( n32996 , n32987 , n32995 );
not ( n32997 , n32996 );
nand ( n32998 , n32997 , n383163 );
or ( n32999 , n383900 , n32998 );
nand ( n33000 , n32999 , RI15b4c0f8_460);
and ( n33001 , n32996 , RI15b4c080_459);
and ( n33002 , n383915 , n18057 );
nor ( n33003 , n33001 , n33002 );
nand ( n33004 , n33000 , n33003 );
buf ( n33005 , n33004 );
buf ( n33006 , n380940 );
buf ( n33007 , n386563 );
not ( n33008 , RI15b62da8_1238);
not ( n33009 , n19608 );
or ( n33010 , n33008 , n33009 );
not ( n33011 , n386805 );
and ( n33012 , n33011 , n386809 );
not ( n33013 , n33011 );
and ( n33014 , n33013 , RI15b62da8_1238);
nor ( n33015 , n33012 , n33014 );
and ( n33016 , n380237 , n33015 );
not ( n33017 , n19356 );
buf ( n33018 , n18744 );
not ( n33019 , n19309 );
not ( n33020 , n19322 );
not ( n33021 , n33020 );
not ( n33022 , n19343 );
or ( n33023 , n33021 , n33022 );
nand ( n33024 , n33023 , n19347 );
not ( n33025 , n33024 );
or ( n33026 , n33019 , n33025 );
nand ( n33027 , n33026 , n19352 );
and ( n33028 , n33018 , n33027 );
not ( n33029 , n33018 );
not ( n33030 , n19352 );
not ( n33031 , n33024 );
not ( n33032 , n33031 );
or ( n33033 , n33030 , n33032 );
nand ( n33034 , n33033 , n19309 );
and ( n33035 , n33029 , n33034 );
nor ( n33036 , n33028 , n33035 );
not ( n33037 , n33036 );
or ( n33038 , n33017 , n33037 );
or ( n33039 , n33036 , n19356 );
nand ( n33040 , n33038 , n33039 );
not ( n33041 , n19389 );
and ( n33042 , n33040 , n33041 );
and ( n33043 , n19513 , RI15b63ca8_1270);
nor ( n33044 , n33042 , n33043 );
not ( n33045 , n382561 );
not ( n33046 , n18688 );
and ( n33047 , n33045 , n33046 );
and ( n33048 , n382561 , n18688 );
nor ( n33049 , n33047 , n33048 );
buf ( n33050 , n33018 );
and ( n33051 , n33049 , n33050 );
not ( n33052 , n33049 );
not ( n33053 , n33050 );
and ( n33054 , n33052 , n33053 );
nor ( n33055 , n33051 , n33054 );
not ( n33056 , n19284 );
and ( n33057 , n33055 , n33056 );
not ( n33058 , n33018 );
not ( n33059 , n19462 );
not ( n33060 , n382579 );
or ( n33061 , n33059 , n33060 );
or ( n33062 , n382575 , n19470 );
nand ( n33063 , n33062 , n19444 );
nand ( n33064 , n33063 , n19450 );
nand ( n33065 , n33061 , n33064 );
not ( n33066 , n33065 );
or ( n33067 , n33058 , n33066 );
or ( n33068 , n33065 , n33050 );
nand ( n33069 , n33067 , n33068 );
and ( n33070 , n33069 , n22761 );
nor ( n33071 , n33057 , n33070 );
nand ( n33072 , n33044 , n33071 );
nor ( n33073 , n22775 , n386811 );
nor ( n33074 , n33016 , n33072 , n33073 );
nand ( n33075 , n33010 , n33074 );
buf ( n33076 , n33075 );
buf ( n33077 , n380203 );
buf ( n33078 , RI15b475f8_300);
or ( n33079 , n381907 , n380909 );
not ( n33080 , n380928 );
and ( n33081 , n33080 , RI15b41dd8_112);
or ( n33082 , n381917 , n380915 );
not ( n33083 , n380933 );
and ( n33084 , n33083 , n381923 );
and ( n33085 , n381926 , n380931 );
nor ( n33086 , n33084 , n33085 );
nand ( n33087 , n33082 , n33086 );
nor ( n33088 , n33081 , n33087 );
nand ( n33089 , n33079 , n33088 );
buf ( n33090 , n33089 );
buf ( n33091 , n382071 );
buf ( n33092 , n381006 );
buf ( n33093 , n380940 );
buf ( n33094 , n384218 );
buf ( n33095 , n22005 );
not ( n33096 , RI15b606c0_1155);
or ( n33097 , n31037 , n22435 );
nand ( n33098 , n33097 , n385188 );
not ( n33099 , n33098 );
or ( n33100 , n33096 , n33099 );
not ( n33101 , n22442 );
nand ( n33102 , n33101 , n31038 );
and ( n33103 , n33102 , RI15b3fab0_37);
not ( n33104 , n31044 );
nor ( n33105 , n33103 , n33104 );
nand ( n33106 , n33100 , n33105 );
buf ( n33107 , n33106 );
buf ( n33108 , n30992 );
buf ( n33109 , n383868 );
not ( n33110 , n383886 );
nand ( n33111 , n33109 , n33110 );
not ( n33112 , n33111 );
not ( n33113 , n33112 );
not ( n33114 , n384122 );
or ( n33115 , n33113 , n33114 );
nand ( n33116 , n385004 , n21337 );
not ( n33117 , n33116 );
and ( n33118 , n384164 , n33117 );
not ( n33119 , n385008 );
and ( n33120 , n33116 , n33111 , n33119 );
nor ( n33121 , n33120 , n21764 );
buf ( n33122 , n383894 );
nor ( n33123 , n385012 , n33122 );
or ( n33124 , n33121 , n33123 );
nand ( n33125 , n33124 , n18154 );
or ( n33126 , n385016 , n383865 );
nand ( n33127 , n33125 , n33126 );
and ( n33128 , n33127 , n383901 );
or ( n33129 , n33128 , n20902 );
buf ( n33130 , n384185 );
not ( n33131 , n33130 );
not ( n33132 , n33126 );
nor ( n33133 , n33123 , n33132 );
or ( n33134 , n33121 , n33133 );
or ( n33135 , n33131 , n33134 );
or ( n33136 , n33126 , n384193 );
nand ( n33137 , n33129 , n33135 , n33136 );
nor ( n33138 , n33118 , n33137 );
nand ( n33139 , n33115 , n33138 );
buf ( n33140 , n33139 );
buf ( n33141 , n31979 );
buf ( n33142 , n22343 );
buf ( n33143 , n386563 );
buf ( n33144 , n32676 );
not ( n33145 , n382285 );
or ( n33146 , n382093 , n33145 );
or ( n33147 , n33145 , n382091 );
nand ( n33148 , n33147 , RI15b4b360_431);
nand ( n33149 , n33146 , n33148 );
nand ( n33150 , n32962 , n33149 );
nand ( n33151 , n382447 , n382080 );
not ( n33152 , n33151 );
not ( n33153 , n382474 );
or ( n33154 , n33152 , n33153 );
nand ( n33155 , n33154 , n32856 );
nor ( n33156 , n32856 , n382447 );
nand ( n33157 , n382488 , n33156 );
and ( n33158 , n382523 , RI15b4b360_431);
buf ( n33159 , n382528 );
and ( n33160 , n33159 , RI15b45168_222);
nor ( n33161 , n33158 , n33160 );
nand ( n33162 , n33150 , n33155 , n33157 , n33161 );
buf ( n33163 , n33162 );
buf ( n33164 , n380906 );
not ( n33165 , n380909 );
not ( n33166 , n33165 );
buf ( n33167 , n384943 );
not ( n33168 , n33167 );
not ( n33169 , n33168 );
nor ( n33170 , n384950 , n380965 );
not ( n33171 , n33170 );
or ( n33172 , n33169 , n33171 );
nand ( n33173 , n33172 , n22097 );
not ( n33174 , n33173 );
not ( n33175 , n33174 );
or ( n33176 , n33166 , n33175 );
not ( n33177 , n22058 );
nand ( n33178 , n33177 , RI15b666d8_1360);
not ( n33179 , n33178 );
not ( n33180 , RI15b66318_1352);
and ( n33181 , n33179 , n33180 );
and ( n33182 , n33178 , RI15b66318_1352);
nor ( n33183 , n33181 , n33182 );
nand ( n33184 , n33183 , n22097 );
not ( n33185 , n33184 );
nor ( n33186 , n384972 , n384968 );
not ( n33187 , n33186 );
and ( n33188 , n33185 , n33187 );
not ( n33189 , n20637 );
not ( n33190 , n33186 );
or ( n33191 , n33189 , n33190 );
nand ( n33192 , n33191 , n22094 );
not ( n33193 , n33183 );
and ( n33194 , n33192 , n33193 );
nor ( n33195 , n33188 , n33194 );
not ( n33196 , n33195 );
and ( n33197 , n33196 , n380913 );
or ( n33198 , n380928 , n385345 );
or ( n33199 , n22241 , n380933 );
buf ( n33200 , n20591 );
nand ( n33201 , n33200 , n381925 );
or ( n33202 , n380926 , n33201 );
nand ( n33203 , n33198 , n33199 , n33202 );
nor ( n33204 , n33197 , n33203 );
nand ( n33205 , n33176 , n33204 );
buf ( n33206 , n33205 );
buf ( n33207 , n384203 );
buf ( n33208 , n22406 );
buf ( n33209 , n17499 );
buf ( n33210 , n380942 );
buf ( n33211 , n18101 );
not ( n33212 , n33211 );
or ( n33213 , n379984 , n33212 );
not ( n33214 , n385161 );
or ( n33215 , n383160 , n33214 );
nand ( n33216 , n33215 , RI15b542d0_737);
nand ( n33217 , n33213 , n33216 , n383165 );
buf ( n33218 , n33217 );
nand ( n33219 , n382974 , n380757 );
not ( n33220 , n33219 );
not ( n33221 , n33220 );
not ( n33222 , n381589 );
or ( n33223 , n33221 , n33222 );
not ( n33224 , n381541 );
nand ( n33225 , n382981 , n33224 );
not ( n33226 , n33225 );
and ( n33227 , n381596 , n33226 );
and ( n33228 , n33225 , n33219 , n380751 );
nor ( n33229 , n33228 , n19630 );
buf ( n33230 , n381493 );
not ( n33231 , n33230 );
nor ( n33232 , n382988 , n33231 );
or ( n33233 , n33229 , n33232 );
nand ( n33234 , n33233 , n19595 );
or ( n33235 , n382992 , n380728 );
nand ( n33236 , n33234 , n33235 );
and ( n33237 , n33236 , n380775 );
or ( n33238 , n33237 , n18708 );
not ( n33239 , n33235 );
nor ( n33240 , n33232 , n33239 );
or ( n33241 , n33229 , n33240 );
or ( n33242 , n382998 , n33241 );
or ( n33243 , n33235 , n381621 );
nand ( n33244 , n33238 , n33242 , n33243 );
nor ( n33245 , n33227 , n33244 );
nand ( n33246 , n33223 , n33245 );
buf ( n33247 , n33246 );
buf ( n33248 , n17499 );
buf ( n33249 , n383174 );
buf ( n33250 , RI15b3ea48_2);
buf ( n33251 , n33250 );
buf ( n33252 , n379844 );
not ( n33253 , n32035 );
nand ( n33254 , n32901 , n33253 );
not ( n33255 , n32912 );
or ( n33256 , n33254 , n33255 );
nand ( n33257 , n32902 , n382080 );
not ( n33258 , n33257 );
or ( n33259 , n33258 , n32024 );
nand ( n33260 , n33259 , n33255 );
buf ( n33261 , n32904 );
not ( n33262 , n33261 );
not ( n33263 , n382495 );
or ( n33264 , n33262 , n33263 );
or ( n33265 , n382495 , n33261 );
nand ( n33266 , n33264 , n33265 );
and ( n33267 , n32963 , n33266 );
and ( n33268 , n382523 , RI15b4bcc0_451);
and ( n33269 , n33159 , RI15b45ac8_242);
nor ( n33270 , n33268 , n33269 );
not ( n33271 , n33270 );
nor ( n33272 , n33267 , n33271 );
nand ( n33273 , n33256 , n33260 , n33272 );
buf ( n33274 , n33273 );
buf ( n33275 , n379802 );
buf ( n33276 , n19653 );
buf ( n33277 , n380203 );
buf ( n33278 , n379847 );
or ( n33279 , n22102 , n32165 );
and ( n33280 , n22203 , n32170 );
not ( n33281 , RI15b43548_162);
or ( n33282 , n32183 , n33281 );
or ( n33283 , n22293 , n32187 );
or ( n33284 , n32181 , n22299 );
nand ( n33285 , n33282 , n33283 , n33284 );
nor ( n33286 , n33280 , n33285 );
nand ( n33287 , n33279 , n33286 );
buf ( n33288 , n33287 );
buf ( n33289 , n380942 );
buf ( n33290 , n382052 );
buf ( n33291 , n381707 );
not ( n33292 , n17576 );
buf ( n33293 , n22516 );
not ( n33294 , n22522 );
nor ( n33295 , n33293 , n33294 );
and ( n33296 , n33292 , n33295 );
and ( n33297 , n18188 , n22617 );
nor ( n33298 , n33297 , n18179 );
or ( n33299 , n33298 , n22835 );
not ( n33300 , n22586 );
or ( n33301 , n33300 , n18079 );
nand ( n33302 , n33301 , n18104 );
nand ( n33303 , n33302 , RI15b562b0_805);
nor ( n33304 , n18197 , RI15b562b0_805);
and ( n33305 , n33300 , n33304 );
not ( n33306 , RI15b58038_868);
or ( n33307 , n22617 , n33306 , RI15b580b0_869);
or ( n33308 , n22835 , RI15b58038_868);
nand ( n33309 , n33307 , n33308 );
and ( n33310 , n18188 , n33309 );
and ( n33311 , n18219 , RI15b571b0_837);
nor ( n33312 , n33305 , n33310 , n33311 );
nand ( n33313 , n33299 , n33303 , n33312 );
nor ( n33314 , n33296 , n33313 );
nand ( n33315 , n33293 , n17507 );
not ( n33316 , n33315 );
not ( n33317 , n17565 );
or ( n33318 , n33316 , n33317 );
nand ( n33319 , n33318 , n33294 );
nand ( n33320 , n33314 , n33319 );
buf ( n33321 , n33320 );
and ( n33322 , n21788 , RI15b56df0_829);
not ( n33323 , n21900 );
buf ( n33324 , n21768 );
and ( n33325 , n33323 , n33324 );
not ( n33326 , n21894 );
and ( n33327 , n33326 , n21898 );
not ( n33328 , n33326 );
and ( n33329 , n33328 , RI15b56df0_829);
nor ( n33330 , n33327 , n33329 );
and ( n33331 , n33330 , n384113 );
nor ( n33332 , n33322 , n33325 , n33331 );
nand ( n33333 , n385154 , n33332 );
buf ( n33334 , n33333 );
buf ( n33335 , n379893 );
buf ( n33336 , n381081 );
buf ( n33337 , n22406 );
or ( n33338 , n31771 , n18235 );
not ( n33339 , n32378 );
and ( n33340 , n33339 , n19370 );
and ( n33341 , n32386 , n18371 );
and ( n33342 , n31778 , n19409 );
nor ( n33343 , n33340 , n33341 , n33342 );
nand ( n33344 , n33338 , n22766 , n33343 );
buf ( n33345 , n33344 );
buf ( n33346 , n22406 );
not ( n33347 , n383129 );
nand ( n33348 , n383137 , n33347 );
not ( n33349 , n33348 );
not ( n33350 , n381460 );
and ( n33351 , n33349 , n33350 );
not ( n33352 , n384184 );
nor ( n33353 , n381400 , n33352 );
nor ( n33354 , n33351 , n33353 );
nand ( n33355 , n381484 , RI15b527a0_679);
or ( n33356 , n33347 , n381423 );
nand ( n33357 , n33356 , n381450 );
not ( n33358 , n383137 );
nand ( n33359 , n33357 , n33358 );
nand ( n33360 , n33354 , n33355 , n33359 );
buf ( n33361 , n33360 );
buf ( n33362 , n380203 );
buf ( n33363 , n382052 );
buf ( n33364 , n22655 );
not ( n33365 , n32165 );
not ( n33366 , n33365 );
not ( n33367 , n33167 );
nand ( n33368 , n33367 , n33170 );
nand ( n33369 , n33368 , n22097 );
not ( n33370 , n33369 );
not ( n33371 , n33370 );
or ( n33372 , n33366 , n33371 );
and ( n33373 , n33196 , n32170 );
not ( n33374 , RI15b436b0_165);
or ( n33375 , n32183 , n33374 );
or ( n33376 , n22241 , n32187 );
or ( n33377 , n32181 , n33201 );
nand ( n33378 , n33375 , n33376 , n33377 );
nor ( n33379 , n33373 , n33378 );
nand ( n33380 , n33372 , n33379 );
buf ( n33381 , n33380 );
buf ( n33382 , RI15b3e9d0_1);
buf ( n33383 , n33382 );
buf ( n33384 , n22408 );
buf ( n33385 , n22716 );
buf ( n33386 , n22788 );
and ( n33387 , n382895 , n382897 );
not ( n33388 , n33387 );
not ( n33389 , n381572 );
not ( n33390 , n381577 );
not ( n33391 , n33390 );
or ( n33392 , n33389 , n33391 );
nand ( n33393 , n33392 , n380686 );
buf ( n33394 , n381578 );
and ( n33395 , n33393 , n33394 );
not ( n33396 , n381578 );
nand ( n33397 , n380698 , n33396 );
nor ( n33398 , n33390 , n33397 );
nor ( n33399 , n33395 , n33398 );
not ( n33400 , n33399 );
not ( n33401 , n33400 );
or ( n33402 , n33388 , n33401 );
not ( n33403 , n382921 );
nand ( n33404 , n33403 , n382929 );
not ( n33405 , n380494 );
nand ( n33406 , n33405 , n380607 );
not ( n33407 , n33406 );
and ( n33408 , n33404 , n33407 , n381522 );
not ( n33409 , n386594 );
buf ( n33410 , n382920 );
nand ( n33411 , n33409 , n33406 , n33410 , n382922 );
or ( n33412 , n33411 , n382917 );
or ( n33413 , n382926 , n380493 );
nand ( n33414 , n33412 , n33413 );
or ( n33415 , n33408 , n33414 );
nand ( n33416 , n381526 , n380737 );
not ( n33417 , n33416 );
and ( n33418 , n33415 , n33417 );
not ( n33419 , n33387 );
and ( n33420 , n33416 , n33419 , n381531 );
nor ( n33421 , n33420 , n19630 );
nor ( n33422 , n381534 , n382941 );
or ( n33423 , n33421 , n33422 );
nand ( n33424 , n33423 , n19595 );
not ( n33425 , n381493 );
or ( n33426 , n381539 , n33425 );
nand ( n33427 , n33424 , n33426 );
and ( n33428 , n33427 , n380775 );
not ( n33429 , RI15b5b698_984);
or ( n33430 , n33428 , n33429 );
buf ( n33431 , n384858 );
buf ( n33432 , n33431 );
buf ( n33433 , n33432 );
not ( n33434 , n33433 );
not ( n33435 , n33422 );
not ( n33436 , n33426 );
not ( n33437 , n33436 );
and ( n33438 , n33435 , n33437 );
nor ( n33439 , n33438 , n33421 );
not ( n33440 , n33439 );
or ( n33441 , n33434 , n33440 );
not ( n33442 , n18919 );
nand ( n33443 , n33442 , n380789 );
or ( n33444 , n33426 , n33443 );
nand ( n33445 , n33430 , n33441 , n33444 );
nor ( n33446 , n33418 , n33445 );
nand ( n33447 , n33402 , n33446 );
buf ( n33448 , n33447 );
not ( n33449 , RI15b53808_714);
not ( n33450 , n383170 );
or ( n33451 , n33449 , n33450 );
not ( n33452 , n385166 );
and ( n33453 , n33452 , n18101 );
not ( n33454 , n33453 );
nor ( n33455 , n381447 , n381458 );
not ( n33456 , n381453 );
nand ( n33457 , n33456 , n383009 );
nand ( n33458 , n33457 , RI15b55770_781);
and ( n33459 , n33458 , RI15b54d20_759);
not ( n33460 , n33458 );
and ( n33461 , n33460 , n382643 );
nor ( n33462 , n33459 , n33461 );
nand ( n33463 , n33455 , n33462 );
or ( n33464 , n33454 , n33463 );
or ( n33465 , n33454 , RI15b55770_781);
nand ( n33466 , n33464 , n33465 );
not ( n33467 , RI15b54d98_760);
not ( n33468 , n33457 );
nand ( n33469 , n33468 , n382643 );
nand ( n33470 , n33469 , RI15b55770_781);
not ( n33471 , n33470 );
or ( n33472 , n33467 , n33471 );
or ( n33473 , n33470 , RI15b54d98_760);
nand ( n33474 , n33472 , n33473 );
and ( n33475 , n33466 , n33474 );
and ( n33476 , n33453 , RI15b55770_781);
not ( n33477 , n33463 );
nor ( n33478 , n33477 , n33474 );
and ( n33479 , n33476 , n33478 );
and ( n33480 , n383147 , RI15b53088_698);
nor ( n33481 , n33475 , n33479 , n33480 );
nand ( n33482 , n33451 , n33481 );
buf ( n33483 , n33482 );
not ( n33484 , RI15b617a0_1191);
nand ( n33485 , n32345 , n33484 );
nor ( n33486 , n33485 , RI15b61818_1192);
not ( n33487 , RI15b61890_1193);
nand ( n33488 , n33486 , n33487 );
not ( n33489 , n33488 );
not ( n33490 , n33489 );
nand ( n33491 , n33490 , RI15b61908_1194);
not ( n33492 , RI15b61980_1195);
and ( n33493 , n33491 , n33492 );
not ( n33494 , n33491 );
and ( n33495 , n33494 , RI15b61980_1195);
nor ( n33496 , n33493 , n33495 );
not ( n33497 , n33496 );
not ( n33498 , RI15b61908_1194);
not ( n33499 , n33490 );
not ( n33500 , n33499 );
or ( n33501 , n33498 , n33500 );
not ( n33502 , n33499 );
not ( n33503 , RI15b61908_1194);
nand ( n33504 , n33502 , n33503 );
nand ( n33505 , n33501 , n33504 );
not ( n33506 , n33505 );
nand ( n33507 , n33497 , n33506 );
not ( n33508 , n33507 );
and ( n33509 , n33499 , RI15b61980_1195);
nor ( n33510 , n33503 , RI15b61980_1195);
nor ( n33511 , n33509 , n33510 );
nand ( n33512 , n33511 , n33504 );
not ( n33513 , n33512 );
not ( n33514 , RI15b619f8_1196);
nor ( n33515 , RI15b61908_1194 , RI15b61980_1195);
and ( n33516 , n33489 , n33515 );
not ( n33517 , n33516 );
or ( n33518 , n33514 , n33517 );
or ( n33519 , n33516 , RI15b619f8_1196);
nand ( n33520 , n33518 , n33519 );
not ( n33521 , n33520 );
not ( n33522 , n33521 );
or ( n33523 , n33513 , n33522 );
not ( n33524 , n33516 );
not ( n33525 , n33524 );
not ( n33526 , n33491 );
nand ( n33527 , n33526 , RI15b61980_1195);
not ( n33528 , n33527 );
or ( n33529 , n33525 , n33528 );
nand ( n33530 , n33529 , n33520 );
nand ( n33531 , n33523 , n33530 );
not ( n33532 , n33531 );
not ( n33533 , n33532 );
or ( n33534 , n33508 , n33533 );
or ( n33535 , n33532 , n33507 );
nand ( n33536 , n33534 , n33535 );
and ( n33537 , RI15b61bd8_1200 , n33536 );
not ( n33538 , RI15b61bd8_1200);
and ( n33539 , n33538 , RI15b619f8_1196);
nor ( n33540 , n33537 , n33539 );
buf ( n33541 , n33540 );
and ( n33542 , n383523 , RI15b61980_1195);
not ( n33543 , n383523 );
not ( n33544 , n33506 );
not ( n33545 , n33496 );
or ( n33546 , n33544 , n33545 );
or ( n33547 , n33496 , n33506 );
nand ( n33548 , n33546 , n33547 );
and ( n33549 , n33543 , n33548 );
nor ( n33550 , n33542 , n33549 );
not ( n33551 , n33499 );
nand ( n33552 , n33551 , RI15b61bd8_1200);
not ( n33553 , n33552 );
buf ( n33554 , n33486 );
nor ( n33555 , n33554 , n33487 );
not ( n33556 , n33555 );
and ( n33557 , n33553 , n33556 );
and ( n33558 , n383523 , RI15b61890_1193);
nor ( n33559 , n33557 , n33558 );
nand ( n33560 , n32338 , n32352 );
not ( n33561 , RI15b61818_1192);
buf ( n33562 , n33485 );
nand ( n33563 , n33562 , RI15b61bd8_1200);
not ( n33564 , n33563 );
or ( n33565 , n33561 , n33564 );
or ( n33566 , n33563 , RI15b61818_1192);
nand ( n33567 , n33565 , n33566 );
nor ( n33568 , n33560 , n33567 );
nand ( n33569 , n33559 , n33568 );
and ( n33570 , n33552 , n33503 );
not ( n33571 , n33552 );
and ( n33572 , n33571 , RI15b61908_1194);
nor ( n33573 , n33570 , n33572 );
nor ( n33574 , n33569 , n33573 );
nand ( n33575 , n33550 , n33574 );
not ( n33576 , n33575 );
buf ( n33577 , n383500 );
buf ( n33578 , n33577 );
not ( n33579 , n33578 );
buf ( n33580 , n33579 );
buf ( n33581 , n33580 );
buf ( n33582 , n33581 );
and ( n33583 , n33576 , n33582 );
or ( n33584 , n384924 , n383589 );
not ( n33585 , n33584 );
nor ( n33586 , n33583 , n33585 );
or ( n33587 , n33541 , n33586 );
or ( n33588 , n384933 , n383589 );
nor ( n33589 , n33576 , n33588 );
nand ( n33590 , n33541 , n33589 );
and ( n33591 , n383601 , RI15b60468_1150);
and ( n33592 , n383607 , RI15b5ee60_1103);
nor ( n33593 , n33591 , n33592 );
nand ( n33594 , n33587 , n33590 , n33593 );
buf ( n33595 , n33594 );
buf ( n33596 , n31979 );
nand ( n33597 , n33109 , n384056 );
or ( n33598 , n31006 , n33597 );
nand ( n33599 , n385004 , n383887 );
not ( n33600 , n33599 );
and ( n33601 , n31016 , n33600 );
and ( n33602 , n33599 , n33597 , n33119 );
nor ( n33603 , n33602 , n21764 );
nor ( n33604 , n385012 , n383865 );
or ( n33605 , n33603 , n33604 );
nand ( n33606 , n33605 , n18154 );
or ( n33607 , n385016 , n383832 );
nand ( n33608 , n33606 , n33607 );
and ( n33609 , n33608 , n383901 );
or ( n33610 , n33609 , n20993 );
not ( n33611 , n31020 );
not ( n33612 , n33611 );
not ( n33613 , n33607 );
nor ( n33614 , n33604 , n33613 );
or ( n33615 , n33603 , n33614 );
or ( n33616 , n33612 , n33615 );
or ( n33617 , n33607 , n31024 );
nand ( n33618 , n33610 , n33616 , n33617 );
nor ( n33619 , n33601 , n33618 );
nand ( n33620 , n33598 , n33619 );
buf ( n33621 , n33620 );
buf ( n33622 , n384996 );
buf ( n33623 , n380203 );
nor ( n33624 , n21320 , n21329 );
not ( n33625 , n33624 );
and ( n33626 , n33625 , n381773 );
not ( n33627 , n33625 );
and ( n33628 , n33627 , n381772 );
nor ( n33629 , n33626 , n33628 );
not ( n33630 , n21361 );
not ( n33631 , n33630 );
and ( n33632 , n33629 , n33631 );
nor ( n33633 , n21537 , n21542 );
not ( n33634 , n33633 );
not ( n33635 , n381742 );
and ( n33636 , n33634 , n33635 );
and ( n33637 , n33633 , n381742 );
nor ( n33638 , n33636 , n33637 );
buf ( n33639 , n21564 );
not ( n33640 , n33639 );
or ( n33641 , n33638 , n33640 );
or ( n33642 , n21737 , n381798 );
nand ( n33643 , n33642 , n381799 );
buf ( n33644 , n385134 );
and ( n33645 , n33643 , n33644 );
and ( n33646 , n21751 , RI15b58038_868);
nor ( n33647 , n33645 , n33646 );
nand ( n33648 , n33641 , n33647 );
nor ( n33649 , n33632 , n33648 );
and ( n33650 , n385164 , RI15b509a0_615);
not ( n33651 , n385174 );
buf ( n33652 , n33651 );
or ( n33653 , n33652 , n381798 );
or ( n33654 , n381773 , n385170 );
or ( n33655 , n381742 , n385178 );
nand ( n33656 , n33653 , n33654 , n33655 );
nor ( n33657 , n33650 , n33656 );
nand ( n33658 , n33649 , n33657 );
buf ( n33659 , n33658 );
buf ( n33660 , n381566 );
buf ( n33661 , n382071 );
not ( n33662 , n379665 );
not ( n33663 , n379565 );
and ( n33664 , n379412 , n379791 );
buf ( n33665 , n33664 );
and ( n33666 , n33663 , n379595 , n379584 , n33665 );
and ( n33667 , n379617 , n379627 );
and ( n33668 , n33666 , n33667 , n379636 );
nand ( n33669 , n33662 , n33668 );
not ( n33670 , n379699 );
nand ( n33671 , n33670 , n379654 );
nor ( n33672 , n33669 , n33671 );
not ( n33673 , n379718 );
and ( n33674 , n33672 , n33673 );
not ( n33675 , n379767 );
nand ( n33676 , n33674 , n33675 );
buf ( n33677 , n379739 );
not ( n33678 , n33677 );
and ( n33679 , n33676 , n33678 );
not ( n33680 , n33676 );
and ( n33681 , n33680 , n33677 );
nor ( n33682 , n33679 , n33681 );
not ( n33683 , n33682 );
not ( n33684 , n33669 );
not ( n33685 , n379673 );
and ( n33686 , n379698 , n33685 );
nand ( n33687 , n33684 , n33686 );
not ( n33688 , n33687 );
not ( n33689 , n379685 );
nor ( n33690 , n33689 , n379668 );
buf ( n33691 , n33690 );
not ( n33692 , n33691 );
and ( n33693 , n33688 , n33692 );
and ( n33694 , n33687 , n33691 );
nor ( n33695 , n33693 , n33694 );
not ( n33696 , n33669 );
not ( n33697 , n379698 );
nand ( n33698 , n33696 , n33697 );
buf ( n33699 , n33685 );
buf ( n33700 , n33699 );
not ( n33701 , n33700 );
not ( n33702 , n33669 );
or ( n33703 , n33701 , n33702 );
not ( n33704 , n33699 );
nand ( n33705 , n33704 , n379698 );
nand ( n33706 , n33703 , n33705 );
not ( n33707 , n33706 );
nand ( n33708 , n33698 , n33707 );
not ( n33709 , n379665 );
buf ( n33710 , n33668 );
not ( n33711 , n33710 );
or ( n33712 , n33709 , n33711 );
or ( n33713 , n33710 , n379665 );
nand ( n33714 , n33712 , n33713 );
not ( n33715 , n33714 );
buf ( n33716 , n33666 );
nand ( n33717 , n33716 , n379618 );
and ( n33718 , n33717 , n379627 );
not ( n33719 , n33717 );
not ( n33720 , n379627 );
and ( n33721 , n33719 , n33720 );
nor ( n33722 , n33718 , n33721 );
buf ( n33723 , n379609 );
not ( n33724 , n33723 );
nand ( n33725 , n33716 , n33724 );
not ( n33726 , n379616 );
and ( n33727 , n33725 , n33726 );
not ( n33728 , n33725 );
and ( n33729 , n33728 , n379616 );
nor ( n33730 , n33727 , n33729 );
nand ( n33731 , n379483 , n33664 );
not ( n33732 , n33731 );
not ( n33733 , n379551 );
not ( n33734 , n379507 );
nor ( n33735 , n33733 , n33734 );
buf ( n33736 , n379497 );
not ( n33737 , n33736 );
not ( n33738 , n33737 );
nand ( n33739 , n33732 , n33735 , n33738 );
not ( n33740 , n379537 );
buf ( n33741 , n33740 );
not ( n33742 , n33741 );
or ( n33743 , n33739 , n33742 );
nor ( n33744 , n33741 , n379589 );
nand ( n33745 , n33739 , n33744 );
nand ( n33746 , n33743 , n33745 , n379535 );
not ( n33747 , n33735 );
not ( n33748 , n33737 );
or ( n33749 , n33731 , n33747 , n33748 );
nand ( n33750 , n33749 , n379493 );
and ( n33751 , n33732 , n33735 );
nand ( n33752 , n33738 , RI15b648d8_1296);
nor ( n33753 , n33751 , n33752 );
nor ( n33754 , n33750 , n33753 );
nand ( n33755 , n33733 , n379507 );
or ( n33756 , n33731 , n33755 );
nand ( n33757 , n379483 , n379507 );
buf ( n33758 , n33757 );
nor ( n33759 , n33664 , n379589 );
or ( n33760 , n33758 , n33759 );
buf ( n33761 , n33733 );
not ( n33762 , n33761 );
nand ( n33763 , n33760 , n33762 );
not ( n33764 , n379548 );
nand ( n33765 , n33756 , n33763 , n33764 );
or ( n33766 , n379507 , n379589 );
nand ( n33767 , n33732 , n33766 );
nor ( n33768 , n33765 , n33767 );
nand ( n33769 , n33754 , n33768 );
nor ( n33770 , n33746 , n33769 );
not ( n33771 , n33757 );
nor ( n33772 , n33740 , n33733 );
nand ( n33773 , n33771 , n33772 , n33736 );
not ( n33774 , n33773 );
not ( n33775 , n33774 );
buf ( n33776 , n379525 );
not ( n33777 , n33776 );
nand ( n33778 , n33777 , n33665 );
or ( n33779 , n33775 , n33778 );
and ( n33780 , n33776 , n33759 );
not ( n33781 , n379523 );
nor ( n33782 , n33780 , n33781 );
nand ( n33783 , n33779 , n33782 );
nor ( n33784 , n33777 , n379589 );
and ( n33785 , n33775 , n33784 );
nor ( n33786 , n33783 , n33785 );
nand ( n33787 , n33770 , n33786 );
buf ( n33788 , n379564 );
not ( n33789 , n33788 );
not ( n33790 , n33789 );
not ( n33791 , n33774 );
nand ( n33792 , n33776 , n33665 );
nor ( n33793 , n33791 , n33792 );
not ( n33794 , n33793 );
or ( n33795 , n33790 , n33794 );
or ( n33796 , n33793 , n33789 );
nand ( n33797 , n33795 , n33796 );
nor ( n33798 , n33787 , n33797 );
nand ( n33799 , n33722 , n33730 , n33798 );
nand ( n33800 , n33716 , n33667 );
and ( n33801 , n33800 , n379636 );
not ( n33802 , n33800 );
and ( n33803 , n33802 , n379637 );
nor ( n33804 , n33801 , n33803 );
not ( n33805 , n33716 );
not ( n33806 , n33724 );
not ( n33807 , n33806 );
and ( n33808 , n33805 , n33807 );
and ( n33809 , n33716 , n33806 );
nor ( n33810 , n33808 , n33809 );
not ( n33811 , n379596 );
not ( n33812 , n33663 );
not ( n33813 , n33665 );
nor ( n33814 , n33812 , n33813 );
buf ( n33815 , n379584 );
nand ( n33816 , n33814 , n33815 );
not ( n33817 , n33816 );
not ( n33818 , n33817 );
or ( n33819 , n33811 , n33818 );
or ( n33820 , n33817 , n379596 );
nand ( n33821 , n33819 , n33820 );
not ( n33822 , n33814 );
not ( n33823 , n33815 );
not ( n33824 , n33823 );
and ( n33825 , n33822 , n33824 );
not ( n33826 , n33822 );
and ( n33827 , n33826 , n33823 );
nor ( n33828 , n33825 , n33827 );
nand ( n33829 , n33793 , n33788 );
nand ( n33830 , n379513 , n379476 );
not ( n33831 , n33830 );
and ( n33832 , n33829 , n33831 );
not ( n33833 , n33829 );
and ( n33834 , n33833 , n33830 );
nor ( n33835 , n33832 , n33834 );
nand ( n33836 , n33828 , n33835 );
nor ( n33837 , n33821 , n33836 );
nand ( n33838 , n33804 , n33810 , n33837 );
nor ( n33839 , n33799 , n33838 );
nand ( n33840 , n33715 , n33839 );
nor ( n33841 , n33708 , n33840 );
nand ( n33842 , n33695 , n33841 );
not ( n33843 , n33842 );
not ( n33844 , n379766 );
nand ( n33845 , n33674 , n33844 );
not ( n33846 , n33845 );
nor ( n33847 , n33674 , n33844 );
nor ( n33848 , n33846 , n33847 );
buf ( n33849 , n379716 );
not ( n33850 , n33849 );
not ( n33851 , n33672 );
not ( n33852 , n33851 );
not ( n33853 , n33852 );
or ( n33854 , n33850 , n33853 );
not ( n33855 , n33669 );
and ( n33856 , n33690 , n33686 );
nand ( n33857 , n33855 , n33856 );
and ( n33858 , n33857 , n379684 );
not ( n33859 , n33857 );
not ( n33860 , n379684 );
and ( n33861 , n33859 , n33860 );
nor ( n33862 , n33858 , n33861 );
nand ( n33863 , n33854 , n33862 );
buf ( n33864 , n379707 );
nor ( n33865 , n33864 , n33849 );
not ( n33866 , n33865 );
not ( n33867 , n33669 );
nand ( n33868 , n33867 , n33670 );
buf ( n33869 , n379654 );
and ( n33870 , n33868 , n33869 );
not ( n33871 , n33868 );
not ( n33872 , n33869 );
and ( n33873 , n33871 , n33872 );
nor ( n33874 , n33870 , n33873 );
nand ( n33875 , n33851 , n33864 );
nand ( n33876 , n33866 , n33874 , n33875 );
nor ( n33877 , n33863 , n33876 );
nand ( n33878 , n33843 , n33848 , n33877 );
not ( n33879 , n33676 );
buf ( n33880 , n379754 );
or ( n33881 , n33674 , n33880 );
not ( n33882 , n33880 );
nand ( n33883 , n33882 , n33844 );
nand ( n33884 , n33881 , n33883 );
nor ( n33885 , n33879 , n33884 );
nor ( n33886 , n33878 , n33885 );
nand ( n33887 , n33683 , n33886 );
not ( n33888 , n33887 );
not ( n33889 , n33676 );
nand ( n33890 , n33889 , n33677 );
and ( n33891 , n33890 , n379731 );
not ( n33892 , n33890 );
not ( n33893 , n379731 );
and ( n33894 , n33892 , n33893 );
nor ( n33895 , n33891 , n33894 );
nand ( n33896 , n33888 , n33895 );
not ( n33897 , n33896 );
not ( n33898 , n33897 );
and ( n33899 , n33674 , n379768 );
buf ( n33900 , n33899 );
not ( n33901 , n33900 );
not ( n33902 , n379463 );
nor ( n33903 , n33901 , n33902 );
not ( n33904 , n33903 );
and ( n33905 , n33898 , n33904 );
not ( n33906 , n33896 );
not ( n33907 , n33900 );
buf ( n33908 , n379456 );
not ( n33909 , n379462 );
nor ( n33910 , n33908 , n33909 );
nand ( n33911 , n33907 , n33910 );
and ( n33912 , n33906 , n33911 );
nor ( n33913 , n33905 , n33912 );
buf ( n33914 , n33908 );
or ( n33915 , n33913 , n33914 );
nor ( n33916 , n33902 , n379773 );
not ( n33917 , n33916 );
not ( n33918 , n33899 );
or ( n33919 , n33917 , n33918 );
nand ( n33920 , n33919 , RI15b648d8_1296);
buf ( n33921 , n33920 );
buf ( n33922 , n33921 );
not ( n33923 , n33922 );
buf ( n33924 , n33923 );
not ( n33925 , n33924 );
not ( n33926 , n33925 );
nand ( n33927 , n33915 , n33926 );
buf ( n33928 , n33921 );
not ( n33929 , n33928 );
not ( n33930 , n33929 );
not ( n33931 , n33886 );
buf ( n33932 , n33682 );
and ( n33933 , n33931 , n33932 );
not ( n33934 , n33931 );
not ( n33935 , n33932 );
and ( n33936 , n33934 , n33935 );
nor ( n33937 , n33933 , n33936 );
not ( n33938 , n33937 );
or ( n33939 , n33930 , n33938 );
nand ( n33940 , n379589 , RI15b646f8_1292);
nand ( n33941 , n33939 , n33940 );
buf ( n33942 , n33878 );
not ( n33943 , n33885 );
xor ( n33944 , n33942 , n33943 );
not ( n33945 , n33923 );
or ( n33946 , n33944 , n33945 );
or ( n33947 , n379448 , RI15b648d8_1296);
nand ( n33948 , n33946 , n33947 );
nor ( n33949 , n33941 , n33948 );
not ( n33950 , n33895 );
and ( n33951 , n33887 , n33950 );
not ( n33952 , n33887 );
and ( n33953 , n33952 , n33895 );
nor ( n33954 , n33951 , n33953 );
buf ( n33955 , n33922 );
not ( n33956 , n33955 );
and ( n33957 , n33954 , n33956 );
not ( n33958 , RI15b64770_1293);
nor ( n33959 , n33958 , RI15b648d8_1296);
nor ( n33960 , n33957 , n33959 );
and ( n33961 , n33949 , n33960 );
not ( n33962 , n33849 );
buf ( n33963 , n33962 );
not ( n33964 , n33963 );
buf ( n33965 , n33852 );
not ( n33966 , n33965 );
or ( n33967 , n33964 , n33966 );
buf ( n33968 , n33963 );
or ( n33969 , n33965 , n33968 );
nand ( n33970 , n33967 , n33969 );
not ( n33971 , n33970 );
buf ( n33972 , n33862 );
not ( n33973 , n33972 );
nor ( n33974 , n33842 , n33973 );
buf ( n33975 , n33874 );
nand ( n33976 , n33974 , n33975 );
not ( n33977 , n33976 );
or ( n33978 , n33971 , n33977 );
buf ( n33979 , n33976 );
or ( n33980 , n33979 , n33970 );
nand ( n33981 , n33978 , n33980 );
and ( n33982 , n33981 , n33923 );
nor ( n33983 , n379711 , RI15b648d8_1296);
nor ( n33984 , n33982 , n33983 );
not ( n33985 , n33922 );
buf ( n33986 , n33975 );
not ( n33987 , n33986 );
and ( n33988 , n33974 , n33987 );
not ( n33989 , n33974 );
and ( n33990 , n33989 , n33986 );
nor ( n33991 , n33988 , n33990 );
not ( n33992 , n33991 );
and ( n33993 , n33985 , n33992 );
and ( n33994 , n379589 , RI15b644a0_1287);
nor ( n33995 , n33993 , n33994 );
nand ( n33996 , n33984 , n33995 );
buf ( n33997 , n33921 );
not ( n33998 , n33810 );
not ( n33999 , n33998 );
and ( n34000 , n33798 , n33835 );
buf ( n34001 , n33828 );
nand ( n34002 , n34000 , n34001 );
nor ( n34003 , n34002 , n33821 );
nand ( n34004 , n33999 , n34003 );
not ( n34005 , n34004 );
not ( n34006 , n34005 );
not ( n34007 , n33730 );
not ( n34008 , n34007 );
and ( n34009 , n34006 , n34008 );
and ( n34010 , n34005 , n34007 );
nor ( n34011 , n34009 , n34010 );
or ( n34012 , n33997 , n34011 );
not ( n34013 , n379613 );
nand ( n34014 , n34012 , n34013 );
not ( n34015 , n34014 );
buf ( n34016 , n33700 );
buf ( n34017 , n34016 );
not ( n34018 , n34017 );
buf ( n34019 , n34018 );
not ( n34020 , n34019 );
not ( n34021 , n34020 );
buf ( n34022 , n33840 );
not ( n34023 , n34022 );
not ( n34024 , n34023 );
or ( n34025 , n34021 , n34024 );
buf ( n34026 , n33696 );
not ( n34027 , n34026 );
and ( n34028 , n34027 , n34022 );
not ( n34029 , n34027 );
and ( n34030 , n34029 , n34019 );
nor ( n34031 , n34028 , n34030 );
nand ( n34032 , n34025 , n34031 );
and ( n34033 , n34032 , n33697 );
buf ( n34034 , n33687 );
not ( n34035 , n34022 );
or ( n34036 , n34034 , n34035 );
not ( n34037 , n34022 );
not ( n34038 , n33705 );
nand ( n34039 , n34037 , n34027 , n34038 );
nand ( n34040 , n34036 , n34039 );
nor ( n34041 , n34033 , n34040 );
or ( n34042 , n33928 , n34041 );
nand ( n34043 , n34042 , n379696 );
not ( n34044 , n34043 );
not ( n34045 , n33922 );
buf ( n34046 , n33722 );
not ( n34047 , n34046 );
not ( n34048 , n34047 );
nor ( n34049 , n34004 , n34007 );
buf ( n34050 , n34049 );
not ( n34051 , n34050 );
or ( n34052 , n34048 , n34051 );
buf ( n34053 , n34050 );
or ( n34054 , n34053 , n34047 );
nand ( n34055 , n34052 , n34054 );
and ( n34056 , n34045 , n34055 );
not ( n34057 , n379624 );
nor ( n34058 , n34056 , n34057 );
nand ( n34059 , n34015 , n34044 , n34058 );
nor ( n34060 , n33996 , n34059 );
not ( n34061 , n34002 );
not ( n34062 , n34061 );
not ( n34063 , n33821 );
and ( n34064 , n34062 , n34063 );
and ( n34065 , n34061 , n33821 );
nor ( n34066 , n34064 , n34065 );
or ( n34067 , n33928 , n34066 );
nor ( n34068 , n379591 , RI15b648d8_1296);
not ( n34069 , n34068 );
nand ( n34070 , n34067 , n34069 );
buf ( n34071 , n33921 );
buf ( n34072 , n34003 );
not ( n34073 , n34072 );
not ( n34074 , n33998 );
and ( n34075 , n34073 , n34074 );
and ( n34076 , n34072 , n33998 );
nor ( n34077 , n34075 , n34076 );
or ( n34078 , n34071 , n34077 );
nand ( n34079 , n34078 , n379608 );
nor ( n34080 , n34070 , n34079 );
not ( n34081 , n33786 );
not ( n34082 , n33770 );
not ( n34083 , n34082 );
or ( n34084 , n34081 , n34083 );
or ( n34085 , n34082 , n33786 );
nand ( n34086 , n34084 , n34085 );
not ( n34087 , n34086 );
not ( n34088 , n33921 );
not ( n34089 , n34088 );
or ( n34090 , n34087 , n34089 );
nand ( n34091 , n34090 , n379523 );
not ( n34092 , n33746 );
buf ( n34093 , n33754 );
or ( n34094 , n34092 , n34093 );
nand ( n34095 , n34094 , n34082 );
buf ( n34096 , n33768 );
buf ( n34097 , n34096 );
buf ( n34098 , n34097 );
nand ( n34099 , n34095 , n34098 );
nor ( n34100 , n34091 , n34099 );
buf ( n34101 , n33921 );
buf ( n34102 , n33839 );
not ( n34103 , n34102 );
not ( n34104 , n33714 );
and ( n34105 , n34103 , n34104 );
and ( n34106 , n34102 , n33714 );
nor ( n34107 , n34105 , n34106 );
or ( n34108 , n34101 , n34107 );
not ( n34109 , n379663 );
nand ( n34110 , n34108 , n34109 );
not ( n34111 , n33804 );
not ( n34112 , n34111 );
and ( n34113 , n34049 , n34046 );
not ( n34114 , n34113 );
or ( n34115 , n34112 , n34114 );
or ( n34116 , n34113 , n34111 );
nand ( n34117 , n34115 , n34116 );
not ( n34118 , n34117 );
not ( n34119 , n34088 );
or ( n34120 , n34118 , n34119 );
nand ( n34121 , n379589 , RI15b641d0_1281);
nand ( n34122 , n34120 , n34121 );
nor ( n34123 , n34110 , n34122 );
buf ( n34124 , n34123 );
not ( n34125 , n34000 );
not ( n34126 , n34001 );
not ( n34127 , n34126 );
and ( n34128 , n34125 , n34127 );
and ( n34129 , n34000 , n34126 );
nor ( n34130 , n34128 , n34129 );
or ( n34131 , n33928 , n34130 );
nand ( n34132 , n34131 , n379582 );
not ( n34133 , n33787 );
not ( n34134 , n34133 );
not ( n34135 , n33797 );
and ( n34136 , n34134 , n34135 );
and ( n34137 , n34133 , n33797 );
nor ( n34138 , n34136 , n34137 );
or ( n34139 , n33921 , n34138 );
nand ( n34140 , n34139 , n379558 );
not ( n34141 , n34140 );
not ( n34142 , n34141 );
nor ( n34143 , n34132 , n34142 );
and ( n34144 , n34080 , n34100 , n34124 , n34143 );
nand ( n34145 , n33927 , n33961 , n34060 , n34144 );
xor ( n34146 , n379462 , n33900 );
xnor ( n34147 , n34146 , n33896 );
not ( n34148 , n33955 );
and ( n34149 , n34147 , n34148 );
nor ( n34150 , n379451 , RI15b648d8_1296);
nor ( n34151 , n34149 , n34150 );
not ( n34152 , n33864 );
buf ( n34153 , n34152 );
and ( n34154 , n33965 , n34153 );
not ( n34155 , n33965 );
nor ( n34156 , n34152 , n33962 );
and ( n34157 , n34155 , n34156 );
nor ( n34158 , n34154 , n34157 );
nor ( n34159 , n33976 , n34158 );
not ( n34160 , n34159 );
not ( n34161 , n33968 );
not ( n34162 , n34161 );
not ( n34163 , n34153 );
or ( n34164 , n34162 , n34163 );
not ( n34165 , n33674 );
nand ( n34166 , n34164 , n34165 );
nand ( n34167 , n33976 , n34166 );
not ( n34168 , n33965 );
nand ( n34169 , n34168 , n33865 );
nand ( n34170 , n34160 , n34167 , n34169 );
not ( n34171 , n34071 );
and ( n34172 , n34170 , n34171 );
nor ( n34173 , n379445 , RI15b648d8_1296);
nor ( n34174 , n34172 , n34173 );
not ( n34175 , n33848 );
not ( n34176 , n33842 );
buf ( n34177 , n33877 );
nand ( n34178 , n34176 , n34177 );
not ( n34179 , n34178 );
or ( n34180 , n34175 , n34179 );
buf ( n34181 , n33845 );
nand ( n34182 , n34180 , n34181 );
not ( n34183 , n34182 );
not ( n34184 , n33921 );
not ( n34185 , n34184 );
or ( n34186 , n34183 , n34185 );
nand ( n34187 , n379589 , RI15b64608_1290);
nand ( n34188 , n34186 , n34187 );
xnor ( n34189 , n34093 , n34097 );
or ( n34190 , n33921 , n34189 );
nand ( n34191 , n34190 , n379493 );
not ( n34192 , n34191 );
nand ( n34193 , n379589 , RI15b64860_1295);
nand ( n34194 , n34192 , n34193 );
not ( n34195 , n34026 );
not ( n34196 , n34195 );
not ( n34197 , n34018 );
and ( n34198 , n34196 , n34197 );
not ( n34199 , n34026 );
and ( n34200 , n34199 , n34018 );
nor ( n34201 , n34198 , n34200 );
and ( n34202 , n34201 , n34035 );
not ( n34203 , n34201 );
not ( n34204 , n34023 );
and ( n34205 , n34203 , n34204 );
nor ( n34206 , n34202 , n34205 );
or ( n34207 , n34101 , n34206 );
nand ( n34208 , n34207 , n379672 );
buf ( n34209 , n34208 );
nor ( n34210 , n34188 , n34194 , n34209 );
buf ( n34211 , n33842 );
not ( n34212 , n34211 );
buf ( n34213 , n33972 );
not ( n34214 , n34213 );
and ( n34215 , n34212 , n34214 );
and ( n34216 , n34211 , n34213 );
nor ( n34217 , n34215 , n34216 );
or ( n34218 , n34071 , n34217 );
nand ( n34219 , n379589 , RI15b64428_1286);
nand ( n34220 , n34218 , n34219 );
not ( n34221 , n33695 );
buf ( n34222 , n33841 );
and ( n34223 , n34221 , n34222 );
not ( n34224 , n34221 );
not ( n34225 , n34222 );
and ( n34226 , n34224 , n34225 );
nor ( n34227 , n34223 , n34226 );
or ( n34228 , n34071 , n34227 );
nand ( n34229 , n379589 , RI15b643b0_1285);
nand ( n34230 , n34228 , n34229 );
nor ( n34231 , n34220 , n34230 );
buf ( n34232 , n33798 );
not ( n34233 , n34232 );
not ( n34234 , n33835 );
not ( n34235 , n34234 );
and ( n34236 , n34233 , n34235 );
and ( n34237 , n34232 , n34234 );
nor ( n34238 , n34236 , n34237 );
or ( n34239 , n33997 , n34238 );
not ( n34240 , n379512 );
nand ( n34241 , n34239 , n34240 );
not ( n34242 , n34241 );
and ( n34243 , n34174 , n34210 , n34231 , n34242 );
nand ( n34244 , n34151 , n34243 );
nor ( n34245 , n34145 , n34244 );
buf ( n34246 , n33926 );
not ( n34247 , n34246 );
nor ( n34248 , n34245 , n34247 );
and ( n34249 , n34248 , n379785 );
not ( n34250 , n34249 );
not ( n34251 , n34250 );
not ( n34252 , n33922 );
and ( n34253 , n34091 , n34252 );
not ( n34254 , n34091 );
and ( n34255 , n34254 , n34071 );
nor ( n34256 , n34253 , n34255 );
or ( n34257 , n34092 , n34098 );
not ( n34258 , n34095 );
nand ( n34259 , n34257 , n34258 );
not ( n34260 , n34259 );
not ( n34261 , n34184 );
or ( n34262 , n34260 , n34261 );
nand ( n34263 , n34262 , n379535 );
not ( n34264 , n34208 );
and ( n34265 , n34263 , n34264 , n34141 );
nand ( n34266 , n34256 , n34265 );
nor ( n34267 , n34241 , n34132 );
nand ( n34268 , n34080 , n34267 );
nor ( n34269 , n34266 , n34268 );
buf ( n34270 , n33813 );
not ( n34271 , n34270 );
nand ( n34272 , n34271 , n33766 );
nor ( n34273 , n33921 , n34272 );
not ( n34274 , n33765 );
not ( n34275 , n33767 );
nor ( n34276 , n34274 , n34275 );
or ( n34277 , n34276 , n34096 );
nand ( n34278 , n34277 , n33764 );
not ( n34279 , n379483 );
nor ( n34280 , n34278 , n34279 );
nand ( n34281 , n34273 , n34280 );
nor ( n34282 , n34281 , n34191 );
and ( n34283 , n34123 , n34282 );
not ( n34284 , n34188 );
and ( n34285 , n34283 , n34174 , n34231 , n34284 );
nand ( n34286 , n34060 , n34269 , n34285 );
buf ( n34287 , n34286 );
buf ( n34288 , n33948 );
not ( n34289 , n34288 );
nand ( n34290 , n34287 , n34289 );
not ( n34291 , n34290 );
and ( n34292 , n34251 , n34291 );
or ( n34293 , n34145 , n34244 );
nand ( n34294 , n34293 , n34246 );
and ( n34295 , n34294 , n379785 );
not ( n34296 , n34295 );
not ( n34297 , n34287 );
nand ( n34298 , n34297 , n379785 );
nand ( n34299 , n34296 , n34298 );
not ( n34300 , n34289 );
and ( n34301 , n34299 , n34300 );
nor ( n34302 , n34292 , n34301 );
not ( n34303 , n33761 );
nand ( n34304 , n379779 , n34303 );
not ( n34305 , n34304 );
not ( n34306 , n34279 );
nand ( n34307 , n34306 , n379779 );
and ( n34308 , n33766 , n379412 );
nand ( n34309 , n379779 , n34308 );
nor ( n34310 , n34307 , n34309 );
nand ( n34311 , n34305 , n34310 );
not ( n34312 , n33784 );
and ( n34313 , n34312 , n379523 );
nor ( n34314 , n33773 , n379413 );
nor ( n34315 , n34313 , n34314 );
not ( n34316 , n34315 );
not ( n34317 , n34316 );
and ( n34318 , n34314 , n33776 );
and ( n34319 , n34318 , n379523 );
not ( n34320 , n34319 );
not ( n34321 , n34320 );
or ( n34322 , n34317 , n34321 );
nand ( n34323 , n34322 , n379779 );
not ( n34324 , n34320 );
not ( n34325 , n33789 );
not ( n34326 , n34318 );
or ( n34327 , n34325 , n34326 );
nand ( n34328 , n34327 , n379558 );
nand ( n34329 , n33788 , RI15b648d8_1296);
nor ( n34330 , n34318 , n34329 );
nor ( n34331 , n34328 , n34330 );
buf ( n34332 , n34331 );
not ( n34333 , n34332 );
or ( n34334 , n34324 , n34333 );
or ( n34335 , n34332 , n34320 );
nand ( n34336 , n34334 , n34335 );
nor ( n34337 , n34323 , n34336 );
nand ( n34338 , n34331 , n34319 );
nand ( n34339 , n34318 , n33788 );
nor ( n34340 , n34339 , n33831 );
not ( n34341 , n34340 );
nor ( n34342 , n33830 , n379589 );
nand ( n34343 , n34339 , n34342 );
nand ( n34344 , n34341 , n34343 , n34240 );
nor ( n34345 , n34338 , n34344 );
not ( n34346 , n379566 );
and ( n34347 , n34346 , n33823 );
not ( n34348 , n34346 );
not ( n34349 , n33823 );
and ( n34350 , n34348 , n34349 );
nor ( n34351 , n34347 , n34350 );
and ( n34352 , n34351 , RI15b648d8_1296);
not ( n34353 , n379582 );
nor ( n34354 , n34352 , n34353 );
and ( n34355 , n34345 , n34354 );
not ( n34356 , n379616 );
not ( n34357 , n379597 );
nor ( n34358 , n34357 , n33723 );
not ( n34359 , n34358 );
or ( n34360 , n34356 , n34359 );
nand ( n34361 , n34360 , n34013 );
nand ( n34362 , n33726 , RI15b648d8_1296);
nor ( n34363 , n34358 , n34362 );
nor ( n34364 , n34361 , n34363 );
not ( n34365 , n33723 );
not ( n34366 , n34357 );
not ( n34367 , n34366 );
or ( n34368 , n34365 , n34367 );
not ( n34369 , n34357 );
not ( n34370 , n33724 );
or ( n34371 , n34369 , n34370 );
nand ( n34372 , n34368 , n34371 );
and ( n34373 , n34372 , RI15b648d8_1296);
not ( n34374 , n379608 );
nor ( n34375 , n34373 , n34374 );
buf ( n34376 , n379585 );
and ( n34377 , n34376 , n379596 );
not ( n34378 , n34376 );
and ( n34379 , n34378 , n379595 );
nor ( n34380 , n34377 , n34379 );
and ( n34381 , n34380 , RI15b648d8_1296);
nor ( n34382 , n34381 , n34068 );
and ( n34383 , n34364 , n34375 , n34382 );
nand ( n34384 , n34355 , n34383 );
buf ( n34385 , n379619 );
and ( n34386 , n34385 , n33720 );
nor ( n34387 , n34386 , n34057 );
not ( n34388 , n34385 );
nor ( n34389 , n33720 , n379589 );
nand ( n34390 , n34388 , n34389 );
nand ( n34391 , n34387 , n34390 );
nor ( n34392 , n34384 , n34391 );
nor ( n34393 , n379637 , n379589 );
not ( n34394 , n34393 );
buf ( n34395 , n379628 );
not ( n34396 , n34395 );
or ( n34397 , n34394 , n34396 );
nand ( n34398 , n34397 , n34121 );
nor ( n34399 , n34395 , n379636 );
nor ( n34400 , n34398 , n34399 );
and ( n34401 , n34392 , n34400 );
not ( n34402 , n379665 );
buf ( n34403 , n379638 );
not ( n34404 , n34403 );
or ( n34405 , n34402 , n34404 );
or ( n34406 , n34403 , n379665 );
nand ( n34407 , n34405 , n34406 );
and ( n34408 , n34407 , RI15b648d8_1296);
nor ( n34409 , n34408 , n379663 );
nand ( n34410 , n34401 , n34409 );
not ( n34411 , n34410 );
nand ( n34412 , n34403 , n379666 );
nor ( n34413 , n34412 , n379589 );
not ( n34414 , n34017 );
and ( n34415 , n34413 , n34414 );
not ( n34416 , n34016 );
nor ( n34417 , n34416 , n379589 );
not ( n34418 , n34417 );
not ( n34419 , n34412 );
or ( n34420 , n34418 , n34419 );
nand ( n34421 , n34420 , n379672 );
nor ( n34422 , n34415 , n34421 );
not ( n34423 , n34422 );
and ( n34424 , n34411 , n34423 );
and ( n34425 , n34410 , n34422 );
nor ( n34426 , n34424 , n34425 );
buf ( n34427 , n33742 );
and ( n34428 , n379779 , n34427 );
not ( n34429 , n34409 );
not ( n34430 , n34429 );
not ( n34431 , n34401 );
or ( n34432 , n34430 , n34431 );
or ( n34433 , n34401 , n34429 );
nand ( n34434 , n34432 , n34433 );
buf ( n34435 , n34382 );
nand ( n34436 , n34355 , n34435 );
buf ( n34437 , n34375 );
and ( n34438 , n34436 , n34437 );
not ( n34439 , n34436 );
not ( n34440 , n34437 );
and ( n34441 , n34439 , n34440 );
nor ( n34442 , n34438 , n34441 );
not ( n34443 , n34391 );
and ( n34444 , n34384 , n34443 );
not ( n34445 , n34384 );
and ( n34446 , n34445 , n34391 );
nor ( n34447 , n34444 , n34446 );
not ( n34448 , n34355 );
not ( n34449 , n34435 );
not ( n34450 , n34449 );
and ( n34451 , n34448 , n34450 );
and ( n34452 , n34355 , n34449 );
nor ( n34453 , n34451 , n34452 );
buf ( n34454 , n34354 );
not ( n34455 , n34454 );
not ( n34456 , n34345 );
not ( n34457 , n34456 );
or ( n34458 , n34455 , n34457 );
or ( n34459 , n34456 , n34454 );
nand ( n34460 , n34458 , n34459 );
not ( n34461 , n34338 );
not ( n34462 , n34461 );
buf ( n34463 , n34344 );
not ( n34464 , n34463 );
and ( n34465 , n34462 , n34464 );
and ( n34466 , n34461 , n34463 );
nor ( n34467 , n34465 , n34466 );
buf ( n34468 , n33748 );
nand ( n34469 , n34467 , n34468 );
nor ( n34470 , n34460 , n34469 );
and ( n34471 , n34453 , n34470 );
nand ( n34472 , n34442 , n34447 , n34471 );
not ( n34473 , n34472 );
buf ( n34474 , n34392 );
not ( n34475 , n34474 );
not ( n34476 , n34400 );
not ( n34477 , n34476 );
and ( n34478 , n34475 , n34477 );
and ( n34479 , n34474 , n34476 );
nor ( n34480 , n34478 , n34479 );
not ( n34481 , n34436 );
nand ( n34482 , n34481 , n34437 );
buf ( n34483 , n34364 );
and ( n34484 , n34482 , n34483 );
not ( n34485 , n34482 );
not ( n34486 , n34483 );
and ( n34487 , n34485 , n34486 );
nor ( n34488 , n34484 , n34487 );
nand ( n34489 , n34473 , n34480 , n34488 );
nor ( n34490 , n34434 , n34489 );
nand ( n34491 , n34337 , n34426 , n34428 , n34490 );
nor ( n34492 , n34311 , n34491 );
not ( n34493 , n34410 );
nand ( n34494 , n34493 , n34422 );
not ( n34495 , n34494 );
not ( n34496 , n34495 );
not ( n34497 , n34017 );
not ( n34498 , n34412 );
not ( n34499 , n34498 );
or ( n34500 , n34497 , n34499 );
nor ( n34501 , n33697 , n379589 );
nand ( n34502 , n34500 , n34501 );
and ( n34503 , n34502 , n379696 );
not ( n34504 , n34018 );
nand ( n34505 , n34413 , n34504 , n33697 );
nand ( n34506 , n34503 , n34505 );
not ( n34507 , n34506 );
and ( n34508 , n34496 , n34507 );
and ( n34509 , n34495 , n34506 );
nor ( n34510 , n34508 , n34509 );
and ( n34511 , n34492 , n34510 );
nor ( n34512 , n34494 , n34506 );
buf ( n34513 , n34512 );
not ( n34514 , n34513 );
not ( n34515 , n33686 );
or ( n34516 , n34412 , n34515 );
buf ( n34517 , n33691 );
not ( n34518 , n34517 );
nor ( n34519 , n34518 , n379589 );
nand ( n34520 , n34516 , n34519 );
and ( n34521 , n34520 , n34229 );
nor ( n34522 , n34517 , n34515 );
nand ( n34523 , n34413 , n34522 );
nand ( n34524 , n34521 , n34523 );
not ( n34525 , n34524 );
and ( n34526 , n34514 , n34525 );
and ( n34527 , n34513 , n34524 );
nor ( n34528 , n34526 , n34527 );
nand ( n34529 , n34511 , n34528 );
not ( n34530 , n34524 );
nand ( n34531 , n34530 , n34512 );
and ( n34532 , n33856 , n33860 );
nand ( n34533 , n34413 , n34532 );
not ( n34534 , n33856 );
not ( n34535 , n34498 );
or ( n34536 , n34534 , n34535 );
nand ( n34537 , n34536 , n379684 );
nand ( n34538 , n34533 , n34537 );
and ( n34539 , n34531 , n34538 );
not ( n34540 , n34531 );
not ( n34541 , n34538 );
and ( n34542 , n34540 , n34541 );
nor ( n34543 , n34539 , n34542 );
nor ( n34544 , n34529 , n34543 );
nor ( n34545 , n34531 , n34538 );
not ( n34546 , n34545 );
nand ( n34547 , n34498 , n33670 );
buf ( n34548 , n33872 );
not ( n34549 , n34548 );
and ( n34550 , n34547 , n34549 );
not ( n34551 , n34547 );
and ( n34552 , n34551 , n34548 );
or ( n34553 , n34550 , n34552 );
not ( n34554 , n34553 );
and ( n34555 , n34546 , n34554 );
and ( n34556 , n34545 , n34553 );
nor ( n34557 , n34555 , n34556 );
nand ( n34558 , n34544 , n34557 );
buf ( n34559 , n379701 );
buf ( n34560 , n34559 );
not ( n34561 , n34161 );
buf ( n34562 , n34561 );
xor ( n34563 , n34560 , n34562 );
or ( n34564 , n34538 , n34553 );
nor ( n34565 , n34531 , n34564 );
not ( n34566 , n34565 );
xnor ( n34567 , n34563 , n34566 );
nor ( n34568 , n34558 , n34567 );
and ( n34569 , n34560 , n34156 );
nor ( n34570 , n34569 , n33865 );
not ( n34571 , n34570 );
not ( n34572 , n34571 );
not ( n34573 , n34566 );
not ( n34574 , n34573 );
or ( n34575 , n34572 , n34574 );
not ( n34576 , n34153 );
nor ( n34577 , n34559 , n34576 );
not ( n34578 , n34562 );
nand ( n34579 , n34577 , n34578 );
nand ( n34580 , n34575 , n34579 );
not ( n34581 , n34576 );
and ( n34582 , n34560 , n34581 );
buf ( n34583 , n379719 );
buf ( n34584 , n34583 );
buf ( n34585 , n34584 );
nor ( n34586 , n34582 , n34585 );
nor ( n34587 , n34573 , n34586 );
nor ( n34588 , n34580 , n34587 );
nand ( n34589 , n34568 , n34588 );
buf ( n34590 , n34585 );
xor ( n34591 , n33844 , n34590 );
and ( n34592 , n34559 , n34561 );
nor ( n34593 , n34592 , n34577 , n34156 );
nand ( n34594 , n34565 , n34593 );
not ( n34595 , n34594 );
not ( n34596 , n34595 );
xnor ( n34597 , n34591 , n34596 );
nor ( n34598 , n34589 , n34597 );
not ( n34599 , n34595 );
buf ( n34600 , n33880 );
nand ( n34601 , n34600 , n33844 );
or ( n34602 , n34585 , n34601 );
not ( n34603 , n34600 );
nand ( n34604 , n34584 , n34603 );
nand ( n34605 , n34602 , n34604 );
not ( n34606 , n34605 );
or ( n34607 , n34599 , n34606 );
or ( n34608 , n34584 , n33844 );
not ( n34609 , n34603 );
or ( n34610 , n34608 , n34609 );
nand ( n34611 , n34607 , n34610 );
not ( n34612 , n34599 );
nand ( n34613 , n34583 , n33675 );
and ( n34614 , n34613 , n33883 );
nor ( n34615 , n34612 , n34614 );
nor ( n34616 , n34611 , n34615 );
and ( n34617 , n34598 , n34616 );
not ( n34618 , n34617 );
nand ( n34619 , n34604 , n34608 , n34601 );
nor ( n34620 , n34594 , n34619 );
not ( n34621 , n34620 );
buf ( n34622 , n33677 );
buf ( n34623 , n34622 );
and ( n34624 , n34613 , n34623 );
not ( n34625 , n34613 );
not ( n34626 , n34623 );
and ( n34627 , n34625 , n34626 );
nor ( n34628 , n34624 , n34627 );
and ( n34629 , n34621 , n34628 );
not ( n34630 , n34612 );
not ( n34631 , n34630 );
or ( n34632 , n34585 , n33883 );
nand ( n34633 , n34632 , n34613 );
not ( n34634 , n34633 );
nor ( n34635 , n34634 , n34628 );
and ( n34636 , n34631 , n34635 );
nor ( n34637 , n34629 , n34636 );
not ( n34638 , n34637 );
and ( n34639 , n34618 , n34638 );
not ( n34640 , n34618 );
and ( n34641 , n34640 , n34637 );
nor ( n34642 , n34639 , n34641 );
buf ( n34643 , n379780 );
buf ( n34644 , n34643 );
not ( n34645 , n34644 );
not ( n34646 , n34645 );
buf ( n34647 , n34646 );
nand ( n34648 , n34642 , n34647 );
and ( n34649 , n379783 , RI15b646f8_1292);
buf ( n34650 , n379796 );
buf ( n34651 , n34650 );
and ( n34652 , n34651 , RI15b5e500_1083);
nor ( n34653 , n34649 , n34652 );
nand ( n34654 , n34302 , n34648 , n34653 );
buf ( n34655 , n34654 );
buf ( n34656 , n379802 );
not ( n34657 , n17507 );
not ( n34658 , n21827 );
not ( n34659 , n34658 );
or ( n34660 , n34657 , n34659 );
nand ( n34661 , n34660 , n17565 );
nand ( n34662 , n34661 , n21835 );
nor ( n34663 , n34658 , n21835 );
nand ( n34664 , n17578 , n34663 );
not ( n34665 , RI15b578b8_852);
or ( n34666 , n21922 , n21927 );
nand ( n34667 , n34666 , n21946 );
not ( n34668 , n34667 );
or ( n34669 , n34665 , n34668 );
not ( n34670 , n21955 );
and ( n34671 , n21949 , n34670 );
nor ( n34672 , n34671 , n379860 );
or ( n34673 , n34672 , n379956 );
nand ( n34674 , n34669 , n34673 );
and ( n34675 , n34674 , n18077 );
or ( n34676 , n22601 , n34670 , RI15b55ab8_788);
and ( n34677 , n18177 , RI15b578b8_852);
and ( n34678 , n18219 , RI15b569b8_820);
nor ( n34679 , n34677 , n34678 , n21751 );
nand ( n34680 , n34676 , n34679 );
not ( n34681 , n21927 );
nor ( n34682 , n18189 , n34681 , RI15b578b8_852);
nor ( n34683 , n34675 , n34680 , n34682 );
nand ( n34684 , n34662 , n34664 , n34683 );
buf ( n34685 , n34684 );
buf ( n34686 , n379895 );
buf ( n34687 , n20663 );
or ( n34688 , n18179 , n18188 );
nand ( n34689 , n34688 , RI15b575e8_846);
nand ( n34690 , n18079 , n18102 );
and ( n34691 , n34690 , RI15b557e8_782);
or ( n34692 , n379924 , RI15b50e50_625);
or ( n34693 , n18219 , n17507 );
nand ( n34694 , n34693 , RI15b566e8_814);
nand ( n34695 , n34692 , n34694 );
nor ( n34696 , n34691 , n34695 );
nand ( n34697 , n34689 , n34696 );
buf ( n34698 , n34697 );
buf ( n34699 , n379847 );
buf ( n34700 , n33382 );
buf ( n34701 , n380942 );
or ( n34702 , n386588 , n33219 );
and ( n34703 , n386600 , n33226 );
not ( n34704 , RI15b5a9f0_957);
or ( n34705 , n33237 , n34704 );
buf ( n34706 , n386617 );
or ( n34707 , n34706 , n33241 );
or ( n34708 , n33235 , n386627 );
nand ( n34709 , n34705 , n34707 , n34708 );
nor ( n34710 , n34703 , n34709 );
nand ( n34711 , n34702 , n34710 );
buf ( n34712 , n34711 );
buf ( n34713 , n18226 );
not ( n34714 , RI15b54618_744);
nor ( n34715 , RI15b54690_745 , RI15b54708_746);
not ( n34716 , RI15b575e8_846);
nand ( n34717 , n34714 , n34715 , n34716 );
and ( n34718 , RI15b54618_744 , RI15b54690_745);
nor ( n34719 , n34718 , RI15b54708_746);
nand ( n34720 , n34719 , RI15b57660_847);
nand ( n34721 , n34717 , n34720 );
buf ( n34722 , n34721 );
buf ( n34723 , n381490 );
buf ( n34724 , RI15b46fe0_287);
buf ( n34725 , n22738 );
buf ( n34726 , n30992 );
nand ( n34727 , n30890 , n386425 );
not ( n34728 , n386419 );
nor ( n34729 , n34727 , n34728 );
and ( n34730 , n34729 , n386414 );
buf ( n34731 , n386409 );
nand ( n34732 , n34730 , n34731 );
not ( n34733 , n386388 );
nor ( n34734 , n34732 , n34733 );
buf ( n34735 , n386376 );
nand ( n34736 , n34734 , n34735 );
not ( n34737 , n386398 );
nor ( n34738 , n34736 , n34737 );
buf ( n34739 , n386383 );
nand ( n34740 , n34738 , n34739 );
not ( n34741 , n386404 );
nor ( n34742 , n34740 , n34741 );
buf ( n34743 , n386393 );
nand ( n34744 , n34742 , n34743 );
not ( n34745 , n34744 );
nor ( n34746 , n34745 , n386446 );
not ( n34747 , n34746 );
not ( n34748 , n386446 );
nor ( n34749 , n34744 , n34748 );
not ( n34750 , n34749 );
nand ( n34751 , n34747 , n34750 );
nand ( n34752 , n34751 , n386500 );
nand ( n34753 , n386174 , n386210 );
not ( n34754 , n386202 );
nor ( n34755 , n34753 , n34754 );
not ( n34756 , n386194 );
nand ( n34757 , n34755 , n34756 );
nor ( n34758 , n34757 , n386186 );
not ( n34759 , n34758 );
and ( n34760 , n34759 , n386198 );
not ( n34761 , n34759 );
not ( n34762 , n386198 );
and ( n34763 , n34761 , n34762 );
nor ( n34764 , n34760 , n34763 );
not ( n34765 , n386261 );
not ( n34766 , n34765 );
not ( n34767 , n34766 );
and ( n34768 , n34764 , n34767 );
not ( n34769 , n385902 );
buf ( n34770 , n385836 );
nor ( n34771 , n34770 , n385891 );
nand ( n34772 , n34769 , n34771 );
buf ( n34773 , n34772 );
not ( n34774 , n385906 );
and ( n34775 , n34773 , n34774 );
not ( n34776 , n34773 );
and ( n34777 , n34776 , n385906 );
nor ( n34778 , n34775 , n34777 );
buf ( n34779 , n30873 );
not ( n34780 , n34779 );
or ( n34781 , n34778 , n34780 );
not ( n34782 , n22396 );
not ( n34783 , n34782 );
not ( n34784 , n34783 );
buf ( n34785 , n34784 );
or ( n34786 , n34785 , n382119 );
nand ( n34787 , n34781 , n34786 );
nor ( n34788 , n34768 , n34787 );
nand ( n34789 , n34752 , n34788 );
not ( n34790 , n34789 );
or ( n34791 , n20638 , n19841 );
buf ( n34792 , n19675 );
not ( n34793 , n34792 );
not ( n34794 , n34793 );
nand ( n34795 , n34794 , n20637 );
and ( n34796 , n30907 , n34795 );
nand ( n34797 , n20637 , n19824 );
and ( n34798 , n34796 , n34797 );
nand ( n34799 , n34791 , n34798 );
and ( n34800 , n34799 , RI15b4ab68_414);
or ( n34801 , n34792 , n20638 , n19824 );
or ( n34802 , n34801 , n19686 , RI15b4ab68_414);
buf ( n34803 , n19846 );
or ( n34804 , n34803 , n22216 );
nand ( n34805 , n34802 , n34804 );
nor ( n34806 , n34800 , n34805 );
nand ( n34807 , n34790 , n34806 );
buf ( n34808 , n34807 );
buf ( n34809 , n32160 );
buf ( n34810 , n22421 );
not ( n34811 , n34810 );
not ( n34812 , n34811 );
and ( n34813 , n34812 , RI15b64338_1284);
buf ( n34814 , n22455 );
not ( n34815 , n34814 );
not ( n34816 , n34815 );
not ( n34817 , n34816 );
buf ( n34818 , n386982 );
not ( n34819 , n34818 );
or ( n34820 , n34817 , n34819 );
and ( n34821 , n22434 , n22418 , n22445 );
and ( n34822 , n22455 , n383406 );
nor ( n34823 , n34821 , n34822 );
nand ( n34824 , n34820 , n34823 );
and ( n34825 , n34824 , RI15b62538_1220);
nand ( n34826 , n22455 , RI15b62ad8_1232);
or ( n34827 , n34818 , n34826 , RI15b62538_1220);
not ( n34828 , n387037 );
and ( n34829 , n34828 , RI15b64338_1284);
not ( n34830 , n34828 );
and ( n34831 , n34830 , n379437 );
nor ( n34832 , n34829 , n34831 );
not ( n34833 , n22449 );
or ( n34834 , n34832 , n34833 );
nand ( n34835 , n34827 , n34834 );
nor ( n34836 , n34813 , n34825 , n34835 );
or ( n34837 , n34836 , n19200 );
buf ( n34838 , n386886 );
and ( n34839 , n34838 , n19628 );
nor ( n34840 , n34839 , n386944 );
or ( n34841 , n386892 , n34840 );
not ( n34842 , n34838 );
buf ( n34843 , n383464 );
not ( n34844 , n34843 );
and ( n34845 , n34842 , n34844 , n386892 );
or ( n34846 , n22424 , n379437 );
or ( n34847 , n383441 , n19598 );
nand ( n34848 , n34846 , n34847 , n19512 );
nor ( n34849 , n34845 , n34848 );
nand ( n34850 , n34837 , n34841 , n34849 );
buf ( n34851 , n34850 );
buf ( n34852 , n380903 );
not ( n34853 , n31507 );
nor ( n34854 , n379337 , n34853 );
not ( n34855 , n31509 );
nand ( n34856 , n34854 , n34855 );
buf ( n34857 , n31501 );
not ( n34858 , n34857 );
nor ( n34859 , n34856 , n34858 );
buf ( n34860 , n34859 );
not ( n34861 , n34860 );
not ( n34862 , n31485 );
and ( n34863 , n34861 , n34862 );
buf ( n34864 , n34860 );
and ( n34865 , n34864 , n31485 );
nor ( n34866 , n34863 , n34865 );
not ( n34867 , n31599 );
or ( n34868 , n34866 , n34867 );
not ( n34869 , n379391 );
not ( n34870 , n31624 );
not ( n34871 , n34870 );
or ( n34872 , n34869 , n34871 );
nand ( n34873 , n34872 , n31700 );
and ( n34874 , n34873 , n31629 );
not ( n34875 , n31706 );
or ( n34876 , n34875 , n34870 , n31629 );
and ( n34877 , n379394 , RI15b57930_853);
and ( n34878 , n379398 , RI15b51738_644);
nor ( n34879 , n34877 , n34878 );
nand ( n34880 , n34876 , n34879 );
nor ( n34881 , n34874 , n34880 );
nand ( n34882 , n34868 , n34881 );
buf ( n34883 , n34882 );
buf ( n34884 , n379844 );
not ( n34885 , n385188 );
and ( n34886 , n34885 , RI15b60918_1160);
not ( n34887 , n379794 );
and ( n34888 , n34887 , RI15b5d768_1054);
nor ( n34889 , n34886 , n34888 );
not ( n34890 , n34889 );
buf ( n34891 , n34890 );
buf ( n34892 , n20665 );
not ( n34893 , n33611 );
or ( n34894 , n32430 , n34893 );
nand ( n34895 , n381417 , n381362 );
not ( n34896 , n382634 );
not ( n34897 , n34896 );
not ( n34898 , n382626 );
or ( n34899 , n34897 , n34898 );
nand ( n34900 , n34899 , n382679 );
and ( n34901 , n34900 , RI15b54a50_753);
or ( n34902 , n32458 , n34896 , RI15b54a50_753);
buf ( n34903 , n21391 );
not ( n34904 , n34903 );
not ( n34905 , n34904 );
buf ( n34906 , n34905 );
not ( n34907 , n34906 );
not ( n34908 , n34907 );
or ( n34909 , n382886 , n34908 );
nand ( n34910 , n34902 , n34909 );
nor ( n34911 , n34901 , n34910 );
and ( n34912 , n34895 , n34911 );
nand ( n34913 , n34894 , n34912 );
buf ( n34914 , n34913 );
buf ( n34915 , n380203 );
not ( n34916 , n32064 );
not ( n34917 , n381589 );
or ( n34918 , n34916 , n34917 );
and ( n34919 , n381596 , n32070 );
or ( n34920 , n32081 , n18717 );
or ( n34921 , n32420 , n32086 );
or ( n34922 , n32079 , n381621 );
nand ( n34923 , n34920 , n34921 , n34922 );
nor ( n34924 , n34919 , n34923 );
nand ( n34925 , n34918 , n34924 );
buf ( n34926 , n34925 );
buf ( n34927 , n22009 );
buf ( n34928 , n379847 );
buf ( n34929 , n22653 );
nand ( n34930 , n379825 , n385220 );
not ( n34931 , n34930 );
nor ( n34932 , n381953 , RI15b48b88_346);
nor ( n34933 , RI15b48c00_347 , RI15b48c78_348);
and ( n34934 , n34932 , n34933 );
not ( n34935 , RI15b48cf0_349);
and ( n34936 , n34934 , n34935 );
not ( n34937 , RI15b48d68_350);
nand ( n34938 , n34936 , n34937 );
nor ( n34939 , n34938 , RI15b48de0_351);
nor ( n34940 , RI15b48e58_352 , RI15b48ed0_353);
nand ( n34941 , n34939 , n34940 );
nand ( n34942 , n34941 , RI15b49308_362);
not ( n34943 , n34942 );
not ( n34944 , RI15b48f48_354);
and ( n34945 , n34943 , n34944 );
and ( n34946 , n34942 , RI15b48f48_354);
nor ( n34947 , n34945 , n34946 );
not ( n34948 , RI15b48e58_352);
not ( n34949 , n34948 );
not ( n34950 , n34939 );
or ( n34951 , n34949 , n34950 );
nand ( n34952 , n34951 , RI15b49308_362);
not ( n34953 , n34952 );
not ( n34954 , RI15b48ed0_353);
and ( n34955 , n34953 , n34954 );
and ( n34956 , n34952 , RI15b48ed0_353);
nor ( n34957 , n34955 , n34956 );
buf ( n34958 , n34932 );
nor ( n34959 , n34958 , n381954 );
not ( n34960 , RI15b48c00_347);
and ( n34961 , n34959 , n34960 );
not ( n34962 , n34959 );
and ( n34963 , n34962 , RI15b48c00_347);
nor ( n34964 , n34961 , n34963 );
nand ( n34965 , n34947 , n34957 , n34964 );
not ( n34966 , n34941 );
not ( n34967 , RI15b48f48_354);
and ( n34968 , n34966 , n34967 );
not ( n34969 , RI15b48fc0_355);
nor ( n34970 , n34968 , n34969 );
not ( n34971 , n34939 );
nor ( n34972 , n381954 , RI15b48e58_352);
and ( n34973 , n34971 , n34972 );
not ( n34974 , n34971 );
and ( n34975 , n34974 , RI15b48e58_352);
or ( n34976 , n34973 , n34975 );
and ( n34977 , n34958 , n34960 );
nor ( n34978 , n34977 , n381954 );
not ( n34979 , RI15b48c78_348);
not ( n34980 , RI15b48de0_351);
nand ( n34981 , n34979 , n34935 , n34980 , n34937 );
or ( n34982 , n34978 , n34981 );
nand ( n34983 , RI15b48d68_350 , RI15b48de0_351);
not ( n34984 , n34983 );
nand ( n34985 , n34978 , n34984 , RI15b48c78_348 , RI15b48cf0_349);
nand ( n34986 , n34982 , n34985 );
and ( n34987 , RI15b490b0_357 , RI15b49128_358 , RI15b49038_356 , RI15b49290_361);
nand ( n34988 , n34986 , n34987 , RI15b491a0_359 , RI15b49218_360);
nor ( n34989 , n34976 , n34988 );
nand ( n34990 , n34970 , n34989 );
or ( n34991 , n34965 , n34990 );
nand ( n34992 , n34991 , RI15b49308_362);
not ( n34993 , n34992 );
nand ( n34994 , n34993 , n34964 );
not ( n34995 , n34994 );
and ( n34996 , n34931 , n34995 );
nand ( n34997 , n34968 , n34969 );
nor ( n34998 , n34997 , RI15b49038_356);
not ( n34999 , RI15b490b0_357);
nand ( n35000 , n34998 , n34999 );
nor ( n35001 , n35000 , RI15b49128_358);
not ( n35002 , RI15b491a0_359);
nand ( n35003 , n35001 , n35002 );
and ( n35004 , n35003 , RI15b49218_360);
not ( n35005 , n35003 );
not ( n35006 , RI15b49218_360);
and ( n35007 , n35005 , n35006 );
nor ( n35008 , n35004 , n35007 );
not ( n35009 , n34992 );
buf ( n35010 , n35009 );
not ( n35011 , n35010 );
not ( n35012 , n35011 );
and ( n35013 , n35008 , n35012 );
nor ( n35014 , n35006 , RI15b49308_362);
nor ( n35015 , n35013 , n35014 );
not ( n35016 , n35010 );
not ( n35017 , n35000 );
and ( n35018 , n35017 , RI15b49128_358);
not ( n35019 , n35017 );
not ( n35020 , RI15b49128_358);
and ( n35021 , n35019 , n35020 );
nor ( n35022 , n35018 , n35021 );
or ( n35023 , n35016 , n35022 );
or ( n35024 , n35020 , RI15b49308_362);
nand ( n35025 , n35023 , n35024 );
not ( n35026 , n35010 );
not ( n35027 , RI15b49038_356);
and ( n35028 , n34997 , n35027 );
not ( n35029 , n34997 );
and ( n35030 , n35029 , RI15b49038_356);
nor ( n35031 , n35028 , n35030 );
or ( n35032 , n35026 , n35031 );
or ( n35033 , n35027 , RI15b49308_362);
nand ( n35034 , n35032 , n35033 );
nor ( n35035 , n35025 , n35034 );
not ( n35036 , n35001 );
and ( n35037 , n35036 , RI15b491a0_359);
not ( n35038 , n35036 );
and ( n35039 , n35038 , n35002 );
nor ( n35040 , n35037 , n35039 );
nand ( n35041 , n35040 , n35010 );
nand ( n35042 , n381954 , RI15b491a0_359);
and ( n35043 , n35041 , n35042 );
and ( n35044 , n35015 , n35035 , n35043 );
not ( n35045 , n35003 );
nand ( n35046 , n35045 , n35006 );
and ( n35047 , n35046 , RI15b49290_361);
not ( n35048 , n35046 );
not ( n35049 , RI15b49290_361);
and ( n35050 , n35048 , n35049 );
nor ( n35051 , n35047 , n35050 );
buf ( n35052 , n35012 );
and ( n35053 , n35051 , n35052 );
nor ( n35054 , n35049 , RI15b49308_362);
nor ( n35055 , n35053 , n35054 );
not ( n35056 , n34998 );
and ( n35057 , n35056 , RI15b490b0_357);
not ( n35058 , n35056 );
and ( n35059 , n35058 , n34999 );
nor ( n35060 , n35057 , n35059 );
nand ( n35061 , n35010 , n35060 );
nand ( n35062 , n381954 , RI15b490b0_357);
and ( n35063 , n35061 , n35062 );
not ( n35064 , n34970 );
nand ( n35065 , n35010 , n34997 , n35064 );
nand ( n35066 , n381954 , RI15b48fc0_355);
and ( n35067 , n35065 , n35066 );
buf ( n35068 , n35009 );
not ( n35069 , RI15b48de0_351);
not ( n35070 , n34938 );
not ( n35071 , n35070 );
or ( n35072 , n35069 , n35071 );
or ( n35073 , n35070 , RI15b48de0_351);
nand ( n35074 , n35072 , n35073 );
and ( n35075 , n35068 , n35074 );
nor ( n35076 , n34980 , RI15b49308_362);
nor ( n35077 , n35075 , n35076 );
not ( n35078 , RI15b48d68_350);
not ( n35079 , n34936 );
or ( n35080 , n35078 , n35079 );
or ( n35081 , n34936 , RI15b48d68_350);
nand ( n35082 , n35080 , n35081 );
not ( n35083 , n35082 );
not ( n35084 , n35009 );
or ( n35085 , n35083 , n35084 );
nand ( n35086 , n381954 , RI15b48d68_350);
nand ( n35087 , n35085 , n35086 );
not ( n35088 , n35087 );
and ( n35089 , n35063 , n35067 , n35077 , n35088 );
not ( n35090 , n34992 );
and ( n35091 , n34934 , RI15b48cf0_349);
not ( n35092 , n34934 );
and ( n35093 , n35092 , n34935 );
nor ( n35094 , n35091 , n35093 );
not ( n35095 , n35094 );
and ( n35096 , n35090 , n35095 );
and ( n35097 , n381954 , RI15b48cf0_349);
nor ( n35098 , n35096 , n35097 );
not ( n35099 , n34965 );
not ( n35100 , n34948 );
not ( n35101 , RI15b49308_362);
and ( n35102 , n35100 , n35101 );
nor ( n35103 , n35102 , n34976 );
not ( n35104 , n34978 );
and ( n35105 , n35104 , n34979 );
not ( n35106 , n35104 );
and ( n35107 , n35106 , RI15b48c78_348);
nor ( n35108 , n35105 , n35107 );
not ( n35109 , n35108 );
and ( n35110 , n35098 , n35099 , n35103 , n35109 );
nand ( n35111 , n35044 , n35055 , n35089 , n35110 );
buf ( n35112 , n35052 );
nand ( n35113 , n35111 , n35112 );
and ( n35114 , n35113 , n34931 );
nor ( n35115 , n34996 , n35114 );
or ( n35116 , n35115 , n35109 );
or ( n35117 , n35113 , n34930 );
not ( n35118 , n35117 );
nor ( n35119 , n34995 , n35108 );
and ( n35120 , n35118 , n35119 );
and ( n35121 , n20631 , RI15b460e0_255);
nor ( n35122 , n35120 , n35121 );
nand ( n35123 , n385213 , RI15b476e8_302);
nand ( n35124 , n35116 , n35122 , n35123 );
buf ( n35125 , n35124 );
buf ( n35126 , n385195 );
buf ( n35127 , n22404 );
buf ( n35128 , n385195 );
not ( n35129 , RI15b53c40_723);
not ( n35130 , n383170 );
or ( n35131 , n35129 , n35130 );
not ( n35132 , n383111 );
or ( n35133 , n35132 , n383152 );
nand ( n35134 , n35133 , n383157 );
not ( n35135 , n383095 );
and ( n35136 , n35134 , n35135 );
not ( n35137 , n35132 );
nor ( n35138 , n35137 , n35135 );
and ( n35139 , n35138 , n383143 );
and ( n35140 , n383147 , RI15b52638_676);
nor ( n35141 , n35136 , n35139 , n35140 );
nand ( n35142 , n35131 , n35141 );
buf ( n35143 , n35142 );
nand ( n35144 , n382974 , n380737 );
not ( n35145 , n35144 );
not ( n35146 , n35145 );
not ( n35147 , n382912 );
or ( n35148 , n35146 , n35147 );
nand ( n35149 , n382981 , n381493 );
not ( n35150 , n35149 );
and ( n35151 , n382931 , n35150 );
and ( n35152 , n35149 , n35144 , n32684 );
nor ( n35153 , n35152 , n19630 );
not ( n35154 , n33224 );
nor ( n35155 , n382988 , n35154 );
or ( n35156 , n35153 , n35155 );
nand ( n35157 , n35156 , n19595 );
or ( n35158 , n382992 , n380756 );
nand ( n35159 , n35157 , n35158 );
and ( n35160 , n35159 , n380775 );
or ( n35161 , n35160 , n19063 );
buf ( n35162 , n382957 );
not ( n35163 , n35162 );
not ( n35164 , n35158 );
nor ( n35165 , n35155 , n35164 );
or ( n35166 , n35153 , n35165 );
or ( n35167 , n35163 , n35166 );
or ( n35168 , n35158 , n382967 );
nand ( n35169 , n35161 , n35167 , n35168 );
nor ( n35170 , n35151 , n35169 );
nand ( n35171 , n35148 , n35170 );
buf ( n35172 , n35171 );
buf ( n35173 , n382537 );
buf ( n35174 , n382067 );
not ( n35175 , RI15b659b8_1332);
nand ( n35176 , n379821 , n386547 );
not ( n35177 , n35176 );
or ( n35178 , n35175 , n35177 );
nand ( n35179 , n379835 , n22278 );
or ( n35180 , n381031 , n385201 );
and ( n35181 , n381035 , n386530 );
nand ( n35182 , n381039 , n20501 );
nor ( n35183 , n35181 , n35182 , n381073 );
nand ( n35184 , n35180 , n381050 , n35183 );
nor ( n35185 , n385202 , n379818 );
or ( n35186 , n35184 , n35185 );
buf ( n35187 , n35186 );
nand ( n35188 , n35187 , RI15b485e8_334);
buf ( n35189 , n385756 );
not ( n35190 , n35189 );
buf ( n35191 , n35190 );
not ( n35192 , n35191 );
and ( n35193 , n386554 , n35192 );
buf ( n35194 , n386510 );
not ( n35195 , n35194 );
not ( n35196 , n35195 );
not ( n35197 , RI15b485e8_334);
nand ( n35198 , RI15b48480_331 , RI15b484f8_332);
not ( n35199 , RI15b48570_333);
nor ( n35200 , n35198 , n35199 );
not ( n35201 , n35200 );
not ( n35202 , n35201 );
or ( n35203 , n35197 , n35202 );
or ( n35204 , n35201 , RI15b485e8_334);
nand ( n35205 , n35203 , n35204 );
and ( n35206 , n35196 , n35205 );
nor ( n35207 , n35193 , n35206 );
and ( n35208 , n35179 , n35188 , n35207 );
nand ( n35209 , n35178 , n35208 );
buf ( n35210 , n35209 );
buf ( n35211 , n381490 );
buf ( n35212 , n32672 );
not ( n35213 , n381014 );
not ( n35214 , RI15b45f78_252);
nor ( n35215 , n35214 , RI15b45e88_250 , RI15b45f00_251 , RI15b45ff0_253);
nor ( n35216 , RI15b44e98_216 , RI15b44f10_217 , RI15b44f88_218 , RI15b45000_219);
nand ( n35217 , n35213 , n35215 , n35216 );
buf ( n35218 , n35217 );
buf ( n35219 , n30992 );
buf ( n35220 , n22655 );
or ( n35221 , n386588 , n32681 );
not ( n35222 , n32683 );
and ( n35223 , n386600 , n35222 );
not ( n35224 , RI15b5a630_949);
or ( n35225 , n32692 , n35224 );
or ( n35226 , n34706 , n32699 );
or ( n35227 , n32690 , n386627 );
nand ( n35228 , n35225 , n35226 , n35227 );
nor ( n35229 , n35223 , n35228 );
nand ( n35230 , n35221 , n35229 );
buf ( n35231 , n35230 );
buf ( n35232 , n31719 );
nor ( n35233 , RI15b54780_747 , RI15b547f8_748);
nand ( n35234 , n35233 , RI15b54870_749);
or ( n35235 , n35234 , RI15b3fa38_36);
nand ( n35236 , RI15b3f9c0_35 , RI15b54870_749);
or ( n35237 , n35236 , n35233 );
or ( n35238 , n385032 , n18094 , RI15b547f8_748 , RI15b54258_736);
nand ( n35239 , n35235 , n35237 , n35238 );
or ( n35240 , RI15b3f9c0_35 , RI15b54258_736);
not ( n35241 , RI15b3fa38_36);
nand ( n35242 , n35240 , n35241 , RI15b54780_747);
and ( n35243 , n35242 , n379339 );
not ( n35244 , n18072 );
nand ( n35245 , n35244 , RI15b547f8_748);
nor ( n35246 , n35243 , n35245 );
or ( n35247 , n35239 , n35246 , n379391 );
buf ( n35248 , n35247 );
buf ( n35249 , n382065 );
not ( n35250 , n384518 );
not ( n35251 , n384523 );
and ( n35252 , n387116 , n35251 );
not ( n35253 , n35252 );
or ( n35254 , n35250 , n35253 );
or ( n35255 , n35252 , n384518 );
nand ( n35256 , n35254 , n35255 );
and ( n35257 , n35256 , n31959 );
not ( n35258 , n384392 );
not ( n35259 , n387129 );
or ( n35260 , n35259 , n384295 );
not ( n35261 , n32537 );
nand ( n35262 , n35260 , n35261 );
not ( n35263 , n35262 );
or ( n35264 , n35258 , n35263 );
not ( n35265 , n384416 );
not ( n35266 , n35265 );
nand ( n35267 , n387138 , n384421 );
not ( n35268 , n35267 );
not ( n35269 , n35268 );
or ( n35270 , n35266 , n35269 );
or ( n35271 , n35268 , n35265 );
nand ( n35272 , n35270 , n35271 );
buf ( n35273 , n384493 );
and ( n35274 , n35272 , n35273 );
and ( n35275 , n19513 , RI15b63f78_1276);
nor ( n35276 , n35274 , n35275 );
nand ( n35277 , n35264 , n35276 );
nor ( n35278 , n35257 , n35277 );
and ( n35279 , n19608 , RI15b63078_1244);
not ( n35280 , n386831 );
and ( n35281 , n35280 , n19630 );
not ( n35282 , n386826 );
and ( n35283 , n35282 , n383446 );
not ( n35284 , n35282 );
and ( n35285 , n35284 , RI15b63078_1244);
nor ( n35286 , n35283 , n35285 );
and ( n35287 , n35286 , n31964 );
nor ( n35288 , n35279 , n35281 , n35287 );
nand ( n35289 , n35278 , n35288 );
buf ( n35290 , n35289 );
buf ( n35291 , n386563 );
buf ( n35292 , n22738 );
buf ( n35293 , n19919 );
not ( n35294 , n35293 );
not ( n35295 , n35294 );
not ( n35296 , n19898 );
or ( n35297 , n35295 , n35296 );
nand ( n35298 , n35297 , n19940 );
nand ( n35299 , n35298 , n19715 );
buf ( n35300 , n19996 );
nor ( n35301 , n35300 , n20502 );
or ( n35302 , n35301 , n20521 );
nand ( n35303 , n35302 , RI15b4a028_390);
not ( n35304 , n19898 );
not ( n35305 , n22368 );
nor ( n35306 , n35305 , n19715 );
nand ( n35307 , n35304 , n35306 );
nor ( n35308 , n20529 , RI15b4a028_390);
and ( n35309 , n35300 , n35308 );
not ( n35310 , n20557 );
and ( n35311 , n20646 , n35310 );
nor ( n35312 , n35311 , n20641 );
or ( n35313 , n35312 , n382143 );
or ( n35314 , n35310 , n382135 , RI15b4be28_454);
or ( n35315 , n382143 , RI15b4bdb0_453);
nand ( n35316 , n35314 , n35315 );
and ( n35317 , n20646 , n35316 );
and ( n35318 , n32620 , RI15b4af28_422);
nor ( n35319 , n35317 , n35318 );
nand ( n35320 , n35313 , n35319 );
nor ( n35321 , n35309 , n35320 );
nand ( n35322 , n35299 , n35303 , n35307 , n35321 );
buf ( n35323 , n35322 );
buf ( n35324 , n382537 );
buf ( n35325 , n22714 );
or ( n35326 , n381015 , n22037 );
not ( n35327 , n35213 );
nand ( n35328 , n35327 , RI15b53b50_721);
nand ( n35329 , n35326 , n35328 );
buf ( n35330 , n35329 );
buf ( n35331 , n22740 );
buf ( n35332 , n32672 );
not ( n35333 , n35187 );
or ( n35334 , n35333 , n34948 );
not ( n35335 , n386547 );
and ( n35336 , n35335 , RI15b66228_1350);
not ( n35337 , n34948 );
nand ( n35338 , n35200 , RI15b485e8_334);
not ( n35339 , RI15b48660_335);
nor ( n35340 , n35338 , n35339 );
nand ( n35341 , n35340 , RI15b486d8_336);
not ( n35342 , n35341 );
nand ( n35343 , n35342 , RI15b48750_337);
not ( n35344 , n35343 );
and ( n35345 , n35344 , RI15b487c8_338);
nand ( n35346 , n35345 , RI15b48840_339);
not ( n35347 , RI15b488b8_340);
nor ( n35348 , n35346 , n35347 );
and ( n35349 , n35348 , RI15b48930_341);
and ( n35350 , n35349 , RI15b489a8_342);
nand ( n35351 , n35350 , RI15b48a20_343);
nand ( n35352 , RI15b48a98_344 , RI15b48b10_345);
nor ( n35353 , n35351 , n35352 );
and ( n35354 , n35353 , RI15b48b88_346);
nand ( n35355 , n35354 , RI15b48c00_347);
nor ( n35356 , n35355 , n34979 );
nand ( n35357 , n35356 , RI15b48cf0_349);
nor ( n35358 , n35357 , n34983 );
not ( n35359 , n35358 );
or ( n35360 , n35337 , n35359 );
or ( n35361 , n35358 , n34948 );
nand ( n35362 , n35360 , n35361 );
buf ( n35363 , n35194 );
and ( n35364 , n35362 , n35363 );
not ( n35365 , n20055 );
not ( n35366 , n385998 );
or ( n35367 , n35365 , n35366 );
not ( n35368 , n383374 );
nand ( n35369 , n385471 , n35368 );
nand ( n35370 , n35367 , n35369 );
nand ( n35371 , n381046 , n35370 );
not ( n35372 , n32779 );
nor ( n35373 , n35371 , n35372 );
and ( n35374 , n35373 , RI15b435c0_163);
not ( n35375 , n35371 );
and ( n35376 , n35375 , n32784 );
and ( n35377 , n35376 , RI15b43980_171);
not ( n35378 , n385263 );
not ( n35379 , n35378 );
not ( n35380 , n35379 );
or ( n35381 , n35371 , n35380 );
or ( n35382 , n35381 , n20337 );
not ( n35383 , n32745 );
nor ( n35384 , n35371 , n35383 );
not ( n35385 , n35384 );
or ( n35386 , n20334 , n35385 );
not ( n35387 , n381046 );
not ( n35388 , n32729 );
and ( n35389 , n35379 , n35388 );
not ( n35390 , n35389 );
nor ( n35391 , n35387 , n35390 );
and ( n35392 , n35391 , RI15b42300_123);
not ( n35393 , n385344 );
buf ( n35394 , n35393 );
buf ( n35395 , n35394 );
buf ( n35396 , n35395 );
and ( n35397 , n35396 , RI15b426c0_131);
nand ( n35398 , n385989 , n35368 );
not ( n35399 , n35398 );
buf ( n35400 , n35399 );
buf ( n35401 , n35400 );
and ( n35402 , n35401 , RI15b40140_51);
not ( n35403 , n385992 );
not ( n35404 , n383374 );
and ( n35405 , n35403 , n35404 );
buf ( n35406 , n35405 );
buf ( n35407 , n35406 );
and ( n35408 , n35407 , RI15b40500_59);
nor ( n35409 , n35397 , n35402 , n35408 );
not ( n35410 , n20110 );
and ( n35411 , n35410 , RI15b40c80_75);
not ( n35412 , n20019 );
and ( n35413 , n35412 , RI15b41f40_115);
nor ( n35414 , n35411 , n35413 );
not ( n35415 , n20092 );
and ( n35416 , n35415 , RI15b42a80_139);
and ( n35417 , n383378 , RI15b408c0_67);
nor ( n35418 , n35416 , n35417 );
and ( n35419 , n35409 , n35414 , n35418 );
nor ( n35420 , n35419 , n381060 );
nor ( n35421 , n35392 , n35420 );
not ( n35422 , n20026 );
nand ( n35423 , n381046 , n35422 );
not ( n35424 , n35423 );
not ( n35425 , n385457 );
and ( n35426 , n35424 , n35425 );
buf ( n35427 , n20098 );
buf ( n35428 , n35427 );
buf ( n35429 , n35428 );
buf ( n35430 , n35429 );
not ( n35431 , n35430 );
not ( n35432 , n35431 );
nand ( n35433 , n381046 , n35432 );
nor ( n35434 , n35433 , n385452 );
nor ( n35435 , n35426 , n35434 );
not ( n35436 , n20105 );
buf ( n35437 , n35436 );
buf ( n35438 , n35437 );
buf ( n35439 , n35438 );
not ( n35440 , n35439 );
not ( n35441 , n35440 );
nand ( n35442 , n381046 , n35441 );
not ( n35443 , n35442 );
not ( n35444 , RI15b41040_83);
not ( n35445 , n35444 );
and ( n35446 , n35443 , n35445 );
not ( n35447 , n35378 );
and ( n35448 , n35447 , n20104 );
nand ( n35449 , n381046 , n35448 );
nor ( n35450 , n35449 , n20363 );
nor ( n35451 , n35446 , n35450 );
and ( n35452 , n35421 , n35435 , n35451 );
nand ( n35453 , n35382 , n35386 , n35452 );
nor ( n35454 , n35374 , n35377 , n35453 );
buf ( n35455 , n381036 );
buf ( n35456 , n35455 );
nor ( n35457 , n35454 , n35456 );
nor ( n35458 , n35336 , n35364 , n35457 );
and ( n35459 , n379820 , n22254 );
and ( n35460 , n35459 , n22252 );
and ( n35461 , n379820 , RI15b666d8_1360);
and ( n35462 , n35461 , RI15b65aa8_1334);
nor ( n35463 , n35460 , n35462 );
nand ( n35464 , n35334 , n35458 , n35463 );
buf ( n35465 , n35464 );
buf ( n35466 , n19655 );
buf ( n35467 , n381021 );
buf ( n35468 , n31030 );
buf ( n35469 , n383867 );
not ( n35470 , n35469 );
buf ( n35471 , n35470 );
not ( n35472 , n35471 );
not ( n35473 , n35472 );
not ( n35474 , n35473 );
not ( n35475 , n384726 );
or ( n35476 , n35474 , n35475 );
not ( n35477 , n384736 );
and ( n35478 , n383875 , n384055 );
and ( n35479 , n384165 , n35478 );
and ( n35480 , n35477 , n35479 );
not ( n35481 , n35479 );
and ( n35482 , n35481 , n35469 , n384741 );
nor ( n35483 , n35482 , n21764 );
or ( n35484 , n35483 , n383833 );
nand ( n35485 , n35484 , n18154 );
nand ( n35486 , n383819 , n384178 );
and ( n35487 , n35485 , n35486 );
nor ( n35488 , n35487 , n383902 );
or ( n35489 , n35488 , n20737 );
not ( n35490 , n384752 );
not ( n35491 , n35490 );
not ( n35492 , n383833 );
not ( n35493 , n35486 );
not ( n35494 , n35493 );
and ( n35495 , n35492 , n35494 );
nor ( n35496 , n35495 , n35483 );
not ( n35497 , n35496 );
or ( n35498 , n35491 , n35497 );
or ( n35499 , n35486 , n384759 );
nand ( n35500 , n35489 , n35498 , n35499 );
nor ( n35501 , n35480 , n35500 );
nand ( n35502 , n35476 , n35501 );
buf ( n35503 , n35502 );
buf ( n35504 , n379403 );
not ( n35505 , RI15b60dc8_1170);
or ( n35506 , n31091 , n35505 );
buf ( n35507 , n31777 );
and ( n35508 , n35507 , n18630 );
buf ( n35509 , n383588 );
not ( n35510 , n35509 );
or ( n35511 , n35510 , n384904 , n386616 );
not ( n35512 , n31078 );
and ( n35513 , n35505 , RI15b60d50_1169);
not ( n35514 , RI15b60d50_1169);
and ( n35515 , n35514 , RI15b60dc8_1170);
nor ( n35516 , n35513 , n35515 );
or ( n35517 , n35512 , n35516 );
nand ( n35518 , n35511 , n35517 );
nor ( n35519 , n35508 , n35518 );
nand ( n35520 , n35506 , n35519 );
buf ( n35521 , n35520 );
buf ( n35522 , n22653 );
not ( n35523 , n35213 );
or ( n35524 , n35523 , n22047 );
buf ( n35525 , n381014 );
nand ( n35526 , n35525 , RI15b53da8_726);
nand ( n35527 , n35524 , n35526 );
buf ( n35528 , n35527 );
buf ( n35529 , n381707 );
buf ( n35530 , n382067 );
buf ( n35531 , n386762 );
not ( n35532 , n35187 );
or ( n35533 , n35532 , n34960 );
buf ( n35534 , n35456 );
and ( n35535 , n35373 , RI15b43368_158);
and ( n35536 , n35376 , RI15b43728_166);
not ( n35537 , n35381 );
and ( n35538 , n35537 , RI15b42fa8_150);
and ( n35539 , n35384 , RI15b42be8_142);
nor ( n35540 , n35538 , n35539 );
not ( n35541 , n35449 );
and ( n35542 , n35541 , RI15b411a8_86);
not ( n35543 , n35442 );
and ( n35544 , n35543 , RI15b40de8_78);
nor ( n35545 , n35542 , n35544 );
not ( n35546 , n35423 );
and ( n35547 , n35546 , RI15b41928_102);
not ( n35548 , n35433 );
and ( n35549 , n35548 , RI15b41568_94);
nor ( n35550 , n35547 , n35549 );
and ( n35551 , n35391 , RI15b420a8_118);
buf ( n35552 , n35407 );
buf ( n35553 , n35552 );
and ( n35554 , n35553 , RI15b402a8_54);
buf ( n35555 , n35396 );
and ( n35556 , n35555 , RI15b42468_126);
buf ( n35557 , n35401 );
and ( n35558 , n35557 , RI15b3fee8_46);
nor ( n35559 , n35554 , n35556 , n35558 );
and ( n35560 , n35410 , RI15b40a28_70);
and ( n35561 , n35412 , RI15b41ce8_110);
nor ( n35562 , n35560 , n35561 );
and ( n35563 , n35415 , RI15b42828_134);
and ( n35564 , n383379 , RI15b40668_62);
nor ( n35565 , n35563 , n35564 );
and ( n35566 , n35559 , n35562 , n35565 );
not ( n35567 , n386530 );
not ( n35568 , n35567 );
nor ( n35569 , n35566 , n35568 );
nor ( n35570 , n35551 , n35569 );
nand ( n35571 , n35540 , n35545 , n35550 , n35570 );
nor ( n35572 , n35535 , n35536 , n35571 );
or ( n35573 , n35534 , n35572 );
and ( n35574 , n35335 , RI15b65fd0_1345);
not ( n35575 , n34960 );
not ( n35576 , n35354 );
or ( n35577 , n35575 , n35576 );
or ( n35578 , n35354 , n34960 );
nand ( n35579 , n35577 , n35578 );
not ( n35580 , n35195 );
and ( n35581 , n35579 , n35580 );
not ( n35582 , RI15b65850_1329);
nor ( n35583 , n379819 , n35582 );
nor ( n35584 , n35574 , n35581 , n35583 );
nand ( n35585 , n35533 , n35573 , n35584 );
buf ( n35586 , n35585 );
buf ( n35587 , n381081 );
not ( n35588 , RI15b65aa8_1334);
not ( n35589 , n35176 );
or ( n35590 , n35588 , n35589 );
nand ( n35591 , n379835 , n22252 );
nand ( n35592 , n35187 , RI15b486d8_336);
buf ( n35593 , n385493 );
buf ( n35594 , n35593 );
and ( n35595 , n386554 , n35594 );
not ( n35596 , RI15b486d8_336);
not ( n35597 , n35340 );
not ( n35598 , n35597 );
or ( n35599 , n35596 , n35598 );
or ( n35600 , n35597 , RI15b486d8_336);
nand ( n35601 , n35599 , n35600 );
and ( n35602 , n35196 , n35601 );
nor ( n35603 , n35595 , n35602 );
and ( n35604 , n35591 , n35592 , n35603 );
nand ( n35605 , n35590 , n35604 );
buf ( n35606 , n35605 );
buf ( n35607 , n380906 );
buf ( n35608 , n19655 );
buf ( n35609 , n32255 );
buf ( n35610 , n31719 );
not ( n35611 , n32244 );
buf ( n35612 , n35611 );
buf ( n35613 , n380942 );
not ( n35614 , RI15b5f9a0_1127);
not ( n35615 , n383601 );
or ( n35616 , n35614 , n35615 );
and ( n35617 , n383505 , RI15b60f30_1173);
and ( n35618 , n383607 , RI15b5f220_1111);
nor ( n35619 , n35617 , n35618 );
nand ( n35620 , n35616 , n35619 );
buf ( n35621 , n35620 );
or ( n35622 , n384703 , n383886 );
or ( n35623 , n31149 , n35622 );
nand ( n35624 , n383876 , n21337 );
not ( n35625 , n35624 );
and ( n35626 , n31161 , n35625 );
and ( n35627 , n35624 , n35622 , n384741 );
nor ( n35628 , n35627 , n21764 );
buf ( n35629 , n33122 );
nor ( n35630 , n383885 , n35629 );
or ( n35631 , n35628 , n35630 );
nand ( n35632 , n35631 , n18154 );
or ( n35633 , n383893 , n383865 );
nand ( n35634 , n35632 , n35633 );
and ( n35635 , n35634 , n383901 );
not ( n35636 , RI15b4f500_571);
or ( n35637 , n35635 , n35636 );
not ( n35638 , n35633 );
nor ( n35639 , n35630 , n35638 );
or ( n35640 , n35628 , n35639 );
or ( n35641 , n31179 , n35640 );
or ( n35642 , n35633 , n31184 );
nand ( n35643 , n35637 , n35641 , n35642 );
nor ( n35644 , n35626 , n35643 );
nand ( n35645 , n35623 , n35644 );
buf ( n35646 , n35645 );
buf ( n35647 , n30992 );
buf ( n35648 , n379893 );
buf ( n35649 , RI15b3ea48_2);
buf ( n35650 , n35649 );
buf ( n35651 , RI15b3ea48_2);
buf ( n35652 , n35651 );
buf ( n35653 , n381566 );
buf ( n35654 , n386762 );
not ( n35655 , RI15b47328_294);
not ( n35656 , n385213 );
or ( n35657 , n35655 , n35656 );
and ( n35658 , n385221 , RI15b488b8_340);
and ( n35659 , n20631 , RI15b46ba8_278);
nor ( n35660 , n35658 , n35659 );
nand ( n35661 , n35657 , n35660 );
buf ( n35662 , n35661 );
buf ( n35663 , n386760 );
and ( n35664 , n22646 , RI15b45a50_241);
and ( n35665 , n22648 , RI15b51eb8_660);
nor ( n35666 , n35664 , n35665 );
not ( n35667 , n35666 );
buf ( n35668 , n35667 );
buf ( n35669 , n384218 );
buf ( n35670 , n22005 );
and ( n35671 , n381525 , n32068 );
not ( n35672 , n32069 );
nor ( n35673 , n35671 , n35672 );
not ( n35674 , n19642 );
or ( n35675 , n35673 , n35674 );
or ( n35676 , n22775 , n382896 );
buf ( n35677 , n18858 );
and ( n35678 , n19257 , n35677 );
nor ( n35679 , n35678 , n19594 , RI15b5d498_1048);
not ( n35680 , n19594 );
and ( n35681 , n35680 , RI15b584e8_878);
nor ( n35682 , n35679 , n35681 );
or ( n35683 , n35682 , RI15b584e8_878);
nand ( n35684 , n35683 , n380774 );
and ( n35685 , n35684 , RI15b586c8_882);
and ( n35686 , n380789 , n380211 );
nor ( n35687 , n35685 , n35686 );
nand ( n35688 , n35675 , n35676 , n35687 );
buf ( n35689 , n35688 );
not ( n35690 , n21742 );
not ( n35691 , n21607 );
buf ( n35692 , n21399 );
and ( n35693 , n35692 , n21414 );
not ( n35694 , n35693 );
and ( n35695 , n35691 , n35694 );
and ( n35696 , n21607 , n35693 );
nor ( n35697 , n35695 , n35696 );
or ( n35698 , n35690 , n35697 );
not ( n35699 , n32456 );
and ( n35700 , n35699 , n21097 );
and ( n35701 , n32456 , n21096 );
nor ( n35702 , n35700 , n35701 );
not ( n35703 , n35702 );
buf ( n35704 , n21206 );
buf ( n35705 , n35704 );
not ( n35706 , n35705 );
or ( n35707 , n35703 , n35706 );
or ( n35708 , n35705 , n35702 );
nand ( n35709 , n35707 , n35708 );
and ( n35710 , n21353 , n35709 );
not ( n35711 , n35693 );
not ( n35712 , n21410 );
not ( n35713 , n35712 );
or ( n35714 , n35711 , n35713 );
or ( n35715 , n35693 , n35712 );
nand ( n35716 , n35714 , n35715 );
and ( n35717 , n21558 , n35716 );
and ( n35718 , n21751 , RI15b576d8_848);
nor ( n35719 , n35710 , n35717 , n35718 );
nand ( n35720 , n35698 , n35719 );
or ( n35721 , n21789 , n379901 );
and ( n35722 , n21766 , n379908 );
and ( n35723 , n383854 , n379901 );
nor ( n35724 , n35722 , n35723 );
nand ( n35725 , n35721 , n35724 );
or ( n35726 , n35720 , n35725 );
buf ( n35727 , n35726 );
or ( n35728 , n382679 , n383022 );
not ( n35729 , n386668 );
not ( n35730 , n35729 );
not ( n35731 , n21556 );
nor ( n35732 , n35731 , n382863 );
and ( n35733 , n35732 , RI15b4c968_478);
and ( n35734 , n379990 , n380128 );
and ( n35735 , n35734 , RI15b4fde8_590);
buf ( n35736 , n379991 );
and ( n35737 , n380061 , RI15b4eee8_558);
and ( n35738 , n382841 , RI15b4dc28_518);
not ( n35739 , n380132 );
and ( n35740 , n35739 , RI15b4d4a8_502);
nor ( n35741 , n35737 , n35738 , n35740 );
and ( n35742 , n382838 , RI15b4dfe8_526);
and ( n35743 , n382856 , RI15b4eb28_550);
nor ( n35744 , n35742 , n35743 );
and ( n35745 , n382826 , RI15b4d868_510);
and ( n35746 , n382849 , RI15b4e768_542);
nor ( n35747 , n35745 , n35746 );
not ( n35748 , n380102 );
nand ( n35749 , n35748 , RI15b4e3a8_534);
nand ( n35750 , n35741 , n35744 , n35747 , n35749 );
and ( n35751 , n35736 , n35750 );
nor ( n35752 , n35733 , n35735 , n35751 );
not ( n35753 , n382540 );
and ( n35754 , n35753 , n380123 );
and ( n35755 , n35754 , RI15b4f668_574);
and ( n35756 , n382541 , n380125 );
and ( n35757 , n35756 , RI15b4fa28_582);
nor ( n35758 , n35755 , n35757 );
and ( n35759 , n21556 , n380099 );
and ( n35760 , n35759 , RI15b4f2a8_566);
and ( n35761 , n35753 , n380115 );
and ( n35762 , n35761 , RI15b4c5a8_470);
nor ( n35763 , n35760 , n35762 );
and ( n35764 , n379991 , n382834 );
and ( n35765 , n35764 , RI15b4d0e8_494);
and ( n35766 , n379991 , n379879 );
and ( n35767 , n35766 , RI15b4cd28_486);
nor ( n35768 , n35765 , n35767 );
and ( n35769 , n35752 , n35758 , n35763 , n35768 );
or ( n35770 , n35730 , n35769 );
and ( n35771 , n382659 , n383022 );
not ( n35772 , n382659 );
and ( n35773 , n35772 , RI15b552c0_771);
nor ( n35774 , n35771 , n35773 );
and ( n35775 , n35774 , n382626 );
buf ( n35776 , n381339 );
not ( n35777 , n35776 );
nor ( n35778 , n381400 , n35777 );
nor ( n35779 , n382691 , n383651 );
nor ( n35780 , n35775 , n35778 , n35779 );
nand ( n35781 , n35728 , n35770 , n35780 );
buf ( n35782 , n35781 );
not ( n35783 , n380756 );
and ( n35784 , n386589 , n35783 );
not ( n35785 , n35784 );
not ( n35786 , n382912 );
or ( n35787 , n35785 , n35786 );
not ( n35788 , n381541 );
nand ( n35789 , n382932 , n35788 );
not ( n35790 , n35789 );
and ( n35791 , n382931 , n35790 );
not ( n35792 , n35784 );
and ( n35793 , n35789 , n35792 , n382937 );
nor ( n35794 , n35793 , n19630 );
not ( n35795 , n33230 );
not ( n35796 , n35795 );
not ( n35797 , n35796 );
nor ( n35798 , n382940 , n35797 );
or ( n35799 , n35794 , n35798 );
nand ( n35800 , n35799 , n19595 );
or ( n35801 , n382945 , n380728 );
nand ( n35802 , n35800 , n35801 );
and ( n35803 , n35802 , n380775 );
or ( n35804 , n35803 , n18513 );
not ( n35805 , n382958 );
not ( n35806 , n35798 );
not ( n35807 , n35801 );
not ( n35808 , n35807 );
and ( n35809 , n35806 , n35808 );
nor ( n35810 , n35809 , n35794 );
not ( n35811 , n35810 );
or ( n35812 , n35805 , n35811 );
or ( n35813 , n35801 , n382967 );
nand ( n35814 , n35804 , n35812 , n35813 );
nor ( n35815 , n35791 , n35814 );
nand ( n35816 , n35787 , n35815 );
buf ( n35817 , n35816 );
buf ( n35818 , n380940 );
buf ( n35819 , n22009 );
buf ( n35820 , n22408 );
buf ( n35821 , n22005 );
buf ( n35822 , n385112 );
or ( n35823 , n22315 , n32165 );
and ( n35824 , n22326 , n32170 );
not ( n35825 , RI15b434d0_161);
or ( n35826 , n32183 , n35825 );
or ( n35827 , n22334 , n32187 );
or ( n35828 , n32181 , n22336 );
nand ( n35829 , n35826 , n35827 , n35828 );
nor ( n35830 , n35824 , n35829 );
nand ( n35831 , n35823 , n35830 );
buf ( n35832 , n35831 );
buf ( n35833 , n382069 );
buf ( n35834 , n386563 );
buf ( n35835 , n18226 );
buf ( n35836 , n382069 );
not ( n35837 , n32121 );
not ( n35838 , n33173 );
not ( n35839 , n35838 );
or ( n35840 , n35837 , n35839 );
and ( n35841 , n33196 , n22211 );
not ( n35842 , RI15b409b0_69);
or ( n35843 , n22237 , n35842 );
or ( n35844 , n22241 , n22296 );
or ( n35845 , n22228 , n33201 );
nand ( n35846 , n35843 , n35844 , n35845 );
nor ( n35847 , n35841 , n35846 );
nand ( n35848 , n35840 , n35847 );
buf ( n35849 , n35848 );
not ( n35850 , n20638 );
not ( n35851 , n381899 );
nand ( n35852 , n35850 , n35851 );
or ( n35853 , n35852 , n22151 );
and ( n35854 , n381909 , RI15b40668_62);
or ( n35855 , n35582 , n22296 );
or ( n35856 , n20576 , n22298 );
or ( n35857 , n35856 , n22228 );
or ( n35858 , n22175 , n20638 );
or ( n35859 , n22213 , n35858 );
nand ( n35860 , n35855 , n35857 , n35859 );
nor ( n35861 , n35854 , n35860 );
nand ( n35862 , n35853 , n35861 );
buf ( n35863 , n35862 );
buf ( n35864 , n384218 );
buf ( n35865 , n381707 );
buf ( n35866 , n379895 );
buf ( n35867 , n386563 );
buf ( n35868 , n384996 );
or ( n35869 , n22149 , n380925 );
or ( n35870 , n32259 , n35869 );
nand ( n35871 , n22208 , n22134 );
not ( n35872 , n35871 );
and ( n35873 , n384983 , n35872 );
and ( n35874 , n35869 , n35871 , n19912 );
nor ( n35875 , n35874 , n22217 );
not ( n35876 , n32180 );
not ( n35877 , n35876 );
buf ( n35878 , n35877 );
nor ( n35879 , n22219 , n35878 );
or ( n35880 , n35875 , n35879 );
nand ( n35881 , n35880 , n20623 );
or ( n35882 , n22224 , n22150 );
and ( n35883 , n35881 , n35882 );
nor ( n35884 , n35883 , n22236 );
or ( n35885 , n35884 , n385381 );
not ( n35886 , n35882 );
nor ( n35887 , n35879 , n35886 );
or ( n35888 , n35875 , n35887 );
or ( n35889 , n22022 , n35888 );
or ( n35890 , n35882 , n384988 );
nand ( n35891 , n35885 , n35889 , n35890 );
nor ( n35892 , n35873 , n35891 );
nand ( n35893 , n35870 , n35892 );
buf ( n35894 , n35893 );
or ( n35895 , n22149 , n32180 );
not ( n35896 , n35895 );
not ( n35897 , n35896 );
not ( n35898 , n32129 );
or ( n35899 , n35897 , n35898 );
nand ( n35900 , n22208 , n32164 );
and ( n35901 , n35895 , n35900 , n19912 );
nor ( n35902 , n35901 , n22217 );
buf ( n35903 , n22210 );
buf ( n35904 , n35903 );
not ( n35905 , n35904 );
nor ( n35906 , n22219 , n35905 );
or ( n35907 , n35902 , n35906 );
nand ( n35908 , n35907 , n20623 );
or ( n35909 , n22224 , n22133 );
and ( n35910 , n35908 , n35909 );
nor ( n35911 , n35910 , n22236 );
not ( n35912 , n35911 );
and ( n35913 , n35912 , RI15b40320_55);
or ( n35914 , n32141 , n35900 );
not ( n35915 , n35909 );
nor ( n35916 , n35906 , n35915 );
or ( n35917 , n35902 , n35916 );
or ( n35918 , n32148 , n35917 );
or ( n35919 , n35909 , n32150 );
nand ( n35920 , n35914 , n35918 , n35919 );
nor ( n35921 , n35913 , n35920 );
nand ( n35922 , n35899 , n35921 );
buf ( n35923 , n35922 );
buf ( n35924 , n381006 );
buf ( n35925 , n379802 );
buf ( n35926 , n30992 );
buf ( n35927 , n384203 );
buf ( n35928 , n384218 );
nand ( n35929 , n22143 , n22147 );
or ( n35930 , n35929 , n22133 );
or ( n35931 , n380968 , n35930 );
not ( n35932 , n380911 );
not ( n35933 , n22130 );
nand ( n35934 , n35932 , n35933 );
not ( n35935 , n35934 );
and ( n35936 , n380986 , n35935 );
and ( n35937 , n35930 , n35934 , n19912 );
nor ( n35938 , n35937 , n22217 );
buf ( n35939 , n22116 );
nor ( n35940 , n35939 , n380919 );
or ( n35941 , n35938 , n35940 );
nand ( n35942 , n35941 , n20623 );
nand ( n35943 , n22223 , RI15b3fd80_43);
or ( n35944 , n35943 , n380925 );
and ( n35945 , n35942 , n35944 );
nor ( n35946 , n35945 , n22236 );
or ( n35947 , n35946 , n35444 );
not ( n35948 , n35944 );
nor ( n35949 , n35940 , n35948 );
or ( n35950 , n35938 , n35949 );
or ( n35951 , n380994 , n35950 );
or ( n35952 , n35944 , n380996 );
nand ( n35953 , n35947 , n35951 , n35952 );
nor ( n35954 , n35936 , n35953 );
nand ( n35955 , n35931 , n35954 );
buf ( n35956 , n35955 );
or ( n35957 , n22149 , n22133 );
or ( n35958 , n381907 , n35957 );
nand ( n35959 , n35932 , n380912 );
and ( n35960 , n35957 , n35959 , n19912 );
nor ( n35961 , n35960 , n22217 );
nor ( n35962 , n22219 , n380919 );
or ( n35963 , n35961 , n35962 );
nand ( n35964 , n35963 , n20623 );
or ( n35965 , n22224 , n380925 );
and ( n35966 , n35964 , n35965 );
nor ( n35967 , n35966 , n22236 );
not ( n35968 , n35967 );
and ( n35969 , n35968 , RI15b3ffd8_48);
or ( n35970 , n381917 , n35959 );
not ( n35971 , n35965 );
nor ( n35972 , n35962 , n35971 );
or ( n35973 , n35961 , n35972 );
not ( n35974 , n35973 );
and ( n35975 , n35974 , n381923 );
and ( n35976 , n381926 , n35971 );
nor ( n35977 , n35975 , n35976 );
nand ( n35978 , n35970 , n35977 );
nor ( n35979 , n35969 , n35978 );
nand ( n35980 , n35958 , n35979 );
buf ( n35981 , n35980 );
buf ( n35982 , n35651 );
and ( n35983 , n381492 , n35783 );
not ( n35984 , n35983 );
or ( n35985 , n386588 , n35984 );
nand ( n35986 , n381526 , n35788 );
not ( n35987 , n35986 );
and ( n35988 , n386600 , n35987 );
and ( n35989 , n35986 , n35984 , n381531 );
nor ( n35990 , n35989 , n19630 );
nor ( n35991 , n381534 , n35797 );
or ( n35992 , n35990 , n35991 );
nand ( n35993 , n35992 , n19595 );
or ( n35994 , n381539 , n380728 );
nand ( n35995 , n35993 , n35994 );
and ( n35996 , n35995 , n380775 );
or ( n35997 , n35996 , n18625 );
not ( n35998 , n35991 );
not ( n35999 , n35994 );
not ( n36000 , n35999 );
and ( n36001 , n35998 , n36000 );
nor ( n36002 , n36001 , n35990 );
not ( n36003 , n36002 );
or ( n36004 , n34706 , n36003 );
or ( n36005 , n35994 , n386627 );
nand ( n36006 , n35997 , n36004 , n36005 );
nor ( n36007 , n35988 , n36006 );
nand ( n36008 , n35985 , n36007 );
buf ( n36009 , n36008 );
buf ( n36010 , n21800 );
not ( n36011 , RI15b535b0_709);
not ( n36012 , n383170 );
or ( n36013 , n36011 , n36012 );
and ( n36014 , n33453 , RI15b54b40_755);
and ( n36015 , n383147 , RI15b52e30_693);
nor ( n36016 , n36014 , n36015 );
nand ( n36017 , n36013 , n36016 );
buf ( n36018 , n36017 );
buf ( n36019 , n32981 );
buf ( n36020 , n382049 );
and ( n36021 , n32747 , RI15b42b70_141);
not ( n36022 , n32749 );
buf ( n36023 , n36022 );
and ( n36024 , n32753 , RI15b418b0_101);
and ( n36025 , n32762 , RI15b414f0_93);
nor ( n36026 , n36024 , n36025 );
and ( n36027 , n32755 , RI15b41c70_109);
and ( n36028 , n32759 , RI15b41130_85);
nor ( n36029 , n36027 , n36028 );
and ( n36030 , n32771 , RI15b43a70_173);
and ( n36031 , n32773 , RI15b42f30_149);
nor ( n36032 , n36030 , n36031 );
and ( n36033 , n32766 , RI15b436b0_165);
and ( n36034 , n32768 , RI15b432f0_157);
nor ( n36035 , n36033 , n36034 );
nand ( n36036 , n36026 , n36029 , n36032 , n36035 );
and ( n36037 , n36023 , n36036 );
and ( n36038 , n32781 , RI15b405f0_61);
nor ( n36039 , n36021 , n36037 , n36038 );
and ( n36040 , n32785 , RI15b427b0_133);
and ( n36041 , n32787 , RI15b423f0_125);
nor ( n36042 , n36040 , n36041 );
and ( n36043 , n32792 , RI15b40230_53);
and ( n36044 , n32794 , RI15b42030_117);
nor ( n36045 , n36043 , n36044 );
and ( n36046 , n32797 , RI15b409b0_69);
and ( n36047 , n32800 , RI15b40d70_77);
nor ( n36048 , n36046 , n36047 );
nand ( n36049 , n36039 , n36042 , n36045 , n36048 );
not ( n36050 , n36049 );
buf ( n36051 , n32805 );
or ( n36052 , n36050 , n36051 );
and ( n36053 , n381055 , RI15b49a88_378);
not ( n36054 , RI15b49a88_378);
nand ( n36055 , n32823 , RI15b49920_375);
not ( n36056 , RI15b49998_376);
nor ( n36057 , n36055 , n36056 );
and ( n36058 , n36057 , RI15b49a10_377);
not ( n36059 , n36058 );
not ( n36060 , n36059 );
or ( n36061 , n36054 , n36060 );
or ( n36062 , n36059 , RI15b49a88_378);
nand ( n36063 , n36061 , n36062 );
buf ( n36064 , n381075 );
and ( n36065 , n36063 , n36064 );
nor ( n36066 , n36053 , n36065 );
nand ( n36067 , n36052 , n36066 );
buf ( n36068 , n36067 );
not ( n36069 , RI15b53e20_727);
not ( n36070 , n32244 );
or ( n36071 , n36069 , n36070 );
and ( n36072 , n32247 , RI15b65418_1320);
and ( n36073 , n32249 , RI15b60288_1146);
nor ( n36074 , n36072 , n36073 );
nand ( n36075 , n36071 , n36074 );
buf ( n36076 , n36075 );
buf ( n36077 , n381081 );
buf ( n36078 , n20663 );
buf ( n36079 , n20665 );
buf ( n36080 , n20665 );
buf ( n36081 , n22788 );
or ( n36082 , n35929 , n22227 );
or ( n36083 , n22102 , n36082 );
and ( n36084 , n22132 , n32163 );
and ( n36085 , n22203 , n36084 );
not ( n36086 , n36084 );
and ( n36087 , n36082 , n36086 , n19912 );
nor ( n36088 , n36087 , n22217 );
nor ( n36089 , n35939 , n35905 );
or ( n36090 , n36088 , n36089 );
nand ( n36091 , n36090 , n20623 );
or ( n36092 , n35943 , n22133 );
and ( n36093 , n36091 , n36092 );
nor ( n36094 , n36093 , n22236 );
or ( n36095 , n36094 , n385517 );
not ( n36096 , n36092 );
nor ( n36097 , n36089 , n36096 );
or ( n36098 , n36088 , n36097 );
or ( n36099 , n22293 , n36098 );
or ( n36100 , n36092 , n22299 );
nand ( n36101 , n36095 , n36099 , n36100 );
nor ( n36102 , n36085 , n36101 );
nand ( n36103 , n36083 , n36102 );
buf ( n36104 , n36103 );
buf ( n36105 , n22714 );
or ( n36106 , n22298 , RI15b3fc90_41);
not ( n36107 , n385999 );
not ( n36108 , n35368 );
or ( n36109 , n36107 , n36108 );
nand ( n36110 , n36109 , n20626 , n20008 );
nand ( n36111 , n36110 , n385209 );
or ( n36112 , n22235 , n36111 );
nand ( n36113 , n36112 , RI15b3fc90_41);
nand ( n36114 , n20626 , RI15b3fc18_40);
nand ( n36115 , n36106 , n36113 , n36114 );
buf ( n36116 , n36115 );
buf ( n36117 , n380906 );
buf ( n36118 , n379844 );
nand ( n36119 , n35851 , n20637 );
nand ( n36120 , n22147 , n22209 );
or ( n36121 , n22143 , n36120 );
or ( n36122 , n36119 , n36121 );
and ( n36123 , n32168 , n22134 );
not ( n36124 , n36123 );
and ( n36125 , n36121 , n36124 , n19912 );
nor ( n36126 , n36125 , n22217 );
nor ( n36127 , n32175 , n35877 );
or ( n36128 , n36126 , n36127 );
nand ( n36129 , n36128 , n20623 );
or ( n36130 , n22105 , n380923 );
and ( n36131 , n36129 , n36130 );
nor ( n36132 , n36131 , n22236 );
not ( n36133 , n36132 );
and ( n36134 , n36133 , RI15b43728_166);
or ( n36135 , n35856 , n36130 );
not ( n36136 , n36130 );
or ( n36137 , n36127 , n36136 );
not ( n36138 , n36126 );
nand ( n36139 , n36137 , n36138 );
or ( n36140 , n35582 , n36139 );
or ( n36141 , n36124 , n35858 );
nand ( n36142 , n36135 , n36140 , n36141 );
nor ( n36143 , n36134 , n36142 );
nand ( n36144 , n36122 , n36143 );
buf ( n36145 , n36144 );
buf ( n36146 , n382537 );
buf ( n36147 , n383498 );
not ( n36148 , n385130 );
nor ( n36149 , n36148 , n21699 );
not ( n36150 , n36149 );
not ( n36151 , n21699 );
nor ( n36152 , n385129 , n36151 );
not ( n36153 , n36152 );
nand ( n36154 , n36150 , n36153 );
nand ( n36155 , n36154 , n21748 );
not ( n36156 , n21301 );
not ( n36157 , n21294 );
not ( n36158 , n36157 );
or ( n36159 , n36156 , n36158 );
or ( n36160 , n36157 , n21301 );
nand ( n36161 , n36159 , n36160 );
buf ( n36162 , n21357 );
and ( n36163 , n36161 , n36162 );
not ( n36164 , n21511 );
not ( n36165 , n36164 );
not ( n36166 , n21515 );
and ( n36167 , n36165 , n36166 );
and ( n36168 , n36164 , n21515 );
nor ( n36169 , n36167 , n36168 );
or ( n36170 , n36169 , n385148 );
or ( n36171 , n21750 , n21986 );
nand ( n36172 , n36170 , n36171 );
nor ( n36173 , n36163 , n36172 );
nand ( n36174 , n36155 , n36173 );
not ( n36175 , n36174 );
and ( n36176 , n385164 , RI15b506d0_609);
or ( n36177 , n21301 , n385170 );
not ( n36178 , n385174 );
or ( n36179 , n36178 , n21699 );
or ( n36180 , n21515 , n385178 );
nand ( n36181 , n36177 , n36179 , n36180 );
nor ( n36182 , n36176 , n36181 );
nand ( n36183 , n36175 , n36182 );
buf ( n36184 , n36183 );
buf ( n36185 , n384203 );
or ( n36186 , n385188 , RI15b608a0_1159);
not ( n36187 , n379794 );
and ( n36188 , n36187 , RI15b5e7d0_1089);
nor ( n36189 , n36188 , n33104 );
nand ( n36190 , n36186 , n36189 );
buf ( n36191 , n36190 );
buf ( n36192 , n20665 );
and ( n36193 , n22646 , RI15b45780_235);
and ( n36194 , n22648 , RI15b51be8_654);
nor ( n36195 , n36193 , n36194 );
not ( n36196 , n36195 );
buf ( n36197 , n36196 );
buf ( n36198 , n381004 );
buf ( n36199 , n382065 );
or ( n36200 , n35929 , n22150 );
or ( n36201 , n22315 , n36200 );
and ( n36202 , n22132 , n32169 );
and ( n36203 , n22326 , n36202 );
not ( n36204 , n36202 );
and ( n36205 , n36200 , n36204 , n19912 );
nor ( n36206 , n36205 , n22217 );
nor ( n36207 , n35939 , n22133 );
or ( n36208 , n36206 , n36207 );
nand ( n36209 , n36208 , n20623 );
or ( n36210 , n35943 , n22227 );
and ( n36211 , n36209 , n36210 );
nor ( n36212 , n36211 , n22236 );
not ( n36213 , RI15b416d0_97);
or ( n36214 , n36212 , n36213 );
not ( n36215 , n36210 );
nor ( n36216 , n36207 , n36215 );
or ( n36217 , n36206 , n36216 );
or ( n36218 , n22334 , n36217 );
or ( n36219 , n36210 , n22336 );
nand ( n36220 , n36214 , n36218 , n36219 );
nor ( n36221 , n36203 , n36220 );
nand ( n36222 , n36201 , n36221 );
buf ( n36223 , n36222 );
buf ( n36224 , n383174 );
buf ( n36225 , n30992 );
buf ( n36226 , n22714 );
buf ( n36227 , RI15b5e1b8_1076);
not ( n36228 , RI15b61c50_1201);
or ( n36229 , n384021 , n36228 );
or ( n36230 , n18955 , n386747 );
or ( n36231 , RI15b61c50_1201 , n384024 );
nand ( n36232 , n36229 , n36230 , n36231 );
buf ( n36233 , n36232 );
buf ( n36234 , n380942 );
buf ( n36235 , n19653 );
not ( n36236 , n383777 );
buf ( n36237 , n383854 );
nand ( n36238 , n36236 , n36237 );
nand ( n36239 , n31162 , n383866 );
or ( n36240 , n36238 , n36239 );
not ( n36241 , RI15b4d250_497);
nand ( n36242 , n383841 , n383843 );
and ( n36243 , n36239 , n36242 , n385009 );
nor ( n36244 , n36243 , n21764 );
nor ( n36245 , n31168 , n383888 );
or ( n36246 , n36244 , n36245 );
nand ( n36247 , n36246 , n18154 );
or ( n36248 , n31172 , n383894 );
and ( n36249 , n36247 , n36248 );
nor ( n36250 , n36249 , n383902 );
or ( n36251 , n36241 , n36250 );
not ( n36252 , n36248 );
nor ( n36253 , n36245 , n36252 );
or ( n36254 , n36244 , n36253 );
not ( n36255 , n36254 );
not ( n36256 , n32709 );
buf ( n36257 , n36256 );
and ( n36258 , n36255 , n36257 );
not ( n36259 , n36242 );
and ( n36260 , n383803 , n36259 );
and ( n36261 , n17991 , n383915 );
and ( n36262 , n36261 , n36252 );
nor ( n36263 , n36258 , n36260 , n36262 );
nand ( n36264 , n36240 , n36251 , n36263 );
buf ( n36265 , n36264 );
not ( n36266 , n381406 );
or ( n36267 , n36266 , n32452 );
not ( n36268 , n32401 );
buf ( n36269 , n36268 );
nand ( n36270 , n36269 , RI15b549d8_752);
and ( n36271 , n32454 , n36270 );
nand ( n36272 , n381486 , RI15b52cc8_690);
nand ( n36273 , n36267 , n36271 , n36272 );
buf ( n36274 , n36273 );
nand ( n36275 , n381492 , n380737 );
not ( n36276 , n36275 );
not ( n36277 , n36276 );
not ( n36278 , n33400 );
or ( n36279 , n36277 , n36278 );
not ( n36280 , n32068 );
nand ( n36281 , n36280 , n382980 );
not ( n36282 , n36281 );
and ( n36283 , n33415 , n36282 );
and ( n36284 , n36281 , n36275 , n32072 );
nor ( n36285 , n36284 , n19630 );
nor ( n36286 , n381534 , n35154 );
or ( n36287 , n36285 , n36286 );
nand ( n36288 , n36287 , n19595 );
or ( n36289 , n380207 , n381538 );
nand ( n36290 , n36288 , n36289 );
and ( n36291 , n36290 , n380775 );
or ( n36292 , n36291 , n18457 );
not ( n36293 , n33432 );
not ( n36294 , n36289 );
nor ( n36295 , n36286 , n36294 );
or ( n36296 , n36285 , n36295 );
or ( n36297 , n36293 , n36296 );
or ( n36298 , n36289 , n33443 );
nand ( n36299 , n36292 , n36297 , n36298 );
nor ( n36300 , n36283 , n36299 );
nand ( n36301 , n36279 , n36300 );
buf ( n36302 , n36301 );
buf ( n36303 , n380903 );
buf ( n36304 , n386762 );
buf ( n36305 , RI15b5df60_1071);
or ( n36306 , n22142 , n36120 );
or ( n36307 , n381907 , n36306 );
not ( n36308 , n381917 );
not ( n36309 , n22135 );
and ( n36310 , n36308 , n36309 );
and ( n36311 , n36306 , n22135 , n19912 );
nor ( n36312 , n36311 , n22217 );
or ( n36313 , n36312 , n22119 );
nand ( n36314 , n36313 , n20623 );
not ( n36315 , n22223 );
or ( n36316 , n22105 , n36315 );
and ( n36317 , n36314 , n36316 );
nor ( n36318 , n36317 , n22236 );
not ( n36319 , RI15b41a18_104);
or ( n36320 , n36318 , n36319 );
not ( n36321 , n381923 );
not ( n36322 , n36316 );
or ( n36323 , n22119 , n36322 );
not ( n36324 , n36312 );
nand ( n36325 , n36323 , n36324 );
or ( n36326 , n36321 , n36325 );
not ( n36327 , n381926 );
or ( n36328 , n36316 , n36327 );
nand ( n36329 , n36320 , n36326 , n36328 );
nor ( n36330 , n36310 , n36329 );
nand ( n36331 , n36307 , n36330 );
buf ( n36332 , n36331 );
buf ( n36333 , n33382 );
buf ( n36334 , n31979 );
buf ( n36335 , n383174 );
buf ( n36336 , n381004 );
buf ( n36337 , n382065 );
buf ( n36338 , n384203 );
not ( n36339 , RI15b525c0_675);
not ( n36340 , n32397 );
or ( n36341 , n36339 , n36340 );
not ( n36342 , n381422 );
or ( n36343 , n383110 , n36342 );
nand ( n36344 , n36343 , n381450 );
and ( n36345 , n36344 , n383102 );
not ( n36346 , n381461 );
not ( n36347 , n383110 );
nor ( n36348 , n36347 , n383102 );
not ( n36349 , n36348 );
or ( n36350 , n36346 , n36349 );
nand ( n36351 , n381401 , n31177 );
nand ( n36352 , n36350 , n36351 );
nor ( n36353 , n36345 , n36352 );
nand ( n36354 , n36341 , n36353 );
buf ( n36355 , n36354 );
not ( n36356 , n31793 );
not ( n36357 , n384518 );
and ( n36358 , n36356 , n36357 );
or ( n36359 , n31771 , n384413 );
or ( n36360 , n384295 , n32378 );
or ( n36361 , n35265 , n31779 );
nand ( n36362 , n36359 , n36360 , n36361 );
nor ( n36363 , n36358 , n36362 );
nand ( n36364 , n35278 , n36363 );
buf ( n36365 , n36364 );
buf ( n36366 , n380903 );
buf ( n36367 , RI15b47418_296);
not ( n36368 , n33165 );
not ( n36369 , n32129 );
or ( n36370 , n36368 , n36369 );
and ( n36371 , n33080 , RI15b41d60_111);
or ( n36372 , n32141 , n380915 );
or ( n36373 , n32148 , n380933 );
or ( n36374 , n380926 , n32150 );
nand ( n36375 , n36372 , n36373 , n36374 );
nor ( n36376 , n36371 , n36375 );
nand ( n36377 , n36370 , n36376 );
buf ( n36378 , n36377 );
buf ( n36379 , n19653 );
buf ( n36380 , n17499 );
buf ( n36381 , n384996 );
buf ( n36382 , n22406 );
or ( n36383 , n380001 , n18081 );
buf ( n36384 , n380009 );
and ( n36385 , n36384 , RI15b4c440_467);
and ( n36386 , n379951 , n18081 );
not ( n36387 , n379951 );
and ( n36388 , n36387 , RI15b558d8_784);
nor ( n36389 , n36386 , n36388 );
and ( n36390 , n379949 , n36389 );
nor ( n36391 , n36385 , n36390 );
nand ( n36392 , n36383 , n36391 );
buf ( n36393 , n36392 );
nand ( n36394 , n381568 , n380737 );
not ( n36395 , n36394 );
not ( n36396 , n36395 );
not ( n36397 , n381507 );
or ( n36398 , n36396 , n36397 );
not ( n36399 , n380743 );
nand ( n36400 , n36399 , n381493 );
not ( n36401 , n36400 );
and ( n36402 , n381524 , n36401 );
and ( n36403 , n36400 , n36394 , n382985 );
nor ( n36404 , n36403 , n19630 );
nor ( n36405 , n380755 , n35154 );
or ( n36406 , n36404 , n36405 );
nand ( n36407 , n36406 , n19595 );
or ( n36408 , n380764 , n380756 );
nand ( n36409 , n36407 , n36408 );
and ( n36410 , n36409 , n380775 );
or ( n36411 , n36410 , n18417 );
not ( n36412 , n381549 );
buf ( n36413 , n36412 );
not ( n36414 , n36408 );
nor ( n36415 , n36405 , n36414 );
or ( n36416 , n36404 , n36415 );
or ( n36417 , n36413 , n36416 );
or ( n36418 , n36408 , n381560 );
nand ( n36419 , n36411 , n36417 , n36418 );
nor ( n36420 , n36402 , n36419 );
nand ( n36421 , n36398 , n36420 );
buf ( n36422 , n36421 );
buf ( n36423 , n386760 );
buf ( n36424 , n383498 );
not ( n36425 , n381726 );
nand ( n36426 , n36425 , n381753 );
and ( n36427 , n381722 , RI15b50b80_619);
nand ( n36428 , n381714 , RI15b50b08_618);
nor ( n36429 , n36428 , RI15b50b80_619);
not ( n36430 , n36429 );
not ( n36431 , n381718 );
or ( n36432 , n36430 , n36431 );
and ( n36433 , n36428 , RI15b50b80_619);
not ( n36434 , n36433 );
nand ( n36435 , n36432 , n36434 );
nor ( n36436 , n36427 , n36435 );
and ( n36437 , n36426 , n36436 );
not ( n36438 , n36426 );
not ( n36439 , n36436 );
and ( n36440 , n36438 , n36439 );
nor ( n36441 , n36437 , n36440 );
not ( n36442 , n22687 );
buf ( n36443 , n36442 );
and ( n36444 , n36441 , n36443 );
nor ( n36445 , n21750 , n22839 );
nor ( n36446 , n36444 , n36445 );
nor ( n36447 , n381779 , n381784 );
not ( n36448 , n36447 );
and ( n36449 , n20692 , RI15b50b80_619);
and ( n36450 , n20691 , n36429 );
nor ( n36451 , n36449 , n36450 , n36433 );
and ( n36452 , n36448 , n36451 );
not ( n36453 , n36448 );
not ( n36454 , n36451 );
and ( n36455 , n36453 , n36454 );
nor ( n36456 , n36452 , n36455 );
buf ( n36457 , n36162 );
nand ( n36458 , n36456 , n36457 );
buf ( n36459 , n381806 );
not ( n36460 , n36459 );
and ( n36461 , n36460 , n36429 );
and ( n36462 , n36459 , RI15b50b80_619);
nor ( n36463 , n36461 , n36462 , n36433 );
nor ( n36464 , n381821 , n36463 );
not ( n36465 , n36464 );
and ( n36466 , n381820 , n36463 );
not ( n36467 , n36466 );
nand ( n36468 , n36465 , n36467 );
nand ( n36469 , n36468 , n21748 );
and ( n36470 , n36446 , n36458 , n36469 );
and ( n36471 , n385164 , RI15b50b80_619);
buf ( n36472 , n385172 );
buf ( n36473 , n36472 );
not ( n36474 , n36473 );
or ( n36475 , n36474 , n36463 );
or ( n36476 , n36451 , n385170 );
or ( n36477 , n36436 , n385178 );
nand ( n36478 , n36475 , n36476 , n36477 );
nor ( n36479 , n36471 , n36478 );
nand ( n36480 , n36470 , n36479 );
buf ( n36481 , n36480 );
buf ( n36482 , n386760 );
buf ( n36483 , n380903 );
buf ( n36484 , n34269 );
not ( n36485 , n34283 );
buf ( n36486 , n34059 );
nor ( n36487 , n36485 , n36486 );
nand ( n36488 , n36484 , n36487 );
not ( n36489 , n34231 );
nor ( n36490 , n36488 , n36489 );
buf ( n36491 , n36490 );
nand ( n36492 , n36491 , n379785 );
not ( n36493 , n36492 );
not ( n36494 , n34295 );
not ( n36495 , n36494 );
not ( n36496 , n36495 );
not ( n36497 , n36496 );
or ( n36498 , n36493 , n36497 );
not ( n36499 , n33995 );
nand ( n36500 , n36498 , n36499 );
not ( n36501 , n34249 );
not ( n36502 , n36501 );
nor ( n36503 , n36491 , n36499 );
nand ( n36504 , n36502 , n36503 );
buf ( n36505 , n34558 );
buf ( n36506 , n34567 );
and ( n36507 , n36505 , n36506 );
not ( n36508 , n36505 );
not ( n36509 , n36506 );
and ( n36510 , n36508 , n36509 );
nor ( n36511 , n36507 , n36510 );
buf ( n36512 , n34644 );
buf ( n36513 , n36512 );
and ( n36514 , n36511 , n36513 );
not ( n36515 , RI15b5e320_1079);
not ( n36516 , n34651 );
or ( n36517 , n36515 , n36516 );
not ( n36518 , n379783 );
or ( n36519 , n36518 , n379711 );
nand ( n36520 , n36517 , n36519 );
nor ( n36521 , n36514 , n36520 );
nand ( n36522 , n36500 , n36504 , n36521 );
buf ( n36523 , n36522 );
or ( n36524 , n31149 , n35472 );
and ( n36525 , n31161 , n35479 );
not ( n36526 , RI15b4de80_523);
or ( n36527 , n35488 , n36526 );
or ( n36528 , n31179 , n35497 );
or ( n36529 , n35486 , n31184 );
nand ( n36530 , n36527 , n36528 , n36529 );
nor ( n36531 , n36525 , n36530 );
nand ( n36532 , n36524 , n36531 );
buf ( n36533 , n36532 );
or ( n36534 , n31053 , n36412 );
nand ( n36535 , n384907 , n384870 );
not ( n36536 , n31091 );
and ( n36537 , n36536 , RI15b61020_1175);
buf ( n36538 , n35507 );
and ( n36539 , n36538 , n382589 );
not ( n36540 , n31082 );
not ( n36541 , n36540 );
not ( n36542 , RI15b61020_1175);
not ( n36543 , n31066 );
not ( n36544 , n36543 );
or ( n36545 , n36542 , n36544 );
or ( n36546 , n36543 , RI15b61020_1175);
nand ( n36547 , n36545 , n36546 );
and ( n36548 , n36541 , n36547 );
nor ( n36549 , n36537 , n36539 , n36548 );
nand ( n36550 , n36534 , n36535 , n36549 );
buf ( n36551 , n36550 );
buf ( n36552 , n379802 );
buf ( n36553 , n387159 );
buf ( n36554 , n382067 );
buf ( n36555 , n34263 );
and ( n36556 , n34282 , n36555 );
buf ( n36557 , n34256 );
nand ( n36558 , n36556 , n36557 );
buf ( n36559 , n34142 );
nor ( n36560 , n36558 , n36559 );
buf ( n36561 , n34268 );
buf ( n36562 , n34014 );
nor ( n36563 , n36561 , n36562 );
nand ( n36564 , n36560 , n36563 );
not ( n36565 , n34058 );
nor ( n36566 , n36564 , n36565 );
buf ( n36567 , n34124 );
nand ( n36568 , n36566 , n36567 );
buf ( n36569 , n34209 );
nor ( n36570 , n36568 , n36569 );
nand ( n36571 , n36570 , n379785 );
not ( n36572 , n36571 );
not ( n36573 , n36494 );
not ( n36574 , n36573 );
not ( n36575 , n36574 );
or ( n36576 , n36572 , n36575 );
buf ( n36577 , n34044 );
not ( n36578 , n36577 );
nand ( n36579 , n36576 , n36578 );
not ( n36580 , n36501 );
not ( n36581 , n36570 );
nand ( n36582 , n36580 , n36581 , n36577 );
not ( n36583 , n34528 );
not ( n36584 , n34511 );
not ( n36585 , n36584 );
or ( n36586 , n36583 , n36585 );
or ( n36587 , n36584 , n34528 );
nand ( n36588 , n36586 , n36587 );
and ( n36589 , n36588 , n34646 );
and ( n36590 , n379783 , RI15b643b0_1285);
and ( n36591 , n34651 , RI15b5e1b8_1076);
nor ( n36592 , n36590 , n36591 );
not ( n36593 , n36592 );
nor ( n36594 , n36589 , n36593 );
nand ( n36595 , n36579 , n36582 , n36594 );
buf ( n36596 , n36595 );
buf ( n36597 , n381006 );
buf ( n36598 , n22408 );
and ( n36599 , n381722 , RI15b50bf8_620);
not ( n36600 , n36428 );
and ( n36601 , n36600 , RI15b50b80_619);
not ( n36602 , n36601 );
nor ( n36603 , n36602 , RI15b50bf8_620);
not ( n36604 , n36603 );
not ( n36605 , n381718 );
or ( n36606 , n36604 , n36605 );
not ( n36607 , RI15b50bf8_620);
nor ( n36608 , n36601 , n36607 );
not ( n36609 , n36608 );
nand ( n36610 , n36606 , n36609 );
nor ( n36611 , n36599 , n36610 );
not ( n36612 , n36611 );
nor ( n36613 , n36426 , n36436 );
nand ( n36614 , n36612 , n36613 );
buf ( n36615 , n381722 );
and ( n36616 , n36615 , RI15b50c70_621);
nand ( n36617 , n36601 , RI15b50bf8_620);
nor ( n36618 , n36617 , RI15b50c70_621);
not ( n36619 , n36618 );
not ( n36620 , n381747 );
or ( n36621 , n36619 , n36620 );
nand ( n36622 , n36617 , RI15b50c70_621);
nand ( n36623 , n36621 , n36622 );
nor ( n36624 , n36616 , n36623 );
nor ( n36625 , n36614 , n36624 );
not ( n36626 , n36625 );
buf ( n36627 , n381720 );
buf ( n36628 , n36627 );
not ( n36629 , n36628 );
and ( n36630 , n36629 , RI15b50ce8_622);
not ( n36631 , n36617 );
and ( n36632 , n36631 , RI15b50c70_621);
not ( n36633 , n36632 );
nor ( n36634 , n36633 , RI15b50ce8_622);
and ( n36635 , n36627 , n36634 );
not ( n36636 , RI15b50ce8_622);
nor ( n36637 , n36632 , n36636 );
nor ( n36638 , n36635 , n36637 );
not ( n36639 , n36638 );
nor ( n36640 , n36630 , n36639 );
and ( n36641 , n36626 , n36640 );
not ( n36642 , n36626 );
not ( n36643 , n36640 );
and ( n36644 , n36642 , n36643 );
nor ( n36645 , n36641 , n36644 );
and ( n36646 , n36645 , n21564 );
nor ( n36647 , n21750 , n22623 );
nor ( n36648 , n36646 , n36647 );
and ( n36649 , n36447 , n36454 );
and ( n36650 , n20692 , RI15b50bf8_620);
and ( n36651 , n20691 , n36603 );
nor ( n36652 , n36650 , n36651 , n36608 );
not ( n36653 , n36652 );
nand ( n36654 , n36649 , n36653 );
and ( n36655 , n20692 , RI15b50c70_621);
and ( n36656 , n20691 , n36618 );
not ( n36657 , n36622 );
nor ( n36658 , n36655 , n36656 , n36657 );
nor ( n36659 , n36654 , n36658 );
not ( n36660 , n36659 );
and ( n36661 , n36634 , n20691 );
and ( n36662 , n20692 , RI15b50ce8_622);
nor ( n36663 , n36661 , n36662 , n36637 );
and ( n36664 , n36660 , n36663 );
not ( n36665 , n36660 );
not ( n36666 , n36663 );
and ( n36667 , n36665 , n36666 );
nor ( n36668 , n36664 , n36667 );
nand ( n36669 , n36668 , n21361 );
not ( n36670 , n36459 );
and ( n36671 , n36670 , n36603 );
and ( n36672 , n36459 , RI15b50bf8_620);
nor ( n36673 , n36671 , n36672 , n36608 );
nand ( n36674 , n36466 , n36673 );
and ( n36675 , n36670 , n36618 );
and ( n36676 , n36459 , RI15b50c70_621);
nor ( n36677 , n36675 , n36676 , n36657 );
not ( n36678 , n36677 );
nor ( n36679 , n36674 , n36678 );
buf ( n36680 , n36459 );
not ( n36681 , n36680 );
and ( n36682 , n36681 , n36634 );
and ( n36683 , n36680 , RI15b50ce8_622);
nor ( n36684 , n36682 , n36683 , n36637 );
nor ( n36685 , n36679 , n36684 );
not ( n36686 , n36685 );
nand ( n36687 , n36679 , n36684 );
nand ( n36688 , n36686 , n36687 );
buf ( n36689 , n33644 );
nand ( n36690 , n36688 , n36689 );
and ( n36691 , n36648 , n36669 , n36690 );
and ( n36692 , n385164 , RI15b50ce8_622);
not ( n36693 , n385174 );
buf ( n36694 , n36693 );
or ( n36695 , n36694 , n36684 );
or ( n36696 , n36663 , n385170 );
or ( n36697 , n36640 , n385178 );
nand ( n36698 , n36695 , n36696 , n36697 );
nor ( n36699 , n36692 , n36698 );
nand ( n36700 , n36691 , n36699 );
buf ( n36701 , n36700 );
buf ( n36702 , n32676 );
buf ( n36703 , n383613 );
buf ( n36704 , RI15b3ea48_2);
buf ( n36705 , n36704 );
buf ( n36706 , n382067 );
nand ( n36707 , n20606 , n386552 );
nand ( n36708 , n20586 , n20601 , n36707 );
and ( n36709 , RI15b449e8_206 , n36708 );
not ( n36710 , RI15b449e8_206);
nand ( n36711 , n20606 , n381061 );
nand ( n36712 , n20609 , n36711 );
and ( n36713 , n36710 , n36712 );
nor ( n36714 , n36709 , n36713 );
buf ( n36715 , n32164 );
nand ( n36716 , n36714 , n36715 );
and ( n36717 , n36716 , n20417 );
not ( n36718 , n36717 );
not ( n36719 , RI15b3fc90_41);
not ( n36720 , n36714 );
or ( n36721 , n36719 , n36720 );
nand ( n36722 , n36721 , n20423 );
not ( n36723 , n385261 );
not ( n36724 , n36723 );
nand ( n36725 , n36724 , n36712 );
not ( n36726 , n386527 );
nand ( n36727 , n20580 , n379828 );
and ( n36728 , n36726 , n36727 , n36707 , n386255 );
and ( n36729 , RI15b44a60_207 , n36728 );
not ( n36730 , RI15b44a60_207);
nand ( n36731 , n20580 , n379818 );
and ( n36732 , n386545 , n36731 );
and ( n36733 , n36730 , n36732 );
or ( n36734 , n36729 , n36733 );
and ( n36735 , n36725 , n36734 );
nand ( n36736 , n36722 , n36735 );
not ( n36737 , n36736 );
or ( n36738 , n36718 , n36737 );
buf ( n36739 , n385272 );
buf ( n36740 , n36739 );
and ( n36741 , n20608 , n36740 );
not ( n36742 , RI15b44ad8_208);
or ( n36743 , n36728 , n36742 );
or ( n36744 , n32741 , n36732 );
or ( n36745 , n36739 , n36711 );
nand ( n36746 , n36743 , n36744 , n36745 );
nor ( n36747 , n36741 , n36746 );
nand ( n36748 , n36738 , n36747 );
not ( n36749 , n36716 );
not ( n36750 , n36736 );
or ( n36751 , n36749 , n36750 );
nand ( n36752 , n36751 , RI15b3fd80_43);
nand ( n36753 , n36748 , n36752 );
or ( n36754 , n36753 , n36315 );
not ( n36755 , n20492 );
not ( n36756 , n385201 );
or ( n36757 , n36755 , n36756 );
nand ( n36758 , n385204 , n20516 );
nand ( n36759 , n36757 , n36758 );
nand ( n36760 , n36759 , RI15b44c40_211);
not ( n36761 , n383369 );
or ( n36762 , n20586 , n36761 );
not ( n36763 , n386522 );
nand ( n36764 , n36760 , n36762 , n36763 , n36707 );
or ( n36765 , n381024 , n386010 );
nand ( n36766 , n36759 , n383370 , RI15b3fc18_40);
not ( n36767 , n386257 );
nand ( n36768 , n36765 , n36766 , n36767 );
nor ( n36769 , n36764 , n36768 );
nand ( n36770 , n36754 , n36769 );
nand ( n36771 , n36770 , n20501 );
and ( n36772 , n20634 , n20492 );
not ( n36773 , n36108 );
nand ( n36774 , n35335 , n36773 , RI15b44a60_207);
not ( n36775 , n36774 );
nor ( n36776 , n36772 , n36775 );
nand ( n36777 , n36771 , n36776 );
not ( n36778 , n36753 );
nand ( n36779 , n36778 , n20461 );
and ( n36780 , n36747 , n36315 );
and ( n36781 , n36779 , n36780 );
buf ( n36782 , n385278 );
or ( n36783 , n20609 , n36782 );
not ( n36784 , RI15b44b50_209);
or ( n36785 , n36784 , n36728 );
or ( n36786 , n36732 , n32735 );
not ( n36787 , n36711 );
or ( n36788 , n35372 , RI15b44b50_209);
not ( n36789 , n35388 );
nand ( n36790 , n36788 , n36789 );
and ( n36791 , n36787 , n36790 );
and ( n36792 , n20606 , n385334 );
nor ( n36793 , n36791 , n36792 );
nand ( n36794 , n36786 , n36793 );
not ( n36795 , n36794 );
nand ( n36796 , n36783 , n36785 , n36795 );
nand ( n36797 , n36796 , n20501 );
nor ( n36798 , n36781 , n36797 );
nor ( n36799 , n36777 , n36798 );
not ( n36800 , n20584 );
or ( n36801 , n36800 , n20517 );
and ( n36802 , n36801 , n20501 );
and ( n36803 , n20631 , n20491 );
or ( n36804 , n20621 , n20491 );
nand ( n36805 , n36804 , n32619 , n36114 );
nor ( n36806 , n36803 , n36805 , n22233 );
not ( n36807 , n36111 );
nand ( n36808 , n36806 , n36807 , n386502 );
nor ( n36809 , n36802 , n385203 , n36808 );
nand ( n36810 , n36799 , n36809 );
buf ( n36811 , n36810 );
buf ( n36812 , n381872 );
or ( n36813 , n380908 , n22227 );
or ( n36814 , n36119 , n36813 );
nand ( n36815 , n22140 , n32164 );
and ( n36816 , n36813 , n36815 , n19912 );
nor ( n36817 , n36816 , n22217 );
not ( n36818 , n35904 );
nor ( n36819 , n380918 , n36818 );
or ( n36820 , n36817 , n36819 );
nand ( n36821 , n36820 , n20623 );
or ( n36822 , n380924 , n22133 );
and ( n36823 , n36821 , n36822 );
nor ( n36824 , n36823 , n22236 );
not ( n36825 , n36824 );
and ( n36826 , n36825 , RI15b420a8_118);
or ( n36827 , n35856 , n36822 );
not ( n36828 , n36822 );
nor ( n36829 , n36819 , n36828 );
or ( n36830 , n36817 , n36829 );
or ( n36831 , n35582 , n36830 );
or ( n36832 , n36815 , n35858 );
nand ( n36833 , n36827 , n36831 , n36832 );
nor ( n36834 , n36826 , n36833 );
nand ( n36835 , n36814 , n36834 );
buf ( n36836 , n36835 );
buf ( n36837 , n385195 );
buf ( n36838 , n379403 );
buf ( n36839 , n17499 );
buf ( n36840 , n19653 );
buf ( n36841 , n19655 );
not ( n36842 , RI15b4c080_459);
and ( n36843 , n32996 , n36842 );
nor ( n36844 , n36843 , n383900 );
not ( n36845 , n36844 );
nor ( n36846 , n36845 , n21774 );
or ( n36847 , n36846 , n18062 );
not ( n36848 , n21764 );
or ( n36849 , RI15b4c170_461 , n36848 );
nor ( n36850 , n21337 , n383866 );
or ( n36851 , n36850 , n383916 );
nand ( n36852 , n36847 , n36849 , n36851 );
buf ( n36853 , n36852 );
buf ( n36854 , RI15b3e9d0_1);
buf ( n36855 , n36854 );
buf ( n36856 , n381021 );
not ( n36857 , RI15b62d30_1237);
not ( n36858 , n19608 );
or ( n36859 , n36857 , n36858 );
buf ( n36860 , n386803 );
and ( n36861 , n19630 , n36860 );
buf ( n36862 , n386797 );
not ( n36863 , RI15b62d30_1237);
and ( n36864 , n36862 , n36863 );
not ( n36865 , n36862 );
and ( n36866 , n36865 , RI15b62d30_1237);
nor ( n36867 , n36864 , n36866 );
and ( n36868 , n19645 , n36867 );
buf ( n36869 , n18682 );
not ( n36870 , n18678 );
or ( n36871 , n18674 , n36870 );
nand ( n36872 , n36871 , n18552 );
and ( n36873 , n36869 , n36872 );
not ( n36874 , n36869 );
and ( n36875 , n36874 , n18679 );
nor ( n36876 , n36873 , n36875 );
not ( n36877 , n36876 );
not ( n36878 , n18451 );
and ( n36879 , n36877 , n36878 );
and ( n36880 , n36876 , n18451 );
nor ( n36881 , n36879 , n36880 );
or ( n36882 , n36881 , n19283 );
not ( n36883 , n382575 );
nand ( n36884 , n19444 , n382578 );
not ( n36885 , n36884 );
and ( n36886 , n36883 , n36885 );
and ( n36887 , n382575 , n36884 );
nor ( n36888 , n36886 , n36887 );
or ( n36889 , n22760 , n36888 );
and ( n36890 , n19308 , n18682 );
not ( n36891 , n19308 );
and ( n36892 , n36891 , n18509 );
nor ( n36893 , n36890 , n36892 );
not ( n36894 , n36893 );
not ( n36895 , n33024 );
or ( n36896 , n36894 , n36895 );
or ( n36897 , n33024 , n36893 );
nand ( n36898 , n36896 , n36897 );
and ( n36899 , n36898 , n19387 );
and ( n36900 , n19513 , RI15b63c30_1269);
nor ( n36901 , n36899 , n36900 );
nand ( n36902 , n36882 , n36889 , n36901 );
nor ( n36903 , n36861 , n36868 , n36902 );
nand ( n36904 , n36859 , n36903 );
buf ( n36905 , n36904 );
buf ( n36906 , n22009 );
buf ( n36907 , n384700 );
buf ( n36908 , n386563 );
and ( n36909 , n34931 , n20493 );
or ( n36910 , n20621 , n20492 );
or ( n36911 , n20630 , n20491 );
nand ( n36912 , n36910 , n36911 );
not ( n36913 , n19921 );
nor ( n36914 , n36909 , n36912 , n36913 );
nand ( n36915 , n36799 , n36914 );
buf ( n36916 , n36915 );
buf ( n36917 , n381707 );
buf ( n36918 , n380865 );
buf ( n36919 , n19651 );
buf ( n36920 , n385195 );
buf ( n36921 , n384218 );
and ( n36922 , n379822 , RI15b65b20_1335);
and ( n36923 , n379825 , RI15b48750_337);
nor ( n36924 , n36922 , n36923 );
nand ( n36925 , n379832 , RI15b46a40_275);
not ( n36926 , n22259 );
nand ( n36927 , n379835 , n36926 );
nand ( n36928 , n36924 , n36925 , n36927 );
buf ( n36929 , n36928 );
nor ( n36930 , n384108 , n384076 );
not ( n36931 , n36930 );
not ( n36932 , n386695 );
not ( n36933 , n384114 );
or ( n36934 , n36932 , n36933 );
nand ( n36935 , n36934 , n384076 );
nand ( n36936 , n36931 , n36935 );
not ( n36937 , n36936 );
or ( n36938 , n36937 , n385002 );
nor ( n36939 , n383851 , n382703 );
not ( n36940 , n36939 );
not ( n36941 , n384155 );
or ( n36942 , n36940 , n36941 );
nand ( n36943 , n384153 , n384710 );
and ( n36944 , n36943 , n384146 );
nor ( n36945 , n36944 , n384147 );
nand ( n36946 , n36942 , n36945 );
and ( n36947 , n36946 , n385006 );
not ( n36948 , RI15b4e3a8_534);
or ( n36949 , n385019 , n36948 );
buf ( n36950 , n35776 );
buf ( n36951 , n36950 );
not ( n36952 , n36951 );
or ( n36953 , n36952 , n385023 );
not ( n36954 , n18107 );
or ( n36955 , n36954 , n383916 );
or ( n36956 , n385017 , n36955 );
nand ( n36957 , n36949 , n36953 , n36956 );
nor ( n36958 , n36947 , n36957 );
nand ( n36959 , n36938 , n36958 );
buf ( n36960 , n36959 );
buf ( n36961 , n382071 );
buf ( n36962 , n381004 );
buf ( n36963 , n31719 );
and ( n36964 , n33098 , RI15b60af8_1164);
and ( n36965 , n31038 , n22443 );
nor ( n36966 , n36965 , RI15b3fab0_37);
nor ( n36967 , n36964 , n36966 );
not ( n36968 , n36967 );
buf ( n36969 , n36968 );
buf ( n36970 , n35649 );
buf ( n36971 , n33250 );
buf ( n36972 , n384218 );
or ( n36973 , n381907 , n35930 );
not ( n36974 , n35946 );
and ( n36975 , n36974 , RI15b40ed8_80);
or ( n36976 , n381917 , n35934 );
not ( n36977 , n35950 );
and ( n36978 , n36977 , n381923 );
and ( n36979 , n381926 , n35948 );
nor ( n36980 , n36978 , n36979 );
nand ( n36981 , n36976 , n36980 );
nor ( n36982 , n36975 , n36981 );
nand ( n36983 , n36973 , n36982 );
buf ( n36984 , n36983 );
or ( n36985 , n380968 , n35957 );
not ( n36986 , n35959 );
and ( n36987 , n380986 , n36986 );
not ( n36988 , RI15b40140_51);
or ( n36989 , n35967 , n36988 );
or ( n36990 , n380994 , n35973 );
or ( n36991 , n35965 , n380996 );
nand ( n36992 , n36989 , n36990 , n36991 );
nor ( n36993 , n36987 , n36992 );
nand ( n36994 , n36985 , n36993 );
buf ( n36995 , n36994 );
buf ( n36996 , n381006 );
buf ( n36997 , n32255 );
nor ( n36998 , n382080 , n382510 );
not ( n36999 , n36998 );
and ( n37000 , n36999 , RI15b47f58_320);
buf ( n37001 , n382525 );
and ( n37002 , n37001 , RI15b45f78_252);
nor ( n37003 , n37000 , n37002 );
not ( n37004 , n37003 );
buf ( n37005 , n37004 );
buf ( n37006 , n22009 );
buf ( n37007 , n31719 );
buf ( n37008 , n31979 );
not ( n37009 , n36813 );
not ( n37010 , n37009 );
not ( n37011 , n33174 );
or ( n37012 , n37010 , n37011 );
not ( n37013 , n36815 );
and ( n37014 , n33196 , n37013 );
not ( n37015 , RI15b423f0_125);
or ( n37016 , n36824 , n37015 );
or ( n37017 , n22241 , n36830 );
or ( n37018 , n36822 , n33201 );
nand ( n37019 , n37016 , n37017 , n37018 );
nor ( n37020 , n37014 , n37019 );
nand ( n37021 , n37012 , n37020 );
buf ( n37022 , n37021 );
buf ( n37023 , n382069 );
buf ( n37024 , n35649 );
buf ( n37025 , n19651 );
buf ( n37026 , n17499 );
buf ( n37027 , n387159 );
not ( n37028 , RI15b4b270_429);
or ( n37029 , n20613 , n37028 );
buf ( n37030 , n19954 );
not ( n37031 , n37030 );
not ( n37032 , n31806 );
or ( n37033 , n37031 , n37032 );
nand ( n37034 , n37033 , n380875 );
and ( n37035 , n37034 , RI15b49470_365);
or ( n37036 , n19722 , n19729 );
or ( n37037 , RI15b4a2f8_396 , RI15b4a370_397);
nand ( n37038 , n37036 , n37037 );
and ( n37039 , n22368 , n37038 );
nor ( n37040 , n37035 , n37039 );
and ( n37041 , n19939 , n32201 );
or ( n37042 , n20529 , n37030 , RI15b49470_365);
or ( n37043 , n382158 , RI15b4b270_429);
not ( n37044 , RI15b4b270_429);
or ( n37045 , n37044 , RI15b4b1f8_428);
nand ( n37046 , n37043 , n37045 );
and ( n37047 , n20566 , n37046 );
nand ( n37048 , n379830 , n379824 );
not ( n37049 , n36740 );
or ( n37050 , n37048 , n37049 );
not ( n37051 , RI15b4b270_429);
or ( n37052 , n37051 , n20639 );
nor ( n37053 , n19915 , RI15b4a280_395);
and ( n37054 , n37053 , n32199 );
and ( n37055 , n20652 , RI15b4a370_397);
nor ( n37056 , n37054 , n37055 );
nand ( n37057 , n37050 , n37052 , n37056 );
nor ( n37058 , n37047 , n37057 );
nand ( n37059 , n37042 , n37058 );
nor ( n37060 , n37041 , n37059 );
nand ( n37061 , n37029 , n37040 , n37060 );
buf ( n37062 , n37061 );
buf ( n37063 , n380942 );
or ( n37064 , n22473 , n386794 );
nand ( n37065 , n37064 , n383474 );
nand ( n37066 , n37065 , n36860 );
not ( n37067 , n36860 );
not ( n37068 , n34843 );
nand ( n37069 , n37067 , n37068 , n386794 );
not ( n37070 , RI15b63c30_1269);
buf ( n37071 , n387021 );
not ( n37072 , n37071 );
not ( n37073 , n37072 );
not ( n37074 , n22449 );
or ( n37075 , n37073 , n37074 );
nand ( n37076 , n37075 , n34811 );
not ( n37077 , n37076 );
or ( n37078 , n37070 , n37077 );
not ( n37079 , n386959 );
not ( n37080 , n37079 );
not ( n37081 , n34814 );
or ( n37082 , n37080 , n37081 );
nand ( n37083 , n37082 , n34823 );
and ( n37084 , n37083 , RI15b61e30_1205);
nor ( n37085 , n34826 , n37079 , RI15b61e30_1205);
or ( n37086 , n34833 , n37072 , RI15b63c30_1269);
or ( n37087 , n22470 , n31753 , n18859 );
nand ( n37088 , n37086 , n37087 );
nor ( n37089 , n37084 , n37085 , n37088 );
nand ( n37090 , n37078 , n37089 );
nand ( n37091 , n37090 , n19201 );
and ( n37092 , n22423 , RI15b63c30_1269);
and ( n37093 , n19599 , RI15b62d30_1237);
nor ( n37094 , n37092 , n37093 , n19513 );
nand ( n37095 , n37066 , n37069 , n37091 , n37094 );
buf ( n37096 , n37095 );
buf ( n37097 , n386762 );
buf ( n37098 , n22408 );
and ( n37099 , n22646 , RI15b45168_222);
and ( n37100 , n22648 , RI15b515d0_641);
nor ( n37101 , n37099 , n37100 );
not ( n37102 , n37101 );
buf ( n37103 , n37102 );
buf ( n37104 , n20663 );
buf ( n37105 , n22740 );
buf ( n37106 , n381490 );
not ( n37107 , RI15b4a118_392);
not ( n37108 , n37107 );
not ( n37109 , n36064 );
buf ( n37110 , n37109 );
buf ( n37111 , n37110 );
not ( n37112 , n37111 );
buf ( n37113 , n37112 );
buf ( n37114 , n37113 );
not ( n37115 , n37114 );
or ( n37116 , n37108 , n37115 );
not ( n37117 , n37113 );
nand ( n37118 , n36058 , RI15b49a88_378);
nor ( n37119 , n37118 , n32614 );
nand ( n37120 , n37119 , RI15b49b78_380);
not ( n37121 , RI15b49bf0_381);
nor ( n37122 , n37120 , n37121 );
nand ( n37123 , n37122 , RI15b49c68_382);
nor ( n37124 , n37123 , n19985 );
nand ( n37125 , n37124 , RI15b49d58_384);
nor ( n37126 , n37125 , n19988 );
nand ( n37127 , n37126 , RI15b49e48_386);
not ( n37128 , RI15b49ec0_387);
nor ( n37129 , n37127 , n37128 );
nand ( n37130 , n37129 , RI15b49f38_388);
nor ( n37131 , n37130 , n19995 );
nand ( n37132 , n37131 , RI15b4a028_390);
not ( n37133 , n37132 );
or ( n37134 , n37117 , n37133 );
nand ( n37135 , n37134 , n381056 );
nor ( n37136 , n37111 , RI15b4a0a0_391);
nor ( n37137 , n37135 , n37136 );
nand ( n37138 , n37116 , n37137 );
not ( n37139 , n37138 );
not ( n37140 , RI15b4a190_393);
or ( n37141 , n37139 , n37140 );
not ( n37142 , RI15b414f0_93);
not ( n37143 , n35448 );
or ( n37144 , n37142 , n37143 );
nand ( n37145 , n35389 , RI15b423f0_125);
nand ( n37146 , n37144 , n37145 );
and ( n37147 , n35405 , RI15b405f0_61);
and ( n37148 , n383375 , RI15b409b0_69);
and ( n37149 , n35427 , RI15b418b0_101);
nor ( n37150 , n37147 , n37148 , n37149 );
and ( n37151 , n35393 , RI15b427b0_133);
and ( n37152 , n35415 , RI15b42b70_141);
and ( n37153 , n35412 , RI15b42030_117);
nor ( n37154 , n37151 , n37152 , n37153 );
and ( n37155 , n35436 , RI15b41130_85);
and ( n37156 , n35399 , RI15b40230_53);
nor ( n37157 , n37155 , n37156 );
and ( n37158 , n35410 , RI15b40d70_77);
and ( n37159 , n35422 , RI15b41c70_109);
nor ( n37160 , n37158 , n37159 );
nand ( n37161 , n37150 , n37154 , n37157 , n37160 );
or ( n37162 , n35378 , n20119 );
and ( n37163 , n385989 , RI15b42f30_149);
and ( n37164 , n386002 , RI15b436b0_165);
and ( n37165 , n385471 , RI15b43a70_173);
nor ( n37166 , n37163 , n37164 , n37165 );
nand ( n37167 , n37162 , n37166 );
and ( n37168 , n37167 , n35370 );
nor ( n37169 , n37146 , n37161 , n37168 );
not ( n37170 , n37169 );
nand ( n37171 , n35436 , RI15b411a8_86);
nand ( n37172 , n35399 , RI15b402a8_54);
not ( n37173 , n20041 );
and ( n37174 , n37173 , RI15b41568_94);
buf ( n37175 , n20036 );
and ( n37176 , n37175 , RI15b42468_126);
nor ( n37177 , n37174 , n37176 );
not ( n37178 , n20060 );
nand ( n37179 , n37178 , RI15b43368_158);
nand ( n37180 , n37171 , n37172 , n37177 , n37179 );
nand ( n37181 , n35393 , RI15b42828_134);
nand ( n37182 , n35412 , RI15b420a8_118);
nand ( n37183 , n35410 , RI15b40de8_78);
nand ( n37184 , n35422 , RI15b41ce8_110);
nand ( n37185 , n37181 , n37182 , n37183 , n37184 );
nor ( n37186 , n37180 , n37185 );
not ( n37187 , n385339 );
and ( n37188 , n37187 , RI15b43728_166);
and ( n37189 , n383376 , RI15b40a28_70);
nor ( n37190 , n37188 , n37189 );
and ( n37191 , n35415 , RI15b42be8_142);
not ( n37192 , n20056 );
and ( n37193 , n37192 , RI15b42fa8_150);
and ( n37194 , n35405 , RI15b40668_62);
nor ( n37195 , n37191 , n37193 , n37194 );
and ( n37196 , n35428 , RI15b41928_102);
not ( n37197 , n35369 );
and ( n37198 , n37197 , RI15b3fee8_46);
nor ( n37199 , n37196 , n37198 );
nand ( n37200 , n37186 , n37190 , n37195 , n37199 );
nand ( n37201 , n37170 , n37200 );
and ( n37202 , n35400 , RI15b40320_55);
and ( n37203 , n37173 , RI15b415e0_95);
buf ( n37204 , n37175 );
and ( n37205 , n37204 , RI15b424e0_127);
nor ( n37206 , n37202 , n37203 , n37205 );
and ( n37207 , n35412 , RI15b42120_119);
and ( n37208 , n35394 , RI15b428a0_135);
nor ( n37209 , n37207 , n37208 );
and ( n37210 , n35437 , RI15b41220_87);
and ( n37211 , n37178 , RI15b433e0_159);
nor ( n37212 , n37210 , n37211 );
and ( n37213 , n35410 , RI15b40e60_79);
and ( n37214 , n35422 , RI15b41d60_111);
nor ( n37215 , n37213 , n37214 );
nand ( n37216 , n37206 , n37209 , n37212 , n37215 );
and ( n37217 , n37192 , RI15b43020_151);
and ( n37218 , n35406 , RI15b406e0_63);
and ( n37219 , n35415 , RI15b42c60_143);
nor ( n37220 , n37217 , n37218 , n37219 );
buf ( n37221 , n37187 );
and ( n37222 , n37221 , RI15b437a0_167);
and ( n37223 , n383377 , RI15b40aa0_71);
nor ( n37224 , n37222 , n37223 );
and ( n37225 , n35429 , RI15b419a0_103);
and ( n37226 , n37197 , RI15b3ff60_47);
nor ( n37227 , n37225 , n37226 );
nand ( n37228 , n37220 , n37224 , n37227 );
nor ( n37229 , n37216 , n37228 );
or ( n37230 , n37201 , n37229 );
not ( n37231 , n37230 );
and ( n37232 , n35401 , RI15b40398_56);
and ( n37233 , n37173 , RI15b41658_96);
buf ( n37234 , n37204 );
and ( n37235 , n37234 , RI15b42558_128);
nor ( n37236 , n37232 , n37233 , n37235 );
and ( n37237 , n35438 , RI15b41298_88);
and ( n37238 , n37178 , RI15b43458_160);
nor ( n37239 , n37237 , n37238 );
and ( n37240 , n35412 , RI15b42198_120);
and ( n37241 , n35395 , RI15b42918_136);
nor ( n37242 , n37240 , n37241 );
and ( n37243 , n35410 , RI15b40ed8_80);
and ( n37244 , n35422 , RI15b41dd8_112);
nor ( n37245 , n37243 , n37244 );
and ( n37246 , n37236 , n37239 , n37242 , n37245 );
and ( n37247 , n37192 , RI15b43098_152);
and ( n37248 , n35407 , RI15b40758_64);
and ( n37249 , n35415 , RI15b42cd8_144);
nor ( n37250 , n37247 , n37248 , n37249 );
buf ( n37251 , n37221 );
and ( n37252 , n37251 , RI15b43818_168);
and ( n37253 , n383378 , RI15b40b18_72);
nor ( n37254 , n37252 , n37253 );
and ( n37255 , n35430 , RI15b41a18_104);
and ( n37256 , n37197 , RI15b3ffd8_48);
nor ( n37257 , n37255 , n37256 );
nand ( n37258 , n37246 , n37250 , n37254 , n37257 );
nand ( n37259 , n37231 , n37258 );
and ( n37260 , n35557 , RI15b40410_57);
and ( n37261 , n37173 , RI15b416d0_97);
buf ( n37262 , n37234 );
and ( n37263 , n37262 , RI15b425d0_129);
nor ( n37264 , n37260 , n37261 , n37263 );
and ( n37265 , n35439 , RI15b41310_89);
and ( n37266 , n37178 , RI15b434d0_161);
nor ( n37267 , n37265 , n37266 );
and ( n37268 , n35412 , RI15b42210_121);
and ( n37269 , n35396 , RI15b42990_137);
nor ( n37270 , n37268 , n37269 );
and ( n37271 , n35410 , RI15b40f50_81);
and ( n37272 , n35422 , RI15b41e50_113);
nor ( n37273 , n37271 , n37272 );
nand ( n37274 , n37264 , n37267 , n37270 , n37273 );
and ( n37275 , n37192 , RI15b43110_153);
and ( n37276 , n35552 , RI15b407d0_65);
and ( n37277 , n35415 , RI15b42d50_145);
nor ( n37278 , n37275 , n37276 , n37277 );
buf ( n37279 , n37251 );
and ( n37280 , n37279 , RI15b43890_169);
and ( n37281 , n383378 , RI15b40b90_73);
nor ( n37282 , n37280 , n37281 );
and ( n37283 , n35430 , RI15b41a90_105);
and ( n37284 , n37197 , RI15b40050_49);
nor ( n37285 , n37283 , n37284 );
nand ( n37286 , n37278 , n37282 , n37285 );
nor ( n37287 , n37274 , n37286 );
or ( n37288 , n37259 , n37287 );
not ( n37289 , n37288 );
and ( n37290 , n35557 , RI15b40488_58);
and ( n37291 , n37173 , RI15b41748_98);
and ( n37292 , n37262 , RI15b42648_130);
nor ( n37293 , n37290 , n37291 , n37292 );
not ( n37294 , n35440 );
and ( n37295 , n37294 , RI15b41388_90);
and ( n37296 , n37178 , RI15b43548_162);
nor ( n37297 , n37295 , n37296 );
and ( n37298 , n35410 , RI15b40fc8_82);
and ( n37299 , RI15b41ec8_114 , n35422 );
nor ( n37300 , n37298 , n37299 );
and ( n37301 , n35412 , RI15b42288_122);
buf ( n37302 , n35396 );
and ( n37303 , n37302 , RI15b42a08_138);
nor ( n37304 , n37301 , n37303 );
nand ( n37305 , n37293 , n37297 , n37300 , n37304 );
not ( n37306 , n37305 );
and ( n37307 , n35553 , RI15b40848_66);
and ( n37308 , n35415 , RI15b42dc8_146);
and ( n37309 , n37192 , RI15b43188_154);
nor ( n37310 , n37307 , n37308 , n37309 );
not ( n37311 , n35431 );
buf ( n37312 , n37311 );
and ( n37313 , n37312 , RI15b41b08_106);
and ( n37314 , n37197 , RI15b400c8_50);
nor ( n37315 , n37313 , n37314 );
buf ( n37316 , n37279 );
and ( n37317 , n37316 , RI15b43908_170);
and ( n37318 , n383379 , RI15b40c08_74);
nor ( n37319 , n37317 , n37318 );
nand ( n37320 , n37306 , n37310 , n37315 , n37319 );
nand ( n37321 , n37289 , n37320 );
buf ( n37322 , n35557 );
buf ( n37323 , n37322 );
and ( n37324 , n37323 , RI15b40500_59);
and ( n37325 , n37173 , RI15b417c0_99);
buf ( n37326 , n37262 );
and ( n37327 , n37326 , RI15b426c0_131);
nor ( n37328 , n37324 , n37325 , n37327 );
buf ( n37329 , n35441 );
and ( n37330 , n37329 , RI15b41400_91);
and ( n37331 , n37178 , RI15b435c0_163);
nor ( n37332 , n37330 , n37331 );
and ( n37333 , n35410 , RI15b41040_83);
and ( n37334 , n35422 , RI15b41f40_115);
nor ( n37335 , n37333 , n37334 );
and ( n37336 , n35412 , RI15b42300_123);
buf ( n37337 , n37302 );
and ( n37338 , n37337 , RI15b42a80_139);
nor ( n37339 , n37336 , n37338 );
nand ( n37340 , n37328 , n37332 , n37335 , n37339 );
and ( n37341 , n37192 , RI15b43200_155);
buf ( n37342 , n35553 );
and ( n37343 , n37342 , RI15b408c0_67);
and ( n37344 , n35415 , RI15b42e40_147);
nor ( n37345 , n37341 , n37343 , n37344 );
buf ( n37346 , n37316 );
and ( n37347 , n37346 , RI15b43980_171);
and ( n37348 , n383380 , RI15b40c80_75);
nor ( n37349 , n37347 , n37348 );
buf ( n37350 , n37312 );
and ( n37351 , n37350 , RI15b41b80_107);
and ( n37352 , n37197 , RI15b40140_51);
nor ( n37353 , n37351 , n37352 );
nand ( n37354 , n37345 , n37349 , n37353 );
nor ( n37355 , n37340 , n37354 );
nor ( n37356 , n37321 , n37355 );
and ( n37357 , n37323 , RI15b40578_60);
and ( n37358 , n37173 , RI15b41838_100);
and ( n37359 , n37326 , RI15b42738_132);
nor ( n37360 , n37357 , n37358 , n37359 );
and ( n37361 , n37329 , RI15b41478_92);
and ( n37362 , n37178 , RI15b43638_164);
nor ( n37363 , n37361 , n37362 );
and ( n37364 , n35410 , RI15b410b8_84);
and ( n37365 , n35422 , RI15b41fb8_116);
nor ( n37366 , n37364 , n37365 );
and ( n37367 , n35412 , RI15b42378_124);
and ( n37368 , n37337 , RI15b42af8_140);
nor ( n37369 , n37367 , n37368 );
nand ( n37370 , n37360 , n37363 , n37366 , n37369 );
not ( n37371 , n37370 );
and ( n37372 , n37192 , RI15b43278_156);
buf ( n37373 , n37342 );
and ( n37374 , n37373 , RI15b40938_68);
and ( n37375 , n35415 , RI15b42eb8_148);
nor ( n37376 , n37372 , n37374 , n37375 );
buf ( n37377 , n37350 );
and ( n37378 , n37377 , RI15b41bf8_108);
and ( n37379 , n37197 , RI15b401b8_52);
nor ( n37380 , n37378 , n37379 );
buf ( n37381 , n37346 );
and ( n37382 , n37381 , RI15b439f8_172);
not ( n37383 , n383382 );
and ( n37384 , n37383 , RI15b40cf8_76);
nor ( n37385 , n37382 , n37384 );
nand ( n37386 , n37371 , n37376 , n37380 , n37385 );
nand ( n37387 , n37356 , n37386 );
not ( n37388 , n37387 );
and ( n37389 , n37329 , RI15b414f0_93);
and ( n37390 , n37178 , RI15b436b0_165);
nor ( n37391 , n37389 , n37390 );
and ( n37392 , n37323 , RI15b405f0_61);
and ( n37393 , n37173 , RI15b418b0_101);
and ( n37394 , n37326 , RI15b427b0_133);
nor ( n37395 , n37392 , n37393 , n37394 );
and ( n37396 , n35410 , RI15b41130_85);
and ( n37397 , n35422 , RI15b42030_117);
nor ( n37398 , n37396 , n37397 );
and ( n37399 , n35412 , RI15b423f0_125);
and ( n37400 , n37337 , RI15b42b70_141);
nor ( n37401 , n37399 , n37400 );
nand ( n37402 , n37391 , n37395 , n37398 , n37401 );
not ( n37403 , n37402 );
and ( n37404 , n37192 , RI15b432f0_157);
and ( n37405 , n37373 , RI15b409b0_69);
and ( n37406 , n35415 , RI15b42f30_149);
nor ( n37407 , n37404 , n37405 , n37406 );
and ( n37408 , n37377 , RI15b41c70_109);
and ( n37409 , n37197 , RI15b40230_53);
nor ( n37410 , n37408 , n37409 );
and ( n37411 , n37381 , RI15b43a70_173);
and ( n37412 , n383384 , RI15b40d70_77);
nor ( n37413 , n37411 , n37412 );
nand ( n37414 , n37403 , n37407 , n37410 , n37413 );
not ( n37415 , n37414 );
and ( n37416 , n37388 , n37415 );
and ( n37417 , n37387 , n37414 );
nor ( n37418 , n37416 , n37417 );
not ( n37419 , n37418 );
not ( n37420 , n381062 );
and ( n37421 , n37419 , n37420 );
not ( n37422 , n37132 );
not ( n37423 , n37113 );
not ( n37424 , RI15b4a0a0_391);
nor ( n37425 , n37423 , n37424 );
and ( n37426 , n37422 , n37425 );
nor ( n37427 , n37107 , RI15b4a190_393);
and ( n37428 , n37426 , n37427 );
nor ( n37429 , n37421 , n37428 );
nand ( n37430 , n37141 , n37429 );
buf ( n37431 , n37430 );
buf ( n37432 , n382049 );
not ( n37433 , RI15b53718_712);
not ( n37434 , n32244 );
or ( n37435 , n37433 , n37434 );
and ( n37436 , n32247 , RI15b64d10_1305);
and ( n37437 , n32249 , RI15b5fb80_1131);
nor ( n37438 , n37436 , n37437 );
nand ( n37439 , n37435 , n37438 );
buf ( n37440 , n37439 );
buf ( n37441 , n22009 );
buf ( n37442 , n386730 );
not ( n37443 , n37442 );
or ( n37444 , n32430 , n37443 );
nand ( n37445 , n381417 , n381355 );
and ( n37446 , n34900 , RI15b54ac8_754);
buf ( n37447 , n21624 );
and ( n37448 , n382885 , n37447 );
buf ( n37449 , n382626 );
not ( n37450 , RI15b54a50_753);
or ( n37451 , n34896 , n37450 , RI15b54ac8_754);
not ( n37452 , RI15b54ac8_754);
or ( n37453 , n37452 , RI15b54a50_753);
nand ( n37454 , n37451 , n37453 );
and ( n37455 , n37449 , n37454 );
nor ( n37456 , n37446 , n37448 , n37455 );
and ( n37457 , n37445 , n37456 );
nand ( n37458 , n37444 , n37457 );
buf ( n37459 , n37458 );
buf ( n37460 , n22408 );
not ( n37461 , n32064 );
not ( n37462 , n33400 );
or ( n37463 , n37461 , n37462 );
and ( n37464 , n33415 , n32070 );
or ( n37465 , n32081 , n18488 );
or ( n37466 , n36293 , n32086 );
or ( n37467 , n32079 , n33443 );
nand ( n37468 , n37465 , n37466 , n37467 );
nor ( n37469 , n37464 , n37468 );
nand ( n37470 , n37463 , n37469 );
buf ( n37471 , n37470 );
buf ( n37472 , n382065 );
and ( n37473 , n22646 , RI15b45d20_247);
and ( n37474 , n22648 , RI15b52188_666);
nor ( n37475 , n37473 , n37474 );
not ( n37476 , n37475 );
buf ( n37477 , n37476 );
not ( n37478 , n384960 );
or ( n37479 , n37478 , n36200 );
and ( n37480 , n384983 , n36202 );
or ( n37481 , n36212 , n385392 );
or ( n37482 , n22022 , n36217 );
or ( n37483 , n36210 , n384988 );
nand ( n37484 , n37481 , n37482 , n37483 );
nor ( n37485 , n37480 , n37484 );
nand ( n37486 , n37479 , n37485 );
buf ( n37487 , n37486 );
buf ( n37488 , n383345 );
buf ( n37489 , n19653 );
buf ( n37490 , n32271 );
buf ( n37491 , n383613 );
buf ( n37492 , n379844 );
buf ( n37493 , n22740 );
buf ( n37494 , n380903 );
or ( n37495 , n380908 , n22150 );
or ( n37496 , n384961 , n37495 );
nand ( n37497 , n22140 , n35903 );
not ( n37498 , n37497 );
and ( n37499 , n384983 , n37498 );
and ( n37500 , n37495 , n37497 , n19912 );
nor ( n37501 , n37500 , n22217 );
nor ( n37502 , n380918 , n22133 );
or ( n37503 , n37501 , n37502 );
nand ( n37504 , n37503 , n20623 );
or ( n37505 , n380924 , n32180 );
and ( n37506 , n37504 , n37505 );
nor ( n37507 , n37506 , n22236 );
not ( n37508 , RI15b42738_132);
or ( n37509 , n37507 , n37508 );
not ( n37510 , n37505 );
nor ( n37511 , n37502 , n37510 );
or ( n37512 , n37501 , n37511 );
or ( n37513 , n22022 , n37512 );
or ( n37514 , n37505 , n384988 );
nand ( n37515 , n37509 , n37513 , n37514 );
nor ( n37516 , n37499 , n37515 );
nand ( n37517 , n37496 , n37516 );
buf ( n37518 , n37517 );
buf ( n37519 , n386760 );
nand ( n37520 , n381406 , n35490 );
not ( n37521 , n381384 );
nand ( n37522 , n381417 , n37521 );
nand ( n37523 , n381486 , RI15b52f20_695);
not ( n37524 , n381439 );
not ( n37525 , n36268 );
or ( n37526 , n37524 , n37525 );
nand ( n37527 , n37526 , n381450 );
not ( n37528 , n381446 );
and ( n37529 , n37527 , n37528 );
nor ( n37530 , n381439 , n37528 );
and ( n37531 , n381461 , n37530 );
nor ( n37532 , n37529 , n37531 );
nand ( n37533 , n37520 , n37522 , n37523 , n37532 );
buf ( n37534 , n37533 );
not ( n37535 , n381494 );
not ( n37536 , n380703 );
or ( n37537 , n37535 , n37536 );
and ( n37538 , n380719 , n381528 );
not ( n37539 , RI15b5bf80_1003);
or ( n37540 , n381544 , n37539 );
buf ( n37541 , n380780 );
not ( n37542 , n37541 );
or ( n37543 , n37542 , n381557 );
or ( n37544 , n381542 , n380790 );
nand ( n37545 , n37540 , n37543 , n37544 );
nor ( n37546 , n37538 , n37545 );
nand ( n37547 , n37537 , n37546 );
buf ( n37548 , n37547 );
buf ( n37549 , n22404 );
buf ( n37550 , n31719 );
buf ( n37551 , n32672 );
buf ( n37552 , n22653 );
not ( n37553 , n386536 );
buf ( n37554 , n383371 );
or ( n37555 , n37553 , n37554 );
or ( n37556 , n385203 , n386534 );
nand ( n37557 , n37556 , RI15b47ee0_319);
and ( n37558 , n20416 , n379824 );
nor ( n37559 , n37558 , n22232 );
nand ( n37560 , n37555 , n37557 , n37559 );
buf ( n37561 , n37560 );
buf ( n37562 , n31033 );
buf ( n37563 , n379844 );
buf ( n37564 , n384203 );
buf ( n37565 , n19655 );
nor ( n37566 , RI15b54780_747 , RI15b54870_749);
nor ( n37567 , n379391 , n37566 );
or ( n37568 , n37567 , RI15b543c0_739);
not ( n37569 , n379396 );
and ( n37570 , n37569 , RI15b52368_670);
and ( n37571 , n35233 , n379339 );
nor ( n37572 , n37570 , n37571 );
nand ( n37573 , n37568 , n37572 );
buf ( n37574 , n37573 );
not ( n37575 , n384274 );
not ( n37576 , n37575 );
not ( n37577 , n32540 );
nand ( n37578 , n37577 , n384283 );
not ( n37579 , n37578 );
or ( n37580 , n37576 , n37579 );
buf ( n37581 , n32541 );
not ( n37582 , n37581 );
nand ( n37583 , n37580 , n37582 );
and ( n37584 , n37583 , n31921 );
not ( n37585 , n32555 );
not ( n37586 , n37585 );
not ( n37587 , n384582 );
not ( n37588 , n37587 );
and ( n37589 , n37586 , n37588 );
and ( n37590 , n37585 , n37587 );
nor ( n37591 , n37589 , n37590 );
or ( n37592 , n37591 , n31958 );
not ( n37593 , n384446 );
not ( n37594 , n37593 );
not ( n37595 , n384443 );
or ( n37596 , n37594 , n37595 );
or ( n37597 , n384443 , n37593 );
nand ( n37598 , n37596 , n37597 );
buf ( n37599 , n380838 );
and ( n37600 , n37598 , n37599 );
and ( n37601 , n19513 , RI15b641d0_1281);
nor ( n37602 , n37600 , n37601 );
nand ( n37603 , n37592 , n37602 );
nor ( n37604 , n37584 , n37603 );
or ( n37605 , n384398 , n31751 );
nand ( n37606 , n37605 , n31771 );
and ( n37607 , n37606 , RI15b5cb38_1028);
and ( n37608 , n31792 , n384582 );
or ( n37609 , n31779 , n384448 , RI15b5cb38_1028);
not ( n37610 , n32377 );
not ( n37611 , n37610 );
or ( n37612 , n37611 , n384274 );
nand ( n37613 , n37609 , n37612 );
nor ( n37614 , n37607 , n37608 , n37613 );
nand ( n37615 , n37604 , n37614 );
buf ( n37616 , n37615 );
buf ( n37617 , n381004 );
not ( n37618 , n32680 );
not ( n37619 , n380645 );
nand ( n37620 , n380624 , n37619 );
not ( n37621 , n37620 );
nand ( n37622 , n380683 , n380648 );
nand ( n37623 , n37621 , n37622 );
not ( n37624 , n37622 );
nand ( n37625 , n37620 , n37624 );
not ( n37626 , n381496 );
not ( n37627 , n37626 );
nand ( n37628 , n37623 , n37625 , n37627 );
not ( n37629 , n37628 );
not ( n37630 , n37629 );
or ( n37631 , n37618 , n37630 );
nand ( n37632 , n33410 , n381522 );
nor ( n37633 , n382919 , n37632 );
or ( n37634 , n382917 , n386594 , n382920 );
or ( n37635 , n382926 , n380597 );
nand ( n37636 , n37634 , n37635 );
or ( n37637 , n37633 , n37636 );
and ( n37638 , n37637 , n35222 );
or ( n37639 , n32692 , n18979 );
buf ( n37640 , n380321 );
not ( n37641 , n37640 );
buf ( n37642 , n37641 );
buf ( n37643 , n37642 );
not ( n37644 , n37643 );
or ( n37645 , n37644 , n32699 );
nand ( n37646 , n19519 , n380789 );
or ( n37647 , n32690 , n37646 );
nand ( n37648 , n37639 , n37645 , n37647 );
nor ( n37649 , n37638 , n37648 );
nand ( n37650 , n37631 , n37649 );
buf ( n37651 , n37650 );
buf ( n37652 , n22007 );
or ( n37653 , n385032 , n379340 );
and ( n37654 , n35236 , RI15b54258_736 , RI15b54780_747);
nor ( n37655 , n37654 , n18096 );
nand ( n37656 , n37653 , n35245 , n37655 );
buf ( n37657 , n37656 );
buf ( n37658 , n379802 );
buf ( n37659 , n382069 );
buf ( n37660 , n381566 );
buf ( n37661 , n381021 );
buf ( n37662 , n18226 );
or ( n37663 , n380908 , n380925 );
or ( n37664 , n380968 , n37663 );
nand ( n37665 , n22140 , n22134 );
not ( n37666 , n37665 );
and ( n37667 , n380986 , n37666 );
and ( n37668 , n37663 , n37665 , n19912 );
nor ( n37669 , n37668 , n22217 );
nor ( n37670 , n380918 , n35878 );
or ( n37671 , n37669 , n37670 );
nand ( n37672 , n37671 , n20623 );
or ( n37673 , n380924 , n22150 );
and ( n37674 , n37672 , n37673 );
nor ( n37675 , n37674 , n22236 );
or ( n37676 , n37675 , n385475 );
not ( n37677 , n37673 );
nor ( n37678 , n37670 , n37677 );
or ( n37679 , n37669 , n37678 );
or ( n37680 , n380994 , n37679 );
or ( n37681 , n37673 , n380996 );
nand ( n37682 , n37676 , n37680 , n37681 );
nor ( n37683 , n37667 , n37682 );
nand ( n37684 , n37664 , n37683 );
buf ( n37685 , n37684 );
buf ( n37686 , n32672 );
buf ( n37687 , n381566 );
buf ( n37688 , n33250 );
and ( n37689 , n36764 , n20501 );
and ( n37690 , n20519 , RI15b44c40_211);
nor ( n37691 , n37689 , n37690 );
not ( n37692 , n37691 );
buf ( n37693 , n37692 );
buf ( n37694 , n382067 );
buf ( n37695 , n379893 );
buf ( n37696 , n381566 );
nand ( n37697 , n18116 , n21556 );
nand ( n37698 , n381467 , n37697 );
nand ( n37699 , n37698 , n18077 , n21402 );
not ( n37700 , n18126 );
or ( n37701 , n18122 , n382542 );
not ( n37702 , n37701 );
or ( n37703 , n37700 , n37702 );
nand ( n37704 , n37703 , n18077 );
or ( n37705 , n18185 , n381476 );
nand ( n37706 , n37705 , n18077 );
nand ( n37707 , n37706 , n385161 );
not ( n37708 , n37707 );
nand ( n37709 , n37704 , n37708 , n381481 , n18164 );
nand ( n37710 , n37709 , RI15b4ff50_593);
or ( n37711 , n21198 , RI15b4ff50_593);
not ( n37712 , n21203 );
nand ( n37713 , n37711 , n37712 );
and ( n37714 , n21559 , n37713 );
and ( n37715 , n21751 , RI15b575e8_846);
nor ( n37716 , n37714 , n37715 );
not ( n37717 , n381472 );
not ( n37718 , n21403 );
or ( n37719 , n21349 , n37718 );
or ( n37720 , n21402 , n21350 );
nand ( n37721 , n21603 , RI15b4ff50_593);
nand ( n37722 , n37719 , n37720 , n37721 );
nand ( n37723 , n37717 , n37722 );
nand ( n37724 , n37699 , n37710 , n37716 , n37723 );
buf ( n37725 , n37724 );
not ( n37726 , n33575 );
nand ( n37727 , n33540 , n37726 );
not ( n37728 , n37727 );
and ( n37729 , n383523 , RI15b61a70_1197);
not ( n37730 , n383523 );
nor ( n37731 , n33531 , n33507 );
not ( n37732 , n37731 );
buf ( n37733 , n33520 );
not ( n37734 , n37733 );
not ( n37735 , n37734 );
not ( n37736 , n33516 );
nor ( n37737 , RI15b619f8_1196 , RI15b61a70_1197);
nand ( n37738 , n33516 , n37737 );
nand ( n37739 , RI15b619f8_1196 , RI15b61a70_1197);
and ( n37740 , n37738 , n37739 );
not ( n37741 , n37740 );
or ( n37742 , n37736 , n37741 );
nor ( n37743 , n33527 , RI15b61a70_1197);
not ( n37744 , n37743 );
not ( n37745 , n37738 );
or ( n37746 , n37744 , n37745 );
nand ( n37747 , n33512 , RI15b61a70_1197);
nand ( n37748 , n37746 , n37747 );
not ( n37749 , n37748 );
nand ( n37750 , n37742 , n37749 );
not ( n37751 , n37750 );
or ( n37752 , n37735 , n37751 );
not ( n37753 , RI15b61a70_1197);
not ( n37754 , n33524 );
or ( n37755 , n37753 , n37754 );
nand ( n37756 , n37755 , n37740 );
and ( n37757 , n37756 , n37733 );
buf ( n37758 , n37738 );
not ( n37759 , n37758 );
buf ( n37760 , n33512 );
and ( n37761 , n37759 , n37760 );
nor ( n37762 , n37757 , n37761 );
nand ( n37763 , n37752 , n37762 );
not ( n37764 , n37763 );
or ( n37765 , n37732 , n37764 );
nor ( n37766 , n33531 , n33507 );
or ( n37767 , n37766 , n37763 );
nand ( n37768 , n37765 , n37767 );
and ( n37769 , n37730 , n37768 );
nor ( n37770 , n37729 , n37769 );
nand ( n37771 , n37728 , n37770 );
buf ( n37772 , n384922 );
buf ( n37773 , n37772 );
not ( n37774 , n37773 );
not ( n37775 , n37774 );
not ( n37776 , n37775 );
buf ( n37777 , n37776 );
nor ( n37778 , n37771 , n37777 );
not ( n37779 , n32343 );
not ( n37780 , n37779 );
not ( n37781 , n37780 );
buf ( n37782 , n37781 );
buf ( n37783 , n37782 );
or ( n37784 , n37778 , n37783 );
not ( n37785 , RI15b61ae8_1198);
buf ( n37786 , n37758 );
nand ( n37787 , n37786 , RI15b61bd8_1200);
not ( n37788 , n37787 );
or ( n37789 , n37785 , n37788 );
or ( n37790 , n37787 , RI15b61ae8_1198);
nand ( n37791 , n37789 , n37790 );
buf ( n37792 , n37791 );
nand ( n37793 , n37784 , n37792 );
nor ( n37794 , n37791 , n384933 );
not ( n37795 , n37794 );
not ( n37796 , n37771 );
or ( n37797 , n37795 , n37796 );
and ( n37798 , n384918 , RI15b5ef50_1105);
buf ( n37799 , n384782 );
nand ( n37800 , n384906 , n37799 );
not ( n37801 , n37800 );
nor ( n37802 , n37798 , n37801 );
nand ( n37803 , n37797 , n37802 );
not ( n37804 , n37803 );
nand ( n37805 , n37793 , n37804 );
buf ( n37806 , n37805 );
buf ( n37807 , n381004 );
not ( n37808 , n37772 );
not ( n37809 , n33560 );
not ( n37810 , n37809 );
or ( n37811 , n37808 , n37810 );
nand ( n37812 , n37811 , n32343 );
nand ( n37813 , n37812 , n33567 );
nor ( n37814 , n37809 , n33567 );
nand ( n37815 , n37814 , n384934 );
nand ( n37816 , n384918 , RI15b5ec80_1099);
nand ( n37817 , n384906 , n380779 );
nand ( n37818 , n37813 , n37815 , n37816 , n37817 );
buf ( n37819 , n37818 );
buf ( n37820 , n379893 );
or ( n37821 , n385163 , n20911 );
not ( n37822 , n21586 );
not ( n37823 , n21599 );
not ( n37824 , n37823 );
buf ( n37825 , n21620 );
not ( n37826 , n37825 );
or ( n37827 , n37824 , n37826 );
nand ( n37828 , n37827 , n21625 );
not ( n37829 , n21629 );
or ( n37830 , n37828 , n37829 );
nand ( n37831 , n37830 , n21582 );
buf ( n37832 , n20908 );
buf ( n37833 , n37832 );
not ( n37834 , n37833 );
not ( n37835 , n37834 );
and ( n37836 , n37831 , n37835 );
not ( n37837 , n21582 );
not ( n37838 , n37828 );
or ( n37839 , n37837 , n37838 );
nand ( n37840 , n37839 , n21629 );
and ( n37841 , n37840 , n37834 );
nor ( n37842 , n37836 , n37841 );
not ( n37843 , n37842 );
or ( n37844 , n37822 , n37843 );
or ( n37845 , n37842 , n21586 );
nand ( n37846 , n37844 , n37845 );
and ( n37847 , n37846 , n21746 );
not ( n37848 , n22667 );
not ( n37849 , n37833 );
and ( n37850 , n21428 , n37849 );
not ( n37851 , n21428 );
and ( n37852 , n37851 , n37833 );
nor ( n37853 , n37850 , n37852 );
not ( n37854 , n37853 );
and ( n37855 , n37848 , n37854 );
and ( n37856 , n22667 , n37853 );
nor ( n37857 , n37855 , n37856 );
or ( n37858 , n37857 , n21561 );
not ( n37859 , n20919 );
buf ( n37860 , n21223 );
not ( n37861 , n21227 );
or ( n37862 , n37860 , n37861 );
nand ( n37863 , n37862 , n20963 );
and ( n37864 , n37863 , n37832 );
not ( n37865 , n37832 );
and ( n37866 , n21228 , n37865 );
nor ( n37867 , n37864 , n37866 );
not ( n37868 , n37867 );
or ( n37869 , n37859 , n37868 );
or ( n37870 , n37867 , n20919 );
nand ( n37871 , n37869 , n37870 );
and ( n37872 , n37871 , n21355 );
and ( n37873 , n21751 , RI15b578b8_852);
nor ( n37874 , n37872 , n37873 );
nand ( n37875 , n37858 , n37874 );
nor ( n37876 , n37847 , n37875 );
not ( n37877 , n36472 );
not ( n37878 , n37877 );
and ( n37879 , n37878 , n21586 );
and ( n37880 , n32368 , n20919 );
and ( n37881 , n385177 , n21428 );
nor ( n37882 , n37879 , n37880 , n37881 );
nand ( n37883 , n37821 , n37876 , n37882 );
buf ( n37884 , n37883 );
buf ( n37885 , n17499 );
nand ( n37886 , n21836 , n17507 );
not ( n37887 , n37886 );
not ( n37888 , n17565 );
or ( n37889 , n37887 , n37888 );
nand ( n37890 , n37889 , n21810 );
nor ( n37891 , n21836 , n21810 );
nand ( n37892 , n385056 , n37891 );
not ( n37893 , RI15b57930_853);
not ( n37894 , n34667 );
or ( n37895 , n37893 , n37894 );
buf ( n37896 , n21956 );
not ( n37897 , n37896 );
or ( n37898 , n18074 , n37897 );
nand ( n37899 , n37898 , n21979 );
and ( n37900 , n37899 , RI15b55b30_789);
or ( n37901 , n21982 , n37896 , RI15b55b30_789);
and ( n37902 , n21927 , n379110 , RI15b578b8_852);
and ( n37903 , n379108 , RI15b57930_853);
nor ( n37904 , n37902 , n37903 );
or ( n37905 , n21922 , n37904 );
nand ( n37906 , n37901 , n37905 );
nor ( n37907 , n37900 , n37906 );
nand ( n37908 , n37895 , n37907 );
and ( n37909 , n37908 , n18077 );
or ( n37910 , n18178 , n379110 );
or ( n37911 , n21803 , n18218 );
nand ( n37912 , n37910 , n37911 , n21750 );
nor ( n37913 , n37909 , n37912 );
nand ( n37914 , n37890 , n37892 , n37913 );
buf ( n37915 , n37914 );
buf ( n37916 , n22007 );
buf ( n37917 , n36704 );
nand ( n37918 , n36659 , n36666 );
nand ( n37919 , n36632 , RI15b50ce8_622);
nor ( n37920 , n37919 , RI15b50d60_623);
and ( n37921 , n37920 , n20691 );
and ( n37922 , n20692 , RI15b50d60_623);
and ( n37923 , n37919 , RI15b50d60_623);
nor ( n37924 , n37921 , n37922 , n37923 );
nor ( n37925 , n37918 , n37924 );
not ( n37926 , n37925 );
not ( n37927 , RI15b50dd8_624);
or ( n37928 , n20691 , n37927 );
not ( n37929 , RI15b50d60_623);
nor ( n37930 , n37919 , n37929 );
nand ( n37931 , n37930 , n37927 );
or ( n37932 , n20692 , n37931 );
not ( n37933 , n37930 );
nand ( n37934 , n37933 , RI15b50dd8_624);
nand ( n37935 , n37928 , n37932 , n37934 );
not ( n37936 , n37935 );
and ( n37937 , n37926 , n37936 );
and ( n37938 , n37925 , n37935 );
nor ( n37939 , n37937 , n37938 );
buf ( n37940 , n22679 );
or ( n37941 , n37939 , n37940 );
not ( n37942 , n36680 );
buf ( n37943 , n37942 );
or ( n37944 , n37943 , n37927 );
not ( n37945 , n37943 );
or ( n37946 , n37945 , n37931 );
nand ( n37947 , n37944 , n37946 , n37934 );
not ( n37948 , n37947 );
not ( n37949 , n36687 );
and ( n37950 , n37942 , n37920 );
and ( n37951 , n36680 , RI15b50d60_623);
nor ( n37952 , n37950 , n37951 , n37923 );
nand ( n37953 , n37949 , n37952 );
not ( n37954 , n37953 );
not ( n37955 , n37954 );
or ( n37956 , n37948 , n37955 );
or ( n37957 , n37954 , n37947 );
nand ( n37958 , n37956 , n37957 );
and ( n37959 , n37958 , n37940 );
nor ( n37960 , n37959 , n21351 );
nand ( n37961 , n37941 , n37960 );
nand ( n37962 , n36625 , n36643 );
not ( n37963 , n37962 );
buf ( n37964 , n36615 );
not ( n37965 , n37964 );
and ( n37966 , n37965 , n37920 );
and ( n37967 , n37964 , RI15b50d60_623);
nor ( n37968 , n37966 , n37967 , n37923 );
not ( n37969 , n37968 );
nand ( n37970 , n37963 , n37969 );
not ( n37971 , n37931 );
and ( n37972 , n37971 , n36628 );
and ( n37973 , n37964 , RI15b50dd8_624);
not ( n37974 , n37934 );
nor ( n37975 , n37972 , n37973 , n37974 );
and ( n37976 , n37970 , n37975 );
not ( n37977 , n37970 );
not ( n37978 , n37975 );
and ( n37979 , n37977 , n37978 );
nor ( n37980 , n37976 , n37979 );
not ( n37981 , n33639 );
not ( n37982 , n37981 );
and ( n37983 , n37980 , n37982 );
nor ( n37984 , n21750 , n22605 );
nor ( n37985 , n37983 , n37984 );
and ( n37986 , n17562 , n18170 );
not ( n37987 , n17523 );
and ( n37988 , n21793 , n37987 , RI15b57480_843);
buf ( n37989 , n22704 );
not ( n37990 , n37989 );
or ( n37991 , n37988 , n37990 );
nand ( n37992 , n37991 , n21789 );
and ( n37993 , n37992 , RI15b57570_845);
or ( n37994 , n17558 , RI15b574f8_844);
nand ( n37995 , n37988 , n17558 , RI15b574f8_844);
nand ( n37996 , n37994 , n37995 );
buf ( n37997 , n384127 );
and ( n37998 , n37996 , n37997 );
nor ( n37999 , n37986 , n37993 , n37998 );
and ( n38000 , n379898 , n37999 );
nand ( n38001 , n37961 , n37985 , n38000 );
buf ( n38002 , n38001 );
buf ( n38003 , n33382 );
buf ( n38004 , RI15b5e410_1081);
buf ( n38005 , n383498 );
buf ( n38006 , n379847 );
not ( n38007 , n380235 );
not ( n38008 , n381507 );
or ( n38009 , n38007 , n38008 );
and ( n38010 , n381524 , n380745 );
or ( n38011 , n380776 , n18425 );
not ( n38012 , n32477 );
or ( n38013 , n38012 , n380785 );
or ( n38014 , n380768 , n381560 );
nand ( n38015 , n38011 , n38013 , n38014 );
nor ( n38016 , n38010 , n38015 );
nand ( n38017 , n38009 , n38016 );
buf ( n38018 , n38017 );
nand ( n38019 , n380002 , RI15b56418_808);
nand ( n38020 , n22592 , RI15b563a0_807);
nor ( n38021 , n379980 , n38020 );
nor ( n38022 , n22592 , RI15b563a0_807);
or ( n38023 , n38021 , n38022 );
nand ( n38024 , n38023 , n379949 );
not ( n38025 , n382744 );
not ( n38026 , n382706 );
or ( n38027 , n38025 , n38026 );
or ( n38028 , n382706 , n382744 );
nand ( n38029 , n38027 , n38028 );
nand ( n38030 , n380012 , n38029 );
nand ( n38031 , n38019 , n38024 , n38030 );
buf ( n38032 , n38031 );
buf ( n38033 , n379844 );
buf ( n38034 , n382052 );
buf ( n38035 , n22479 );
or ( n38036 , n381056 , n32812 );
or ( n38037 , n20287 , n381062 );
and ( n38038 , n32811 , RI15b49560_367);
not ( n38039 , n32811 );
and ( n38040 , n38039 , n32812 );
nor ( n38041 , n38038 , n38040 );
or ( n38042 , n38041 , n381077 );
nand ( n38043 , n38036 , n38037 , n38042 );
buf ( n38044 , n38043 );
buf ( n38045 , n381081 );
buf ( n38046 , n387159 );
buf ( n38047 , n381014 );
and ( n38048 , n38047 , RI15b53448_706);
not ( n38049 , n381014 );
and ( n38050 , n38049 , RI15b65940_1331);
nor ( n38051 , n38048 , n38050 );
not ( n38052 , n38051 );
buf ( n38053 , n38052 );
buf ( n38054 , n381566 );
buf ( n38055 , n382065 );
buf ( n38056 , n387159 );
and ( n38057 , n20634 , n20491 );
nor ( n38058 , n38057 , n20635 );
nand ( n38059 , n20638 , n20519 , n20630 , n38058 );
buf ( n38060 , n38059 );
buf ( n38061 , n22714 );
buf ( n38062 , n384203 );
buf ( n38063 , n381872 );
buf ( n38064 , n379844 );
nand ( n38065 , n32162 , n22134 );
or ( n38066 , n22102 , n38065 );
and ( n38067 , n380911 , n35933 );
and ( n38068 , n22203 , n38067 );
not ( n38069 , n38067 );
and ( n38070 , n38065 , n38069 , n19912 );
nor ( n38071 , n38070 , n22217 );
nor ( n38072 , n32175 , n380919 );
or ( n38073 , n38071 , n38072 );
nand ( n38074 , n38073 , n20623 );
or ( n38075 , n32179 , n380925 );
and ( n38076 , n38074 , n38075 );
nor ( n38077 , n38076 , n22236 );
or ( n38078 , n38077 , n20273 );
not ( n38079 , n38075 );
nor ( n38080 , n38072 , n38079 );
or ( n38081 , n38071 , n38080 );
or ( n38082 , n22293 , n38081 );
or ( n38083 , n38075 , n22299 );
nand ( n38084 , n38078 , n38082 , n38083 );
nor ( n38085 , n38068 , n38084 );
nand ( n38086 , n38066 , n38085 );
buf ( n38087 , n38086 );
buf ( n38088 , n382069 );
buf ( n38089 , RI15b5dd08_1066);
and ( n38090 , n34812 , RI15b64068_1278);
not ( n38091 , n386973 );
not ( n38092 , n38091 );
buf ( n38093 , n34814 );
not ( n38094 , n38093 );
or ( n38095 , n38092 , n38094 );
nand ( n38096 , n38095 , n34823 );
and ( n38097 , n38096 , RI15b62268_1214);
or ( n38098 , n34826 , n38091 , RI15b62268_1214);
not ( n38099 , n387032 );
not ( n38100 , n38099 );
not ( n38101 , RI15b64068_1278);
and ( n38102 , n38100 , n38101 );
and ( n38103 , n38099 , RI15b64068_1278);
nor ( n38104 , n38102 , n38103 );
or ( n38105 , n34833 , n38104 );
nand ( n38106 , n38098 , n38105 );
nor ( n38107 , n38090 , n38097 , n38106 );
or ( n38108 , n38107 , n19200 );
buf ( n38109 , n386844 );
not ( n38110 , n386839 );
not ( n38111 , n38110 );
not ( n38112 , n22473 );
and ( n38113 , n38111 , n38112 );
not ( n38114 , n383474 );
nor ( n38115 , n38113 , n38114 );
or ( n38116 , n38109 , n38115 );
not ( n38117 , n383464 );
and ( n38118 , n38117 , n38109 , n38110 );
not ( n38119 , RI15b64068_1278);
or ( n38120 , n22424 , n38119 );
or ( n38121 , n386842 , n19598 );
nand ( n38122 , n38120 , n38121 , n19512 );
nor ( n38123 , n38118 , n38122 );
nand ( n38124 , n38108 , n38116 , n38123 );
buf ( n38125 , n38124 );
buf ( n38126 , n381707 );
buf ( n38127 , n380865 );
buf ( n38128 , n386229 );
not ( n38129 , n38128 );
not ( n38130 , n386049 );
and ( n38131 , n38129 , n38130 );
and ( n38132 , n38128 , n386049 );
nor ( n38133 , n38131 , n38132 );
not ( n38134 , n386262 );
or ( n38135 , n38133 , n38134 );
not ( n38136 , n386479 );
buf ( n38137 , n386475 );
nand ( n38138 , n38137 , n386478 );
nand ( n38139 , n38136 , n38138 );
and ( n38140 , n38139 , n386500 );
nor ( n38141 , n384692 , n382130 );
nor ( n38142 , n38140 , n38141 );
nand ( n38143 , n38135 , n38142 );
not ( n38144 , n385924 );
and ( n38145 , n38144 , n385936 );
not ( n38146 , n38144 );
and ( n38147 , n38146 , n385935 );
nor ( n38148 , n38145 , n38147 );
not ( n38149 , n386018 );
nor ( n38150 , n38148 , n38149 );
nor ( n38151 , n38143 , n38150 );
not ( n38152 , n20637 );
not ( n38153 , n19884 );
or ( n38154 , n38152 , n38153 );
nand ( n38155 , n38154 , n34798 );
and ( n38156 , n38155 , RI15b4ae38_420);
or ( n38157 , n34801 , n19884 , RI15b4ae38_420);
or ( n38158 , n19890 , n22216 );
nand ( n38159 , n38157 , n38158 );
nor ( n38160 , n38156 , n38159 );
nand ( n38161 , n38151 , n38160 );
buf ( n38162 , n38161 );
buf ( n38163 , n382049 );
buf ( n38164 , n387159 );
buf ( n38165 , n381490 );
buf ( n38166 , n380865 );
not ( n38167 , n34826 );
not ( n38168 , RI15b62a60_1231);
nand ( n38169 , n38167 , n38168 );
nor ( n38170 , n387002 , n38169 );
not ( n38171 , RI15b648d8_1296);
and ( n38172 , n30852 , RI15b64860_1295);
not ( n38173 , n38172 );
or ( n38174 , n38171 , n38173 );
nand ( n38175 , n38174 , n22449 );
nor ( n38176 , n38172 , RI15b648d8_1296);
nor ( n38177 , n38175 , n38176 );
or ( n38178 , n38170 , n38177 );
nand ( n38179 , n38178 , n19201 );
not ( n38180 , n387010 );
nand ( n38181 , n38180 , n387014 );
and ( n38182 , n22426 , RI15b648d8_1296);
not ( n38183 , n22466 );
and ( n38184 , n38183 , RI15b62ad8_1232);
and ( n38185 , n19599 , RI15b639d8_1264);
nor ( n38186 , n38182 , n38184 , n38185 );
nand ( n38187 , n38179 , n38181 , n38186 );
buf ( n38188 , n38187 );
buf ( n38189 , n386563 );
not ( n38190 , n385796 );
not ( n38191 , n30867 );
or ( n38192 , n38190 , n38191 );
or ( n38193 , n30867 , n385796 );
nand ( n38194 , n38192 , n38193 );
and ( n38195 , n38194 , n386017 );
not ( n38196 , n386134 );
and ( n38197 , n386061 , n386012 );
not ( n38198 , n386061 );
not ( n38199 , n386012 );
and ( n38200 , n38198 , n38199 );
nor ( n38201 , n38197 , n38200 );
not ( n38202 , n38201 );
and ( n38203 , n38196 , n38202 );
and ( n38204 , n386134 , n38201 );
nor ( n38205 , n38203 , n38204 );
or ( n38206 , n38205 , n386260 );
xnor ( n38207 , n386362 , n386368 );
or ( n38208 , n38207 , n386499 );
not ( n38209 , n22395 );
or ( n38210 , n382099 , n38209 );
nand ( n38211 , n38206 , n38208 , n38210 );
nor ( n38212 , n38195 , n38211 );
and ( n38213 , n30908 , RI15b4a5c8_402);
or ( n38214 , n19764 , n22216 );
not ( n38215 , n19758 );
and ( n38216 , n38215 , RI15b4a5c8_402);
not ( n38217 , n38215 );
and ( n38218 , n38217 , n19762 );
nor ( n38219 , n38216 , n38218 );
or ( n38220 , n38219 , n20638 );
nand ( n38221 , n38214 , n38220 );
nor ( n38222 , n38213 , n38221 );
nand ( n38223 , n38212 , n38222 );
buf ( n38224 , n38223 );
buf ( n38225 , n19651 );
buf ( n38226 , n384218 );
buf ( n38227 , n20665 );
buf ( n38228 , n383498 );
or ( n38229 , n381907 , n36082 );
not ( n38230 , n36094 );
and ( n38231 , n38230 , RI15b41298_88);
or ( n38232 , n381917 , n36086 );
not ( n38233 , n36098 );
and ( n38234 , n38233 , n381923 );
and ( n38235 , n381926 , n36096 );
nor ( n38236 , n38234 , n38235 );
nand ( n38237 , n38232 , n38236 );
nor ( n38238 , n38231 , n38237 );
nand ( n38239 , n38229 , n38238 );
buf ( n38240 , n38239 );
and ( n38241 , n22148 , n35903 );
not ( n38242 , n35903 );
and ( n38243 , n22147 , n38242 );
nor ( n38244 , n38241 , n38243 );
or ( n38245 , n38244 , n20638 );
or ( n38246 , n36110 , RI15b3fc18_40);
not ( n38247 , n22235 );
nand ( n38248 , n38246 , n38247 );
and ( n38249 , n38248 , RI15b3fd80_43);
not ( n38250 , n22207 );
and ( n38251 , n22217 , n38250 );
and ( n38252 , n381925 , n22115 );
nor ( n38253 , n38249 , n38251 , n38252 );
nand ( n38254 , n38245 , n38253 );
buf ( n38255 , n38254 );
buf ( n38256 , n30992 );
buf ( n38257 , n382065 );
buf ( n38258 , n379802 );
or ( n38259 , n37478 , n36082 );
and ( n38260 , n384983 , n36084 );
not ( n38261 , RI15b41478_92);
or ( n38262 , n36094 , n38261 );
or ( n38263 , n22022 , n36098 );
or ( n38264 , n36092 , n384988 );
nand ( n38265 , n38262 , n38263 , n38264 );
nor ( n38266 , n38260 , n38265 );
nand ( n38267 , n38259 , n38266 );
buf ( n38268 , n38267 );
buf ( n38269 , n385195 );
buf ( n38270 , n31979 );
buf ( n38271 , RI15b45ff0_253);
buf ( n38272 , n379844 );
buf ( n38273 , n22007 );
buf ( n38274 , n32160 );
buf ( n38275 , n383345 );
or ( n38276 , n22315 , n37495 );
and ( n38277 , n22326 , n37498 );
not ( n38278 , RI15b425d0_129);
or ( n38279 , n37507 , n38278 );
or ( n38280 , n22334 , n37512 );
or ( n38281 , n37505 , n22336 );
nand ( n38282 , n38279 , n38280 , n38281 );
nor ( n38283 , n38277 , n38282 );
nand ( n38284 , n38276 , n38283 );
buf ( n38285 , n38284 );
not ( n38286 , n383318 );
nor ( n38287 , n38286 , n383152 );
not ( n38288 , n383157 );
or ( n38289 , n38287 , n38288 );
buf ( n38290 , n383306 );
not ( n38291 , n38290 );
nand ( n38292 , n38289 , n38291 );
nand ( n38293 , n38290 , n38286 , n383143 );
and ( n38294 , n383170 , RI15b54000_731);
and ( n38295 , n383147 , RI15b529f8_684);
nor ( n38296 , n38294 , n38295 );
nand ( n38297 , n38292 , n38293 , n38296 );
buf ( n38298 , n38297 );
buf ( n38299 , n22007 );
buf ( n38300 , n379802 );
buf ( n38301 , n382069 );
not ( n38302 , n382976 );
not ( n38303 , n382912 );
or ( n38304 , n38302 , n38303 );
and ( n38305 , n382931 , n382983 );
or ( n38306 , n382995 , n19072 );
not ( n38307 , n382958 );
or ( n38308 , n38307 , n383001 );
or ( n38309 , n382993 , n382967 );
nand ( n38310 , n38306 , n38308 , n38309 );
nor ( n38311 , n38305 , n38310 );
nand ( n38312 , n38304 , n38311 );
buf ( n38313 , n38312 );
buf ( n38314 , n18226 );
buf ( n38315 , n22479 );
not ( n38316 , RI15b55c98_792);
not ( n38317 , n380000 );
or ( n38318 , n38316 , n38317 );
and ( n38319 , n381636 , RI15b4e9c0_547);
and ( n38320 , n381639 , RI15b4e600_539);
nor ( n38321 , n38319 , n38320 );
and ( n38322 , n381643 , RI15b4ed80_555);
buf ( n38323 , n380007 );
and ( n38324 , n381651 , RI15b4dac0_515);
and ( n38325 , n381657 , RI15b4fc80_587);
nor ( n38326 , n38324 , n38325 );
and ( n38327 , n381661 , RI15b4f8c0_579);
and ( n38328 , n381663 , RI15b4f140_563);
nor ( n38329 , n38327 , n38328 );
and ( n38330 , n381667 , RI15b4d340_499);
and ( n38331 , n381669 , RI15b4d700_507);
nor ( n38332 , n38330 , n38331 );
and ( n38333 , n381672 , RI15b4de80_523);
and ( n38334 , n381674 , RI15b4f500_571);
nor ( n38335 , n38333 , n38334 );
nand ( n38336 , n38326 , n38329 , n38332 , n38335 );
and ( n38337 , n38323 , n38336 );
and ( n38338 , n381680 , RI15b4c800_475);
nor ( n38339 , n38322 , n38337 , n38338 );
and ( n38340 , n381684 , RI15b4c440_467);
and ( n38341 , n381686 , RI15b4e240_531);
nor ( n38342 , n38340 , n38341 );
and ( n38343 , n381689 , RI15b4cbc0_483);
and ( n38344 , n381691 , RI15b4cf80_491);
nor ( n38345 , n38343 , n38344 );
nand ( n38346 , n38321 , n38339 , n38342 , n38345 );
not ( n38347 , n381695 );
and ( n38348 , n38346 , n38347 );
not ( n38349 , RI15b55c98_792);
not ( n38350 , n379961 );
not ( n38351 , n38350 );
or ( n38352 , n38349 , n38351 );
or ( n38353 , n38350 , RI15b55c98_792);
nand ( n38354 , n38352 , n38353 );
and ( n38355 , n379949 , n38354 );
nor ( n38356 , n38348 , n38355 );
nand ( n38357 , n38318 , n38356 );
buf ( n38358 , n38357 );
not ( n38359 , n381570 );
not ( n38360 , n381507 );
or ( n38361 , n38359 , n38360 );
and ( n38362 , n381524 , n381599 );
or ( n38363 , n381609 , n18420 );
or ( n38364 , n32478 , n381619 );
or ( n38365 , n381607 , n381560 );
nand ( n38366 , n38363 , n38364 , n38365 );
nor ( n38367 , n38362 , n38366 );
nand ( n38368 , n38361 , n38367 );
buf ( n38369 , n38368 );
buf ( n38370 , n22343 );
buf ( n38371 , n22005 );
buf ( n38372 , n17499 );
nand ( n38373 , n32162 , n35876 );
or ( n38374 , n22315 , n38373 );
and ( n38375 , n32168 , n32163 );
and ( n38376 , n22326 , n38375 );
not ( n38377 , n38375 );
and ( n38378 , n38373 , n38377 , n19912 );
nor ( n38379 , n38378 , n22217 );
nor ( n38380 , n32175 , n36818 );
or ( n38381 , n38379 , n38380 );
nand ( n38382 , n38381 , n20623 );
or ( n38383 , n32179 , n22133 );
and ( n38384 , n38382 , n38383 );
nor ( n38385 , n38384 , n22236 );
or ( n38386 , n38385 , n20169 );
not ( n38387 , n38383 );
nor ( n38388 , n38380 , n38387 );
or ( n38389 , n38379 , n38388 );
or ( n38390 , n22334 , n38389 );
or ( n38391 , n38383 , n22336 );
nand ( n38392 , n38386 , n38390 , n38391 );
nor ( n38393 , n38376 , n38392 );
nand ( n38394 , n38374 , n38393 );
buf ( n38395 , n38394 );
buf ( n38396 , n383613 );
buf ( n38397 , n20663 );
or ( n38398 , n36937 , n35622 );
and ( n38399 , n36946 , n35625 );
not ( n38400 , RI15b4f668_574);
or ( n38401 , n35635 , n38400 );
buf ( n38402 , n36950 );
not ( n38403 , n38402 );
or ( n38404 , n38403 , n35640 );
or ( n38405 , n35633 , n36955 );
nand ( n38406 , n38401 , n38404 , n38405 );
nor ( n38407 , n38399 , n38406 );
nand ( n38408 , n38398 , n38407 );
buf ( n38409 , n38408 );
not ( n38410 , RI15b5f838_1124);
not ( n38411 , n383601 );
or ( n38412 , n38410 , n38411 );
and ( n38413 , n383505 , RI15b60dc8_1170);
and ( n38414 , n383607 , RI15b5f0b8_1108);
nor ( n38415 , n38413 , n38414 );
nand ( n38416 , n38412 , n38415 );
buf ( n38417 , n38416 );
buf ( n38418 , n22740 );
buf ( n38419 , n22007 );
buf ( n38420 , n22655 );
buf ( n38421 , n22653 );
buf ( n38422 , n382052 );
buf ( n38423 , n32255 );
not ( n38424 , RI15b53880_715);
not ( n38425 , n32244 );
or ( n38426 , n38424 , n38425 );
and ( n38427 , n32247 , RI15b64e78_1308);
and ( n38428 , n32249 , RI15b5fce8_1134);
nor ( n38429 , n38427 , n38428 );
nand ( n38430 , n38426 , n38429 );
buf ( n38431 , n38430 );
buf ( n38432 , n19655 );
not ( n38433 , n37131 );
not ( n38434 , RI15b4a028_390);
and ( n38435 , n38433 , n38434 );
not ( n38436 , n38433 );
and ( n38437 , n38436 , RI15b4a028_390);
nor ( n38438 , n38435 , n38437 );
nand ( n38439 , n38438 , n37114 );
and ( n38440 , n381055 , RI15b4a028_390);
not ( n38441 , n37320 );
not ( n38442 , n37288 );
or ( n38443 , n38441 , n38442 );
or ( n38444 , n37288 , n37320 );
nand ( n38445 , n38443 , n38444 );
and ( n38446 , n386555 , n38445 );
nor ( n38447 , n38440 , n38446 );
nand ( n38448 , n38439 , n38447 );
buf ( n38449 , n38448 );
buf ( n38450 , n22404 );
buf ( n38451 , n22738 );
buf ( n38452 , n30992 );
buf ( n38453 , n31033 );
not ( n38454 , RI15b658c8_1330);
not ( n38455 , n35176 );
or ( n38456 , n38454 , n38455 );
nand ( n38457 , n35187 , RI15b484f8_332);
buf ( n38458 , n385696 );
and ( n38459 , n386554 , n38458 );
not ( n38460 , RI15b48480_331);
or ( n38461 , n38460 , RI15b484f8_332);
not ( n38462 , RI15b484f8_332);
or ( n38463 , n38462 , RI15b48480_331);
nand ( n38464 , n38461 , n38463 );
and ( n38465 , n35363 , n38464 );
nor ( n38466 , n38459 , n38465 );
and ( n38467 , n379841 , n38457 , n38466 );
nand ( n38468 , n38456 , n38467 );
buf ( n38469 , n38468 );
not ( n38470 , n384025 );
and ( n38471 , n384039 , RI15b62100_1211);
nor ( n38472 , n386970 , n386972 );
nand ( n38473 , n38471 , n38472 );
not ( n38474 , RI15b62268_1214);
nor ( n38475 , n38473 , n38474 );
and ( n38476 , n38475 , RI15b622e0_1215);
and ( n38477 , n38476 , RI15b62358_1216);
nand ( n38478 , n38477 , RI15b623d0_1217);
nor ( n38479 , n38478 , n386980 );
and ( n38480 , n38479 , RI15b624c0_1219);
nand ( n38481 , n38480 , RI15b62538_1220 , RI15b625b0_1221);
not ( n38482 , RI15b62628_1222);
nor ( n38483 , n38481 , n38482 );
nand ( n38484 , n38483 , RI15b626a0_1223);
nor ( n38485 , n38484 , n386990 );
and ( n38486 , n38485 , RI15b62790_1225);
nand ( n38487 , n38486 , RI15b62808_1226);
nor ( n38488 , n38487 , n386995 );
nand ( n38489 , n38488 , RI15b628f8_1228);
not ( n38490 , n38489 );
or ( n38491 , n38470 , n38490 );
nand ( n38492 , n38491 , n384021 );
nor ( n38493 , n384024 , RI15b62970_1229);
nor ( n38494 , n38492 , n38493 );
or ( n38495 , n38494 , n387001 );
not ( n38496 , n38489 );
not ( n38497 , n38496 );
nand ( n38498 , n384025 , RI15b62970_1229);
nor ( n38499 , n38497 , n38498 );
nand ( n38500 , n38499 , n387001 );
buf ( n38501 , n18812 );
and ( n38502 , n19266 , n38501 );
and ( n38503 , n38502 , RI15b59c58_928);
not ( n38504 , n383938 );
not ( n38505 , n38504 );
and ( n38506 , n18789 , n38505 );
and ( n38507 , n38506 , RI15b5be18_1000);
nor ( n38508 , n38503 , n38507 );
and ( n38509 , n18789 , n38501 );
and ( n38510 , n38509 , RI15b5a018_936);
not ( n38511 , n38504 );
and ( n38512 , n19266 , n38511 );
and ( n38513 , n38512 , RI15b5ba58_992);
nor ( n38514 , n38510 , n38513 );
and ( n38515 , n19274 , n38501 );
and ( n38516 , n38515 , RI15b5a3d8_944);
not ( n38517 , n18794 );
and ( n38518 , n38517 , RI15b5ab58_960);
nor ( n38519 , n38516 , n38518 );
buf ( n38520 , n18835 );
buf ( n38521 , n38520 );
buf ( n38522 , n38521 );
buf ( n38523 , n38522 );
and ( n38524 , n38523 , RI15b5b2d8_976);
and ( n38525 , n19274 , n38511 );
and ( n38526 , n38525 , RI15b5c1d8_1008);
nor ( n38527 , n38524 , n38526 );
nand ( n38528 , n38508 , n38514 , n38519 , n38527 );
and ( n38529 , n19256 , n38505 );
and ( n38530 , n38529 , RI15b5b698_984);
not ( n38531 , n18843 );
and ( n38532 , n38531 , RI15b5af18_968);
nor ( n38533 , n38530 , n38532 );
and ( n38534 , n19256 , n38501 );
and ( n38535 , n38534 , RI15b59898_920);
not ( n38536 , n18849 );
and ( n38537 , n38536 , RI15b5a798_952);
nor ( n38538 , n38535 , n38537 );
not ( n38539 , n18864 );
and ( n38540 , n38539 , RI15b58998_888);
not ( n38541 , n18859 );
and ( n38542 , n38541 , RI15b594d8_912);
nor ( n38543 , n38540 , n38542 );
not ( n38544 , n18807 );
and ( n38545 , n38544 , RI15b58d58_896);
buf ( n38546 , n18799 );
buf ( n38547 , n38546 );
buf ( n38548 , n38547 );
buf ( n38549 , n38548 );
and ( n38550 , n38549 , RI15b59118_904);
nor ( n38551 , n38545 , n38550 );
nand ( n38552 , n38533 , n38538 , n38543 , n38551 );
nor ( n38553 , n38528 , n38552 );
not ( n38554 , n38553 );
and ( n38555 , n38502 , RI15b59a78_924);
and ( n38556 , n38506 , RI15b5bc38_996);
nor ( n38557 , n38555 , n38556 );
and ( n38558 , n38509 , RI15b59e38_932);
and ( n38559 , n38512 , RI15b5b878_988);
nor ( n38560 , n38558 , n38559 );
and ( n38561 , n38515 , RI15b5a1f8_940);
and ( n38562 , n38517 , RI15b5a978_956);
nor ( n38563 , n38561 , n38562 );
and ( n38564 , n38520 , RI15b5b0f8_972);
and ( n38565 , n38525 , RI15b5bff8_1004);
nor ( n38566 , n38564 , n38565 );
nand ( n38567 , n38557 , n38560 , n38563 , n38566 );
and ( n38568 , n38529 , RI15b5b4b8_980);
and ( n38569 , n38531 , RI15b5ad38_964);
nor ( n38570 , n38568 , n38569 );
and ( n38571 , n38534 , RI15b596b8_916);
and ( n38572 , n38536 , RI15b5a5b8_948);
nor ( n38573 , n38571 , n38572 );
and ( n38574 , n38539 , RI15b587b8_884);
and ( n38575 , n38541 , RI15b592f8_908);
nor ( n38576 , n38574 , n38575 );
and ( n38577 , n38544 , RI15b58b78_892);
and ( n38578 , n38546 , RI15b58f38_900);
nor ( n38579 , n38577 , n38578 );
nand ( n38580 , n38570 , n38573 , n38576 , n38579 );
nor ( n38581 , n38567 , n38580 );
not ( n38582 , n38581 );
buf ( n38583 , n18775 );
not ( n38584 , n38583 );
not ( n38585 , n18258 );
and ( n38586 , n38584 , n38585 );
not ( n38587 , RI15b5d420_1047);
not ( n38588 , n18775 );
or ( n38589 , n38587 , n38588 );
not ( n38590 , n383937 );
nand ( n38591 , n38589 , n38590 );
nor ( n38592 , n38586 , n38591 );
not ( n38593 , n38583 );
not ( n38594 , RI15b5d3a8_1046);
and ( n38595 , n38593 , n38594 );
and ( n38596 , n18927 , RI15b5d3a8_1046);
nor ( n38597 , n38595 , n38596 );
not ( n38598 , n38597 );
nand ( n38599 , n38592 , n38598 );
buf ( n38600 , n18290 );
not ( n38601 , n38600 );
not ( n38602 , n38601 );
nor ( n38603 , n38599 , n38602 );
and ( n38604 , n38603 , RI15b5a540_947);
buf ( n38605 , n18618 );
not ( n38606 , n38605 );
nor ( n38607 , n38599 , n38606 );
and ( n38608 , n38607 , RI15b5a180_939);
buf ( n38609 , n18375 );
not ( n38610 , n38609 );
not ( n38611 , n19031 );
and ( n38612 , n38610 , n38611 );
not ( n38613 , RI15b59280_907);
not ( n38614 , n18618 );
or ( n38615 , n38613 , n38614 );
buf ( n38616 , n18250 );
nand ( n38617 , n38616 , RI15b58ec0_899);
nand ( n38618 , n38615 , n38617 );
nor ( n38619 , n38612 , n38618 );
nand ( n38620 , n38592 , n38597 );
or ( n38621 , n38619 , n38620 );
nor ( n38622 , n38592 , n38597 );
nand ( n38623 , n38622 , n38601 , RI15b5c340_1011);
nand ( n38624 , n38621 , n38623 );
nor ( n38625 , n38604 , n38608 , n38624 );
buf ( n38626 , n38616 );
not ( n38627 , n38626 );
nor ( n38628 , n38599 , n38627 );
and ( n38629 , n38628 , RI15b59dc0_931);
buf ( n38630 , n38609 );
nor ( n38631 , n38599 , n38630 );
and ( n38632 , n38631 , RI15b59a00_923);
not ( n38633 , RI15b5b800_987);
not ( n38634 , n18376 );
or ( n38635 , n38633 , n38634 );
not ( n38636 , n37539 );
nand ( n38637 , n38636 , n18618 );
nand ( n38638 , n38635 , n38637 );
and ( n38639 , n38616 , RI15b5bbc0_995);
nor ( n38640 , n38638 , n38639 );
not ( n38641 , n38622 );
or ( n38642 , n38640 , n38641 );
not ( n38643 , n38600 );
nand ( n38644 , n38643 , RI15b59640_915);
or ( n38645 , n38620 , n38644 );
nand ( n38646 , n38642 , n38645 );
nor ( n38647 , n38629 , n38632 , n38646 );
not ( n38648 , n38592 );
nand ( n38649 , n38648 , n38597 );
not ( n38650 , n38649 );
buf ( n38651 , n38600 );
not ( n38652 , n38651 );
nand ( n38653 , n38650 , n38652 );
not ( n38654 , n38653 );
and ( n38655 , n38654 , RI15b5b440_979);
not ( n38656 , n38605 );
nor ( n38657 , n38649 , n38656 );
and ( n38658 , n38657 , RI15b5b080_971);
nor ( n38659 , n38655 , n38658 );
and ( n38660 , n38650 , n38626 );
and ( n38661 , n38660 , RI15b5acc0_963);
nor ( n38662 , n38649 , n38630 );
and ( n38663 , n38662 , RI15b5a900_955);
nor ( n38664 , n38661 , n38663 );
nand ( n38665 , n38625 , n38647 , n38659 , n38664 );
nand ( n38666 , n38582 , n38665 );
and ( n38667 , n38502 , RI15b59af0_925);
and ( n38668 , n38506 , RI15b5bcb0_997);
nor ( n38669 , n38667 , n38668 );
and ( n38670 , n38509 , RI15b59eb0_933);
and ( n38671 , n38512 , RI15b5b8f0_989);
nor ( n38672 , n38670 , n38671 );
and ( n38673 , n38515 , RI15b5a270_941);
and ( n38674 , n38517 , RI15b5a9f0_957);
nor ( n38675 , n38673 , n38674 );
and ( n38676 , n38521 , RI15b5b170_973);
and ( n38677 , n38525 , RI15b5c070_1005);
nor ( n38678 , n38676 , n38677 );
nand ( n38679 , n38669 , n38672 , n38675 , n38678 );
and ( n38680 , n38529 , RI15b5b530_981);
and ( n38681 , n38531 , RI15b5adb0_965);
nor ( n38682 , n38680 , n38681 );
and ( n38683 , n38534 , RI15b59730_917);
and ( n38684 , n38536 , RI15b5a630_949);
nor ( n38685 , n38683 , n38684 );
and ( n38686 , n38539 , RI15b58830_885);
and ( n38687 , n38541 , RI15b59370_909);
nor ( n38688 , n38686 , n38687 );
and ( n38689 , n38544 , RI15b58bf0_893);
and ( n38690 , n38547 , RI15b58fb0_901);
nor ( n38691 , n38689 , n38690 );
nand ( n38692 , n38682 , n38685 , n38688 , n38691 );
nor ( n38693 , n38679 , n38692 );
nor ( n38694 , n38666 , n38693 );
and ( n38695 , n38502 , RI15b59b68_926);
and ( n38696 , n38506 , RI15b5bd28_998);
nor ( n38697 , n38695 , n38696 );
and ( n38698 , n38509 , RI15b59f28_934);
and ( n38699 , n38512 , RI15b5b968_990);
nor ( n38700 , n38698 , n38699 );
and ( n38701 , n38515 , RI15b5a2e8_942);
and ( n38702 , n38517 , RI15b5aa68_958);
nor ( n38703 , n38701 , n38702 );
and ( n38704 , n38521 , RI15b5b1e8_974);
and ( n38705 , n38525 , RI15b5c0e8_1006);
nor ( n38706 , n38704 , n38705 );
nand ( n38707 , n38697 , n38700 , n38703 , n38706 );
and ( n38708 , n38529 , RI15b5b5a8_982);
and ( n38709 , n38531 , RI15b5ae28_966);
nor ( n38710 , n38708 , n38709 );
and ( n38711 , n38534 , RI15b597a8_918);
and ( n38712 , n38536 , RI15b5a6a8_950);
nor ( n38713 , n38711 , n38712 );
and ( n38714 , n38539 , RI15b588a8_886);
and ( n38715 , n38541 , RI15b593e8_910);
nor ( n38716 , n38714 , n38715 );
and ( n38717 , n38544 , RI15b58c68_894);
and ( n38718 , n38547 , RI15b59028_902);
nor ( n38719 , n38717 , n38718 );
nand ( n38720 , n38710 , n38713 , n38716 , n38719 );
nor ( n38721 , n38707 , n38720 );
not ( n38722 , n38721 );
and ( n38723 , n38694 , n38722 );
and ( n38724 , n38502 , RI15b59be0_927);
and ( n38725 , n38506 , RI15b5bda0_999);
nor ( n38726 , n38724 , n38725 );
and ( n38727 , n38509 , RI15b59fa0_935);
and ( n38728 , n38512 , RI15b5b9e0_991);
nor ( n38729 , n38727 , n38728 );
and ( n38730 , n38515 , RI15b5a360_943);
and ( n38731 , n38517 , RI15b5aae0_959);
nor ( n38732 , n38730 , n38731 );
and ( n38733 , n38522 , RI15b5b260_975);
and ( n38734 , n38525 , RI15b5c160_1007);
nor ( n38735 , n38733 , n38734 );
nand ( n38736 , n38726 , n38729 , n38732 , n38735 );
and ( n38737 , n38529 , RI15b5b620_983);
and ( n38738 , n38531 , RI15b5aea0_967);
nor ( n38739 , n38737 , n38738 );
and ( n38740 , n38534 , RI15b59820_919);
and ( n38741 , n38536 , RI15b5a720_951);
nor ( n38742 , n38740 , n38741 );
and ( n38743 , n38539 , RI15b58920_887);
and ( n38744 , n38541 , RI15b59460_911);
nor ( n38745 , n38743 , n38744 );
and ( n38746 , n38544 , RI15b58ce0_895);
and ( n38747 , n38548 , RI15b590a0_903);
nor ( n38748 , n38746 , n38747 );
nand ( n38749 , n38739 , n38742 , n38745 , n38748 );
nor ( n38750 , n38736 , n38749 );
not ( n38751 , n38750 );
and ( n38752 , n38723 , n38751 );
nand ( n38753 , n38554 , n38752 );
and ( n38754 , n38502 , RI15b59cd0_929);
and ( n38755 , n38506 , RI15b5be90_1001);
nor ( n38756 , n38754 , n38755 );
and ( n38757 , n38509 , RI15b5a090_937);
and ( n38758 , n38512 , RI15b5bad0_993);
nor ( n38759 , n38757 , n38758 );
and ( n38760 , n38515 , RI15b5a450_945);
and ( n38761 , n38517 , RI15b5abd0_961);
nor ( n38762 , n38760 , n38761 );
buf ( n38763 , n38523 );
and ( n38764 , n38763 , RI15b5b350_977);
and ( n38765 , n38525 , RI15b5c250_1009);
nor ( n38766 , n38764 , n38765 );
nand ( n38767 , n38756 , n38759 , n38762 , n38766 );
and ( n38768 , n38529 , RI15b5b710_985);
and ( n38769 , n38531 , RI15b5af90_969);
nor ( n38770 , n38768 , n38769 );
and ( n38771 , n38534 , RI15b59910_921);
and ( n38772 , n38536 , RI15b5a810_953);
nor ( n38773 , n38771 , n38772 );
and ( n38774 , n38539 , RI15b58a10_889);
and ( n38775 , n38541 , RI15b59550_913);
nor ( n38776 , n38774 , n38775 );
and ( n38777 , n38544 , RI15b58dd0_897);
buf ( n38778 , n38549 );
and ( n38779 , n38778 , RI15b59190_905);
nor ( n38780 , n38777 , n38779 );
nand ( n38781 , n38770 , n38773 , n38776 , n38780 );
nor ( n38782 , n38767 , n38781 );
nor ( n38783 , n38753 , n38782 );
not ( n38784 , n38783 );
and ( n38785 , n38502 , RI15b59d48_930);
and ( n38786 , n38509 , RI15b5a108_938);
nor ( n38787 , n38785 , n38786 );
and ( n38788 , n38512 , RI15b5bb48_994);
and ( n38789 , n38506 , RI15b5bf08_1002);
nor ( n38790 , n38788 , n38789 );
and ( n38791 , n38515 , RI15b5a4c8_946);
and ( n38792 , n38517 , RI15b5ac48_962);
nor ( n38793 , n38791 , n38792 );
buf ( n38794 , n38763 );
and ( n38795 , n38794 , RI15b5b3c8_978);
and ( n38796 , n38525 , RI15b5c2c8_1010);
nor ( n38797 , n38795 , n38796 );
nand ( n38798 , n38787 , n38790 , n38793 , n38797 );
and ( n38799 , n38529 , RI15b5b788_986);
and ( n38800 , n38531 , RI15b5b008_970);
nor ( n38801 , n38799 , n38800 );
and ( n38802 , n38534 , RI15b59988_922);
and ( n38803 , n38539 , RI15b58a88_890);
nor ( n38804 , n38802 , n38803 );
and ( n38805 , n38536 , RI15b5a888_954);
and ( n38806 , n38541 , RI15b595c8_914);
nor ( n38807 , n38805 , n38806 );
and ( n38808 , n38544 , RI15b58e48_898);
buf ( n38809 , n38778 );
and ( n38810 , n38809 , RI15b59208_906);
nor ( n38811 , n38808 , n38810 );
nand ( n38812 , n38801 , n38804 , n38807 , n38811 );
nor ( n38813 , n38798 , n38812 );
not ( n38814 , n38813 );
and ( n38815 , n38784 , n38814 );
and ( n38816 , n38783 , n38813 );
nor ( n38817 , n38815 , n38816 );
or ( n38818 , n38817 , n386747 );
nand ( n38819 , n38495 , n38500 , n38818 );
buf ( n38820 , n38819 );
buf ( n38821 , n381021 );
buf ( n38822 , n382069 );
buf ( n38823 , n385000 );
not ( n38824 , n385001 );
nand ( n38825 , n38823 , n38824 );
or ( n38826 , n31006 , n38825 );
nand ( n38827 , n384167 , n383866 );
not ( n38828 , n38827 );
and ( n38829 , n31016 , n38828 );
and ( n38830 , n38827 , n38825 , n33119 );
nor ( n38831 , n38830 , n21764 );
nor ( n38832 , n384173 , n383888 );
or ( n38833 , n38831 , n38832 );
nand ( n38834 , n38833 , n18154 );
or ( n38835 , n384179 , n383894 );
nand ( n38836 , n38834 , n38835 );
and ( n38837 , n38836 , n383901 );
or ( n38838 , n38837 , n17723 );
not ( n38839 , n38835 );
nor ( n38840 , n38832 , n38839 );
or ( n38841 , n38831 , n38840 );
or ( n38842 , n31022 , n38841 );
or ( n38843 , n38835 , n31024 );
nand ( n38844 , n38838 , n38842 , n38843 );
nor ( n38845 , n38829 , n38844 );
nand ( n38846 , n38826 , n38845 );
buf ( n38847 , n38846 );
buf ( n38848 , n22009 );
buf ( n38849 , n384199 );
buf ( n38850 , n383498 );
buf ( n38851 , n22404 );
buf ( n38852 , n17499 );
buf ( n38853 , n382073 );
not ( n38854 , n382030 );
not ( n38855 , n382017 );
or ( n38856 , n38854 , n38855 );
or ( n38857 , n382017 , n382030 );
nand ( n38858 , n38856 , n38857 );
and ( n38859 , n379822 , n38858 );
nor ( n38860 , n379834 , n382025 );
nor ( n38861 , n38859 , n38860 );
nand ( n38862 , n379832 , RI15b46d10_281);
nand ( n38863 , n379825 , RI15b48a20_343);
nand ( n38864 , n38861 , n38862 , n38863 );
buf ( n38865 , n38864 );
buf ( n38866 , n22005 );
buf ( n38867 , n385197 );
or ( n38868 , n381907 , n32165 );
not ( n38869 , n32183 );
and ( n38870 , n38869 , RI15b43458_160);
or ( n38871 , n381917 , n32172 );
not ( n38872 , n32187 );
and ( n38873 , n38872 , n381923 );
and ( n38874 , n381926 , n32185 );
nor ( n38875 , n38873 , n38874 );
nand ( n38876 , n38871 , n38875 );
nor ( n38877 , n38870 , n38876 );
nand ( n38878 , n38868 , n38877 );
buf ( n38879 , n38878 );
buf ( n38880 , n22406 );
buf ( n38881 , n381021 );
and ( n38882 , n31770 , RI15b5c610_1017);
or ( n38883 , n31782 , n19313 );
and ( n38884 , n32386 , n18688 );
and ( n38885 , n31778 , n19450 );
nor ( n38886 , n38884 , n38885 );
nand ( n38887 , n38883 , n38886 );
nor ( n38888 , n38882 , n33072 , n38887 );
not ( n38889 , n38888 );
buf ( n38890 , n38889 );
buf ( n38891 , n21800 );
buf ( n38892 , n383087 );
not ( n38893 , n38892 );
buf ( n38894 , n383140 );
nor ( n38895 , n38893 , n38894 );
nand ( n38896 , n38895 , n381461 );
not ( n38897 , n381423 );
not ( n38898 , n38897 );
not ( n38899 , n38894 );
or ( n38900 , n38898 , n38899 );
nand ( n38901 , n38900 , n381450 );
not ( n38902 , n38892 );
nand ( n38903 , n38901 , n38902 );
nand ( n38904 , n381485 , RI15b52890_681);
nor ( n38905 , n381400 , n381408 );
not ( n38906 , n38905 );
nand ( n38907 , n38896 , n38903 , n38904 , n38906 );
buf ( n38908 , n38907 );
buf ( n38909 , n379893 );
buf ( n38910 , n32538 );
or ( n38911 , n32537 , n38910 );
not ( n38912 , n32539 );
nand ( n38913 , n38911 , n38912 );
and ( n38914 , n38913 , n384391 );
nor ( n38915 , n35267 , n35265 );
not ( n38916 , n38915 );
not ( n38917 , n384433 );
and ( n38918 , n38916 , n38917 );
and ( n38919 , n38915 , n384433 );
nor ( n38920 , n38918 , n38919 );
not ( n38921 , n384492 );
or ( n38922 , n38920 , n38921 );
xor ( n38923 , n384526 , n384558 );
and ( n38924 , n38923 , n19286 );
and ( n38925 , n19513 , RI15b63ff0_1277);
nor ( n38926 , n38924 , n38925 );
nand ( n38927 , n38922 , n38926 );
nor ( n38928 , n38914 , n38927 );
and ( n38929 , n384634 , RI15b630f0_1245);
and ( n38930 , n386838 , n19630 );
and ( n38931 , n384631 , n384636 );
nor ( n38932 , n38929 , n38930 , n38931 );
nand ( n38933 , n38928 , n38932 );
buf ( n38934 , n38933 );
buf ( n38935 , n22402 );
buf ( n38936 , n22716 );
buf ( n38937 , n19891 );
not ( n38938 , n19920 );
nor ( n38939 , n38937 , n38938 );
not ( n38940 , n22350 );
or ( n38941 , n38939 , n38940 );
nand ( n38942 , n38941 , n19897 );
buf ( n38943 , n19994 );
not ( n38944 , n38943 );
nor ( n38945 , n38944 , n20502 );
or ( n38946 , n38945 , n20521 );
nand ( n38947 , n38946 , RI15b49fb0_389);
nand ( n38948 , n32511 , n19995 );
nor ( n38949 , n38943 , n38948 );
nor ( n38950 , n35312 , n382135 );
or ( n38951 , n22354 , n35310 , RI15b4bdb0_453);
or ( n38952 , n22390 , n19696 );
nand ( n38953 , n38951 , n38952 );
nor ( n38954 , n38949 , n38950 , n38953 );
nor ( n38955 , n20525 , n19897 );
nand ( n38956 , n38937 , n38955 );
nand ( n38957 , n38942 , n38947 , n38954 , n38956 );
buf ( n38958 , n38957 );
buf ( n38959 , n32676 );
buf ( n38960 , n380906 );
buf ( n38961 , n22788 );
buf ( n38962 , n383613 );
or ( n38963 , n31149 , n383845 );
and ( n38964 , n31161 , n383878 );
not ( n38965 , RI15b4f140_563);
or ( n38966 , n383903 , n38965 );
or ( n38967 , n32452 , n383911 );
or ( n38968 , n383895 , n31184 );
nand ( n38969 , n38966 , n38967 , n38968 );
nor ( n38970 , n38964 , n38969 );
nand ( n38971 , n38963 , n38970 );
buf ( n38972 , n38971 );
buf ( n38973 , n32981 );
not ( n38974 , n383504 );
not ( n38975 , n38974 );
not ( n38976 , n383566 );
and ( n38977 , n38975 , n38976 );
nor ( n38978 , n38977 , n383577 );
not ( n38979 , n383574 );
or ( n38980 , n38978 , n38979 );
and ( n38981 , n383601 , RI15b5fd60_1135);
and ( n38982 , n383566 , n38979 );
and ( n38983 , n383603 , n38982 );
and ( n38984 , n383607 , RI15b5f5e0_1119);
nor ( n38985 , n38981 , n38983 , n38984 );
nand ( n38986 , n38980 , n38985 );
buf ( n38987 , n38986 );
not ( n38988 , n19918 );
not ( n38989 , n38988 );
buf ( n38990 , n19781 );
not ( n38991 , n38990 );
or ( n38992 , n38989 , n38991 );
nand ( n38993 , n38992 , n22350 );
not ( n38994 , n19788 );
and ( n38995 , n38993 , n38994 );
buf ( n38996 , n380882 );
buf ( n38997 , n20540 );
or ( n38998 , n38996 , n38997 , RI15b4b630_437);
not ( n38999 , n19968 );
or ( n39000 , n22362 , n38999 , RI15b49830_373);
nand ( n39001 , n38998 , n39000 );
nor ( n39002 , n38995 , n39001 );
not ( n39003 , n38994 );
not ( n39004 , n38990 );
nand ( n39005 , n39003 , n383353 , n39004 );
and ( n39006 , n20565 , n38997 );
nor ( n39007 , n39006 , n22372 );
not ( n39008 , RI15b4b630_437);
or ( n39009 , n39007 , n39008 );
and ( n39010 , n22378 , n38999 );
nor ( n39011 , n39010 , n22383 );
or ( n39012 , n39011 , n32821 );
nand ( n39013 , n39009 , n39012 );
nand ( n39014 , n39013 , n20501 );
and ( n39015 , n22388 , RI15b4b630_437);
and ( n39016 , n32621 , RI15b4a730_405);
nor ( n39017 , n39015 , n39016 , n383396 );
nand ( n39018 , n39002 , n39005 , n39014 , n39017 );
buf ( n39019 , n39018 );
buf ( n39020 , n19651 );
buf ( n39021 , n22479 );
buf ( n39022 , n380865 );
buf ( n39023 , n32271 );
not ( n39024 , n31903 );
buf ( n39025 , n31899 );
not ( n39026 , n39025 );
or ( n39027 , n39024 , n39026 );
not ( n39028 , n31904 );
nand ( n39029 , n39027 , n39028 );
buf ( n39030 , n384392 );
nand ( n39031 , n39029 , n39030 );
not ( n39032 , n31850 );
and ( n39033 , n39032 , n31857 );
not ( n39034 , n39032 );
and ( n39035 , n39034 , n31858 );
nor ( n39036 , n39033 , n39035 );
not ( n39037 , n31883 );
nand ( n39038 , n39036 , n39037 );
not ( n39039 , n31941 );
not ( n39040 , n31944 );
and ( n39041 , n39039 , n39040 );
not ( n39042 , n39039 );
and ( n39043 , n39042 , n31944 );
nor ( n39044 , n39041 , n39043 );
not ( n39045 , n387122 );
and ( n39046 , n39044 , n39045 );
nor ( n39047 , n19512 , n33958 );
nor ( n39048 , n39046 , n39047 );
and ( n39049 , n39031 , n39038 , n39048 );
not ( n39050 , n381497 );
or ( n39051 , n383427 , n39050 );
nand ( n39052 , n39051 , n384642 );
nand ( n39053 , n39052 , RI15b63870_1261);
and ( n39054 , n384655 , n383427 , n386926 );
and ( n39055 , n386930 , n19630 );
nor ( n39056 , n39054 , n39055 );
nand ( n39057 , n39049 , n39053 , n39056 );
buf ( n39058 , n39057 );
buf ( n39059 , n32271 );
buf ( n39060 , n22343 );
not ( n39061 , n21446 );
not ( n39062 , n39061 );
buf ( n39063 , n21226 );
not ( n39064 , n39063 );
not ( n39065 , n39064 );
not ( n39066 , n39065 );
not ( n39067 , n22663 );
or ( n39068 , n39066 , n39067 );
not ( n39069 , n22660 );
and ( n39070 , n39069 , n21453 );
not ( n39071 , n22661 );
nor ( n39072 , n39070 , n39071 );
or ( n39073 , n39072 , n39065 );
nand ( n39074 , n39068 , n39073 );
not ( n39075 , n39074 );
or ( n39076 , n39062 , n39075 );
or ( n39077 , n39074 , n39061 );
nand ( n39078 , n39076 , n39077 );
and ( n39079 , n39078 , n22685 );
not ( n39080 , n37828 );
and ( n39081 , n39064 , n21580 );
not ( n39082 , n39063 );
nor ( n39083 , n39082 , n21580 );
nor ( n39084 , n39081 , n39083 );
not ( n39085 , n39084 );
and ( n39086 , n39080 , n39085 );
and ( n39087 , n37828 , n39084 );
nor ( n39088 , n39086 , n39087 );
or ( n39089 , n39088 , n21744 );
nand ( n39090 , n21227 , n20963 );
not ( n39091 , n39090 );
buf ( n39092 , n37860 );
not ( n39093 , n39092 );
or ( n39094 , n39091 , n39093 );
or ( n39095 , n39092 , n39090 );
nand ( n39096 , n39094 , n39095 );
and ( n39097 , n21354 , n39096 );
and ( n39098 , n21751 , RI15b57840_851);
nor ( n39099 , n39097 , n39098 );
nand ( n39100 , n39089 , n39099 );
nor ( n39101 , n39079 , n39100 );
and ( n39102 , n21788 , RI15b56940_819);
buf ( n39103 , n21766 );
and ( n39104 , n39103 , n21813 );
not ( n39105 , RI15b56940_819);
not ( n39106 , n17527 );
not ( n39107 , n39106 );
or ( n39108 , n39105 , n39107 );
or ( n39109 , n39106 , RI15b56940_819);
nand ( n39110 , n39108 , n39109 );
and ( n39111 , n21794 , n39110 );
nor ( n39112 , n39102 , n39104 , n39111 );
nand ( n39113 , n39101 , n39112 );
buf ( n39114 , n39113 );
not ( n39115 , RI15b584e8_878);
or ( n39116 , n35682 , n39115 );
or ( n39117 , RI15b58560_879 , n380788 );
not ( n39118 , n380774 );
not ( n39119 , n35682 );
nor ( n39120 , n39119 , n383598 );
not ( n39121 , n39120 );
or ( n39122 , n39118 , n39121 );
nand ( n39123 , n39122 , RI15b58560_879);
nand ( n39124 , n39116 , n39117 , n39123 );
buf ( n39125 , n39124 );
buf ( n39126 , n32672 );
and ( n39127 , n22646 , RI15b454b0_229);
and ( n39128 , n22648 , RI15b51918_648);
nor ( n39129 , n39127 , n39128 );
not ( n39130 , n39129 );
buf ( n39131 , n39130 );
buf ( n39132 , n383498 );
buf ( n39133 , n386760 );
not ( n39134 , n38065 );
not ( n39135 , n39134 );
not ( n39136 , n33370 );
or ( n39137 , n39135 , n39136 );
and ( n39138 , n33196 , n38067 );
or ( n39139 , n38077 , n385341 );
or ( n39140 , n22241 , n38081 );
or ( n39141 , n38075 , n33201 );
nand ( n39142 , n39139 , n39140 , n39141 );
nor ( n39143 , n39138 , n39142 );
nand ( n39144 , n39137 , n39143 );
buf ( n39145 , n39144 );
buf ( n39146 , n383613 );
buf ( n39147 , n381872 );
buf ( n39148 , n20663 );
buf ( n39149 , n33382 );
not ( n39150 , n36121 );
not ( n39151 , n39150 );
not ( n39152 , n32129 );
or ( n39153 , n39151 , n39152 );
and ( n39154 , n36133 , RI15b437a0_167);
or ( n39155 , n32141 , n36124 );
not ( n39156 , n36139 );
not ( n39157 , n32148 );
and ( n39158 , n39156 , n39157 );
not ( n39159 , n32150 );
and ( n39160 , n39159 , n36136 );
nor ( n39161 , n39158 , n39160 );
nand ( n39162 , n39155 , n39161 );
nor ( n39163 , n39154 , n39162 );
nand ( n39164 , n39153 , n39163 );
buf ( n39165 , n39164 );
buf ( n39166 , n379844 );
buf ( n39167 , n383498 );
buf ( n39168 , n36560 );
buf ( n39169 , n34242 );
nand ( n39170 , n39168 , n39169 );
buf ( n39171 , n34132 );
nor ( n39172 , n39170 , n39171 );
buf ( n39173 , n39172 );
nand ( n39174 , n39173 , n379785 );
not ( n39175 , n39174 );
not ( n39176 , n36496 );
or ( n39177 , n39175 , n39176 );
buf ( n39178 , n34070 );
buf ( n39179 , n39178 );
buf ( n39180 , n39179 );
nand ( n39181 , n39177 , n39180 );
nor ( n39182 , n39173 , n39179 );
nand ( n39183 , n36502 , n39182 );
buf ( n39184 , n34468 );
not ( n39185 , n39184 );
nor ( n39186 , n34311 , n39185 );
buf ( n39187 , n34428 );
and ( n39188 , n39186 , n39187 );
buf ( n39189 , n34337 );
nand ( n39190 , n39188 , n39189 );
not ( n39191 , n34467 );
nor ( n39192 , n39190 , n39191 );
not ( n39193 , n34460 );
and ( n39194 , n39192 , n39193 );
buf ( n39195 , n34453 );
nand ( n39196 , n39194 , n39195 );
buf ( n39197 , n39196 );
buf ( n39198 , n34442 );
not ( n39199 , n39198 );
and ( n39200 , n39197 , n39199 );
not ( n39201 , n39197 );
buf ( n39202 , n39198 );
and ( n39203 , n39201 , n39202 );
nor ( n39204 , n39200 , n39203 );
and ( n39205 , n39204 , n36513 );
not ( n39206 , RI15b5de70_1069);
not ( n39207 , n34651 );
or ( n39208 , n39206 , n39207 );
not ( n39209 , RI15b64068_1278);
or ( n39210 , n36518 , n39209 );
nand ( n39211 , n39208 , n39210 );
nor ( n39212 , n39205 , n39211 );
nand ( n39213 , n39181 , n39183 , n39212 );
buf ( n39214 , n39213 );
not ( n39215 , RI15b50fb8_628);
nor ( n39216 , n39215 , n381632 );
and ( n39217 , n382692 , n39216 );
and ( n39218 , n18156 , n36842 );
nor ( n39219 , n39218 , n18219 );
nand ( n39220 , n383165 , n39219 , n383163 , n18169 );
and ( n39221 , n39220 , RI15b51030_629);
nor ( n39222 , n39217 , n39221 );
not ( n39223 , n39222 );
buf ( n39224 , n39223 );
buf ( n39225 , n384203 );
buf ( n39226 , n379802 );
buf ( n39227 , n32255 );
buf ( n39228 , n19651 );
buf ( n39229 , n384203 );
buf ( n39230 , n383345 );
and ( n39231 , n379822 , RI15b65940_1331);
and ( n39232 , n379825 , RI15b48570_333);
nor ( n39233 , n39231 , n39232 );
nand ( n39234 , n379832 , RI15b46860_271);
nand ( n39235 , n379835 , n22283 );
nand ( n39236 , n39233 , n39234 , n39235 );
buf ( n39237 , n39236 );
buf ( n39238 , n383613 );
buf ( n39239 , n32981 );
buf ( n39240 , n380903 );
or ( n39241 , n22315 , n37663 );
and ( n39242 , n22326 , n37666 );
or ( n39243 , n37675 , n385574 );
or ( n39244 , n22334 , n37679 );
or ( n39245 , n37673 , n22336 );
nand ( n39246 , n39243 , n39244 , n39245 );
nor ( n39247 , n39242 , n39246 );
nand ( n39248 , n39241 , n39247 );
buf ( n39249 , n39248 );
buf ( n39250 , n379802 );
buf ( n39251 , n380865 );
buf ( n39252 , n380940 );
buf ( n39253 , n22714 );
or ( n39254 , n20627 , RI15b3fc18_40);
nand ( n39255 , n39254 , n385209 );
nor ( n39256 , n22232 , n39255 , n22234 );
or ( n39257 , n39256 , n20008 );
nand ( n39258 , n39257 , n36774 );
buf ( n39259 , n39258 );
buf ( n39260 , n32160 );
buf ( n39261 , n22716 );
buf ( n39262 , n32255 );
buf ( n39263 , n22714 );
not ( n39264 , n381014 );
not ( n39265 , n39264 );
or ( n39266 , n39265 , n22254 );
nand ( n39267 , n35525 , RI15b541e0_735);
nand ( n39268 , n39266 , n39267 );
buf ( n39269 , n39268 );
not ( n39270 , RI15b65b98_1336);
not ( n39271 , n35176 );
or ( n39272 , n39270 , n39271 );
nand ( n39273 , n379835 , n22245 );
nand ( n39274 , n35187 , RI15b487c8_338);
buf ( n39275 , n38199 );
and ( n39276 , n386554 , n39275 );
not ( n39277 , RI15b487c8_338);
not ( n39278 , n35343 );
or ( n39279 , n39277 , n39278 );
or ( n39280 , n35343 , RI15b487c8_338);
nand ( n39281 , n39279 , n39280 );
and ( n39282 , n35363 , n39281 );
nor ( n39283 , n39276 , n39282 );
and ( n39284 , n39273 , n39274 , n39283 );
nand ( n39285 , n39272 , n39284 );
buf ( n39286 , n39285 );
buf ( n39287 , n31033 );
buf ( n39288 , n382052 );
buf ( n39289 , n22343 );
nor ( n39290 , n386513 , n386556 );
or ( n39291 , n39290 , RI15b43ae8_174);
or ( n39292 , n379830 , n20510 );
nand ( n39293 , n39292 , n20501 );
not ( n39294 , n379817 );
nand ( n39295 , n30902 , n386535 , n39293 , n39294 );
and ( n39296 , n39295 , RI15b43ae8_174);
buf ( n39297 , n386302 );
not ( n39298 , n39297 );
nand ( n39299 , n39298 , RI15b43ae8_174);
or ( n39300 , n381050 , n39299 );
buf ( n39301 , n39297 );
or ( n39302 , n39301 , RI15b43ae8_174);
nand ( n39303 , n39302 , n385739 );
and ( n39304 , n386258 , n39303 );
and ( n39305 , n22393 , RI15b4b180_427);
buf ( n39306 , n386104 );
and ( n39307 , n386011 , n39306 );
nor ( n39308 , n39304 , n39305 , n39307 );
nand ( n39309 , n39300 , n39308 );
nor ( n39310 , n39296 , n39309 );
nand ( n39311 , n39291 , n39310 );
buf ( n39312 , n39311 );
buf ( n39313 , n379847 );
buf ( n39314 , n380203 );
buf ( n39315 , n17499 );
buf ( n39316 , n382052 );
not ( n39317 , n37663 );
not ( n39318 , n39317 );
not ( n39319 , n33369 );
not ( n39320 , n39319 );
or ( n39321 , n39318 , n39320 );
and ( n39322 , n33196 , n37666 );
not ( n39323 , RI15b42b70_141);
or ( n39324 , n37675 , n39323 );
or ( n39325 , n22241 , n37679 );
or ( n39326 , n37673 , n33201 );
nand ( n39327 , n39324 , n39325 , n39326 );
nor ( n39328 , n39322 , n39327 );
nand ( n39329 , n39321 , n39328 );
buf ( n39330 , n39329 );
buf ( n39331 , n384203 );
buf ( n39332 , n20665 );
buf ( n39333 , n384810 );
not ( n39334 , n39333 );
not ( n39335 , n39334 );
or ( n39336 , n31053 , n39335 );
not ( n39337 , n384815 );
nand ( n39338 , n384907 , n39337 );
and ( n39339 , n36536 , RI15b61188_1178);
and ( n39340 , n383945 , RI15b58830_885);
and ( n39341 , n383949 , RI15b5a630_949);
nor ( n39342 , n39340 , n39341 );
and ( n39343 , n383955 , RI15b5adb0_965);
and ( n39344 , n383960 , RI15b5a9f0_957);
nor ( n39345 , n39343 , n39344 );
and ( n39346 , n383965 , RI15b5b170_973);
and ( n39347 , n383970 , RI15b59eb0_933);
and ( n39348 , n383972 , RI15b5a270_941);
nor ( n39349 , n39347 , n39348 );
and ( n39350 , n383975 , RI15b59730_917);
and ( n39351 , n383977 , RI15b59af0_925);
nor ( n39352 , n39350 , n39351 );
and ( n39353 , n383982 , RI15b5bcb0_997);
and ( n39354 , n383984 , RI15b5b8f0_989);
nor ( n39355 , n39353 , n39354 );
and ( n39356 , n383987 , RI15b5c070_1005);
and ( n39357 , n383989 , RI15b5b530_981);
nor ( n39358 , n39356 , n39357 );
nand ( n39359 , n39349 , n39352 , n39355 , n39358 );
and ( n39360 , n383968 , n39359 );
and ( n39361 , n383994 , RI15b58bf0_893);
nor ( n39362 , n39346 , n39360 , n39361 );
and ( n39363 , n383997 , RI15b58fb0_901);
and ( n39364 , n383999 , RI15b59370_909);
nor ( n39365 , n39363 , n39364 );
nand ( n39366 , n39342 , n39345 , n39362 , n39365 );
not ( n39367 , n31122 );
buf ( n39368 , n39367 );
and ( n39369 , n39366 , n39368 );
not ( n39370 , RI15b61188_1178);
not ( n39371 , n31070 );
not ( n39372 , n39371 );
or ( n39373 , n39370 , n39372 );
or ( n39374 , n39371 , RI15b61188_1178);
nand ( n39375 , n39373 , n39374 );
and ( n39376 , n36541 , n39375 );
nor ( n39377 , n39339 , n39369 , n39376 );
nand ( n39378 , n39336 , n39338 , n39377 );
buf ( n39379 , n39378 );
not ( n39380 , n31151 );
not ( n39381 , n39380 );
not ( n39382 , n384726 );
or ( n39383 , n39381 , n39382 );
and ( n39384 , n384737 , n31164 );
or ( n39385 , n31175 , n17741 );
not ( n39386 , n35490 );
or ( n39387 , n39386 , n31182 );
or ( n39388 , n31173 , n384759 );
nand ( n39389 , n39385 , n39387 , n39388 );
nor ( n39390 , n39384 , n39389 );
nand ( n39391 , n39383 , n39390 );
buf ( n39392 , n39391 );
buf ( n39393 , n20665 );
buf ( n39394 , n382073 );
buf ( n39395 , n30992 );
buf ( n39396 , n22479 );
and ( n39397 , n32747 , RI15b428a0_135);
and ( n39398 , n32753 , RI15b415e0_95);
and ( n39399 , n32755 , RI15b419a0_103);
nor ( n39400 , n39398 , n39399 );
and ( n39401 , n32759 , RI15b40e60_79);
and ( n39402 , n32762 , RI15b41220_87);
nor ( n39403 , n39401 , n39402 );
and ( n39404 , n32766 , RI15b433e0_159);
and ( n39405 , n32768 , RI15b43020_151);
nor ( n39406 , n39404 , n39405 );
and ( n39407 , n32771 , RI15b437a0_167);
and ( n39408 , n32773 , RI15b42c60_143);
nor ( n39409 , n39407 , n39408 );
nand ( n39410 , n39400 , n39403 , n39406 , n39409 );
and ( n39411 , n36022 , n39410 );
and ( n39412 , n32781 , RI15b40320_55);
nor ( n39413 , n39397 , n39411 , n39412 );
and ( n39414 , n32785 , RI15b424e0_127);
and ( n39415 , n32787 , RI15b42120_119);
nor ( n39416 , n39414 , n39415 );
and ( n39417 , n32792 , RI15b3ff60_47);
and ( n39418 , n32794 , RI15b41d60_111);
nor ( n39419 , n39417 , n39418 );
and ( n39420 , n32797 , RI15b406e0_63);
and ( n39421 , n32800 , RI15b40aa0_71);
nor ( n39422 , n39420 , n39421 );
nand ( n39423 , n39413 , n39416 , n39419 , n39422 );
not ( n39424 , n39423 );
or ( n39425 , n39424 , n32807 );
and ( n39426 , n381055 , RI15b497b8_372);
not ( n39427 , RI15b497b8_372);
not ( n39428 , n32818 );
or ( n39429 , n39427 , n39428 );
or ( n39430 , n32818 , RI15b497b8_372);
nand ( n39431 , n39429 , n39430 );
and ( n39432 , n381076 , n39431 );
nor ( n39433 , n39426 , n39432 );
nand ( n39434 , n39425 , n39433 );
buf ( n39435 , n39434 );
buf ( n39436 , n382065 );
buf ( n39437 , n387159 );
buf ( n39438 , n32160 );
not ( n39439 , RI15b540f0_733);
not ( n39440 , n32244 );
or ( n39441 , n39439 , n39440 );
and ( n39442 , n32247 , RI15b656e8_1326);
and ( n39443 , n32249 , RI15b60558_1152);
nor ( n39444 , n39442 , n39443 );
nand ( n39445 , n39441 , n39444 );
buf ( n39446 , n39445 );
buf ( n39447 , n30992 );
buf ( n39448 , n20665 );
or ( n39449 , n35852 , n35869 );
not ( n39450 , n35884 );
and ( n39451 , n39450 , RI15b40a28_70);
or ( n39452 , n35582 , n35888 );
or ( n39453 , n35856 , n35882 );
or ( n39454 , n35871 , n35858 );
nand ( n39455 , n39452 , n39453 , n39454 );
nor ( n39456 , n39451 , n39455 );
nand ( n39457 , n39449 , n39456 );
buf ( n39458 , n39457 );
not ( n39459 , n35896 );
not ( n39460 , n33174 );
or ( n39461 , n39459 , n39460 );
not ( n39462 , n35900 );
and ( n39463 , n33196 , n39462 );
or ( n39464 , n35911 , n385292 );
or ( n39465 , n22241 , n35917 );
or ( n39466 , n35909 , n33201 );
nand ( n39467 , n39464 , n39465 , n39466 );
nor ( n39468 , n39463 , n39467 );
nand ( n39469 , n39461 , n39468 );
buf ( n39470 , n39469 );
buf ( n39471 , n381566 );
buf ( n39472 , n22005 );
buf ( n39473 , n386760 );
not ( n39474 , RI15b47490_297);
not ( n39475 , n385213 );
or ( n39476 , n39474 , n39475 );
and ( n39477 , n385221 , RI15b48a20_343);
and ( n39478 , n20631 , RI15b46d10_281);
nor ( n39479 , n39477 , n39478 );
nand ( n39480 , n39476 , n39479 );
buf ( n39481 , n39480 );
buf ( n39482 , n380865 );
buf ( n39483 , n383174 );
buf ( n39484 , n386563 );
buf ( n39485 , n379403 );
buf ( n39486 , n22738 );
buf ( n39487 , n381872 );
buf ( n39488 , n386532 );
buf ( n39489 , n31719 );
buf ( n39490 , n381004 );
buf ( n39491 , n381490 );
not ( n39492 , RI15b471c0_291);
not ( n39493 , n385213 );
or ( n39494 , n39492 , n39493 );
and ( n39495 , n385221 , RI15b48750_337);
and ( n39496 , n20631 , RI15b46a40_275);
nor ( n39497 , n39495 , n39496 );
nand ( n39498 , n39494 , n39497 );
buf ( n39499 , n39498 );
buf ( n39500 , n32160 );
buf ( n39501 , n380203 );
buf ( n39502 , n22343 );
not ( n39503 , n386514 );
or ( n39504 , n39503 , n386368 );
and ( n39505 , n386540 , RI15b43e30_181);
and ( n39506 , n386549 , n385368 );
and ( n39507 , n386556 , n386061 );
nor ( n39508 , n39505 , n39506 , n39507 );
nand ( n39509 , n39504 , n38212 , n39508 );
buf ( n39510 , n39509 );
buf ( n39511 , n379847 );
buf ( n39512 , n32160 );
buf ( n39513 , n22007 );
buf ( n39514 , n379844 );
or ( n39515 , n386588 , n382936 );
and ( n39516 , n386600 , n382934 );
not ( n39517 , RI15b59730_917);
or ( n39518 , n382949 , n39517 );
or ( n39519 , n34706 , n382965 );
or ( n39520 , n382947 , n386627 );
nand ( n39521 , n39518 , n39519 , n39520 );
nor ( n39522 , n39516 , n39521 );
nand ( n39523 , n39515 , n39522 );
buf ( n39524 , n39523 );
not ( n39525 , n382683 );
buf ( n39526 , n382629 );
not ( n39527 , n39526 );
not ( n39528 , n39527 );
or ( n39529 , n39525 , n39528 );
nand ( n39530 , n39529 , n382682 );
not ( n39531 , n39527 );
nor ( n39532 , n39531 , RI15b556f8_780);
nor ( n39533 , n39530 , n39532 );
not ( n39534 , RI15b55770_781);
or ( n39535 , n39533 , n39534 );
not ( n39536 , RI15b55770_781);
not ( n39537 , RI15b556f8_780);
nor ( n39538 , n382683 , n39537 );
and ( n39539 , n382688 , n39536 , n39538 );
nor ( n39540 , n382691 , n384711 );
nor ( n39541 , n39539 , n39540 );
nand ( n39542 , n39535 , n39541 );
buf ( n39543 , n39542 );
buf ( n39544 , n22009 );
buf ( n39545 , n22007 );
buf ( n39546 , n379893 );
buf ( n39547 , n384357 );
nor ( n39548 , n32546 , n39547 );
not ( n39549 , n39548 );
buf ( n39550 , n39547 );
nand ( n39551 , n32546 , n39550 );
nand ( n39552 , n39549 , n39551 );
nand ( n39553 , n39552 , n39030 );
not ( n39554 , n32626 );
not ( n39555 , n384592 );
and ( n39556 , n39554 , n39555 );
not ( n39557 , n39554 );
and ( n39558 , n39557 , n384592 );
nor ( n39559 , n39556 , n39558 );
and ( n39560 , n39559 , n387123 );
not ( n39561 , n32641 );
not ( n39562 , n32638 );
and ( n39563 , n39561 , n39562 );
and ( n39564 , n32641 , n32638 );
nor ( n39565 , n39563 , n39564 );
or ( n39566 , n39565 , n384494 );
or ( n39567 , n19512 , n379437 );
nand ( n39568 , n39566 , n39567 );
nor ( n39569 , n39560 , n39568 );
nand ( n39570 , n39553 , n39569 );
not ( n39571 , n39570 );
and ( n39572 , n31792 , n384592 );
buf ( n39573 , n37610 );
not ( n39574 , n39573 );
or ( n39575 , n39547 , n39574 );
or ( n39576 , n31771 , n384351 );
or ( n39577 , n32638 , n31779 );
nand ( n39578 , n39575 , n39576 , n39577 );
nor ( n39579 , n39572 , n39578 );
nand ( n39580 , n39571 , n39579 );
buf ( n39581 , n39580 );
buf ( n39582 , n21800 );
nand ( n39583 , n31426 , n31429 );
not ( n39584 , n379291 );
buf ( n39585 , n379301 );
and ( n39586 , n39584 , n39585 );
not ( n39587 , n39584 );
not ( n39588 , n39585 );
and ( n39589 , n39587 , n39588 );
nor ( n39590 , n39586 , n39589 );
not ( n39591 , n39590 );
nor ( n39592 , n39583 , n39591 );
buf ( n39593 , n379302 );
buf ( n39594 , n39593 );
not ( n39595 , n39594 );
buf ( n39596 , n31685 );
not ( n39597 , n39596 );
and ( n39598 , n39595 , n39597 );
and ( n39599 , n39594 , n39596 );
nor ( n39600 , n39598 , n39599 );
and ( n39601 , n39592 , n39600 );
not ( n39602 , n39593 );
nand ( n39603 , n39602 , n39596 );
not ( n39604 , n379330 );
and ( n39605 , n39603 , n39604 );
or ( n39606 , n39603 , n39604 );
nand ( n39607 , n39606 , n379327 );
nor ( n39608 , n39605 , n39607 );
and ( n39609 , n39601 , n39608 );
not ( n39610 , n39603 );
nand ( n39611 , n39610 , n39604 );
not ( n39612 , n379319 );
and ( n39613 , n39611 , n39612 );
nor ( n39614 , n39613 , n379334 );
not ( n39615 , n39614 );
and ( n39616 , n39609 , n39615 );
not ( n39617 , n39609 );
and ( n39618 , n39617 , n39614 );
nor ( n39619 , n39616 , n39618 );
not ( n39620 , n39619 );
not ( n39621 , n39608 );
not ( n39622 , n39601 );
not ( n39623 , n39622 );
or ( n39624 , n39621 , n39623 );
or ( n39625 , n39622 , n39608 );
nand ( n39626 , n39624 , n39625 );
nor ( n39627 , n39583 , n39591 );
not ( n39628 , n39627 );
not ( n39629 , n39628 );
not ( n39630 , n39600 );
and ( n39631 , n39629 , n39630 );
and ( n39632 , n39628 , n39600 );
nor ( n39633 , n39631 , n39632 );
not ( n39634 , n39590 );
not ( n39635 , n39583 );
or ( n39636 , n39634 , n39635 );
buf ( n39637 , n39583 );
or ( n39638 , n39637 , n39590 );
nand ( n39639 , n39636 , n39638 );
not ( n39640 , n31592 );
nand ( n39641 , n39640 , n31434 );
nor ( n39642 , n39639 , n39641 );
nand ( n39643 , n39633 , n39642 );
nor ( n39644 , n39626 , n39643 );
nand ( n39645 , n39620 , n39644 );
nand ( n39646 , n39609 , n39615 );
not ( n39647 , n379334 );
not ( n39648 , n379045 );
and ( n39649 , n39647 , n39648 );
and ( n39650 , n379334 , n379045 );
nor ( n39651 , n39649 , n39650 );
and ( n39652 , n39646 , n39651 );
not ( n39653 , n39646 );
not ( n39654 , n39651 );
and ( n39655 , n39653 , n39654 );
nor ( n39656 , n39652 , n39655 );
not ( n39657 , n39656 );
and ( n39658 , n39645 , n39657 );
not ( n39659 , n39645 );
and ( n39660 , n39659 , n39656 );
nor ( n39661 , n39658 , n39660 );
buf ( n39662 , n31602 );
not ( n39663 , n39662 );
or ( n39664 , n39661 , n39663 );
not ( n39665 , n379391 );
nand ( n39666 , n31665 , n31679 );
nor ( n39667 , n39666 , n31676 );
not ( n39668 , n31695 );
and ( n39669 , n39667 , n39668 );
nand ( n39670 , n39669 , n31687 );
nor ( n39671 , n39670 , n31672 );
buf ( n39672 , n39671 );
not ( n39673 , n39672 );
or ( n39674 , n39665 , n39673 );
nand ( n39675 , n39674 , n31700 );
and ( n39676 , n39675 , n39612 );
not ( n39677 , n31708 );
buf ( n39678 , n39677 );
not ( n39679 , n39678 );
nand ( n39680 , n39679 , n379319 );
or ( n39681 , n39672 , n39680 );
and ( n39682 , n379394 , RI15b583f8_876);
buf ( n39683 , n31712 );
and ( n39684 , n39683 , RI15b52200_667);
nor ( n39685 , n39682 , n39684 );
nand ( n39686 , n39681 , n39685 );
nor ( n39687 , n39676 , n39686 );
nand ( n39688 , n39664 , n39687 );
buf ( n39689 , n39688 );
buf ( n39690 , n385112 );
nand ( n39691 , n384054 , n33110 );
or ( n39692 , n31149 , n39691 );
nand ( n39693 , n384167 , n21337 );
not ( n39694 , n39693 );
and ( n39695 , n31161 , n39694 );
and ( n39696 , n39693 , n39691 , n383882 );
nor ( n39697 , n39696 , n21764 );
nor ( n39698 , n384173 , n33122 );
or ( n39699 , n39697 , n39698 );
nand ( n39700 , n39699 , n18154 );
or ( n39701 , n383865 , n384179 );
nand ( n39702 , n39700 , n39701 );
and ( n39703 , n39702 , n383901 );
or ( n39704 , n39703 , n17645 );
not ( n39705 , n39701 );
nor ( n39706 , n39698 , n39705 );
or ( n39707 , n39697 , n39706 );
or ( n39708 , n31179 , n39707 );
or ( n39709 , n39701 , n31184 );
nand ( n39710 , n39704 , n39708 , n39709 );
nor ( n39711 , n39695 , n39710 );
nand ( n39712 , n39692 , n39711 );
buf ( n39713 , n39712 );
buf ( n39714 , n383968 );
and ( n39715 , n38654 , RI15b5b3c8_978);
buf ( n39716 , n38657 );
buf ( n39717 , n39716 );
and ( n39718 , n39717 , RI15b5b008_970);
nor ( n39719 , n39715 , n39718 );
buf ( n39720 , n38660 );
buf ( n39721 , n39720 );
and ( n39722 , n39721 , RI15b5ac48_962);
buf ( n39723 , n38662 );
buf ( n39724 , n39723 );
and ( n39725 , n39724 , RI15b5a888_954);
nor ( n39726 , n39722 , n39725 );
buf ( n39727 , n38603 );
buf ( n39728 , n39727 );
and ( n39729 , n39728 , RI15b5a4c8_946);
buf ( n39730 , n38607 );
buf ( n39731 , n39730 );
and ( n39732 , n39731 , RI15b5a108_938);
nor ( n39733 , n39729 , n39732 );
buf ( n39734 , n38628 );
buf ( n39735 , n39734 );
and ( n39736 , n39735 , RI15b59d48_930);
buf ( n39737 , n38631 );
buf ( n39738 , n39737 );
and ( n39739 , n39738 , RI15b59988_922);
nor ( n39740 , n39736 , n39739 );
nand ( n39741 , n39719 , n39726 , n39733 , n39740 );
and ( n39742 , n39714 , n39741 );
not ( n39743 , n19494 );
nor ( n39744 , n39743 , n38620 );
buf ( n39745 , n38626 );
and ( n39746 , n39744 , n39745 );
and ( n39747 , n39746 , RI15b58e48_898);
not ( n39748 , n38641 );
nand ( n39749 , n19494 , n39748 );
buf ( n39750 , n38651 );
nor ( n39751 , n39749 , n39750 );
and ( n39752 , n39751 , RI15b5c2c8_1010);
nor ( n39753 , n39742 , n39747 , n39752 );
not ( n39754 , n38656 );
not ( n39755 , n39754 );
nor ( n39756 , n39749 , n39755 );
and ( n39757 , n39756 , RI15b5bf08_1002);
not ( n39758 , n39745 );
nor ( n39759 , n39749 , n39758 );
and ( n39760 , n39759 , RI15b5bb48_994);
nor ( n39761 , n39757 , n39760 );
not ( n39762 , n39750 );
and ( n39763 , n39744 , n39762 );
and ( n39764 , n39763 , RI15b595c8_914);
and ( n39765 , n39744 , n39754 );
and ( n39766 , n39765 , RI15b59208_906);
nor ( n39767 , n39764 , n39766 );
not ( n39768 , n38630 );
and ( n39769 , n39744 , n39768 );
and ( n39770 , n39769 , RI15b58a88_890);
not ( n39771 , n39749 );
and ( n39772 , n39771 , n39768 );
and ( n39773 , n39772 , RI15b5b788_986);
nor ( n39774 , n39770 , n39773 );
and ( n39775 , n39753 , n39761 , n39767 , n39774 );
not ( n39776 , n383929 );
not ( n39777 , n39776 );
or ( n39778 , n39775 , n39777 );
or ( n39779 , n386988 , n384021 );
not ( n39780 , n38483 );
and ( n39781 , n39780 , RI15b626a0_1223);
not ( n39782 , n39780 );
and ( n39783 , n39782 , n386988 );
nor ( n39784 , n39781 , n39783 );
or ( n39785 , n384024 , n39784 );
nand ( n39786 , n39778 , n39779 , n39785 );
buf ( n39787 , n39786 );
buf ( n39788 , n22738 );
buf ( n39789 , n22653 );
buf ( n39790 , n382073 );
not ( n39791 , n39178 );
nand ( n39792 , n39791 , n39172 );
nor ( n39793 , n39792 , n385039 );
buf ( n39794 , n34079 );
not ( n39795 , n39794 );
nand ( n39796 , n39793 , n39795 );
not ( n39797 , n39796 );
not ( n39798 , n36573 );
not ( n39799 , n39798 );
or ( n39800 , n39797 , n39799 );
buf ( n39801 , n36562 );
nand ( n39802 , n39800 , n39801 );
not ( n39803 , n34488 );
not ( n39804 , n39803 );
nor ( n39805 , n39196 , n39199 );
nand ( n39806 , n39804 , n39805 );
buf ( n39807 , n39806 );
not ( n39808 , n34447 );
and ( n39809 , n39807 , n39808 );
not ( n39810 , n39807 );
and ( n39811 , n39810 , n34447 );
nor ( n39812 , n39809 , n39811 );
not ( n39813 , n34645 );
buf ( n39814 , n39813 );
and ( n39815 , n39812 , n39814 );
not ( n39816 , RI15b5df60_1071);
not ( n39817 , n34651 );
or ( n39818 , n39816 , n39817 );
or ( n39819 , n36518 , n379431 );
nand ( n39820 , n39818 , n39819 );
nor ( n39821 , n39815 , n39820 );
not ( n39822 , n39792 );
not ( n39823 , n39794 );
nand ( n39824 , n39822 , n39823 );
not ( n39825 , n39801 );
nand ( n39826 , n36580 , n39824 , n39825 );
nand ( n39827 , n39802 , n39821 , n39826 );
buf ( n39828 , n39827 );
buf ( n39829 , n22408 );
not ( n39830 , n379925 );
not ( n39831 , n39830 );
not ( n39832 , n37697 );
not ( n39833 , n39832 );
or ( n39834 , n39831 , n39833 );
or ( n39835 , n381467 , n379926 );
nand ( n39836 , n39834 , n39835 );
and ( n39837 , n18060 , RI15b50f40_627);
not ( n39838 , n17603 );
nor ( n39839 , n39837 , n39838 );
nor ( n39840 , n32366 , n39839 );
not ( n39841 , n21555 );
not ( n39842 , n18116 );
or ( n39843 , n39841 , n39842 );
nand ( n39844 , n39843 , n21784 );
nor ( n39845 , n385156 , n39844 );
not ( n39846 , RI15b50f40_627);
nor ( n39847 , n39845 , n39846 );
nor ( n39848 , n39836 , n39840 , n39847 );
or ( n39849 , n39848 , n18078 );
and ( n39850 , n39220 , RI15b50f40_627);
and ( n39851 , n383915 , n379927 );
or ( n39852 , n21407 , n37927 );
or ( n39853 , n21364 , RI15b50dd8_624);
nand ( n39854 , n39852 , n39853 );
and ( n39855 , n32986 , n39854 );
nor ( n39856 , n39850 , n39851 , n39855 );
nand ( n39857 , n39849 , n39856 );
buf ( n39858 , n39857 );
buf ( n39859 , n383345 );
or ( n39860 , n35852 , n380909 );
and ( n39861 , n33080 , RI15b41ce8_110);
or ( n39862 , n35856 , n380926 );
or ( n39863 , n35582 , n380933 );
or ( n39864 , n380915 , n35858 );
nand ( n39865 , n39862 , n39863 , n39864 );
nor ( n39866 , n39861 , n39865 );
nand ( n39867 , n39860 , n39866 );
buf ( n39868 , n39867 );
buf ( n39869 , n382071 );
buf ( n39870 , n382537 );
buf ( n39871 , n384996 );
buf ( n39872 , n380903 );
buf ( n39873 , RI15b47238_292);
buf ( n39874 , n382069 );
not ( n39875 , n36951 );
or ( n39876 , n32430 , n39875 );
nand ( n39877 , n381417 , n381341 );
and ( n39878 , n386637 , RI15b54b40_755);
and ( n39879 , n382885 , n39065 );
not ( n39880 , RI15b54b40_755);
not ( n39881 , n382636 );
or ( n39882 , n39880 , n39881 );
or ( n39883 , n382636 , RI15b54b40_755);
nand ( n39884 , n39882 , n39883 );
and ( n39885 , n37449 , n39884 );
nor ( n39886 , n39878 , n39879 , n39885 );
and ( n39887 , n39877 , n39886 );
nand ( n39888 , n39876 , n39887 );
buf ( n39889 , n39888 );
buf ( n39890 , n383498 );
not ( n39891 , n32063 );
not ( n39892 , n39891 );
not ( n39893 , n382912 );
or ( n39894 , n39892 , n39893 );
and ( n39895 , n382931 , n32070 );
not ( n39896 , RI15b5a360_943);
or ( n39897 , n32081 , n39896 );
or ( n39898 , n382959 , n32086 );
or ( n39899 , n32079 , n382967 );
nand ( n39900 , n39897 , n39898 , n39899 );
nor ( n39901 , n39895 , n39900 );
nand ( n39902 , n39894 , n39901 );
buf ( n39903 , n39902 );
buf ( n39904 , n383345 );
buf ( n39905 , n385197 );
not ( n39906 , n38486 );
and ( n39907 , n39906 , RI15b62808_1226);
not ( n39908 , n39906 );
and ( n39909 , n39908 , n386993 );
nor ( n39910 , n39907 , n39909 );
or ( n39911 , n39910 , n384024 );
and ( n39912 , n384022 , RI15b62808_1226);
not ( n39913 , n38721 );
buf ( n39914 , n38694 );
not ( n39915 , n39914 );
or ( n39916 , n39913 , n39915 );
or ( n39917 , n39914 , n38721 );
nand ( n39918 , n39916 , n39917 );
and ( n39919 , n386746 , n39918 );
nor ( n39920 , n39912 , n39919 );
nand ( n39921 , n39911 , n39920 );
buf ( n39922 , n39921 );
not ( n39923 , n38825 );
not ( n39924 , n39923 );
not ( n39925 , n384726 );
or ( n39926 , n39924 , n39925 );
and ( n39927 , n35477 , n38828 );
or ( n39928 , n38837 , n17765 );
or ( n39929 , n39386 , n38841 );
or ( n39930 , n38835 , n384759 );
nand ( n39931 , n39928 , n39929 , n39930 );
nor ( n39932 , n39927 , n39931 );
nand ( n39933 , n39926 , n39932 );
buf ( n39934 , n39933 );
buf ( n39935 , n19655 );
buf ( n39936 , n384199 );
buf ( n39937 , n386563 );
buf ( n39938 , n379893 );
not ( n39939 , n385815 );
not ( n39940 , n39939 );
not ( n39941 , n39275 );
not ( n39942 , n39941 );
not ( n39943 , n30868 );
or ( n39944 , n39942 , n39943 );
nor ( n39945 , n30867 , n385368 );
nor ( n39946 , n39945 , n385808 );
nand ( n39947 , n39944 , n39946 );
not ( n39948 , n385822 );
nor ( n39949 , n39947 , n39948 );
nand ( n39950 , n39940 , n39949 );
not ( n39951 , n385795 );
nor ( n39952 , n39950 , n39951 );
nand ( n39953 , n39952 , n385791 );
and ( n39954 , n39953 , n385779 );
not ( n39955 , n39953 );
not ( n39956 , n385779 );
and ( n39957 , n39955 , n39956 );
nor ( n39958 , n39954 , n39957 );
not ( n39959 , n386020 );
nor ( n39960 , n39958 , n39959 );
buf ( n39961 , n386147 );
not ( n39962 , n386162 );
nand ( n39963 , n39961 , n39962 );
nor ( n39964 , n39963 , n386158 );
not ( n39965 , n386153 );
and ( n39966 , n39964 , n39965 );
nand ( n39967 , n39966 , n386172 );
and ( n39968 , n39967 , n386167 );
not ( n39969 , n39967 );
not ( n39970 , n386167 );
and ( n39971 , n39969 , n39970 );
nor ( n39972 , n39968 , n39971 );
buf ( n39973 , n386262 );
buf ( n39974 , n39973 );
not ( n39975 , n39974 );
or ( n39976 , n39972 , n39975 );
buf ( n39977 , n34736 );
not ( n39978 , n39977 );
not ( n39979 , n39978 );
buf ( n39980 , n34734 );
not ( n39981 , n39980 );
not ( n39982 , n34735 );
nand ( n39983 , n39981 , n39982 );
nand ( n39984 , n39979 , n39983 );
nand ( n39985 , n39984 , n386500 );
nand ( n39986 , n39976 , n39985 );
buf ( n39987 , n34783 );
buf ( n39988 , n39987 );
not ( n39989 , n39988 );
nor ( n39990 , n39989 , n20547 );
nor ( n39991 , n39960 , n39986 , n39990 );
and ( n39992 , n386517 , n39982 );
or ( n39993 , n386541 , n385251 );
or ( n39994 , n39956 , n386550 );
or ( n39995 , n39970 , n386557 );
nand ( n39996 , n39993 , n39994 , n39995 );
nor ( n39997 , n39992 , n39996 );
nand ( n39998 , n39991 , n39997 );
buf ( n39999 , n39998 );
buf ( n40000 , n32160 );
buf ( n40001 , n22655 );
buf ( n40002 , n386760 );
buf ( n40003 , n382065 );
buf ( n40004 , n22714 );
buf ( n40005 , n382067 );
not ( n40006 , n382509 );
nand ( n40007 , n40006 , RI15b48318_328);
nand ( n40008 , n36998 , n40007 );
and ( n40009 , n40008 , RI15b482a0_327);
buf ( n40010 , n40009 );
buf ( n40011 , n22404 );
or ( n40012 , n383180 , n33419 );
not ( n40013 , n33428 );
and ( n40014 , n40013 , RI15b5b4b8_980);
or ( n40015 , n383184 , n33416 );
buf ( n40016 , n383186 );
not ( n40017 , n40016 );
and ( n40018 , n33439 , n40017 );
not ( n40019 , n383192 );
and ( n40020 , n40019 , n33436 );
nor ( n40021 , n40018 , n40020 );
nand ( n40022 , n40015 , n40021 );
nor ( n40023 , n40014 , n40022 );
nand ( n40024 , n40012 , n40023 );
buf ( n40025 , n40024 );
not ( n40026 , RI15b539e8_718);
not ( n40027 , n383170 );
or ( n40028 , n40026 , n40027 );
not ( n40029 , RI15b54f00_763);
not ( n40030 , n383011 );
not ( n40031 , n40030 );
nand ( n40032 , n40031 , n382646 );
not ( n40033 , n40032 );
nand ( n40034 , n40033 , n383012 );
nand ( n40035 , n40034 , RI15b55770_781);
not ( n40036 , n40035 );
or ( n40037 , n40029 , n40036 );
or ( n40038 , n40035 , RI15b54f00_763);
nand ( n40039 , n40037 , n40038 );
not ( n40040 , n40039 );
not ( n40041 , RI15b54e88_762);
nand ( n40042 , n40032 , RI15b55770_781);
not ( n40043 , n40042 );
or ( n40044 , n40041 , n40043 );
or ( n40045 , n40042 , RI15b54e88_762);
nand ( n40046 , n40044 , n40045 );
not ( n40047 , RI15b54e10_761);
nand ( n40048 , n40030 , RI15b55770_781);
not ( n40049 , n40048 );
or ( n40050 , n40047 , n40049 );
or ( n40051 , n40048 , RI15b54e10_761);
nand ( n40052 , n40050 , n40051 );
not ( n40053 , n40052 );
nor ( n40054 , n33474 , n33463 );
nand ( n40055 , n40053 , n40054 );
nor ( n40056 , n40046 , n40055 );
nand ( n40057 , n40040 , n40056 );
or ( n40058 , n33454 , n40057 );
nand ( n40059 , n40058 , n33465 );
buf ( n40060 , n383045 );
not ( n40061 , RI15b55770_781);
nor ( n40062 , n40060 , n40061 );
and ( n40063 , n40062 , RI15b54f78_764);
not ( n40064 , n40062 );
and ( n40065 , n40064 , n383015 );
nor ( n40066 , n40063 , n40065 );
and ( n40067 , n40059 , n40066 );
not ( n40068 , n40057 );
nor ( n40069 , n40068 , n40066 );
and ( n40070 , n33476 , n40069 );
and ( n40071 , n383147 , RI15b53268_702);
nor ( n40072 , n40067 , n40070 , n40071 );
nand ( n40073 , n40028 , n40072 );
buf ( n40074 , n40073 );
buf ( n40075 , n385112 );
buf ( n40076 , n385195 );
buf ( n40077 , n385195 );
buf ( n40078 , n22406 );
buf ( n40079 , n383345 );
buf ( n40080 , n384199 );
not ( n40081 , n37009 );
not ( n40082 , n32129 );
or ( n40083 , n40081 , n40082 );
and ( n40084 , n36825 , RI15b42120_119);
or ( n40085 , n32141 , n36815 );
or ( n40086 , n32148 , n36830 );
or ( n40087 , n36822 , n32150 );
nand ( n40088 , n40085 , n40086 , n40087 );
nor ( n40089 , n40084 , n40088 );
nand ( n40090 , n40083 , n40089 );
buf ( n40091 , n40090 );
buf ( n40092 , n381490 );
buf ( n40093 , n31719 );
not ( n40094 , n386500 );
or ( n40095 , n34749 , n386441 );
nand ( n40096 , n40095 , n386447 );
not ( n40097 , n40096 );
or ( n40098 , n40094 , n40097 );
nand ( n40099 , n34758 , n34762 );
not ( n40100 , n386179 );
and ( n40101 , n40099 , n40100 );
not ( n40102 , n40099 );
and ( n40103 , n40102 , n386179 );
nor ( n40104 , n40101 , n40103 );
and ( n40105 , n40104 , n386264 );
nor ( n40106 , n34772 , n385906 );
not ( n40107 , n40106 );
not ( n40108 , n385877 );
and ( n40109 , n40107 , n40108 );
and ( n40110 , n40106 , n385877 );
nor ( n40111 , n40109 , n40110 );
not ( n40112 , n34779 );
or ( n40113 , n40111 , n40112 );
or ( n40114 , n34785 , n382120 );
nand ( n40115 , n40113 , n40114 );
nor ( n40116 , n40105 , n40115 );
nand ( n40117 , n40098 , n40116 );
not ( n40118 , n40117 );
not ( n40119 , n19848 );
not ( n40120 , n20637 );
or ( n40121 , n40119 , n40120 );
nand ( n40122 , n40121 , n34798 );
and ( n40123 , n40122 , RI15b4abe0_415);
or ( n40124 , n34801 , n19848 , RI15b4abe0_415);
or ( n40125 , n32504 , n22216 );
nand ( n40126 , n40124 , n40125 );
nor ( n40127 , n40123 , n40126 );
nand ( n40128 , n40118 , n40127 );
buf ( n40129 , n40128 );
buf ( n40130 , n382067 );
buf ( n40131 , n386879 );
or ( n40132 , n40131 , n22473 );
buf ( n40133 , n383474 );
nand ( n40134 , n40132 , n40133 );
nand ( n40135 , n40134 , n386885 );
not ( n40136 , n386885 );
nand ( n40137 , n40136 , n387011 , n40131 );
not ( n40138 , n386981 );
and ( n40139 , n40138 , n34816 );
not ( n40140 , n34823 );
nor ( n40141 , n40139 , n40140 );
not ( n40142 , RI15b624c0_1219);
or ( n40143 , n40141 , n40142 );
not ( n40144 , n34810 );
not ( n40145 , n40144 );
and ( n40146 , n40145 , RI15b642c0_1283);
or ( n40147 , n40138 , n34826 , RI15b624c0_1219);
and ( n40148 , n387036 , RI15b642c0_1283);
not ( n40149 , n387036 );
and ( n40150 , n40149 , n379436 );
nor ( n40151 , n40148 , n40150 );
or ( n40152 , n34833 , n40151 );
nand ( n40153 , n40147 , n40152 );
nor ( n40154 , n40146 , n40153 );
nand ( n40155 , n40143 , n40154 );
nand ( n40156 , n40155 , n19201 );
and ( n40157 , n22423 , RI15b642c0_1283);
and ( n40158 , n19599 , RI15b633c0_1251);
nor ( n40159 , n40157 , n40158 , n19513 );
nand ( n40160 , n40135 , n40137 , n40156 , n40159 );
buf ( n40161 , n40160 );
buf ( n40162 , n386762 );
buf ( n40163 , RI15b5e668_1086);
buf ( n40164 , n22343 );
buf ( n40165 , n386513 );
not ( n40166 , n40165 );
or ( n40167 , n40166 , n386313 );
and ( n40168 , n386540 , RI15b43cc8_178);
or ( n40169 , n386550 , n385550 );
or ( n40170 , n386557 , n386087 );
nand ( n40171 , n40169 , n40170 );
nor ( n40172 , n40168 , n40171 );
buf ( n40173 , n385543 );
buf ( n40174 , n40173 );
and ( n40175 , n386313 , n40174 );
not ( n40176 , n386313 );
not ( n40177 , n40174 );
and ( n40178 , n40176 , n40177 );
nor ( n40179 , n40175 , n40178 );
not ( n40180 , n40179 );
not ( n40181 , n386335 );
not ( n40182 , n386339 );
nand ( n40183 , n386308 , n40182 );
not ( n40184 , n40183 );
or ( n40185 , n40181 , n40184 );
nand ( n40186 , n40185 , n386352 );
not ( n40187 , n40186 );
or ( n40188 , n40180 , n40187 );
or ( n40189 , n40186 , n40179 );
nand ( n40190 , n40188 , n40189 );
and ( n40191 , n386500 , n40190 );
not ( n40192 , n385550 );
not ( n40193 , n385758 );
not ( n40194 , n40193 );
or ( n40195 , n40192 , n40194 );
or ( n40196 , n40193 , n385550 );
nand ( n40197 , n40195 , n40196 );
and ( n40198 , n40197 , n40174 );
not ( n40199 , n40197 );
not ( n40200 , n40174 );
and ( n40201 , n40199 , n40200 );
nor ( n40202 , n40198 , n40201 );
or ( n40203 , n386013 , n40202 );
and ( n40204 , n386120 , n40173 );
not ( n40205 , n386120 );
not ( n40206 , n40173 );
and ( n40207 , n40205 , n40206 );
nor ( n40208 , n40204 , n40207 );
and ( n40209 , n40208 , n386087 );
nor ( n40210 , n40208 , n386087 );
nor ( n40211 , n40209 , n40210 );
or ( n40212 , n386259 , n40211 );
or ( n40213 , n383358 , n31821 );
nand ( n40214 , n40203 , n40212 , n40213 );
nor ( n40215 , n40191 , n40214 );
nand ( n40216 , n40167 , n40172 , n40215 );
buf ( n40217 , n40216 );
buf ( n40218 , n36854 );
buf ( n40219 , n22653 );
buf ( n40220 , n22740 );
buf ( n40221 , n31979 );
buf ( n40222 , n385112 );
and ( n40223 , n384166 , n384056 );
and ( n40224 , n383875 , n33122 );
nor ( n40225 , n40223 , n40224 );
not ( n40226 , n21775 );
or ( n40227 , n40225 , n40226 );
or ( n40228 , n17998 , n36844 );
and ( n40229 , n21764 , n383862 );
and ( n40230 , n383915 , n383830 );
nor ( n40231 , n40229 , n40230 );
nand ( n40232 , n40227 , n40228 , n40231 );
buf ( n40233 , n40232 );
buf ( n40234 , n382537 );
buf ( n40235 , n387159 );
not ( n40236 , RI15b62cb8_1236);
or ( n40237 , n19607 , n40236 );
not ( n40238 , n19434 );
or ( n40239 , n19431 , n40238 );
nand ( n40240 , n40239 , n19421 );
buf ( n40241 , n18544 );
buf ( n40242 , n40241 );
not ( n40243 , n40242 );
and ( n40244 , n40240 , n40243 );
and ( n40245 , n19435 , n40242 );
nor ( n40246 , n40244 , n40245 );
not ( n40247 , n40246 );
not ( n40248 , n19456 );
and ( n40249 , n40247 , n40248 );
and ( n40250 , n40246 , n19456 );
nor ( n40251 , n40249 , n40250 );
or ( n40252 , n40251 , n19499 );
and ( n40253 , n19343 , n40243 );
not ( n40254 , n19343 );
and ( n40255 , n40254 , n40242 );
nor ( n40256 , n40253 , n40255 );
not ( n40257 , n40256 );
not ( n40258 , n19321 );
and ( n40259 , n40257 , n40258 );
and ( n40260 , n40256 , n19321 );
nor ( n40261 , n40259 , n40260 );
or ( n40262 , n40261 , n19388 );
not ( n40263 , n19282 );
not ( n40264 , n18674 );
not ( n40265 , n40264 );
not ( n40266 , n18550 );
not ( n40267 , n40241 );
or ( n40268 , n40266 , n40267 );
or ( n40269 , n40241 , n18550 );
nand ( n40270 , n40268 , n40269 );
not ( n40271 , n40270 );
and ( n40272 , n40265 , n40271 );
and ( n40273 , n40264 , n40270 );
nor ( n40274 , n40272 , n40273 );
not ( n40275 , n40274 );
and ( n40276 , n40263 , n40275 );
and ( n40277 , n19513 , RI15b63bb8_1268);
nor ( n40278 , n40276 , n40277 );
nand ( n40279 , n40252 , n40262 , n40278 );
or ( n40280 , n22775 , n386792 );
not ( n40281 , n19644 );
and ( n40282 , n40236 , RI15b62c40_1235);
and ( n40283 , n383476 , RI15b62cb8_1236);
nor ( n40284 , n40282 , n40283 );
or ( n40285 , n40281 , n40284 );
nand ( n40286 , n40280 , n40285 );
nor ( n40287 , n40279 , n40286 );
nand ( n40288 , n40237 , n40287 );
buf ( n40289 , n40288 );
buf ( n40290 , n382065 );
not ( n40291 , n32680 );
not ( n40292 , n382912 );
or ( n40293 , n40291 , n40292 );
and ( n40294 , n382931 , n35222 );
or ( n40295 , n32692 , n19066 );
not ( n40296 , n35162 );
or ( n40297 , n40296 , n32699 );
or ( n40298 , n32690 , n382967 );
nand ( n40299 , n40295 , n40297 , n40298 );
nor ( n40300 , n40294 , n40299 );
nand ( n40301 , n40293 , n40300 );
buf ( n40302 , n40301 );
buf ( n40303 , n380203 );
or ( n40304 , n379396 , RI15b54258_736);
not ( n40305 , n379340 );
and ( n40306 , n35244 , n40305 );
not ( n40307 , RI15b3fa38_36);
not ( n40308 , n35233 );
or ( n40309 , n40307 , n40308 );
and ( n40310 , RI15b3f9c0_35 , RI15b54780_747 , RI15b547f8_748);
nor ( n40311 , n40310 , n37566 );
nand ( n40312 , n40309 , n40311 );
nor ( n40313 , n35236 , RI15b547f8_748);
nor ( n40314 , n40306 , n40312 , n40313 );
nand ( n40315 , n40304 , n40314 );
buf ( n40316 , n40315 );
buf ( n40317 , n384996 );
buf ( n40318 , n381006 );
buf ( n40319 , n379895 );
or ( n40320 , n386588 , n380747 );
and ( n40321 , n386600 , n380745 );
or ( n40322 , n380776 , n19153 );
or ( n40323 , n386618 , n380785 );
or ( n40324 , n380768 , n386627 );
nand ( n40325 , n40322 , n40323 , n40324 );
nor ( n40326 , n40321 , n40325 );
nand ( n40327 , n40320 , n40326 );
buf ( n40328 , n40327 );
not ( n40329 , n22598 );
not ( n40330 , n379949 );
or ( n40331 , n40329 , n40330 );
not ( n40332 , n379949 );
nand ( n40333 , RI15b563a0_807 , RI15b56418_808);
nor ( n40334 , n379980 , n40333 );
nand ( n40335 , n40334 , RI15b56490_809);
not ( n40336 , n40335 );
or ( n40337 , n40332 , n40336 );
nand ( n40338 , n40337 , n380001 );
nor ( n40339 , n379948 , RI15b56508_810);
nor ( n40340 , n40338 , n40339 );
nand ( n40341 , n40331 , n40340 );
nor ( n40342 , n379948 , RI15b565f8_812);
nor ( n40343 , n40341 , n40342 );
or ( n40344 , n40343 , n18084 );
not ( n40345 , n40335 );
not ( n40346 , n40345 );
nand ( n40347 , n379949 , RI15b56508_810);
nor ( n40348 , n40346 , n40347 );
not ( n40349 , RI15b565f8_812);
nor ( n40350 , n40349 , n22598 , RI15b56670_813);
nand ( n40351 , n40348 , n40350 );
nand ( n40352 , n40344 , n40351 );
buf ( n40353 , n40352 );
buf ( n40354 , RI15b5dab0_1061);
buf ( n40355 , n382537 );
buf ( n40356 , n18226 );
buf ( n40357 , n22740 );
buf ( n40358 , n22343 );
buf ( n40359 , n381081 );
not ( n40360 , n40099 );
nand ( n40361 , n40360 , n386179 );
not ( n40362 , n386222 );
and ( n40363 , n40361 , n40362 );
not ( n40364 , n40361 );
and ( n40365 , n40364 , n386222 );
nor ( n40366 , n40363 , n40365 );
not ( n40367 , n386265 );
and ( n40368 , n40366 , n40367 );
not ( n40369 , n385877 );
nand ( n40370 , n40369 , n40106 );
not ( n40371 , n40370 );
not ( n40372 , n40371 );
not ( n40373 , n385870 );
and ( n40374 , n40372 , n40373 );
and ( n40375 , n40371 , n385870 );
nor ( n40376 , n40374 , n40375 );
not ( n40377 , n386019 );
or ( n40378 , n40376 , n40377 );
not ( n40379 , n386457 );
not ( n40380 , n386456 );
not ( n40381 , n40380 );
nand ( n40382 , n40381 , n386447 );
nand ( n40383 , n40379 , n40382 );
and ( n40384 , n40383 , n386500 );
and ( n40385 , n39987 , RI15b4bb58_448);
nor ( n40386 , n40384 , n40385 );
nand ( n40387 , n40378 , n40386 );
nor ( n40388 , n40368 , n40387 );
buf ( n40389 , n386514 );
not ( n40390 , n40389 );
not ( n40391 , n40390 );
not ( n40392 , n40380 );
and ( n40393 , n40391 , n40392 );
or ( n40394 , n386541 , n385860 );
or ( n40395 , n385870 , n386550 );
or ( n40396 , n40362 , n386557 );
nand ( n40397 , n40394 , n40395 , n40396 );
nor ( n40398 , n40393 , n40397 );
nand ( n40399 , n40388 , n40398 );
buf ( n40400 , n40399 );
buf ( n40401 , n384218 );
not ( n40402 , n21892 );
nor ( n40403 , n21886 , n40402 );
and ( n40404 , n33292 , n40403 );
buf ( n40405 , n21939 );
or ( n40406 , n21922 , n40405 );
nand ( n40407 , n40406 , n21946 );
and ( n40408 , n40407 , RI15b57c78_860);
not ( n40409 , n21968 );
not ( n40410 , n21949 );
or ( n40411 , n40409 , n40410 );
nand ( n40412 , n40411 , n21979 );
and ( n40413 , n40412 , RI15b55e78_796);
nor ( n40414 , n40408 , n40413 );
or ( n40415 , n40414 , n18078 );
and ( n40416 , n18188 , n40405 , n21940 );
or ( n40417 , n22601 , n21968 , RI15b55e78_796);
and ( n40418 , n18177 , RI15b57c78_860);
and ( n40419 , n18219 , RI15b56d78_828);
nor ( n40420 , n40418 , n40419 , n21751 );
nand ( n40421 , n40417 , n40420 );
nor ( n40422 , n40416 , n40421 );
nand ( n40423 , n40415 , n40422 );
nor ( n40424 , n40404 , n40423 );
not ( n40425 , n17507 );
not ( n40426 , n21886 );
or ( n40427 , n40425 , n40426 );
nand ( n40428 , n40427 , n17565 );
nand ( n40429 , n40428 , n40402 );
nand ( n40430 , n40424 , n40429 );
buf ( n40431 , n40430 );
buf ( n40432 , n22007 );
buf ( n40433 , n19651 );
buf ( n40434 , n381745 );
and ( n40435 , n40434 , n381752 );
not ( n40436 , n40434 );
not ( n40437 , n381752 );
and ( n40438 , n40436 , n40437 );
nor ( n40439 , n40435 , n40438 );
not ( n40440 , n385148 );
and ( n40441 , n40439 , n40440 );
nor ( n40442 , n21750 , n22836 );
nor ( n40443 , n40441 , n40442 );
not ( n40444 , n381775 );
not ( n40445 , n381778 );
and ( n40446 , n40444 , n40445 );
not ( n40447 , n40444 );
and ( n40448 , n40447 , n381778 );
nor ( n40449 , n40446 , n40448 );
nand ( n40450 , n40449 , n36162 );
nor ( n40451 , n381805 , n381810 );
not ( n40452 , n40451 );
nand ( n40453 , n40452 , n381811 );
nand ( n40454 , n40453 , n385134 );
and ( n40455 , n40443 , n40450 , n40454 );
and ( n40456 , n22529 , n33324 );
not ( n40457 , n22704 );
or ( n40458 , n40457 , n17516 );
nand ( n40459 , n40458 , n21790 );
and ( n40460 , n40459 , RI15b57228_838);
and ( n40461 , n17516 , n22525 );
and ( n40462 , n21795 , n40461 );
nor ( n40463 , n40456 , n40460 , n40462 );
nand ( n40464 , n40455 , n40463 );
buf ( n40465 , n40464 );
buf ( n40466 , n381081 );
buf ( n40467 , n33382 );
or ( n40468 , n384703 , n383865 );
or ( n40469 , n386705 , n40468 );
and ( n40470 , n383871 , n35478 );
and ( n40471 , n386716 , n40470 );
not ( n40472 , n40470 );
and ( n40473 , n40472 , n40468 , n33119 );
nor ( n40474 , n40473 , n21764 );
nor ( n40475 , n383885 , n383832 );
or ( n40476 , n40474 , n40475 );
nand ( n40477 , n40476 , n18154 );
nand ( n40478 , n383819 , n383892 );
nand ( n40479 , n40477 , n40478 );
and ( n40480 , n40479 , n383901 );
not ( n40481 , RI15b4fd70_589);
or ( n40482 , n40480 , n40481 );
not ( n40483 , n40478 );
nor ( n40484 , n40475 , n40483 );
or ( n40485 , n40474 , n40484 );
or ( n40486 , n386732 , n40485 );
or ( n40487 , n40478 , n386738 );
nand ( n40488 , n40482 , n40486 , n40487 );
nor ( n40489 , n40471 , n40488 );
nand ( n40490 , n40469 , n40489 );
buf ( n40491 , n40490 );
not ( n40492 , RI15b5f130_1109);
not ( n40493 , n384918 );
or ( n40494 , n40492 , n40493 );
and ( n40495 , n32275 , RI15b60e40_1171);
and ( n40496 , n384906 , n37641 );
nor ( n40497 , n40495 , n40496 );
nand ( n40498 , n40494 , n40497 );
buf ( n40499 , n40498 );
buf ( n40500 , n381872 );
buf ( n40501 , n33250 );
buf ( n40502 , n33250 );
nand ( n40503 , n40144 , n31766 , n19600 );
or ( n40504 , n40503 , n19513 );
nand ( n40505 , n40504 , RI15b608a0_1159);
nand ( n40506 , n40505 , n19590 );
buf ( n40507 , n40506 );
or ( n40508 , n31149 , n33111 );
and ( n40509 , n31161 , n33117 );
not ( n40510 , RI15b4e600_539);
or ( n40511 , n33128 , n40510 );
or ( n40512 , n31179 , n33134 );
or ( n40513 , n33126 , n31184 );
nand ( n40514 , n40511 , n40512 , n40513 );
nor ( n40515 , n40509 , n40514 );
nand ( n40516 , n40508 , n40515 );
buf ( n40517 , n40516 );
buf ( n40518 , n382065 );
not ( n40519 , n383845 );
not ( n40520 , n40519 );
not ( n40521 , n384726 );
or ( n40522 , n40520 , n40521 );
and ( n40523 , n35477 , n383878 );
or ( n40524 , n383903 , n17774 );
not ( n40525 , n384753 );
or ( n40526 , n40525 , n383911 );
or ( n40527 , n383895 , n384759 );
nand ( n40528 , n40524 , n40526 , n40527 );
nor ( n40529 , n40523 , n40528 );
nand ( n40530 , n40522 , n40529 );
buf ( n40531 , n40530 );
buf ( n40532 , n31719 );
buf ( n40533 , n380906 );
and ( n40534 , n383505 , n383522 );
nor ( n40535 , n40534 , n383577 );
or ( n40536 , n40535 , n383529 );
and ( n40537 , n383601 , RI15b5fb08_1130);
and ( n40538 , n383603 , n384936 );
and ( n40539 , n383607 , RI15b5f388_1114);
nor ( n40540 , n40537 , n40538 , n40539 );
nand ( n40541 , n40536 , n40540 );
buf ( n40542 , n40541 );
buf ( n40543 , n380940 );
buf ( n40544 , n36152 );
nor ( n40545 , n40544 , n21646 );
not ( n40546 , n40545 );
and ( n40547 , n36152 , n21646 );
not ( n40548 , n40547 );
nand ( n40549 , n40546 , n40548 );
nand ( n40550 , n40549 , n21748 );
not ( n40551 , n20708 );
buf ( n40552 , n21303 );
not ( n40553 , n40552 );
or ( n40554 , n40551 , n40553 );
or ( n40555 , n40552 , n20708 );
nand ( n40556 , n40554 , n40555 );
not ( n40557 , n21359 );
and ( n40558 , n40556 , n40557 );
not ( n40559 , RI15b57de0_863);
not ( n40560 , n21751 );
or ( n40561 , n40559 , n40560 );
not ( n40562 , n21516 );
and ( n40563 , n40562 , n21520 );
not ( n40564 , n40562 );
and ( n40565 , n40564 , n21521 );
nor ( n40566 , n40563 , n40565 );
not ( n40567 , n21562 );
nand ( n40568 , n40566 , n40567 );
nand ( n40569 , n40561 , n40568 );
nor ( n40570 , n40558 , n40569 );
nand ( n40571 , n40550 , n40570 );
not ( n40572 , n40571 );
and ( n40573 , n385164 , RI15b50748_610);
or ( n40574 , n36474 , n21646 );
or ( n40575 , n20708 , n385170 );
or ( n40576 , n21520 , n385178 );
nand ( n40577 , n40574 , n40575 , n40576 );
nor ( n40578 , n40573 , n40577 );
nand ( n40579 , n40572 , n40578 );
buf ( n40580 , n40579 );
buf ( n40581 , n382071 );
not ( n40582 , RI15b5e758_1088);
not ( n40583 , n379795 );
or ( n40584 , n40582 , n40583 );
or ( n40585 , n385188 , RI15b607b0_1157);
nand ( n40586 , n40584 , n40585 );
buf ( n40587 , n40586 );
buf ( n40588 , n20665 );
buf ( n40589 , n22007 );
or ( n40590 , n31006 , n31151 );
and ( n40591 , n31016 , n31164 );
or ( n40592 , n31175 , n17702 );
not ( n40593 , n31021 );
or ( n40594 , n40593 , n31182 );
or ( n40595 , n31173 , n31024 );
nand ( n40596 , n40592 , n40594 , n40595 );
nor ( n40597 , n40591 , n40596 );
nand ( n40598 , n40590 , n40597 );
buf ( n40599 , n40598 );
buf ( n40600 , n384218 );
buf ( n40601 , n31979 );
buf ( n40602 , n37799 );
not ( n40603 , n40602 );
or ( n40604 , n31053 , n40603 );
not ( n40605 , n384786 );
nand ( n40606 , n384907 , n40605 );
and ( n40607 , n31092 , RI15b61368_1182);
and ( n40608 , n383945 , RI15b58a10_889);
and ( n40609 , n383949 , RI15b5a810_953);
nor ( n40610 , n40608 , n40609 );
and ( n40611 , n383955 , RI15b5af90_969);
and ( n40612 , n383960 , RI15b5abd0_961);
nor ( n40613 , n40611 , n40612 );
and ( n40614 , n383965 , RI15b5b350_977);
and ( n40615 , n383970 , RI15b5a090_937);
and ( n40616 , n383972 , RI15b5a450_945);
nor ( n40617 , n40615 , n40616 );
and ( n40618 , n383975 , RI15b59910_921);
and ( n40619 , n383977 , RI15b59cd0_929);
nor ( n40620 , n40618 , n40619 );
and ( n40621 , n383982 , RI15b5be90_1001);
and ( n40622 , n383984 , RI15b5bad0_993);
nor ( n40623 , n40621 , n40622 );
and ( n40624 , n383987 , RI15b5c250_1009);
and ( n40625 , n383989 , RI15b5b710_985);
nor ( n40626 , n40624 , n40625 );
nand ( n40627 , n40617 , n40620 , n40623 , n40626 );
and ( n40628 , n383968 , n40627 );
and ( n40629 , n383994 , RI15b58dd0_897);
nor ( n40630 , n40614 , n40628 , n40629 );
and ( n40631 , n383997 , RI15b59190_905);
and ( n40632 , n383999 , RI15b59550_913);
nor ( n40633 , n40631 , n40632 );
nand ( n40634 , n40610 , n40613 , n40630 , n40633 );
and ( n40635 , n40634 , n31125 );
not ( n40636 , n36540 );
nor ( n40637 , n31076 , RI15b61368_1182);
and ( n40638 , n40636 , n40637 );
nor ( n40639 , n40607 , n40635 , n40638 );
nand ( n40640 , n40604 , n40606 , n40639 );
buf ( n40641 , n40640 );
not ( n40642 , n33924 );
or ( n40643 , n40642 , n34278 );
nand ( n40644 , n40643 , n33764 );
not ( n40645 , n40644 );
not ( n40646 , RI15b63c30_1269);
not ( n40647 , n379589 );
or ( n40648 , n40646 , n40647 );
or ( n40649 , n33928 , n34279 );
nand ( n40650 , n40648 , n40649 );
buf ( n40651 , n34273 );
nand ( n40652 , n40650 , n40651 );
not ( n40653 , n40652 );
or ( n40654 , n40645 , n40653 );
or ( n40655 , n40652 , n40644 );
nand ( n40656 , n40654 , n40655 );
nand ( n40657 , n40656 , n379785 );
buf ( n40658 , n34311 );
buf ( n40659 , n39184 );
not ( n40660 , n40659 );
and ( n40661 , n40658 , n40660 );
not ( n40662 , n40658 );
and ( n40663 , n40662 , n40659 );
nor ( n40664 , n40661 , n40663 );
and ( n40665 , n40664 , n379780 );
not ( n40666 , RI15b5db28_1062);
not ( n40667 , n379796 );
or ( n40668 , n40666 , n40667 );
or ( n40669 , n36518 , n379492 );
nand ( n40670 , n40668 , n40669 );
nor ( n40671 , n40665 , n40670 );
nand ( n40672 , n40657 , n40671 );
buf ( n40673 , n40672 );
nand ( n40674 , n31667 , n379341 );
and ( n40675 , n40674 , RI15b544b0_741);
and ( n40676 , n37569 , RI15b51378_636);
nor ( n40677 , n40675 , n40676 );
not ( n40678 , n40677 );
buf ( n40679 , n40678 );
buf ( n40680 , n385197 );
buf ( n40681 , n383174 );
buf ( n40682 , n380903 );
or ( n40683 , n31793 , n384502 );
not ( n40684 , n384378 );
nand ( n40685 , n384372 , n384377 );
nand ( n40686 , n40684 , n40685 );
not ( n40687 , n22750 );
nand ( n40688 , n40686 , n40687 );
not ( n40689 , n384479 );
not ( n40690 , n40689 );
not ( n40691 , n384475 );
or ( n40692 , n40690 , n40691 );
or ( n40693 , n384475 , n40689 );
nand ( n40694 , n40692 , n40693 );
nand ( n40695 , n40694 , n37599 );
not ( n40696 , n19512 );
not ( n40697 , n379711 );
and ( n40698 , n40696 , n40697 );
not ( n40699 , n384502 );
not ( n40700 , n384597 );
or ( n40701 , n40699 , n40700 );
or ( n40702 , n384597 , n384502 );
nand ( n40703 , n40701 , n40702 );
and ( n40704 , n40703 , n380811 );
nor ( n40705 , n40698 , n40704 );
nand ( n40706 , n40688 , n40695 , n40705 );
not ( n40707 , n40706 );
and ( n40708 , n31770 , RI15b5ce80_1035);
and ( n40709 , n37610 , n384377 );
and ( n40710 , n31778 , n40689 );
nor ( n40711 , n40708 , n40709 , n40710 );
nand ( n40712 , n40683 , n40707 , n40711 );
buf ( n40713 , n40712 );
buf ( n40714 , n382049 );
buf ( n40715 , n39639 );
not ( n40716 , n39641 );
xor ( n40717 , n40715 , n40716 );
not ( n40718 , n31601 );
or ( n40719 , n40717 , n40718 );
not ( n40720 , n379391 );
not ( n40721 , n39666 );
not ( n40722 , n40721 );
or ( n40723 , n40720 , n40722 );
nand ( n40724 , n40723 , n31700 );
and ( n40725 , n40724 , n31676 );
or ( n40726 , n40721 , n31709 , n31676 );
and ( n40727 , n379394 , RI15b58218_872);
and ( n40728 , n31712 , RI15b52020_663);
nor ( n40729 , n40727 , n40728 );
nand ( n40730 , n40726 , n40729 );
nor ( n40731 , n40725 , n40730 );
nand ( n40732 , n40719 , n40731 );
buf ( n40733 , n40732 );
buf ( n40734 , n386760 );
buf ( n40735 , n382052 );
buf ( n40736 , n380906 );
buf ( n40737 , n384996 );
not ( n40738 , n385961 );
not ( n40739 , n40738 );
not ( n40740 , n385970 );
and ( n40741 , n40739 , n40740 );
and ( n40742 , n40738 , n385970 );
nor ( n40743 , n40741 , n40742 );
nor ( n40744 , n40743 , n40377 );
not ( n40745 , n386236 );
not ( n40746 , n40745 );
not ( n40747 , n386240 );
and ( n40748 , n40746 , n40747 );
and ( n40749 , n40745 , n386240 );
nor ( n40750 , n40748 , n40749 );
not ( n40751 , n386263 );
not ( n40752 , n40751 );
or ( n40753 , n40750 , n40752 );
not ( n40754 , n386492 );
buf ( n40755 , n386488 );
nand ( n40756 , n40755 , n386491 );
nand ( n40757 , n40754 , n40756 );
and ( n40758 , n40757 , n386500 );
buf ( n40759 , n34782 );
nor ( n40760 , n40759 , n387178 );
nor ( n40761 , n40758 , n40760 );
nand ( n40762 , n40753 , n40761 );
nor ( n40763 , n40744 , n40762 );
not ( n40764 , n386516 );
and ( n40765 , n40764 , n386491 );
or ( n40766 , n386541 , n385974 );
or ( n40767 , n385970 , n386550 );
or ( n40768 , n386557 , n386240 );
nand ( n40769 , n40766 , n40767 , n40768 );
nor ( n40770 , n40765 , n40769 );
nand ( n40771 , n40763 , n40770 );
buf ( n40772 , n40771 );
buf ( n40773 , n37727 );
buf ( n40774 , n33582 );
not ( n40775 , n40774 );
nor ( n40776 , n40773 , n40775 );
or ( n40777 , n40776 , n33585 );
buf ( n40778 , n37770 );
not ( n40779 , n40778 );
nand ( n40780 , n40777 , n40779 );
not ( n40781 , n33588 );
nand ( n40782 , n40778 , n40773 , n40781 );
and ( n40783 , n383601 , RI15b604e0_1151);
and ( n40784 , n383607 , RI15b5eed8_1104);
nor ( n40785 , n40783 , n40784 );
nand ( n40786 , n40780 , n40782 , n40785 );
buf ( n40787 , n40786 );
buf ( n40788 , n22714 );
or ( n40789 , n31149 , n33597 );
and ( n40790 , n31161 , n33600 );
not ( n40791 , RI15b4e9c0_547);
or ( n40792 , n33609 , n40791 );
or ( n40793 , n32452 , n33615 );
or ( n40794 , n33607 , n31184 );
nand ( n40795 , n40792 , n40793 , n40794 );
nor ( n40796 , n40790 , n40795 );
nand ( n40797 , n40789 , n40796 );
buf ( n40798 , n40797 );
buf ( n40799 , n380942 );
buf ( n40800 , n385195 );
buf ( n40801 , n39168 );
nand ( n40802 , n40801 , n379785 );
not ( n40803 , n40802 );
not ( n40804 , n36496 );
or ( n40805 , n40803 , n40804 );
not ( n40806 , n39169 );
buf ( n40807 , n40806 );
nand ( n40808 , n40805 , n40807 );
not ( n40809 , n36501 );
nor ( n40810 , n40801 , n40806 );
nand ( n40811 , n40809 , n40810 );
buf ( n40812 , n39192 );
not ( n40813 , n40812 );
and ( n40814 , n40813 , n34460 );
not ( n40815 , n40813 );
and ( n40816 , n40815 , n39193 );
nor ( n40817 , n40814 , n40816 );
and ( n40818 , n40817 , n36513 );
not ( n40819 , RI15b5dd80_1067);
not ( n40820 , n34651 );
or ( n40821 , n40819 , n40820 );
or ( n40822 , n36518 , n379573 );
nand ( n40823 , n40821 , n40822 );
nor ( n40824 , n40818 , n40823 );
nand ( n40825 , n40808 , n40811 , n40824 );
buf ( n40826 , n40825 );
not ( n40827 , RI15b4c0f8_460);
and ( n40828 , n37698 , n20731 );
not ( n40829 , n39844 );
not ( n40830 , n18145 );
and ( n40831 , n40829 , n40830 , n18126 );
nor ( n40832 , n40831 , n20731 );
nor ( n40833 , n40828 , n40832 );
not ( n40834 , n40833 );
or ( n40835 , n40827 , n40834 );
nand ( n40836 , n40835 , n18062 );
not ( n40837 , n39845 );
and ( n40838 , n40837 , RI15b50ec8_626);
or ( n40839 , n32367 , RI15b50ec8_626);
nand ( n40840 , n37698 , n385101 );
nand ( n40841 , n40839 , n40840 );
nor ( n40842 , n40838 , n40841 );
and ( n40843 , n40836 , n40842 );
not ( n40844 , n383888 );
and ( n40845 , n40833 , n40844 );
nor ( n40846 , n40843 , n40845 );
not ( n40847 , n39848 );
and ( n40848 , n40847 , RI15b4c1e8_462);
not ( n40849 , n40847 );
and ( n40850 , n40849 , n17998 );
nor ( n40851 , n40848 , n40850 );
or ( n40852 , n40846 , n40851 );
nand ( n40853 , n40847 , n384178 );
not ( n40854 , n381467 );
nand ( n40855 , n40854 , n18214 );
nor ( n40856 , n17622 , RI15b50f40_627);
or ( n40857 , n40837 , n40856 );
nand ( n40858 , n40857 , RI15b50fb8_628);
or ( n40859 , n32366 , n381633 );
not ( n40860 , n40856 );
not ( n40861 , RI15b50fb8_628);
nand ( n40862 , n40860 , n39832 , n40861 );
nand ( n40863 , n40855 , n40858 , n40859 , n40862 );
nand ( n40864 , n40863 , n17998 , n384177 );
nand ( n40865 , n40853 , n40864 , n384179 );
nand ( n40866 , n40852 , n40865 );
not ( n40867 , n384178 );
not ( n40868 , n40867 );
not ( n40869 , n39848 );
or ( n40870 , n40868 , n40869 );
nand ( n40871 , n40870 , n40863 );
and ( n40872 , n382548 , RI15b510a8_630);
or ( n40873 , n40830 , n21977 );
or ( n40874 , n21350 , n18130 );
nand ( n40875 , n40873 , n40874 , n37701 );
nor ( n40876 , n40872 , n40875 );
not ( n40877 , n18139 );
and ( n40878 , n18182 , n40877 , n39216 );
nor ( n40879 , n40878 , n382550 );
and ( n40880 , n40871 , n40876 , n40879 );
nand ( n40881 , n40866 , n40880 );
nand ( n40882 , n40881 , n18077 );
buf ( n40883 , n381475 );
nand ( n40884 , n379984 , n18141 );
or ( n40885 , n40884 , n18099 );
nand ( n40886 , n40885 , n18077 );
nand ( n40887 , n40883 , n40886 );
and ( n40888 , n383147 , n18072 );
and ( n40889 , n18164 , n18165 );
nor ( n40890 , n40889 , n18072 );
nor ( n40891 , n40888 , n40890 , n383898 );
not ( n40892 , n32998 );
nand ( n40893 , n40891 , n40892 , n21750 );
nor ( n40894 , n40887 , n40893 );
nand ( n40895 , n40882 , n40894 );
buf ( n40896 , n40895 );
buf ( n40897 , n383498 );
buf ( n40898 , n383345 );
not ( n40899 , RI15b55a40_787);
not ( n40900 , n380000 );
or ( n40901 , n40899 , n40900 );
and ( n40902 , n36384 , RI15b4c5a8_470);
not ( n40903 , RI15b55a40_787);
not ( n40904 , n379954 );
not ( n40905 , n40904 );
or ( n40906 , n40903 , n40905 );
or ( n40907 , n40904 , RI15b55a40_787);
nand ( n40908 , n40906 , n40907 );
and ( n40909 , n379949 , n40908 );
nor ( n40910 , n40902 , n40909 );
nand ( n40911 , n40901 , n40910 );
buf ( n40912 , n40911 );
not ( n40913 , n36395 );
not ( n40914 , n382912 );
or ( n40915 , n40913 , n40914 );
and ( n40916 , n382931 , n36401 );
or ( n40917 , n36410 , n19081 );
or ( n40918 , n35805 , n36416 );
or ( n40919 , n36408 , n382967 );
nand ( n40920 , n40917 , n40918 , n40919 );
nor ( n40921 , n40916 , n40920 );
nand ( n40922 , n40915 , n40921 );
buf ( n40923 , n40922 );
buf ( n40924 , n22005 );
buf ( n40925 , n385112 );
buf ( n40926 , n381004 );
not ( n40927 , n19201 );
nand ( n40928 , n19533 , n19497 );
not ( n40929 , n40928 );
nor ( n40930 , n19558 , n19533 );
nor ( n40931 , n40929 , n40930 );
buf ( n40932 , n18281 );
or ( n40933 , n40931 , n40932 );
or ( n40934 , n32385 , RI15b5d330_1045);
nand ( n40935 , n19533 , n19496 );
and ( n40936 , n31754 , n40935 );
nand ( n40937 , n40936 , n31759 , n19148 );
nand ( n40938 , n40937 , RI15b5d330_1045);
nand ( n40939 , n40933 , n40934 , n40938 );
not ( n40940 , n40939 );
or ( n40941 , n40927 , n40940 );
nand ( n40942 , n35680 , n39115 );
nand ( n40943 , n31766 , n380773 , n19598 , n40942 );
not ( n40944 , n40943 );
or ( n40945 , n40944 , n18302 );
not ( n40946 , n19331 );
not ( n40947 , RI15b5d240_1043);
and ( n40948 , n40946 , n40947 );
and ( n40949 , n19293 , RI15b5d240_1043);
nor ( n40950 , n40948 , n40949 );
not ( n40951 , n35681 );
or ( n40952 , n40950 , n40951 );
buf ( n40953 , n40932 );
or ( n40954 , n40953 , n380788 );
nand ( n40955 , n40945 , n40952 , n40954 );
not ( n40956 , n40955 );
nand ( n40957 , n40941 , n40956 );
buf ( n40958 , n40957 );
buf ( n40959 , n382537 );
buf ( n40960 , n385195 );
buf ( n40961 , n31640 );
nand ( n40962 , n40961 , n379374 );
nor ( n40963 , n40962 , n31644 );
and ( n40964 , n40963 , n31304 );
nand ( n40965 , n40964 , n379168 );
nor ( n40966 , n40965 , n31201 );
not ( n40967 , n40966 );
nor ( n40968 , n40967 , n31667 );
or ( n40969 , n40968 , n31699 );
nand ( n40970 , n40969 , n379192 );
not ( n40971 , n31706 );
buf ( n40972 , n40971 );
nor ( n40973 , n40972 , n379192 );
and ( n40974 , n40967 , n40973 );
not ( n40975 , n31549 );
not ( n40976 , n31543 );
not ( n40977 , n40976 );
or ( n40978 , n40975 , n40977 );
or ( n40979 , n40976 , n31549 );
nand ( n40980 , n40978 , n40979 );
not ( n40981 , n40980 );
not ( n40982 , n31599 );
or ( n40983 , n40981 , n40982 );
and ( n40984 , n379394 , RI15b57d68_862);
and ( n40985 , n31712 , RI15b51b70_653);
nor ( n40986 , n40984 , n40985 );
nand ( n40987 , n40983 , n40986 );
nor ( n40988 , n40974 , n40987 );
nand ( n40989 , n40970 , n40988 );
buf ( n40990 , n40989 );
buf ( n40991 , n32160 );
buf ( n40992 , n21800 );
buf ( n40993 , n381707 );
buf ( n40994 , n384218 );
nor ( n40995 , n34994 , n35108 );
nand ( n40996 , n40995 , n35098 );
nor ( n40997 , n40996 , n35087 );
and ( n40998 , n40997 , n35077 );
nand ( n40999 , n40998 , n35103 );
not ( n41000 , n34957 );
nor ( n41001 , n40999 , n41000 );
not ( n41002 , n41001 );
not ( n41003 , n34947 );
not ( n41004 , n35011 );
and ( n41005 , n41003 , n41004 );
not ( n41006 , n41003 );
and ( n41007 , n41006 , n35011 );
nor ( n41008 , n41005 , n41007 );
not ( n41009 , n41008 );
and ( n41010 , n41002 , n41009 );
not ( n41011 , n41002 );
and ( n41012 , n41011 , n41008 );
nor ( n41013 , n41010 , n41012 );
not ( n41014 , n41013 );
not ( n41015 , n379825 );
or ( n41016 , n41014 , n41015 );
buf ( n41017 , n379832 );
nand ( n41018 , n41017 , RI15b463b0_261);
and ( n41019 , n35459 , n22245 );
and ( n41020 , n35461 , RI15b65b98_1336);
nor ( n41021 , n41019 , n41020 );
nand ( n41022 , n41016 , n41018 , n41021 );
buf ( n41023 , n41022 );
buf ( n41024 , n379893 );
buf ( n41025 , n384996 );
nand ( n41026 , n41001 , n41008 );
buf ( n41027 , n41026 );
not ( n41028 , n41027 );
not ( n41029 , n41015 );
and ( n41030 , n41028 , n41029 );
not ( n41031 , n41015 );
nand ( n41032 , n41031 , n35113 );
not ( n41033 , n41032 );
nor ( n41034 , n41030 , n41033 );
or ( n41035 , n41034 , n35067 );
or ( n41036 , n35113 , n41015 );
not ( n41037 , n41036 );
nand ( n41038 , n41037 , n41027 , n35067 );
nand ( n41039 , n41017 , RI15b46428_262);
not ( n41040 , n382000 );
or ( n41041 , n22287 , n41040 );
or ( n41042 , n32143 , n382000 );
nand ( n41043 , n41041 , n41042 );
and ( n41044 , n35461 , n41043 );
and ( n41045 , n35459 , n41040 );
nor ( n41046 , n41044 , n41045 );
and ( n41047 , n41038 , n41039 , n41046 );
nand ( n41048 , n41035 , n41047 );
buf ( n41049 , n41048 );
buf ( n41050 , n382049 );
buf ( n41051 , n381021 );
buf ( n41052 , n22740 );
not ( n41053 , n383930 );
and ( n41054 , n383945 , RI15b58b00_891);
and ( n41055 , n383949 , RI15b5a900_955);
nor ( n41056 , n41054 , n41055 );
and ( n41057 , n383955 , RI15b5b080_971);
and ( n41058 , n383960 , RI15b5acc0_963);
nor ( n41059 , n41057 , n41058 );
and ( n41060 , n383965 , RI15b5b440_979);
and ( n41061 , n383970 , RI15b5a180_939);
and ( n41062 , n383977 , RI15b59dc0_931);
nor ( n41063 , n41061 , n41062 );
and ( n41064 , n383972 , RI15b5a540_947);
and ( n41065 , n383975 , RI15b59a00_923);
nor ( n41066 , n41064 , n41065 );
and ( n41067 , n383987 , RI15b5c340_1011);
and ( n41068 , n383989 , RI15b5b800_987);
nor ( n41069 , n41067 , n41068 );
and ( n41070 , n383982 , RI15b5bf80_1003);
and ( n41071 , n383984 , RI15b5bbc0_995);
nor ( n41072 , n41070 , n41071 );
nand ( n41073 , n41063 , n41066 , n41069 , n41072 );
and ( n41074 , n383967 , n41073 );
and ( n41075 , n383994 , RI15b58ec0_899);
nor ( n41076 , n41060 , n41074 , n41075 );
and ( n41077 , n383997 , RI15b59280_907);
and ( n41078 , n383999 , RI15b59640_915);
nor ( n41079 , n41077 , n41078 );
nand ( n41080 , n41056 , n41059 , n41076 , n41079 );
not ( n41081 , n41080 );
or ( n41082 , n41053 , n41081 );
and ( n41083 , n384022 , RI15b62358_1216);
not ( n41084 , RI15b62358_1216);
not ( n41085 , n38476 );
not ( n41086 , n41085 );
or ( n41087 , n41084 , n41086 );
or ( n41088 , n41085 , RI15b62358_1216);
nand ( n41089 , n41087 , n41088 );
and ( n41090 , n384025 , n41089 );
nor ( n41091 , n41083 , n41090 );
nand ( n41092 , n41082 , n41091 );
buf ( n41093 , n41092 );
buf ( n41094 , n379847 );
buf ( n41095 , n382069 );
or ( n41096 , n383814 , n384057 );
and ( n41097 , n383857 , n384169 );
or ( n41098 , n384182 , n21148 );
not ( n41099 , n383907 );
or ( n41100 , n41099 , n384190 );
or ( n41101 , n384180 , n383917 );
nand ( n41102 , n41098 , n41100 , n41101 );
nor ( n41103 , n41097 , n41102 );
nand ( n41104 , n41096 , n41103 );
buf ( n41105 , n41104 );
buf ( n41106 , n22402 );
buf ( n41107 , n383345 );
not ( n41108 , n21837 );
nor ( n41109 , n41108 , n21846 );
and ( n41110 , n379855 , n41109 );
not ( n41111 , n21958 );
not ( n41112 , n21949 );
or ( n41113 , n41111 , n41112 );
nand ( n41114 , n41113 , n21979 );
and ( n41115 , n41114 , RI15b55ba8_790);
and ( n41116 , n18150 , RI15b579a8_854);
or ( n41117 , n21982 , n21958 , RI15b55ba8_790);
not ( n41118 , n21929 );
not ( n41119 , RI15b579a8_854);
and ( n41120 , n41118 , n41119 );
and ( n41121 , n21929 , RI15b579a8_854);
nor ( n41122 , n41120 , n41121 );
or ( n41123 , n21922 , n41122 );
nand ( n41124 , n41117 , n41123 );
nor ( n41125 , n41115 , n41116 , n41124 );
or ( n41126 , n41125 , n18078 );
and ( n41127 , n18177 , RI15b579a8_854);
and ( n41128 , n18219 , RI15b56aa8_822);
nor ( n41129 , n41127 , n41128 , n21751 );
nand ( n41130 , n41126 , n41129 );
nor ( n41131 , n41110 , n41130 );
not ( n41132 , n17507 );
not ( n41133 , n41108 );
or ( n41134 , n41132 , n41133 );
nand ( n41135 , n41134 , n17565 );
nand ( n41136 , n41135 , n21846 );
nand ( n41137 , n41131 , n41136 );
buf ( n41138 , n41137 );
buf ( n41139 , n381707 );
buf ( n41140 , n381707 );
not ( n41141 , n37924 );
and ( n41142 , n37918 , n41141 );
not ( n41143 , n37918 );
and ( n41144 , n41143 , n37924 );
nor ( n41145 , n41142 , n41144 );
nor ( n41146 , n41145 , n33630 );
and ( n41147 , n37962 , n37969 );
not ( n41148 , n37962 );
and ( n41149 , n41148 , n37968 );
nor ( n41150 , n41147 , n41149 );
nor ( n41151 , n41150 , n33640 );
not ( n41152 , n37952 );
not ( n41153 , n41152 );
not ( n41154 , n36687 );
or ( n41155 , n41153 , n41154 );
nand ( n41156 , n41155 , n37953 );
nand ( n41157 , n41156 , n36689 );
nand ( n41158 , n21751 , RI15b583f8_876);
nand ( n41159 , n41157 , n41158 );
nor ( n41160 , n41146 , n41151 , n41159 );
not ( n41161 , n22573 );
and ( n41162 , n41161 , n21771 );
and ( n41163 , n37992 , RI15b574f8_844);
not ( n41164 , n37997 );
nor ( n41165 , n41164 , RI15b574f8_844);
and ( n41166 , n37988 , n41165 );
nor ( n41167 , n41162 , n41163 , n41166 );
nand ( n41168 , n41160 , n41167 );
buf ( n41169 , n41168 );
buf ( n41170 , n36854 );
buf ( n41171 , n33382 );
nand ( n41172 , n384907 , n384848 );
not ( n41173 , n384913 );
nand ( n41174 , n41173 , n381614 );
nand ( n41175 , n384918 , RI15b5f298_1112);
nand ( n41176 , n37773 , RI15b60fa8_1174);
nand ( n41177 , n41172 , n41174 , n41175 , n41176 );
buf ( n41178 , n41177 );
or ( n41179 , n383814 , n40468 );
and ( n41180 , n383857 , n40470 );
or ( n41181 , n40480 , n21142 );
not ( n41182 , n383907 );
or ( n41183 , n41182 , n40485 );
or ( n41184 , n40478 , n383917 );
nand ( n41185 , n41181 , n41183 , n41184 );
nor ( n41186 , n41180 , n41185 );
nand ( n41187 , n41179 , n41186 );
buf ( n41188 , n41187 );
buf ( n41189 , n382071 );
buf ( n41190 , n380865 );
nand ( n41191 , n40966 , n379191 );
nor ( n41192 , n41191 , n31667 );
or ( n41193 , n41192 , n31699 );
nand ( n41194 , n41193 , n31648 );
not ( n41195 , n31706 );
nor ( n41196 , n41195 , n31648 );
and ( n41197 , n41191 , n41196 );
buf ( n41198 , n31550 );
not ( n41199 , n31557 );
and ( n41200 , n41198 , n41199 );
not ( n41201 , n41198 );
and ( n41202 , n41201 , n31557 );
nor ( n41203 , n41200 , n41202 );
or ( n41204 , n31600 , n41203 );
and ( n41205 , n379394 , RI15b57de0_863);
buf ( n41206 , n379398 );
and ( n41207 , n41206 , RI15b51be8_654);
nor ( n41208 , n41205 , n41207 );
nand ( n41209 , n41204 , n41208 );
nor ( n41210 , n41197 , n41209 );
nand ( n41211 , n41194 , n41210 );
buf ( n41212 , n41211 );
buf ( n41213 , n384203 );
and ( n41214 , n19559 , n40935 );
and ( n41215 , RI15b5d2b8_1044 , n41214 );
not ( n41216 , RI15b5d2b8_1044);
and ( n41217 , n41216 , n40931 );
nor ( n41218 , n41215 , n41217 );
not ( n41219 , n41218 );
or ( n41220 , n41219 , n19200 );
and ( n41221 , n40943 , RI15b5d2b8_1044);
and ( n41222 , n380789 , n18249 );
and ( n41223 , n35681 , n19336 );
nor ( n41224 , n41221 , n41222 , n41223 );
nand ( n41225 , n41220 , n41224 );
buf ( n41226 , n41225 );
buf ( n41227 , n381081 );
buf ( n41228 , n379802 );
buf ( n41229 , n31979 );
not ( n41230 , n39256 );
and ( n41231 , n41230 , RI15b44b50_209);
and ( n41232 , n381925 , n385300 );
nor ( n41233 , n41231 , n41232 );
nand ( n41234 , n36797 , n41233 );
buf ( n41235 , n41234 );
buf ( n41236 , n32160 );
buf ( n41237 , n20663 );
buf ( n41238 , n35651 );
buf ( n41239 , n381004 );
not ( n41240 , n385922 );
buf ( n41241 , n385914 );
not ( n41242 , n41241 );
or ( n41243 , n41240 , n41242 );
or ( n41244 , n41241 , n385922 );
nand ( n41245 , n41243 , n41244 );
and ( n41246 , n41245 , n34779 );
not ( n41247 , n386224 );
not ( n41248 , n41247 );
not ( n41249 , n386228 );
and ( n41250 , n41248 , n41249 );
and ( n41251 , n41247 , n386228 );
nor ( n41252 , n41250 , n41251 );
not ( n41253 , n386262 );
or ( n41254 , n41252 , n41253 );
not ( n41255 , n386300 );
not ( n41256 , n386474 );
not ( n41257 , n41256 );
or ( n41258 , n41255 , n41257 );
nand ( n41259 , n41258 , n38137 );
and ( n41260 , n41259 , n386500 );
not ( n41261 , RI15b4bcc0_451);
nor ( n41262 , n38209 , n41261 );
nor ( n41263 , n41260 , n41262 );
nand ( n41264 , n41254 , n41263 );
nor ( n41265 , n41246 , n41264 );
not ( n41266 , n40165 );
not ( n41267 , n41266 );
and ( n41268 , n41267 , n386300 );
or ( n41269 , n386541 , n385926 );
or ( n41270 , n385922 , n386550 );
or ( n41271 , n386228 , n386557 );
nand ( n41272 , n41269 , n41270 , n41271 );
nor ( n41273 , n41268 , n41272 );
nand ( n41274 , n41265 , n41273 );
buf ( n41275 , n41274 );
buf ( n41276 , n22716 );
and ( n41277 , n39950 , n39951 );
not ( n41278 , n39950 );
and ( n41279 , n41278 , n385795 );
nor ( n41280 , n41277 , n41279 );
and ( n41281 , n41280 , n386020 );
not ( n41282 , n40751 );
not ( n41283 , n386153 );
not ( n41284 , n39964 );
or ( n41285 , n41283 , n41284 );
or ( n41286 , n39964 , n386153 );
nand ( n41287 , n41285 , n41286 );
not ( n41288 , n41287 );
or ( n41289 , n41282 , n41288 );
not ( n41290 , n34731 );
not ( n41291 , n41290 );
not ( n41292 , n34730 );
not ( n41293 , n41292 );
not ( n41294 , n41293 );
not ( n41295 , n41294 );
or ( n41296 , n41291 , n41295 );
buf ( n41297 , n34732 );
nand ( n41298 , n41296 , n41297 );
and ( n41299 , n41298 , n386500 );
not ( n41300 , n38209 );
buf ( n41301 , n41300 );
buf ( n41302 , n41301 );
and ( n41303 , n41302 , RI15b4b720_439);
nor ( n41304 , n41299 , n41303 );
nand ( n41305 , n41289 , n41304 );
nor ( n41306 , n41281 , n41305 );
buf ( n41307 , n41266 );
buf ( n41308 , n41307 );
not ( n41309 , n41308 );
and ( n41310 , n41309 , n41290 );
or ( n41311 , n386541 , n385787 );
or ( n41312 , n39951 , n386550 );
or ( n41313 , n386153 , n386557 );
nand ( n41314 , n41311 , n41312 , n41313 );
nor ( n41315 , n41310 , n41314 );
nand ( n41316 , n41306 , n41315 );
buf ( n41317 , n41316 );
buf ( n41318 , n22740 );
buf ( n41319 , n22738 );
buf ( n41320 , n22343 );
buf ( n41321 , n18226 );
or ( n41322 , n36937 , n35472 );
and ( n41323 , n36946 , n35479 );
not ( n41324 , RI15b4dfe8_526);
or ( n41325 , n35488 , n41324 );
not ( n41326 , n38402 );
or ( n41327 , n41326 , n35497 );
or ( n41328 , n35486 , n36955 );
nand ( n41329 , n41325 , n41327 , n41328 );
nor ( n41330 , n41323 , n41329 );
nand ( n41331 , n41322 , n41330 );
buf ( n41332 , n41331 );
or ( n41333 , n31053 , n38307 );
not ( n41334 , n384832 );
nand ( n41335 , n384907 , n41334 );
not ( n41336 , n31127 );
or ( n41337 , n41336 , n31062 );
nand ( n41338 , n41337 , n31091 );
and ( n41339 , n41338 , RI15b60eb8_1172);
buf ( n41340 , n31081 );
not ( n41341 , n31062 );
or ( n41342 , n41340 , n41341 , RI15b60eb8_1172);
not ( n41343 , n36538 );
not ( n41344 , n40243 );
or ( n41345 , n41343 , n41344 );
nand ( n41346 , n41342 , n41345 );
nor ( n41347 , n41339 , n41346 );
nand ( n41348 , n41333 , n41335 , n41347 );
buf ( n41349 , n41348 );
buf ( n41350 , n22009 );
buf ( n41351 , n382067 );
buf ( n41352 , n33250 );
and ( n41353 , n40937 , RI15b5d3a8_1046);
or ( n41354 , n32385 , n383943 );
or ( n41355 , n383484 , n40928 );
nand ( n41356 , n40930 , n383484 );
nand ( n41357 , n41354 , n41355 , n41356 );
nor ( n41358 , n41353 , n41357 );
or ( n41359 , n41358 , n19200 );
and ( n41360 , n40943 , RI15b5d3a8_1046);
and ( n41361 , n380789 , n383485 );
or ( n41362 , n19331 , n40947 );
buf ( n41363 , n19303 );
or ( n41364 , n41363 , RI15b5d240_1043);
nand ( n41365 , n41362 , n41364 );
and ( n41366 , n35681 , n41365 );
nor ( n41367 , n41360 , n41361 , n41366 );
nand ( n41368 , n41359 , n41367 );
buf ( n41369 , n41368 );
buf ( n41370 , n35651 );
buf ( n41371 , n40965 );
nor ( n41372 , n41371 , n31667 );
or ( n41373 , n41372 , n31699 );
nand ( n41374 , n41373 , n31201 );
nor ( n41375 , n41195 , n31201 );
and ( n41376 , n41371 , n41375 );
not ( n41377 , n31542 );
buf ( n41378 , n31535 );
not ( n41379 , n41378 );
not ( n41380 , n41379 );
or ( n41381 , n41377 , n41380 );
or ( n41382 , n41379 , n31542 );
nand ( n41383 , n41381 , n41382 );
not ( n41384 , n41383 );
not ( n41385 , n31599 );
or ( n41386 , n41384 , n41385 );
and ( n41387 , n379394 , RI15b57cf0_861);
and ( n41388 , n41206 , RI15b51af8_652);
nor ( n41389 , n41387 , n41388 );
nand ( n41390 , n41386 , n41389 );
nor ( n41391 , n41376 , n41390 );
nand ( n41392 , n41374 , n41391 );
buf ( n41393 , n41392 );
buf ( n41394 , n380865 );
buf ( n41395 , n379895 );
buf ( n41396 , n379847 );
not ( n41397 , n33365 );
not ( n41398 , n32129 );
or ( n41399 , n41397 , n41398 );
and ( n41400 , n38869 , RI15b433e0_159);
or ( n41401 , n32141 , n32172 );
or ( n41402 , n32148 , n32187 );
or ( n41403 , n32181 , n32150 );
nand ( n41404 , n41401 , n41402 , n41403 );
nor ( n41405 , n41400 , n41404 );
nand ( n41406 , n41399 , n41405 );
buf ( n41407 , n41406 );
buf ( n41408 , n379844 );
buf ( n41409 , n32981 );
not ( n41410 , RI15b61818_1192);
or ( n41411 , n31091 , n41410 );
nor ( n41412 , n383584 , n31130 );
nand ( n41413 , n31075 , n41412 );
nor ( n41414 , n41413 , n32280 );
and ( n41415 , n41414 , RI15b614d0_1185);
nand ( n41416 , n41415 , RI15b61548_1186);
nor ( n41417 , n41416 , n32309 );
nand ( n41418 , n41417 , RI15b61638_1188);
not ( n41419 , n41418 );
nand ( n41420 , n41419 , RI15b616b0_1189);
nand ( n41421 , RI15b61728_1190 , RI15b617a0_1191);
nor ( n41422 , n41420 , n41421 );
not ( n41423 , n41422 );
and ( n41424 , n41423 , n41410 );
not ( n41425 , n41423 );
and ( n41426 , n41425 , RI15b61818_1192);
nor ( n41427 , n41424 , n41426 );
and ( n41428 , n41427 , n31082 );
or ( n41429 , n31052 , n380480 );
nand ( n41430 , n41429 , n37817 );
not ( n41431 , n35507 );
not ( n41432 , n38665 );
not ( n41433 , n38581 );
and ( n41434 , n41432 , n41433 );
and ( n41435 , n38665 , n38581 );
nor ( n41436 , n41434 , n41435 );
nor ( n41437 , n41431 , n41436 );
nor ( n41438 , n41428 , n41430 , n41437 );
nand ( n41439 , n41411 , n41438 );
buf ( n41440 , n41439 );
buf ( n41441 , n383498 );
buf ( n41442 , n20663 );
or ( n41443 , n31150 , n383886 );
or ( n41444 , n383814 , n41443 );
nand ( n41445 , n31162 , n21337 );
not ( n41446 , n41445 );
and ( n41447 , n383857 , n41446 );
and ( n41448 , n41445 , n41443 , n385009 );
nor ( n41449 , n41448 , n21764 );
nor ( n41450 , n31168 , n35629 );
or ( n41451 , n41449 , n41450 );
nand ( n41452 , n41451 , n18154 );
or ( n41453 , n383865 , n31172 );
and ( n41454 , n41452 , n41453 );
nor ( n41455 , n41454 , n383902 );
not ( n41456 , RI15b4d688_506);
or ( n41457 , n41455 , n41456 );
not ( n41458 , n383907 );
not ( n41459 , n41453 );
nor ( n41460 , n41450 , n41459 );
or ( n41461 , n41449 , n41460 );
or ( n41462 , n41458 , n41461 );
or ( n41463 , n41453 , n383917 );
nand ( n41464 , n41457 , n41462 , n41463 );
nor ( n41465 , n41447 , n41464 );
nand ( n41466 , n41444 , n41465 );
buf ( n41467 , n41466 );
buf ( n41468 , n33382 );
buf ( n41469 , RI15b47a30_309);
buf ( n41470 , n379895 );
buf ( n41471 , n31033 );
buf ( n41472 , n22655 );
buf ( n41473 , n22738 );
buf ( n41474 , n34738 );
buf ( n41475 , n34739 );
nor ( n41476 , n41474 , n41475 );
not ( n41477 , n41476 );
buf ( n41478 , n34740 );
nand ( n41479 , n41477 , n41478 );
nand ( n41480 , n41479 , n386500 );
buf ( n41481 , n34753 );
and ( n41482 , n41481 , n34754 );
not ( n41483 , n41481 );
and ( n41484 , n41483 , n386202 );
nor ( n41485 , n41482 , n41484 );
and ( n41486 , n41485 , n34765 );
buf ( n41487 , n385835 );
not ( n41488 , n41487 );
not ( n41489 , n385257 );
and ( n41490 , n41488 , n41489 );
and ( n41491 , n41487 , n385257 );
nor ( n41492 , n41490 , n41491 );
not ( n41493 , n386017 );
or ( n41494 , n41492 , n41493 );
nand ( n41495 , n41300 , RI15b4b900_443);
nand ( n41496 , n41494 , n41495 );
nor ( n41497 , n41486 , n41496 );
nand ( n41498 , n41480 , n41497 );
not ( n41499 , n41498 );
not ( n41500 , n41266 );
not ( n41501 , n41475 );
and ( n41502 , n41500 , n41501 );
or ( n41503 , n386541 , n385837 );
or ( n41504 , n385257 , n386550 );
or ( n41505 , n34754 , n386557 );
nand ( n41506 , n41503 , n41504 , n41505 );
nor ( n41507 , n41502 , n41506 );
nand ( n41508 , n41499 , n41507 );
buf ( n41509 , n41508 );
buf ( n41510 , n32160 );
buf ( n41511 , n21800 );
and ( n41512 , n35357 , n35363 );
buf ( n41513 , n35186 );
nor ( n41514 , n41512 , n41513 );
or ( n41515 , n41514 , n34980 );
and ( n41516 , n35537 , RI15b43188_154);
buf ( n41517 , n35384 );
and ( n41518 , n41517 , RI15b42dc8_146);
nor ( n41519 , n41516 , n41518 );
and ( n41520 , n35376 , RI15b43908_170);
and ( n41521 , n35373 , RI15b43548_162);
nor ( n41522 , n41520 , n41521 );
nor ( n41523 , n32749 , n20110 );
and ( n41524 , n41523 , RI15b40c08_74);
nor ( n41525 , n35568 , n383381 );
and ( n41526 , n41525 , RI15b40848_66);
nor ( n41527 , n41524 , n41526 );
nand ( n41528 , n35567 , n37342 );
not ( n41529 , n41528 );
and ( n41530 , n41529 , RI15b40488_58);
nand ( n41531 , n381061 , n37322 );
not ( n41532 , n41531 );
and ( n41533 , n41532 , RI15b400c8_50);
and ( n41534 , n35448 , RI15b41388_90);
and ( n41535 , n37294 , RI15b40fc8_82);
not ( n41536 , n35431 );
and ( n41537 , n41536 , RI15b41748_98);
nor ( n41538 , n41535 , n41537 );
and ( n41539 , n35422 , RI15b41b08_106);
and ( n41540 , n35412 , RI15b41ec8_114);
nor ( n41541 , n41539 , n41540 );
and ( n41542 , n35415 , RI15b42a08_138);
and ( n41543 , n35555 , RI15b42648_130);
nor ( n41544 , n41542 , n41543 );
or ( n41545 , n35390 , n385525 );
nand ( n41546 , n41538 , n41541 , n41544 , n41545 );
nor ( n41547 , n41534 , n41546 );
nor ( n41548 , n32749 , n41547 );
nor ( n41549 , n41530 , n41533 , n41548 );
nand ( n41550 , n41519 , n41522 , n41527 , n41549 );
not ( n41551 , n35455 );
and ( n41552 , n41550 , n41551 );
and ( n41553 , n35335 , RI15b661b0_1349);
or ( n41554 , n35357 , n34937 , RI15b48de0_351);
or ( n41555 , n34980 , RI15b48d68_350);
nand ( n41556 , n41554 , n41555 );
and ( n41557 , n41556 , n35363 );
nor ( n41558 , n41552 , n41553 , n41557 );
and ( n41559 , n35459 , n22266 );
and ( n41560 , n35461 , RI15b65a30_1333);
nor ( n41561 , n41559 , n41560 );
nand ( n41562 , n41515 , n41558 , n41561 );
buf ( n41563 , n41562 );
buf ( n41564 , n381081 );
buf ( n41565 , n381021 );
or ( n41566 , n381015 , n22039 );
nand ( n41567 , n35525 , RI15b53bc8_722);
nand ( n41568 , n41566 , n41567 );
buf ( n41569 , n41568 );
buf ( n41570 , n22653 );
buf ( n41571 , n22406 );
not ( n41572 , n40999 );
nand ( n41573 , n41572 , n379825 );
not ( n41574 , n41573 );
not ( n41575 , n41032 );
or ( n41576 , n41574 , n41575 );
nand ( n41577 , n41576 , n41000 );
not ( n41578 , n41036 );
nor ( n41579 , n41572 , n41000 );
nand ( n41580 , n41578 , n41579 );
buf ( n41581 , n379832 );
buf ( n41582 , n41581 );
nand ( n41583 , n41582 , RI15b46338_260);
and ( n41584 , n35459 , n36926 );
and ( n41585 , n35461 , RI15b65b20_1335);
nor ( n41586 , n41584 , n41585 );
nand ( n41587 , n41577 , n41580 , n41583 , n41586 );
buf ( n41588 , n41587 );
buf ( n41589 , n381006 );
buf ( n41590 , n379893 );
buf ( n41591 , n22408 );
or ( n41592 , n31149 , n41443 );
and ( n41593 , n31161 , n41446 );
or ( n41594 , n41455 , n17653 );
or ( n41595 , n32452 , n41461 );
or ( n41596 , n41453 , n31184 );
nand ( n41597 , n41594 , n41595 , n41596 );
nor ( n41598 , n41593 , n41597 );
nand ( n41599 , n41592 , n41598 );
buf ( n41600 , n41599 );
buf ( n41601 , n384199 );
and ( n41602 , n41420 , n31127 );
nor ( n41603 , n41602 , n36536 );
or ( n41604 , n41603 , n33484 );
or ( n41605 , n31124 , n39775 );
not ( n41606 , RI15b61728_1190);
or ( n41607 , n41420 , n41606 , RI15b617a0_1191);
or ( n41608 , n33484 , RI15b61728_1190);
nand ( n41609 , n41607 , n41608 );
and ( n41610 , n41609 , n31127 );
not ( n41611 , n32358 );
nor ( n41612 , n31052 , n380474 );
nor ( n41613 , n41610 , n41611 , n41612 );
nand ( n41614 , n41604 , n41605 , n41613 );
buf ( n41615 , n41614 );
buf ( n41616 , n33382 );
buf ( n41617 , RI15b47c10_313);
buf ( n41618 , n20665 );
buf ( n41619 , n22738 );
buf ( n41620 , n382073 );
and ( n41621 , n36999 , RI15b48048_322);
and ( n41622 , n37001 , RI15b44e98_216);
nor ( n41623 , n41621 , n41622 );
not ( n41624 , n41623 );
buf ( n41625 , n41624 );
buf ( n41626 , n382067 );
buf ( n41627 , n22653 );
buf ( n41628 , n22655 );
or ( n41629 , n381907 , n36121 );
and ( n41630 , n36308 , n36123 );
not ( n41631 , RI15b43818_168);
or ( n41632 , n36132 , n41631 );
or ( n41633 , n36321 , n36139 );
or ( n41634 , n36130 , n36327 );
nand ( n41635 , n41632 , n41633 , n41634 );
nor ( n41636 , n41630 , n41635 );
nand ( n41637 , n41629 , n41636 );
buf ( n41638 , n41637 );
buf ( n41639 , n385112 );
buf ( n41640 , n32271 );
buf ( n41641 , n379895 );
buf ( n41642 , n380942 );
not ( n41643 , n379825 );
not ( n41644 , n35067 );
nor ( n41645 , n41026 , n41644 );
buf ( n41646 , n41645 );
not ( n41647 , n41646 );
or ( n41648 , n41643 , n41647 );
nand ( n41649 , n41648 , n41032 );
nand ( n41650 , n41649 , n35034 );
not ( n41651 , n41036 );
not ( n41652 , n41646 );
not ( n41653 , n35034 );
nand ( n41654 , n41651 , n41652 , n41653 );
nand ( n41655 , n41582 , RI15b464a0_263);
and ( n41656 , n35461 , n32490 );
not ( n41657 , n381988 );
and ( n41658 , n35459 , n41657 );
nor ( n41659 , n41656 , n41658 );
nand ( n41660 , n41650 , n41654 , n41655 , n41659 );
buf ( n41661 , n41660 );
buf ( n41662 , n32672 );
buf ( n41663 , n384199 );
buf ( n41664 , n32271 );
or ( n41665 , n385163 , n20916 );
and ( n41666 , n36472 , n21580 );
and ( n41667 , n32368 , n20926 );
and ( n41668 , n385177 , n39061 );
nor ( n41669 , n41666 , n41667 , n41668 );
nand ( n41670 , n41665 , n41669 , n39101 );
buf ( n41671 , n41670 );
buf ( n41672 , n33382 );
not ( n41673 , n33559 );
nor ( n41674 , n41673 , n33568 );
nand ( n41675 , n41674 , n384934 );
not ( n41676 , n37772 );
not ( n41677 , n33568 );
or ( n41678 , n41676 , n41677 );
nand ( n41679 , n41678 , n32343 );
nand ( n41680 , n41679 , n41673 );
nand ( n41681 , n384918 , RI15b5ecf8_1100);
buf ( n41682 , n384823 );
nand ( n41683 , n384906 , n41682 );
nand ( n41684 , n41675 , n41680 , n41681 , n41683 );
buf ( n41685 , n41684 );
not ( n41686 , RI15b53628_710);
not ( n41687 , n383170 );
or ( n41688 , n41686 , n41687 );
xor ( n41689 , n381437 , n381438 );
and ( n41690 , n33453 , n41689 );
and ( n41691 , n383147 , RI15b52ea8_694);
nor ( n41692 , n41690 , n41691 );
nand ( n41693 , n41688 , n41692 );
buf ( n41694 , n41693 );
buf ( n41695 , n385195 );
buf ( n41696 , n32672 );
or ( n41697 , n383180 , n35984 );
not ( n41698 , n35996 );
and ( n41699 , n41698 , RI15b5b878_988);
or ( n41700 , n383184 , n35986 );
not ( n41701 , n40016 );
and ( n41702 , n36002 , n41701 );
and ( n41703 , n40019 , n35999 );
nor ( n41704 , n41702 , n41703 );
nand ( n41705 , n41700 , n41704 );
nor ( n41706 , n41699 , n41705 );
nand ( n41707 , n41697 , n41706 );
buf ( n41708 , n41707 );
buf ( n41709 , n22404 );
and ( n41710 , n38047 , RI15b53f88_730);
and ( n41711 , n35213 , RI15b66480_1355);
nor ( n41712 , n41710 , n41711 );
not ( n41713 , n41712 );
buf ( n41714 , n41713 );
buf ( n41715 , n41551 );
and ( n41716 , n32803 , n41715 );
and ( n41717 , n35335 , RI15b65df0_1341);
not ( n41718 , RI15b48a20_343);
not ( n41719 , n35350 );
not ( n41720 , n41719 );
or ( n41721 , n41718 , n41720 );
or ( n41722 , n41719 , RI15b48a20_343);
nand ( n41723 , n41721 , n41722 );
and ( n41724 , n35363 , n41723 );
nor ( n41725 , n41716 , n41717 , n41724 );
buf ( n41726 , n41513 );
nand ( n41727 , n41726 , RI15b48a20_343);
nand ( n41728 , n38861 , n41725 , n41727 );
buf ( n41729 , n41728 );
buf ( n41730 , n22716 );
buf ( n41731 , n22653 );
buf ( n41732 , n31033 );
not ( n41733 , RI15b61890_1193);
nand ( n41734 , n41422 , RI15b61818_1192);
nand ( n41735 , n41734 , n31080 );
nand ( n41736 , n41735 , n31091 );
not ( n41737 , n41736 );
or ( n41738 , n41733 , n41737 );
and ( n41739 , n38666 , n38693 );
not ( n41740 , n39714 );
nor ( n41741 , n41739 , n39914 , n41740 );
and ( n41742 , n41741 , n39368 );
not ( n41743 , n41734 );
nor ( n41744 , n31079 , RI15b61890_1193);
and ( n41745 , n41743 , n41744 );
or ( n41746 , n31052 , n380461 );
nand ( n41747 , n41746 , n41683 );
nor ( n41748 , n41742 , n41745 , n41747 );
nand ( n41749 , n41738 , n41748 );
buf ( n41750 , n41749 );
buf ( n41751 , n384199 );
or ( n41752 , n36238 , n41445 );
or ( n41753 , n17974 , n41455 );
not ( n41754 , n41461 );
and ( n41755 , n41754 , n32711 );
not ( n41756 , n41443 );
and ( n41757 , n383803 , n41756 );
and ( n41758 , n36261 , n41459 );
nor ( n41759 , n41755 , n41757 , n41758 );
nand ( n41760 , n41752 , n41753 , n41759 );
buf ( n41761 , n41760 );
buf ( n41762 , n22408 );
buf ( n41763 , RI15b47850_305);
buf ( n41764 , n386760 );
not ( n41765 , n384327 );
not ( n41766 , n41765 );
not ( n41767 , n32539 );
not ( n41768 , n41767 );
or ( n41769 , n41766 , n41768 );
not ( n41770 , n41767 );
nand ( n41771 , n41770 , n384327 );
nand ( n41772 , n41769 , n41771 );
and ( n41773 , n41772 , n384392 );
not ( n41774 , n38915 );
nor ( n41775 , n41774 , n384433 );
not ( n41776 , n41775 );
not ( n41777 , n384429 );
and ( n41778 , n41776 , n41777 );
and ( n41779 , n41775 , n384429 );
nor ( n41780 , n41778 , n41779 );
or ( n41781 , n41780 , n384494 );
not ( n41782 , n384550 );
not ( n41783 , n32552 );
not ( n41784 , n41783 );
or ( n41785 , n41782 , n41784 );
or ( n41786 , n41783 , n384550 );
nand ( n41787 , n41785 , n41786 );
and ( n41788 , n41787 , n380811 );
and ( n41789 , n19513 , RI15b64068_1278);
nor ( n41790 , n41788 , n41789 );
nand ( n41791 , n41781 , n41790 );
nor ( n41792 , n41773 , n41791 );
or ( n41793 , n32581 , n386842 );
or ( n41794 , n22775 , n38109 );
or ( n41795 , RI15b63168_1246 , n384652 );
nand ( n41796 , n41793 , n41794 , n41795 );
not ( n41797 , n41796 );
nand ( n41798 , n41792 , n41797 );
buf ( n41799 , n41798 );
buf ( n41800 , n19651 );
buf ( n41801 , n382537 );
not ( n41802 , n19883 );
nor ( n41803 , n41802 , n19922 );
not ( n41804 , n19942 );
or ( n41805 , n41803 , n41804 );
not ( n41806 , n19890 );
nand ( n41807 , n41805 , n41806 );
buf ( n41808 , n19992 );
not ( n41809 , n41808 );
nor ( n41810 , n41809 , n20502 );
or ( n41811 , n41810 , n20521 );
nand ( n41812 , n41811 , RI15b49f38_388);
or ( n41813 , n41808 , n20529 , RI15b49f38_388);
or ( n41814 , n382130 , RI15b4bcc0_451);
nand ( n41815 , n20556 , n382130 , RI15b4bcc0_451);
nand ( n41816 , n41814 , n41815 );
and ( n41817 , n20647 , n41816 );
and ( n41818 , n20656 , RI15b4ae38_420);
nor ( n41819 , n41817 , n41818 );
nand ( n41820 , n41813 , n41819 );
not ( n41821 , n38996 );
not ( n41822 , n20556 );
and ( n41823 , n41821 , n41822 );
nor ( n41824 , n41823 , n20641 );
nor ( n41825 , n41824 , n382130 );
nor ( n41826 , n41820 , n41825 );
buf ( n41827 , n380871 );
not ( n41828 , n41827 );
nand ( n41829 , n41802 , n41828 , n19890 );
nand ( n41830 , n41807 , n41812 , n41826 , n41829 );
buf ( n41831 , n41830 );
buf ( n41832 , n384700 );
buf ( n41833 , n36704 );
not ( n41834 , RI15b47670_301);
not ( n41835 , n385213 );
or ( n41836 , n41834 , n41835 );
not ( n41837 , n34930 );
not ( n41838 , n34964 );
and ( n41839 , n41837 , n41838 );
and ( n41840 , n20631 , RI15b46068_254);
nor ( n41841 , n41839 , n41840 );
nand ( n41842 , n41836 , n41841 );
buf ( n41843 , n41842 );
buf ( n41844 , n380903 );
buf ( n41845 , n22404 );
buf ( n41846 , n383345 );
buf ( n41847 , n22740 );
buf ( n41848 , n384700 );
buf ( n41849 , n22788 );
not ( n41850 , RI15b524d0_673);
not ( n41851 , n32397 );
or ( n41852 , n41850 , n41851 );
not ( n41853 , n381424 );
not ( n41854 , n383052 );
and ( n41855 , n41853 , n41854 );
not ( n41856 , n32709 );
nand ( n41857 , n381401 , n41856 );
not ( n41858 , n41857 );
nor ( n41859 , n41855 , n41858 );
nand ( n41860 , n41852 , n41859 );
buf ( n41861 , n41860 );
and ( n41862 , n31792 , n384550 );
not ( n41863 , RI15b5c9d0_1025);
or ( n41864 , n31771 , n41863 );
or ( n41865 , n384327 , n37611 );
or ( n41866 , n384429 , n31779 );
nand ( n41867 , n41864 , n41865 , n41866 );
nor ( n41868 , n41862 , n41867 );
nand ( n41869 , n41792 , n41868 );
buf ( n41870 , n41869 );
buf ( n41871 , n22408 );
not ( n41872 , n386590 );
not ( n41873 , n33400 );
or ( n41874 , n41872 , n41873 );
and ( n41875 , n33415 , n386603 );
or ( n41876 , n386612 , n18492 );
or ( n41877 , n36293 , n386624 );
or ( n41878 , n386610 , n33443 );
nand ( n41879 , n41876 , n41877 , n41878 );
nor ( n41880 , n41875 , n41879 );
nand ( n41881 , n41874 , n41880 );
buf ( n41882 , n41881 );
buf ( n41883 , n382049 );
buf ( n41884 , n384218 );
buf ( n41885 , n381240 );
buf ( n41886 , n41885 );
or ( n41887 , n32430 , n41886 );
not ( n41888 , n381275 );
nand ( n41889 , n381417 , n41888 );
and ( n41890 , n386637 , RI15b54e88_762);
and ( n41891 , n381636 , RI15b4eab0_549);
and ( n41892 , n381639 , RI15b4e6f0_541);
nor ( n41893 , n41891 , n41892 );
and ( n41894 , n381643 , RI15b4ee70_557);
not ( n41895 , n381650 );
not ( n41896 , n41895 );
and ( n41897 , n41896 , RI15b4dbb0_517);
and ( n41898 , n381657 , RI15b4fd70_589);
nor ( n41899 , n41897 , n41898 );
and ( n41900 , n381661 , RI15b4f9b0_581);
and ( n41901 , n381663 , RI15b4f230_565);
nor ( n41902 , n41900 , n41901 );
and ( n41903 , n381667 , RI15b4d430_501);
and ( n41904 , n381669 , RI15b4d7f0_509);
nor ( n41905 , n41903 , n41904 );
and ( n41906 , n381672 , RI15b4df70_525);
and ( n41907 , n381674 , RI15b4f5f0_573);
nor ( n41908 , n41906 , n41907 );
nand ( n41909 , n41899 , n41902 , n41905 , n41908 );
and ( n41910 , n381646 , n41909 );
and ( n41911 , n381680 , RI15b4c8f0_477);
nor ( n41912 , n41894 , n41910 , n41911 );
and ( n41913 , n381684 , RI15b4c530_469);
and ( n41914 , n381686 , RI15b4e330_533);
nor ( n41915 , n41913 , n41914 );
and ( n41916 , n381689 , RI15b4ccb0_485);
and ( n41917 , n381691 , RI15b4d070_493);
nor ( n41918 , n41916 , n41917 );
nand ( n41919 , n41893 , n41912 , n41915 , n41918 );
and ( n41920 , n41919 , n32437 );
not ( n41921 , RI15b54e88_762);
not ( n41922 , n382647 );
not ( n41923 , n41922 );
or ( n41924 , n41921 , n41923 );
or ( n41925 , n41922 , RI15b54e88_762);
nand ( n41926 , n41924 , n41925 );
and ( n41927 , n382627 , n41926 );
nor ( n41928 , n41890 , n41920 , n41927 );
and ( n41929 , n41889 , n41928 );
nand ( n41930 , n41887 , n41929 );
buf ( n41931 , n41930 );
buf ( n41932 , n383928 );
not ( n41933 , n41932 );
not ( n41934 , n41933 );
buf ( n41935 , n383967 );
and ( n41936 , n38654 , RI15b5b170_973);
and ( n41937 , n39717 , RI15b5adb0_965);
nor ( n41938 , n41936 , n41937 );
and ( n41939 , n39721 , RI15b5a9f0_957);
and ( n41940 , n39724 , RI15b5a630_949);
nor ( n41941 , n41939 , n41940 );
and ( n41942 , n39728 , RI15b5a270_941);
and ( n41943 , n39731 , RI15b59eb0_933);
nor ( n41944 , n41942 , n41943 );
and ( n41945 , n39735 , RI15b59af0_925);
and ( n41946 , n39738 , RI15b59730_917);
nor ( n41947 , n41945 , n41946 );
nand ( n41948 , n41938 , n41941 , n41944 , n41947 );
and ( n41949 , n41935 , n41948 );
and ( n41950 , n39746 , RI15b58bf0_893);
and ( n41951 , n39751 , RI15b5c070_1005);
nor ( n41952 , n41949 , n41950 , n41951 );
and ( n41953 , n39756 , RI15b5bcb0_997);
and ( n41954 , n39759 , RI15b5b8f0_989);
nor ( n41955 , n41953 , n41954 );
and ( n41956 , n39763 , RI15b59370_909);
and ( n41957 , n39765 , RI15b58fb0_901);
nor ( n41958 , n41956 , n41957 );
and ( n41959 , n39769 , RI15b58830_885);
and ( n41960 , n39772 , RI15b5b530_981);
nor ( n41961 , n41959 , n41960 );
nand ( n41962 , n41952 , n41955 , n41958 , n41961 );
not ( n41963 , n41962 );
or ( n41964 , n41934 , n41963 );
and ( n41965 , n384022 , RI15b62448_1218);
not ( n41966 , RI15b62448_1218);
not ( n41967 , n38478 );
or ( n41968 , n41966 , n41967 );
or ( n41969 , n38478 , RI15b62448_1218);
nand ( n41970 , n41968 , n41969 );
and ( n41971 , n41970 , n384025 );
nor ( n41972 , n41965 , n41971 );
nand ( n41973 , n41964 , n41972 );
buf ( n41974 , n41973 );
buf ( n41975 , n22740 );
buf ( n41976 , n36854 );
buf ( n41977 , n385112 );
buf ( n41978 , n381021 );
not ( n41979 , n39691 );
not ( n41980 , n41979 );
not ( n41981 , n384726 );
or ( n41982 , n41980 , n41981 );
and ( n41983 , n384737 , n39694 );
or ( n41984 , n39703 , n17755 );
or ( n41985 , n384754 , n39707 );
or ( n41986 , n39701 , n384759 );
nand ( n41987 , n41984 , n41985 , n41986 );
nor ( n41988 , n41983 , n41987 );
nand ( n41989 , n41982 , n41988 );
buf ( n41990 , n41989 );
not ( n41991 , n41853 );
not ( n41992 , n41991 );
not ( n41993 , n41992 );
not ( n41994 , n383320 );
or ( n41995 , n41993 , n41994 );
nand ( n41996 , n41995 , n381450 );
not ( n41997 , n383326 );
nand ( n41998 , n41996 , n41997 );
not ( n41999 , n383320 );
nor ( n42000 , n41997 , n381460 );
and ( n42001 , n41999 , n42000 );
not ( n42002 , RI15b52ae8_686);
not ( n42003 , n32397 );
or ( n42004 , n42002 , n42003 );
not ( n42005 , n382889 );
nand ( n42006 , n42004 , n42005 );
nor ( n42007 , n42001 , n42006 );
nand ( n42008 , n41998 , n42007 );
buf ( n42009 , n42008 );
and ( n42010 , n40930 , n19336 );
not ( n42011 , n19429 );
or ( n42012 , n42011 , n19280 );
and ( n42013 , n19280 , RI15b5c3b8_1012);
buf ( n42014 , n18666 );
nor ( n42015 , n42014 , n19336 );
nor ( n42016 , n42013 , n42015 );
nand ( n42017 , n42012 , n42016 );
and ( n42018 , n19194 , n42017 );
not ( n42019 , n19549 );
nand ( n42020 , n42019 , n22470 , n19556 );
and ( n42021 , n42020 , RI15b5c3b8_1012);
nor ( n42022 , n42010 , n42018 , n42021 );
or ( n42023 , n42022 , n19200 );
and ( n42024 , n31778 , n19336 );
not ( n42025 , RI15b5c3b8_1012);
not ( n42026 , n31767 );
or ( n42027 , n42025 , n42026 );
buf ( n42028 , n42014 );
or ( n42029 , n42028 , RI15b5c3b8_1012);
not ( n42030 , n18667 );
nand ( n42031 , n42029 , n42030 );
and ( n42032 , n19498 , n42031 );
and ( n42033 , n19513 , RI15b63a50_1265);
nor ( n42034 , n42032 , n42033 );
nand ( n42035 , n42027 , n42034 );
nor ( n42036 , n42024 , n42035 );
nand ( n42037 , n42023 , n42036 );
buf ( n42038 , n42037 );
buf ( n42039 , n383174 );
buf ( n42040 , n32672 );
buf ( n42041 , n22738 );
buf ( n42042 , n31558 );
and ( n42043 , n42042 , n31565 );
not ( n42044 , n42042 );
not ( n42045 , n31565 );
and ( n42046 , n42044 , n42045 );
nor ( n42047 , n42043 , n42046 );
nand ( n42048 , n42047 , n31599 );
not ( n42049 , n31652 );
and ( n42050 , n42049 , n379391 );
or ( n42051 , n42050 , n31699 );
nand ( n42052 , n42051 , n31330 );
or ( n42053 , n42049 , n31705 );
not ( n42054 , n42053 );
nand ( n42055 , n42054 , n379218 );
and ( n42056 , n379394 , RI15b57e58_864);
and ( n42057 , n31712 , RI15b51c60_655);
nor ( n42058 , n42056 , n42057 );
nand ( n42059 , n42048 , n42052 , n42055 , n42058 );
buf ( n42060 , n42059 );
buf ( n42061 , n35649 );
or ( n42062 , n384244 , n40947 );
nor ( n42063 , n31871 , n31925 , RI15b5d240_1043);
and ( n42064 , n384244 , n42063 );
not ( n42065 , n31871 );
not ( n42066 , n31925 );
and ( n42067 , n42065 , n42066 );
nor ( n42068 , n42067 , n40947 );
nor ( n42069 , n42064 , n42068 );
nand ( n42070 , n42062 , n42069 );
not ( n42071 , n42070 );
not ( n42072 , n31919 );
or ( n42073 , n42071 , n42072 );
or ( n42074 , n31919 , n42070 );
nand ( n42075 , n42073 , n42074 );
buf ( n42076 , n31923 );
and ( n42077 , n42075 , n42076 );
or ( n42078 , n384600 , n40947 );
and ( n42079 , n384600 , n42063 );
nor ( n42080 , n42079 , n42068 );
nand ( n42081 , n42078 , n42080 );
not ( n42082 , n42081 );
not ( n42083 , n31953 );
nand ( n42084 , n42083 , n31928 );
not ( n42085 , n42084 );
or ( n42086 , n42082 , n42085 );
or ( n42087 , n42084 , n42081 );
nand ( n42088 , n42086 , n42087 );
buf ( n42089 , n31960 );
and ( n42090 , n42088 , n42089 );
nor ( n42091 , n42077 , n42090 );
not ( n42092 , n31775 );
or ( n42093 , n42092 , n40947 );
nand ( n42094 , n42092 , n42063 );
not ( n42095 , n42068 );
nand ( n42096 , n42093 , n42094 , n42095 );
not ( n42097 , n42096 );
buf ( n42098 , n31859 );
not ( n42099 , n31882 );
or ( n42100 , n42098 , n42099 );
nor ( n42101 , n31866 , n31876 );
or ( n42102 , n42101 , n42099 );
nand ( n42103 , n42100 , n42102 );
not ( n42104 , n42103 );
or ( n42105 , n42097 , n42104 );
not ( n42106 , n42101 );
nor ( n42107 , n42106 , n42096 );
and ( n42108 , n42098 , n42107 , n31884 );
nor ( n42109 , n19512 , n379589 );
nor ( n42110 , n42108 , n42109 );
nand ( n42111 , n42105 , n42110 );
not ( n42112 , n42081 );
not ( n42113 , n31792 );
or ( n42114 , n42112 , n42113 );
not ( n42115 , n32378 );
buf ( n42116 , n42115 );
not ( n42117 , n42116 );
not ( n42118 , n42117 );
and ( n42119 , n42070 , n42118 );
and ( n42120 , n42096 , n31778 );
and ( n42121 , n31770 , RI15b5d240_1043);
nor ( n42122 , n42119 , n42120 , n42121 );
nand ( n42123 , n42114 , n42122 );
nor ( n42124 , n42111 , n42123 );
nand ( n42125 , n42091 , n42124 );
buf ( n42126 , n42125 );
buf ( n42127 , n387159 );
buf ( n42128 , n386760 );
not ( n42129 , n382512 );
nor ( n42130 , n382088 , n383358 );
or ( n42131 , n42130 , n382213 );
nand ( n42132 , n42131 , n382450 );
or ( n42133 , n42132 , n33145 );
xor ( n42134 , RI15b4b360_431 , n382088 );
not ( n42135 , n42134 );
or ( n42136 , n33145 , n42135 );
nand ( n42137 , n42136 , n382269 );
nand ( n42138 , n42133 , n42137 );
nand ( n42139 , n42129 , n42138 );
not ( n42140 , n382080 );
not ( n42141 , n382448 );
buf ( n42142 , n42141 );
not ( n42143 , n42142 );
or ( n42144 , n42140 , n42143 );
nand ( n42145 , n42144 , n382474 );
buf ( n42146 , n32835 );
not ( n42147 , n42146 );
nand ( n42148 , n42145 , n42147 );
not ( n42149 , n32035 );
not ( n42150 , n42142 );
nand ( n42151 , n42149 , n42146 , n42150 );
and ( n42152 , n382523 , RI15b4b3d8_432);
buf ( n42153 , n382528 );
and ( n42154 , n42153 , RI15b451e0_223);
nor ( n42155 , n42152 , n42154 );
nand ( n42156 , n42139 , n42148 , n42151 , n42155 );
buf ( n42157 , n42156 );
buf ( n42158 , n384996 );
buf ( n42159 , n22714 );
not ( n42160 , n379346 );
not ( n42161 , n379343 );
or ( n42162 , n42160 , n42161 );
and ( n42163 , n379394 , RI15b576d8_848);
and ( n42164 , n379398 , RI15b514e0_639);
and ( n42165 , n379391 , n379365 );
nor ( n42166 , n42163 , n42164 , n42165 );
nand ( n42167 , n42162 , n42166 );
buf ( n42168 , n42167 );
nor ( n42169 , n33955 , n379791 );
and ( n42170 , n42169 , n379413 );
not ( n42171 , n42169 );
and ( n42172 , n42171 , n379412 );
nor ( n42173 , n42170 , n42172 );
nand ( n42174 , n42173 , n379785 );
or ( n42175 , n33766 , n379413 );
or ( n42176 , n379412 , n33734 );
nand ( n42177 , n42175 , n42176 );
and ( n42178 , n379780 , n42177 );
and ( n42179 , n379783 , RI15b63bb8_1268);
and ( n42180 , n379796 , RI15b5d9c0_1059);
nor ( n42181 , n42179 , n42180 );
not ( n42182 , n42181 );
nor ( n42183 , n42178 , n42182 );
nand ( n42184 , n42174 , n42183 );
buf ( n42185 , n42184 );
buf ( n42186 , n379844 );
buf ( n42187 , n383174 );
not ( n42188 , n34814 );
buf ( n42189 , n386967 );
not ( n42190 , n42189 );
or ( n42191 , n42188 , n42190 );
nand ( n42192 , n42191 , n34823 );
and ( n42193 , n42192 , RI15b62088_1210);
and ( n42194 , n34812 , RI15b63e88_1274);
or ( n42195 , n34826 , n42189 , RI15b62088_1210);
not ( n42196 , n387027 );
not ( n42197 , n42196 );
not ( n42198 , RI15b63e88_1274);
and ( n42199 , n42197 , n42198 );
and ( n42200 , n42196 , RI15b63e88_1274);
nor ( n42201 , n42199 , n42200 );
or ( n42202 , n34833 , n42201 );
nand ( n42203 , n42195 , n42202 );
nor ( n42204 , n42193 , n42194 , n42203 );
or ( n42205 , n42204 , n19200 );
not ( n42206 , n386815 );
not ( n42207 , n42206 );
not ( n42208 , n22473 );
and ( n42209 , n42207 , n42208 );
nor ( n42210 , n42209 , n38114 );
or ( n42211 , n380852 , n42210 );
and ( n42212 , n387011 , n42206 , n380852 );
or ( n42213 , n22424 , n379556 );
or ( n42214 , n380850 , n19598 );
nand ( n42215 , n42213 , n42214 , n19512 );
nor ( n42216 , n42212 , n42215 );
nand ( n42217 , n42205 , n42211 , n42216 );
buf ( n42218 , n42217 );
buf ( n42219 , n32676 );
not ( n42220 , n20637 );
not ( n42221 , n19700 );
or ( n42222 , n42220 , n42221 );
nand ( n42223 , n42222 , n34798 );
and ( n42224 , n42223 , RI15b4b018_424);
or ( n42225 , n34801 , n19700 , RI15b4b018_424);
not ( n42226 , n19706 );
or ( n42227 , n42226 , n22216 );
nand ( n42228 , n42225 , n42227 );
nor ( n42229 , n42224 , n42228 );
nand ( n42230 , n386506 , n42229 );
buf ( n42231 , n42230 );
buf ( n42232 , n386762 );
buf ( n42233 , n386563 );
and ( n42234 , n22646 , RI15b45ac8_242);
and ( n42235 , n22648 , RI15b51f30_661);
nor ( n42236 , n42234 , n42235 );
not ( n42237 , n42236 );
buf ( n42238 , n42237 );
buf ( n42239 , n382071 );
not ( n42240 , RI15b53b50_721);
not ( n42241 , n383170 );
or ( n42242 , n42240 , n42241 );
or ( n42243 , n383152 , n41854 );
nand ( n42244 , n42243 , n383157 );
not ( n42245 , n383109 );
and ( n42246 , n42244 , n42245 );
nor ( n42247 , n42245 , n383052 );
and ( n42248 , n383143 , n42247 );
and ( n42249 , n383147 , RI15b52548_674);
nor ( n42250 , n42246 , n42248 , n42249 );
nand ( n42251 , n42242 , n42250 );
buf ( n42252 , n42251 );
not ( n42253 , n35145 );
not ( n42254 , n381589 );
or ( n42255 , n42253 , n42254 );
and ( n42256 , n381596 , n35150 );
or ( n42257 , n35160 , n18698 );
not ( n42258 , n32419 );
or ( n42259 , n42258 , n35166 );
or ( n42260 , n35158 , n381621 );
nand ( n42261 , n42257 , n42259 , n42260 );
nor ( n42262 , n42256 , n42261 );
nand ( n42263 , n42255 , n42262 );
buf ( n42264 , n42263 );
buf ( n42265 , n385112 );
buf ( n42266 , n383174 );
buf ( n42267 , n22408 );
or ( n42268 , n36119 , n36082 );
and ( n42269 , n38230 , RI15b411a8_86);
or ( n42270 , n35582 , n36098 );
or ( n42271 , n35856 , n36092 );
or ( n42272 , n36086 , n35858 );
nand ( n42273 , n42270 , n42271 , n42272 );
nor ( n42274 , n42269 , n42273 );
nand ( n42275 , n42268 , n42274 );
buf ( n42276 , n42275 );
and ( n42277 , n38248 , RI15b3fe70_45);
buf ( n42278 , n42277 );
buf ( n42279 , n30992 );
buf ( n42280 , n386760 );
buf ( n42281 , n22009 );
not ( n42282 , RI15b53bc8_722);
not ( n42283 , n32244 );
or ( n42284 , n42282 , n42283 );
and ( n42285 , n32247 , RI15b651c0_1315);
and ( n42286 , n32249 , RI15b60030_1141);
nor ( n42287 , n42285 , n42286 );
nand ( n42288 , n42284 , n42287 );
buf ( n42289 , n42288 );
buf ( n42290 , n386563 );
buf ( n42291 , n22479 );
buf ( n42292 , n386762 );
buf ( n42293 , n32981 );
or ( n42294 , n381056 , n19985 );
not ( n42295 , n41550 );
or ( n42296 , n32807 , n42295 );
and ( n42297 , n37123 , RI15b49ce0_383);
not ( n42298 , n37123 );
and ( n42299 , n42298 , n19985 );
nor ( n42300 , n42297 , n42299 );
or ( n42301 , n37110 , n42300 );
nand ( n42302 , n42294 , n42296 , n42301 );
buf ( n42303 , n42302 );
buf ( n42304 , n22402 );
buf ( n42305 , n22716 );
buf ( n42306 , n19839 );
and ( n42307 , n42306 , n19920 );
nor ( n42308 , n42307 , n38940 );
or ( n42309 , n42308 , n34803 );
not ( n42310 , n42306 );
nand ( n42311 , n380870 , n42310 , n34803 );
and ( n42312 , n20641 , RI15b4ba68_446);
buf ( n42313 , n19982 );
and ( n42314 , n42313 , n31806 );
nor ( n42315 , n42314 , n31809 );
or ( n42316 , n42315 , n19983 );
not ( n42317 , n20552 );
and ( n42318 , n42317 , RI15b4ba68_446);
not ( n42319 , n42317 );
and ( n42320 , n42319 , n382119 );
nor ( n42321 , n42318 , n42320 );
or ( n42322 , n42321 , n22354 );
not ( n42323 , n42313 );
and ( n42324 , n42323 , n22361 , n19983 );
buf ( n42325 , n20652 );
not ( n42326 , n42325 );
or ( n42327 , n42326 , n19687 );
not ( n42328 , n22394 );
nand ( n42329 , n42327 , n42328 );
nor ( n42330 , n42324 , n42329 );
nand ( n42331 , n42316 , n42322 , n42330 );
nor ( n42332 , n42312 , n42331 );
nand ( n42333 , n42309 , n42311 , n42332 );
buf ( n42334 , n42333 );
buf ( n42335 , n384700 );
buf ( n42336 , n32271 );
not ( n42337 , n383440 );
not ( n42338 , n381497 );
or ( n42339 , n42337 , n42338 );
nand ( n42340 , n42339 , n32582 );
and ( n42341 , n42340 , RI15b63438_1252);
or ( n42342 , n384652 , n383440 , RI15b63438_1252);
or ( n42343 , n386892 , n22775 );
nand ( n42344 , n42342 , n42343 );
nor ( n42345 , n42341 , n42344 );
nand ( n42346 , n39571 , n42345 );
buf ( n42347 , n42346 );
buf ( n42348 , n381872 );
buf ( n42349 , n386563 );
buf ( n42350 , n385112 );
not ( n42351 , n383930 );
and ( n42352 , n383945 , RI15b587b8_884);
and ( n42353 , n383949 , RI15b5a5b8_948);
nor ( n42354 , n42352 , n42353 );
and ( n42355 , n383955 , RI15b5ad38_964);
and ( n42356 , n383960 , RI15b5a978_956);
nor ( n42357 , n42355 , n42356 );
and ( n42358 , n383965 , RI15b5b0f8_972);
and ( n42359 , n383970 , RI15b59e38_932);
and ( n42360 , n383972 , RI15b5a1f8_940);
nor ( n42361 , n42359 , n42360 );
and ( n42362 , n383975 , RI15b596b8_916);
and ( n42363 , n383977 , RI15b59a78_924);
nor ( n42364 , n42362 , n42363 );
and ( n42365 , n383982 , RI15b5bc38_996);
and ( n42366 , n383984 , RI15b5b878_988);
nor ( n42367 , n42365 , n42366 );
and ( n42368 , n383987 , RI15b5bff8_1004);
and ( n42369 , n383989 , RI15b5b4b8_980);
nor ( n42370 , n42368 , n42369 );
nand ( n42371 , n42361 , n42364 , n42367 , n42370 );
and ( n42372 , n383968 , n42371 );
and ( n42373 , n383994 , RI15b58b78_892);
nor ( n42374 , n42358 , n42372 , n42373 );
and ( n42375 , n383997 , RI15b58f38_900);
and ( n42376 , n383999 , RI15b592f8_908);
nor ( n42377 , n42375 , n42376 );
nand ( n42378 , n42354 , n42357 , n42374 , n42377 );
not ( n42379 , n42378 );
or ( n42380 , n42351 , n42379 );
and ( n42381 , n384022 , RI15b62010_1209);
not ( n42382 , RI15b62010_1209);
not ( n42383 , n384036 );
not ( n42384 , n42383 );
or ( n42385 , n42382 , n42384 );
or ( n42386 , n42383 , RI15b62010_1209);
nand ( n42387 , n42385 , n42386 );
and ( n42388 , n384025 , n42387 );
nor ( n42389 , n42381 , n42388 );
nand ( n42390 , n42380 , n42389 );
buf ( n42391 , n42390 );
and ( n42392 , n22646 , RI15b457f8_236);
and ( n42393 , n22648 , RI15b51c60_655);
nor ( n42394 , n42392 , n42393 );
not ( n42395 , n42394 );
buf ( n42396 , n42395 );
or ( n42397 , n36238 , n386717 );
not ( n42398 , n386727 );
and ( n42399 , n42398 , RI15b4ce90_489);
or ( n42400 , n386735 , n32710 );
or ( n42401 , n386706 , n383802 );
not ( n42402 , n36261 );
or ( n42403 , n386725 , n42402 );
nand ( n42404 , n42400 , n42401 , n42403 );
nor ( n42405 , n42399 , n42404 );
nand ( n42406 , n42397 , n42405 );
buf ( n42407 , n42406 );
or ( n42408 , n36119 , n36200 );
not ( n42409 , n36212 );
and ( n42410 , n42409 , RI15b41568_94);
or ( n42411 , n35582 , n36217 );
or ( n42412 , n35856 , n36210 );
or ( n42413 , n36204 , n35858 );
nand ( n42414 , n42411 , n42412 , n42413 );
nor ( n42415 , n42410 , n42414 );
nand ( n42416 , n42408 , n42415 );
buf ( n42417 , n42416 );
buf ( n42418 , n383174 );
buf ( n42419 , n30992 );
and ( n42420 , n22646 , RI15b451e0_223);
and ( n42421 , n22648 , RI15b51648_642);
nor ( n42422 , n42420 , n42421 );
not ( n42423 , n42422 );
buf ( n42424 , n42423 );
buf ( n42425 , n381566 );
buf ( n42426 , n381006 );
buf ( n42427 , n379844 );
buf ( n42428 , n22740 );
buf ( n42429 , n19651 );
buf ( n42430 , n21800 );
not ( n42431 , n382057 );
buf ( n42432 , n382277 );
not ( n42433 , n42432 );
or ( n42434 , n42431 , n42433 );
not ( n42435 , n382058 );
not ( n42436 , n382062 );
or ( n42437 , n42435 , n42436 );
nand ( n42438 , n42437 , RI15b4b180_427);
nand ( n42439 , n42434 , n42438 );
buf ( n42440 , n42439 );
not ( n42441 , n19201 );
not ( n42442 , RI15b5d420_1047);
not ( n42443 , n40937 );
or ( n42444 , n42442 , n42443 );
buf ( n42445 , n18262 );
buf ( n42446 , n42445 );
and ( n42447 , n40930 , n42446 );
or ( n42448 , n32385 , n383941 );
not ( n42449 , n40928 );
not ( n42450 , n383959 );
or ( n42451 , n42450 , RI15b5d420_1047);
nand ( n42452 , n42451 , n18258 );
and ( n42453 , n42449 , n42452 );
not ( n42454 , n383939 );
and ( n42455 , n42450 , n42454 );
nor ( n42456 , n42453 , n42455 );
nand ( n42457 , n42448 , n42456 );
nor ( n42458 , n42447 , n42457 );
nand ( n42459 , n42444 , n42458 );
not ( n42460 , n42459 );
or ( n42461 , n42441 , n42460 );
and ( n42462 , n40943 , RI15b5d420_1047);
and ( n42463 , n380789 , n42446 );
nor ( n42464 , n42462 , n42463 );
nand ( n42465 , n42461 , n42464 );
buf ( n42466 , n42465 );
buf ( n42467 , n384203 );
not ( n42468 , n40964 );
nor ( n42469 , n42468 , n31667 );
or ( n42470 , n42469 , n31699 );
nand ( n42471 , n42470 , n379167 );
not ( n42472 , n31534 );
not ( n42473 , n31526 );
not ( n42474 , n42473 );
or ( n42475 , n42472 , n42474 );
or ( n42476 , n42473 , n31534 );
nand ( n42477 , n42475 , n42476 );
and ( n42478 , n31599 , n42477 );
not ( n42479 , RI15b51a80_651);
not ( n42480 , n379398 );
or ( n42481 , n42479 , n42480 );
not ( n42482 , n379394 );
or ( n42483 , n42482 , n21940 );
nand ( n42484 , n42481 , n42483 );
nor ( n42485 , n42478 , n42484 );
nand ( n42486 , n42468 , n31708 , n379168 );
nand ( n42487 , n42471 , n42485 , n42486 );
buf ( n42488 , n42487 );
buf ( n42489 , n36854 );
buf ( n42490 , n34857 );
not ( n42491 , n42490 );
not ( n42492 , n34856 );
or ( n42493 , n42491 , n42492 );
or ( n42494 , n34856 , n42490 );
nand ( n42495 , n42493 , n42494 );
nand ( n42496 , n42495 , n31599 );
not ( n42497 , n31618 );
not ( n42498 , n31623 );
not ( n42499 , n42498 );
or ( n42500 , n42497 , n42499 );
or ( n42501 , n42498 , n31618 );
nand ( n42502 , n42500 , n42501 );
and ( n42503 , n42502 , n379391 );
and ( n42504 , n379394 , RI15b578b8_852);
and ( n42505 , n379398 , RI15b516c0_643);
nor ( n42506 , n42503 , n42504 , n42505 );
nand ( n42507 , n42496 , n42506 );
buf ( n42508 , n42507 );
buf ( n42509 , n379847 );
and ( n42510 , n34885 , RI15b60990_1161);
and ( n42511 , n34887 , RI15b5d7e0_1055);
nor ( n42512 , n42510 , n42511 );
not ( n42513 , n42512 );
buf ( n42514 , n42513 );
buf ( n42515 , n380903 );
buf ( n42516 , n22007 );
buf ( n42517 , n18226 );
buf ( n42518 , n382069 );
not ( n42519 , n21723 );
not ( n42520 , n42519 );
nand ( n42521 , n40547 , n21652 );
not ( n42522 , n42521 );
nand ( n42523 , n42522 , n21674 );
not ( n42524 , n42523 );
or ( n42525 , n42520 , n42524 );
nand ( n42526 , n42525 , n21725 );
and ( n42527 , n42526 , n36689 );
not ( n42528 , n21319 );
not ( n42529 , n20696 );
and ( n42530 , n42528 , n42529 );
and ( n42531 , n21319 , n20696 );
nor ( n42532 , n42530 , n42531 );
not ( n42533 , n21360 );
or ( n42534 , n42532 , n42533 );
not ( n42535 , n21382 );
not ( n42536 , n21536 );
or ( n42537 , n42535 , n42536 );
or ( n42538 , n21536 , n21382 );
nand ( n42539 , n42537 , n42538 );
not ( n42540 , n22688 );
not ( n42541 , n42540 );
and ( n42542 , n42539 , n42541 );
nor ( n42543 , n21750 , n22614 );
nor ( n42544 , n42542 , n42543 );
nand ( n42545 , n42534 , n42544 );
nor ( n42546 , n42527 , n42545 );
and ( n42547 , n21788 , RI15b57048_834);
buf ( n42548 , n21770 );
and ( n42549 , n22507 , n42548 );
and ( n42550 , n17548 , n17549 );
not ( n42551 , n17548 );
and ( n42552 , n42551 , RI15b57048_834);
nor ( n42553 , n42550 , n42552 );
and ( n42554 , n42553 , n384127 );
nor ( n42555 , n42547 , n42549 , n42554 );
nand ( n42556 , n42546 , n42555 );
buf ( n42557 , n42556 );
not ( n42558 , n22490 );
nor ( n42559 , n42558 , n22498 );
and ( n42560 , n33292 , n42559 );
buf ( n42561 , n22609 );
or ( n42562 , n21922 , n42561 );
nand ( n42563 , n42562 , n21946 );
and ( n42564 , n42563 , RI15b57e58_864);
not ( n42565 , n21949 );
not ( n42566 , n22578 );
not ( n42567 , n42566 );
or ( n42568 , n42565 , n42567 );
nand ( n42569 , n42568 , n21979 );
and ( n42570 , n42569 , RI15b56058_800);
nor ( n42571 , n42564 , n42570 );
or ( n42572 , n42571 , n18078 );
and ( n42573 , n18188 , n42561 , n22610 );
or ( n42574 , n22601 , n42566 , RI15b56058_800);
and ( n42575 , n18177 , RI15b57e58_864);
and ( n42576 , n18219 , RI15b56f58_832);
nor ( n42577 , n42575 , n42576 , n21751 );
nand ( n42578 , n42574 , n42577 );
nor ( n42579 , n42573 , n42578 );
nand ( n42580 , n42572 , n42579 );
nor ( n42581 , n42560 , n42580 );
not ( n42582 , n17507 );
not ( n42583 , n42558 );
or ( n42584 , n42582 , n42583 );
nand ( n42585 , n42584 , n17565 );
nand ( n42586 , n42585 , n22498 );
nand ( n42587 , n42581 , n42586 );
buf ( n42588 , n42587 );
buf ( n42589 , n379844 );
buf ( n42590 , n22788 );
or ( n42591 , n31006 , n41443 );
and ( n42592 , n31016 , n41446 );
or ( n42593 , n41455 , n20979 );
or ( n42594 , n31022 , n41461 );
or ( n42595 , n41453 , n31024 );
nand ( n42596 , n42593 , n42594 , n42595 );
nor ( n42597 , n42592 , n42596 );
nand ( n42598 , n42591 , n42597 );
buf ( n42599 , n42598 );
buf ( n42600 , n19653 );
or ( n42601 , n41603 , n41606 );
and ( n42602 , n38654 , RI15b5b350_977);
buf ( n42603 , n39716 );
and ( n42604 , n42603 , RI15b5af90_969);
nor ( n42605 , n42602 , n42604 );
buf ( n42606 , n39720 );
and ( n42607 , n42606 , RI15b5abd0_961);
buf ( n42608 , n39723 );
and ( n42609 , n42608 , RI15b5a810_953);
nor ( n42610 , n42607 , n42609 );
buf ( n42611 , n39727 );
and ( n42612 , n42611 , RI15b5a450_945);
buf ( n42613 , n39730 );
and ( n42614 , n42613 , RI15b5a090_937);
nor ( n42615 , n42612 , n42614 );
buf ( n42616 , n39734 );
and ( n42617 , n42616 , RI15b59cd0_929);
buf ( n42618 , n39737 );
and ( n42619 , n42618 , RI15b59910_921);
nor ( n42620 , n42617 , n42619 );
nand ( n42621 , n42605 , n42610 , n42615 , n42620 );
and ( n42622 , n41935 , n42621 );
and ( n42623 , n39746 , RI15b58dd0_897);
and ( n42624 , n39751 , RI15b5c250_1009);
nor ( n42625 , n42622 , n42623 , n42624 );
and ( n42626 , n39756 , RI15b5be90_1001);
and ( n42627 , n39759 , RI15b5bad0_993);
nor ( n42628 , n42626 , n42627 );
and ( n42629 , n39763 , RI15b59550_913);
and ( n42630 , n39765 , RI15b59190_905);
nor ( n42631 , n42629 , n42630 );
and ( n42632 , n39769 , RI15b58a10_889);
and ( n42633 , n39772 , RI15b5b710_985);
nor ( n42634 , n42632 , n42633 );
nand ( n42635 , n42625 , n42628 , n42631 , n42634 );
and ( n42636 , n42635 , n31123 );
or ( n42637 , n41420 , n31079 , RI15b61728_1190);
not ( n42638 , n380632 );
or ( n42639 , n31052 , n42638 );
nand ( n42640 , n42637 , n42639 );
not ( n42641 , n384906 );
not ( n42642 , n381613 );
nor ( n42643 , n42641 , n42642 );
nor ( n42644 , n42636 , n42640 , n42643 );
nand ( n42645 , n42601 , n42644 );
buf ( n42646 , n42645 );
buf ( n42647 , n384218 );
buf ( n42648 , n31033 );
not ( n42649 , RI15b53ad8_720);
not ( n42650 , n32244 );
or ( n42651 , n42649 , n42650 );
and ( n42652 , n32247 , RI15b650d0_1313);
and ( n42653 , n32249 , RI15b5ff40_1139);
nor ( n42654 , n42652 , n42653 );
nand ( n42655 , n42651 , n42654 );
buf ( n42656 , n42655 );
buf ( n42657 , n19655 );
buf ( n42658 , n382049 );
or ( n42659 , n19988 , n381056 );
and ( n42660 , n35537 , RI15b43278_156);
and ( n42661 , n35373 , RI15b43638_164);
nor ( n42662 , n42660 , n42661 );
and ( n42663 , n35376 , RI15b439f8_172);
and ( n42664 , n35391 , RI15b42378_124);
and ( n42665 , n37302 , RI15b42738_132);
and ( n42666 , n35415 , RI15b42af8_140);
and ( n42667 , n35412 , RI15b41fb8_116);
nor ( n42668 , n42665 , n42666 , n42667 );
or ( n42669 , n35568 , n42668 );
or ( n42670 , n41531 , n20409 );
nand ( n42671 , n42669 , n42670 );
nor ( n42672 , n42664 , n42671 );
and ( n42673 , n35541 , RI15b41478_92);
and ( n42674 , n35546 , RI15b41bf8_108);
nor ( n42675 , n42673 , n42674 );
and ( n42676 , n35543 , RI15b410b8_84);
and ( n42677 , n35548 , RI15b41838_100);
nor ( n42678 , n42676 , n42677 );
nand ( n42679 , n42672 , n42675 , n42678 );
nor ( n42680 , n42663 , n42679 );
nand ( n42681 , n41517 , RI15b42eb8_148);
and ( n42682 , n41525 , RI15b40938_68);
and ( n42683 , n41523 , RI15b40cf8_76);
and ( n42684 , n41529 , RI15b40578_60);
nor ( n42685 , n42682 , n42683 , n42684 );
nand ( n42686 , n42662 , n42680 , n42681 , n42685 );
not ( n42687 , n42686 );
buf ( n42688 , n32807 );
or ( n42689 , n42687 , n42688 );
buf ( n42690 , n37110 );
and ( n42691 , n37125 , RI15b49dd0_385);
not ( n42692 , n37125 );
and ( n42693 , n42692 , n19988 );
nor ( n42694 , n42691 , n42693 );
or ( n42695 , n42690 , n42694 );
nand ( n42696 , n42659 , n42689 , n42695 );
buf ( n42697 , n42696 );
buf ( n42698 , n35651 );
buf ( n42699 , n19653 );
buf ( n42700 , n31996 );
nor ( n42701 , n31990 , n42700 );
not ( n42702 , n32009 );
nand ( n42703 , n42701 , n42702 );
nor ( n42704 , n42703 , n382079 );
or ( n42705 , n42704 , n32024 );
buf ( n42706 , n32001 );
nand ( n42707 , n42705 , n42706 );
not ( n42708 , n42703 );
not ( n42709 , n42708 );
nor ( n42710 , n32924 , n42706 );
and ( n42711 , n42709 , n42710 );
buf ( n42712 , n32039 );
not ( n42713 , n42712 );
not ( n42714 , n32010 );
and ( n42715 , n42713 , n42714 );
and ( n42716 , n42712 , n32010 );
nor ( n42717 , n42715 , n42716 );
or ( n42718 , n382513 , n42717 );
and ( n42719 , n382523 , RI15b4b720_439);
buf ( n42720 , n382529 );
and ( n42721 , n42720 , RI15b45528_230);
nor ( n42722 , n42719 , n42721 );
nand ( n42723 , n42718 , n42722 );
nor ( n42724 , n42711 , n42723 );
nand ( n42725 , n42707 , n42724 );
buf ( n42726 , n42725 );
buf ( n42727 , n22479 );
buf ( n42728 , n384218 );
buf ( n42729 , n384199 );
buf ( n42730 , n32160 );
buf ( n42731 , n32255 );
or ( n42732 , n22216 , RI15b4a2f8_396);
or ( n42733 , n30908 , n20637 );
nand ( n42734 , n42733 , RI15b4a2f8_396);
not ( n42735 , n39306 );
or ( n42736 , n386106 , RI15b43ae8_174);
or ( n42737 , n38458 , n386022 );
nand ( n42738 , n42736 , n42737 , n386112 );
not ( n42739 , n42738 );
or ( n42740 , n42735 , n42739 );
or ( n42741 , n42738 , n39306 );
nand ( n42742 , n42740 , n42741 );
and ( n42743 , n386258 , n42742 );
and ( n42744 , n22393 , RI15b4b1f8_428);
not ( n42745 , n39299 );
not ( n42746 , n42738 );
or ( n42747 , n42745 , n42746 );
or ( n42748 , n42738 , n39299 );
nand ( n42749 , n42747 , n42748 );
and ( n42750 , n386011 , n42749 );
nor ( n42751 , n42743 , n42744 , n42750 );
nand ( n42752 , n42732 , n42734 , n42751 );
buf ( n42753 , n42752 );
buf ( n42754 , n22479 );
not ( n42755 , RI15b535b0_709);
not ( n42756 , n32244 );
or ( n42757 , n42755 , n42756 );
and ( n42758 , n32247 , RI15b64ba8_1302);
and ( n42759 , n32249 , RI15b5fa18_1128);
nor ( n42760 , n42758 , n42759 );
nand ( n42761 , n42757 , n42760 );
buf ( n42762 , n42761 );
buf ( n42763 , n32981 );
buf ( n42764 , n31033 );
not ( n42765 , n383929 );
not ( n42766 , n42765 );
not ( n42767 , n40634 );
or ( n42768 , n42766 , n42767 );
and ( n42769 , n384022 , RI15b62268_1214);
not ( n42770 , RI15b62268_1214);
not ( n42771 , n38473 );
or ( n42772 , n42770 , n42771 );
or ( n42773 , n38473 , RI15b62268_1214);
nand ( n42774 , n42772 , n42773 );
and ( n42775 , n384025 , n42774 );
nor ( n42776 , n42769 , n42775 );
nand ( n42777 , n42768 , n42776 );
buf ( n42778 , n42777 );
buf ( n42779 , n383345 );
buf ( n42780 , RI15b5e8c0_1091);
or ( n42781 , n31006 , n384057 );
and ( n42782 , n31016 , n384169 );
or ( n42783 , n384182 , n20971 );
or ( n42784 , n31022 , n384190 );
or ( n42785 , n384180 , n31024 );
nand ( n42786 , n42783 , n42784 , n42785 );
nor ( n42787 , n42782 , n42786 );
nand ( n42788 , n42781 , n42787 );
buf ( n42789 , n42788 );
buf ( n42790 , n382073 );
not ( n42791 , RI15b53358_704);
not ( n42792 , n32244 );
or ( n42793 , n42791 , n42792 );
and ( n42794 , n32247 , RI15b64950_1297);
and ( n42795 , n32249 , RI15b5f7c0_1123);
nor ( n42796 , n42794 , n42795 );
nand ( n42797 , n42793 , n42796 );
buf ( n42798 , n42797 );
buf ( n42799 , n380942 );
buf ( n42800 , n20663 );
not ( n42801 , RI15b4a550_401);
not ( n42802 , n30908 );
or ( n42803 , n42801 , n42802 );
and ( n42804 , n22217 , n19756 );
buf ( n42805 , n19751 );
and ( n42806 , n42805 , n19662 );
not ( n42807 , n42805 );
and ( n42808 , n42807 , RI15b4a550_401);
nor ( n42809 , n42806 , n42808 );
and ( n42810 , n20637 , n42809 );
not ( n42811 , n386080 );
buf ( n42812 , n386125 );
not ( n42813 , n42812 );
not ( n42814 , n386129 );
and ( n42815 , n42813 , n42814 );
not ( n42816 , n386075 );
nor ( n42817 , n42815 , n42816 );
buf ( n42818 , n385768 );
or ( n42819 , n42817 , n42818 );
and ( n42820 , n42812 , n386075 );
nor ( n42821 , n42820 , n386129 );
not ( n42822 , n42818 );
or ( n42823 , n42821 , n42822 );
nand ( n42824 , n42819 , n42823 );
not ( n42825 , n42824 );
or ( n42826 , n42811 , n42825 );
or ( n42827 , n42824 , n386080 );
nand ( n42828 , n42826 , n42827 );
not ( n42829 , n386260 );
and ( n42830 , n42828 , n42829 );
not ( n42831 , n386358 );
not ( n42832 , n386314 );
not ( n42833 , n42832 );
nand ( n42834 , n42833 , n40186 );
buf ( n42835 , n386356 );
nand ( n42836 , n42834 , n42835 );
not ( n42837 , n42836 );
or ( n42838 , n42831 , n42837 );
nand ( n42839 , n42838 , n386345 );
not ( n42840 , n42839 );
not ( n42841 , n386343 );
nand ( n42842 , n42841 , n386348 );
not ( n42843 , n42842 );
and ( n42844 , n42840 , n42843 );
and ( n42845 , n42839 , n42842 );
nor ( n42846 , n42844 , n42845 );
nor ( n42847 , n42846 , n386499 );
nor ( n42848 , n42830 , n42847 );
and ( n42849 , n385769 , n385433 );
not ( n42850 , n42849 );
not ( n42851 , n385766 );
not ( n42852 , n42851 );
or ( n42853 , n42850 , n42852 );
or ( n42854 , n42851 , n42849 );
nand ( n42855 , n42853 , n42854 );
and ( n42856 , n42855 , n386015 );
and ( n42857 , n22395 , RI15b4b450_433);
nor ( n42858 , n42856 , n42857 );
nand ( n42859 , n42848 , n42858 );
nor ( n42860 , n42804 , n42810 , n42859 );
nand ( n42861 , n42803 , n42860 );
buf ( n42862 , n42861 );
buf ( n42863 , n387159 );
buf ( n42864 , n22738 );
buf ( n42865 , n22402 );
buf ( n42866 , n382049 );
not ( n42867 , n40998 );
or ( n42868 , n42867 , n41015 );
nand ( n42869 , n42868 , n41032 );
not ( n42870 , n35103 );
nand ( n42871 , n42869 , n42870 );
not ( n42872 , n42867 );
nor ( n42873 , n42872 , n42870 );
nand ( n42874 , n41578 , n42873 );
nand ( n42875 , n41582 , RI15b462c0_259);
nand ( n42876 , n42871 , n42874 , n42875 , n35463 );
buf ( n42877 , n42876 );
buf ( n42878 , n22343 );
buf ( n42879 , n36704 );
buf ( n42880 , n386762 );
buf ( n42881 , n35649 );
buf ( n42882 , n379895 );
buf ( n42883 , n380942 );
buf ( n42884 , n22508 );
nor ( n42885 , n42884 , n21763 );
and ( n42886 , n33292 , n42885 );
not ( n42887 , n22613 );
and ( n42888 , n18188 , n42887 );
nor ( n42889 , n42888 , n379916 );
or ( n42890 , n42889 , n22615 );
not ( n42891 , n18086 );
not ( n42892 , n22583 );
not ( n42893 , n42892 );
or ( n42894 , n42891 , n42893 );
nand ( n42895 , n42894 , n18104 );
and ( n42896 , n42895 , RI15b561c0_803);
or ( n42897 , n42887 , n22614 , RI15b57fc0_867);
or ( n42898 , n22615 , RI15b57f48_866);
nand ( n42899 , n42897 , n42898 );
and ( n42900 , n18188 , n42899 );
or ( n42901 , n42892 , n18197 , RI15b561c0_803);
and ( n42902 , n18177 , RI15b57fc0_867);
and ( n42903 , n18219 , RI15b570c0_835);
nor ( n42904 , n42902 , n42903 );
nand ( n42905 , n42901 , n42904 );
nor ( n42906 , n42896 , n42900 , n42905 );
nand ( n42907 , n42890 , n42906 );
nor ( n42908 , n42886 , n42907 );
nand ( n42909 , n42884 , n17507 );
not ( n42910 , n42909 );
not ( n42911 , n17565 );
or ( n42912 , n42910 , n42911 );
nand ( n42913 , n42912 , n21763 );
nand ( n42914 , n42908 , n42913 );
buf ( n42915 , n42914 );
and ( n42916 , n21788 , RI15b56ee0_831);
buf ( n42917 , n21769 );
and ( n42918 , n21919 , n42917 );
not ( n42919 , n21912 );
and ( n42920 , n42919 , n21916 );
not ( n42921 , n42919 );
and ( n42922 , n42921 , RI15b56ee0_831);
nor ( n42923 , n42920 , n42922 );
and ( n42924 , n42923 , n384127 );
nor ( n42925 , n42916 , n42918 , n42924 );
nand ( n42926 , n40572 , n42925 );
buf ( n42927 , n42926 );
buf ( n42928 , n30992 );
buf ( n42929 , n22009 );
not ( n42930 , n35869 );
not ( n42931 , n42930 );
not ( n42932 , n32129 );
or ( n42933 , n42931 , n42932 );
and ( n42934 , n39450 , RI15b40aa0_71);
or ( n42935 , n32141 , n35871 );
or ( n42936 , n32148 , n35888 );
or ( n42937 , n35882 , n32150 );
nand ( n42938 , n42935 , n42936 , n42937 );
nor ( n42939 , n42934 , n42938 );
nand ( n42940 , n42933 , n42939 );
buf ( n42941 , n42940 );
not ( n42942 , n384960 );
or ( n42943 , n42942 , n35895 );
and ( n42944 , n384983 , n39462 );
not ( n42945 , RI15b40578_60);
or ( n42946 , n35911 , n42945 );
or ( n42947 , n22022 , n35917 );
or ( n42948 , n35909 , n384988 );
nand ( n42949 , n42946 , n42947 , n42948 );
nor ( n42950 , n42944 , n42949 );
nand ( n42951 , n42943 , n42950 );
buf ( n42952 , n42951 );
buf ( n42953 , n381566 );
buf ( n42954 , n383498 );
or ( n42955 , n383180 , n36275 );
not ( n42956 , n36291 );
and ( n42957 , n42956 , RI15b5bff8_1004);
or ( n42958 , n383184 , n36281 );
not ( n42959 , n36296 );
and ( n42960 , n42959 , n41701 );
and ( n42961 , n40019 , n36294 );
nor ( n42962 , n42960 , n42961 );
nand ( n42963 , n42958 , n42962 );
nor ( n42964 , n42957 , n42963 );
nand ( n42965 , n42955 , n42964 );
buf ( n42966 , n42965 );
buf ( n42967 , n21800 );
buf ( n42968 , n22788 );
not ( n42969 , n381406 );
not ( n42970 , n33130 );
or ( n42971 , n42969 , n42970 );
nand ( n42972 , n381417 , n381331 );
nand ( n42973 , n36269 , n41689 );
and ( n42974 , n42972 , n42973 );
nand ( n42975 , n381486 , RI15b52ea8_694);
nand ( n42976 , n42971 , n42974 , n42975 );
buf ( n42977 , n42976 );
buf ( n42978 , n20665 );
or ( n42979 , n32430 , n42970 );
and ( n42980 , n386637 , RI15b54bb8_756);
and ( n42981 , n382885 , n37835 );
not ( n42982 , RI15b54bb8_756);
not ( n42983 , n382638 );
not ( n42984 , n42983 );
or ( n42985 , n42982 , n42984 );
or ( n42986 , n42983 , RI15b54bb8_756);
nand ( n42987 , n42985 , n42986 );
and ( n42988 , n37449 , n42987 );
nor ( n42989 , n42980 , n42981 , n42988 );
and ( n42990 , n42972 , n42989 );
nand ( n42991 , n42979 , n42990 );
buf ( n42992 , n42991 );
buf ( n42993 , n32271 );
not ( n42994 , n39891 );
not ( n42995 , n37629 );
or ( n42996 , n42994 , n42995 );
and ( n42997 , n37637 , n32070 );
not ( n42998 , RI15b5a2e8_942);
or ( n42999 , n32081 , n42998 );
buf ( n43000 , n37642 );
not ( n43001 , n43000 );
or ( n43002 , n43001 , n32086 );
or ( n43003 , n32079 , n37646 );
nand ( n43004 , n42999 , n43002 , n43003 );
nor ( n43005 , n42997 , n43004 );
nand ( n43006 , n42996 , n43005 );
buf ( n43007 , n43006 );
buf ( n43008 , n385112 );
buf ( n43009 , n385195 );
not ( n43010 , n34719 );
not ( n43011 , n22801 );
nor ( n43012 , n43010 , n43011 );
buf ( n43013 , n43012 );
buf ( n43014 , n384218 );
buf ( n43015 , n383345 );
not ( n43016 , n33220 );
not ( n43017 , n37629 );
or ( n43018 , n43016 , n43017 );
and ( n43019 , n37637 , n33226 );
or ( n43020 , n33237 , n18975 );
or ( n43021 , n37644 , n33241 );
or ( n43022 , n33235 , n37646 );
nand ( n43023 , n43020 , n43021 , n43022 );
nor ( n43024 , n43019 , n43023 );
nand ( n43025 , n43018 , n43024 );
buf ( n43026 , n43025 );
buf ( n43027 , n382071 );
buf ( n43028 , n32255 );
not ( n43029 , n31982 );
nor ( n43030 , n43029 , n382079 );
or ( n43031 , n43030 , n382475 );
nand ( n43032 , n43031 , n31988 );
nor ( n43033 , n382487 , n31988 );
nand ( n43034 , n43029 , n43033 );
not ( n43035 , n382512 );
or ( n43036 , n382514 , n382516 );
not ( n43037 , n43036 );
buf ( n43038 , n31992 );
not ( n43039 , n43038 );
and ( n43040 , n43037 , n43039 );
and ( n43041 , n43036 , n43038 );
nor ( n43042 , n43040 , n43041 );
not ( n43043 , n43042 );
and ( n43044 , n43035 , n43043 );
not ( n43045 , RI15b453c0_227);
not ( n43046 , n382528 );
or ( n43047 , n43045 , n43046 );
not ( n43048 , n382523 );
not ( n43049 , RI15b4b5b8_436);
or ( n43050 , n43048 , n43049 );
nand ( n43051 , n43047 , n43050 );
nor ( n43052 , n43044 , n43051 );
nand ( n43053 , n43034 , n43052 );
not ( n43054 , n43053 );
nand ( n43055 , n43032 , n43054 );
buf ( n43056 , n43055 );
buf ( n43057 , n382069 );
buf ( n43058 , n31030 );
nor ( n43059 , n41736 , n41744 );
or ( n43060 , n43059 , n33503 );
nor ( n43061 , n35512 , n33487 );
and ( n43062 , n41743 , n43061 );
not ( n43063 , n43062 );
or ( n43064 , RI15b61908_1194 , n43063 );
and ( n43065 , n36538 , n39918 );
nor ( n43066 , n42641 , n39333 );
nor ( n43067 , n31052 , n380468 );
nor ( n43068 , n43065 , n43066 , n43067 );
nand ( n43069 , n43060 , n43064 , n43068 );
buf ( n43070 , n43069 );
buf ( n43071 , n384199 );
not ( n43072 , n36259 );
not ( n43073 , n384726 );
or ( n43074 , n43072 , n43073 );
not ( n43075 , n36239 );
and ( n43076 , n35477 , n43075 );
or ( n43077 , n36250 , n20771 );
or ( n43078 , n40525 , n36254 );
or ( n43079 , n36248 , n384759 );
nand ( n43080 , n43077 , n43078 , n43079 );
nor ( n43081 , n43076 , n43080 );
nand ( n43082 , n43074 , n43081 );
buf ( n43083 , n43082 );
buf ( n43084 , n22408 );
buf ( n43085 , RI15b47670_301);
buf ( n43086 , n386760 );
buf ( n43087 , n380906 );
and ( n43088 , n32899 , n32037 , n42141 );
and ( n43089 , n32837 , n43088 );
not ( n43090 , n32855 );
nand ( n43091 , n43089 , n43090 );
not ( n43092 , n32852 );
nor ( n43093 , n43091 , n43092 );
buf ( n43094 , n43093 );
not ( n43095 , n43094 );
nor ( n43096 , n43095 , n382079 );
not ( n43097 , n32023 );
buf ( n43098 , n43097 );
buf ( n43099 , n43098 );
or ( n43100 , n43096 , n43099 );
nand ( n43101 , n43100 , n32884 );
buf ( n43102 , n43094 );
not ( n43103 , n43102 );
not ( n43104 , n32941 );
nor ( n43105 , n43104 , n32884 );
and ( n43106 , n43103 , n43105 );
buf ( n43107 , n382513 );
buf ( n43108 , n382378 );
not ( n43109 , n43108 );
not ( n43110 , n32885 );
and ( n43111 , n43109 , n43110 );
and ( n43112 , n43108 , n32885 );
nor ( n43113 , n43111 , n43112 );
or ( n43114 , n43107 , n43113 );
and ( n43115 , n382523 , RI15b4ba68_446);
buf ( n43116 , n382529 );
and ( n43117 , n43116 , RI15b45870_237);
nor ( n43118 , n43115 , n43117 );
nand ( n43119 , n43114 , n43118 );
nor ( n43120 , n43106 , n43119 );
nand ( n43121 , n43101 , n43120 );
buf ( n43122 , n43121 );
buf ( n43123 , n384996 );
buf ( n43124 , n382049 );
buf ( n43125 , n382073 );
buf ( n43126 , n19651 );
buf ( n43127 , n22005 );
not ( n43128 , n39317 );
not ( n43129 , n32129 );
or ( n43130 , n43128 , n43129 );
not ( n43131 , n37675 );
and ( n43132 , n43131 , RI15b428a0_135);
or ( n43133 , n32141 , n37665 );
or ( n43134 , n32148 , n37679 );
or ( n43135 , n37673 , n32150 );
nand ( n43136 , n43133 , n43134 , n43135 );
nor ( n43137 , n43132 , n43136 );
nand ( n43138 , n43130 , n43137 );
buf ( n43139 , n43138 );
buf ( n43140 , n383345 );
buf ( n43141 , n22406 );
buf ( n43142 , n20663 );
buf ( n43143 , n20665 );
and ( n43144 , n41645 , n41653 );
not ( n43145 , n43144 );
nor ( n43146 , n43145 , n41015 );
or ( n43147 , n43146 , n41033 );
not ( n43148 , n35063 );
nand ( n43149 , n43147 , n43148 );
and ( n43150 , n43145 , n41578 , n35063 );
not ( n43151 , RI15b46518_264);
not ( n43152 , n379832 );
or ( n43153 , n43151 , n43152 );
not ( n43154 , n382002 );
not ( n43155 , n381980 );
or ( n43156 , n43154 , n43155 );
or ( n43157 , n381980 , n382002 );
nand ( n43158 , n43156 , n43157 );
and ( n43159 , n35461 , n43158 );
and ( n43160 , n35459 , n381975 );
nor ( n43161 , n43159 , n43160 );
nand ( n43162 , n43153 , n43161 );
nor ( n43163 , n43150 , n43162 );
nand ( n43164 , n43149 , n43163 );
buf ( n43165 , n43164 );
buf ( n43166 , n32672 );
buf ( n43167 , n22740 );
buf ( n43168 , n380940 );
buf ( n43169 , n384996 );
buf ( n43170 , n380203 );
buf ( n43171 , RI15b47058_288);
not ( n43172 , n36306 );
not ( n43173 , n43172 );
not ( n43174 , n39319 );
or ( n43175 , n43173 , n43174 );
and ( n43176 , n33196 , n36309 );
not ( n43177 , RI15b41c70_109);
or ( n43178 , n36318 , n43177 );
or ( n43179 , n22241 , n36325 );
or ( n43180 , n36316 , n33201 );
nand ( n43181 , n43178 , n43179 , n43180 );
nor ( n43182 , n43176 , n43181 );
nand ( n43183 , n43175 , n43182 );
buf ( n43184 , n43183 );
buf ( n43185 , n384199 );
buf ( n43186 , n19651 );
nor ( n43187 , RI15b606c0_1155 , RI15b60b70_1165);
not ( n43188 , n43187 );
buf ( n43189 , n379405 );
not ( n43190 , n43189 );
or ( n43191 , n43188 , n43190 );
not ( n43192 , RI15b60af8_1164);
nand ( n43193 , n43192 , n43187 );
not ( n43194 , n43193 );
and ( n43195 , RI15b606c0_1155 , RI15b60af8_1164);
nor ( n43196 , n43195 , RI15b60b70_1165);
nand ( n43197 , n43196 , RI15b63ac8_1266);
not ( n43198 , n43197 );
or ( n43199 , n43194 , n43198 );
nand ( n43200 , n43199 , RI15b63a50_1265);
nand ( n43201 , n43191 , n43200 );
buf ( n43202 , n43201 );
not ( n43203 , n385002 );
not ( n43204 , n43203 );
not ( n43205 , n384726 );
or ( n43206 , n43204 , n43205 );
and ( n43207 , n35477 , n385006 );
or ( n43208 , n385019 , n380103 );
or ( n43209 , n40525 , n385023 );
or ( n43210 , n385017 , n384759 );
nand ( n43211 , n43208 , n43209 , n43210 );
nor ( n43212 , n43207 , n43211 );
nand ( n43213 , n43206 , n43212 );
buf ( n43214 , n43213 );
buf ( n43215 , n381004 );
buf ( n43216 , n22714 );
buf ( n43217 , n20665 );
buf ( n43218 , n383498 );
not ( n43219 , n33996 );
nand ( n43220 , n43219 , n36490 );
not ( n43221 , n34174 );
nor ( n43222 , n43220 , n43221 );
nand ( n43223 , n43222 , n379785 );
not ( n43224 , n43223 );
not ( n43225 , n39798 );
or ( n43226 , n43224 , n43225 );
buf ( n43227 , n34188 );
nand ( n43228 , n43226 , n43227 );
not ( n43229 , n34250 );
not ( n43230 , n43222 );
not ( n43231 , n43227 );
nand ( n43232 , n43229 , n43230 , n43231 );
buf ( n43233 , n34616 );
not ( n43234 , n43233 );
buf ( n43235 , n34598 );
not ( n43236 , n43235 );
not ( n43237 , n43236 );
or ( n43238 , n43234 , n43237 );
or ( n43239 , n43236 , n43233 );
nand ( n43240 , n43238 , n43239 );
buf ( n43241 , n34645 );
not ( n43242 , n43241 );
nand ( n43243 , n43240 , n43242 );
and ( n43244 , n379783 , RI15b64680_1291);
and ( n43245 , n34651 , RI15b5e488_1082);
nor ( n43246 , n43244 , n43245 );
nand ( n43247 , n43228 , n43232 , n43243 , n43246 );
buf ( n43248 , n43247 );
not ( n43249 , n381769 );
and ( n43250 , n33624 , n381772 );
not ( n43251 , n43250 );
or ( n43252 , n43249 , n43251 );
or ( n43253 , n43250 , n381769 );
nand ( n43254 , n43252 , n43253 );
and ( n43255 , n43254 , n33631 );
not ( n43256 , n381742 );
nand ( n43257 , n43256 , n33633 );
and ( n43258 , n43257 , n381737 );
not ( n43259 , n43257 );
and ( n43260 , n43259 , n381736 );
nor ( n43261 , n43258 , n43260 );
or ( n43262 , n43261 , n37981 );
not ( n43263 , n381799 );
or ( n43264 , n43263 , n381803 );
not ( n43265 , n381805 );
nand ( n43266 , n43264 , n43265 );
buf ( n43267 , n21748 );
and ( n43268 , n43266 , n43267 );
and ( n43269 , n21751 , RI15b580b0_869);
nor ( n43270 , n43268 , n43269 );
nand ( n43271 , n43262 , n43270 );
nor ( n43272 , n43255 , n43271 );
and ( n43273 , n385164 , RI15b50a18_616);
or ( n43274 , n33652 , n381803 );
or ( n43275 , n381769 , n385170 );
or ( n43276 , n381736 , n385178 );
nand ( n43277 , n43274 , n43275 , n43276 );
nor ( n43278 , n43273 , n43277 );
nand ( n43279 , n43272 , n43278 );
buf ( n43280 , n43279 );
not ( n43281 , n32680 );
not ( n43282 , n33400 );
or ( n43283 , n43281 , n43282 );
and ( n43284 , n33415 , n35222 );
or ( n43285 , n32692 , n18468 );
or ( n43286 , n36293 , n32699 );
or ( n43287 , n32690 , n33443 );
nand ( n43288 , n43285 , n43286 , n43287 );
nor ( n43289 , n43284 , n43288 );
nand ( n43290 , n43283 , n43289 );
buf ( n43291 , n43290 );
buf ( n43292 , n383174 );
not ( n43293 , n40674 );
nand ( n43294 , n379340 , RI15b54780_747);
nand ( n43295 , n43293 , n43294 );
and ( n43296 , n43295 , RI15b54708_746);
buf ( n43297 , n43296 );
buf ( n43298 , n20665 );
buf ( n43299 , n385112 );
buf ( n43300 , n22005 );
or ( n43301 , n40833 , n18078 );
and ( n43302 , n39220 , RI15b50e50_625);
and ( n43303 , n383915 , n20731 );
and ( n43304 , n32986 , n21402 );
nor ( n43305 , n43302 , n43303 , n43304 );
nand ( n43306 , n43301 , n43305 );
buf ( n43307 , n43306 );
nor ( n43308 , n39806 , n39808 );
buf ( n43309 , n34480 );
nand ( n43310 , n43308 , n43309 );
buf ( n43311 , n43310 );
buf ( n43312 , n34434 );
not ( n43313 , n43312 );
xor ( n43314 , n43311 , n43313 );
not ( n43315 , n39814 );
or ( n43316 , n43314 , n43315 );
not ( n43317 , n36494 );
and ( n43318 , n36566 , n379785 );
nor ( n43319 , n43317 , n43318 );
not ( n43320 , n43319 );
not ( n43321 , n34122 );
not ( n43322 , n43321 );
and ( n43323 , n43320 , n43322 );
not ( n43324 , n36566 );
nand ( n43325 , n43324 , n43321 );
or ( n43326 , n36501 , n43325 );
and ( n43327 , n379783 , RI15b64248_1282);
and ( n43328 , n34651 , RI15b5e050_1073);
nor ( n43329 , n43327 , n43328 );
nand ( n43330 , n43326 , n43329 );
nor ( n43331 , n43323 , n43330 );
nand ( n43332 , n43316 , n43331 );
buf ( n43333 , n43332 );
buf ( n43334 , n17499 );
not ( n43335 , n39134 );
not ( n43336 , n32129 );
or ( n43337 , n43335 , n43336 );
not ( n43338 , n38077 );
and ( n43339 , n43338 , RI15b42c60_143);
or ( n43340 , n32141 , n38069 );
or ( n43341 , n32148 , n38081 );
or ( n43342 , n38075 , n32150 );
nand ( n43343 , n43340 , n43341 , n43342 );
nor ( n43344 , n43339 , n43343 );
nand ( n43345 , n43337 , n43344 );
buf ( n43346 , n43345 );
buf ( n43347 , n22005 );
buf ( n43348 , n379403 );
buf ( n43349 , RI15b3e9d0_1);
buf ( n43350 , n43349 );
buf ( n43351 , n19651 );
buf ( n43352 , n382069 );
buf ( n43353 , n17499 );
buf ( n43354 , n382073 );
or ( n43355 , n381907 , n36813 );
and ( n43356 , n36825 , RI15b42198_120);
or ( n43357 , n381917 , n36815 );
not ( n43358 , n36830 );
and ( n43359 , n43358 , n381923 );
and ( n43360 , n381926 , n36828 );
nor ( n43361 , n43359 , n43360 );
nand ( n43362 , n43357 , n43361 );
nor ( n43363 , n43356 , n43362 );
nand ( n43364 , n43355 , n43363 );
buf ( n43365 , n43364 );
buf ( n43366 , n383174 );
buf ( n43367 , n31979 );
buf ( n43368 , n17499 );
or ( n43369 , n31006 , n386706 );
and ( n43370 , n31016 , n386718 );
or ( n43371 , n386727 , n20976 );
or ( n43372 , n34893 , n386735 );
or ( n43373 , n386725 , n31024 );
nand ( n43374 , n43371 , n43372 , n43373 );
nor ( n43375 , n43370 , n43374 );
nand ( n43376 , n43369 , n43375 );
buf ( n43377 , n43376 );
and ( n43378 , n22646 , RI15b45d98_248);
and ( n43379 , n22648 , RI15b52200_667);
nor ( n43380 , n43378 , n43379 );
not ( n43381 , n43380 );
buf ( n43382 , n43381 );
or ( n43383 , n384021 , n386961 );
or ( n43384 , n18732 , n386747 );
not ( n43385 , n384032 );
and ( n43386 , n43385 , RI15b61ea8_1206);
not ( n43387 , n43385 );
and ( n43388 , n43387 , n386961 );
nor ( n43389 , n43386 , n43388 );
or ( n43390 , n43389 , n384024 );
nand ( n43391 , n43383 , n43384 , n43390 );
buf ( n43392 , n43391 );
buf ( n43393 , n384199 );
buf ( n43394 , n380906 );
buf ( n43395 , n383345 );
not ( n43396 , n386706 );
not ( n43397 , n43396 );
not ( n43398 , n384726 );
or ( n43399 , n43397 , n43398 );
and ( n43400 , n384737 , n386718 );
or ( n43401 , n386727 , n20837 );
or ( n43402 , n40525 , n386735 );
or ( n43403 , n386725 , n384759 );
nand ( n43404 , n43401 , n43402 , n43403 );
nor ( n43405 , n43400 , n43404 );
nand ( n43406 , n43399 , n43405 );
buf ( n43407 , n43406 );
buf ( n43408 , RI15b5dfd8_1072);
buf ( n43409 , n22714 );
and ( n43410 , n384022 , RI15b61cc8_1202);
and ( n43411 , n386746 , RI15b58830_885);
and ( n43412 , RI15b61cc8_1202 , RI15b61c50_1201);
not ( n43413 , RI15b61cc8_1202);
and ( n43414 , n43413 , n36228 );
nor ( n43415 , n43412 , n43414 );
and ( n43416 , n384025 , n43415 );
nor ( n43417 , n43410 , n43411 , n43416 );
not ( n43418 , n43417 );
buf ( n43419 , n43418 );
nor ( n43420 , n33257 , n33255 );
nand ( n43421 , n43420 , n32909 );
not ( n43422 , n43421 );
or ( n43423 , n43422 , n32958 );
not ( n43424 , n32919 );
nand ( n43425 , n43423 , n43424 );
not ( n43426 , n32919 );
not ( n43427 , n32036 );
not ( n43428 , n32913 );
or ( n43429 , n43427 , n43428 );
nand ( n43430 , n43429 , n33254 );
not ( n43431 , n43430 );
or ( n43432 , n43426 , n43431 );
not ( n43433 , n382513 );
not ( n43434 , n32920 );
not ( n43435 , n43434 );
not ( n43436 , n382497 );
or ( n43437 , n43435 , n43436 );
or ( n43438 , n382497 , n43434 );
nand ( n43439 , n43437 , n43438 );
and ( n43440 , n43433 , n43439 );
and ( n43441 , n382523 , RI15b4bdb0_453);
and ( n43442 , n42153 , RI15b45bb8_244);
nor ( n43443 , n43441 , n43442 );
not ( n43444 , n43443 );
nor ( n43445 , n43440 , n43444 );
nand ( n43446 , n43432 , n43445 );
not ( n43447 , n43446 );
nand ( n43448 , n43425 , n43447 );
buf ( n43449 , n43448 );
buf ( n43450 , n22009 );
buf ( n43451 , n384199 );
buf ( n43452 , n33250 );
buf ( n43453 , n386762 );
or ( n43454 , n381056 , n19960 );
or ( n43455 , n36988 , n381062 );
not ( n43456 , n32813 );
and ( n43457 , n43456 , RI15b495d8_368);
not ( n43458 , n43456 );
and ( n43459 , n43458 , n19960 );
nor ( n43460 , n43457 , n43459 );
not ( n43461 , n36064 );
or ( n43462 , n43460 , n43461 );
nand ( n43463 , n43454 , n43455 , n43462 );
buf ( n43464 , n43463 );
buf ( n43465 , n382049 );
buf ( n43466 , n382073 );
or ( n43467 , n381015 , n379836 );
nand ( n43468 , n35525 , RI15b533d0_705);
nand ( n43469 , n43467 , n43468 );
buf ( n43470 , n43469 );
buf ( n43471 , n32160 );
buf ( n43472 , n19655 );
buf ( n43473 , n380940 );
not ( n43474 , n31572 );
not ( n43475 , n43474 );
buf ( n43476 , n31566 );
not ( n43477 , n43476 );
or ( n43478 , n43475 , n43477 );
or ( n43479 , n43476 , n43474 );
nand ( n43480 , n43478 , n43479 );
nand ( n43481 , n43480 , n31599 );
nand ( n43482 , n42050 , n379218 );
nand ( n43483 , n43482 , n31700 );
not ( n43484 , n379206 );
nand ( n43485 , n43483 , n43484 );
not ( n43486 , n31330 );
not ( n43487 , n31706 );
or ( n43488 , n43486 , n43487 );
nand ( n43489 , n43488 , n42053 );
nand ( n43490 , n43489 , n379206 );
and ( n43491 , n379394 , RI15b57ed0_865);
and ( n43492 , n31712 , RI15b51cd8_656);
nor ( n43493 , n43491 , n43492 );
nand ( n43494 , n43481 , n43485 , n43490 , n43493 );
buf ( n43495 , n43494 );
buf ( n43496 , n35649 );
and ( n43497 , n31792 , n31928 );
or ( n43498 , n31916 , n42117 );
or ( n43499 , n31771 , n31925 );
or ( n43500 , n31779 , n31876 );
nand ( n43501 , n43498 , n43499 , n43500 );
nor ( n43502 , n43497 , n43501 );
nand ( n43503 , n31963 , n43502 );
buf ( n43504 , n43503 );
buf ( n43505 , n382537 );
buf ( n43506 , n33250 );
buf ( n43507 , n31033 );
or ( n43508 , n385219 , RI15b3fa38_36);
nor ( n43509 , n382076 , RI15b48390_329 , RI15b47e68_318);
and ( n43510 , n43509 , RI15b3f9c0_35);
or ( n43511 , RI15b3f9c0_35 , RI15b47e68_318);
nand ( n43512 , n43511 , n35241 , RI15b48318_328);
and ( n43513 , n43512 , n382078 );
nand ( n43514 , n20492 , RI15b48390_329);
nor ( n43515 , n43513 , n43514 );
nand ( n43516 , RI15b3f9c0_35 , RI15b48408_330);
nor ( n43517 , n385218 , n43516 );
nor ( n43518 , n43510 , n43515 , n43517 );
nand ( n43519 , n43508 , n43518 , n382079 );
buf ( n43520 , n43519 );
buf ( n43521 , n386762 );
not ( n43522 , n380235 );
not ( n43523 , n381589 );
or ( n43524 , n43522 , n43523 );
and ( n43525 , n381596 , n380745 );
or ( n43526 , n380776 , n18732 );
or ( n43527 , n381616 , n380785 );
or ( n43528 , n380768 , n381621 );
nand ( n43529 , n43526 , n43527 , n43528 );
nor ( n43530 , n43525 , n43529 );
nand ( n43531 , n43524 , n43530 );
buf ( n43532 , n43531 );
not ( n43533 , n40334 );
not ( n43534 , RI15b56490_809);
and ( n43535 , n43533 , n43534 );
not ( n43536 , n43533 );
and ( n43537 , n43536 , RI15b56490_809);
nor ( n43538 , n43535 , n43537 );
nand ( n43539 , n43538 , n379949 );
and ( n43540 , n380000 , RI15b56490_809);
not ( n43541 , n382745 );
not ( n43542 , n382785 );
and ( n43543 , n43541 , n43542 );
and ( n43544 , n382745 , n382785 );
nor ( n43545 , n43543 , n43544 );
not ( n43546 , n43545 );
and ( n43547 , n380012 , n43546 );
nor ( n43548 , n43540 , n43547 );
nand ( n43549 , n43539 , n43548 );
buf ( n43550 , n43549 );
buf ( n43551 , n379847 );
buf ( n43552 , RI15b5e230_1077);
buf ( n43553 , n22005 );
buf ( n43554 , n19655 );
buf ( n43555 , n19653 );
buf ( n43556 , n385112 );
not ( n43557 , n35478 );
and ( n43558 , n383871 , n43557 );
nor ( n43559 , n43558 , n35479 );
not ( n43560 , n21776 );
or ( n43561 , n43559 , n43560 );
not ( n43562 , n21765 );
or ( n43563 , n43562 , n383841 );
and ( n43564 , n36845 , RI15b4c260_463);
and ( n43565 , n383915 , n383823 );
nor ( n43566 , n43564 , n43565 );
nand ( n43567 , n43561 , n43563 , n43566 );
buf ( n43568 , n43567 );
buf ( n43569 , n386760 );
buf ( n43570 , n387159 );
or ( n43571 , n19607 , n383476 );
and ( n43572 , n19630 , n383480 );
and ( n43573 , n19644 , n383476 );
not ( n43574 , n19338 );
nand ( n43575 , n19421 , n19434 );
not ( n43576 , n43575 );
not ( n43577 , n43576 );
and ( n43578 , n43574 , n43577 );
and ( n43579 , n19338 , n43576 );
nor ( n43580 , n43578 , n43579 );
or ( n43581 , n19388 , n43580 );
and ( n43582 , n18670 , n18591 );
not ( n43583 , n18669 );
or ( n43584 , n43583 , n18667 );
nand ( n43585 , n43584 , n18632 );
and ( n43586 , n43585 , n18590 );
nor ( n43587 , n43582 , n43586 );
not ( n43588 , n43587 );
not ( n43589 , n18595 );
and ( n43590 , n43588 , n43589 );
and ( n43591 , n43587 , n18595 );
nor ( n43592 , n43590 , n43591 );
or ( n43593 , n19283 , n43592 );
not ( n43594 , n43575 );
not ( n43595 , n19431 );
or ( n43596 , n43594 , n43595 );
or ( n43597 , n19431 , n43575 );
nand ( n43598 , n43596 , n43597 );
and ( n43599 , n43598 , n19498 );
and ( n43600 , n19513 , RI15b63b40_1267);
nor ( n43601 , n43599 , n43600 );
nand ( n43602 , n43581 , n43593 , n43601 );
nor ( n43603 , n43572 , n43573 , n43602 );
nand ( n43604 , n43571 , n43603 );
buf ( n43605 , n43604 );
or ( n43606 , n36937 , n33111 );
and ( n43607 , n36946 , n33117 );
or ( n43608 , n33128 , n17819 );
or ( n43609 , n39875 , n33134 );
or ( n43610 , n33126 , n36955 );
nand ( n43611 , n43608 , n43609 , n43610 );
nor ( n43612 , n43607 , n43611 );
nand ( n43613 , n43606 , n43612 );
buf ( n43614 , n43613 );
buf ( n43615 , n381566 );
and ( n43616 , n383607 , n22428 );
nor ( n43617 , n43616 , n383413 , n383596 );
or ( n43618 , n43617 , n385033 );
not ( n43619 , n31757 );
not ( n43620 , n383501 );
or ( n43621 , n43619 , n43620 );
not ( n43622 , n31756 );
nand ( n43623 , n43621 , n43622 );
and ( n43624 , n43623 , n22462 );
not ( n43625 , n31757 );
not ( n43626 , n19627 );
and ( n43627 , n43625 , n43626 );
nor ( n43628 , n43627 , n384921 );
nor ( n43629 , n43624 , n43628 , n383595 );
nand ( n43630 , n43618 , n43629 );
buf ( n43631 , n43630 );
buf ( n43632 , n380203 );
buf ( n43633 , n22714 );
buf ( n43634 , n381566 );
buf ( n43635 , n31979 );
or ( n43636 , n36747 , n20519 );
not ( n43637 , RI15b44ad8_208);
or ( n43638 , n39256 , n43637 );
or ( n43639 , n37049 , n22298 );
and ( n43640 , n386110 , RI15b44970_205);
not ( n43641 , RI15b44970_205);
and ( n43642 , n386066 , n43641 );
nor ( n43643 , n43640 , n43642 );
or ( n43644 , n43643 , n36114 );
nand ( n43645 , n43638 , n43639 , n43644 );
not ( n43646 , n43645 );
nand ( n43647 , n43636 , n43646 );
buf ( n43648 , n43647 );
buf ( n43649 , n35651 );
buf ( n43650 , n32676 );
buf ( n43651 , n22005 );
buf ( n43652 , n380940 );
or ( n43653 , n383180 , n386591 );
not ( n43654 , n386612 );
and ( n43655 , n43654 , RI15b59e38_932);
or ( n43656 , n383184 , n386602 );
and ( n43657 , n386623 , n41701 );
and ( n43658 , n40019 , n386620 );
nor ( n43659 , n43657 , n43658 );
nand ( n43660 , n43656 , n43659 );
nor ( n43661 , n43655 , n43660 );
nand ( n43662 , n43653 , n43661 );
buf ( n43663 , n43662 );
or ( n43664 , n382679 , n383016 );
and ( n43665 , n35732 , RI15b4c710_473);
and ( n43666 , n35734 , RI15b4fb90_585);
and ( n43667 , n380061 , RI15b4ec90_553);
and ( n43668 , n382793 , RI15b4d9d0_513);
and ( n43669 , n35739 , RI15b4d250_497);
nor ( n43670 , n43667 , n43668 , n43669 );
not ( n43671 , n41895 );
and ( n43672 , n43671 , RI15b4dd90_521);
and ( n43673 , n382806 , RI15b4e8d0_545);
nor ( n43674 , n43672 , n43673 );
and ( n43675 , n382780 , RI15b4d610_505);
and ( n43676 , n382801 , RI15b4e510_537);
nor ( n43677 , n43675 , n43676 );
nand ( n43678 , n35748 , RI15b4e150_529);
nand ( n43679 , n43670 , n43674 , n43677 , n43678 );
and ( n43680 , n379991 , n43679 );
nor ( n43681 , n43665 , n43666 , n43680 );
and ( n43682 , n35754 , RI15b4f410_569);
and ( n43683 , n35756 , RI15b4f7d0_577);
nor ( n43684 , n43682 , n43683 );
and ( n43685 , n35759 , RI15b4f050_561);
and ( n43686 , n35761 , RI15b4c350_465);
nor ( n43687 , n43685 , n43686 );
and ( n43688 , n35764 , RI15b4ce90_489);
and ( n43689 , n35766 , RI15b4cad0_481);
nor ( n43690 , n43688 , n43689 );
nand ( n43691 , n43681 , n43684 , n43687 , n43690 );
and ( n43692 , n43691 , n35729 );
or ( n43693 , n382691 , n383700 );
not ( n43694 , n382652 );
and ( n43695 , n43694 , RI15b55068_766);
not ( n43696 , n43694 );
and ( n43697 , n43696 , n383016 );
nor ( n43698 , n43695 , n43697 );
not ( n43699 , n382624 );
or ( n43700 , n43698 , n43699 );
nand ( n43701 , n43693 , n43700 , n41857 );
nor ( n43702 , n43692 , n43701 );
nand ( n43703 , n43664 , n43702 );
buf ( n43704 , n43703 );
buf ( n43705 , n383345 );
not ( n43706 , RI15b53880_715);
not ( n43707 , n383170 );
or ( n43708 , n43706 , n43707 );
not ( n43709 , n40054 );
not ( n43710 , n33453 );
or ( n43711 , n43709 , n43710 );
nand ( n43712 , n43711 , n33465 );
and ( n43713 , n43712 , n40052 );
nor ( n43714 , n40054 , n40052 );
and ( n43715 , n33476 , n43714 );
and ( n43716 , n383147 , RI15b53100_699);
nor ( n43717 , n43713 , n43715 , n43716 );
nand ( n43718 , n43708 , n43717 );
buf ( n43719 , n43718 );
buf ( n43720 , n380940 );
buf ( n43721 , n384203 );
not ( n43722 , n33387 );
not ( n43723 , n382912 );
or ( n43724 , n43722 , n43723 );
and ( n43725 , n382931 , n33417 );
not ( n43726 , RI15b5b620_983);
or ( n43727 , n33428 , n43726 );
or ( n43728 , n35163 , n33440 );
or ( n43729 , n33426 , n382967 );
nand ( n43730 , n43727 , n43728 , n43729 );
nor ( n43731 , n43725 , n43730 );
nand ( n43732 , n43724 , n43731 );
buf ( n43733 , n43732 );
buf ( n43734 , n22740 );
buf ( n43735 , n33382 );
buf ( n43736 , n379893 );
buf ( n43737 , n21800 );
or ( n43738 , n32525 , n386534 );
nand ( n43739 , n43738 , RI15b47f58_320);
nand ( n43740 , n43739 , n41015 , n37559 );
buf ( n43741 , n43740 );
buf ( n43742 , n386812 );
or ( n43743 , n43742 , n22473 );
nand ( n43744 , n43743 , n383474 );
nand ( n43745 , n43744 , n382612 );
not ( n43746 , n382612 );
nand ( n43747 , n43746 , n37068 , n43742 );
not ( n43748 , n34815 );
buf ( n43749 , n386962 );
and ( n43750 , n43748 , n43749 );
nor ( n43751 , n43750 , n40140 );
or ( n43752 , n43751 , n386963 );
and ( n43753 , n40145 , RI15b63d20_1271);
or ( n43754 , n34826 , n43749 , RI15b61f20_1207);
not ( n43755 , n387023 );
not ( n43756 , RI15b63d20_1271);
and ( n43757 , n43755 , n43756 );
and ( n43758 , n387023 , RI15b63d20_1271);
nor ( n43759 , n43757 , n43758 );
or ( n43760 , n34833 , n43759 );
nand ( n43761 , n43754 , n43760 );
nor ( n43762 , n43753 , n43761 );
nand ( n43763 , n43752 , n43762 );
nand ( n43764 , n43763 , n19201 );
and ( n43765 , n22423 , RI15b63d20_1271);
and ( n43766 , n19599 , RI15b62e20_1239);
nor ( n43767 , n43765 , n43766 , n19513 );
nand ( n43768 , n43745 , n43747 , n43764 , n43767 );
buf ( n43769 , n43768 );
buf ( n43770 , n386762 );
buf ( n43771 , n35649 );
and ( n43772 , n22646 , RI15b45528_230);
and ( n43773 , n22648 , RI15b51990_649);
nor ( n43774 , n43772 , n43773 );
not ( n43775 , n43774 );
buf ( n43776 , n43775 );
buf ( n43777 , n382073 );
or ( n43778 , n20641 , n20568 );
nand ( n43779 , n43778 , RI15b4b180_427);
not ( n43780 , n20520 );
nand ( n43781 , n43780 , n20502 );
and ( n43782 , n43781 , RI15b49380_363);
or ( n43783 , n37048 , RI15b449e8_206);
not ( n43784 , n19934 );
or ( n43785 , n43784 , n20654 );
nand ( n43786 , n43785 , RI15b4a280_395);
nand ( n43787 , n43783 , n43786 );
nor ( n43788 , n43782 , n43787 );
nand ( n43789 , n43779 , n43788 );
buf ( n43790 , n43789 );
buf ( n43791 , n381081 );
buf ( n43792 , n383174 );
or ( n43793 , n386705 , n41443 );
and ( n43794 , n386716 , n41446 );
not ( n43795 , RI15b4d7f0_509);
or ( n43796 , n41455 , n43795 );
or ( n43797 , n386732 , n41461 );
or ( n43798 , n41453 , n386738 );
nand ( n43799 , n43796 , n43797 , n43798 );
nor ( n43800 , n43794 , n43799 );
nand ( n43801 , n43793 , n43800 );
buf ( n43802 , n43801 );
buf ( n43803 , n19653 );
or ( n43804 , n31091 , n32329 );
and ( n43805 , n38654 , RI15b5b2d8_976);
and ( n43806 , n39716 , RI15b5af18_968);
nor ( n43807 , n43805 , n43806 );
and ( n43808 , n39720 , RI15b5ab58_960);
and ( n43809 , n39723 , RI15b5a798_952);
nor ( n43810 , n43808 , n43809 );
and ( n43811 , n39727 , RI15b5a3d8_944);
and ( n43812 , n39730 , RI15b5a018_936);
nor ( n43813 , n43811 , n43812 );
and ( n43814 , n39734 , RI15b59c58_928);
and ( n43815 , n39737 , RI15b59898_920);
nor ( n43816 , n43814 , n43815 );
nand ( n43817 , n43807 , n43810 , n43813 , n43816 );
and ( n43818 , n383967 , n43817 );
and ( n43819 , n39746 , RI15b58d58_896);
and ( n43820 , n39751 , RI15b5c1d8_1008);
nor ( n43821 , n43818 , n43819 , n43820 );
and ( n43822 , n39756 , RI15b5be18_1000);
and ( n43823 , n39759 , RI15b5ba58_992);
nor ( n43824 , n43822 , n43823 );
and ( n43825 , n39763 , RI15b594d8_912);
and ( n43826 , n39765 , RI15b59118_904);
nor ( n43827 , n43825 , n43826 );
and ( n43828 , n39769 , RI15b58998_888);
and ( n43829 , n39772 , RI15b5b698_984);
nor ( n43830 , n43828 , n43829 );
nand ( n43831 , n43821 , n43824 , n43827 , n43830 );
and ( n43832 , n43831 , n31121 );
or ( n43833 , n31052 , n380630 );
and ( n43834 , n41418 , RI15b616b0_1189);
not ( n43835 , n41418 );
and ( n43836 , n43835 , n32329 );
nor ( n43837 , n43834 , n43836 );
not ( n43838 , n31078 );
or ( n43839 , n43837 , n43838 );
nand ( n43840 , n43833 , n43839 );
not ( n43841 , n33431 );
nor ( n43842 , n42641 , n43841 );
nor ( n43843 , n43832 , n43840 , n43842 );
nand ( n43844 , n43804 , n43843 );
buf ( n43845 , n43844 );
buf ( n43846 , n33382 );
buf ( n43847 , n383498 );
buf ( n43848 , n383613 );
or ( n43849 , n382679 , n382657 );
and ( n43850 , n380061 , RI15b4edf8_556);
and ( n43851 , n382836 , RI15b4def8_524);
and ( n43852 , n380115 , RI15b4c4b8_468);
nor ( n43853 , n43850 , n43851 , n43852 );
and ( n43854 , n35739 , RI15b4d3b8_500);
or ( n43855 , n382800 , n21013 );
or ( n43856 , n17716 , n382812 );
and ( n43857 , n382758 , RI15b4ea38_548);
and ( n43858 , n379876 , RI15b4cc38_484);
nor ( n43859 , n43857 , n43858 );
nand ( n43860 , n43855 , n43856 , n43859 );
nor ( n43861 , n43854 , n43860 );
and ( n43862 , n382841 , RI15b4db38_516);
and ( n43863 , n382788 , RI15b4cff8_492);
and ( n43864 , n382824 , RI15b4d778_508);
nor ( n43865 , n43862 , n43863 , n43864 );
nand ( n43866 , n35748 , RI15b4e2b8_532);
nand ( n43867 , n43853 , n43861 , n43865 , n43866 );
and ( n43868 , n35736 , n43867 );
and ( n43869 , n35759 , RI15b4f1b8_564);
and ( n43870 , n35734 , RI15b4fcf8_588);
nor ( n43871 , n43868 , n43869 , n43870 );
and ( n43872 , n35754 , RI15b4f578_572);
and ( n43873 , n35756 , RI15b4f938_580);
nor ( n43874 , n43872 , n43873 );
nand ( n43875 , n43871 , n43874 );
and ( n43876 , n43875 , n386667 );
or ( n43877 , n382691 , n383637 );
and ( n43878 , n382656 , RI15b551d0_769);
not ( n43879 , n382656 );
and ( n43880 , n43879 , n382657 );
nor ( n43881 , n43878 , n43880 );
or ( n43882 , n43881 , n43699 );
nand ( n43883 , n43877 , n43882 );
nor ( n43884 , n381400 , n31019 );
nor ( n43885 , n43876 , n43883 , n43884 );
nand ( n43886 , n43849 , n43885 );
buf ( n43887 , n43886 );
not ( n43888 , n35784 );
not ( n43889 , n381589 );
or ( n43890 , n43888 , n43889 );
and ( n43891 , n381596 , n35790 );
not ( n43892 , RI15b59cd0_929);
or ( n43893 , n35803 , n43892 );
or ( n43894 , n381616 , n35811 );
or ( n43895 , n35801 , n381621 );
nand ( n43896 , n43893 , n43894 , n43895 );
nor ( n43897 , n43891 , n43896 );
nand ( n43898 , n43890 , n43897 );
buf ( n43899 , n43898 );
buf ( n43900 , n20665 );
not ( n43901 , RI15b55c20_791);
not ( n43902 , n380000 );
or ( n43903 , n43901 , n43902 );
and ( n43904 , n381636 , RI15b4e948_546);
and ( n43905 , n381639 , RI15b4e588_538);
nor ( n43906 , n43904 , n43905 );
and ( n43907 , n381643 , RI15b4ed08_554);
and ( n43908 , n41896 , RI15b4da48_514);
and ( n43909 , n382852 , RI15b4fc08_586);
nor ( n43910 , n43908 , n43909 );
and ( n43911 , n381661 , RI15b4f848_578);
and ( n43912 , n381663 , RI15b4f0c8_562);
nor ( n43913 , n43911 , n43912 );
and ( n43914 , n381667 , RI15b4d2c8_498);
and ( n43915 , n381669 , RI15b4d688_506);
nor ( n43916 , n43914 , n43915 );
and ( n43917 , n381672 , RI15b4de08_522);
and ( n43918 , n381674 , RI15b4f488_570);
nor ( n43919 , n43917 , n43918 );
nand ( n43920 , n43910 , n43913 , n43916 , n43919 );
and ( n43921 , n38323 , n43920 );
and ( n43922 , n381680 , RI15b4c788_474);
nor ( n43923 , n43907 , n43921 , n43922 );
and ( n43924 , n381684 , RI15b4c3c8_466);
and ( n43925 , n381686 , RI15b4e1c8_530);
nor ( n43926 , n43924 , n43925 );
and ( n43927 , n381689 , RI15b4cb48_482);
and ( n43928 , n381691 , RI15b4cf08_490);
nor ( n43929 , n43927 , n43928 );
nand ( n43930 , n43906 , n43923 , n43926 , n43929 );
not ( n43931 , n381695 );
and ( n43932 , n43930 , n43931 );
not ( n43933 , RI15b55c20_791);
not ( n43934 , n379959 );
or ( n43935 , n43933 , n43934 );
or ( n43936 , n379959 , RI15b55c20_791);
nand ( n43937 , n43935 , n43936 );
and ( n43938 , n379949 , n43937 );
nor ( n43939 , n43932 , n43938 );
nand ( n43940 , n43903 , n43939 );
buf ( n43941 , n43940 );
not ( n43942 , n381570 );
not ( n43943 , n380703 );
or ( n43944 , n43942 , n43943 );
and ( n43945 , n380719 , n381599 );
or ( n43946 , n381609 , n19034 );
or ( n43947 , n380782 , n381619 );
or ( n43948 , n381607 , n380790 );
nand ( n43949 , n43946 , n43947 , n43948 );
nor ( n43950 , n43945 , n43949 );
nand ( n43951 , n43944 , n43950 );
buf ( n43952 , n43951 );
buf ( n43953 , n384218 );
buf ( n43954 , n385195 );
buf ( n43955 , n22738 );
buf ( n43956 , n383613 );
buf ( n43957 , n22714 );
buf ( n43958 , n381707 );
buf ( n43959 , n32255 );
nor ( n43960 , RI15b48318_328 , RI15b48408_330);
nor ( n43961 , n382080 , n43960 );
or ( n43962 , n43961 , RI15b47fd0_321);
and ( n43963 , n37001 , RI15b45f00_251);
and ( n43964 , n385218 , n382078 );
nor ( n43965 , n43963 , n43964 );
nand ( n43966 , n43962 , n43965 );
buf ( n43967 , n43966 );
nand ( n43968 , n35677 , RI15b5d330_1045);
or ( n43969 , n31052 , n43968 );
not ( n43970 , RI15b5d498_1048);
or ( n43971 , n40944 , n43970 );
nand ( n43972 , n43969 , n43971 );
buf ( n43973 , n43972 );
buf ( n43974 , n385195 );
not ( n43975 , n31479 );
not ( n43976 , n43975 );
not ( n43977 , n31494 );
nand ( n43978 , n34859 , n43977 );
not ( n43979 , n379338 );
buf ( n43980 , n31483 );
nand ( n43981 , n43979 , n43980 );
nor ( n43982 , n43978 , n43981 );
nand ( n43983 , n43976 , n43982 );
buf ( n43984 , n31522 );
not ( n43985 , n43984 );
nor ( n43986 , n43983 , n43985 );
buf ( n43987 , n31474 );
not ( n43988 , n43987 );
nand ( n43989 , n43986 , n43988 );
not ( n43990 , n31467 );
and ( n43991 , n43989 , n43990 );
not ( n43992 , n43989 );
and ( n43993 , n43992 , n31467 );
nor ( n43994 , n43991 , n43993 );
nand ( n43995 , n43994 , n31601 );
not ( n43996 , n379391 );
not ( n43997 , n40963 );
or ( n43998 , n43996 , n43997 );
nand ( n43999 , n43998 , n31700 );
and ( n44000 , n43999 , n379158 );
or ( n44001 , n40963 , n31709 , n379158 );
and ( n44002 , n379394 , RI15b57c00_859);
and ( n44003 , n31712 , RI15b51a08_650);
nor ( n44004 , n44002 , n44003 );
nand ( n44005 , n44001 , n44004 );
nor ( n44006 , n44000 , n44005 );
nand ( n44007 , n43995 , n44006 );
buf ( n44008 , n44007 );
buf ( n44009 , n19655 );
buf ( n44010 , n20665 );
not ( n44011 , n42930 );
not ( n44012 , n35838 );
or ( n44013 , n44011 , n44012 );
and ( n44014 , n33196 , n35872 );
not ( n44015 , RI15b40d70_77);
or ( n44016 , n35884 , n44015 );
or ( n44017 , n22241 , n35888 );
or ( n44018 , n35882 , n33201 );
nand ( n44019 , n44016 , n44017 , n44018 );
nor ( n44020 , n44014 , n44019 );
nand ( n44021 , n44013 , n44020 );
buf ( n44022 , n44021 );
or ( n44023 , n35852 , n35895 );
and ( n44024 , n35912 , RI15b402a8_54);
or ( n44025 , n35582 , n35917 );
or ( n44026 , n35856 , n35909 );
or ( n44027 , n35900 , n35858 );
nand ( n44028 , n44025 , n44026 , n44027 );
nor ( n44029 , n44024 , n44028 );
nand ( n44030 , n44023 , n44029 );
buf ( n44031 , n44030 );
buf ( n44032 , n384218 );
buf ( n44033 , n383498 );
buf ( n44034 , n30992 );
not ( n44035 , n384807 );
nand ( n44036 , n384907 , n44035 );
not ( n44037 , n384913 );
not ( n44038 , n384802 );
buf ( n44039 , n44038 );
nand ( n44040 , n44037 , n44039 );
nand ( n44041 , n384918 , RI15b5f5e0_1119);
not ( n44042 , n384922 );
or ( n44043 , n44042 , n383566 );
not ( n44044 , n384927 );
nand ( n44045 , n44043 , n44044 );
and ( n44046 , n44045 , n383574 );
and ( n44047 , n384934 , n38982 );
nor ( n44048 , n44046 , n44047 );
nand ( n44049 , n44036 , n44040 , n44041 , n44048 );
buf ( n44050 , n44049 );
buf ( n44051 , n35651 );
buf ( n44052 , n33382 );
buf ( n44053 , n19651 );
or ( n44054 , n31149 , n384704 );
and ( n44055 , n31161 , n384739 );
or ( n44056 , n384749 , n17678 );
or ( n44057 , n31179 , n384757 );
or ( n44058 , n384747 , n31184 );
nand ( n44059 , n44056 , n44057 , n44058 );
nor ( n44060 , n44055 , n44059 );
nand ( n44061 , n44054 , n44060 );
buf ( n44062 , n44061 );
buf ( n44063 , n22714 );
buf ( n44064 , n43091 );
buf ( n44065 , n44064 );
nor ( n44066 , n44065 , n382079 );
or ( n44067 , n44066 , n32958 );
nand ( n44068 , n44067 , n32851 );
nor ( n44069 , n43104 , n32851 );
and ( n44070 , n44065 , n44069 );
not ( n44071 , n382513 );
not ( n44072 , n44071 );
or ( n44073 , n382347 , n382366 );
not ( n44074 , n44073 );
not ( n44075 , n32841 );
and ( n44076 , n44074 , n44075 );
and ( n44077 , n44073 , n32841 );
nor ( n44078 , n44076 , n44077 );
or ( n44079 , n44072 , n44078 );
and ( n44080 , n382523 , RI15b4b978_444);
and ( n44081 , n32974 , RI15b45780_235);
nor ( n44082 , n44080 , n44081 );
nand ( n44083 , n44079 , n44082 );
nor ( n44084 , n44070 , n44083 );
nand ( n44085 , n44068 , n44084 );
buf ( n44086 , n44085 );
buf ( n44087 , n22479 );
buf ( n44088 , n384996 );
buf ( n44089 , n31979 );
buf ( n44090 , n31719 );
buf ( n44091 , n383556 );
buf ( n44092 , n44091 );
and ( n44093 , n383505 , n44092 );
nor ( n44094 , n44093 , n383577 );
or ( n44095 , n44094 , n383565 );
and ( n44096 , n383601 , RI15b5fce8_1134);
not ( n44097 , n383565 );
nor ( n44098 , n44097 , n44091 );
and ( n44099 , n383603 , n44098 );
and ( n44100 , n383607 , RI15b5f568_1118);
nor ( n44101 , n44096 , n44099 , n44100 );
nand ( n44102 , n44095 , n44101 );
buf ( n44103 , n44102 );
buf ( n44104 , n35649 );
buf ( n44105 , n379403 );
or ( n44106 , n31006 , n383845 );
and ( n44107 , n31016 , n383878 );
or ( n44108 , n383903 , n21004 );
not ( n44109 , n33611 );
or ( n44110 , n44109 , n383911 );
or ( n44111 , n383895 , n31024 );
nand ( n44112 , n44108 , n44110 , n44111 );
nor ( n44113 , n44107 , n44112 );
nand ( n44114 , n44106 , n44113 );
buf ( n44115 , n44114 );
buf ( n44116 , n382049 );
buf ( n44117 , n22402 );
and ( n44118 , n36999 , RI15b480c0_323);
and ( n44119 , n37001 , RI15b44f10_217);
nor ( n44120 , n44118 , n44119 );
not ( n44121 , n44120 );
buf ( n44122 , n44121 );
buf ( n44123 , n380906 );
buf ( n44124 , n379403 );
buf ( n44125 , n17499 );
buf ( n44126 , n382071 );
buf ( n44127 , n384203 );
buf ( n44128 , n381566 );
buf ( n44129 , RI15b5dd80_1067);
not ( n44130 , n43172 );
not ( n44131 , n32129 );
or ( n44132 , n44130 , n44131 );
not ( n44133 , n36318 );
and ( n44134 , n44133 , RI15b419a0_103);
or ( n44135 , n32141 , n22135 );
not ( n44136 , n36325 );
and ( n44137 , n44136 , n39157 );
and ( n44138 , n39159 , n36322 );
nor ( n44139 , n44137 , n44138 );
nand ( n44140 , n44135 , n44139 );
nor ( n44141 , n44134 , n44140 );
nand ( n44142 , n44132 , n44141 );
buf ( n44143 , n44142 );
buf ( n44144 , n384218 );
buf ( n44145 , n31719 );
buf ( n44146 , n20663 );
buf ( n44147 , n386762 );
or ( n44148 , n32955 , n32958 );
nand ( n44149 , n44148 , n32938 );
not ( n44150 , n32945 );
not ( n44151 , n32926 );
or ( n44152 , n44150 , n44151 );
nand ( n44153 , n44152 , n32937 );
not ( n44154 , n382505 );
not ( n44155 , n382504 );
not ( n44156 , n44155 );
or ( n44157 , n44154 , n44156 );
or ( n44158 , n44155 , n382505 );
nand ( n44159 , n44157 , n44158 );
and ( n44160 , n32965 , n44159 );
and ( n44161 , n382523 , RI15b4bf18_456);
and ( n44162 , n32975 , RI15b45d20_247);
nor ( n44163 , n44160 , n44161 , n44162 );
nand ( n44164 , n44149 , n44153 , n44163 );
buf ( n44165 , n44164 );
buf ( n44166 , n32892 );
nand ( n44167 , n43093 , n44166 );
not ( n44168 , n32035 );
and ( n44169 , n44167 , n44168 );
not ( n44170 , n44169 );
buf ( n44171 , n32863 );
not ( n44172 , n44171 );
not ( n44173 , n44172 );
or ( n44174 , n44170 , n44173 );
nor ( n44175 , n44167 , n382079 );
or ( n44176 , n44175 , n32024 );
nand ( n44177 , n44176 , n44173 );
buf ( n44178 , n32864 );
not ( n44179 , n44178 );
buf ( n44180 , n382390 );
buf ( n44181 , n32859 );
nand ( n44182 , n44180 , n44181 );
not ( n44183 , n44182 );
or ( n44184 , n44179 , n44183 );
or ( n44185 , n44182 , n44178 );
nand ( n44186 , n44184 , n44185 );
and ( n44187 , n43433 , n44186 );
and ( n44188 , n382523 , RI15b4bb58_448);
and ( n44189 , n42720 , RI15b45960_239);
nor ( n44190 , n44188 , n44189 );
not ( n44191 , n44190 );
nor ( n44192 , n44187 , n44191 );
nand ( n44193 , n44174 , n44177 , n44192 );
buf ( n44194 , n44193 );
buf ( n44195 , n31979 );
buf ( n44196 , n384218 );
buf ( n44197 , n384700 );
buf ( n44198 , n31979 );
buf ( n44199 , n380203 );
buf ( n44200 , n381490 );
or ( n44201 , n31771 , n18546 );
not ( n44202 , n31781 );
or ( n44203 , n19321 , n44202 );
and ( n44204 , n31778 , n19456 );
and ( n44205 , n32386 , n18550 );
nor ( n44206 , n44204 , n44205 , n40279 );
nand ( n44207 , n44201 , n44203 , n44206 );
buf ( n44208 , n44207 );
not ( n44209 , n383317 );
nand ( n44210 , n44209 , n381461 );
buf ( n44211 , n383316 );
not ( n44212 , n44211 );
or ( n44213 , n44210 , n44212 );
not ( n44214 , n36268 );
or ( n44215 , n44209 , n44214 );
nand ( n44216 , n44215 , n381450 );
not ( n44217 , n44211 );
nand ( n44218 , n44216 , n44217 );
and ( n44219 , n381484 , RI15b52980_683);
buf ( n44220 , n381276 );
nor ( n44221 , n381400 , n44220 );
nor ( n44222 , n44219 , n44221 );
nand ( n44223 , n44213 , n44218 , n44222 );
buf ( n44224 , n44223 );
buf ( n44225 , n383345 );
or ( n44226 , n36119 , n32165 );
and ( n44227 , n38869 , RI15b43368_158);
or ( n44228 , n35856 , n32181 );
or ( n44229 , n35582 , n32187 );
or ( n44230 , n32172 , n35858 );
nand ( n44231 , n44228 , n44229 , n44230 );
nor ( n44232 , n44227 , n44231 );
nand ( n44233 , n44226 , n44232 );
buf ( n44234 , n44233 );
buf ( n44235 , n385197 );
buf ( n44236 , n32981 );
buf ( n44237 , n383498 );
not ( n44238 , RI15b53cb8_724);
not ( n44239 , n32244 );
or ( n44240 , n44238 , n44239 );
and ( n44241 , n32247 , RI15b652b0_1317);
and ( n44242 , n32249 , RI15b60120_1143);
nor ( n44243 , n44241 , n44242 );
nand ( n44244 , n44240 , n44243 );
buf ( n44245 , n44244 );
buf ( n44246 , n35651 );
buf ( n44247 , n32676 );
buf ( n44248 , n22404 );
buf ( n44249 , n382052 );
or ( n44250 , n381056 , n37121 );
and ( n44251 , n35373 , RI15b43458_160);
and ( n44252 , n35376 , RI15b43818_168);
and ( n44253 , n35537 , RI15b43098_152);
and ( n44254 , n35384 , RI15b42cd8_144);
nor ( n44255 , n44253 , n44254 );
and ( n44256 , n35391 , RI15b42198_120);
and ( n44257 , n35546 , RI15b41a18_104);
nor ( n44258 , n44256 , n44257 );
and ( n44259 , n35541 , RI15b41298_88);
and ( n44260 , n35543 , RI15b40ed8_80);
nor ( n44261 , n44259 , n44260 );
and ( n44262 , n35548 , RI15b41658_96);
and ( n44263 , n35396 , RI15b42558_128);
and ( n44264 , n35401 , RI15b3ffd8_48);
and ( n44265 , n35407 , RI15b40398_56);
nor ( n44266 , n44263 , n44264 , n44265 );
and ( n44267 , n35410 , RI15b40b18_72);
and ( n44268 , n35412 , RI15b41dd8_112);
nor ( n44269 , n44267 , n44268 );
and ( n44270 , n35415 , RI15b42918_136);
and ( n44271 , n383378 , RI15b40758_64);
nor ( n44272 , n44270 , n44271 );
and ( n44273 , n44266 , n44269 , n44272 );
nor ( n44274 , n44273 , n381047 );
nor ( n44275 , n44262 , n44274 );
and ( n44276 , n44258 , n44261 , n44275 );
nand ( n44277 , n44255 , n44276 );
nor ( n44278 , n44251 , n44252 , n44277 );
or ( n44279 , n32805 , n44278 );
and ( n44280 , n37120 , RI15b49bf0_381);
not ( n44281 , n37120 );
and ( n44282 , n44281 , n37121 );
nor ( n44283 , n44280 , n44282 );
or ( n44284 , n37109 , n44283 );
nand ( n44285 , n44250 , n44279 , n44284 );
buf ( n44286 , n44285 );
not ( n44287 , n384798 );
nand ( n44288 , n384907 , n44287 );
buf ( n44289 , n384793 );
not ( n44290 , n44289 );
nand ( n44291 , n384914 , n44290 );
nand ( n44292 , n384918 , RI15b5f4f0_1117);
or ( n44293 , n44042 , n383547 );
nand ( n44294 , n44293 , n44044 );
and ( n44295 , n44294 , n383555 );
not ( n44296 , n383555 );
and ( n44297 , n383547 , n44296 );
and ( n44298 , n384934 , n44297 );
nor ( n44299 , n44295 , n44298 );
nand ( n44300 , n44288 , n44291 , n44292 , n44299 );
buf ( n44301 , n44300 );
buf ( n44302 , n384996 );
or ( n44303 , n386705 , n384704 );
and ( n44304 , n386716 , n384739 );
or ( n44305 , n384749 , n17867 );
not ( n44306 , n386731 );
or ( n44307 , n44306 , n384757 );
or ( n44308 , n384747 , n386738 );
nand ( n44309 , n44305 , n44307 , n44308 );
nor ( n44310 , n44304 , n44309 );
nand ( n44311 , n44303 , n44310 );
buf ( n44312 , n44311 );
buf ( n44313 , n381707 );
buf ( n44314 , n31979 );
buf ( n44315 , n21800 );
buf ( n44316 , n40997 );
not ( n44317 , n44316 );
or ( n44318 , n44317 , n41015 );
nand ( n44319 , n44318 , n41032 );
not ( n44320 , n35077 );
nand ( n44321 , n44319 , n44320 );
nor ( n44322 , n44316 , n44320 );
nand ( n44323 , n41578 , n44322 );
nand ( n44324 , n41582 , RI15b46248_258);
nand ( n44325 , n44321 , n44323 , n44324 , n41561 );
buf ( n44326 , n44325 );
buf ( n44327 , n20665 );
buf ( n44328 , n18226 );
buf ( n44329 , n21847 );
not ( n44330 , n21853 );
nor ( n44331 , n44329 , n44330 );
and ( n44332 , n21802 , n44331 );
or ( n44333 , n18074 , n21960 );
nand ( n44334 , n44333 , n21979 );
and ( n44335 , n44334 , RI15b55c20_791);
and ( n44336 , n18150 , RI15b57a20_855);
not ( n44337 , n21960 );
or ( n44338 , n21982 , n44337 , RI15b55c20_791);
and ( n44339 , n21931 , n379136 );
not ( n44340 , n21931 );
and ( n44341 , n44340 , RI15b57a20_855);
nor ( n44342 , n44339 , n44341 );
or ( n44343 , n21922 , n44342 );
nand ( n44344 , n44338 , n44343 );
nor ( n44345 , n44335 , n44336 , n44344 );
or ( n44346 , n44345 , n18078 );
and ( n44347 , n18177 , RI15b57a20_855);
and ( n44348 , n18219 , RI15b56b20_823);
nor ( n44349 , n44347 , n44348 , n21751 );
nand ( n44350 , n44346 , n44349 );
nor ( n44351 , n44332 , n44350 );
nand ( n44352 , n44329 , n17507 );
not ( n44353 , n44352 );
not ( n44354 , n17565 );
or ( n44355 , n44353 , n44354 );
nand ( n44356 , n44355 , n44330 );
nand ( n44357 , n44351 , n44356 );
buf ( n44358 , n44357 );
buf ( n44359 , n382071 );
buf ( n44360 , n382071 );
not ( n44361 , n37989 );
not ( n44362 , n17523 );
or ( n44363 , n44361 , n44362 );
nand ( n44364 , n44363 , n21790 );
and ( n44365 , n44364 , RI15b57480_843);
and ( n44366 , n22564 , n21771 );
nor ( n44367 , n17523 , RI15b57480_843);
and ( n44368 , n21795 , n44367 );
nor ( n44369 , n44365 , n44366 , n44368 );
nand ( n44370 , n36691 , n44369 );
buf ( n44371 , n44370 );
buf ( n44372 , n380865 );
buf ( n44373 , n17499 );
buf ( n44374 , n380203 );
not ( n44375 , n34295 );
not ( n44376 , n44375 );
nor ( n44377 , n34286 , n34288 );
not ( n44378 , n33941 );
and ( n44379 , n44377 , n44378 );
buf ( n44380 , n33960 );
nand ( n44381 , n44379 , n44380 );
buf ( n44382 , n34151 );
not ( n44383 , n44382 );
nor ( n44384 , n44381 , n44383 );
nand ( n44385 , n44384 , n379785 );
not ( n44386 , n44385 );
or ( n44387 , n44376 , n44386 );
and ( n44388 , n33927 , n34193 );
not ( n44389 , n44388 );
nand ( n44390 , n44387 , n44389 );
not ( n44391 , n44384 );
nand ( n44392 , n34249 , n44391 , n44388 );
and ( n44393 , n34651 , RI15b5e6e0_1087);
nor ( n44394 , n44393 , n34644 );
nand ( n44395 , n44390 , n44392 , n44394 );
buf ( n44396 , n44395 );
buf ( n44397 , n384996 );
nor ( n44398 , n40547 , n21652 );
not ( n44399 , n44398 );
not ( n44400 , n42522 );
nand ( n44401 , n44399 , n44400 );
nand ( n44402 , n44401 , n33644 );
and ( n44403 , n21304 , n21311 );
not ( n44404 , n21304 );
and ( n44405 , n44404 , n381764 );
nor ( n44406 , n44403 , n44405 );
and ( n44407 , n44406 , n21360 );
not ( n44408 , RI15b57e58_864);
not ( n44409 , n21751 );
or ( n44410 , n44408 , n44409 );
buf ( n44411 , n21523 );
not ( n44412 , n44411 );
not ( n44413 , n21527 );
and ( n44414 , n44412 , n44413 );
and ( n44415 , n44411 , n21527 );
nor ( n44416 , n44414 , n44415 );
or ( n44417 , n44416 , n42540 );
nand ( n44418 , n44410 , n44417 );
nor ( n44419 , n44407 , n44418 );
nand ( n44420 , n44402 , n44419 );
not ( n44421 , n44420 );
and ( n44422 , n385164 , RI15b507c0_611);
not ( n44423 , n385174 );
or ( n44424 , n44423 , n21652 );
or ( n44425 , n21311 , n385170 );
or ( n44426 , n21527 , n385178 );
nand ( n44427 , n44424 , n44425 , n44426 );
nor ( n44428 , n44422 , n44427 );
nand ( n44429 , n44421 , n44428 );
buf ( n44430 , n44429 );
buf ( n44431 , n381014 );
or ( n44432 , n44431 , n380965 );
nand ( n44433 , n35525 , RI15b540f0_733);
nand ( n44434 , n44432 , n44433 );
buf ( n44435 , n44434 );
and ( n44436 , n39423 , n41715 );
and ( n44437 , n35335 , RI15b65c88_1338);
not ( n44438 , RI15b488b8_340);
not ( n44439 , n35346 );
or ( n44440 , n44438 , n44439 );
or ( n44441 , n35346 , RI15b488b8_340);
nand ( n44442 , n44440 , n44441 );
and ( n44443 , n35363 , n44442 );
nor ( n44444 , n44436 , n44437 , n44443 );
nand ( n44445 , n41726 , RI15b488b8_340);
nand ( n44446 , n32493 , n44444 , n44445 );
buf ( n44447 , n44446 );
buf ( n44448 , n380940 );
buf ( n44449 , n380906 );
buf ( n44450 , n19653 );
buf ( n44451 , n386762 );
not ( n44452 , RI15b61980_1195);
nand ( n44453 , n31128 , n33503 );
and ( n44454 , n43059 , n44453 );
not ( n44455 , n44454 );
not ( n44456 , n44455 );
or ( n44457 , n44452 , n44456 );
and ( n44458 , n43062 , n33510 );
buf ( n44459 , n41431 );
not ( n44460 , n38723 );
not ( n44461 , n38750 );
and ( n44462 , n44460 , n44461 );
and ( n44463 , n38723 , n38750 );
nor ( n44464 , n44462 , n44463 );
or ( n44465 , n44459 , n44464 );
or ( n44466 , n31052 , n380597 );
nand ( n44467 , n44465 , n44466 );
nor ( n44468 , n42641 , n44289 );
nor ( n44469 , n44458 , n44467 , n44468 );
nand ( n44470 , n44457 , n44469 );
buf ( n44471 , n44470 );
buf ( n44472 , n19653 );
not ( n44473 , n36259 );
not ( n44474 , n384122 );
or ( n44475 , n44473 , n44474 );
and ( n44476 , n384164 , n43075 );
or ( n44477 , n36250 , n20870 );
or ( n44478 , n384187 , n36254 );
or ( n44479 , n36248 , n384193 );
nand ( n44480 , n44477 , n44478 , n44479 );
nor ( n44481 , n44476 , n44480 );
nand ( n44482 , n44475 , n44481 );
buf ( n44483 , n44482 );
buf ( n44484 , n380203 );
buf ( n44485 , RI15b47490_297);
buf ( n44486 , n17499 );
nand ( n44487 , n379816 , n382040 );
and ( n44488 , n382033 , n44487 , n379812 );
nor ( n44489 , n382032 , n382040 );
or ( n44490 , n44489 , n379812 , n22254 );
nand ( n44491 , n44490 , n379820 );
nor ( n44492 , n44488 , n44491 );
not ( n44493 , n44492 );
nand ( n44494 , n35187 , RI15b48b88_346);
not ( n44495 , n35456 );
nand ( n44496 , n36049 , n44495 );
and ( n44497 , n35335 , RI15b65f58_1344);
not ( n44498 , RI15b48b88_346);
not ( n44499 , n35353 );
not ( n44500 , n44499 );
or ( n44501 , n44498 , n44500 );
or ( n44502 , n44499 , RI15b48b88_346);
nand ( n44503 , n44501 , n44502 );
buf ( n44504 , n35363 );
and ( n44505 , n44503 , n44504 );
nor ( n44506 , n44497 , n44505 );
nand ( n44507 , n44493 , n44494 , n44496 , n44506 );
buf ( n44508 , n44507 );
buf ( n44509 , n386760 );
or ( n44510 , n381015 , n22059 );
nand ( n44511 , n381017 , RI15b53e20_727);
nand ( n44512 , n44510 , n44511 );
buf ( n44513 , n44512 );
buf ( n44514 , n19653 );
buf ( n44515 , n380906 );
buf ( n44516 , n32676 );
buf ( n44517 , n380903 );
buf ( n44518 , n384199 );
buf ( n44519 , n379802 );
or ( n44520 , n35852 , n37495 );
not ( n44521 , n37507 );
and ( n44522 , n44521 , RI15b42468_126);
or ( n44523 , n35856 , n37505 );
or ( n44524 , n35582 , n37512 );
or ( n44525 , n37497 , n35858 );
nand ( n44526 , n44523 , n44524 , n44525 );
nor ( n44527 , n44522 , n44526 );
nand ( n44528 , n44520 , n44527 );
buf ( n44529 , n44528 );
buf ( n44530 , n33382 );
not ( n44531 , n19857 );
not ( n44532 , n20637 );
or ( n44533 , n44531 , n44532 );
nand ( n44534 , n44533 , n34798 );
and ( n44535 , n44534 , RI15b4ac58_416);
or ( n44536 , n34801 , n19857 , RI15b4ac58_416);
or ( n44537 , n19860 , n22216 );
nand ( n44538 , n44536 , n44537 );
nor ( n44539 , n44535 , n44538 );
nand ( n44540 , n40388 , n44539 );
buf ( n44541 , n44540 );
buf ( n44542 , n32981 );
buf ( n44543 , n32255 );
not ( n44544 , n387035 );
not ( n44545 , n44544 );
not ( n44546 , n22449 );
or ( n44547 , n44545 , n44546 );
nand ( n44548 , n44547 , n34811 );
and ( n44549 , n44548 , RI15b64248_1282);
not ( n44550 , n34814 );
buf ( n44551 , n386979 );
not ( n44552 , n44551 );
or ( n44553 , n44550 , n44552 );
nand ( n44554 , n44553 , n34823 );
and ( n44555 , n44554 , RI15b62448_1218);
or ( n44556 , n34826 , n44551 , RI15b62448_1218);
and ( n44557 , n379632 , RI15b64248_1282);
nor ( n44558 , n44544 , n379632 , RI15b64248_1282);
nor ( n44559 , n44557 , n44558 );
or ( n44560 , n34833 , n44559 );
nand ( n44561 , n44556 , n44560 );
nor ( n44562 , n44549 , n44555 , n44561 );
or ( n44563 , n44562 , n19200 );
not ( n44564 , n386871 );
not ( n44565 , n44564 );
not ( n44566 , n22473 );
and ( n44567 , n44565 , n44566 );
not ( n44568 , n383474 );
nor ( n44569 , n44567 , n44568 );
or ( n44570 , n386878 , n44569 );
and ( n44571 , n38117 , n44564 , n386878 );
or ( n44572 , n22424 , n379662 );
or ( n44573 , n386876 , n19598 );
nand ( n44574 , n44572 , n44573 , n19512 );
nor ( n44575 , n44571 , n44574 );
nand ( n44576 , n44563 , n44570 , n44575 );
buf ( n44577 , n44576 );
buf ( n44578 , RI15b5e488_1082);
buf ( n44579 , n384700 );
buf ( n44580 , n22714 );
buf ( n44581 , n22716 );
not ( n44582 , n20545 );
and ( n44583 , n20565 , n44582 );
nor ( n44584 , n44583 , n22372 );
not ( n44585 , n44584 );
and ( n44586 , n44585 , RI15b4b888_442);
buf ( n44587 , n19976 );
not ( n44588 , n44587 );
not ( n44589 , n22377 );
or ( n44590 , n44588 , n44589 );
nand ( n44591 , n44590 , n383364 );
and ( n44592 , n44591 , RI15b49a88_378);
or ( n44593 , n22359 , n44587 , RI15b49a88_378);
and ( n44594 , n20547 , RI15b4b888_442);
nor ( n44595 , n44582 , n20547 , RI15b4b888_442);
nor ( n44596 , n44594 , n44595 );
or ( n44597 , n20564 , n44596 );
nand ( n44598 , n44593 , n44597 );
nor ( n44599 , n44586 , n44592 , n44598 );
or ( n44600 , n44599 , n20519 );
buf ( n44601 , n19822 );
not ( n44602 , n19815 );
not ( n44603 , n44602 );
not ( n44604 , n19918 );
and ( n44605 , n44603 , n44604 );
nor ( n44606 , n44605 , n384684 );
or ( n44607 , n44601 , n44606 );
and ( n44608 , n384687 , n44602 , n44601 );
or ( n44609 , n20639 , n20546 );
or ( n44610 , n19820 , n22390 );
nand ( n44611 , n44609 , n44610 , n384692 );
nor ( n44612 , n44608 , n44611 );
nand ( n44613 , n44600 , n44607 , n44612 );
buf ( n44614 , n44613 );
and ( n44615 , n19646 , n383419 );
nor ( n44616 , n384641 , n44615 );
or ( n44617 , n44616 , n383420 );
or ( n44618 , n31971 , n383419 , RI15b63618_1256);
nand ( n44619 , n386912 , n19630 );
nand ( n44620 , n44618 , n44619 );
nor ( n44621 , n40706 , n44620 );
nand ( n44622 , n44617 , n44621 );
buf ( n44623 , n44622 );
buf ( n44624 , n22738 );
buf ( n44625 , n31719 );
buf ( n44626 , n19651 );
or ( n44627 , n22315 , n36121 );
and ( n44628 , n22326 , n36123 );
or ( n44629 , n36132 , n20175 );
or ( n44630 , n22334 , n36139 );
or ( n44631 , n36130 , n22336 );
nand ( n44632 , n44629 , n44630 , n44631 );
nor ( n44633 , n44628 , n44632 );
nand ( n44634 , n44627 , n44633 );
buf ( n44635 , n44634 );
buf ( n44636 , n33382 );
buf ( n44637 , n379895 );
buf ( n44638 , n22653 );
buf ( n44639 , n22655 );
buf ( n44640 , n381566 );
or ( n44641 , n18167 , n18072 );
nand ( n44642 , n44641 , n18151 , n21786 );
nand ( n44643 , n44642 , RI15b54258_736);
or ( n44644 , n18097 , n17505 );
not ( n44645 , n36342 );
nand ( n44646 , n44644 , n44645 );
and ( n44647 , n40884 , n33211 , n35244 );
nor ( n44648 , n44647 , n383166 );
nand ( n44649 , n18204 , n383913 , n382546 );
nand ( n44650 , n44643 , n44646 , n44648 , n44649 );
buf ( n44651 , n44650 );
not ( n44652 , n33220 );
not ( n44653 , n381507 );
or ( n44654 , n44652 , n44653 );
and ( n44655 , n381524 , n33226 );
or ( n44656 , n33237 , n18400 );
or ( n44657 , n36413 , n33241 );
or ( n44658 , n33235 , n381560 );
nand ( n44659 , n44656 , n44657 , n44658 );
nor ( n44660 , n44655 , n44659 );
nand ( n44661 , n44654 , n44660 );
buf ( n44662 , n44661 );
buf ( n44663 , n381006 );
buf ( n44664 , n22007 );
buf ( n44665 , n32981 );
buf ( n44666 , n22716 );
buf ( n44667 , n381004 );
buf ( n44668 , n22007 );
not ( n44669 , n41267 );
or ( n44670 , n44669 , n386419 );
not ( n44671 , n385822 );
not ( n44672 , n39947 );
or ( n44673 , n44671 , n44672 );
or ( n44674 , n39947 , n385822 );
nand ( n44675 , n44673 , n44674 );
and ( n44676 , n44675 , n386019 );
not ( n44677 , n39961 );
not ( n44678 , n386162 );
and ( n44679 , n44677 , n44678 );
and ( n44680 , n39961 , n386162 );
nor ( n44681 , n44679 , n44680 );
or ( n44682 , n44681 , n386261 );
buf ( n44683 , n34727 );
and ( n44684 , n44683 , n34728 );
buf ( n44685 , n34729 );
nor ( n44686 , n44684 , n44685 );
or ( n44687 , n44686 , n386499 );
not ( n44688 , RI15b4b630_437);
or ( n44689 , n40759 , n44688 );
nand ( n44690 , n44682 , n44687 , n44689 );
nor ( n44691 , n44676 , n44690 );
and ( n44692 , n386540 , RI15b43f98_184);
and ( n44693 , n386549 , n385822 );
and ( n44694 , n386556 , n39962 );
nor ( n44695 , n44692 , n44693 , n44694 );
nand ( n44696 , n44670 , n44691 , n44695 );
buf ( n44697 , n44696 );
buf ( n44698 , n22343 );
buf ( n44699 , n382065 );
not ( n44700 , n22552 );
nor ( n44701 , n44700 , n17506 );
or ( n44702 , n44701 , n379905 );
not ( n44703 , n22558 );
nand ( n44704 , n44702 , n44703 );
not ( n44705 , n22594 );
nor ( n44706 , n44705 , n18079 );
or ( n44707 , n44706 , n18103 );
nand ( n44708 , n44707 , RI15b56508_810);
nor ( n44709 , n18197 , RI15b56508_810);
and ( n44710 , n44705 , n44709 );
not ( n44711 , n18188 );
not ( n44712 , n22621 );
or ( n44713 , n44711 , n44712 );
nand ( n44714 , n44713 , n22604 );
and ( n44715 , n44714 , RI15b58308_874);
or ( n44716 , n18189 , n22621 , RI15b58308_874);
or ( n44717 , n18218 , n22556 );
nand ( n44718 , n44716 , n44717 );
nor ( n44719 , n44715 , n44718 );
not ( n44720 , n44719 );
nor ( n44721 , n44710 , n44720 );
nor ( n44722 , n17576 , n44703 );
nand ( n44723 , n44700 , n44722 );
nand ( n44724 , n44704 , n44708 , n44721 , n44723 );
buf ( n44725 , n44724 );
buf ( n44726 , n386563 );
buf ( n44727 , n380203 );
buf ( n44728 , n385115 );
or ( n44729 , n44728 , n385116 );
buf ( n44730 , n385117 );
not ( n44731 , n44730 );
nand ( n44732 , n44729 , n44731 );
and ( n44733 , n44732 , n385133 );
buf ( n44734 , n21257 );
not ( n44735 , n21282 );
and ( n44736 , n44734 , n44735 );
not ( n44737 , n44734 );
and ( n44738 , n44737 , n21282 );
nor ( n44739 , n44736 , n44738 );
not ( n44740 , n21354 );
or ( n44741 , n44739 , n44740 );
not ( n44742 , n21494 );
not ( n44743 , n44742 );
buf ( n44744 , n21479 );
not ( n44745 , n44744 );
or ( n44746 , n44743 , n44745 );
or ( n44747 , n44744 , n44742 );
nand ( n44748 , n44746 , n44747 );
not ( n44749 , n21560 );
and ( n44750 , n44748 , n44749 );
and ( n44751 , n21751 , RI15b57a98_856);
nor ( n44752 , n44750 , n44751 );
nand ( n44753 , n44741 , n44752 );
nor ( n44754 , n44733 , n44753 );
and ( n44755 , n21788 , RI15b56b98_824);
not ( n44756 , n21861 );
and ( n44757 , n44756 , n21768 );
not ( n44758 , n21855 );
and ( n44759 , n44758 , n21859 );
not ( n44760 , n44758 );
and ( n44761 , n44760 , RI15b56b98_824);
nor ( n44762 , n44759 , n44761 );
and ( n44763 , n44762 , n22704 );
nor ( n44764 , n44755 , n44757 , n44763 );
nand ( n44765 , n44754 , n44764 );
buf ( n44766 , n44765 );
buf ( n44767 , n381872 );
buf ( n44768 , n383345 );
nand ( n44769 , n43144 , n35063 );
buf ( n44770 , n44769 );
nor ( n44771 , n44770 , n41015 );
or ( n44772 , n44771 , n41033 );
buf ( n44773 , n35025 );
buf ( n44774 , n44773 );
buf ( n44775 , n44774 );
nand ( n44776 , n44772 , n44775 );
nor ( n44777 , n41036 , n44774 );
and ( n44778 , n44770 , n44777 );
not ( n44779 , RI15b46590_265);
not ( n44780 , n41017 );
or ( n44781 , n44779 , n44780 );
not ( n44782 , n382016 );
not ( n44783 , n44782 );
not ( n44784 , n382003 );
or ( n44785 , n44783 , n44784 );
or ( n44786 , n382003 , n44782 );
nand ( n44787 , n44785 , n44786 );
and ( n44788 , n35461 , n44787 );
not ( n44789 , n382012 );
and ( n44790 , n35459 , n44789 );
nor ( n44791 , n44788 , n44790 );
nand ( n44792 , n44781 , n44791 );
nor ( n44793 , n44778 , n44792 );
nand ( n44794 , n44776 , n44793 );
buf ( n44795 , n44794 );
buf ( n44796 , n32672 );
buf ( n44797 , n22402 );
not ( n44798 , n41991 );
nand ( n44799 , n44798 , n18098 );
and ( n44800 , n40882 , n44799 );
not ( n44801 , n40830 );
and ( n44802 , n44801 , n18077 );
nor ( n44803 , n44802 , n383147 );
nand ( n44804 , n40883 , n44803 );
and ( n44805 , n44804 , RI15b51210_633);
or ( n44806 , n18169 , n35244 );
not ( n44807 , n37989 );
nand ( n44808 , n44806 , n44807 , n18171 );
nor ( n44809 , n44805 , n44808 );
nand ( n44810 , n44800 , n44809 );
buf ( n44811 , n44810 );
buf ( n44812 , n32271 );
buf ( n44813 , n386760 );
not ( n44814 , n39188 );
not ( n44815 , n44814 );
buf ( n44816 , n34323 );
not ( n44817 , n44816 );
nand ( n44818 , n44815 , n44817 );
and ( n44819 , n44818 , n34336 );
not ( n44820 , n44818 );
not ( n44821 , n34336 );
and ( n44822 , n44820 , n44821 );
nor ( n44823 , n44819 , n44822 );
nand ( n44824 , n44823 , n34643 );
not ( n44825 , n36556 );
not ( n44826 , n44825 );
not ( n44827 , n36557 );
or ( n44828 , n44826 , n44827 );
or ( n44829 , n36557 , n44825 );
nand ( n44830 , n44828 , n44829 );
nand ( n44831 , n44830 , n379785 );
and ( n44832 , n379783 , RI15b63e88_1274);
and ( n44833 , n34650 , RI15b5dc90_1065);
nor ( n44834 , n44832 , n44833 );
nand ( n44835 , n44824 , n44831 , n44834 );
buf ( n44836 , n44835 );
buf ( n44837 , n22740 );
not ( n44838 , RI15b539e8_718);
not ( n44839 , n32244 );
or ( n44840 , n44838 , n44839 );
and ( n44841 , n32247 , RI15b64fe0_1311);
and ( n44842 , n32249 , RI15b5fe50_1137);
nor ( n44843 , n44841 , n44842 );
nand ( n44844 , n44840 , n44843 );
buf ( n44845 , n44844 );
buf ( n44846 , n32255 );
buf ( n44847 , n32255 );
and ( n44848 , n37127 , n37128 );
not ( n44849 , n37127 );
and ( n44850 , n44849 , RI15b49ec0_387);
nor ( n44851 , n44848 , n44850 );
nand ( n44852 , n44851 , n37112 );
and ( n44853 , n381055 , RI15b49ec0_387);
and ( n44854 , n37201 , n37229 );
buf ( n44855 , n36023 );
not ( n44856 , n44855 );
not ( n44857 , n37230 );
nor ( n44858 , n44854 , n44856 , n44857 );
not ( n44859 , n42688 );
and ( n44860 , n44858 , n44859 );
nor ( n44861 , n44853 , n44860 );
nand ( n44862 , n44852 , n44861 );
buf ( n44863 , n44862 );
buf ( n44864 , n32981 );
buf ( n44865 , n379893 );
buf ( n44866 , n386762 );
not ( n44867 , RI15b52c50_689);
not ( n44868 , n381485 );
or ( n44869 , n44867 , n44868 );
or ( n44870 , n381423 , RI15b548e8_750);
nand ( n44871 , n44870 , n381450 , n381460 );
and ( n44872 , n44871 , RI15b54960_751);
nand ( n44873 , n381401 , n383905 );
not ( n44874 , n44873 );
nor ( n44875 , n44872 , n44874 );
nand ( n44876 , n44869 , n44875 );
buf ( n44877 , n44876 );
not ( n44878 , n36276 );
not ( n44879 , n381589 );
or ( n44880 , n44878 , n44879 );
and ( n44881 , n381596 , n36282 );
or ( n44882 , n36291 , n18691 );
or ( n44883 , n32420 , n36296 );
or ( n44884 , n36289 , n381621 );
nand ( n44885 , n44882 , n44883 , n44884 );
nor ( n44886 , n44881 , n44885 );
nand ( n44887 , n44880 , n44886 );
buf ( n44888 , n44887 );
buf ( n44889 , n381490 );
buf ( n44890 , n382537 );
buf ( n44891 , n19651 );
buf ( n44892 , n22408 );
not ( n44893 , n41652 );
and ( n44894 , n44893 , n34931 );
nor ( n44895 , n44894 , n35114 );
or ( n44896 , n44895 , n41653 );
and ( n44897 , n41652 , n35118 , n41653 );
and ( n44898 , n20631 , RI15b464a0_263);
nor ( n44899 , n44897 , n44898 );
nand ( n44900 , n385213 , RI15b47aa8_310);
nand ( n44901 , n44896 , n44899 , n44900 );
buf ( n44902 , n44901 );
buf ( n44903 , n31033 );
buf ( n44904 , n22655 );
buf ( n44905 , n382537 );
buf ( n44906 , n34742 );
buf ( n44907 , n34743 );
nor ( n44908 , n44906 , n44907 );
not ( n44909 , n44908 );
nand ( n44910 , n44909 , n34744 );
nand ( n44911 , n44910 , n386500 );
buf ( n44912 , n34757 );
and ( n44913 , n44912 , n386186 );
not ( n44914 , n44912 );
not ( n44915 , n386186 );
and ( n44916 , n44914 , n44915 );
nor ( n44917 , n44913 , n44916 );
and ( n44918 , n44917 , n34767 );
buf ( n44919 , n34771 );
not ( n44920 , n44919 );
not ( n44921 , n385902 );
and ( n44922 , n44920 , n44921 );
and ( n44923 , n44919 , n385902 );
nor ( n44924 , n44922 , n44923 );
or ( n44925 , n44924 , n38149 );
not ( n44926 , n39987 );
or ( n44927 , n44926 , n382117 );
nand ( n44928 , n44925 , n44927 );
nor ( n44929 , n44918 , n44928 );
nand ( n44930 , n44911 , n44929 );
not ( n44931 , n44930 );
not ( n44932 , n41307 );
not ( n44933 , n44907 );
and ( n44934 , n44932 , n44933 );
or ( n44935 , n386541 , n385893 );
or ( n44936 , n385902 , n386550 );
or ( n44937 , n386186 , n386557 );
nand ( n44938 , n44935 , n44936 , n44937 );
nor ( n44939 , n44934 , n44938 );
nand ( n44940 , n44931 , n44939 );
buf ( n44941 , n44940 );
buf ( n44942 , n379893 );
buf ( n44943 , n36854 );
or ( n44944 , n386588 , n382975 );
and ( n44945 , n386600 , n382983 );
not ( n44946 , RI15b5adb0_965);
or ( n44947 , n382995 , n44946 );
or ( n44948 , n34706 , n383001 );
or ( n44949 , n382993 , n386627 );
nand ( n44950 , n44947 , n44948 , n44949 );
nor ( n44951 , n44945 , n44950 );
nand ( n44952 , n44944 , n44951 );
buf ( n44953 , n44952 );
not ( n44954 , n383153 );
not ( n44955 , n383320 );
or ( n44956 , n44954 , n44955 );
nand ( n44957 , n44956 , n383157 );
nand ( n44958 , n44957 , n41997 );
nor ( n44959 , n41997 , n383144 );
and ( n44960 , n41999 , n44959 );
not ( n44961 , RI15b52ae8_686);
not ( n44962 , n383147 );
or ( n44963 , n44961 , n44962 );
nand ( n44964 , n383170 , RI15b540f0_733);
nand ( n44965 , n44963 , n44964 );
nor ( n44966 , n44960 , n44965 );
nand ( n44967 , n44958 , n44966 );
buf ( n44968 , n44967 );
buf ( n44969 , n379847 );
buf ( n44970 , n380903 );
buf ( n44971 , n36854 );
buf ( n44972 , n32672 );
buf ( n44973 , n32271 );
nor ( n44974 , n43145 , n34930 );
or ( n44975 , n44974 , n35114 );
nand ( n44976 , n44975 , n43148 );
nor ( n44977 , n35117 , n43148 );
and ( n44978 , n43145 , n44977 );
and ( n44979 , n20631 , RI15b46518_264);
nor ( n44980 , n44978 , n44979 );
nand ( n44981 , n385213 , RI15b47b20_311);
nand ( n44982 , n44976 , n44980 , n44981 );
buf ( n44983 , n44982 );
buf ( n44984 , n382052 );
not ( n44985 , n38480 );
and ( n44986 , n44985 , n384025 );
nor ( n44987 , n44986 , n384022 );
or ( n44988 , n44987 , n386983 );
and ( n44989 , n38480 , n384025 , n386983 );
and ( n44990 , n38654 , RI15b5b260_975);
and ( n44991 , n42603 , RI15b5aea0_967);
nor ( n44992 , n44990 , n44991 );
and ( n44993 , n42606 , RI15b5aae0_959);
and ( n44994 , n42608 , RI15b5a720_951);
nor ( n44995 , n44993 , n44994 );
and ( n44996 , n42611 , RI15b5a360_943);
and ( n44997 , n42613 , RI15b59fa0_935);
nor ( n44998 , n44996 , n44997 );
and ( n44999 , n42616 , RI15b59be0_927);
and ( n45000 , n42618 , RI15b59820_919);
nor ( n45001 , n44999 , n45000 );
nand ( n45002 , n44992 , n44995 , n44998 , n45001 );
and ( n45003 , n41935 , n45002 );
and ( n45004 , n39746 , RI15b58ce0_895);
and ( n45005 , n39751 , RI15b5c160_1007);
nor ( n45006 , n45003 , n45004 , n45005 );
and ( n45007 , n39756 , RI15b5bda0_999);
and ( n45008 , n39759 , RI15b5b9e0_991);
nor ( n45009 , n45007 , n45008 );
and ( n45010 , n39763 , RI15b59460_911);
and ( n45011 , n39765 , RI15b590a0_903);
nor ( n45012 , n45010 , n45011 );
and ( n45013 , n39769 , RI15b58920_887);
and ( n45014 , n39772 , RI15b5b620_983);
nor ( n45015 , n45013 , n45014 );
nand ( n45016 , n45006 , n45009 , n45012 , n45015 );
and ( n45017 , n45016 , n39776 );
nor ( n45018 , n44989 , n45017 );
nand ( n45019 , n44988 , n45018 );
buf ( n45020 , n45019 );
buf ( n45021 , n22740 );
buf ( n45022 , n22738 );
buf ( n45023 , n385112 );
buf ( n45024 , n382071 );
or ( n45025 , n36937 , n39691 );
and ( n45026 , n36946 , n39694 );
or ( n45027 , n39703 , n17803 );
or ( n45028 , n38403 , n39707 );
or ( n45029 , n39701 , n36955 );
nand ( n45030 , n45027 , n45028 , n45029 );
nor ( n45031 , n45026 , n45030 );
nand ( n45032 , n45025 , n45031 );
buf ( n45033 , n45032 );
or ( n45034 , n381907 , n38373 );
not ( n45035 , n38385 );
and ( n45036 , n45035 , RI15b43098_152);
or ( n45037 , n381917 , n38377 );
not ( n45038 , n38389 );
and ( n45039 , n45038 , n381923 );
and ( n45040 , n381926 , n38387 );
nor ( n45041 , n45039 , n45040 );
nand ( n45042 , n45037 , n45041 );
nor ( n45043 , n45036 , n45042 );
nand ( n45044 , n45034 , n45043 );
buf ( n45045 , n45044 );
buf ( n45046 , n380940 );
buf ( n45047 , n20663 );
buf ( n45048 , n382071 );
buf ( n45049 , n385197 );
buf ( n45050 , n32160 );
buf ( n45051 , n386760 );
not ( n45052 , n31806 );
not ( n45053 , n19991 );
not ( n45054 , n45053 );
or ( n45055 , n45052 , n45054 );
nand ( n45056 , n45055 , n380875 );
and ( n45057 , n45056 , RI15b49ec0_387);
or ( n45058 , n45053 , n20529 , RI15b49ec0_387);
and ( n45059 , n20647 , n20556 , n41261 );
and ( n45060 , n20656 , RI15b4adc0_419);
nor ( n45061 , n45059 , n45060 );
nand ( n45062 , n45058 , n45061 );
nor ( n45063 , n41824 , n41261 );
nor ( n45064 , n45057 , n45062 , n45063 );
not ( n45065 , n19876 );
nor ( n45066 , n45065 , n19922 );
or ( n45067 , n45066 , n41804 );
not ( n45068 , n19882 );
nand ( n45069 , n45067 , n45068 );
not ( n45070 , n41827 );
nand ( n45071 , n45065 , n45070 , n19882 );
nand ( n45072 , n45064 , n45069 , n45071 );
buf ( n45073 , n45072 );
buf ( n45074 , n22406 );
buf ( n45075 , n379893 );
not ( n45076 , n384318 );
not ( n45077 , n45076 );
not ( n45078 , n41771 );
or ( n45079 , n45077 , n45078 );
nand ( n45080 , n45079 , n32540 );
and ( n45081 , n45080 , n384392 );
xnor ( n45082 , n32553 , n384565 );
not ( n45083 , n380811 );
or ( n45084 , n45082 , n45083 );
not ( n45085 , n384441 );
not ( n45086 , n45085 );
not ( n45087 , n384435 );
or ( n45088 , n45086 , n45087 );
or ( n45089 , n384435 , n45085 );
nand ( n45090 , n45088 , n45089 );
and ( n45091 , n45090 , n384492 );
and ( n45092 , n19513 , RI15b640e0_1279);
nor ( n45093 , n45091 , n45092 );
nand ( n45094 , n45084 , n45093 );
nor ( n45095 , n45081 , n45094 );
or ( n45096 , n381593 , RI15b63168_1246);
nand ( n45097 , n45096 , n32581 );
and ( n45098 , n45097 , RI15b631e0_1247);
or ( n45099 , n384652 , n386842 , RI15b631e0_1247);
not ( n45100 , n386852 );
nand ( n45101 , n45100 , n19630 );
nand ( n45102 , n45099 , n45101 );
nor ( n45103 , n45098 , n45102 );
nand ( n45104 , n45095 , n45103 );
buf ( n45105 , n45104 );
not ( n45106 , n40468 );
not ( n45107 , n45106 );
not ( n45108 , n384726 );
or ( n45109 , n45107 , n45108 );
and ( n45110 , n384737 , n40470 );
or ( n45111 , n40480 , n20799 );
or ( n45112 , n384754 , n40485 );
or ( n45113 , n40478 , n384759 );
nand ( n45114 , n45111 , n45112 , n45113 );
nor ( n45115 , n45110 , n45114 );
nand ( n45116 , n45109 , n45115 );
buf ( n45117 , n45116 );
not ( n45118 , n37777 );
not ( n45119 , n45118 );
nor ( n45120 , n37771 , n37791 );
not ( n45121 , n45120 );
or ( n45122 , n45119 , n45121 );
not ( n45123 , n37783 );
nand ( n45124 , n45122 , n45123 );
not ( n45125 , RI15b61ae8_1198);
not ( n45126 , n45125 );
not ( n45127 , n37786 );
not ( n45128 , n45127 );
or ( n45129 , n45126 , n45128 );
nand ( n45130 , n45129 , RI15b61bd8_1200);
not ( n45131 , RI15b61b60_1199);
and ( n45132 , n45130 , n45131 );
not ( n45133 , n45130 );
and ( n45134 , n45133 , RI15b61b60_1199);
nor ( n45135 , n45132 , n45134 );
nand ( n45136 , n45124 , n45135 );
not ( n45137 , n45120 );
nor ( n45138 , n45135 , n384933 );
and ( n45139 , n45137 , n45138 );
not ( n45140 , RI15b5efc8_1106);
not ( n45141 , n384918 );
or ( n45142 , n45140 , n45141 );
not ( n45143 , n31054 );
nand ( n45144 , n384906 , n45143 );
nand ( n45145 , n45142 , n45144 );
nor ( n45146 , n45139 , n45145 );
nand ( n45147 , n45136 , n45146 );
buf ( n45148 , n45147 );
buf ( n45149 , n35649 );
buf ( n45150 , n381566 );
buf ( n45151 , n32672 );
not ( n45152 , n31841 );
not ( n45153 , n31832 );
not ( n45154 , n45153 );
or ( n45155 , n45152 , n45154 );
or ( n45156 , n45153 , n31841 );
nand ( n45157 , n45155 , n45156 );
buf ( n45158 , n35273 );
nand ( n45159 , n45157 , n45158 );
nor ( n45160 , n384388 , n31891 );
not ( n45161 , n45160 );
not ( n45162 , n31892 );
nand ( n45163 , n45161 , n45162 );
nand ( n45164 , n45163 , n31921 );
not ( n45165 , n31930 );
not ( n45166 , n31933 );
and ( n45167 , n45165 , n45166 );
not ( n45168 , n45165 );
and ( n45169 , n45168 , n31933 );
nor ( n45170 , n45167 , n45169 );
and ( n45171 , n45170 , n387121 );
nor ( n45172 , n19512 , n379448 );
nor ( n45173 , n45171 , n45172 );
and ( n45174 , n45159 , n45164 , n45173 );
not ( n45175 , n381572 );
or ( n45176 , n45175 , n383424 );
nand ( n45177 , n45176 , n384642 );
nand ( n45178 , n45177 , RI15b63780_1259);
and ( n45179 , n384655 , n383424 , n386767 );
and ( n45180 , n386771 , n19630 );
nor ( n45181 , n45179 , n45180 );
nand ( n45182 , n45174 , n45178 , n45181 );
buf ( n45183 , n45182 );
not ( n45184 , n32594 );
buf ( n45185 , n19798 );
not ( n45186 , n45185 );
or ( n45187 , n45184 , n45186 );
nand ( n45188 , n45187 , n22350 );
not ( n45189 , n19804 );
and ( n45190 , n45188 , n45189 );
or ( n45191 , n38996 , n20543 , RI15b4b720_439);
buf ( n45192 , n19971 );
or ( n45193 , n22362 , n45192 , RI15b49920_375);
nand ( n45194 , n45191 , n45193 );
nor ( n45195 , n45190 , n45194 );
not ( n45196 , n45189 );
not ( n45197 , n45185 );
nand ( n45198 , n45196 , n22368 , n45197 );
or ( n45199 , n384662 , n382109 );
and ( n45200 , n22378 , n45192 );
nor ( n45201 , n45200 , n22383 );
or ( n45202 , n45201 , n19972 );
nand ( n45203 , n45199 , n45202 );
nand ( n45204 , n45203 , n20501 );
and ( n45205 , n22388 , RI15b4b720_439);
and ( n45206 , n32621 , RI15b4a820_407);
nor ( n45207 , n45205 , n45206 , n383396 );
nand ( n45208 , n45195 , n45198 , n45204 , n45207 );
buf ( n45209 , n45208 );
buf ( n45210 , n22716 );
buf ( n45211 , n22402 );
buf ( n45212 , n383174 );
buf ( n45213 , n22406 );
buf ( n45214 , n22343 );
buf ( n45215 , n36704 );
buf ( n45216 , n22538 );
nor ( n45217 , n45216 , n17506 );
or ( n45218 , n45217 , n379905 );
nand ( n45219 , n45218 , n22544 );
not ( n45220 , n22591 );
nor ( n45221 , n45220 , n18079 );
or ( n45222 , n45221 , n18103 );
nand ( n45223 , n45222 , RI15b56418_808);
not ( n45224 , n22544 );
nand ( n45225 , n45216 , n379855 , n45224 );
nor ( n45226 , n18197 , RI15b56418_808);
and ( n45227 , n45220 , n45226 );
not ( n45228 , n22620 );
not ( n45229 , n18189 );
and ( n45230 , n45228 , n45229 );
nor ( n45231 , n45230 , n18179 );
or ( n45232 , n45231 , n22839 );
and ( n45233 , n18188 , n22620 , n22839 );
and ( n45234 , n18219 , RI15b57318_840);
nor ( n45235 , n45233 , n45234 );
nand ( n45236 , n45232 , n45235 );
nor ( n45237 , n45227 , n45236 );
nand ( n45238 , n45219 , n45223 , n45225 , n45237 );
buf ( n45239 , n45238 );
not ( n45240 , n385120 );
buf ( n45241 , n385119 );
not ( n45242 , n45241 );
or ( n45243 , n45240 , n45242 );
buf ( n45244 , n385121 );
not ( n45245 , n45244 );
nand ( n45246 , n45243 , n45245 );
and ( n45247 , n45246 , n385135 );
not ( n45248 , n21276 );
nor ( n45249 , n44734 , n21282 );
nand ( n45250 , n45248 , n45249 );
not ( n45251 , n21270 );
and ( n45252 , n45250 , n45251 );
not ( n45253 , n45250 );
and ( n45254 , n45253 , n21270 );
nor ( n45255 , n45252 , n45254 );
or ( n45256 , n45255 , n21358 );
not ( n45257 , n21484 );
not ( n45258 , n45257 );
nand ( n45259 , n44744 , n21494 );
not ( n45260 , n21490 );
nor ( n45261 , n45259 , n45260 );
not ( n45262 , n45261 );
or ( n45263 , n45258 , n45262 );
or ( n45264 , n45261 , n45257 );
nand ( n45265 , n45263 , n45264 );
and ( n45266 , n45265 , n22686 );
and ( n45267 , n21751 , RI15b57b88_858);
nor ( n45268 , n45266 , n45267 );
nand ( n45269 , n45256 , n45268 );
nor ( n45270 , n45247 , n45269 );
and ( n45271 , n21788 , RI15b56c88_826);
not ( n45272 , n21878 );
and ( n45273 , n45272 , n21769 );
not ( n45274 , n21872 );
and ( n45275 , n45274 , n21876 );
not ( n45276 , n45274 );
and ( n45277 , n45276 , RI15b56c88_826);
nor ( n45278 , n45275 , n45277 );
and ( n45279 , n45278 , n384113 );
nor ( n45280 , n45271 , n45273 , n45279 );
nand ( n45281 , n45270 , n45280 );
buf ( n45282 , n45281 );
buf ( n45283 , n32271 );
buf ( n45284 , n32271 );
buf ( n45285 , n382537 );
and ( n45286 , n379822 , RI15b659b8_1332);
and ( n45287 , n379825 , RI15b485e8_334);
nor ( n45288 , n45286 , n45287 );
nand ( n45289 , n379832 , RI15b468d8_272);
nand ( n45290 , n45288 , n45289 , n35179 );
buf ( n45291 , n45290 );
buf ( n45292 , n380865 );
buf ( n45293 , n382052 );
buf ( n45294 , n382065 );
buf ( n45295 , n31573 );
not ( n45296 , n45295 );
buf ( n45297 , n31580 );
not ( n45298 , n45297 );
and ( n45299 , n45296 , n45298 );
not ( n45300 , n45296 );
and ( n45301 , n45300 , n45297 );
nor ( n45302 , n45299 , n45301 );
not ( n45303 , n31599 );
not ( n45304 , n45303 );
nand ( n45305 , n45302 , n45304 );
not ( n45306 , n31357 );
nand ( n45307 , n42050 , n45306 );
nand ( n45308 , n45307 , n31700 );
nand ( n45309 , n45308 , n379229 );
or ( n45310 , n40971 , n45306 );
nand ( n45311 , n45310 , n42053 );
nand ( n45312 , n45311 , n31358 );
and ( n45313 , n379394 , RI15b57f48_866);
and ( n45314 , n31712 , RI15b51d50_657);
nor ( n45315 , n45313 , n45314 );
nand ( n45316 , n45305 , n45309 , n45312 , n45315 );
buf ( n45317 , n45316 );
buf ( n45318 , n35649 );
not ( n45319 , n31866 );
not ( n45320 , n31859 );
or ( n45321 , n45319 , n45320 );
or ( n45322 , n31859 , n31866 );
nand ( n45323 , n45321 , n45322 );
nand ( n45324 , n45323 , n31884 );
not ( n45325 , n31951 );
not ( n45326 , n31945 );
or ( n45327 , n45325 , n45326 );
or ( n45328 , n31945 , n31951 );
nand ( n45329 , n45327 , n45328 );
and ( n45330 , n45329 , n39045 );
nor ( n45331 , n19512 , n379451 );
nor ( n45332 , n45330 , n45331 );
nor ( n45333 , n31904 , n31910 );
not ( n45334 , n45333 );
nand ( n45335 , n45334 , n31911 );
nand ( n45336 , n45335 , n32549 );
and ( n45337 , n45324 , n45332 , n45336 );
and ( n45338 , n31792 , n31952 );
or ( n45339 , n31910 , n42117 );
not ( n45340 , RI15b5d150_1041);
or ( n45341 , n31771 , n45340 );
or ( n45342 , n31779 , n31866 );
nand ( n45343 , n45339 , n45341 , n45342 );
nor ( n45344 , n45338 , n45343 );
nand ( n45345 , n45337 , n45344 );
buf ( n45346 , n45345 );
buf ( n45347 , n22479 );
buf ( n45348 , n32981 );
buf ( n45349 , n387159 );
buf ( n45350 , n382049 );
and ( n45351 , n32747 , RI15b42a80_139);
not ( n45352 , n32749 );
and ( n45353 , n32753 , RI15b417c0_99);
and ( n45354 , n32762 , RI15b41400_91);
nor ( n45355 , n45353 , n45354 );
and ( n45356 , n32755 , RI15b41b80_107);
and ( n45357 , n32759 , RI15b41040_83);
nor ( n45358 , n45356 , n45357 );
and ( n45359 , n32766 , RI15b435c0_163);
and ( n45360 , n32768 , RI15b43200_155);
nor ( n45361 , n45359 , n45360 );
and ( n45362 , n32771 , RI15b43980_171);
and ( n45363 , n32773 , RI15b42e40_147);
nor ( n45364 , n45362 , n45363 );
nand ( n45365 , n45355 , n45358 , n45361 , n45364 );
and ( n45366 , n45352 , n45365 );
and ( n45367 , n32781 , RI15b40500_59);
nor ( n45368 , n45351 , n45366 , n45367 );
and ( n45369 , n32785 , RI15b426c0_131);
and ( n45370 , n32787 , RI15b42300_123);
nor ( n45371 , n45369 , n45370 );
and ( n45372 , n32792 , RI15b40140_51);
and ( n45373 , n32794 , RI15b41f40_115);
nor ( n45374 , n45372 , n45373 );
and ( n45375 , n32797 , RI15b408c0_67);
and ( n45376 , n32800 , RI15b40c80_75);
nor ( n45377 , n45375 , n45376 );
nand ( n45378 , n45368 , n45371 , n45374 , n45377 );
not ( n45379 , n45378 );
not ( n45380 , n32806 );
or ( n45381 , n45379 , n45380 );
and ( n45382 , n381055 , RI15b49998_376);
not ( n45383 , RI15b49998_376);
not ( n45384 , n36055 );
or ( n45385 , n45383 , n45384 );
or ( n45386 , n36055 , RI15b49998_376);
nand ( n45387 , n45385 , n45386 );
and ( n45388 , n381076 , n45387 );
nor ( n45389 , n45382 , n45388 );
nand ( n45390 , n45381 , n45389 );
buf ( n45391 , n45390 );
not ( n45392 , RI15b53f10_729);
not ( n45393 , n32244 );
or ( n45394 , n45392 , n45393 );
and ( n45395 , n32247 , RI15b65508_1322);
and ( n45396 , n32249 , RI15b60378_1148);
nor ( n45397 , n45395 , n45396 );
nand ( n45398 , n45394 , n45397 );
buf ( n45399 , n45398 );
buf ( n45400 , n386762 );
buf ( n45401 , n379847 );
buf ( n45402 , n387159 );
and ( n45403 , n35118 , n41027 , n35067 );
and ( n45404 , n20631 , RI15b46428_262);
nor ( n45405 , n45403 , n45404 );
nor ( n45406 , n41027 , n34930 );
or ( n45407 , n35114 , n45406 );
nand ( n45408 , n45407 , n41644 );
nand ( n45409 , n385213 , RI15b47a30_309);
nand ( n45410 , n45405 , n45408 , n45409 );
buf ( n45411 , n45410 );
buf ( n45412 , n385195 );
buf ( n45413 , n385197 );
buf ( n45414 , n381021 );
not ( n45415 , n38492 );
or ( n45416 , n45415 , n386998 );
not ( n45417 , n38753 );
not ( n45418 , n45417 );
not ( n45419 , n38782 );
and ( n45420 , n45418 , n45419 );
and ( n45421 , n45417 , n38782 );
nor ( n45422 , n45420 , n45421 );
not ( n45423 , n45422 );
not ( n45424 , n386747 );
and ( n45425 , n45423 , n45424 );
and ( n45426 , n38496 , n38493 );
nor ( n45427 , n45425 , n45426 );
nand ( n45428 , n45416 , n45427 );
buf ( n45429 , n45428 );
buf ( n45430 , n381872 );
buf ( n45431 , n385112 );
or ( n45432 , n386705 , n38825 );
and ( n45433 , n386716 , n38828 );
or ( n45434 , n38837 , n17860 );
not ( n45435 , n37442 );
or ( n45436 , n45435 , n38841 );
or ( n45437 , n38835 , n386738 );
nand ( n45438 , n45434 , n45436 , n45437 );
nor ( n45439 , n45433 , n45438 );
nand ( n45440 , n45432 , n45439 );
buf ( n45441 , n45440 );
or ( n45442 , n36937 , n41443 );
and ( n45443 , n36946 , n41446 );
or ( n45444 , n41455 , n17806 );
or ( n45445 , n38403 , n41461 );
or ( n45446 , n41453 , n36955 );
nand ( n45447 , n45444 , n45445 , n45446 );
nor ( n45448 , n45443 , n45447 );
nand ( n45449 , n45442 , n45448 );
buf ( n45450 , n45449 );
buf ( n45451 , n19653 );
or ( n45452 , n31091 , n32320 );
and ( n45453 , n45016 , n39367 );
or ( n45454 , n31052 , n380656 );
not ( n45455 , n31078 );
not ( n45456 , n41417 );
and ( n45457 , n45456 , RI15b61638_1188);
not ( n45458 , n45456 );
and ( n45459 , n45458 , n32320 );
nor ( n45460 , n45457 , n45459 );
or ( n45461 , n45455 , n45460 );
nand ( n45462 , n384906 , n382956 );
nand ( n45463 , n45454 , n45461 , n45462 );
nor ( n45464 , n45453 , n45463 );
nand ( n45465 , n45452 , n45464 );
buf ( n45466 , n45465 );
buf ( n45467 , n382065 );
buf ( n45468 , n384203 );
buf ( n45469 , n33382 );
buf ( n45470 , n20665 );
and ( n45471 , n382668 , RI15b55518_776);
not ( n45472 , n382668 );
and ( n45473 , n45472 , n382669 );
nor ( n45474 , n45471 , n45473 );
or ( n45475 , n45474 , n382629 );
nand ( n45476 , n386637 , RI15b55518_776);
and ( n45477 , n382692 , n383784 );
and ( n45478 , n382885 , n38029 );
nor ( n45479 , n45477 , n45478 , n44221 );
nand ( n45480 , n45475 , n45476 , n45479 );
buf ( n45481 , n45480 );
buf ( n45482 , n22408 );
not ( n45483 , n382898 );
not ( n45484 , n381507 );
or ( n45485 , n45483 , n45484 );
and ( n45486 , n381524 , n382934 );
not ( n45487 , RI15b59988_922);
or ( n45488 , n382949 , n45487 );
or ( n45489 , n381551 , n382965 );
or ( n45490 , n382947 , n381560 );
nand ( n45491 , n45488 , n45489 , n45490 );
nor ( n45492 , n45486 , n45491 );
nand ( n45493 , n45485 , n45492 );
buf ( n45494 , n45493 );
not ( n45495 , RI15b50130_597);
or ( n45496 , n385163 , n45495 );
and ( n45497 , n36472 , n21597 );
not ( n45498 , n21098 );
and ( n45499 , n35704 , n45498 );
buf ( n45500 , n21211 );
nor ( n45501 , n45499 , n45500 );
buf ( n45502 , n21214 );
not ( n45503 , n45502 );
and ( n45504 , n45501 , n45503 );
buf ( n45505 , n21023 );
not ( n45506 , n45505 );
nor ( n45507 , n45504 , n45506 );
and ( n45508 , n21219 , n45507 );
not ( n45509 , n21219 );
not ( n45510 , n45501 );
and ( n45511 , n45510 , n45505 );
nor ( n45512 , n45511 , n45502 );
and ( n45513 , n45509 , n45512 );
nor ( n45514 , n45508 , n45513 );
not ( n45515 , n37447 );
and ( n45516 , n45514 , n45515 );
not ( n45517 , n45514 );
and ( n45518 , n45517 , n37447 );
nor ( n45519 , n45516 , n45518 );
or ( n45520 , n45519 , n44740 );
not ( n45521 , n21439 );
not ( n45522 , n39069 );
or ( n45523 , n45521 , n45522 );
or ( n45524 , n39069 , n21439 );
nand ( n45525 , n45523 , n45524 );
not ( n45526 , n37447 );
and ( n45527 , n45525 , n45526 );
not ( n45528 , n45525 );
and ( n45529 , n45528 , n37447 );
nor ( n45530 , n45527 , n45529 );
not ( n45531 , n21559 );
or ( n45532 , n45530 , n45531 );
not ( n45533 , n21625 );
nor ( n45534 , n45533 , n21599 );
not ( n45535 , n45534 );
not ( n45536 , n37825 );
not ( n45537 , n45536 );
or ( n45538 , n45535 , n45537 );
or ( n45539 , n45536 , n45534 );
nand ( n45540 , n45538 , n45539 );
and ( n45541 , n45540 , n21742 );
and ( n45542 , n21751 , RI15b577c8_850);
nor ( n45543 , n45541 , n45542 );
nand ( n45544 , n45520 , n45532 , n45543 );
nor ( n45545 , n45497 , n45544 );
and ( n45546 , n32368 , n21219 );
and ( n45547 , n385177 , n21439 );
nor ( n45548 , n45546 , n45547 );
nand ( n45549 , n45496 , n45545 , n45548 );
buf ( n45550 , n45549 );
not ( n45551 , n37773 );
not ( n45552 , n33569 );
not ( n45553 , n45552 );
or ( n45554 , n45551 , n45553 );
not ( n45555 , n37779 );
nand ( n45556 , n45554 , n45555 );
nand ( n45557 , n45556 , n33573 );
not ( n45558 , n33573 );
nand ( n45559 , n45558 , n384934 );
nor ( n45560 , n45552 , n45559 );
and ( n45561 , n384918 , RI15b5ed70_1101);
nor ( n45562 , n45560 , n45561 , n43066 );
nand ( n45563 , n45557 , n45562 );
buf ( n45564 , n45563 );
buf ( n45565 , n379844 );
buf ( n45566 , n379893 );
buf ( n45567 , n22404 );
buf ( n45568 , n32160 );
buf ( n45569 , RI15b5db28_1062);
buf ( n45570 , n381707 );
buf ( n45571 , n386832 );
or ( n45572 , n45571 , n22473 );
nand ( n45573 , n45572 , n383474 );
nand ( n45574 , n45573 , n386838 );
not ( n45575 , n386838 );
not ( n45576 , n34843 );
nand ( n45577 , n45575 , n45576 , n45571 );
not ( n45578 , n42188 );
buf ( n45579 , n386971 );
and ( n45580 , n45578 , n45579 );
nor ( n45581 , n45580 , n40140 );
or ( n45582 , n45581 , n386972 );
and ( n45583 , n40145 , RI15b63ff0_1277);
or ( n45584 , n34826 , n45579 , RI15b621f0_1213);
not ( n45585 , n387031 );
not ( n45586 , n45585 );
not ( n45587 , RI15b63ff0_1277);
and ( n45588 , n45586 , n45587 );
and ( n45589 , n45585 , RI15b63ff0_1277);
nor ( n45590 , n45588 , n45589 );
or ( n45591 , n34833 , n45590 );
nand ( n45592 , n45584 , n45591 );
nor ( n45593 , n45583 , n45592 );
nand ( n45594 , n45582 , n45593 );
nand ( n45595 , n45594 , n19201 );
and ( n45596 , n22423 , RI15b63ff0_1277);
and ( n45597 , n19599 , RI15b630f0_1245);
nor ( n45598 , n45596 , n45597 , n19513 );
nand ( n45599 , n45574 , n45577 , n45595 , n45598 );
buf ( n45600 , n45599 );
buf ( n45601 , n22738 );
buf ( n45602 , n385937 );
and ( n45603 , n45602 , n385946 );
not ( n45604 , n45602 );
not ( n45605 , n385946 );
and ( n45606 , n45604 , n45605 );
nor ( n45607 , n45603 , n45606 );
and ( n45608 , n45607 , n386019 );
buf ( n45609 , n386230 );
not ( n45610 , n386234 );
and ( n45611 , n45609 , n45610 );
not ( n45612 , n45609 );
and ( n45613 , n45612 , n386234 );
nor ( n45614 , n45611 , n45613 );
or ( n45615 , n45614 , n34766 );
not ( n45616 , n386487 );
not ( n45617 , n386479 );
not ( n45618 , n386486 );
nand ( n45619 , n45617 , n45618 );
nand ( n45620 , n45616 , n45619 );
and ( n45621 , n45620 , n386500 );
nor ( n45622 , n34782 , n382135 );
nor ( n45623 , n45621 , n45622 );
nand ( n45624 , n45615 , n45623 );
nor ( n45625 , n45608 , n45624 );
not ( n45626 , n20637 );
not ( n45627 , n19695 );
or ( n45628 , n45626 , n45627 );
nand ( n45629 , n45628 , n34798 );
and ( n45630 , n45629 , RI15b4aeb0_421);
or ( n45631 , n34801 , n19695 , RI15b4aeb0_421);
not ( n45632 , n19897 );
or ( n45633 , n45632 , n22216 );
nand ( n45634 , n45631 , n45633 );
nor ( n45635 , n45630 , n45634 );
nand ( n45636 , n45625 , n45635 );
buf ( n45637 , n45636 );
buf ( n45638 , n385197 );
buf ( n45639 , n32672 );
buf ( n45640 , n22005 );
nor ( n45641 , n44770 , n34930 );
or ( n45642 , n45641 , n35114 );
nand ( n45643 , n45642 , n44775 );
nor ( n45644 , n35117 , n44774 );
and ( n45645 , n44770 , n45644 );
and ( n45646 , n385213 , RI15b47b98_312);
and ( n45647 , n20631 , RI15b46590_265);
nor ( n45648 , n45646 , n45647 );
not ( n45649 , n45648 );
nor ( n45650 , n45645 , n45649 );
nand ( n45651 , n45643 , n45650 );
buf ( n45652 , n45651 );
buf ( n45653 , n387159 );
buf ( n45654 , n35651 );
buf ( n45655 , n382069 );
buf ( n45656 , n33250 );
or ( n45657 , n36238 , n384738 );
or ( n45658 , n17984 , n384749 );
not ( n45659 , n384757 );
and ( n45660 , n45659 , n36257 );
and ( n45661 , n383803 , n384705 );
and ( n45662 , n36261 , n384755 );
nor ( n45663 , n45660 , n45661 , n45662 );
nand ( n45664 , n45657 , n45658 , n45663 );
buf ( n45665 , n45664 );
nand ( n45666 , n384914 , n31055 );
nand ( n45667 , n384918 , RI15b5f6d0_1121);
nand ( n45668 , n383575 , n383586 );
or ( n45669 , n44042 , n45668 );
nand ( n45670 , n45669 , n44044 );
not ( n45671 , n32278 );
nor ( n45672 , n45671 , n383523 );
and ( n45673 , n45672 , RI15b613e0_1183);
not ( n45674 , n45672 );
and ( n45675 , n45674 , n31130 );
nor ( n45676 , n45673 , n45675 );
and ( n45677 , n45670 , n45676 );
not ( n45678 , n45676 );
and ( n45679 , n45668 , n45678 );
and ( n45680 , n384934 , n45679 );
nor ( n45681 , n45677 , n45680 );
nand ( n45682 , n31059 , n45666 , n45667 , n45681 );
buf ( n45683 , n45682 );
buf ( n45684 , n380903 );
buf ( n45685 , n19651 );
buf ( n45686 , n381006 );
and ( n45687 , n379822 , n43158 );
nor ( n45688 , n379834 , n381978 );
nor ( n45689 , n45687 , n45688 );
nand ( n45690 , n379832 , RI15b46c20_279);
nand ( n45691 , n379825 , RI15b48930_341);
nand ( n45692 , n45689 , n45690 , n45691 );
buf ( n45693 , n45692 );
buf ( n45694 , n382049 );
buf ( n45695 , n22788 );
or ( n45696 , n386588 , n32063 );
and ( n45697 , n386600 , n32070 );
or ( n45698 , n32081 , n19174 );
or ( n45699 , n386618 , n32086 );
or ( n45700 , n32079 , n386627 );
nand ( n45701 , n45698 , n45699 , n45700 );
nor ( n45702 , n45697 , n45701 );
nand ( n45703 , n45696 , n45702 );
buf ( n45704 , n45703 );
buf ( n45705 , n22738 );
buf ( n45706 , n382065 );
or ( n45707 , n32430 , n35491 );
buf ( n45708 , n382639 );
not ( n45709 , n45708 );
not ( n45710 , n382626 );
or ( n45711 , n45709 , n45710 );
nand ( n45712 , n45711 , n382679 );
and ( n45713 , n45712 , RI15b54c30_757);
or ( n45714 , n386674 , n45708 , RI15b54c30_757);
not ( n45715 , n22679 );
or ( n45716 , n382886 , n45715 );
nand ( n45717 , n45714 , n45716 );
nor ( n45718 , n45713 , n45717 );
and ( n45719 , n37522 , n45718 );
nand ( n45720 , n45707 , n45719 );
buf ( n45721 , n45720 );
or ( n45722 , n40936 , n19200 );
not ( n45723 , n31759 );
or ( n45724 , n45723 , n19200 );
nand ( n45725 , n45724 , RI15b5d510_1049);
not ( n45726 , n19573 );
nand ( n45727 , n45722 , n45725 , n45726 );
buf ( n45728 , n45727 );
buf ( n45729 , n22788 );
not ( n45730 , n43986 );
and ( n45731 , n45730 , n43987 );
not ( n45732 , n45730 );
and ( n45733 , n45732 , n43988 );
nor ( n45734 , n45731 , n45733 );
not ( n45735 , n31600 );
nand ( n45736 , n45734 , n45735 );
or ( n45737 , n40962 , n31667 );
nand ( n45738 , n45737 , n31700 );
and ( n45739 , n45738 , n31644 );
not ( n45740 , n40962 );
or ( n45741 , n39677 , n45740 , n31644 );
and ( n45742 , n379394 , RI15b57b88_858);
and ( n45743 , n31712 , RI15b51990_649);
nor ( n45744 , n45742 , n45743 );
nand ( n45745 , n45741 , n45744 );
nor ( n45746 , n45739 , n45745 );
nand ( n45747 , n45736 , n45746 );
buf ( n45748 , n45747 );
buf ( n45749 , n22406 );
or ( n45750 , n383814 , n33597 );
and ( n45751 , n383857 , n33600 );
not ( n45752 , RI15b4e948_546);
or ( n45753 , n33609 , n45752 );
or ( n45754 , n41458 , n33615 );
or ( n45755 , n33607 , n383917 );
nand ( n45756 , n45753 , n45754 , n45755 );
nor ( n45757 , n45751 , n45756 );
nand ( n45758 , n45750 , n45757 );
buf ( n45759 , n45758 );
buf ( n45760 , n380942 );
buf ( n45761 , n383174 );
not ( n45762 , n40774 );
nor ( n45763 , n37771 , n45762 );
or ( n45764 , n45763 , n33585 );
nand ( n45765 , n45764 , n37792 );
nor ( n45766 , n37791 , n33588 );
not ( n45767 , n45766 );
not ( n45768 , n37771 );
or ( n45769 , n45767 , n45768 );
and ( n45770 , n383601 , RI15b60558_1152);
and ( n45771 , n383607 , RI15b5ef50_1105);
nor ( n45772 , n45770 , n45771 );
nand ( n45773 , n45769 , n45772 );
not ( n45774 , n45773 );
nand ( n45775 , n45765 , n45774 );
buf ( n45776 , n45775 );
buf ( n45777 , n33250 );
buf ( n45778 , n379844 );
buf ( n45779 , n380203 );
buf ( n45780 , n382052 );
buf ( n45781 , n22655 );
not ( n45782 , n386111 );
or ( n45783 , n39290 , n45782 );
and ( n45784 , n386540 , RI15b43b60_175);
or ( n45785 , n386550 , RI15b43b60_175);
nand ( n45786 , n45785 , n42751 );
nor ( n45787 , n45784 , n45786 );
nand ( n45788 , n45783 , n45787 );
buf ( n45789 , n45788 );
or ( n45790 , n381907 , n35869 );
and ( n45791 , n39450 , RI15b40b18_72);
or ( n45792 , n381917 , n35871 );
not ( n45793 , n35888 );
and ( n45794 , n45793 , n381923 );
and ( n45795 , n381926 , n35886 );
nor ( n45796 , n45794 , n45795 );
nand ( n45797 , n45792 , n45796 );
nor ( n45798 , n45791 , n45797 );
nand ( n45799 , n45790 , n45798 );
buf ( n45800 , n45799 );
or ( n45801 , n380968 , n35895 );
and ( n45802 , n380986 , n39462 );
not ( n45803 , RI15b40500_59);
or ( n45804 , n35911 , n45803 );
or ( n45805 , n380994 , n35917 );
or ( n45806 , n35909 , n380996 );
nand ( n45807 , n45804 , n45805 , n45806 );
nor ( n45808 , n45802 , n45807 );
nand ( n45809 , n45801 , n45808 );
buf ( n45810 , n45809 );
buf ( n45811 , n22009 );
buf ( n45812 , n35651 );
buf ( n45813 , n22653 );
buf ( n45814 , n384996 );
buf ( n45815 , n379895 );
buf ( n45816 , n380940 );
and ( n45817 , n379822 , RI15b65b98_1336);
and ( n45818 , n379825 , RI15b487c8_338);
nor ( n45819 , n45817 , n45818 );
nand ( n45820 , n379832 , RI15b46ab8_276);
nand ( n45821 , n45819 , n45820 , n39273 );
buf ( n45822 , n45821 );
buf ( n45823 , n380865 );
buf ( n45824 , n381021 );
buf ( n45825 , n379403 );
buf ( n45826 , n18226 );
not ( n45827 , n382664 );
not ( n45828 , n386674 );
and ( n45829 , n45827 , n45828 );
nor ( n45830 , n45829 , n386637 );
or ( n45831 , n45830 , n382666 );
nor ( n45832 , n386674 , RI15b55428_774);
and ( n45833 , n382664 , n45832 );
or ( n45834 , n380167 , n380192 );
nand ( n45835 , n45834 , n35736 , n380193 );
or ( n45836 , n35730 , n45835 );
or ( n45837 , n382691 , n383669 );
nand ( n45838 , n45836 , n45837 );
nor ( n45839 , n45833 , n38905 , n45838 );
nand ( n45840 , n45831 , n45839 );
buf ( n45841 , n45840 );
or ( n45842 , n383180 , n35792 );
not ( n45843 , n35803 );
and ( n45844 , n45843 , RI15b59a78_924);
or ( n45845 , n383184 , n35789 );
and ( n45846 , n35810 , n41701 );
and ( n45847 , n40019 , n35807 );
nor ( n45848 , n45846 , n45847 );
nand ( n45849 , n45845 , n45848 );
nor ( n45850 , n45844 , n45849 );
nand ( n45851 , n45842 , n45850 );
buf ( n45852 , n45851 );
buf ( n45853 , n22655 );
not ( n45854 , n35233 );
nand ( n45855 , n40305 , RI15b54780_747);
nand ( n45856 , n45854 , n45855 );
and ( n45857 , n45856 , RI15b3fab0_37);
and ( n45858 , n37567 , n43294 );
nor ( n45859 , n45858 , n17505 );
nor ( n45860 , n45857 , n45859 , n37571 );
not ( n45861 , n45860 );
buf ( n45862 , n45861 );
buf ( n45863 , n22009 );
buf ( n45864 , n380865 );
not ( n45865 , n32680 );
not ( n45866 , n381589 );
or ( n45867 , n45865 , n45866 );
and ( n45868 , n381596 , n35222 );
or ( n45869 , n32692 , n18705 );
or ( n45870 , n42258 , n32699 );
or ( n45871 , n32690 , n381621 );
nand ( n45872 , n45869 , n45870 , n45871 );
nor ( n45873 , n45868 , n45872 );
nand ( n45874 , n45867 , n45873 );
buf ( n45875 , n45874 );
buf ( n45876 , n22007 );
buf ( n45877 , n31719 );
or ( n45878 , n36735 , n20519 );
or ( n45879 , n39256 , n20425 );
and ( n45880 , n386110 , n43641 );
and ( n45881 , n386066 , RI15b44970_205);
nor ( n45882 , n45880 , n45881 );
or ( n45883 , n45882 , n36114 );
or ( n45884 , n36723 , n22298 );
nand ( n45885 , n45879 , n45883 , n45884 );
not ( n45886 , n45885 );
nand ( n45887 , n45878 , n45886 );
buf ( n45888 , n45887 );
buf ( n45889 , n382067 );
buf ( n45890 , n380865 );
buf ( n45891 , n385197 );
buf ( n45892 , n385112 );
not ( n45893 , n42765 );
and ( n45894 , n383945 , RI15b58920_887);
and ( n45895 , n383949 , RI15b5a720_951);
nor ( n45896 , n45894 , n45895 );
and ( n45897 , n383955 , RI15b5aea0_967);
and ( n45898 , n383960 , RI15b5aae0_959);
nor ( n45899 , n45897 , n45898 );
and ( n45900 , n383965 , RI15b5b260_975);
and ( n45901 , n383970 , RI15b59fa0_935);
and ( n45902 , n383972 , RI15b5a360_943);
nor ( n45903 , n45901 , n45902 );
and ( n45904 , n383975 , RI15b59820_919);
and ( n45905 , n383977 , RI15b59be0_927);
nor ( n45906 , n45904 , n45905 );
and ( n45907 , n383982 , RI15b5bda0_999);
and ( n45908 , n383984 , RI15b5b9e0_991);
nor ( n45909 , n45907 , n45908 );
and ( n45910 , n383987 , RI15b5c160_1007);
and ( n45911 , n383989 , RI15b5b620_983);
nor ( n45912 , n45910 , n45911 );
nand ( n45913 , n45903 , n45906 , n45909 , n45912 );
and ( n45914 , n383968 , n45913 );
and ( n45915 , n383994 , RI15b58ce0_895);
nor ( n45916 , n45900 , n45914 , n45915 );
and ( n45917 , n383997 , RI15b590a0_903);
and ( n45918 , n383999 , RI15b59460_911);
nor ( n45919 , n45917 , n45918 );
nand ( n45920 , n45896 , n45899 , n45916 , n45919 );
not ( n45921 , n45920 );
or ( n45922 , n45893 , n45921 );
not ( n45923 , n38471 );
not ( n45924 , n45923 );
not ( n45925 , n384025 );
or ( n45926 , n45924 , n45925 );
nand ( n45927 , n45926 , n384021 );
and ( n45928 , n45927 , RI15b62178_1212);
nor ( n45929 , n45923 , RI15b62178_1212);
and ( n45930 , n384025 , n45929 );
nor ( n45931 , n45928 , n45930 );
nand ( n45932 , n45922 , n45931 );
buf ( n45933 , n45932 );
and ( n45934 , n22646 , RI15b45258_224);
and ( n45935 , n22648 , RI15b516c0_643);
nor ( n45936 , n45934 , n45935 );
not ( n45937 , n45936 );
buf ( n45938 , n45937 );
or ( n45939 , n36937 , n384057 );
and ( n45940 , n36946 , n384169 );
or ( n45941 , n384182 , n17810 );
or ( n45942 , n36952 , n384190 );
or ( n45943 , n384180 , n36955 );
nand ( n45944 , n45941 , n45942 , n45943 );
nor ( n45945 , n45940 , n45944 );
nand ( n45946 , n45939 , n45945 );
buf ( n45947 , n45946 );
buf ( n45948 , n384199 );
buf ( n45949 , n32981 );
not ( n45950 , RI15b46f68_286);
not ( n45951 , n385213 );
or ( n45952 , n45950 , n45951 );
and ( n45953 , n385221 , RI15b484f8_332);
and ( n45954 , n20631 , RI15b467e8_270);
nor ( n45955 , n45953 , n45954 );
nand ( n45956 , n45952 , n45955 );
buf ( n45957 , n45956 );
buf ( n45958 , n32160 );
buf ( n45959 , n383174 );
buf ( n45960 , n33382 );
buf ( n45961 , n386762 );
buf ( n45962 , n381004 );
buf ( n45963 , n383174 );
buf ( n45964 , RI15b5e6e0_1087);
or ( n45965 , n42942 , n36306 );
and ( n45966 , n384983 , n36309 );
or ( n45967 , n36318 , n385374 );
or ( n45968 , n22022 , n36325 );
or ( n45969 , n36316 , n384988 );
nand ( n45970 , n45967 , n45968 , n45969 );
nor ( n45971 , n45966 , n45970 );
nand ( n45972 , n45965 , n45971 );
buf ( n45973 , n45972 );
buf ( n45974 , n384199 );
buf ( n45975 , n383345 );
buf ( n45976 , n32676 );
not ( n45977 , n17507 );
not ( n45978 , n22565 );
or ( n45979 , n45977 , n45978 );
nand ( n45980 , n45979 , n17565 );
nand ( n45981 , n45980 , n41161 );
nor ( n45982 , n22599 , n18079 );
or ( n45983 , n45982 , n18103 );
nand ( n45984 , n45983 , RI15b565f8_812);
nand ( n45985 , n22566 , n22574 );
nor ( n45986 , n18197 , RI15b565f8_812);
and ( n45987 , n22599 , n45986 );
or ( n45988 , n22604 , n379043 );
xor ( n45989 , RI15b583f8_876 , n22624 );
and ( n45990 , n45989 , n18188 );
and ( n45991 , n18219 , RI15b574f8_844);
nor ( n45992 , n45990 , n45991 );
nand ( n45993 , n45988 , n45992 );
nor ( n45994 , n45987 , n45993 );
nand ( n45995 , n45981 , n45984 , n45985 , n45994 );
buf ( n45996 , n45995 );
buf ( n45997 , RI15b45f78_252);
buf ( n45998 , n22005 );
and ( n45999 , n21573 , n22690 );
not ( n46000 , n21662 );
or ( n46001 , n45999 , n46000 );
buf ( n46002 , n385114 );
nand ( n46003 , n46001 , n46002 );
and ( n46004 , n46003 , n385133 );
buf ( n46005 , n21238 );
not ( n46006 , n46005 );
not ( n46007 , n21254 );
and ( n46008 , n46006 , n46007 );
and ( n46009 , n46005 , n21254 );
nor ( n46010 , n46008 , n46009 );
or ( n46011 , n46010 , n44740 );
not ( n46012 , n21471 );
not ( n46013 , n21467 );
not ( n46014 , n46013 );
or ( n46015 , n46012 , n46014 );
or ( n46016 , n46013 , n21471 );
nand ( n46017 , n46015 , n46016 );
and ( n46018 , n46017 , n21559 );
and ( n46019 , n21751 , RI15b579a8_854);
nor ( n46020 , n46018 , n46019 );
nand ( n46021 , n46011 , n46020 );
nor ( n46022 , n46004 , n46021 );
and ( n46023 , n21788 , RI15b56aa8_822);
and ( n46024 , n21846 , n39103 );
and ( n46025 , n21840 , n21838 );
not ( n46026 , n21840 );
and ( n46027 , n46026 , RI15b56aa8_822);
nor ( n46028 , n46025 , n46027 );
and ( n46029 , n46028 , n21794 );
nor ( n46030 , n46023 , n46024 , n46029 );
nand ( n46031 , n46022 , n46030 );
buf ( n46032 , n46031 );
buf ( n46033 , n22655 );
buf ( n46034 , n381021 );
buf ( n46035 , n22404 );
buf ( n46036 , n40996 );
or ( n46037 , n46036 , n41015 );
nand ( n46038 , n46037 , n41032 );
nand ( n46039 , n46038 , n35087 );
and ( n46040 , n46036 , n35088 );
nand ( n46041 , n41651 , n46040 );
nand ( n46042 , n41582 , RI15b461d0_257);
and ( n46043 , n35459 , n22278 );
and ( n46044 , n35461 , RI15b659b8_1332);
nor ( n46045 , n46043 , n46044 );
nand ( n46046 , n46039 , n46041 , n46042 , n46045 );
buf ( n46047 , n46046 );
buf ( n46048 , n381566 );
buf ( n46049 , n35651 );
buf ( n46050 , n382049 );
buf ( n46051 , n379844 );
buf ( n46052 , n32981 );
not ( n46053 , RI15b479b8_308);
not ( n46054 , n385213 );
or ( n46055 , n46053 , n46054 );
and ( n46056 , n41013 , n34931 );
and ( n46057 , n20631 , RI15b463b0_261);
nor ( n46058 , n46056 , n46057 );
nand ( n46059 , n46055 , n46058 );
buf ( n46060 , n46059 );
buf ( n46061 , n380903 );
or ( n46062 , n36937 , n36242 );
and ( n46063 , n36946 , n43075 );
not ( n46064 , RI15b4d4a8_502);
or ( n46065 , n36250 , n46064 );
or ( n46066 , n41326 , n36254 );
or ( n46067 , n36248 , n36955 );
nand ( n46068 , n46065 , n46066 , n46067 );
nor ( n46069 , n46063 , n46068 );
nand ( n46070 , n46062 , n46069 );
buf ( n46071 , n46070 );
buf ( n46072 , n35649 );
buf ( n46073 , RI15b472b0_293);
buf ( n46074 , n386760 );
nand ( n46075 , n31128 , n33492 );
nand ( n46076 , n44454 , n46075 );
not ( n46077 , n46076 );
not ( n46078 , RI15b619f8_1196);
or ( n46079 , n46077 , n46078 );
nand ( n46080 , n43062 , RI15b61908_1194 , RI15b61980_1195);
or ( n46081 , RI15b619f8_1196 , n46080 );
not ( n46082 , n38553 );
not ( n46083 , n38752 );
or ( n46084 , n46082 , n46083 );
or ( n46085 , n38752 , n38553 );
nand ( n46086 , n46084 , n46085 );
buf ( n46087 , n44459 );
not ( n46088 , n46087 );
and ( n46089 , n46086 , n46088 );
nor ( n46090 , n42641 , n380364 );
nor ( n46091 , n31052 , n380575 );
nor ( n46092 , n46089 , n46090 , n46091 );
nand ( n46093 , n46079 , n46081 , n46092 );
buf ( n46094 , n46093 );
buf ( n46095 , n381707 );
or ( n46096 , n41514 , n34937 );
and ( n46097 , n35537 , RI15b43110_153);
and ( n46098 , n41517 , RI15b42d50_145);
nor ( n46099 , n46097 , n46098 );
and ( n46100 , n35376 , RI15b43890_169);
and ( n46101 , n35373 , RI15b434d0_161);
nor ( n46102 , n46100 , n46101 );
and ( n46103 , n41523 , RI15b40b90_73);
and ( n46104 , n41525 , RI15b407d0_65);
nor ( n46105 , n46103 , n46104 );
or ( n46106 , n41531 , n381058 );
and ( n46107 , n35448 , RI15b41310_89);
and ( n46108 , n35441 , RI15b40f50_81);
and ( n46109 , n37311 , RI15b416d0_97);
nor ( n46110 , n46108 , n46109 );
and ( n46111 , n35422 , RI15b41a90_105);
and ( n46112 , n35412 , RI15b41e50_113);
nor ( n46113 , n46111 , n46112 );
and ( n46114 , n35415 , RI15b42990_137);
and ( n46115 , n35555 , RI15b425d0_129);
nor ( n46116 , n46114 , n46115 );
nand ( n46117 , n46110 , n46113 , n46116 );
not ( n46118 , RI15b42210_121);
nor ( n46119 , n35390 , n46118 );
nor ( n46120 , n46107 , n46117 , n46119 );
or ( n46121 , n46120 , n32749 );
not ( n46122 , RI15b40410_57);
or ( n46123 , n46122 , n41528 );
nand ( n46124 , n46106 , n46121 , n46123 );
not ( n46125 , n46124 );
nand ( n46126 , n46099 , n46102 , n46105 , n46125 );
not ( n46127 , n35456 );
and ( n46128 , n46126 , n46127 );
and ( n46129 , n35335 , RI15b66138_1348);
nor ( n46130 , n35357 , n35195 , RI15b48d68_350);
nor ( n46131 , n46128 , n46129 , n46130 );
nand ( n46132 , n46096 , n46131 , n46045 );
buf ( n46133 , n46132 );
buf ( n46134 , n381081 );
buf ( n46135 , n384199 );
or ( n46136 , n381015 , n22041 );
nand ( n46137 , n35525 , RI15b53c40_723);
nand ( n46138 , n46136 , n46137 );
buf ( n46139 , n46138 );
buf ( n46140 , n380906 );
buf ( n46141 , n22406 );
buf ( n46142 , n22788 );
buf ( n46143 , n33250 );
buf ( n46144 , n384996 );
or ( n46145 , n31006 , n35622 );
and ( n46146 , n31016 , n35625 );
or ( n46147 , n35635 , n21000 );
or ( n46148 , n40593 , n35640 );
or ( n46149 , n35633 , n31024 );
nand ( n46150 , n46147 , n46148 , n46149 );
nor ( n46151 , n46146 , n46150 );
nand ( n46152 , n46145 , n46151 );
buf ( n46153 , n46152 );
not ( n46154 , RI15b5f928_1126);
not ( n46155 , n383601 );
or ( n46156 , n46154 , n46155 );
and ( n46157 , n383505 , RI15b60eb8_1172);
and ( n46158 , n383607 , RI15b5f1a8_1110);
nor ( n46159 , n46157 , n46158 );
nand ( n46160 , n46156 , n46159 );
buf ( n46161 , n46160 );
not ( n46162 , RI15b536a0_711);
not ( n46163 , n383170 );
or ( n46164 , n46162 , n46163 );
not ( n46165 , n381439 );
not ( n46166 , n33453 );
or ( n46167 , n46165 , n46166 );
nand ( n46168 , n46167 , n33465 );
and ( n46169 , n46168 , n37528 );
and ( n46170 , n33476 , n37530 );
and ( n46171 , n383147 , RI15b52f20_695);
nor ( n46172 , n46169 , n46170 , n46171 );
nand ( n46173 , n46164 , n46172 );
buf ( n46174 , n46173 );
buf ( n46175 , n35649 );
buf ( n46176 , n380942 );
not ( n46177 , n33387 );
not ( n46178 , n380703 );
or ( n46179 , n46177 , n46178 );
and ( n46180 , n380719 , n33417 );
not ( n46181 , RI15b5b800_987);
or ( n46182 , n33428 , n46181 );
not ( n46183 , n380781 );
or ( n46184 , n46183 , n33440 );
or ( n46185 , n33426 , n380790 );
nand ( n46186 , n46182 , n46184 , n46185 );
nor ( n46187 , n46180 , n46186 );
nand ( n46188 , n46179 , n46187 );
buf ( n46189 , n46188 );
buf ( n46190 , n379802 );
buf ( n46191 , n382073 );
or ( n46192 , n22315 , n36813 );
and ( n46193 , n22326 , n37013 );
or ( n46194 , n36824 , n46118 );
or ( n46195 , n22334 , n36830 );
or ( n46196 , n36822 , n22336 );
nand ( n46197 , n46194 , n46195 , n46196 );
nor ( n46198 , n46193 , n46197 );
nand ( n46199 , n46192 , n46198 );
buf ( n46200 , n46199 );
buf ( n46201 , n379893 );
buf ( n46202 , n382069 );
buf ( n46203 , n22009 );
buf ( n46204 , n19653 );
not ( n46205 , n44039 );
or ( n46206 , n31053 , n46205 );
not ( n46207 , n31073 );
not ( n46208 , n31081 );
not ( n46209 , n46208 );
or ( n46210 , n46207 , n46209 );
nand ( n46211 , n46210 , n31091 );
and ( n46212 , n46211 , RI15b612f0_1181);
and ( n46213 , n383945 , RI15b58998_888);
and ( n46214 , n383949 , RI15b5a798_952);
nor ( n46215 , n46213 , n46214 );
and ( n46216 , n383955 , RI15b5af18_968);
and ( n46217 , n383960 , RI15b5ab58_960);
nor ( n46218 , n46216 , n46217 );
and ( n46219 , n383965 , RI15b5b2d8_976);
and ( n46220 , n383970 , RI15b5a018_936);
and ( n46221 , n383972 , RI15b5a3d8_944);
nor ( n46222 , n46220 , n46221 );
and ( n46223 , n383975 , RI15b59898_920);
and ( n46224 , n383977 , RI15b59c58_928);
nor ( n46225 , n46223 , n46224 );
and ( n46226 , n383982 , RI15b5be18_1000);
and ( n46227 , n383984 , RI15b5ba58_992);
nor ( n46228 , n46226 , n46227 );
and ( n46229 , n383987 , RI15b5c1d8_1008);
and ( n46230 , n383989 , RI15b5b698_984);
nor ( n46231 , n46229 , n46230 );
nand ( n46232 , n46222 , n46225 , n46228 , n46231 );
and ( n46233 , n383967 , n46232 );
and ( n46234 , n383994 , RI15b58d58_896);
nor ( n46235 , n46219 , n46233 , n46234 );
and ( n46236 , n383997 , RI15b59118_904);
and ( n46237 , n383999 , RI15b594d8_912);
nor ( n46238 , n46236 , n46237 );
nand ( n46239 , n46215 , n46218 , n46235 , n46238 );
and ( n46240 , n46239 , n31125 );
or ( n46241 , n31073 , n383563 , RI15b612f0_1181);
or ( n46242 , n383570 , RI15b61278_1180);
nand ( n46243 , n46241 , n46242 );
and ( n46244 , n40636 , n46243 );
nor ( n46245 , n46212 , n46240 , n46244 );
nand ( n46246 , n46206 , n44036 , n46245 );
buf ( n46247 , n46246 );
buf ( n46248 , n381707 );
or ( n46249 , n386705 , n31151 );
and ( n46250 , n386716 , n31164 );
or ( n46251 , n31175 , n17838 );
or ( n46252 , n45435 , n31182 );
or ( n46253 , n31173 , n386738 );
nand ( n46254 , n46251 , n46252 , n46253 );
nor ( n46255 , n46250 , n46254 );
nand ( n46256 , n46249 , n46255 );
buf ( n46257 , n46256 );
or ( n46258 , n22102 , n35957 );
and ( n46259 , n22203 , n36986 );
or ( n46260 , n35967 , n20287 );
or ( n46261 , n22293 , n35973 );
or ( n46262 , n35965 , n22299 );
nand ( n46263 , n46260 , n46261 , n46262 );
nor ( n46264 , n46259 , n46263 );
nand ( n46265 , n46258 , n46264 );
buf ( n46266 , n46265 );
buf ( n46267 , n384996 );
buf ( n46268 , n379895 );
buf ( n46269 , n381707 );
buf ( n46270 , n22009 );
or ( n46271 , n22315 , n35930 );
and ( n46272 , n22326 , n35935 );
not ( n46273 , RI15b40f50_81);
or ( n46274 , n35946 , n46273 );
or ( n46275 , n22334 , n35950 );
or ( n46276 , n35944 , n22336 );
nand ( n46277 , n46274 , n46275 , n46276 );
nor ( n46278 , n46272 , n46277 );
nand ( n46279 , n46271 , n46278 );
buf ( n46280 , n46279 );
buf ( n46281 , n384203 );
buf ( n46282 , n36488 );
buf ( n46283 , n34230 );
nor ( n46284 , n46282 , n46283 );
nand ( n46285 , n46284 , n379785 );
not ( n46286 , n46285 );
not ( n46287 , n36495 );
not ( n46288 , n46287 );
or ( n46289 , n46286 , n46288 );
buf ( n46290 , n34220 );
buf ( n46291 , n46290 );
nand ( n46292 , n46289 , n46291 );
nor ( n46293 , n46284 , n46290 );
nand ( n46294 , n36580 , n46293 );
buf ( n46295 , n34544 );
not ( n46296 , n46295 );
not ( n46297 , n34557 );
and ( n46298 , n46296 , n46297 );
not ( n46299 , n46296 );
and ( n46300 , n46299 , n34557 );
nor ( n46301 , n46298 , n46300 );
buf ( n46302 , n36512 );
and ( n46303 , n46301 , n46302 );
not ( n46304 , RI15b5e2a8_1078);
not ( n46305 , n34651 );
or ( n46306 , n46304 , n46305 );
or ( n46307 , n36518 , n379708 );
nand ( n46308 , n46306 , n46307 );
nor ( n46309 , n46303 , n46308 );
nand ( n46310 , n46292 , n46294 , n46309 );
buf ( n46311 , n46310 );
not ( n46312 , n36611 );
not ( n46313 , n36613 );
or ( n46314 , n46312 , n46313 );
or ( n46315 , n36613 , n36611 );
nand ( n46316 , n46314 , n46315 );
and ( n46317 , n46316 , n42541 );
nor ( n46318 , n21750 , n379309 );
nor ( n46319 , n46317 , n46318 );
not ( n46320 , n36649 );
and ( n46321 , n46320 , n36652 );
not ( n46322 , n46320 );
and ( n46323 , n46322 , n36653 );
nor ( n46324 , n46321 , n46323 );
nand ( n46325 , n46324 , n36457 );
nor ( n46326 , n36466 , n36673 );
not ( n46327 , n46326 );
nand ( n46328 , n46327 , n36674 );
nand ( n46329 , n46328 , n33644 );
and ( n46330 , n46319 , n46325 , n46329 );
and ( n46331 , n385164 , RI15b50bf8_620);
or ( n46332 , n44423 , n36673 );
or ( n46333 , n36652 , n385170 );
or ( n46334 , n36611 , n385178 );
nand ( n46335 , n46332 , n46333 , n46334 );
nor ( n46336 , n46331 , n46335 );
nand ( n46337 , n46330 , n46336 );
buf ( n46338 , n46337 );
buf ( n46339 , n20665 );
buf ( n46340 , n21611 );
and ( n46341 , n46340 , n34907 );
not ( n46342 , n46340 );
and ( n46343 , n46342 , n34906 );
nor ( n46344 , n46341 , n46343 );
and ( n46345 , n46344 , n21615 );
nor ( n46346 , n46344 , n21615 );
nor ( n46347 , n46345 , n46346 );
or ( n46348 , n21743 , n46347 );
not ( n46349 , n21022 );
not ( n46350 , n46349 );
not ( n46351 , n34903 );
or ( n46352 , n46350 , n46351 );
or ( n46353 , n34905 , n46349 );
nand ( n46354 , n46352 , n46353 );
not ( n46355 , n46354 );
not ( n46356 , n45501 );
or ( n46357 , n46355 , n46356 );
or ( n46358 , n45501 , n46354 );
nand ( n46359 , n46357 , n46358 );
and ( n46360 , n21353 , n46359 );
not ( n46361 , n21387 );
not ( n46362 , n46361 );
not ( n46363 , n21414 );
not ( n46364 , n35712 );
or ( n46365 , n46363 , n46364 );
nand ( n46366 , n46365 , n35692 );
and ( n46367 , n46366 , n34904 );
and ( n46368 , n21415 , n34903 );
nor ( n46369 , n46367 , n46368 );
not ( n46370 , n46369 );
or ( n46371 , n46362 , n46370 );
or ( n46372 , n46369 , n46361 );
nand ( n46373 , n46371 , n46372 );
and ( n46374 , n46373 , n21558 );
and ( n46375 , n21751 , RI15b57750_849);
nor ( n46376 , n46360 , n46374 , n46375 );
nand ( n46377 , n46348 , n46376 );
not ( n46378 , n46377 );
and ( n46379 , n21788 , RI15b56850_817);
and ( n46380 , n39103 , n17573 );
or ( n46381 , n379901 , RI15b56850_817);
not ( n46382 , RI15b56850_817);
or ( n46383 , n46382 , RI15b567d8_816);
nand ( n46384 , n46381 , n46383 );
and ( n46385 , n36237 , n46384 );
nor ( n46386 , n46379 , n46380 , n46385 );
nand ( n46387 , n46378 , n46386 );
buf ( n46388 , n46387 );
and ( n46389 , n380742 , n35796 );
and ( n46390 , n380741 , n35795 );
nor ( n46391 , n46389 , n46390 );
not ( n46392 , n19641 );
or ( n46393 , n46391 , n46392 );
and ( n46394 , n35684 , RI15b58650_881);
and ( n46395 , n380789 , n380754 );
and ( n46396 , n19630 , n380726 );
nor ( n46397 , n46394 , n46395 , n46396 );
nand ( n46398 , n46393 , n46397 );
buf ( n46399 , n46398 );
buf ( n46400 , n32672 );
and ( n46401 , n22646 , RI15b45870_237);
and ( n46402 , n22648 , RI15b51cd8_656);
nor ( n46403 , n46401 , n46402 );
not ( n46404 , n46403 );
buf ( n46405 , n46404 );
buf ( n46406 , n382069 );
buf ( n46407 , n380203 );
buf ( n46408 , n381081 );
not ( n46409 , n39633 );
xor ( n46410 , n46409 , n39642 );
or ( n46411 , n46410 , n31603 );
not ( n46412 , n379391 );
buf ( n46413 , n39667 );
not ( n46414 , n46413 );
or ( n46415 , n46412 , n46414 );
nand ( n46416 , n46415 , n31700 );
and ( n46417 , n46416 , n31695 );
or ( n46418 , n46413 , n39678 , n31695 );
and ( n46419 , n379394 , RI15b58290_873);
and ( n46420 , n39683 , RI15b52098_664);
nor ( n46421 , n46419 , n46420 );
nand ( n46422 , n46418 , n46421 );
nor ( n46423 , n46417 , n46422 );
nand ( n46424 , n46411 , n46423 );
buf ( n46425 , n46424 );
buf ( n46426 , n379893 );
and ( n46427 , n31792 , n384530 );
not ( n46428 , n384259 );
not ( n46429 , n37611 );
not ( n46430 , n46429 );
or ( n46431 , n46428 , n46430 );
or ( n46432 , n31771 , n384240 );
or ( n46433 , n32648 , n31779 );
nand ( n46434 , n46431 , n46432 , n46433 );
nor ( n46435 , n46427 , n46434 );
nand ( n46436 , n32660 , n46435 );
buf ( n46437 , n46436 );
buf ( n46438 , n22714 );
buf ( n46439 , n383174 );
buf ( n46440 , n382069 );
and ( n46441 , n22646 , RI15b45b40_243);
and ( n46442 , n22648 , RI15b51fa8_662);
nor ( n46443 , n46441 , n46442 );
not ( n46444 , n46443 );
buf ( n46445 , n46444 );
or ( n46446 , n380968 , n36200 );
and ( n46447 , n380986 , n36202 );
or ( n46448 , n36212 , n385452 );
or ( n46449 , n380994 , n36217 );
or ( n46450 , n36210 , n380996 );
nand ( n46451 , n46448 , n46449 , n46450 );
nor ( n46452 , n46447 , n46451 );
nand ( n46453 , n46446 , n46452 );
buf ( n46454 , n46453 );
buf ( n46455 , n379802 );
buf ( n46456 , n22402 );
and ( n46457 , n36999 , RI15b48138_324);
and ( n46458 , n37001 , RI15b44f88_218);
nor ( n46459 , n46457 , n46458 );
not ( n46460 , n46459 );
buf ( n46461 , n46460 );
buf ( n46462 , n381707 );
buf ( n46463 , n383613 );
buf ( n46464 , n386760 );
buf ( n46465 , n381004 );
not ( n46466 , n384705 );
not ( n46467 , n384122 );
or ( n46468 , n46466 , n46467 );
and ( n46469 , n384164 , n384739 );
or ( n46470 , n384749 , n20888 );
not ( n46471 , n384186 );
or ( n46472 , n46471 , n384757 );
or ( n46473 , n384747 , n384193 );
nand ( n46474 , n46470 , n46472 , n46473 );
nor ( n46475 , n46469 , n46474 );
nand ( n46476 , n46468 , n46475 );
buf ( n46477 , n46476 );
buf ( n46478 , n18226 );
nand ( n46479 , n384907 , n384825 );
buf ( n46480 , n41682 );
nand ( n46481 , n44037 , n46480 );
nand ( n46482 , n384918 , RI15b5f400_1115);
not ( n46483 , n383530 );
or ( n46484 , n44042 , n46483 );
nand ( n46485 , n46484 , n44044 );
not ( n46486 , n383538 );
and ( n46487 , n46485 , n46486 );
and ( n46488 , n383538 , n46483 );
and ( n46489 , n384934 , n46488 );
nor ( n46490 , n46487 , n46489 );
nand ( n46491 , n46479 , n46481 , n46482 , n46490 );
buf ( n46492 , n46491 );
buf ( n46493 , n380865 );
not ( n46494 , RI15b472b0_293);
not ( n46495 , n385213 );
or ( n46496 , n46494 , n46495 );
and ( n46497 , n385221 , RI15b48840_339);
and ( n46498 , n20631 , RI15b46b30_277);
nor ( n46499 , n46497 , n46498 );
nand ( n46500 , n46496 , n46499 );
buf ( n46501 , n46500 );
buf ( n46502 , n381021 );
buf ( n46503 , n32271 );
buf ( n46504 , n17499 );
buf ( n46505 , n379847 );
buf ( n46506 , n382049 );
buf ( n46507 , n22005 );
not ( n46508 , n34931 );
nor ( n46509 , n44769 , n44773 );
buf ( n46510 , n46509 );
not ( n46511 , n46510 );
or ( n46512 , n46508 , n46511 );
not ( n46513 , n35114 );
nand ( n46514 , n46512 , n46513 );
not ( n46515 , n35043 );
nand ( n46516 , n46514 , n46515 );
not ( n46517 , n46510 );
and ( n46518 , n46517 , n35118 , n35043 );
and ( n46519 , n385213 , RI15b47c10_313);
and ( n46520 , n20631 , RI15b46608_266);
nor ( n46521 , n46519 , n46520 );
not ( n46522 , n46521 );
nor ( n46523 , n46518 , n46522 );
nand ( n46524 , n46516 , n46523 );
buf ( n46525 , n46524 );
buf ( n46526 , n20663 );
buf ( n46527 , n22716 );
buf ( n46528 , n19651 );
or ( n46529 , n22775 , RI15b62bc8_1234);
or ( n46530 , n19608 , n19645 );
nand ( n46531 , n46530 , RI15b62bc8_1234);
or ( n46532 , RI15b5c3b8_1012 , RI15b5c430_1013);
nand ( n46533 , n46532 , n41363 );
and ( n46534 , n18631 , n46533 );
not ( n46535 , n19424 );
nor ( n46536 , n46534 , n46535 );
not ( n46537 , n42015 );
and ( n46538 , n46536 , n46537 );
not ( n46539 , n46536 );
and ( n46540 , n46539 , n42015 );
nor ( n46541 , n46538 , n46540 );
and ( n46542 , n19281 , n46541 );
and ( n46543 , n19513 , RI15b63ac8_1266);
not ( n46544 , n42011 );
not ( n46545 , n46536 );
or ( n46546 , n46544 , n46545 );
or ( n46547 , n46536 , n42011 );
nand ( n46548 , n46546 , n46547 );
and ( n46549 , n19500 , n46548 );
nor ( n46550 , n46542 , n46543 , n46549 );
nand ( n46551 , n46529 , n46531 , n46550 );
buf ( n46552 , n46551 );
buf ( n46553 , n381707 );
buf ( n46554 , n380942 );
nor ( n46555 , n36844 , n384177 );
buf ( n46556 , n46555 );
not ( n46557 , RI15b4a4d8_400);
not ( n46558 , n30908 );
or ( n46559 , n46557 , n46558 );
not ( n46560 , n19742 );
and ( n46561 , n46560 , n19746 );
not ( n46562 , n46560 );
and ( n46563 , n46562 , RI15b4a4d8_400);
nor ( n46564 , n46561 , n46563 );
and ( n46565 , n20637 , n46564 );
not ( n46566 , n386319 );
not ( n46567 , n42836 );
or ( n46568 , n46566 , n46567 );
not ( n46569 , n42835 );
nor ( n46570 , n46569 , n40186 );
or ( n46571 , n46570 , n42832 );
nand ( n46572 , n46571 , n386344 );
nand ( n46573 , n46568 , n46572 );
not ( n46574 , n35594 );
and ( n46575 , n46573 , n46574 );
not ( n46576 , n46573 );
and ( n46577 , n46576 , n35594 );
nor ( n46578 , n46575 , n46577 );
or ( n46579 , n46578 , n386499 );
xor ( n46580 , n385440 , n385493 );
xor ( n46581 , n46580 , n385763 );
and ( n46582 , n386014 , n46581 );
not ( n46583 , n35593 );
and ( n46584 , n46583 , n386128 );
and ( n46585 , n35593 , n386074 );
nor ( n46586 , n46584 , n46585 );
not ( n46587 , n46586 );
not ( n46588 , n42812 );
or ( n46589 , n46587 , n46588 );
or ( n46590 , n42812 , n46586 );
nand ( n46591 , n46589 , n46590 );
and ( n46592 , n46591 , n386258 );
and ( n46593 , n22394 , RI15b4b3d8_432);
nor ( n46594 , n46582 , n46592 , n46593 );
nand ( n46595 , n46579 , n46594 );
nor ( n46596 , n22216 , n19748 );
nor ( n46597 , n46565 , n46595 , n46596 );
nand ( n46598 , n46559 , n46597 );
buf ( n46599 , n46598 );
buf ( n46600 , n22740 );
buf ( n46601 , n19655 );
not ( n46602 , RI15b533d0_705);
not ( n46603 , n32244 );
or ( n46604 , n46602 , n46603 );
and ( n46605 , n32247 , RI15b649c8_1298);
and ( n46606 , n32249 , RI15b5f838_1124);
nor ( n46607 , n46605 , n46606 );
nand ( n46608 , n46604 , n46607 );
buf ( n46609 , n46608 );
buf ( n46610 , n32672 );
buf ( n46611 , n382067 );
buf ( n46612 , n383498 );
buf ( n46613 , n384218 );
not ( n46614 , n379825 );
not ( n46615 , n46510 );
or ( n46616 , n46614 , n46615 );
nand ( n46617 , n46616 , n41032 );
nand ( n46618 , n46617 , n46515 );
and ( n46619 , n46517 , n41651 , n35043 );
not ( n46620 , RI15b46608_266);
not ( n46621 , n379832 );
or ( n46622 , n46620 , n46621 );
and ( n46623 , n38858 , n35461 );
and ( n46624 , n35459 , n382026 );
nor ( n46625 , n46623 , n46624 );
nand ( n46626 , n46622 , n46625 );
nor ( n46627 , n46619 , n46626 );
nand ( n46628 , n46618 , n46627 );
buf ( n46629 , n46628 );
buf ( n46630 , n382049 );
buf ( n46631 , n387159 );
buf ( n46632 , n22655 );
not ( n46633 , n385947 );
and ( n46634 , n46633 , n385960 );
not ( n46635 , n46633 );
and ( n46636 , n46635 , n385959 );
nor ( n46637 , n46634 , n46636 );
not ( n46638 , n386019 );
nor ( n46639 , n46637 , n46638 );
buf ( n46640 , n386235 );
not ( n46641 , n46640 );
not ( n46642 , n386045 );
and ( n46643 , n46641 , n46642 );
and ( n46644 , n46640 , n386045 );
nor ( n46645 , n46643 , n46644 );
not ( n46646 , n39973 );
or ( n46647 , n46645 , n46646 );
not ( n46648 , n386290 );
not ( n46649 , n386487 );
not ( n46650 , n46649 );
or ( n46651 , n46648 , n46650 );
nand ( n46652 , n46651 , n40755 );
and ( n46653 , n46652 , n386500 );
nor ( n46654 , n34784 , n382143 );
nor ( n46655 , n46653 , n46654 );
nand ( n46656 , n46647 , n46655 );
nor ( n46657 , n46639 , n46656 );
and ( n46658 , n40389 , n386290 );
or ( n46659 , n386541 , n386287 );
or ( n46660 , n385959 , n386550 );
or ( n46661 , n386557 , n386045 );
nand ( n46662 , n46659 , n46660 , n46661 );
nor ( n46663 , n46658 , n46662 );
nand ( n46664 , n46657 , n46663 );
buf ( n46665 , n46664 );
buf ( n46666 , n380865 );
buf ( n46667 , n387159 );
buf ( n46668 , n381872 );
buf ( n46669 , n33250 );
and ( n46670 , n33294 , n21771 );
not ( n46671 , n17514 );
not ( n46672 , n37997 );
or ( n46673 , n46671 , n46672 );
nand ( n46674 , n46673 , n21790 );
and ( n46675 , n46674 , RI15b571b0_837);
nor ( n46676 , n17514 , RI15b571b0_837);
and ( n46677 , n21795 , n46676 );
nor ( n46678 , n46670 , n46675 , n46677 );
nand ( n46679 , n43272 , n46678 );
buf ( n46680 , n46679 );
buf ( n46681 , n19655 );
buf ( n46682 , n382065 );
buf ( n46683 , n21893 );
nor ( n46684 , n46683 , n33323 );
and ( n46685 , n379855 , n46684 );
and ( n46686 , n40407 , RI15b57cf0_861);
not ( n46687 , n21970 );
not ( n46688 , n46687 );
not ( n46689 , n21949 );
or ( n46690 , n46688 , n46689 );
nand ( n46691 , n46690 , n21979 );
and ( n46692 , n46691 , RI15b55ef0_797);
or ( n46693 , n21982 , n46687 , RI15b55ef0_797);
and ( n46694 , n40405 , n21941 , RI15b57c78_860);
and ( n46695 , n21940 , RI15b57cf0_861);
nor ( n46696 , n46694 , n46695 );
or ( n46697 , n21922 , n46696 );
nand ( n46698 , n46693 , n46697 );
nor ( n46699 , n46686 , n46692 , n46698 );
or ( n46700 , n46699 , n18078 );
and ( n46701 , n18177 , RI15b57cf0_861);
and ( n46702 , n18219 , RI15b56df0_829);
nor ( n46703 , n46701 , n46702 , n21751 );
nand ( n46704 , n46700 , n46703 );
nor ( n46705 , n46685 , n46704 );
nand ( n46706 , n46683 , n17507 );
not ( n46707 , n46706 );
not ( n46708 , n17565 );
or ( n46709 , n46707 , n46708 );
nand ( n46710 , n46709 , n33323 );
nand ( n46711 , n46705 , n46710 );
buf ( n46712 , n46711 );
buf ( n46713 , n379893 );
buf ( n46714 , n32676 );
buf ( n46715 , n384996 );
buf ( n46716 , n19653 );
buf ( n46717 , n382073 );
nand ( n46718 , n32020 , n32037 );
nor ( n46719 , n46718 , n382079 );
buf ( n46720 , n382474 );
not ( n46721 , n46720 );
or ( n46722 , n46719 , n46721 );
nand ( n46723 , n46722 , n32898 );
nor ( n46724 , n32035 , n32898 );
and ( n46725 , n46718 , n46724 );
not ( n46726 , n382337 );
and ( n46727 , n382338 , RI15b4b888_442);
nor ( n46728 , n46727 , n382348 );
and ( n46729 , n46726 , n46728 );
not ( n46730 , n46726 );
and ( n46731 , n46730 , n382343 );
or ( n46732 , n46729 , n46731 );
or ( n46733 , n382513 , n46732 );
and ( n46734 , n382523 , RI15b4b888_442);
and ( n46735 , n382529 , RI15b45690_233);
nor ( n46736 , n46734 , n46735 );
nand ( n46737 , n46733 , n46736 );
nor ( n46738 , n46725 , n46737 );
nand ( n46739 , n46723 , n46738 );
buf ( n46740 , n46739 );
buf ( n46741 , n380942 );
not ( n46742 , RI15b55608_778);
not ( n46743 , n382680 );
or ( n46744 , n46742 , n46743 );
and ( n46745 , n382685 , n382681 );
not ( n46746 , n382786 );
not ( n46747 , n382831 );
and ( n46748 , n46746 , n46747 );
and ( n46749 , n382786 , n382831 );
nor ( n46750 , n46748 , n46749 );
or ( n46751 , n382886 , n46750 );
or ( n46752 , n383744 , n382691 );
nor ( n46753 , n381400 , n41885 );
not ( n46754 , n46753 );
nand ( n46755 , n46751 , n46752 , n46754 );
nor ( n46756 , n46745 , n46755 );
nand ( n46757 , n46744 , n46756 );
buf ( n46758 , n46757 );
buf ( n46759 , n22007 );
not ( n46760 , n382898 );
not ( n46761 , n33400 );
or ( n46762 , n46760 , n46761 );
and ( n46763 , n33415 , n382934 );
not ( n46764 , RI15b59898_920);
or ( n46765 , n382949 , n46764 );
or ( n46766 , n36293 , n382965 );
or ( n46767 , n382947 , n33443 );
nand ( n46768 , n46765 , n46766 , n46767 );
nor ( n46769 , n46763 , n46768 );
nand ( n46770 , n46762 , n46769 );
buf ( n46771 , n46770 );
buf ( n46772 , n22655 );
not ( n46773 , RI15b53790_713);
not ( n46774 , n32244 );
or ( n46775 , n46773 , n46774 );
and ( n46776 , n32247 , RI15b64d88_1306);
and ( n46777 , n32249 , RI15b5fbf8_1132);
nor ( n46778 , n46776 , n46777 );
nand ( n46779 , n46775 , n46778 );
buf ( n46780 , n46779 );
or ( n46781 , n37137 , n37107 );
not ( n46782 , n37356 );
not ( n46783 , n46782 );
not ( n46784 , n37386 );
and ( n46785 , n46783 , n46784 );
and ( n46786 , n46782 , n37386 );
nor ( n46787 , n46785 , n46786 );
not ( n46788 , n46787 );
not ( n46789 , n381062 );
and ( n46790 , n46788 , n46789 );
and ( n46791 , n37426 , n37107 );
nor ( n46792 , n46790 , n46791 );
nand ( n46793 , n46781 , n46792 );
buf ( n46794 , n46793 );
buf ( n46795 , n384700 );
buf ( n46796 , n35651 );
buf ( n46797 , n20663 );
buf ( n46798 , n22716 );
buf ( n46799 , n384700 );
buf ( n46800 , n387159 );
buf ( n46801 , n35651 );
not ( n46802 , RI15b54078_732);
not ( n46803 , n32244 );
or ( n46804 , n46802 , n46803 );
and ( n46805 , n32247 , RI15b65670_1325);
and ( n46806 , n32249 , RI15b604e0_1151);
nor ( n46807 , n46805 , n46806 );
nand ( n46808 , n46804 , n46807 );
buf ( n46809 , n46808 );
buf ( n46810 , n22479 );
and ( n46811 , n32747 , RI15b42918_136);
not ( n46812 , n32749 );
and ( n46813 , n32753 , RI15b41658_96);
and ( n46814 , n32755 , RI15b41a18_104);
nor ( n46815 , n46813 , n46814 );
and ( n46816 , n32759 , RI15b40ed8_80);
and ( n46817 , n32762 , RI15b41298_88);
nor ( n46818 , n46816 , n46817 );
and ( n46819 , n32766 , RI15b43458_160);
and ( n46820 , n32768 , RI15b43098_152);
nor ( n46821 , n46819 , n46820 );
and ( n46822 , n32771 , RI15b43818_168);
and ( n46823 , n32773 , RI15b42cd8_144);
nor ( n46824 , n46822 , n46823 );
nand ( n46825 , n46815 , n46818 , n46821 , n46824 );
and ( n46826 , n46812 , n46825 );
and ( n46827 , n32781 , RI15b40398_56);
nor ( n46828 , n46811 , n46826 , n46827 );
and ( n46829 , n32785 , RI15b42558_128);
and ( n46830 , n32787 , RI15b42198_120);
nor ( n46831 , n46829 , n46830 );
and ( n46832 , n32792 , RI15b3ffd8_48);
and ( n46833 , n32794 , RI15b41dd8_112);
nor ( n46834 , n46832 , n46833 );
and ( n46835 , n32797 , RI15b40758_64);
and ( n46836 , n32800 , RI15b40b18_72);
nor ( n46837 , n46835 , n46836 );
nand ( n46838 , n46828 , n46831 , n46834 , n46837 );
not ( n46839 , n46838 );
or ( n46840 , n46839 , n36051 );
and ( n46841 , n381055 , RI15b49830_373);
not ( n46842 , RI15b49830_373);
not ( n46843 , n32820 );
or ( n46844 , n46842 , n46843 );
or ( n46845 , n32820 , RI15b49830_373);
nand ( n46846 , n46844 , n46845 );
and ( n46847 , n36064 , n46846 );
nor ( n46848 , n46841 , n46847 );
nand ( n46849 , n46840 , n46848 );
buf ( n46850 , n46849 );
or ( n46851 , n383180 , n35144 );
not ( n46852 , n35160 );
and ( n46853 , n46852 , RI15b5b0f8_972);
or ( n46854 , n383184 , n35149 );
or ( n46855 , n32696 , n35166 );
or ( n46856 , n35158 , n383192 );
nand ( n46857 , n46854 , n46855 , n46856 );
nor ( n46858 , n46853 , n46857 );
nand ( n46859 , n46851 , n46858 );
buf ( n46860 , n46859 );
buf ( n46861 , n380203 );
not ( n46862 , RI15b53da8_726);
not ( n46863 , n383170 );
or ( n46864 , n46862 , n46863 );
or ( n46865 , n33347 , n383152 );
nand ( n46866 , n46865 , n383157 );
and ( n46867 , n46866 , n33358 );
not ( n46868 , RI15b527a0_679);
not ( n46869 , n383147 );
or ( n46870 , n46868 , n46869 );
or ( n46871 , n33348 , n383144 );
nand ( n46872 , n46870 , n46871 );
nor ( n46873 , n46867 , n46872 );
nand ( n46874 , n46864 , n46873 );
buf ( n46875 , n46874 );
buf ( n46876 , n382069 );
buf ( n46877 , n385112 );
buf ( n46878 , n381021 );
not ( n46879 , RI15b46e78_284);
not ( n46880 , n379832 );
or ( n46881 , n46879 , n46880 );
and ( n46882 , n379825 , RI15b48b88_346);
nor ( n46883 , n46882 , n44492 );
nand ( n46884 , n46881 , n46883 );
buf ( n46885 , n46884 );
buf ( n46886 , n22005 );
buf ( n46887 , n32255 );
buf ( n46888 , n383345 );
buf ( n46889 , n381566 );
buf ( n46890 , n380203 );
buf ( n46891 , n382069 );
not ( n46892 , n36395 );
not ( n46893 , n380703 );
or ( n46894 , n46892 , n46893 );
and ( n46895 , n380719 , n36401 );
or ( n46896 , n36410 , n19029 );
or ( n46897 , n380782 , n36416 );
or ( n46898 , n36408 , n380790 );
nand ( n46899 , n46896 , n46897 , n46898 );
nor ( n46900 , n46895 , n46899 );
nand ( n46901 , n46894 , n46900 );
buf ( n46902 , n46901 );
not ( n46903 , RI15b55860_783);
not ( n46904 , n380000 );
or ( n46905 , n46903 , n46904 );
not ( n46906 , n379948 );
not ( n46907 , n385099 );
and ( n46908 , n46906 , n46907 );
and ( n46909 , n380010 , RI15b4c3c8_466);
nor ( n46910 , n46908 , n46909 );
nand ( n46911 , n46905 , n46910 );
buf ( n46912 , n46911 );
buf ( n46913 , n33382 );
or ( n46914 , n22102 , n37495 );
and ( n46915 , n22203 , n37498 );
or ( n46916 , n37507 , n385527 );
or ( n46917 , n22293 , n37512 );
or ( n46918 , n37505 , n22299 );
nand ( n46919 , n46916 , n46917 , n46918 );
nor ( n46920 , n46915 , n46919 );
nand ( n46921 , n46914 , n46920 );
buf ( n46922 , n46921 );
buf ( n46923 , n22343 );
buf ( n46924 , n380203 );
buf ( n46925 , n381021 );
buf ( n46926 , n379844 );
buf ( n46927 , n22788 );
buf ( n46928 , n32160 );
buf ( n46929 , n379847 );
not ( n46930 , RI15b475f8_300);
not ( n46931 , n385213 );
or ( n46932 , n46930 , n46931 );
and ( n46933 , n385221 , RI15b48b88_346);
and ( n46934 , n20631 , RI15b46e78_284);
nor ( n46935 , n46933 , n46934 );
nand ( n46936 , n46932 , n46935 );
buf ( n46937 , n46936 );
buf ( n46938 , n32255 );
buf ( n46939 , n22788 );
or ( n46940 , n36266 , n39875 );
nand ( n46941 , n36269 , RI15b54b40_755);
and ( n46942 , n39877 , n46941 );
nand ( n46943 , n381486 , RI15b52e30_693);
nand ( n46944 , n46940 , n46942 , n46943 );
buf ( n46945 , n46944 );
or ( n46946 , n386588 , n36275 );
and ( n46947 , n386600 , n36282 );
not ( n46948 , RI15b5c070_1005);
or ( n46949 , n36291 , n46948 );
or ( n46950 , n386618 , n36296 );
or ( n46951 , n36289 , n386627 );
nand ( n46952 , n46949 , n46950 , n46951 );
nor ( n46953 , n46947 , n46952 );
nand ( n46954 , n46946 , n46953 );
buf ( n46955 , n46954 );
buf ( n46956 , n380940 );
buf ( n46957 , n22653 );
buf ( n46958 , n22408 );
buf ( n46959 , n385197 );
not ( n46960 , n38373 );
not ( n46961 , n46960 );
not ( n46962 , n39319 );
or ( n46963 , n46961 , n46962 );
and ( n46964 , n33196 , n38375 );
or ( n46965 , n38385 , n20119 );
or ( n46966 , n22241 , n38389 );
or ( n46967 , n38383 , n33201 );
nand ( n46968 , n46965 , n46966 , n46967 );
nor ( n46969 , n46964 , n46968 );
nand ( n46970 , n46963 , n46969 );
buf ( n46971 , n46970 );
not ( n46972 , RI15b47058_288);
not ( n46973 , n385213 );
or ( n46974 , n46972 , n46973 );
and ( n46975 , n385221 , RI15b485e8_334);
and ( n46976 , n20631 , RI15b468d8_272);
nor ( n46977 , n46975 , n46976 );
nand ( n46978 , n46974 , n46977 );
buf ( n46979 , n46978 );
buf ( n46980 , n32160 );
buf ( n46981 , n22005 );
buf ( n46982 , n379847 );
buf ( n46983 , n386762 );
buf ( n46984 , n382065 );
buf ( n46985 , n381081 );
buf ( n46986 , n382071 );
not ( n46987 , n32869 );
and ( n46988 , n32941 , n46987 );
nor ( n46989 , n44169 , n46988 );
or ( n46990 , n46989 , n32874 );
not ( n46991 , n44167 );
nor ( n46992 , n44171 , n382079 );
nand ( n46993 , n46991 , n46992 );
buf ( n46994 , n32868 );
or ( n46995 , n46993 , n46994 );
not ( n46996 , n32024 );
nand ( n46997 , n46995 , n46996 );
nand ( n46998 , n46997 , n32874 );
not ( n46999 , n43107 );
xor ( n47000 , n382421 , n382430 );
and ( n47001 , n46999 , n47000 );
and ( n47002 , n382523 , RI15b4bc48_450);
and ( n47003 , n43116 , RI15b45a50_241);
nor ( n47004 , n47002 , n47003 );
not ( n47005 , n47004 );
nor ( n47006 , n47001 , n47005 );
nand ( n47007 , n46990 , n46998 , n47006 );
buf ( n47008 , n47007 );
buf ( n47009 , n382073 );
buf ( n47010 , n22404 );
buf ( n47011 , n383174 );
buf ( n47012 , n386563 );
buf ( n47013 , n43349 );
not ( n47014 , RI15b47418_296);
not ( n47015 , n385213 );
or ( n47016 , n47014 , n47015 );
and ( n47017 , n385221 , RI15b489a8_342);
and ( n47018 , n20631 , RI15b46c98_280);
nor ( n47019 , n47017 , n47018 );
nand ( n47020 , n47016 , n47019 );
buf ( n47021 , n47020 );
buf ( n47022 , n384700 );
nor ( n47023 , n45296 , n45298 );
not ( n47024 , n47023 );
buf ( n47025 , n31458 );
not ( n47026 , n47025 );
and ( n47027 , n47024 , n47026 );
not ( n47028 , n47024 );
not ( n47029 , n47026 );
and ( n47030 , n47028 , n47029 );
nor ( n47031 , n47027 , n47030 );
nand ( n47032 , n47031 , n45735 );
or ( n47033 , n31707 , n379230 );
nand ( n47034 , n47033 , n42053 );
not ( n47035 , n31655 );
and ( n47036 , n47034 , n47035 );
and ( n47037 , n379394 , RI15b57fc0_867);
buf ( n47038 , n379398 );
and ( n47039 , n47038 , RI15b51dc8_658);
nor ( n47040 , n47037 , n47039 );
not ( n47041 , n47040 );
nor ( n47042 , n47036 , n47041 );
not ( n47043 , n379230 );
not ( n47044 , n42050 );
or ( n47045 , n47043 , n47044 );
nand ( n47046 , n47045 , n31700 );
nand ( n47047 , n47046 , n31655 );
nand ( n47048 , n47032 , n47042 , n47047 );
buf ( n47049 , n47048 );
buf ( n47050 , n384203 );
and ( n47051 , n31792 , n31944 );
and ( n47052 , n31770 , RI15b5d0d8_1040);
and ( n47053 , n42116 , n31903 );
and ( n47054 , n31858 , n31778 );
nor ( n47055 , n47052 , n47053 , n47054 );
not ( n47056 , n47055 );
nor ( n47057 , n47051 , n47056 );
nand ( n47058 , n39049 , n47057 );
buf ( n47059 , n47058 );
not ( n47060 , n382976 );
not ( n47061 , n381507 );
or ( n47062 , n47060 , n47061 );
and ( n47063 , n381524 , n382983 );
or ( n47064 , n382995 , n18380 );
or ( n47065 , n32478 , n383001 );
or ( n47066 , n382993 , n381560 );
nand ( n47067 , n47064 , n47065 , n47066 );
nor ( n47068 , n47063 , n47067 );
nand ( n47069 , n47062 , n47068 );
buf ( n47070 , n47069 );
nand ( n47071 , n38895 , n383143 );
not ( n47072 , n383153 );
not ( n47073 , n38894 );
or ( n47074 , n47072 , n47073 );
nand ( n47075 , n47074 , n383157 );
nand ( n47076 , n47075 , n38902 );
nand ( n47077 , n383170 , RI15b53e98_728);
nand ( n47078 , n383147 , RI15b52890_681);
nand ( n47079 , n47071 , n47076 , n47077 , n47078 );
buf ( n47080 , n47079 );
buf ( n47081 , n380903 );
buf ( n47082 , n379844 );
buf ( n47083 , n22406 );
buf ( n47084 , n19651 );
buf ( n47085 , n382071 );
or ( n47086 , n31006 , n35472 );
and ( n47087 , n31016 , n35479 );
or ( n47088 , n35488 , n20966 );
or ( n47089 , n34893 , n35497 );
or ( n47090 , n35486 , n31024 );
nand ( n47091 , n47088 , n47089 , n47090 );
nor ( n47092 , n47087 , n47091 );
nand ( n47093 , n47086 , n47092 );
buf ( n47094 , n47093 );
or ( n47095 , n31053 , n381615 );
and ( n47096 , n36536 , RI15b60fa8_1174);
not ( n47097 , n33050 );
and ( n47098 , n36538 , n47097 );
not ( n47099 , RI15b60fa8_1174);
not ( n47100 , n31064 );
or ( n47101 , n47099 , n47100 );
or ( n47102 , n31064 , RI15b60fa8_1174);
nand ( n47103 , n47101 , n47102 );
and ( n47104 , n40636 , n47103 );
nor ( n47105 , n47096 , n47098 , n47104 );
nand ( n47106 , n47095 , n41172 , n47105 );
buf ( n47107 , n47106 );
buf ( n47108 , n22343 );
not ( n47109 , n35957 );
not ( n47110 , n47109 );
not ( n47111 , n32129 );
or ( n47112 , n47110 , n47111 );
and ( n47113 , n35968 , RI15b3ff60_47);
or ( n47114 , n32141 , n35959 );
or ( n47115 , n32148 , n35973 );
or ( n47116 , n35965 , n32150 );
nand ( n47117 , n47114 , n47115 , n47116 );
nor ( n47118 , n47113 , n47117 );
nand ( n47119 , n47112 , n47118 );
buf ( n47120 , n47119 );
buf ( n47121 , n20665 );
buf ( n47122 , n382067 );
buf ( n47123 , n22007 );
buf ( n47124 , n20665 );
or ( n47125 , n42942 , n35930 );
and ( n47126 , n384983 , n35935 );
not ( n47127 , RI15b410b8_84);
or ( n47128 , n35946 , n47127 );
or ( n47129 , n22022 , n35950 );
or ( n47130 , n35944 , n384988 );
nand ( n47131 , n47128 , n47129 , n47130 );
nor ( n47132 , n47126 , n47131 );
nand ( n47133 , n47125 , n47132 );
buf ( n47134 , n47133 );
or ( n47135 , n42942 , n38065 );
and ( n47136 , n384983 , n38067 );
or ( n47137 , n38077 , n20395 );
or ( n47138 , n22022 , n38081 );
or ( n47139 , n38075 , n384988 );
nand ( n47140 , n47137 , n47138 , n47139 );
nor ( n47141 , n47136 , n47140 );
nand ( n47142 , n47135 , n47141 );
buf ( n47143 , n47142 );
buf ( n47144 , n22009 );
buf ( n47145 , n22402 );
buf ( n47146 , n382071 );
buf ( n47147 , n43349 );
buf ( n47148 , n31979 );
buf ( n47149 , n19653 );
not ( n47150 , n46480 );
or ( n47151 , n31053 , n47150 );
and ( n47152 , n36536 , RI15b61110_1177);
and ( n47153 , n42378 , n39368 );
not ( n47154 , n41340 );
not ( n47155 , RI15b61110_1177);
not ( n47156 , n31069 );
or ( n47157 , n47155 , n47156 );
or ( n47158 , n31069 , RI15b61110_1177);
nand ( n47159 , n47157 , n47158 );
and ( n47160 , n47154 , n47159 );
nor ( n47161 , n47152 , n47153 , n47160 );
nand ( n47162 , n47151 , n46479 , n47161 );
buf ( n47163 , n47162 );
or ( n47164 , n36238 , n35481 );
or ( n47165 , n21164 , n35488 );
and ( n47166 , n35496 , n36256 );
and ( n47167 , n383803 , n35470 );
and ( n47168 , n36261 , n35493 );
nor ( n47169 , n47166 , n47167 , n47168 );
nand ( n47170 , n47164 , n47165 , n47169 );
buf ( n47171 , n47170 );
buf ( n47172 , n384996 );
buf ( n47173 , n30992 );
and ( n47174 , n22646 , RI15b455a0_231);
and ( n47175 , n22648 , RI15b51a08_650);
nor ( n47176 , n47174 , n47175 );
not ( n47177 , n47176 );
buf ( n47178 , n47177 );
buf ( n47179 , n379802 );
buf ( n47180 , n20665 );
or ( n47181 , n381907 , n36200 );
and ( n47182 , n42409 , RI15b41658_96);
or ( n47183 , n381917 , n36204 );
not ( n47184 , n36217 );
and ( n47185 , n47184 , n381923 );
and ( n47186 , n381926 , n36215 );
nor ( n47187 , n47185 , n47186 );
nand ( n47188 , n47183 , n47187 );
nor ( n47189 , n47182 , n47188 );
nand ( n47190 , n47181 , n47189 );
buf ( n47191 , n47190 );
buf ( n47192 , n383174 );
buf ( n47193 , n31979 );
or ( n47194 , n31091 , n32309 );
buf ( n47195 , n31121 );
not ( n47196 , n47195 );
and ( n47197 , n38654 , RI15b5b1e8_974);
and ( n47198 , n39717 , RI15b5ae28_966);
nor ( n47199 , n47197 , n47198 );
and ( n47200 , n39721 , RI15b5aa68_958);
and ( n47201 , n39724 , RI15b5a6a8_950);
nor ( n47202 , n47200 , n47201 );
and ( n47203 , n39728 , RI15b5a2e8_942);
and ( n47204 , n39731 , RI15b59f28_934);
nor ( n47205 , n47203 , n47204 );
and ( n47206 , n39735 , RI15b59b68_926);
and ( n47207 , n39738 , RI15b597a8_918);
nor ( n47208 , n47206 , n47207 );
nand ( n47209 , n47199 , n47202 , n47205 , n47208 );
and ( n47210 , n383968 , n47209 );
and ( n47211 , n39746 , RI15b58c68_894);
and ( n47212 , n39751 , RI15b5c0e8_1006);
nor ( n47213 , n47210 , n47211 , n47212 );
and ( n47214 , n39756 , RI15b5bd28_998);
and ( n47215 , n39759 , RI15b5b968_990);
nor ( n47216 , n47214 , n47215 );
and ( n47217 , n39763 , RI15b593e8_910);
and ( n47218 , n39765 , RI15b59028_902);
nor ( n47219 , n47217 , n47218 );
and ( n47220 , n39769 , RI15b588a8_886);
and ( n47221 , n39772 , RI15b5b5a8_982);
nor ( n47222 , n47220 , n47221 );
and ( n47223 , n47213 , n47216 , n47219 , n47222 );
or ( n47224 , n47196 , n47223 );
or ( n47225 , n31052 , n380622 );
and ( n47226 , n41416 , RI15b615c0_1187);
not ( n47227 , n41416 );
and ( n47228 , n47227 , n32309 );
nor ( n47229 , n47226 , n47228 );
or ( n47230 , n47229 , n43838 );
nand ( n47231 , n47225 , n47230 );
nor ( n47232 , n47231 , n40496 );
nand ( n47233 , n47194 , n47224 , n47232 );
buf ( n47234 , n47233 );
buf ( n47235 , n381006 );
buf ( n47236 , n380203 );
not ( n47237 , n41756 );
not ( n47238 , n384122 );
or ( n47239 , n47237 , n47238 );
and ( n47240 , n384164 , n41446 );
or ( n47241 , n41455 , n17900 );
or ( n47242 , n384187 , n41461 );
or ( n47243 , n41453 , n384193 );
nand ( n47244 , n47241 , n47242 , n47243 );
nor ( n47245 , n47240 , n47244 );
nand ( n47246 , n47239 , n47245 );
buf ( n47247 , n47246 );
buf ( n47248 , n22007 );
not ( n47249 , n36624 );
not ( n47250 , n36614 );
not ( n47251 , n47250 );
or ( n47252 , n47249 , n47251 );
or ( n47253 , n47250 , n36624 );
nand ( n47254 , n47252 , n47253 );
and ( n47255 , n47254 , n21564 );
nor ( n47256 , n21750 , n22622 );
nor ( n47257 , n47255 , n47256 );
and ( n47258 , n36654 , n36658 );
not ( n47259 , n36654 );
not ( n47260 , n36658 );
and ( n47261 , n47259 , n47260 );
nor ( n47262 , n47258 , n47261 );
not ( n47263 , n21359 );
nand ( n47264 , n47262 , n47263 );
not ( n47265 , n36674 );
nor ( n47266 , n47265 , n36677 );
not ( n47267 , n47266 );
not ( n47268 , n36679 );
nand ( n47269 , n47267 , n47268 );
nand ( n47270 , n47269 , n33644 );
and ( n47271 , n47257 , n47264 , n47270 );
and ( n47272 , n44703 , n42548 );
not ( n47273 , n384127 );
or ( n47274 , n17522 , n47273 );
nand ( n47275 , n47274 , n21790 );
and ( n47276 , n47275 , RI15b57408_842);
and ( n47277 , n17522 , n22556 );
and ( n47278 , n21795 , n47277 );
nor ( n47279 , n47272 , n47276 , n47278 );
nand ( n47280 , n47271 , n47279 );
buf ( n47281 , n47280 );
buf ( n47282 , n32676 );
buf ( n47283 , n382537 );
nor ( n47284 , n21854 , n44756 );
and ( n47285 , n379855 , n47284 );
buf ( n47286 , n21961 );
not ( n47287 , n47286 );
not ( n47288 , n21949 );
or ( n47289 , n47287 , n47288 );
nand ( n47290 , n47289 , n21979 );
and ( n47291 , n47290 , RI15b55c98_792);
and ( n47292 , n18150 , RI15b57a98_856);
or ( n47293 , n21982 , n47286 , RI15b55c98_792);
not ( n47294 , n21932 );
not ( n47295 , n47294 );
not ( n47296 , RI15b57a98_856);
and ( n47297 , n47295 , n47296 );
and ( n47298 , n47294 , RI15b57a98_856);
nor ( n47299 , n47297 , n47298 );
or ( n47300 , n21922 , n47299 );
nand ( n47301 , n47293 , n47300 );
nor ( n47302 , n47291 , n47292 , n47301 );
or ( n47303 , n47302 , n18078 );
and ( n47304 , n18177 , RI15b57a98_856);
and ( n47305 , n18219 , RI15b56b98_824);
nor ( n47306 , n47304 , n47305 , n21751 );
nand ( n47307 , n47303 , n47306 );
nor ( n47308 , n47285 , n47307 );
not ( n47309 , n17507 );
not ( n47310 , n21854 );
or ( n47311 , n47309 , n47310 );
nand ( n47312 , n47311 , n17565 );
nand ( n47313 , n47312 , n44756 );
nand ( n47314 , n47308 , n47313 );
buf ( n47315 , n47314 );
buf ( n47316 , n32271 );
buf ( n47317 , n384203 );
buf ( n47318 , n382052 );
buf ( n47319 , n22655 );
or ( n47320 , n22102 , n36121 );
and ( n47321 , n22203 , n36123 );
not ( n47322 , RI15b43908_170);
or ( n47323 , n36132 , n47322 );
or ( n47324 , n22293 , n36139 );
or ( n47325 , n36130 , n22299 );
nand ( n47326 , n47323 , n47324 , n47325 );
nor ( n47327 , n47321 , n47326 );
nand ( n47328 , n47320 , n47327 );
buf ( n47329 , n47328 );
buf ( n47330 , n381004 );
buf ( n47331 , n22343 );
buf ( n47332 , n379895 );
not ( n47333 , n22523 );
nor ( n47334 , n47333 , n22529 );
and ( n47335 , n21802 , n47334 );
not ( n47336 , RI15b56328_806);
not ( n47337 , n18086 );
not ( n47338 , n22588 );
not ( n47339 , n47338 );
or ( n47340 , n47337 , n47339 );
nand ( n47341 , n47340 , n18104 );
not ( n47342 , n47341 );
or ( n47343 , n47336 , n47342 );
not ( n47344 , RI15b56328_806);
nand ( n47345 , n18198 , n47344 );
nor ( n47346 , n47338 , n47345 );
not ( n47347 , n22619 );
and ( n47348 , n18188 , n47347 );
nor ( n47349 , n47348 , n18179 );
nor ( n47350 , n47349 , n22836 );
or ( n47351 , n18189 , n47347 , RI15b58128_870);
or ( n47352 , n18218 , n22525 );
nand ( n47353 , n47351 , n47352 );
nor ( n47354 , n47346 , n47350 , n47353 );
nand ( n47355 , n47343 , n47354 );
nor ( n47356 , n47335 , n47355 );
not ( n47357 , n17507 );
not ( n47358 , n47333 );
or ( n47359 , n47357 , n47358 );
nand ( n47360 , n47359 , n17565 );
nand ( n47361 , n47360 , n22529 );
nand ( n47362 , n47356 , n47361 );
buf ( n47363 , n47362 );
buf ( n47364 , n385122 );
not ( n47365 , n47364 );
nor ( n47366 , n47365 , n21710 );
not ( n47367 , n47366 );
not ( n47368 , n385125 );
nand ( n47369 , n47367 , n47368 );
and ( n47370 , n47369 , n43267 );
nor ( n47371 , n45250 , n21270 );
nand ( n47372 , n47371 , n21291 );
or ( n47373 , n47372 , n21264 );
nand ( n47374 , n47373 , n36457 );
and ( n47375 , n47372 , n21264 );
or ( n47376 , n47374 , n47375 );
not ( n47377 , n21499 );
and ( n47378 , n45261 , n21484 );
not ( n47379 , n21503 );
and ( n47380 , n47378 , n47379 );
not ( n47381 , n47380 );
or ( n47382 , n47377 , n47381 );
or ( n47383 , n47380 , n21499 );
nand ( n47384 , n47382 , n47383 );
and ( n47385 , n47384 , n36443 );
and ( n47386 , n21751 , RI15b57c78_860);
nor ( n47387 , n47385 , n47386 );
nand ( n47388 , n47376 , n47387 );
nor ( n47389 , n47370 , n47388 );
and ( n47390 , n21788 , RI15b56d78_828);
and ( n47391 , n40402 , n21770 );
not ( n47392 , n21887 );
and ( n47393 , n47392 , n17540 );
not ( n47394 , n47392 );
and ( n47395 , n47394 , RI15b56d78_828);
nor ( n47396 , n47393 , n47395 );
and ( n47397 , n47396 , n384127 );
nor ( n47398 , n47390 , n47391 , n47397 );
nand ( n47399 , n47389 , n47398 );
buf ( n47400 , n47399 );
buf ( n47401 , n35651 );
buf ( n47402 , n22716 );
buf ( n47403 , n32672 );
buf ( n47404 , n381004 );
buf ( n47405 , n22402 );
and ( n47406 , n41572 , n34931 );
nor ( n47407 , n47406 , n35114 );
or ( n47408 , n47407 , n34957 );
and ( n47409 , n35118 , n41579 );
and ( n47410 , n20631 , RI15b46338_260);
nor ( n47411 , n47409 , n47410 );
nand ( n47412 , n385213 , RI15b47940_307);
nand ( n47413 , n47408 , n47411 , n47412 );
buf ( n47414 , n47413 );
buf ( n47415 , n22788 );
not ( n47416 , n383163 );
not ( n47417 , n21789 );
or ( n47418 , n47416 , n47417 );
nand ( n47419 , n47418 , RI15b566e8_814);
not ( n47420 , n37718 );
not ( n47421 , n37721 );
or ( n47422 , n47420 , n47421 );
nand ( n47423 , n47422 , n21740 );
nand ( n47424 , n47419 , n37716 , n47423 );
buf ( n47425 , n47424 );
and ( n47426 , n22646 , RI15b45e10_249);
and ( n47427 , n22648 , RI15b52278_668);
nor ( n47428 , n47426 , n47427 );
not ( n47429 , n47428 );
buf ( n47430 , n47429 );
buf ( n47431 , n22738 );
buf ( n47432 , n381006 );
buf ( n47433 , n35649 );
or ( n47434 , n383180 , n380747 );
not ( n47435 , n380776 );
and ( n47436 , n47435 , RI15b587b8_884);
or ( n47437 , n383184 , n380744 );
or ( n47438 , n32696 , n380785 );
or ( n47439 , n380768 , n383192 );
nand ( n47440 , n47437 , n47438 , n47439 );
nor ( n47441 , n47436 , n47440 );
nand ( n47442 , n47434 , n47441 );
buf ( n47443 , n47442 );
not ( n47444 , n31700 );
nand ( n47445 , n39671 , n379319 );
not ( n47446 , n47445 );
nand ( n47447 , n47446 , n379391 );
not ( n47448 , n47447 );
or ( n47449 , n47444 , n47448 );
not ( n47450 , n379045 );
nand ( n47451 , n47449 , n47450 );
nor ( n47452 , n41195 , n47450 );
not ( n47453 , n47452 );
not ( n47454 , n47445 );
or ( n47455 , n47453 , n47454 );
nand ( n47456 , n31712 , RI15b52278_668);
and ( n47457 , n45303 , n47456 );
nand ( n47458 , n47455 , n47457 );
not ( n47459 , n47458 );
nand ( n47460 , n47451 , n47459 );
buf ( n47461 , n47460 );
buf ( n47462 , n379893 );
buf ( n47463 , n22738 );
and ( n47464 , n31792 , n384595 );
or ( n47465 , n31771 , n384234 );
or ( n47466 , n384348 , n32378 );
or ( n47467 , n32640 , n31779 );
nand ( n47468 , n47465 , n47466 , n47467 );
nor ( n47469 , n47464 , n47468 );
nand ( n47470 , n32577 , n47469 );
buf ( n47471 , n47470 );
buf ( n47472 , n381872 );
not ( n47473 , n383357 );
and ( n47474 , n47473 , RI15b4b3d8_432);
buf ( n47475 , n19959 );
not ( n47476 , n47475 );
not ( n47477 , n22377 );
or ( n47478 , n47476 , n47477 );
nand ( n47479 , n47478 , n383364 );
and ( n47480 , n47479 , RI15b495d8_368);
or ( n47481 , n22359 , n47475 , RI15b495d8_368);
and ( n47482 , n383358 , RI15b4b3d8_432);
nor ( n47483 , n383355 , n383358 , RI15b4b3d8_432);
nor ( n47484 , n47482 , n47483 );
or ( n47485 , n20564 , n47484 );
nand ( n47486 , n47481 , n47485 );
nor ( n47487 , n47474 , n47480 , n47486 );
or ( n47488 , n47487 , n20519 );
not ( n47489 , n19741 );
not ( n47490 , n47489 );
not ( n47491 , n19918 );
and ( n47492 , n47490 , n47491 );
not ( n47493 , n22350 );
nor ( n47494 , n47492 , n47493 );
or ( n47495 , n47494 , n19748 );
and ( n47496 , n383353 , n47489 , n19748 );
or ( n47497 , n20639 , n382253 );
or ( n47498 , n19746 , n22390 );
nand ( n47499 , n47497 , n47498 , n384692 );
nor ( n47500 , n47496 , n47499 );
nand ( n47501 , n47488 , n47495 , n47500 );
buf ( n47502 , n47501 );
buf ( n47503 , n381490 );
buf ( n47504 , n22479 );
or ( n47505 , n22425 , n379787 );
and ( n47506 , n383409 , RI15b61cc8_1202);
not ( n47507 , n383473 );
nor ( n47508 , n47507 , n383490 );
or ( n47509 , n47508 , RI15b62bc8_1234);
and ( n47510 , n22450 , n379787 );
not ( n47511 , n40953 );
and ( n47512 , n22471 , n47511 );
nor ( n47513 , n47510 , n47512 );
nand ( n47514 , n47509 , n47513 );
nor ( n47515 , n47506 , n47514 );
not ( n47516 , n383482 );
and ( n47517 , n47516 , n43415 );
or ( n47518 , n383464 , n383467 );
nand ( n47519 , n47518 , n19598 );
and ( n47520 , n47519 , RI15b62bc8_1234);
nor ( n47521 , n47517 , n47520 );
nand ( n47522 , n47505 , n47515 , n47521 );
buf ( n47523 , n47522 );
buf ( n47524 , n381872 );
buf ( n47525 , n381707 );
buf ( n47526 , n22653 );
not ( n47527 , RI15b5fa90_1129);
not ( n47528 , n383601 );
or ( n47529 , n47527 , n47528 );
xor ( n47530 , n383520 , n383521 );
and ( n47531 , n383505 , n47530 );
and ( n47532 , n383607 , RI15b5f310_1113);
nor ( n47533 , n47531 , n47532 );
nand ( n47534 , n47529 , n47533 );
buf ( n47535 , n47534 );
buf ( n47536 , n22009 );
or ( n47537 , n36238 , n35624 );
not ( n47538 , RI15b4f410_569);
or ( n47539 , n47538 , n35635 );
not ( n47540 , n35640 );
and ( n47541 , n47540 , n32711 );
not ( n47542 , n35622 );
and ( n47543 , n383803 , n47542 );
and ( n47544 , n36261 , n35638 );
nor ( n47545 , n47541 , n47543 , n47544 );
nand ( n47546 , n47537 , n47539 , n47545 );
buf ( n47547 , n47546 );
and ( n47548 , n40674 , RI15b54348_738);
not ( n47549 , n379396 );
and ( n47550 , n47549 , RI15b523e0_671);
nor ( n47551 , n47548 , n47550 );
not ( n47552 , n47551 );
buf ( n47553 , n47552 );
not ( n47554 , n384283 );
not ( n47555 , n47554 );
not ( n47556 , n32540 );
or ( n47557 , n47555 , n47556 );
nand ( n47558 , n47557 , n37578 );
and ( n47559 , n47558 , n384392 );
buf ( n47560 , n32554 );
not ( n47561 , n47560 );
not ( n47562 , n384570 );
and ( n47563 , n47561 , n47562 );
and ( n47564 , n47560 , n384570 );
nor ( n47565 , n47563 , n47564 );
not ( n47566 , n19287 );
or ( n47567 , n47565 , n47566 );
not ( n47568 , n384409 );
not ( n47569 , n384442 );
or ( n47570 , n47568 , n47569 );
or ( n47571 , n384442 , n384409 );
nand ( n47572 , n47570 , n47571 );
and ( n47573 , n47572 , n37599 );
and ( n47574 , n19513 , RI15b64158_1280);
nor ( n47575 , n47573 , n47574 );
nand ( n47576 , n47567 , n47575 );
nor ( n47577 , n47559 , n47576 );
not ( n47578 , n31793 );
not ( n47579 , n384570 );
and ( n47580 , n47578 , n47579 );
or ( n47581 , n31771 , n384279 );
and ( n47582 , n42115 , n47554 );
not ( n47583 , n384409 );
and ( n47584 , n31778 , n47583 );
nor ( n47585 , n47582 , n47584 );
nand ( n47586 , n47581 , n47585 );
nor ( n47587 , n47580 , n47586 );
nand ( n47588 , n47577 , n47587 );
buf ( n47589 , n47588 );
buf ( n47590 , n384203 );
buf ( n47591 , n32255 );
not ( n47592 , n382287 );
xor ( n47593 , n382261 , n47592 );
nand ( n47594 , n44071 , n47593 );
not ( n47595 , n382080 );
buf ( n47596 , n382449 );
not ( n47597 , n47596 );
or ( n47598 , n47595 , n47597 );
nand ( n47599 , n47598 , n32023 );
nand ( n47600 , n47599 , n382456 );
not ( n47601 , n47596 );
not ( n47602 , n32035 );
nand ( n47603 , n47601 , n47602 , n382457 );
and ( n47604 , n382523 , RI15b4b450_433);
and ( n47605 , n32974 , RI15b45258_224);
nor ( n47606 , n47604 , n47605 );
nand ( n47607 , n47594 , n47600 , n47603 , n47606 );
buf ( n47608 , n47607 );
buf ( n47609 , n382069 );
buf ( n47610 , n19653 );
buf ( n47611 , n22402 );
buf ( n47612 , n384700 );
and ( n47613 , n34885 , RI15b60a08_1162);
not ( n47614 , n379794 );
and ( n47615 , n47614 , RI15b5d858_1056);
nor ( n47616 , n47613 , n47615 );
not ( n47617 , n47616 );
buf ( n47618 , n47617 );
buf ( n47619 , n22007 );
and ( n47620 , n34854 , n34855 );
not ( n47621 , n34854 );
and ( n47622 , n47621 , n31509 );
nor ( n47623 , n47620 , n47622 );
not ( n47624 , n47623 );
not ( n47625 , n379343 );
or ( n47626 , n47624 , n47625 );
buf ( n47627 , n379369 );
not ( n47628 , n47627 );
not ( n47629 , n31616 );
or ( n47630 , n47629 , n379367 );
nand ( n47631 , n47630 , n379383 );
not ( n47632 , n47631 );
or ( n47633 , n47628 , n47632 );
or ( n47634 , n47631 , n47627 );
nand ( n47635 , n47633 , n47634 );
and ( n47636 , n47635 , n379391 );
and ( n47637 , n379394 , RI15b57840_851);
and ( n47638 , n379398 , RI15b51648_642);
nor ( n47639 , n47636 , n47637 , n47638 );
nand ( n47640 , n47626 , n47639 );
buf ( n47641 , n47640 );
buf ( n47642 , n385112 );
nand ( n47643 , n381568 , n35783 );
not ( n47644 , n47643 );
not ( n47645 , n47644 );
not ( n47646 , n381507 );
or ( n47647 , n47645 , n47646 );
or ( n47648 , n380743 , n381541 );
not ( n47649 , n47648 );
and ( n47650 , n381524 , n47649 );
and ( n47651 , n47648 , n47643 , n381601 );
nor ( n47652 , n47651 , n19630 );
nor ( n47653 , n380755 , n33231 );
or ( n47654 , n47652 , n47653 );
nand ( n47655 , n47654 , n19595 );
or ( n47656 , n380764 , n380728 );
nand ( n47657 , n47655 , n47656 );
and ( n47658 , n47657 , n380775 );
or ( n47659 , n47658 , n18429 );
not ( n47660 , n381550 );
not ( n47661 , n47656 );
nor ( n47662 , n47653 , n47661 );
or ( n47663 , n47652 , n47662 );
or ( n47664 , n47660 , n47663 );
or ( n47665 , n47656 , n381560 );
nand ( n47666 , n47659 , n47664 , n47665 );
nor ( n47667 , n47650 , n47666 );
nand ( n47668 , n47647 , n47667 );
buf ( n47669 , n47668 );
or ( n47670 , n380001 , n379973 );
and ( n47671 , n35734 , RI15b4fc80_587);
and ( n47672 , n380061 , RI15b4ed80_555);
and ( n47673 , n382793 , RI15b4dac0_515);
and ( n47674 , n35739 , RI15b4d340_499);
nor ( n47675 , n47672 , n47673 , n47674 );
and ( n47676 , n381651 , RI15b4de80_523);
and ( n47677 , n382806 , RI15b4e9c0_547);
nor ( n47678 , n47676 , n47677 );
and ( n47679 , n382825 , RI15b4d700_507);
not ( n47680 , n382800 );
and ( n47681 , n47680 , RI15b4e600_539);
nor ( n47682 , n47679 , n47681 );
nand ( n47683 , n35748 , RI15b4e240_531);
nand ( n47684 , n47675 , n47678 , n47682 , n47683 );
and ( n47685 , n381646 , n47684 );
and ( n47686 , n35732 , RI15b4c800_475);
nor ( n47687 , n47671 , n47685 , n47686 );
and ( n47688 , n35754 , RI15b4f500_571);
and ( n47689 , n35756 , RI15b4f8c0_579);
nor ( n47690 , n47688 , n47689 );
and ( n47691 , n35759 , RI15b4f140_563);
and ( n47692 , n35761 , RI15b4c440_467);
nor ( n47693 , n47691 , n47692 );
and ( n47694 , n35764 , RI15b4cf80_491);
and ( n47695 , n35766 , RI15b4cbc0_483);
nor ( n47696 , n47694 , n47695 );
nand ( n47697 , n47687 , n47690 , n47693 , n47696 );
and ( n47698 , n47697 , n381696 );
and ( n47699 , n379972 , n379973 );
not ( n47700 , n379972 );
and ( n47701 , n47700 , RI15b56058_800);
nor ( n47702 , n47699 , n47701 );
and ( n47703 , n47702 , n379949 );
nor ( n47704 , n47698 , n47703 );
nand ( n47705 , n47670 , n47704 );
buf ( n47706 , n47705 );
buf ( n47707 , n383498 );
buf ( n47708 , RI15b47aa8_310);
buf ( n47709 , n384700 );
buf ( n47710 , n17499 );
and ( n47711 , n385164 , RI15b50d60_623);
or ( n47712 , n33652 , n37952 );
or ( n47713 , n37924 , n385170 );
or ( n47714 , n37968 , n385178 );
nand ( n47715 , n47712 , n47713 , n47714 );
nor ( n47716 , n47711 , n47715 );
nand ( n47717 , n41160 , n47716 );
buf ( n47718 , n47717 );
not ( n47719 , n36568 );
nand ( n47720 , n47719 , n379785 );
not ( n47721 , n47720 );
not ( n47722 , n36574 );
or ( n47723 , n47721 , n47722 );
buf ( n47724 , n36569 );
nand ( n47725 , n47723 , n47724 );
nor ( n47726 , n47719 , n36569 );
nand ( n47727 , n36502 , n47726 );
not ( n47728 , n34510 );
not ( n47729 , n47728 );
buf ( n47730 , n34492 );
not ( n47731 , n47730 );
or ( n47732 , n47729 , n47731 );
or ( n47733 , n47730 , n47728 );
nand ( n47734 , n47732 , n47733 );
not ( n47735 , n34645 );
and ( n47736 , n47734 , n47735 );
and ( n47737 , n379783 , RI15b64338_1284);
and ( n47738 , n34651 , RI15b5e140_1075);
nor ( n47739 , n47736 , n47737 , n47738 );
nand ( n47740 , n47725 , n47727 , n47739 );
buf ( n47741 , n47740 );
buf ( n47742 , n33382 );
buf ( n47743 , n32271 );
not ( n47744 , n386590 );
not ( n47745 , n382912 );
or ( n47746 , n47744 , n47745 );
and ( n47747 , n382931 , n386603 );
not ( n47748 , RI15b59fa0_935);
or ( n47749 , n386612 , n47748 );
or ( n47750 , n40296 , n386624 );
or ( n47751 , n386610 , n382967 );
nand ( n47752 , n47749 , n47750 , n47751 );
nor ( n47753 , n47747 , n47752 );
nand ( n47754 , n47746 , n47753 );
buf ( n47755 , n47754 );
buf ( n47756 , n32676 );
buf ( n47757 , n382069 );
buf ( n47758 , n382888 );
or ( n47759 , n32430 , n47758 );
not ( n47760 , n381317 );
nand ( n47761 , n381417 , n47760 );
and ( n47762 , n386637 , RI15b54f00_763);
and ( n47763 , n381636 , RI15b4eb28_550);
and ( n47764 , n381639 , RI15b4e768_542);
nor ( n47765 , n47763 , n47764 );
and ( n47766 , n381643 , RI15b4eee8_558);
and ( n47767 , n41896 , RI15b4dc28_518);
and ( n47768 , n381657 , RI15b4fde8_590);
nor ( n47769 , n47767 , n47768 );
and ( n47770 , n381661 , RI15b4fa28_582);
and ( n47771 , n381663 , RI15b4f2a8_566);
nor ( n47772 , n47770 , n47771 );
and ( n47773 , n381667 , RI15b4d4a8_502);
and ( n47774 , n381669 , RI15b4d868_510);
nor ( n47775 , n47773 , n47774 );
and ( n47776 , n381672 , RI15b4dfe8_526);
and ( n47777 , n381674 , RI15b4f668_574);
nor ( n47778 , n47776 , n47777 );
nand ( n47779 , n47769 , n47772 , n47775 , n47778 );
and ( n47780 , n38323 , n47779 );
and ( n47781 , n381680 , RI15b4c968_478);
nor ( n47782 , n47766 , n47780 , n47781 );
and ( n47783 , n381684 , RI15b4c5a8_470);
and ( n47784 , n381686 , RI15b4e3a8_534);
nor ( n47785 , n47783 , n47784 );
and ( n47786 , n381689 , RI15b4cd28_486);
and ( n47787 , n381691 , RI15b4d0e8_494);
nor ( n47788 , n47786 , n47787 );
nand ( n47789 , n47765 , n47782 , n47785 , n47788 );
and ( n47790 , n47789 , n386671 );
not ( n47791 , RI15b54f00_763);
not ( n47792 , n382648 );
not ( n47793 , n47792 );
or ( n47794 , n47791 , n47793 );
or ( n47795 , n47792 , RI15b54f00_763);
nand ( n47796 , n47794 , n47795 );
and ( n47797 , n32439 , n47796 );
nor ( n47798 , n47762 , n47790 , n47797 );
and ( n47799 , n47761 , n47798 );
nand ( n47800 , n47759 , n47799 );
buf ( n47801 , n47800 );
buf ( n47802 , n22408 );
not ( n47803 , n42459 );
buf ( n47804 , n382941 );
nor ( n47805 , n41218 , n47804 );
nor ( n47806 , n47805 , RI15b58650_881);
not ( n47807 , n47806 );
not ( n47808 , n40939 );
not ( n47809 , RI15b58560_879);
not ( n47810 , n41219 );
or ( n47811 , n47809 , n47810 );
nand ( n47812 , n47811 , n19261 );
nand ( n47813 , n47808 , n47812 );
not ( n47814 , n47813 );
or ( n47815 , n47807 , n47814 );
nand ( n47816 , n47815 , n41358 );
not ( n47817 , n47805 );
not ( n47818 , n47817 );
not ( n47819 , n47813 );
or ( n47820 , n47818 , n47819 );
nand ( n47821 , n47820 , RI15b58650_881);
nand ( n47822 , n47816 , n47821 );
or ( n47823 , n47822 , RI15b58740_883);
and ( n47824 , n41358 , n32078 );
nand ( n47825 , n47823 , n47824 );
not ( n47826 , n47825 );
or ( n47827 , n47803 , n47826 );
not ( n47828 , n47822 );
not ( n47829 , n32078 );
and ( n47830 , n47828 , n47829 );
or ( n47831 , RI15b584e8_878 , RI15b5d510_1049);
nand ( n47832 , n47831 , n45723 );
or ( n47833 , n22469 , n43968 , n22428 );
nand ( n47834 , n47833 , n19148 );
not ( n47835 , n47834 );
nand ( n47836 , n40936 , n47832 , n47835 );
nor ( n47837 , n47830 , n47836 );
nand ( n47838 , n47827 , n47837 );
or ( n47839 , n47838 , n22447 );
nand ( n47840 , n47839 , n19201 );
nand ( n47841 , n19590 , n19577 );
and ( n47842 , n47841 , n22428 );
and ( n47843 , n383607 , n22427 );
nor ( n47844 , n47842 , n47843 );
and ( n47845 , n39120 , n47844 , n19512 , n380772 );
nand ( n47846 , n47840 , n47845 );
buf ( n47847 , n47846 );
buf ( n47848 , n385195 );
and ( n47849 , n43983 , n43985 );
not ( n47850 , n43983 );
and ( n47851 , n47850 , n43984 );
nor ( n47852 , n47849 , n47851 );
nand ( n47853 , n47852 , n31601 );
not ( n47854 , n379391 );
buf ( n47855 , n40961 );
not ( n47856 , n47855 );
or ( n47857 , n47854 , n47856 );
nand ( n47858 , n47857 , n31700 );
and ( n47859 , n47858 , n379145 );
or ( n47860 , n41195 , n47855 , n379145 );
and ( n47861 , n379394 , RI15b57b10_857);
and ( n47862 , n47038 , RI15b51918_648);
nor ( n47863 , n47861 , n47862 );
nand ( n47864 , n47860 , n47863 );
nor ( n47865 , n47859 , n47864 );
nand ( n47866 , n47853 , n47865 );
buf ( n47867 , n47866 );
buf ( n47868 , n379844 );
not ( n47869 , n42521 );
nor ( n47870 , n47869 , n21674 );
not ( n47871 , n47870 );
nand ( n47872 , n47871 , n42523 );
nand ( n47873 , n47872 , n21748 );
not ( n47874 , n21312 );
not ( n47875 , n21318 );
and ( n47876 , n47874 , n47875 );
not ( n47877 , n47874 );
and ( n47878 , n47877 , n21318 );
nor ( n47879 , n47876 , n47878 );
and ( n47880 , n47879 , n47263 );
not ( n47881 , n21529 );
and ( n47882 , n47881 , n21535 );
not ( n47883 , n47881 );
and ( n47884 , n47883 , n21534 );
nor ( n47885 , n47882 , n47884 );
not ( n47886 , n21563 );
or ( n47887 , n47885 , n47886 );
or ( n47888 , n21750 , n22611 );
nand ( n47889 , n47887 , n47888 );
nor ( n47890 , n47880 , n47889 );
nand ( n47891 , n47873 , n47890 );
not ( n47892 , n47891 );
and ( n47893 , n385164 , RI15b50838_612);
or ( n47894 , n36693 , n21674 );
or ( n47895 , n47875 , n385170 );
or ( n47896 , n21534 , n385178 );
nand ( n47897 , n47894 , n47895 , n47896 );
nor ( n47898 , n47893 , n47897 );
nand ( n47899 , n47892 , n47898 );
buf ( n47900 , n47899 );
buf ( n47901 , n18226 );
buf ( n47902 , n384996 );
nand ( n47903 , n34617 , n34637 );
not ( n47904 , n34613 );
nand ( n47905 , n47904 , n34622 );
or ( n47906 , n47905 , n33893 );
xor ( n47907 , n33909 , n47906 );
nand ( n47908 , n34620 , n34628 );
not ( n47909 , n47908 );
and ( n47910 , n47905 , n379731 );
not ( n47911 , n47905 );
and ( n47912 , n47911 , n33893 );
nor ( n47913 , n47910 , n47912 );
nand ( n47914 , n47909 , n47913 );
xnor ( n47915 , n47907 , n47914 );
not ( n47916 , n47915 );
buf ( n47917 , n47908 );
and ( n47918 , n47917 , n47913 );
not ( n47919 , n47913 );
nand ( n47920 , n47919 , n34628 , n34633 );
nor ( n47921 , n34630 , n47920 );
nor ( n47922 , n47918 , n47921 );
buf ( n47923 , n47922 );
nand ( n47924 , n47916 , n47923 );
nor ( n47925 , n47903 , n47924 );
not ( n47926 , n33914 );
not ( n47927 , n47906 );
and ( n47928 , n379462 , n47927 );
not ( n47929 , n379462 );
not ( n47930 , n47914 );
and ( n47931 , n47929 , n47930 );
nor ( n47932 , n47928 , n47931 );
nand ( n47933 , n47914 , n47906 );
nand ( n47934 , n47932 , n47933 );
not ( n47935 , n47934 );
or ( n47936 , n47926 , n47935 );
not ( n47937 , n47930 );
nor ( n47938 , n47906 , n33902 );
and ( n47939 , n47937 , n47938 );
nand ( n47940 , n47906 , n33910 );
nor ( n47941 , n47937 , n47940 );
nor ( n47942 , n47939 , n47941 );
nand ( n47943 , n47936 , n47942 );
not ( n47944 , n47943 );
nand ( n47945 , n47944 , n34646 );
or ( n47946 , n47925 , n47945 );
nand ( n47947 , n47922 , n34644 );
nor ( n47948 , n47915 , n47947 );
nand ( n47949 , n47943 , n47948 );
nor ( n47950 , n47903 , n47949 );
and ( n47951 , n379783 , RI15b64860_1295);
and ( n47952 , n34651 , RI15b5e668_1086);
nor ( n47953 , n47951 , n47952 );
not ( n47954 , n47953 );
nor ( n47955 , n47950 , n47954 );
buf ( n47956 , n44382 );
and ( n47957 , n34249 , n44381 , n47956 );
not ( n47958 , n44381 );
nand ( n47959 , n47958 , n379785 );
nand ( n47960 , n34296 , n47959 );
not ( n47961 , n47956 );
and ( n47962 , n47960 , n47961 );
nor ( n47963 , n47957 , n47962 );
nand ( n47964 , n47946 , n47955 , n47963 );
buf ( n47965 , n47964 );
not ( n47966 , n22373 );
and ( n47967 , n47966 , RI15b4b4c8_434);
not ( n47968 , n19963 );
not ( n47969 , n47968 );
not ( n47970 , n22377 );
or ( n47971 , n47969 , n47970 );
nand ( n47972 , n47971 , n383364 );
and ( n47973 , n47972 , RI15b496c8_370);
or ( n47974 , n22359 , n47968 , RI15b496c8_370);
and ( n47975 , n22374 , RI15b4b4c8_434);
nor ( n47976 , n22356 , n22374 , RI15b4b4c8_434);
nor ( n47977 , n47975 , n47976 );
or ( n47978 , n20564 , n47977 );
nand ( n47979 , n47974 , n47978 );
nor ( n47980 , n47967 , n47973 , n47979 );
or ( n47981 , n47980 , n20519 );
not ( n47982 , n19757 );
not ( n47983 , n47982 );
not ( n47984 , n19918 );
and ( n47985 , n47983 , n47984 );
not ( n47986 , n22350 );
nor ( n47987 , n47985 , n47986 );
or ( n47988 , n19764 , n47987 );
and ( n47989 , n22368 , n47982 , n19764 );
or ( n47990 , n20639 , n382099 );
or ( n47991 , n19762 , n22390 );
nand ( n47992 , n47990 , n47991 , n384692 );
nor ( n47993 , n47989 , n47992 );
nand ( n47994 , n47981 , n47988 , n47993 );
buf ( n47995 , n47994 );
buf ( n47996 , n382073 );
buf ( n47997 , n22479 );
buf ( n47998 , n381081 );
buf ( n47999 , n35651 );
nand ( n48000 , n383432 , n31965 );
and ( n48001 , n384642 , n48000 );
not ( n48002 , RI15b639d8_1264);
nor ( n48003 , n48001 , n48002 );
not ( n48004 , n387012 );
not ( n48005 , n48004 );
or ( n48006 , n31971 , n383432 , RI15b639d8_1264);
or ( n48007 , n383462 , n383597 );
nand ( n48008 , n48006 , n48007 );
or ( n48009 , n48005 , n48008 );
nor ( n48010 , n42111 , n48003 , n48009 );
nand ( n48011 , n42091 , n48010 );
buf ( n48012 , n48011 );
buf ( n48013 , n19651 );
buf ( n48014 , n22479 );
buf ( n48015 , n382049 );
buf ( n48016 , n387159 );
or ( n48017 , n381056 , n32614 );
or ( n48018 , n32805 , n35572 );
and ( n48019 , n37118 , RI15b49b00_379);
not ( n48020 , n37118 );
and ( n48021 , n48020 , n32614 );
nor ( n48022 , n48019 , n48021 );
or ( n48023 , n37109 , n48022 );
nand ( n48024 , n48017 , n48018 , n48023 );
buf ( n48025 , n48024 );
not ( n48026 , RI15b53da8_726);
not ( n48027 , n32244 );
or ( n48028 , n48026 , n48027 );
and ( n48029 , n32247 , RI15b653a0_1319);
and ( n48030 , n32249 , RI15b60210_1145);
nor ( n48031 , n48029 , n48030 );
nand ( n48032 , n48028 , n48031 );
buf ( n48033 , n48032 );
buf ( n48034 , n382052 );
or ( n48035 , n39265 , n35582 );
nand ( n48036 , n381017 , RI15b53358_704);
nand ( n48037 , n48035 , n48036 );
buf ( n48038 , n48037 );
buf ( n48039 , n22653 );
buf ( n48040 , n32255 );
or ( n48041 , n381056 , n19962 );
or ( n48042 , n20409 , n381062 );
not ( n48043 , n32814 );
and ( n48044 , n48043 , RI15b49650_369);
not ( n48045 , n48043 );
and ( n48046 , n48045 , n19962 );
nor ( n48047 , n48044 , n48046 );
or ( n48048 , n48047 , n381077 );
nand ( n48049 , n48041 , n48042 , n48048 );
buf ( n48050 , n48049 );
buf ( n48051 , n384700 );
not ( n48052 , n37495 );
not ( n48053 , n48052 );
not ( n48054 , n33370 );
or ( n48055 , n48053 , n48054 );
and ( n48056 , n33196 , n37498 );
not ( n48057 , RI15b427b0_133);
or ( n48058 , n37507 , n48057 );
or ( n48059 , n22241 , n37512 );
or ( n48060 , n37505 , n33201 );
nand ( n48061 , n48058 , n48059 , n48060 );
nor ( n48062 , n48056 , n48061 );
nand ( n48063 , n48055 , n48062 );
buf ( n48064 , n48063 );
buf ( n48065 , n379847 );
buf ( n48066 , n380942 );
buf ( n48067 , n22740 );
buf ( n48068 , n380903 );
not ( n48069 , n379974 );
and ( n48070 , n48069 , n379949 );
nor ( n48071 , n48070 , n380000 );
or ( n48072 , n48071 , n22580 );
and ( n48073 , n379974 , n379949 , n22580 );
and ( n48074 , n43875 , n38347 );
nor ( n48075 , n48073 , n48074 );
nand ( n48076 , n48072 , n48075 );
buf ( n48077 , n48076 );
buf ( n48078 , RI15b478c8_306);
buf ( n48079 , n379895 );
not ( n48080 , n47644 );
not ( n48081 , n381589 );
or ( n48082 , n48080 , n48081 );
and ( n48083 , n381596 , n47649 );
or ( n48084 , n47658 , n18735 );
or ( n48085 , n32420 , n47663 );
or ( n48086 , n47656 , n381621 );
nand ( n48087 , n48084 , n48085 , n48086 );
nor ( n48088 , n48083 , n48087 );
nand ( n48089 , n48082 , n48088 );
buf ( n48090 , n48089 );
buf ( n48091 , n385197 );
buf ( n48092 , n22479 );
buf ( n48093 , n382071 );
buf ( n48094 , n385112 );
buf ( n48095 , n380940 );
or ( n48096 , n380001 , n21952 );
and ( n48097 , n380010 , RI15b4c530_469);
and ( n48098 , n379953 , n21952 );
not ( n48099 , n379953 );
and ( n48100 , n48099 , RI15b559c8_786);
nor ( n48101 , n48098 , n48100 );
and ( n48102 , n379949 , n48101 );
nor ( n48103 , n48097 , n48102 );
nand ( n48104 , n48096 , n48103 );
buf ( n48105 , n48104 );
not ( n48106 , n36395 );
not ( n48107 , n33400 );
or ( n48108 , n48106 , n48107 );
and ( n48109 , n33415 , n36401 );
or ( n48110 , n36410 , n18463 );
or ( n48111 , n36293 , n36416 );
or ( n48112 , n36408 , n33443 );
nand ( n48113 , n48110 , n48111 , n48112 );
nor ( n48114 , n48109 , n48113 );
nand ( n48115 , n48108 , n48114 );
buf ( n48116 , n48115 );
not ( n48117 , n47644 );
not ( n48118 , n380703 );
or ( n48119 , n48117 , n48118 );
and ( n48120 , n380719 , n47649 );
or ( n48121 , n47658 , n19036 );
or ( n48122 , n380782 , n47663 );
or ( n48123 , n47656 , n380790 );
nand ( n48124 , n48121 , n48122 , n48123 );
nor ( n48125 , n48120 , n48124 );
nand ( n48126 , n48119 , n48125 );
buf ( n48127 , n48126 );
buf ( n48128 , n379895 );
buf ( n48129 , RI15b47c88_314);
not ( n48130 , RI15b55fe0_799);
not ( n48131 , n380000 );
or ( n48132 , n48130 , n48131 );
and ( n48133 , n35734 , RI15b4fc08_586);
and ( n48134 , n380061 , RI15b4ed08_554);
not ( n48135 , n382792 );
and ( n48136 , n48135 , RI15b4da48_514);
and ( n48137 , n35739 , RI15b4d2c8_498);
nor ( n48138 , n48134 , n48136 , n48137 );
and ( n48139 , n43671 , RI15b4de08_522);
and ( n48140 , n382806 , RI15b4e948_546);
nor ( n48141 , n48139 , n48140 );
and ( n48142 , n382780 , RI15b4d688_506);
and ( n48143 , n382801 , RI15b4e588_538);
nor ( n48144 , n48142 , n48143 );
nand ( n48145 , n35748 , RI15b4e1c8_530);
nand ( n48146 , n48138 , n48141 , n48144 , n48145 );
and ( n48147 , n381646 , n48146 );
and ( n48148 , n35732 , RI15b4c788_474);
nor ( n48149 , n48133 , n48147 , n48148 );
and ( n48150 , n35754 , RI15b4f488_570);
and ( n48151 , n35756 , RI15b4f848_578);
nor ( n48152 , n48150 , n48151 );
and ( n48153 , n35759 , RI15b4f0c8_562);
and ( n48154 , n35761 , RI15b4c3c8_466);
nor ( n48155 , n48153 , n48154 );
and ( n48156 , n35764 , RI15b4cf08_490);
and ( n48157 , n35766 , RI15b4cb48_482);
nor ( n48158 , n48156 , n48157 );
nand ( n48159 , n48149 , n48152 , n48155 , n48158 );
and ( n48160 , n48159 , n381696 );
not ( n48161 , RI15b55fe0_799);
not ( n48162 , n379970 );
or ( n48163 , n48161 , n48162 );
or ( n48164 , n379970 , RI15b55fe0_799);
nand ( n48165 , n48163 , n48164 );
and ( n48166 , n48165 , n379949 );
nor ( n48167 , n48160 , n48166 );
nand ( n48168 , n48132 , n48167 );
buf ( n48169 , n48168 );
buf ( n48170 , n22479 );
buf ( n48171 , n381006 );
buf ( n48172 , n383345 );
buf ( n48173 , n32672 );
buf ( n48174 , n18226 );
nand ( n48175 , n46509 , n35043 );
buf ( n48176 , n48175 );
nor ( n48177 , n48176 , n34930 );
or ( n48178 , n48177 , n35114 );
not ( n48179 , n35015 );
nand ( n48180 , n48178 , n48179 );
nor ( n48181 , n35117 , n48179 );
not ( n48182 , n48181 );
not ( n48183 , n48176 );
or ( n48184 , n48182 , n48183 );
and ( n48185 , n385213 , RI15b47c88_314);
and ( n48186 , n20631 , RI15b46680_267);
nor ( n48187 , n48185 , n48186 );
nand ( n48188 , n48184 , n48187 );
not ( n48189 , n48188 );
nand ( n48190 , n48180 , n48189 );
buf ( n48191 , n48190 );
buf ( n48192 , n382073 );
not ( n48193 , n40338 );
or ( n48194 , n48193 , n22595 );
not ( n48195 , n380012 );
not ( n48196 , n48195 );
not ( n48197 , n46750 );
and ( n48198 , n48196 , n48197 );
and ( n48199 , n40345 , n40339 );
nor ( n48200 , n48198 , n48199 );
nand ( n48201 , n48194 , n48200 );
buf ( n48202 , n48201 );
buf ( n48203 , n379847 );
buf ( n48204 , RI15b5e050_1073);
buf ( n48205 , n385197 );
buf ( n48206 , n383498 );
not ( n48207 , n380235 );
not ( n48208 , n33400 );
or ( n48209 , n48207 , n48208 );
and ( n48210 , n33415 , n380745 );
or ( n48211 , n380776 , n18496 );
or ( n48212 , n36293 , n380785 );
or ( n48213 , n380768 , n33443 );
nand ( n48214 , n48211 , n48212 , n48213 );
nor ( n48215 , n48210 , n48214 );
nand ( n48216 , n48209 , n48215 );
buf ( n48217 , n48216 );
buf ( n48218 , n19832 );
or ( n48219 , n48218 , n31799 );
nand ( n48220 , n48219 , n19938 );
nand ( n48221 , n48220 , n19838 );
not ( n48222 , n19838 );
nand ( n48223 , n48222 , n32502 , n48218 );
and ( n48224 , n20641 , RI15b4b9f0_445);
buf ( n48225 , n19981 );
not ( n48226 , n48225 );
and ( n48227 , n48226 , n31806 );
nor ( n48228 , n48227 , n31809 );
or ( n48229 , n48228 , n37121 );
not ( n48230 , n20551 );
and ( n48231 , n48230 , RI15b4b9f0_445);
not ( n48232 , n48230 );
and ( n48233 , n48232 , n382117 );
nor ( n48234 , n48231 , n48233 );
or ( n48235 , n48234 , n22354 );
and ( n48236 , n48225 , n22361 , n37121 );
not ( n48237 , RI15b4aaf0_413);
or ( n48238 , n42326 , n48237 );
nand ( n48239 , n48238 , n31821 );
nor ( n48240 , n48236 , n48239 );
nand ( n48241 , n48229 , n48235 , n48240 );
nor ( n48242 , n48224 , n48241 );
nand ( n48243 , n48221 , n48223 , n48242 );
buf ( n48244 , n48243 );
buf ( n48245 , n22479 );
not ( n48246 , n39551 );
not ( n48247 , n384338 );
or ( n48248 , n48246 , n48247 );
nand ( n48249 , n48248 , n384360 );
and ( n48250 , n48249 , n31923 );
and ( n48251 , n32627 , n384543 );
not ( n48252 , n32627 );
and ( n48253 , n48252 , n32628 );
nor ( n48254 , n48251 , n48253 );
not ( n48255 , n39045 );
or ( n48256 , n48254 , n48255 );
and ( n48257 , n32642 , n32643 );
not ( n48258 , n32642 );
and ( n48259 , n48258 , n384455 );
nor ( n48260 , n48257 , n48259 );
and ( n48261 , n48260 , n31882 );
and ( n48262 , n19513 , RI15b643b0_1285);
nor ( n48263 , n48261 , n48262 );
nand ( n48264 , n48256 , n48263 );
nor ( n48265 , n48250 , n48264 );
and ( n48266 , n384638 , RI15b634b0_1253);
or ( n48267 , n384652 , n383442 , RI15b634b0_1253);
or ( n48268 , n386897 , n22775 );
nand ( n48269 , n48267 , n48268 );
nor ( n48270 , n48266 , n48269 );
nand ( n48271 , n48265 , n48270 );
buf ( n48272 , n48271 );
buf ( n48273 , n18226 );
buf ( n48274 , n19651 );
buf ( n48275 , n380865 );
buf ( n48276 , n22716 );
buf ( n48277 , n32160 );
buf ( n48278 , n32981 );
buf ( n48279 , n382537 );
not ( n48280 , n38485 );
and ( n48281 , n48280 , RI15b62790_1225);
not ( n48282 , n48280 );
not ( n48283 , RI15b62790_1225);
and ( n48284 , n48282 , n48283 );
nor ( n48285 , n48281 , n48284 );
or ( n48286 , n48285 , n384024 );
and ( n48287 , n384022 , RI15b62790_1225);
not ( n48288 , n39777 );
and ( n48289 , n41741 , n48288 );
nor ( n48290 , n48287 , n48289 );
nand ( n48291 , n48286 , n48290 );
buf ( n48292 , n48291 );
or ( n48293 , n36238 , n39693 );
not ( n48294 , n39703 );
and ( n48295 , n48294 , RI15b4c710_473);
not ( n48296 , n36256 );
or ( n48297 , n39707 , n48296 );
or ( n48298 , n39691 , n383802 );
or ( n48299 , n39701 , n42402 );
nand ( n48300 , n48297 , n48298 , n48299 );
nor ( n48301 , n48295 , n48300 );
nand ( n48302 , n48293 , n48301 );
buf ( n48303 , n48302 );
or ( n48304 , n22315 , n38065 );
and ( n48305 , n22326 , n38067 );
not ( n48306 , RI15b42d50_145);
or ( n48307 , n38077 , n48306 );
or ( n48308 , n22334 , n38081 );
or ( n48309 , n38075 , n22336 );
nand ( n48310 , n48307 , n48308 , n48309 );
nor ( n48311 , n48305 , n48310 );
nand ( n48312 , n48304 , n48311 );
buf ( n48313 , n48312 );
buf ( n48314 , n379403 );
buf ( n48315 , n384203 );
buf ( n48316 , n382067 );
buf ( n48317 , n381566 );
buf ( n48318 , n385112 );
buf ( n48319 , n383498 );
buf ( n48320 , n22653 );
buf ( n48321 , n381004 );
or ( n48322 , n40166 , n386319 );
not ( n48323 , n46595 );
and ( n48324 , n386540 , RI15b43d40_179);
and ( n48325 , n386549 , n385440 );
and ( n48326 , n386556 , n386128 );
nor ( n48327 , n48324 , n48325 , n48326 );
nand ( n48328 , n48322 , n48323 , n48327 );
buf ( n48329 , n48328 );
or ( n48330 , n31149 , n385002 );
and ( n48331 , n31161 , n385006 );
not ( n48332 , RI15b4e240_531);
or ( n48333 , n385019 , n48332 );
or ( n48334 , n32452 , n385023 );
or ( n48335 , n385017 , n31184 );
nand ( n48336 , n48333 , n48334 , n48335 );
nor ( n48337 , n48331 , n48336 );
nand ( n48338 , n48330 , n48337 );
buf ( n48339 , n48338 );
buf ( n48340 , n387159 );
buf ( n48341 , n384218 );
buf ( n48342 , n32981 );
and ( n48343 , n22435 , RI15b60cd8_1168);
not ( n48344 , n385035 );
nor ( n48345 , n48343 , n48344 );
or ( n48346 , n22427 , n48345 );
and ( n48347 , n385043 , RI15b60738_1156 , RI15b60be8_1166);
and ( n48348 , n31039 , RI15b3f9c0_35);
nor ( n48349 , n48347 , n48348 );
nand ( n48350 , n48346 , n48349 , n383589 );
buf ( n48351 , n48350 );
not ( n48352 , n31806 );
not ( n48353 , n19989 );
or ( n48354 , n48352 , n48353 );
nand ( n48355 , n48354 , n380875 );
and ( n48356 , n48355 , RI15b49e48_386);
not ( n48357 , n19989 );
nand ( n48358 , n48357 , n32511 , n19990 );
not ( n48359 , n20555 );
or ( n48360 , n48359 , n382125 , RI15b4bc48_450);
or ( n48361 , n382126 , RI15b4bbd0_449);
nand ( n48362 , n48360 , n48361 );
and ( n48363 , n20647 , n48362 );
and ( n48364 , n387180 , RI15b4ad48_418);
nor ( n48365 , n48363 , n48364 );
nand ( n48366 , n48358 , n48365 );
and ( n48367 , n20568 , n48359 );
nor ( n48368 , n48367 , n20641 );
nor ( n48369 , n48368 , n382126 );
nor ( n48370 , n48356 , n48366 , n48369 );
not ( n48371 , n19921 );
not ( n48372 , n48371 );
not ( n48373 , n19869 );
not ( n48374 , n48373 );
or ( n48375 , n48372 , n48374 );
nand ( n48376 , n48375 , n19942 );
nand ( n48377 , n48376 , n19875 );
or ( n48378 , n48373 , n387170 , n19875 );
nand ( n48379 , n48370 , n48377 , n48378 );
buf ( n48380 , n48379 );
buf ( n48381 , n22406 );
buf ( n48382 , n22005 );
or ( n48383 , n384623 , n383435 );
nand ( n48384 , n48383 , n32581 );
and ( n48385 , n48384 , RI15b63258_1248);
or ( n48386 , n384652 , n383434 , RI15b63258_1248);
not ( n48387 , n386862 );
or ( n48388 , n48387 , n22775 );
nand ( n48389 , n48386 , n48388 );
nor ( n48390 , n48385 , n48389 );
nand ( n48391 , n47577 , n48390 );
buf ( n48392 , n48391 );
buf ( n48393 , n382052 );
buf ( n48394 , n381081 );
buf ( n48395 , n22408 );
or ( n48396 , n382679 , n382662 );
and ( n48397 , n382692 , n383725 );
and ( n48398 , n382661 , RI15b55338_772);
not ( n48399 , n382661 );
and ( n48400 , n48399 , n382662 );
nor ( n48401 , n48398 , n48400 );
or ( n48402 , n48401 , n382625 );
not ( n48403 , n386667 );
and ( n48404 , n380123 , RI15b4f6e0_575);
and ( n48405 , n380125 , RI15b4faa0_583);
nor ( n48406 , n48404 , n48405 );
and ( n48407 , n380061 , RI15b4ef60_559);
and ( n48408 , n381650 , RI15b4e060_527);
and ( n48409 , n380115 , RI15b4c620_471);
nor ( n48410 , n48407 , n48408 , n48409 );
and ( n48411 , n382841 , RI15b4dca0_519);
and ( n48412 , n382788 , RI15b4d160_495);
and ( n48413 , n382780 , RI15b4d8e0_511);
nor ( n48414 , n48411 , n48412 , n48413 );
nand ( n48415 , n35748 , RI15b4e420_535);
nand ( n48416 , n48406 , n48410 , n48414 , n48415 );
and ( n48417 , n380128 , RI15b4fe60_591);
and ( n48418 , n380099 , RI15b4f320_567);
nor ( n48419 , n48417 , n48418 );
and ( n48420 , n382849 , RI15b4e7e0_543);
and ( n48421 , n382813 , RI15b4c9e0_479);
nor ( n48422 , n48420 , n48421 );
and ( n48423 , n382856 , RI15b4eba0_551);
and ( n48424 , n379878 , RI15b4cda0_487);
nor ( n48425 , n48423 , n48424 );
nand ( n48426 , n35739 , RI15b4d520_503);
nand ( n48427 , n48419 , n48422 , n48425 , n48426 );
or ( n48428 , n48416 , n48427 );
nand ( n48429 , n48428 , n35736 );
or ( n48430 , n48403 , n48429 );
nand ( n48431 , n48402 , n48430 );
nor ( n48432 , n48397 , n48431 , n33353 );
nand ( n48433 , n48396 , n48432 );
buf ( n48434 , n48433 );
not ( n48435 , n35784 );
not ( n48436 , n37629 );
or ( n48437 , n48435 , n48436 );
and ( n48438 , n37637 , n35790 );
or ( n48439 , n35803 , n18585 );
or ( n48440 , n43001 , n35811 );
or ( n48441 , n35801 , n37646 );
nand ( n48442 , n48439 , n48440 , n48441 );
nor ( n48443 , n48438 , n48442 );
nand ( n48444 , n48437 , n48443 );
buf ( n48445 , n48444 );
buf ( n48446 , n379844 );
buf ( n48447 , n380942 );
buf ( n48448 , n22788 );
not ( n48449 , RI15b53cb8_724);
not ( n48450 , n383170 );
or ( n48451 , n48449 , n48450 );
or ( n48452 , n32400 , n383152 );
nand ( n48453 , n48452 , n383157 );
and ( n48454 , n48453 , n32404 );
and ( n48455 , n32407 , n383143 );
and ( n48456 , n383147 , RI15b526b0_677);
nor ( n48457 , n48454 , n48455 , n48456 );
nand ( n48458 , n48451 , n48457 );
buf ( n48459 , n48458 );
buf ( n48460 , n385112 );
not ( n48461 , n35145 );
not ( n48462 , n37629 );
or ( n48463 , n48461 , n48462 );
and ( n48464 , n37637 , n35150 );
or ( n48465 , n35160 , n18558 );
or ( n48466 , n37644 , n35166 );
or ( n48467 , n35158 , n37646 );
nand ( n48468 , n48465 , n48466 , n48467 );
nor ( n48469 , n48464 , n48468 );
nand ( n48470 , n48463 , n48469 );
buf ( n48471 , n48470 );
buf ( n48472 , n382067 );
buf ( n48473 , n22404 );
not ( n48474 , n386863 );
or ( n48475 , n48474 , n22473 );
nand ( n48476 , n48475 , n383474 );
not ( n48477 , n386870 );
nand ( n48478 , n48476 , n48477 );
not ( n48479 , n48477 );
nand ( n48480 , n48479 , n37068 , n48474 );
not ( n48481 , RI15b641d0_1281);
not ( n48482 , n44548 );
or ( n48483 , n48481 , n48482 );
not ( n48484 , n34814 );
not ( n48485 , n386978 );
not ( n48486 , n48485 );
or ( n48487 , n48484 , n48486 );
nand ( n48488 , n48487 , n34823 );
and ( n48489 , n48488 , RI15b623d0_1217);
or ( n48490 , n34833 , n44544 , RI15b641d0_1281);
or ( n48491 , n34826 , n48485 , RI15b623d0_1217);
nand ( n48492 , n48490 , n48491 );
nor ( n48493 , n48489 , n48492 );
nand ( n48494 , n48483 , n48493 );
nand ( n48495 , n48494 , n19201 );
and ( n48496 , n22423 , RI15b641d0_1281);
and ( n48497 , n19599 , RI15b632d0_1249);
nor ( n48498 , n48496 , n48497 , n19513 );
nand ( n48499 , n48478 , n48480 , n48495 , n48498 );
buf ( n48500 , n48499 );
buf ( n48501 , RI15b5e2a8_1078);
buf ( n48502 , n32676 );
buf ( n48503 , n18226 );
not ( n48504 , n386219 );
not ( n48505 , n48504 );
nor ( n48506 , n40361 , n40362 );
not ( n48507 , n48506 );
or ( n48508 , n48505 , n48507 );
or ( n48509 , n48506 , n48504 );
nand ( n48510 , n48508 , n48509 );
buf ( n48511 , n39975 );
not ( n48512 , n48511 );
and ( n48513 , n48510 , n48512 );
nor ( n48514 , n40370 , n385870 );
buf ( n48515 , n48514 );
not ( n48516 , n48515 );
not ( n48517 , n385912 );
not ( n48518 , n48517 );
and ( n48519 , n48516 , n48518 );
and ( n48520 , n48515 , n48517 );
nor ( n48521 , n48519 , n48520 );
not ( n48522 , n386020 );
or ( n48523 , n48521 , n48522 );
or ( n48524 , n386457 , n386465 );
nand ( n48525 , n48524 , n386466 );
and ( n48526 , n48525 , n386500 );
buf ( n48527 , n41302 );
and ( n48528 , n48527 , RI15b4bbd0_449);
nor ( n48529 , n48526 , n48528 );
nand ( n48530 , n48523 , n48529 );
nor ( n48531 , n48513 , n48530 );
buf ( n48532 , n19862 );
or ( n48533 , n20638 , n48532 );
nand ( n48534 , n48533 , n34798 );
and ( n48535 , n48534 , RI15b4acd0_417);
not ( n48536 , n48532 );
or ( n48537 , n34801 , n48536 , RI15b4acd0_417);
or ( n48538 , n19868 , n22216 );
nand ( n48539 , n48537 , n48538 );
nor ( n48540 , n48535 , n48539 );
nand ( n48541 , n48531 , n48540 );
buf ( n48542 , n48541 );
or ( n48543 , n383180 , n36394 );
not ( n48544 , n36410 );
and ( n48545 , n48544 , RI15b592f8_908);
or ( n48546 , n383184 , n36400 );
or ( n48547 , n383189 , n36416 );
or ( n48548 , n36408 , n383192 );
nand ( n48549 , n48546 , n48547 , n48548 );
nor ( n48550 , n48545 , n48549 );
nand ( n48551 , n48543 , n48550 );
buf ( n48552 , n48551 );
buf ( n48553 , n20665 );
buf ( n48554 , n22005 );
buf ( n48555 , n22716 );
not ( n48556 , RI15b55ba8_790);
not ( n48557 , n380000 );
or ( n48558 , n48556 , n48557 );
and ( n48559 , n381636 , RI15b4e8d0_545);
and ( n48560 , n381639 , RI15b4e510_537);
nor ( n48561 , n48559 , n48560 );
and ( n48562 , n381643 , RI15b4ec90_553);
and ( n48563 , n381651 , RI15b4d9d0_513);
and ( n48564 , n382803 , RI15b4fb90_585);
nor ( n48565 , n48563 , n48564 );
and ( n48566 , n381661 , RI15b4f7d0_577);
and ( n48567 , n381663 , RI15b4f050_561);
nor ( n48568 , n48566 , n48567 );
and ( n48569 , n381667 , RI15b4d250_497);
and ( n48570 , n381669 , RI15b4d610_505);
nor ( n48571 , n48569 , n48570 );
and ( n48572 , n381672 , RI15b4dd90_521);
and ( n48573 , n381674 , RI15b4f410_569);
nor ( n48574 , n48572 , n48573 );
nand ( n48575 , n48565 , n48568 , n48571 , n48574 );
and ( n48576 , n386643 , n48575 );
and ( n48577 , n381680 , RI15b4c710_473);
nor ( n48578 , n48562 , n48576 , n48577 );
and ( n48579 , n381684 , RI15b4c350_465);
and ( n48580 , n381686 , RI15b4e150_529);
nor ( n48581 , n48579 , n48580 );
and ( n48582 , n381689 , RI15b4cad0_481);
and ( n48583 , n381691 , RI15b4ce90_489);
nor ( n48584 , n48582 , n48583 );
nand ( n48585 , n48561 , n48578 , n48581 , n48584 );
and ( n48586 , n48585 , n38347 );
not ( n48587 , RI15b55ba8_790);
not ( n48588 , n379958 );
not ( n48589 , n48588 );
or ( n48590 , n48587 , n48589 );
or ( n48591 , n48588 , RI15b55ba8_790);
nand ( n48592 , n48590 , n48591 );
and ( n48593 , n379949 , n48592 );
nor ( n48594 , n48586 , n48593 );
nand ( n48595 , n48558 , n48594 );
buf ( n48596 , n48595 );
buf ( n48597 , n18226 );
buf ( n48598 , RI15b470d0_289);
buf ( n48599 , n381006 );
not ( n48600 , n41340 );
not ( n48601 , n48600 );
nor ( n48602 , n48601 , RI15b619f8_1196);
nor ( n48603 , n46076 , n48602 );
not ( n48604 , RI15b61a70_1197);
or ( n48605 , n48603 , n48604 );
not ( n48606 , n46080 );
and ( n48607 , n48606 , n48604 , RI15b619f8_1196);
or ( n48608 , n45422 , n44459 );
or ( n48609 , n380493 , n31052 );
nand ( n48610 , n384906 , n44038 );
nand ( n48611 , n48608 , n48609 , n48610 );
nor ( n48612 , n48607 , n48611 );
nand ( n48613 , n48605 , n48612 );
buf ( n48614 , n48613 );
buf ( n48615 , n20663 );
or ( n48616 , n386705 , n36242 );
and ( n48617 , n386716 , n43075 );
not ( n48618 , RI15b4d430_501);
or ( n48619 , n36250 , n48618 );
or ( n48620 , n37443 , n36254 );
or ( n48621 , n36248 , n386738 );
nand ( n48622 , n48619 , n48620 , n48621 );
nor ( n48623 , n48617 , n48622 );
nand ( n48624 , n48616 , n48623 );
buf ( n48625 , n48624 );
buf ( n48626 , n22653 );
buf ( n48627 , n21800 );
buf ( n48628 , n40995 );
not ( n48629 , n48628 );
or ( n48630 , n48629 , n41015 );
nand ( n48631 , n48630 , n41032 );
not ( n48632 , n35098 );
nand ( n48633 , n48631 , n48632 );
nor ( n48634 , n48628 , n48632 );
nand ( n48635 , n41578 , n48634 );
nand ( n48636 , n41582 , RI15b46158_256);
and ( n48637 , n35459 , n22283 );
and ( n48638 , n35461 , RI15b65940_1331);
nor ( n48639 , n48637 , n48638 );
nand ( n48640 , n48633 , n48635 , n48636 , n48639 );
buf ( n48641 , n48640 );
buf ( n48642 , n384218 );
buf ( n48643 , n31719 );
not ( n48644 , n38974 );
not ( n48645 , n383547 );
and ( n48646 , n48644 , n48645 );
nor ( n48647 , n48646 , n383577 );
or ( n48648 , n48647 , n44296 );
and ( n48649 , n383601 , RI15b5fc70_1133);
and ( n48650 , n383603 , n44297 );
and ( n48651 , n383607 , RI15b5f4f0_1117);
nor ( n48652 , n48649 , n48650 , n48651 );
nand ( n48653 , n48648 , n48652 );
buf ( n48654 , n48653 );
buf ( n48655 , n22653 );
buf ( n48656 , n383613 );
or ( n48657 , n386705 , n383845 );
and ( n48658 , n386716 , n383878 );
not ( n48659 , RI15b4f230_565);
or ( n48660 , n383903 , n48659 );
or ( n48661 , n44306 , n383911 );
or ( n48662 , n383895 , n386738 );
nand ( n48663 , n48660 , n48661 , n48662 );
nor ( n48664 , n48658 , n48663 );
nand ( n48665 , n48657 , n48664 );
buf ( n48666 , n48665 );
buf ( n48667 , n22714 );
not ( n48668 , RI15b543c0_739);
nand ( n48669 , n21946 , n385161 , n21750 );
not ( n48670 , n48669 );
or ( n48671 , n48668 , n48670 );
nand ( n48672 , n48671 , n18164 );
buf ( n48673 , n48672 );
buf ( n48674 , n382537 );
buf ( n48675 , n22343 );
not ( n48676 , n33220 );
not ( n48677 , n382912 );
or ( n48678 , n48676 , n48677 );
and ( n48679 , n382931 , n33226 );
or ( n48680 , n33237 , n18523 );
or ( n48681 , n35163 , n33241 );
or ( n48682 , n33235 , n382967 );
nand ( n48683 , n48680 , n48681 , n48682 );
nor ( n48684 , n48679 , n48683 );
nand ( n48685 , n48678 , n48684 );
buf ( n48686 , n48685 );
buf ( n48687 , n383174 );
buf ( n48688 , n381707 );
buf ( n48689 , n22406 );
or ( n48690 , n22372 , n386534 , n22395 );
nand ( n48691 , n48690 , RI15b47fd0_321);
nand ( n48692 , n48691 , n20621 );
buf ( n48693 , n48692 );
buf ( n48694 , n33382 );
buf ( n48695 , n32160 );
not ( n48696 , n43396 );
not ( n48697 , n384122 );
or ( n48698 , n48696 , n48697 );
and ( n48699 , n384164 , n386718 );
or ( n48700 , n386727 , n20864 );
or ( n48701 , n33131 , n386735 );
or ( n48702 , n386725 , n384193 );
nand ( n48703 , n48700 , n48701 , n48702 );
nor ( n48704 , n48699 , n48703 );
nand ( n48705 , n48698 , n48704 );
buf ( n48706 , n48705 );
buf ( n48707 , RI15b5ddf8_1068);
buf ( n48708 , n382073 );
not ( n48709 , RI15b61d40_1203);
or ( n48710 , n384021 , n48709 );
or ( n48711 , n18992 , n386747 );
and ( n48712 , n384027 , RI15b61d40_1203);
not ( n48713 , n384027 );
not ( n48714 , RI15b61d40_1203);
and ( n48715 , n48713 , n48714 );
nor ( n48716 , n48712 , n48715 );
or ( n48717 , n48716 , n384024 );
nand ( n48718 , n48710 , n48711 , n48717 );
buf ( n48719 , n48718 );
buf ( n48720 , n19653 );
buf ( n48721 , n386760 );
buf ( n48722 , n381490 );
buf ( n48723 , n384218 );
or ( n48724 , n32430 , n381409 );
and ( n48725 , n45712 , RI15b54ca8_758);
and ( n48726 , n48585 , n32437 );
or ( n48727 , n45708 , n381442 , RI15b54ca8_758);
or ( n48728 , n383009 , RI15b54c30_757);
nand ( n48729 , n48727 , n48728 );
and ( n48730 , n32439 , n48729 );
nor ( n48731 , n48725 , n48726 , n48730 );
and ( n48732 , n381418 , n48731 );
nand ( n48733 , n48724 , n48732 );
buf ( n48734 , n48733 );
buf ( n48735 , n32271 );
or ( n48736 , n383180 , n32062 );
not ( n48737 , n32081 );
and ( n48738 , n48737 , RI15b5a1f8_940);
or ( n48739 , n383184 , n32069 );
not ( n48740 , n32086 );
and ( n48741 , n48740 , n41701 );
and ( n48742 , n40019 , n32084 );
nor ( n48743 , n48741 , n48742 );
nand ( n48744 , n48739 , n48743 );
nor ( n48745 , n48738 , n48744 );
nand ( n48746 , n48736 , n48745 );
buf ( n48747 , n48746 );
or ( n48748 , n48071 , n22582 );
and ( n48749 , n35734 , RI15b4fd70_589);
and ( n48750 , n35759 , RI15b4f230_565);
and ( n48751 , n381650 , RI15b4df70_525);
and ( n48752 , n48135 , RI15b4dbb0_517);
and ( n48753 , n380115 , RI15b4c530_469);
nor ( n48754 , n48751 , n48752 , n48753 );
and ( n48755 , n382788 , RI15b4d070_493);
and ( n48756 , n382780 , RI15b4d7f0_509);
nor ( n48757 , n48755 , n48756 );
and ( n48758 , n382813 , RI15b4c8f0_477);
and ( n48759 , n379877 , RI15b4ccb0_485);
nor ( n48760 , n48758 , n48759 );
nand ( n48761 , n35739 , RI15b4d430_501);
and ( n48762 , n48754 , n48757 , n48760 , n48761 );
and ( n48763 , n382806 , RI15b4eab0_549);
and ( n48764 , n380061 , RI15b4ee70_557);
and ( n48765 , n47680 , RI15b4e6f0_541);
nor ( n48766 , n48763 , n48764 , n48765 );
nand ( n48767 , n35748 , RI15b4e330_533);
and ( n48768 , n48762 , n48766 , n48767 );
not ( n48769 , n386643 );
nor ( n48770 , n48768 , n48769 );
nor ( n48771 , n48749 , n48750 , n48770 );
and ( n48772 , n35754 , RI15b4f5f0_573);
and ( n48773 , n35756 , RI15b4f9b0_581);
nor ( n48774 , n48772 , n48773 );
nand ( n48775 , n48771 , n48774 );
and ( n48776 , n48775 , n38347 );
or ( n48777 , n48069 , n22580 , RI15b56148_802);
or ( n48778 , n22582 , RI15b560d0_801);
nand ( n48779 , n48777 , n48778 );
and ( n48780 , n48779 , n379949 );
nor ( n48781 , n48776 , n48780 );
nand ( n48782 , n48748 , n48781 );
buf ( n48783 , n48782 );
buf ( n48784 , RI15b476e8_302);
buf ( n48785 , n381872 );
not ( n48786 , n47644 );
not ( n48787 , n33400 );
or ( n48788 , n48786 , n48787 );
and ( n48789 , n33415 , n47649 );
or ( n48790 , n47658 , n18499 );
or ( n48791 , n36293 , n47663 );
or ( n48792 , n47656 , n33443 );
nand ( n48793 , n48790 , n48791 , n48792 );
nor ( n48794 , n48789 , n48793 );
nand ( n48795 , n48788 , n48794 );
buf ( n48796 , n48795 );
buf ( n48797 , n43349 );
buf ( n48798 , n22479 );
buf ( n48799 , n381707 );
buf ( n48800 , n22655 );
nand ( n48801 , n41173 , n382958 );
nand ( n48802 , n384918 , RI15b5f1a8_1110);
nand ( n48803 , n37773 , RI15b60eb8_1172);
nand ( n48804 , n41335 , n48801 , n48802 , n48803 );
buf ( n48805 , n48804 );
or ( n48806 , n31006 , n40468 );
and ( n48807 , n31016 , n40470 );
or ( n48808 , n40480 , n20997 );
or ( n48809 , n34893 , n40485 );
or ( n48810 , n40478 , n31024 );
nand ( n48811 , n48808 , n48809 , n48810 );
nor ( n48812 , n48807 , n48811 );
nand ( n48813 , n48806 , n48812 );
buf ( n48814 , n48813 );
or ( n48815 , n383180 , n381569 );
not ( n48816 , n381609 );
and ( n48817 , n48816 , RI15b58f38_900);
or ( n48818 , n383184 , n381598 );
or ( n48819 , n383189 , n381619 );
or ( n48820 , n381607 , n383192 );
nand ( n48821 , n48818 , n48819 , n48820 );
nor ( n48822 , n48817 , n48821 );
nand ( n48823 , n48815 , n48822 );
buf ( n48824 , n48823 );
buf ( n48825 , n384203 );
not ( n48826 , RI15b55f68_798);
not ( n48827 , n380000 );
or ( n48828 , n48826 , n48827 );
and ( n48829 , n43691 , n381696 );
not ( n48830 , RI15b55f68_798);
not ( n48831 , n379969 );
not ( n48832 , n48831 );
or ( n48833 , n48830 , n48832 );
or ( n48834 , n48831 , RI15b55f68_798);
nand ( n48835 , n48833 , n48834 );
and ( n48836 , n48835 , n379949 );
nor ( n48837 , n48829 , n48836 );
nand ( n48838 , n48828 , n48837 );
buf ( n48839 , n48838 );
buf ( n48840 , n22404 );
buf ( n48841 , n17499 );
buf ( n48842 , n22788 );
not ( n48843 , RI15b53a60_719);
not ( n48844 , n383170 );
or ( n48845 , n48843 , n48844 );
nor ( n48846 , n40057 , n40066 );
not ( n48847 , n48846 );
not ( n48848 , n33453 );
or ( n48849 , n48847 , n48848 );
nand ( n48850 , n48849 , n33465 );
not ( n48851 , n383015 );
not ( n48852 , n40060 );
or ( n48853 , n48851 , n48852 );
nand ( n48854 , n48853 , RI15b55770_781);
and ( n48855 , n48854 , n382651 );
not ( n48856 , n48854 );
and ( n48857 , n48856 , RI15b54ff0_765);
nor ( n48858 , n48855 , n48857 );
and ( n48859 , n48850 , n48858 );
nor ( n48860 , n48846 , n48858 );
and ( n48861 , n33476 , n48860 );
and ( n48862 , n383147 , RI15b532e0_703);
nor ( n48863 , n48859 , n48861 , n48862 );
nand ( n48864 , n48845 , n48863 );
buf ( n48865 , n48864 );
not ( n48866 , n35145 );
not ( n48867 , n380703 );
or ( n48868 , n48866 , n48867 );
and ( n48869 , n380719 , n35150 );
or ( n48870 , n35160 , n19021 );
not ( n48871 , n37541 );
or ( n48872 , n48871 , n35166 );
or ( n48873 , n35158 , n380790 );
nand ( n48874 , n48870 , n48872 , n48873 );
nor ( n48875 , n48869 , n48874 );
nand ( n48876 , n48868 , n48875 );
buf ( n48877 , n48876 );
buf ( n48878 , n379847 );
or ( n48879 , n36714 , n20519 );
or ( n48880 , n39256 , n20429 );
or ( n48881 , RI15b449e8_206 , n22298 );
or ( n48882 , RI15b43ae8_174 , n36114 );
nand ( n48883 , n48880 , n48881 , n48882 );
not ( n48884 , n48883 );
nand ( n48885 , n48879 , n48884 );
buf ( n48886 , n48885 );
buf ( n48887 , n380906 );
buf ( n48888 , n381081 );
buf ( n48889 , n379844 );
buf ( n48890 , n33250 );
not ( n48891 , RI15b538f8_716);
not ( n48892 , n32244 );
or ( n48893 , n48891 , n48892 );
and ( n48894 , n32247 , RI15b64ef0_1309);
and ( n48895 , n32249 , RI15b5fd60_1135);
nor ( n48896 , n48894 , n48895 );
nand ( n48897 , n48893 , n48896 );
buf ( n48898 , n48897 );
buf ( n48899 , n22716 );
and ( n48900 , n37130 , n19995 );
not ( n48901 , n37130 );
and ( n48902 , n48901 , RI15b49fb0_389);
nor ( n48903 , n48900 , n48902 );
nand ( n48904 , n48903 , n37113 );
and ( n48905 , n381055 , RI15b49fb0_389);
and ( n48906 , n37259 , n37287 );
buf ( n48907 , n44855 );
not ( n48908 , n48907 );
not ( n48909 , n37288 );
nor ( n48910 , n48906 , n48908 , n48909 );
buf ( n48911 , n44859 );
and ( n48912 , n48910 , n48911 );
nor ( n48913 , n48905 , n48912 );
nand ( n48914 , n48904 , n48913 );
buf ( n48915 , n48914 );
buf ( n48916 , n382052 );
buf ( n48917 , n31719 );
buf ( n48918 , n21800 );
not ( n48919 , RI15b60120_1143);
not ( n48920 , n383601 );
or ( n48921 , n48919 , n48920 );
buf ( n48922 , n32318 );
or ( n48923 , n48922 , n33577 );
nand ( n48924 , n48923 , n33584 );
and ( n48925 , n48924 , n32327 );
and ( n48926 , n383607 , RI15b5eb18_1096);
not ( n48927 , n32327 );
nand ( n48928 , n48927 , n48922 );
nor ( n48929 , n48928 , n33588 );
nor ( n48930 , n48925 , n48926 , n48929 );
nand ( n48931 , n48921 , n48930 );
buf ( n48932 , n48931 );
buf ( n48933 , n20663 );
buf ( n48934 , n384996 );
buf ( n48935 , n33250 );
nand ( n48936 , n33109 , n383866 );
or ( n48937 , n31149 , n48936 );
nand ( n48938 , n385004 , n384056 );
not ( n48939 , n48938 );
and ( n48940 , n31161 , n48939 );
and ( n48941 , n48938 , n48936 , n383882 );
nor ( n48942 , n48941 , n21764 );
nor ( n48943 , n385012 , n383832 );
or ( n48944 , n48942 , n48943 );
nand ( n48945 , n48944 , n18154 );
or ( n48946 , n385016 , n383886 );
nand ( n48947 , n48945 , n48946 );
and ( n48948 , n48947 , n383901 );
not ( n48949 , RI15b4ed80_555);
or ( n48950 , n48948 , n48949 );
not ( n48951 , n48946 );
nor ( n48952 , n48943 , n48951 );
or ( n48953 , n48942 , n48952 );
or ( n48954 , n31179 , n48953 );
or ( n48955 , n48946 , n31184 );
nand ( n48956 , n48950 , n48954 , n48955 );
nor ( n48957 , n48940 , n48956 );
nand ( n48958 , n48937 , n48957 );
buf ( n48959 , n48958 );
or ( n48960 , n381015 , n22028 );
nand ( n48961 , n381017 , RI15b53808_714);
nand ( n48962 , n48960 , n48961 );
buf ( n48963 , n48962 );
buf ( n48964 , n31033 );
buf ( n48965 , n32981 );
buf ( n48966 , n22479 );
buf ( n48967 , n381081 );
buf ( n48968 , n44504 );
not ( n48969 , n48968 );
nand ( n48970 , n35358 , RI15b48e58_352);
not ( n48971 , n48970 );
nand ( n48972 , n48971 , RI15b48ed0_353);
nand ( n48973 , RI15b48f48_354 , RI15b48fc0_355);
nor ( n48974 , n48972 , n48973 );
and ( n48975 , n48974 , RI15b49038_356);
nand ( n48976 , n48975 , RI15b490b0_357);
not ( n48977 , n48976 );
or ( n48978 , n48969 , n48977 );
buf ( n48979 , n35187 );
buf ( n48980 , n48979 );
not ( n48981 , n48980 );
nand ( n48982 , n48978 , n48981 );
nand ( n48983 , n48982 , RI15b491a0_359);
nand ( n48984 , n35002 , RI15b49128_358);
nor ( n48985 , n48976 , n48984 );
nor ( n48986 , n35002 , RI15b49128_358);
or ( n48987 , n48985 , n48986 );
buf ( n48988 , n35363 );
buf ( n48989 , n48988 );
not ( n48990 , n48989 );
buf ( n48991 , n48990 );
not ( n48992 , n48991 );
nand ( n48993 , n48987 , n48992 );
and ( n48994 , n37321 , n37355 );
not ( n48995 , n48907 );
nor ( n48996 , n48994 , n37356 , n48995 );
not ( n48997 , n35534 );
buf ( n48998 , n48997 );
and ( n48999 , n48996 , n48998 );
and ( n49000 , n35335 , RI15b66570_1357);
nor ( n49001 , n48999 , n49000 );
nand ( n49002 , n48983 , n48993 , n46625 , n49001 );
buf ( n49003 , n49002 );
not ( n49004 , n48504 );
nand ( n49005 , n49004 , n48506 );
not ( n49006 , n386215 );
and ( n49007 , n49005 , n49006 );
not ( n49008 , n49005 );
and ( n49009 , n49008 , n386215 );
nor ( n49010 , n49007 , n49009 );
not ( n49011 , n48511 );
and ( n49012 , n49010 , n49011 );
and ( n49013 , n48514 , n385912 );
not ( n49014 , n49013 );
not ( n49015 , n385858 );
and ( n49016 , n49014 , n49015 );
and ( n49017 , n49013 , n385858 );
nor ( n49018 , n49016 , n49017 );
not ( n49019 , n386020 );
or ( n49020 , n49018 , n49019 );
and ( n49021 , n386466 , n386473 );
nor ( n49022 , n49021 , n386474 );
not ( n49023 , n49022 );
and ( n49024 , n49023 , n386500 );
and ( n49025 , n39988 , RI15b4bc48_450);
nor ( n49026 , n49024 , n49025 );
nand ( n49027 , n49020 , n49026 );
nor ( n49028 , n49012 , n49027 );
not ( n49029 , n41308 );
buf ( n49030 , n49029 );
and ( n49031 , n49030 , n386473 );
not ( n49032 , RI15b445b0_197);
or ( n49033 , n386541 , n49032 );
or ( n49034 , n385858 , n386550 );
or ( n49035 , n49006 , n386557 );
nand ( n49036 , n49033 , n49034 , n49035 );
nor ( n49037 , n49031 , n49036 );
nand ( n49038 , n49028 , n49037 );
buf ( n49039 , n49038 );
buf ( n49040 , n382065 );
buf ( n49041 , n380906 );
buf ( n49042 , n381872 );
buf ( n49043 , n33382 );
buf ( n49044 , n382073 );
or ( n49045 , n36238 , n385005 );
not ( n49046 , n385019 );
and ( n49047 , n49046 , RI15b4e150_529);
or ( n49048 , n385023 , n32710 );
or ( n49049 , n385002 , n383802 );
or ( n49050 , n385017 , n42402 );
nand ( n49051 , n49048 , n49049 , n49050 );
nor ( n49052 , n49047 , n49051 );
nand ( n49053 , n49045 , n49052 );
buf ( n49054 , n49053 );
buf ( n49055 , n379403 );
or ( n49056 , n31091 , n35514 );
and ( n49057 , n35507 , n42028 );
not ( n49058 , n35509 );
or ( n49059 , n49058 , n384904 , n40016 );
or ( n49060 , n35512 , RI15b60d50_1169);
nand ( n49061 , n49059 , n49060 );
nor ( n49062 , n49057 , n49061 );
nand ( n49063 , n49056 , n49062 );
buf ( n49064 , n49063 );
buf ( n49065 , n20663 );
or ( n49066 , n30908 , n385210 );
nand ( n49067 , n49066 , RI15b4a280_395);
not ( n49068 , n39299 );
buf ( n49069 , n386011 );
nand ( n49070 , n49068 , n49069 );
nand ( n49071 , n49067 , n39308 , n49070 );
buf ( n49072 , n49071 );
buf ( n49073 , n32676 );
not ( n49074 , RI15b53628_710);
not ( n49075 , n32244 );
or ( n49076 , n49074 , n49075 );
and ( n49077 , n32247 , RI15b64c20_1303);
and ( n49078 , n32249 , RI15b5fa90_1129);
nor ( n49079 , n49077 , n49078 );
nand ( n49080 , n49076 , n49079 );
buf ( n49081 , n49080 );
buf ( n49082 , n382067 );
buf ( n49083 , n22740 );
buf ( n49084 , n22404 );
buf ( n49085 , n381021 );
buf ( n49086 , n381490 );
nand ( n49087 , RI15b49128_358 , RI15b491a0_359);
nor ( n49088 , n48976 , n49087 );
not ( n49089 , n49088 );
and ( n49090 , n49089 , n35006 );
not ( n49091 , n49089 );
and ( n49092 , n49091 , RI15b49218_360);
nor ( n49093 , n49090 , n49092 );
not ( n49094 , n48992 );
not ( n49095 , n49094 );
nand ( n49096 , n49093 , n49095 );
buf ( n49097 , n48980 );
and ( n49098 , n49097 , RI15b49218_360);
not ( n49099 , n386554 );
or ( n49100 , n46787 , n49099 );
or ( n49101 , n380965 , n386547 );
not ( n49102 , n381968 );
not ( n49103 , n382031 );
or ( n49104 , n49102 , n49103 );
or ( n49105 , n382031 , n381968 );
nand ( n49106 , n49104 , n49105 );
and ( n49107 , n49106 , n35461 );
and ( n49108 , n35459 , RI15b65e68_1342);
nor ( n49109 , n49107 , n49108 );
nand ( n49110 , n49100 , n49101 , n49109 );
nor ( n49111 , n49098 , n49110 );
nand ( n49112 , n49096 , n49111 );
buf ( n49113 , n49112 );
and ( n49114 , n38047 , RI15b53790_713);
and ( n49115 , n38049 , RI15b65c88_1338);
nor ( n49116 , n49114 , n49115 );
not ( n49117 , n49116 );
buf ( n49118 , n49117 );
buf ( n49119 , n381081 );
buf ( n49120 , n31033 );
or ( n49121 , n31771 , n18238 );
not ( n49122 , n31784 );
and ( n49123 , n49122 , n19377 );
and ( n49124 , n32386 , n380796 );
and ( n49125 , n31778 , n19403 );
nor ( n49126 , n49123 , n49124 , n49125 );
nand ( n49127 , n49121 , n19517 , n49126 );
buf ( n49128 , n49127 );
buf ( n49129 , n386762 );
not ( n49130 , RI15b52728_678);
not ( n49131 , n32397 );
or ( n49132 , n49130 , n49131 );
buf ( n49133 , n383121 );
or ( n49134 , n49133 , n36342 );
nand ( n49135 , n49134 , n381450 );
and ( n49136 , n49135 , n383128 );
not ( n49137 , n49133 );
nor ( n49138 , n49137 , n383128 );
and ( n49139 , n49138 , n381461 );
nor ( n49140 , n49136 , n49139 , n35778 );
nand ( n49141 , n49132 , n49140 );
buf ( n49142 , n49141 );
buf ( n49143 , n383174 );
buf ( n49144 , n32981 );
buf ( n49145 , n383613 );
or ( n49146 , n31006 , n48936 );
and ( n49147 , n31016 , n48939 );
or ( n49148 , n48948 , n20990 );
or ( n49149 , n33612 , n48953 );
or ( n49150 , n48946 , n31024 );
nand ( n49151 , n49148 , n49149 , n49150 );
nor ( n49152 , n49147 , n49151 );
nand ( n49153 , n49146 , n49152 );
buf ( n49154 , n49153 );
buf ( n49155 , n33250 );
not ( n49156 , RI15b600a8_1142);
not ( n49157 , n383601 );
or ( n49158 , n49156 , n49157 );
not ( n49159 , n32308 );
or ( n49160 , n49159 , n33577 );
nand ( n49161 , n49160 , n33584 );
not ( n49162 , n32317 );
and ( n49163 , n49161 , n49162 );
not ( n49164 , n49159 );
nor ( n49165 , n49164 , n49162 );
and ( n49166 , n49165 , n40781 );
and ( n49167 , n383607 , RI15b5eaa0_1095);
nor ( n49168 , n49163 , n49166 , n49167 );
nand ( n49169 , n49158 , n49168 );
buf ( n49170 , n49169 );
not ( n49171 , n37773 );
not ( n49172 , n33574 );
or ( n49173 , n49171 , n49172 );
nand ( n49174 , n49173 , n37780 );
buf ( n49175 , n33550 );
not ( n49176 , n49175 );
nand ( n49177 , n49174 , n49176 );
not ( n49178 , n33574 );
nand ( n49179 , n49175 , n49178 , n384934 );
and ( n49180 , n384918 , RI15b5ede8_1102);
nor ( n49181 , n49180 , n44468 );
nand ( n49182 , n49177 , n49179 , n49181 );
buf ( n49183 , n49182 );
buf ( n49184 , n22406 );
buf ( n49185 , n380203 );
or ( n49186 , n385163 , n21020 );
and ( n49187 , n36472 , n21615 );
and ( n49188 , n385177 , n46361 );
nor ( n49189 , n49187 , n49188 );
and ( n49190 , n32368 , n46349 );
nor ( n49191 , n49190 , n46377 );
nand ( n49192 , n49186 , n49189 , n49191 );
buf ( n49193 , n49192 );
buf ( n49194 , n22655 );
buf ( n49195 , n18226 );
not ( n49196 , n47542 );
not ( n49197 , n384122 );
or ( n49198 , n49196 , n49197 );
and ( n49199 , n384164 , n35625 );
or ( n49200 , n35635 , n20881 );
or ( n49201 , n384187 , n35640 );
or ( n49202 , n35633 , n384193 );
nand ( n49203 , n49200 , n49201 , n49202 );
nor ( n49204 , n49199 , n49203 );
nand ( n49205 , n49198 , n49204 );
buf ( n49206 , n49205 );
not ( n49207 , RI15b5f7c0_1123);
not ( n49208 , n383601 );
or ( n49209 , n49207 , n49208 );
and ( n49210 , n383505 , RI15b60d50_1169);
and ( n49211 , n383607 , RI15b5f040_1107);
nor ( n49212 , n49210 , n49211 );
nand ( n49213 , n49209 , n49212 );
buf ( n49214 , n49213 );
buf ( n49215 , n386563 );
buf ( n49216 , n19653 );
buf ( n49217 , n22716 );
not ( n49218 , RI15b45e88_250);
not ( n49219 , n382527 );
or ( n49220 , n49218 , n49219 );
or ( n49221 , n36998 , RI15b47ee0_319);
nand ( n49222 , n49220 , n49221 );
buf ( n49223 , n49222 );
buf ( n49224 , n379403 );
buf ( n49225 , n30992 );
buf ( n49226 , n32676 );
not ( n49227 , n32680 );
not ( n49228 , n381507 );
or ( n49229 , n49227 , n49228 );
and ( n49230 , n381524 , n35222 );
or ( n49231 , n32692 , n18397 );
or ( n49232 , n36413 , n32699 );
or ( n49233 , n32690 , n381560 );
nand ( n49234 , n49231 , n49232 , n49233 );
nor ( n49235 , n49230 , n49234 );
nand ( n49236 , n49229 , n49235 );
buf ( n49237 , n49236 );
buf ( n49238 , n35649 );
and ( n49239 , n43295 , RI15b54618_744);
and ( n49240 , n35234 , n45855 );
nor ( n49241 , n49240 , RI15b3fab0_37);
nor ( n49242 , n49239 , n49241 );
not ( n49243 , n49242 );
buf ( n49244 , n49243 );
buf ( n49245 , n384218 );
buf ( n49246 , n22653 );
buf ( n49247 , n380942 );
nor ( n49248 , n48176 , n41015 );
or ( n49249 , n49248 , n41033 );
nand ( n49250 , n49249 , n48179 );
nor ( n49251 , n41036 , n48179 );
not ( n49252 , n49251 );
not ( n49253 , n48176 );
or ( n49254 , n49252 , n49253 );
and ( n49255 , n41017 , RI15b46680_267);
not ( n49256 , n49109 );
nor ( n49257 , n49255 , n49256 );
nand ( n49258 , n49254 , n49257 );
not ( n49259 , n49258 );
nand ( n49260 , n49250 , n49259 );
buf ( n49261 , n49260 );
buf ( n49262 , n32672 );
buf ( n49263 , n381021 );
not ( n49264 , n382526 );
or ( n49265 , n49264 , RI15b47e68_318);
and ( n49266 , n20492 , n382509 );
not ( n49267 , RI15b3fa38_36);
not ( n49268 , n385218 );
or ( n49269 , n49267 , n49268 );
and ( n49270 , RI15b3f9c0_35 , RI15b48318_328 , RI15b48390_329);
nor ( n49271 , n49270 , n43960 );
nand ( n49272 , n49269 , n49271 );
nor ( n49273 , n43516 , RI15b48390_329);
nor ( n49274 , n49266 , n49272 , n49273 );
nand ( n49275 , n49265 , n49274 );
buf ( n49276 , n49275 );
buf ( n49277 , n21800 );
buf ( n49278 , n19655 );
buf ( n49279 , n386563 );
buf ( n49280 , n22740 );
buf ( n49281 , n35651 );
buf ( n49282 , n22653 );
buf ( n49283 , n383613 );
or ( n49284 , n22315 , n35869 );
and ( n49285 , n22326 , n35872 );
not ( n49286 , RI15b40b90_73);
or ( n49287 , n35884 , n49286 );
or ( n49288 , n22334 , n35888 );
or ( n49289 , n35882 , n22336 );
nand ( n49290 , n49287 , n49288 , n49289 );
nor ( n49291 , n49285 , n49290 );
nand ( n49292 , n49284 , n49291 );
buf ( n49293 , n49292 );
or ( n49294 , n22102 , n35895 );
and ( n49295 , n22203 , n39462 );
not ( n49296 , RI15b40488_58);
or ( n49297 , n35911 , n49296 );
or ( n49298 , n22293 , n35917 );
or ( n49299 , n35909 , n22299 );
nand ( n49300 , n49297 , n49298 , n49299 );
nor ( n49301 , n49295 , n49300 );
nand ( n49302 , n49294 , n49301 );
buf ( n49303 , n49302 );
buf ( n49304 , n20665 );
not ( n49305 , n43220 );
nand ( n49306 , n49305 , n379785 );
not ( n49307 , n49306 );
not ( n49308 , n46287 );
or ( n49309 , n49307 , n49308 );
nand ( n49310 , n49309 , n43221 );
nor ( n49311 , n49305 , n43221 );
nand ( n49312 , n36580 , n49311 );
buf ( n49313 , n34589 );
and ( n49314 , n49313 , n34597 );
not ( n49315 , n49313 );
not ( n49316 , n34597 );
and ( n49317 , n49315 , n49316 );
nor ( n49318 , n49314 , n49317 );
and ( n49319 , n49318 , n46302 );
not ( n49320 , RI15b5e410_1081);
not ( n49321 , n34651 );
or ( n49322 , n49320 , n49321 );
or ( n49323 , n36518 , n379446 );
nand ( n49324 , n49322 , n49323 );
nor ( n49325 , n49319 , n49324 );
nand ( n49326 , n49310 , n49312 , n49325 );
buf ( n49327 , n49326 );
and ( n49328 , n385164 , RI15b50a90_617);
or ( n49329 , n40445 , n385170 );
or ( n49330 , n37877 , n381810 );
or ( n49331 , n381752 , n385178 );
nand ( n49332 , n49329 , n49330 , n49331 );
nor ( n49333 , n49328 , n49332 );
nand ( n49334 , n40455 , n49333 );
buf ( n49335 , n49334 );
buf ( n49336 , n381006 );
buf ( n49337 , n380203 );
buf ( n49338 , n32328 );
and ( n49339 , n49338 , n33579 );
nor ( n49340 , n49339 , n33585 );
or ( n49341 , n49340 , n32337 );
not ( n49342 , n32337 );
nor ( n49343 , n49338 , n49342 );
and ( n49344 , n49343 , n40781 );
and ( n49345 , n383607 , RI15b5eb90_1097);
nor ( n49346 , n49344 , n49345 );
nand ( n49347 , n383601 , RI15b60198_1144);
nand ( n49348 , n49341 , n49346 , n49347 );
buf ( n49349 , n49348 );
buf ( n49350 , n22714 );
or ( n49351 , n383814 , n48936 );
and ( n49352 , n383857 , n48939 );
not ( n49353 , RI15b4ed08_554);
or ( n49354 , n48948 , n49353 );
or ( n49355 , n383908 , n48953 );
or ( n49356 , n48946 , n383917 );
nand ( n49357 , n49354 , n49355 , n49356 );
nor ( n49358 , n49352 , n49357 );
nand ( n49359 , n49351 , n49358 );
buf ( n49360 , n49359 );
buf ( n49361 , n383613 );
buf ( n49362 , n387159 );
not ( n49363 , n43196 );
nor ( n49364 , n49363 , n43189 );
buf ( n49365 , n49364 );
or ( n49366 , n383814 , n33111 );
and ( n49367 , n383857 , n33117 );
or ( n49368 , n33128 , n21125 );
or ( n49369 , n41458 , n33134 );
or ( n49370 , n33126 , n383917 );
nand ( n49371 , n49368 , n49369 , n49370 );
nor ( n49372 , n49367 , n49371 );
nand ( n49373 , n49366 , n49372 );
buf ( n49374 , n49373 );
buf ( n49375 , n382065 );
buf ( n49376 , n31719 );
buf ( n49377 , n31979 );
or ( n49378 , n381015 , n22029 );
nand ( n49379 , n35525 , RI15b53880_715);
nand ( n49380 , n49378 , n49379 );
buf ( n49381 , n49380 );
buf ( n49382 , n31033 );
buf ( n49383 , n21800 );
not ( n49384 , n48982 );
or ( n49385 , n49384 , n35020 );
not ( n49386 , n48976 );
nor ( n49387 , n48990 , RI15b49128_358);
nand ( n49388 , n49386 , n49387 );
and ( n49389 , n386554 , n38445 );
and ( n49390 , n35335 , RI15b664f8_1356);
nor ( n49391 , n49389 , n49390 );
nand ( n49392 , n49388 , n49391 );
not ( n49393 , n44791 );
nor ( n49394 , n49392 , n49393 );
nand ( n49395 , n49385 , n49394 );
buf ( n49396 , n49395 );
buf ( n49397 , n22479 );
buf ( n49398 , n32981 );
buf ( n49399 , n22716 );
buf ( n49400 , n31033 );
buf ( n49401 , n381872 );
buf ( n49402 , n22655 );
or ( n49403 , n386515 , n386431 );
and ( n49404 , n386540 , RI15b43ea8_182);
not ( n49405 , n385807 );
or ( n49406 , n386550 , n49405 );
or ( n49407 , n386557 , n386055 );
nand ( n49408 , n49406 , n49407 );
nor ( n49409 , n49404 , n49408 );
nand ( n49410 , n49403 , n30897 , n49409 );
buf ( n49411 , n49410 );
buf ( n49412 , RI15b45f00_251);
buf ( n49413 , n382052 );
and ( n49414 , n19920 , n19730 );
nor ( n49415 , n49414 , n47493 );
or ( n49416 , n49415 , n19727 );
and ( n49417 , n32525 , RI15b4b2e8_430);
not ( n49418 , n19727 );
nor ( n49419 , n49418 , n19730 );
and ( n49420 , n22368 , n49419 );
nor ( n49421 , n49417 , n49420 );
not ( n49422 , n19956 );
or ( n49423 , n20502 , n49422 );
nand ( n49424 , n49423 , n380875 );
and ( n49425 , n49424 , RI15b494e8_366);
and ( n49426 , n32511 , n49422 , n19957 );
not ( n49427 , n20533 );
not ( n49428 , RI15b4b2e8_430);
and ( n49429 , n49427 , n49428 );
and ( n49430 , n20533 , RI15b4b2e8_430);
nor ( n49431 , n49429 , n49430 );
or ( n49432 , n22354 , n49431 );
or ( n49433 , n36782 , n37048 );
and ( n49434 , n22388 , RI15b4b2e8_430);
not ( n49435 , n20653 );
and ( n49436 , n49435 , RI15b4a3e8_398);
nor ( n49437 , n49434 , n49436 );
nand ( n49438 , n49432 , n49433 , n49437 );
nor ( n49439 , n49425 , n49426 , n49438 );
nand ( n49440 , n49416 , n49421 , n49439 );
buf ( n49441 , n49440 );
buf ( n49442 , n32676 );
buf ( n49443 , n381490 );
buf ( n49444 , n386957 );
or ( n49445 , n383482 , n49444 , RI15b61db8_1204);
buf ( n49446 , n386793 );
nand ( n49447 , n19628 , n49446 );
and ( n49448 , n383473 , n49447 );
or ( n49449 , n49448 , n386792 );
nand ( n49450 , n49445 , n49449 );
not ( n49451 , n49446 );
nand ( n49452 , n49451 , n386792 );
or ( n49453 , n383464 , n49452 );
and ( n49454 , n22471 , n42445 );
and ( n49455 , n22423 , RI15b63bb8_1268);
and ( n49456 , n19599 , RI15b62cb8_1236);
nor ( n49457 , n49454 , n49455 , n49456 );
nand ( n49458 , n49453 , n49457 );
not ( n49459 , n22450 );
not ( n49460 , n387020 );
not ( n49461 , RI15b63bb8_1268);
and ( n49462 , n49460 , n49461 );
and ( n49463 , n387020 , RI15b63bb8_1268);
nor ( n49464 , n49462 , n49463 );
nor ( n49465 , n49459 , n49464 );
nor ( n49466 , n49450 , n49458 , n49465 );
not ( n49467 , n49444 );
not ( n49468 , n383402 );
or ( n49469 , n49467 , n49468 );
nand ( n49470 , n49469 , n383408 );
nand ( n49471 , n49470 , RI15b61db8_1204);
nand ( n49472 , n383413 , RI15b63bb8_1268);
nand ( n49473 , n49466 , n49471 , n49472 );
buf ( n49474 , n49473 );
buf ( n49475 , n22005 );
buf ( n49476 , n33382 );
buf ( n49477 , n32981 );
and ( n49478 , n35118 , n42873 );
and ( n49479 , n20631 , RI15b462c0_259);
nor ( n49480 , n49478 , n49479 );
nor ( n49481 , n42867 , n34930 );
or ( n49482 , n35114 , n49481 );
nand ( n49483 , n49482 , n42870 );
nand ( n49484 , n385213 , RI15b478c8_306);
nand ( n49485 , n49480 , n49483 , n49484 );
buf ( n49486 , n49485 );
buf ( n49487 , n385195 );
buf ( n49488 , n22404 );
buf ( n49489 , n381081 );
not ( n49490 , n382158 );
not ( n49491 , n382057 );
or ( n49492 , n49490 , n49491 );
nand ( n49493 , n49492 , n382059 );
buf ( n49494 , n49493 );
buf ( n49495 , n22406 );
buf ( n49496 , n382067 );
buf ( n49497 , n379895 );
buf ( n49498 , n380906 );
buf ( n49499 , n379403 );
buf ( n49500 , n381490 );
buf ( n49501 , n32160 );
and ( n49502 , n36999 , RI15b481b0_325);
and ( n49503 , n37001 , RI15b45000_219);
nor ( n49504 , n49502 , n49503 );
not ( n49505 , n49504 );
buf ( n49506 , n49505 );
buf ( n49507 , n380903 );
buf ( n49508 , RI15b5e500_1083);
or ( n49509 , n380968 , n36306 );
and ( n49510 , n380986 , n36309 );
or ( n49511 , n36318 , n385457 );
or ( n49512 , n380994 , n36325 );
or ( n49513 , n36316 , n380996 );
nand ( n49514 , n49511 , n49512 , n49513 );
nor ( n49515 , n49510 , n49514 );
nand ( n49516 , n49509 , n49515 );
buf ( n49517 , n49516 );
buf ( n49518 , n384199 );
buf ( n49519 , n384218 );
buf ( n49520 , n379403 );
buf ( n49521 , n22005 );
and ( n49522 , n40674 , RI15b545a0_743);
not ( n49523 , n379396 );
and ( n49524 , n49523 , RI15b51468_638);
nor ( n49525 , n49522 , n49524 );
not ( n49526 , n49525 );
buf ( n49527 , n49526 );
not ( n49528 , n379507 );
not ( n49529 , n33759 );
or ( n49530 , n49528 , n49529 );
buf ( n49531 , n34270 );
or ( n49532 , n33766 , n49531 );
nand ( n49533 , n49530 , n49532 );
not ( n49534 , n49533 );
not ( n49535 , n33925 );
not ( n49536 , n49535 );
or ( n49537 , n49534 , n49536 );
not ( n49538 , n49531 );
or ( n49539 , n33955 , n49538 );
nor ( n49540 , n387019 , RI15b648d8_1296);
nand ( n49541 , n49539 , n49540 );
nand ( n49542 , n49537 , n49541 );
nand ( n49543 , n49542 , n379785 );
buf ( n49544 , n34307 );
and ( n49545 , n34309 , n49544 );
not ( n49546 , n34309 );
not ( n49547 , n49544 );
and ( n49548 , n49546 , n49547 );
nor ( n49549 , n49545 , n49548 );
and ( n49550 , n49549 , n22440 );
not ( n49551 , RI15b5da38_1060);
not ( n49552 , n379796 );
or ( n49553 , n49551 , n49552 );
or ( n49554 , n36518 , n379479 );
nand ( n49555 , n49553 , n49554 );
nor ( n49556 , n49550 , n49555 );
nand ( n49557 , n49543 , n49556 );
buf ( n49558 , n49557 );
buf ( n49559 , n385197 );
and ( n49560 , n22646 , RI15b452d0_225);
and ( n49561 , n22648 , RI15b51738_644);
nor ( n49562 , n49560 , n49561 );
not ( n49563 , n49562 );
buf ( n49564 , n49563 );
buf ( n49565 , n383498 );
buf ( n49566 , n379403 );
and ( n49567 , n21788 , RI15b569b8_820);
and ( n49568 , n21768 , n21835 );
buf ( n49569 , n21829 );
and ( n49570 , n49569 , n17529 );
not ( n49571 , n49569 );
and ( n49572 , n49571 , RI15b569b8_820);
nor ( n49573 , n49570 , n49572 );
and ( n49574 , n22704 , n49573 );
nor ( n49575 , n49567 , n49568 , n49574 );
nand ( n49576 , n37876 , n49575 );
buf ( n49577 , n49576 );
not ( n49578 , n22462 );
not ( n49579 , n45723 );
or ( n49580 , n49578 , n49579 );
nand ( n49581 , n49580 , n19201 );
nand ( n49582 , n49581 , RI15b584e8_878);
not ( n49583 , n19281 );
nand ( n49584 , n49582 , n382570 , n49583 );
buf ( n49585 , n49584 );
buf ( n49586 , n21800 );
or ( n49587 , n386705 , n385002 );
and ( n49588 , n386716 , n385006 );
not ( n49589 , RI15b4e330_533);
or ( n49590 , n385019 , n49589 );
or ( n49591 , n37443 , n385023 );
or ( n49592 , n385017 , n386738 );
nand ( n49593 , n49590 , n49591 , n49592 );
nor ( n49594 , n49588 , n49593 );
nand ( n49595 , n49587 , n49594 );
buf ( n49596 , n49595 );
buf ( n49597 , n19653 );
buf ( n49598 , n383613 );
buf ( n49599 , n31033 );
and ( n49600 , n33098 , RI15b60b70_1165);
buf ( n49601 , n49600 );
buf ( n49602 , n33382 );
buf ( n49603 , n382052 );
buf ( n49604 , n22402 );
buf ( n49605 , n381004 );
or ( n49606 , n31006 , n39691 );
and ( n49607 , n31016 , n39694 );
or ( n49608 , n39703 , n17716 );
or ( n49609 , n33612 , n39707 );
or ( n49610 , n39701 , n31024 );
nand ( n49611 , n49608 , n49609 , n49610 );
nor ( n49612 , n49607 , n49611 );
nand ( n49613 , n49606 , n49612 );
buf ( n49614 , n49613 );
not ( n49615 , n42635 );
or ( n49616 , n49615 , n39777 );
or ( n49617 , n38482 , n384021 );
and ( n49618 , n38481 , RI15b62628_1222);
not ( n49619 , n38481 );
and ( n49620 , n49619 , n38482 );
nor ( n49621 , n49618 , n49620 );
or ( n49622 , n384024 , n49621 );
nand ( n49623 , n49616 , n49617 , n49622 );
buf ( n49624 , n49623 );
buf ( n49625 , n22402 );
buf ( n49626 , n381490 );
nand ( n49627 , n49088 , RI15b49218_360);
and ( n49628 , n49627 , n35049 );
not ( n49629 , n49627 );
and ( n49630 , n49629 , RI15b49290_361);
nor ( n49631 , n49628 , n49630 );
not ( n49632 , n48992 );
not ( n49633 , n49632 );
nand ( n49634 , n49631 , n49633 );
and ( n49635 , n49097 , RI15b49290_361);
or ( n49636 , n37418 , n49099 );
or ( n49637 , n384945 , n386547 );
nand ( n49638 , n379820 , RI15b65ee0_1343);
nand ( n49639 , n49636 , n49637 , n49638 );
nor ( n49640 , n49635 , n49639 );
nand ( n49641 , n49634 , n49640 );
buf ( n49642 , n49641 );
buf ( n49643 , n381490 );
buf ( n49644 , n22653 );
or ( n49645 , n381015 , n22025 );
nand ( n49646 , n35525 , RI15b53718_712);
nand ( n49647 , n49645 , n49646 );
buf ( n49648 , n49647 );
nand ( n49649 , n44209 , n383143 );
nor ( n49650 , n49649 , n44217 );
not ( n49651 , n49650 );
nor ( n49652 , n44209 , n383152 );
or ( n49653 , n49652 , n38288 );
nand ( n49654 , n49653 , n44212 );
nand ( n49655 , n383170 , RI15b53f88_730);
nand ( n49656 , n383147 , RI15b52980_683);
nand ( n49657 , n49651 , n49654 , n49655 , n49656 );
buf ( n49658 , n49657 );
buf ( n49659 , n380903 );
buf ( n49660 , n379847 );
buf ( n49661 , n32672 );
not ( n49662 , n382976 );
not ( n49663 , n33400 );
or ( n49664 , n49662 , n49663 );
and ( n49665 , n33415 , n382983 );
or ( n49666 , n382995 , n18483 );
or ( n49667 , n36293 , n383001 );
or ( n49668 , n382993 , n33443 );
nand ( n49669 , n49666 , n49667 , n49668 );
nor ( n49670 , n49665 , n49669 );
nand ( n49671 , n49664 , n49670 );
buf ( n49672 , n49671 );
or ( n49673 , n31793 , n384523 );
and ( n49674 , n31770 , RI15b5c868_1022);
and ( n49675 , n46429 , n387126 );
and ( n49676 , n31778 , n384421 );
nor ( n49677 , n49674 , n49675 , n49676 );
nand ( n49678 , n49673 , n387147 , n49677 );
buf ( n49679 , n49678 );
buf ( n49680 , n32676 );
buf ( n49681 , n380903 );
not ( n49682 , RI15b52638_676);
not ( n49683 , n32397 );
or ( n49684 , n49682 , n49683 );
or ( n49685 , n35132 , n32401 );
nand ( n49686 , n49685 , n381450 );
and ( n49687 , n49686 , n35135 );
and ( n49688 , n35138 , n381461 );
nor ( n49689 , n49687 , n49688 , n43884 );
nand ( n49690 , n49684 , n49689 );
buf ( n49691 , n49690 );
buf ( n49692 , n382071 );
buf ( n49693 , n381490 );
buf ( n49694 , n379802 );
buf ( n49695 , n381872 );
not ( n49696 , RI15b46d88_282);
not ( n49697 , n379832 );
or ( n49698 , n49696 , n49697 );
and ( n49699 , n379820 , RI15b65e68_1342);
and ( n49700 , n379825 , RI15b48a98_344);
nor ( n49701 , n49699 , n49700 );
nand ( n49702 , n49698 , n49701 );
buf ( n49703 , n49702 );
buf ( n49704 , n19651 );
or ( n49705 , n22102 , n36813 );
and ( n49706 , n22203 , n37013 );
or ( n49707 , n36824 , n385525 );
or ( n49708 , n22293 , n36830 );
or ( n49709 , n36822 , n22299 );
nand ( n49710 , n49707 , n49708 , n49709 );
nor ( n49711 , n49706 , n49710 );
nand ( n49712 , n49705 , n49711 );
buf ( n49713 , n49712 );
buf ( n49714 , n22653 );
buf ( n49715 , n380940 );
buf ( n49716 , n381006 );
buf ( n49717 , n381006 );
buf ( n49718 , n22408 );
buf ( n49719 , n32981 );
buf ( n49720 , n22009 );
or ( n49721 , n36119 , n35930 );
and ( n49722 , n36974 , RI15b40de8_78);
or ( n49723 , n35582 , n35950 );
or ( n49724 , n35856 , n35944 );
or ( n49725 , n35934 , n35858 );
nand ( n49726 , n49723 , n49724 , n49725 );
nor ( n49727 , n49722 , n49726 );
nand ( n49728 , n49721 , n49727 );
buf ( n49729 , n49728 );
not ( n49730 , n47109 );
not ( n49731 , n35838 );
or ( n49732 , n49730 , n49731 );
and ( n49733 , n33196 , n36986 );
not ( n49734 , RI15b40230_53);
or ( n49735 , n35967 , n49734 );
or ( n49736 , n22241 , n35973 );
or ( n49737 , n35965 , n33201 );
nand ( n49738 , n49735 , n49736 , n49737 );
nor ( n49739 , n49733 , n49738 );
nand ( n49740 , n49732 , n49739 );
buf ( n49741 , n49740 );
buf ( n49742 , n31033 );
buf ( n49743 , n383613 );
or ( n49744 , n386705 , n48936 );
and ( n49745 , n386716 , n48939 );
not ( n49746 , RI15b4ee70_557);
or ( n49747 , n48948 , n49746 );
or ( n49748 , n37443 , n48953 );
or ( n49749 , n48946 , n386738 );
nand ( n49750 , n49747 , n49748 , n49749 );
nor ( n49751 , n49745 , n49750 );
nand ( n49752 , n49744 , n49751 );
buf ( n49753 , n49752 );
buf ( n49754 , n380906 );
not ( n49755 , RI15b60030_1141);
not ( n49756 , n383601 );
or ( n49757 , n49755 , n49756 );
or ( n49758 , n32307 , n33577 );
nand ( n49759 , n49758 , n33584 );
and ( n49760 , n49759 , n32289 );
not ( n49761 , n32307 );
nor ( n49762 , n49761 , n32289 );
and ( n49763 , n49762 , n40781 );
and ( n49764 , n383607 , RI15b5ea28_1094);
nor ( n49765 , n49760 , n49763 , n49764 );
nand ( n49766 , n49757 , n49765 );
buf ( n49767 , n49766 );
not ( n49768 , RI15b65a30_1333);
not ( n49769 , n35176 );
or ( n49770 , n49768 , n49769 );
nand ( n49771 , n379835 , n22266 );
nand ( n49772 , n35187 , RI15b48660_335);
not ( n49773 , n40200 );
and ( n49774 , n386554 , n49773 );
not ( n49775 , RI15b48660_335);
not ( n49776 , n35338 );
or ( n49777 , n49775 , n49776 );
or ( n49778 , n35338 , RI15b48660_335);
nand ( n49779 , n49777 , n49778 );
and ( n49780 , n35363 , n49779 );
nor ( n49781 , n49774 , n49780 );
and ( n49782 , n49771 , n49772 , n49781 );
nand ( n49783 , n49770 , n49782 );
buf ( n49784 , n49783 );
buf ( n49785 , n31033 );
buf ( n49786 , n380865 );
buf ( n49787 , n21800 );
buf ( n49788 , n33250 );
buf ( n49789 , n39264 );
buf ( n49790 , n386760 );
not ( n49791 , n386515 );
not ( n49792 , n386441 );
and ( n49793 , n49791 , n49792 );
or ( n49794 , n386541 , n385863 );
or ( n49795 , n385877 , n386550 );
or ( n49796 , n40100 , n386557 );
nand ( n49797 , n49794 , n49795 , n49796 );
nor ( n49798 , n49793 , n49797 );
nand ( n49799 , n40118 , n49798 );
buf ( n49800 , n49799 );
buf ( n49801 , n36704 );
buf ( n49802 , n380906 );
buf ( n49803 , n33382 );
buf ( n49804 , n380942 );
nand ( n49805 , n47023 , n47025 );
not ( n49806 , n49805 );
buf ( n49807 , n31453 );
not ( n49808 , n49807 );
and ( n49809 , n49806 , n49808 );
not ( n49810 , n49806 );
not ( n49811 , n49808 );
and ( n49812 , n49810 , n49811 );
nor ( n49813 , n49809 , n49812 );
not ( n49814 , n31601 );
or ( n49815 , n49813 , n49814 );
nand ( n49816 , n42049 , n31656 );
or ( n49817 , n49816 , n31667 );
nand ( n49818 , n49817 , n31700 );
and ( n49819 , n49818 , n379248 );
not ( n49820 , n49816 );
or ( n49821 , n49820 , n40972 , n379248 );
and ( n49822 , n379394 , RI15b58038_868);
and ( n49823 , n47038 , RI15b51e40_659);
nor ( n49824 , n49822 , n49823 );
nand ( n49825 , n49821 , n49824 );
nor ( n49826 , n49819 , n49825 );
nand ( n49827 , n49815 , n49826 );
buf ( n49828 , n49827 );
buf ( n49829 , n35649 );
nor ( n49830 , n31892 , n31898 );
not ( n49831 , n49830 );
nand ( n49832 , n49831 , n39025 );
buf ( n49833 , n384391 );
nand ( n49834 , n49832 , n49833 );
and ( n49835 , n31842 , n31849 );
not ( n49836 , n31842 );
not ( n49837 , n31849 );
and ( n49838 , n49836 , n49837 );
nor ( n49839 , n49835 , n49838 );
nand ( n49840 , n49839 , n31882 );
and ( n49841 , n31934 , n31940 );
not ( n49842 , n31934 );
not ( n49843 , n31940 );
and ( n49844 , n49842 , n49843 );
nor ( n49845 , n49841 , n49844 );
not ( n49846 , n31958 );
and ( n49847 , n49845 , n49846 );
nor ( n49848 , n19512 , n379720 );
nor ( n49849 , n49847 , n49848 );
and ( n49850 , n49834 , n49840 , n49849 );
and ( n49851 , n31792 , n49843 );
not ( n49852 , RI15b5d060_1039);
or ( n49853 , n31771 , n49852 );
or ( n49854 , n31898 , n32378 );
or ( n49855 , n31779 , n31849 );
nand ( n49856 , n49853 , n49854 , n49855 );
nor ( n49857 , n49851 , n49856 );
nand ( n49858 , n49850 , n49857 );
buf ( n49859 , n49858 );
buf ( n49860 , n384996 );
buf ( n49861 , RI15b5dba0_1063);
or ( n49862 , n36119 , n36306 );
and ( n49863 , n44133 , RI15b41928_102);
or ( n49864 , n35856 , n36316 );
or ( n49865 , n35582 , n36325 );
or ( n49866 , n22135 , n35858 );
nand ( n49867 , n49864 , n49865 , n49866 );
nor ( n49868 , n49863 , n49867 );
nand ( n49869 , n49862 , n49868 );
buf ( n49870 , n49869 );
buf ( n49871 , n382537 );
buf ( n49872 , n382071 );
buf ( n49873 , n22788 );
buf ( n49874 , n22007 );
not ( n49875 , n34281 );
nand ( n49876 , n49875 , n379785 );
not ( n49877 , n49876 );
not ( n49878 , n36496 );
or ( n49879 , n49877 , n49878 );
not ( n49880 , n34192 );
buf ( n49881 , n49880 );
nand ( n49882 , n49879 , n49881 );
nor ( n49883 , n49875 , n49880 );
nand ( n49884 , n36580 , n49883 );
not ( n49885 , n39187 );
not ( n49886 , n49885 );
buf ( n49887 , n39186 );
not ( n49888 , n49887 );
or ( n49889 , n49886 , n49888 );
or ( n49890 , n49887 , n49885 );
nand ( n49891 , n49889 , n49890 );
and ( n49892 , n49891 , n22440 );
and ( n49893 , n379783 , RI15b63d98_1272);
and ( n49894 , n34651 , RI15b5dba0_1063);
nor ( n49895 , n49892 , n49893 , n49894 );
nand ( n49896 , n49882 , n49884 , n49895 );
buf ( n49897 , n49896 );
and ( n49898 , n40674 , RI15b54438_740);
and ( n49899 , n49523 , RI15b51300_635);
nor ( n49900 , n49898 , n49899 );
not ( n49901 , n49900 );
buf ( n49902 , n49901 );
buf ( n49903 , n379847 );
or ( n49904 , n379976 , n380001 );
buf ( n49905 , n43931 );
not ( n49906 , n49905 );
or ( n49907 , n35769 , n49906 );
and ( n49908 , n379975 , RI15b561c0_803);
not ( n49909 , n379975 );
and ( n49910 , n49909 , n379976 );
nor ( n49911 , n49908 , n49910 );
or ( n49912 , n379948 , n49911 );
nand ( n49913 , n49904 , n49907 , n49912 );
buf ( n49914 , n49913 );
buf ( n49915 , RI15b47508_298);
buf ( n49916 , n22408 );
not ( n49917 , n47644 );
not ( n49918 , n382912 );
or ( n49919 , n49917 , n49918 );
and ( n49920 , n382931 , n47649 );
or ( n49921 , n47658 , n18529 );
or ( n49922 , n35805 , n47663 );
or ( n49923 , n47656 , n382967 );
nand ( n49924 , n49921 , n49922 , n49923 );
nor ( n49925 , n49920 , n49924 );
nand ( n49926 , n49919 , n49925 );
buf ( n49927 , n49926 );
buf ( n49928 , n43349 );
buf ( n49929 , n381490 );
buf ( n49930 , n379802 );
buf ( n49931 , n35649 );
not ( n49932 , n41756 );
not ( n49933 , n384726 );
or ( n49934 , n49932 , n49933 );
and ( n49935 , n35477 , n41446 );
or ( n49936 , n41455 , n17758 );
or ( n49937 , n39386 , n41461 );
or ( n49938 , n41453 , n384759 );
nand ( n49939 , n49936 , n49937 , n49938 );
nor ( n49940 , n49935 , n49939 );
nand ( n49941 , n49934 , n49940 );
buf ( n49942 , n49941 );
buf ( n49943 , n19653 );
or ( n49944 , n31091 , n32282 );
and ( n49945 , n41962 , n47195 );
or ( n49946 , n31052 , n386573 );
not ( n49947 , n41415 );
and ( n49948 , n49947 , RI15b61548_1186);
not ( n49949 , n49947 );
and ( n49950 , n49949 , n32282 );
nor ( n49951 , n49948 , n49950 );
or ( n49952 , n49951 , n45455 );
nand ( n49953 , n384906 , n386615 );
nand ( n49954 , n49946 , n49952 , n49953 );
nor ( n49955 , n49945 , n49954 );
nand ( n49956 , n49944 , n49955 );
buf ( n49957 , n49956 );
or ( n49958 , n386588 , n381569 );
and ( n49959 , n386600 , n381599 );
or ( n49960 , n381609 , n19165 );
or ( n49961 , n386618 , n381619 );
or ( n49962 , n381607 , n386627 );
nand ( n49963 , n49960 , n49961 , n49962 );
nor ( n49964 , n49959 , n49963 );
nand ( n49965 , n49958 , n49964 );
buf ( n49966 , n49965 );
buf ( n49967 , n379895 );
not ( n49968 , RI15b55ef0_797);
not ( n49969 , n380000 );
or ( n49970 , n49968 , n49969 );
and ( n49971 , n386666 , n381696 );
not ( n49972 , RI15b55ef0_797);
not ( n49973 , n379967 );
or ( n49974 , n49972 , n49973 );
or ( n49975 , n379967 , RI15b55ef0_797);
nand ( n49976 , n49974 , n49975 );
and ( n49977 , n49976 , n379949 );
nor ( n49978 , n49971 , n49977 );
nand ( n49979 , n49970 , n49978 );
buf ( n49980 , n49979 );
buf ( n49981 , n386762 );
buf ( n49982 , n381006 );
buf ( n49983 , n19774 );
and ( n49984 , n49983 , n19920 );
nor ( n49985 , n49984 , n384684 );
or ( n49986 , n49985 , n19780 );
not ( n49987 , n49983 );
nand ( n49988 , n49987 , n19780 );
or ( n49989 , n49988 , n380869 );
and ( n49990 , n20641 , RI15b4b5b8_436);
not ( n49991 , n20502 );
not ( n49992 , n19966 );
not ( n49993 , n49992 );
and ( n49994 , n49991 , n49993 );
nor ( n49995 , n49994 , n31809 );
or ( n49996 , n49995 , n19967 );
not ( n49997 , n20539 );
not ( n49998 , n49997 );
not ( n49999 , RI15b4b5b8_436);
and ( n50000 , n49998 , n49999 );
and ( n50001 , n49997 , RI15b4b5b8_436);
nor ( n50002 , n50000 , n50001 );
or ( n50003 , n50002 , n22354 );
and ( n50004 , n22361 , n49992 , n19967 );
or ( n50005 , n20653 , n19666 );
nand ( n50006 , n50005 , n42328 );
nor ( n50007 , n50004 , n50006 );
nand ( n50008 , n49996 , n50003 , n50007 );
nor ( n50009 , n49990 , n50008 );
nand ( n50010 , n49986 , n49989 , n50009 );
buf ( n50011 , n50010 );
buf ( n50012 , n382073 );
buf ( n50013 , n384700 );
buf ( n50014 , n22406 );
buf ( n50015 , n22007 );
not ( n50016 , n31965 );
not ( n50017 , n383428 );
or ( n50018 , n50016 , n50017 );
nand ( n50019 , n50018 , n384642 );
nand ( n50020 , n50019 , RI15b638e8_1262);
and ( n50021 , n386938 , n19630 );
nor ( n50022 , n383428 , RI15b638e8_1262);
and ( n50023 , n384655 , n50022 );
nor ( n50024 , n50021 , n50023 );
nand ( n50025 , n45337 , n50020 , n50024 );
buf ( n50026 , n50025 );
not ( n50027 , n33578 );
not ( n50028 , n50027 );
not ( n50029 , n32339 );
or ( n50030 , n50028 , n50029 );
nand ( n50031 , n50030 , n33584 );
nand ( n50032 , n50031 , n32353 );
nand ( n50033 , n32355 , n40781 );
nand ( n50034 , n383601 , RI15b60210_1145);
nand ( n50035 , n383607 , RI15b5ec08_1098);
nand ( n50036 , n50032 , n50033 , n50034 , n50035 );
buf ( n50037 , n50036 );
buf ( n50038 , n30992 );
or ( n50039 , n36238 , n48938 );
not ( n50040 , n48948 );
and ( n50041 , n50040 , RI15b4ec90_553);
or ( n50042 , n48953 , n48296 );
or ( n50043 , n48936 , n383802 );
or ( n50044 , n48946 , n42402 );
nand ( n50045 , n50042 , n50043 , n50044 );
nor ( n50046 , n50041 , n50045 );
nand ( n50047 , n50039 , n50046 );
buf ( n50048 , n50047 );
buf ( n50049 , n382069 );
buf ( n50050 , n19651 );
buf ( n50051 , n382049 );
buf ( n50052 , n383498 );
not ( n50053 , n34931 );
nor ( n50054 , n48175 , n48179 );
not ( n50055 , n50054 );
or ( n50056 , n50053 , n50055 );
nand ( n50057 , n50056 , n46513 );
not ( n50058 , n35055 );
nand ( n50059 , n50057 , n50058 );
not ( n50060 , n50054 );
nor ( n50061 , n35117 , n50058 );
and ( n50062 , n50060 , n50061 );
and ( n50063 , n385213 , RI15b47d00_315);
and ( n50064 , n20631 , RI15b466f8_268);
nor ( n50065 , n50063 , n50064 );
not ( n50066 , n50065 );
nor ( n50067 , n50062 , n50066 );
nand ( n50068 , n50059 , n50067 );
buf ( n50069 , n50068 );
buf ( n50070 , n387159 );
buf ( n50071 , n383345 );
buf ( n50072 , n18226 );
buf ( n50073 , n33382 );
not ( n50074 , n382898 );
not ( n50075 , n37629 );
or ( n50076 , n50074 , n50075 );
and ( n50077 , n37637 , n382934 );
not ( n50078 , RI15b597a8_918);
or ( n50079 , n382949 , n50078 );
not ( n50080 , n43000 );
or ( n50081 , n50080 , n382965 );
or ( n50082 , n382947 , n37646 );
nand ( n50083 , n50079 , n50081 , n50082 );
nor ( n50084 , n50077 , n50083 );
nand ( n50085 , n50076 , n50084 );
buf ( n50086 , n50085 );
not ( n50087 , n39530 );
or ( n50088 , n50087 , n39537 );
nor ( n50089 , n382683 , RI15b556f8_780);
and ( n50090 , n382688 , n50089 );
not ( n50091 , n382832 );
nand ( n50092 , n50091 , n382880 );
not ( n50093 , n50092 );
and ( n50094 , n382834 , RI15b4d598_504);
and ( n50095 , n382838 , RI15b4e498_536);
nor ( n50096 , n50094 , n50095 );
and ( n50097 , n382842 , RI15b4e0d8_528);
and ( n50098 , n382844 , RI15b4d958_512);
and ( n50099 , n382846 , RI15b4e858_544);
nor ( n50100 , n50097 , n50098 , n50099 );
and ( n50101 , n382850 , RI15b4ec18_552);
and ( n50102 , n382853 , RI15b4ca58_480);
nor ( n50103 , n50101 , n50102 );
and ( n50104 , n382857 , RI15b4efd8_560);
and ( n50105 , n379880 , RI15b4d1d8_496);
nor ( n50106 , n50104 , n50105 );
nand ( n50107 , n50096 , n50100 , n50103 , n50106 );
not ( n50108 , n50107 );
and ( n50109 , n382864 , RI15b4ce18_488);
and ( n50110 , n380061 , RI15b4f398_568);
and ( n50111 , n382867 , RI15b4c698_472);
nor ( n50112 , n50109 , n50110 , n50111 );
and ( n50113 , n382870 , RI15b4fb18_584);
and ( n50114 , n382872 , RI15b4f758_576);
nor ( n50115 , n50113 , n50114 );
and ( n50116 , n382875 , RI15b4dd18_520);
and ( n50117 , n382877 , RI15b4fed8_592);
nor ( n50118 , n50116 , n50117 );
nand ( n50119 , n50108 , n50112 , n50115 , n50118 );
not ( n50120 , n50119 );
and ( n50121 , n50093 , n50120 );
and ( n50122 , n50092 , n50119 );
nor ( n50123 , n50121 , n50122 );
or ( n50124 , n50123 , n382886 );
or ( n50125 , n383730 , n382691 );
buf ( n50126 , n381320 );
nor ( n50127 , n381400 , n50126 );
not ( n50128 , n50127 );
nand ( n50129 , n50124 , n50125 , n50128 );
nor ( n50130 , n50090 , n50129 );
nand ( n50131 , n50088 , n50130 );
buf ( n50132 , n50131 );
buf ( n50133 , n381004 );
or ( n50134 , n19608 , n383598 );
nand ( n50135 , n50134 , RI15b62b50_1233);
not ( n50136 , n42011 );
not ( n50137 , n46537 );
or ( n50138 , n50136 , n50137 );
nand ( n50139 , n50138 , n19281 );
nand ( n50140 , n50135 , n42034 , n50139 );
buf ( n50141 , n50140 );
buf ( n50142 , n387159 );
buf ( n50143 , n380942 );
or ( n50144 , n36238 , n38827 );
not ( n50145 , n38837 );
and ( n50146 , n50145 , RI15b4c350_465);
or ( n50147 , n38841 , n32710 );
or ( n50148 , n38825 , n383802 );
or ( n50149 , n38835 , n42402 );
nand ( n50150 , n50147 , n50148 , n50149 );
nor ( n50151 , n50146 , n50150 );
nand ( n50152 , n50144 , n50151 );
buf ( n50153 , n50152 );
buf ( n50154 , n22009 );
buf ( n50155 , n22402 );
buf ( n50156 , n379403 );
and ( n50157 , n21788 , RI15b56fd0_833);
and ( n50158 , n22488 , n21770 );
not ( n50159 , n17547 );
and ( n50160 , n50159 , n22481 );
not ( n50161 , n50159 );
and ( n50162 , n50161 , RI15b56fd0_833);
nor ( n50163 , n50160 , n50162 );
and ( n50164 , n50163 , n384127 );
nor ( n50165 , n50157 , n50158 , n50164 );
nand ( n50166 , n47892 , n50165 );
buf ( n50167 , n50166 );
buf ( n50168 , n22499 );
nor ( n50169 , n50168 , n22488 );
and ( n50170 , n21802 , n50169 );
and ( n50171 , n42563 , RI15b57ed0_865);
not ( n50172 , n21949 );
buf ( n50173 , n22579 );
not ( n50174 , n50173 );
or ( n50175 , n50172 , n50174 );
nand ( n50176 , n50175 , n21979 );
and ( n50177 , n50176 , RI15b560d0_801);
or ( n50178 , n50173 , n21982 , RI15b560d0_801);
and ( n50179 , n42561 , n22611 , RI15b57e58_864);
and ( n50180 , n22610 , RI15b57ed0_865);
nor ( n50181 , n50179 , n50180 );
or ( n50182 , n21922 , n50181 );
nand ( n50183 , n50178 , n50182 );
nor ( n50184 , n50171 , n50177 , n50183 );
or ( n50185 , n50184 , n18078 );
and ( n50186 , n18177 , RI15b57ed0_865);
and ( n50187 , n18219 , RI15b56fd0_833);
nor ( n50188 , n50186 , n50187 , n21751 );
nand ( n50189 , n50185 , n50188 );
nor ( n50190 , n50170 , n50189 );
nand ( n50191 , n50168 , n17507 );
not ( n50192 , n50191 );
not ( n50193 , n17565 );
or ( n50194 , n50192 , n50193 );
nand ( n50195 , n50194 , n22488 );
nand ( n50196 , n50190 , n50195 );
buf ( n50197 , n50196 );
buf ( n50198 , n386762 );
buf ( n50199 , n32271 );
buf ( n50200 , n22007 );
buf ( n50201 , n385195 );
not ( n50202 , n33387 );
not ( n50203 , n37629 );
or ( n50204 , n50202 , n50203 );
and ( n50205 , n37637 , n33417 );
not ( n50206 , RI15b5b5a8_982);
or ( n50207 , n33428 , n50206 );
not ( n50208 , n37643 );
or ( n50209 , n50208 , n33440 );
or ( n50210 , n33426 , n37646 );
nand ( n50211 , n50207 , n50209 , n50210 );
nor ( n50212 , n50205 , n50211 );
nand ( n50213 , n50204 , n50212 );
buf ( n50214 , n50213 );
not ( n50215 , RI15b538f8_716);
not ( n50216 , n383170 );
or ( n50217 , n50215 , n50216 );
or ( n50218 , n33454 , n40055 );
nand ( n50219 , n50218 , n33465 );
and ( n50220 , n50219 , n40046 );
not ( n50221 , n40055 );
nor ( n50222 , n50221 , n40046 );
and ( n50223 , n33476 , n50222 );
and ( n50224 , n383147 , RI15b53178_700);
nor ( n50225 , n50220 , n50223 , n50224 );
nand ( n50226 , n50217 , n50225 );
buf ( n50227 , n50226 );
buf ( n50228 , n22009 );
buf ( n50229 , n22007 );
buf ( n50230 , n379802 );
buf ( n50231 , n380865 );
not ( n50232 , RI15b47148_290);
not ( n50233 , n385213 );
or ( n50234 , n50232 , n50233 );
and ( n50235 , n385221 , RI15b486d8_336);
and ( n50236 , n20631 , RI15b469c8_274);
nor ( n50237 , n50235 , n50236 );
nand ( n50238 , n50234 , n50237 );
buf ( n50239 , n50238 );
buf ( n50240 , n32160 );
or ( n50241 , n35523 , n22030 );
nand ( n50242 , n35525 , RI15b538f8_716);
nand ( n50243 , n50241 , n50242 );
buf ( n50244 , n50243 );
buf ( n50245 , n31719 );
buf ( n50246 , n379844 );
not ( n50247 , n48975 );
and ( n50248 , n50247 , n34999 );
not ( n50249 , n50247 );
and ( n50250 , n50249 , RI15b490b0_357);
nor ( n50251 , n50248 , n50250 );
not ( n50252 , n48991 );
nand ( n50253 , n50251 , n50252 );
nand ( n50254 , n48980 , RI15b490b0_357);
and ( n50255 , n48910 , n48998 );
and ( n50256 , n35335 , RI15b66480_1355);
nor ( n50257 , n50255 , n50256 );
nand ( n50258 , n50253 , n50254 , n43161 , n50257 );
buf ( n50259 , n50258 );
buf ( n50260 , n384700 );
buf ( n50261 , n381872 );
nand ( n50262 , n40503 , RI15b607b0_1157);
or ( n50263 , n22462 , RI15b607b0_1157);
nand ( n50264 , n50263 , n35509 );
nand ( n50265 , n50262 , n50264 , n380773 );
buf ( n50266 , n50265 );
buf ( n50267 , n382065 );
buf ( n50268 , n18226 );
buf ( n50269 , n382071 );
or ( n50270 , n386705 , n33111 );
and ( n50271 , n386716 , n33117 );
not ( n50272 , RI15b4e6f0_541);
or ( n50273 , n33128 , n50272 );
or ( n50274 , n45435 , n33134 );
or ( n50275 , n33126 , n386738 );
nand ( n50276 , n50273 , n50274 , n50275 );
nor ( n50277 , n50271 , n50276 );
nand ( n50278 , n50270 , n50277 );
buf ( n50279 , n50278 );
not ( n50280 , n48052 );
not ( n50281 , n32129 );
or ( n50282 , n50280 , n50281 );
and ( n50283 , n44521 , RI15b424e0_127);
or ( n50284 , n32141 , n37497 );
or ( n50285 , n32148 , n37512 );
or ( n50286 , n37505 , n32150 );
nand ( n50287 , n50284 , n50285 , n50286 );
nor ( n50288 , n50283 , n50287 );
nand ( n50289 , n50282 , n50288 );
buf ( n50290 , n50289 );
buf ( n50291 , n384996 );
buf ( n50292 , n380903 );
buf ( n50293 , n384199 );
buf ( n50294 , n385197 );
buf ( n50295 , n35649 );
and ( n50296 , n22646 , RI15b458e8_238);
and ( n50297 , n22648 , RI15b51d50_657);
nor ( n50298 , n50296 , n50297 );
not ( n50299 , n50298 );
buf ( n50300 , n50299 );
buf ( n50301 , n20663 );
and ( n50302 , n385971 , n385986 );
not ( n50303 , n50302 );
buf ( n50304 , n385939 );
buf ( n50305 , n50304 );
not ( n50306 , n50305 );
and ( n50307 , n50306 , RI15b448f8_204);
nand ( n50308 , n385975 , RI15b44880_203);
nor ( n50309 , n50308 , RI15b448f8_204);
not ( n50310 , n50309 );
not ( n50311 , n50304 );
or ( n50312 , n50310 , n50311 );
nand ( n50313 , n50308 , RI15b448f8_204);
nand ( n50314 , n50312 , n50313 );
nor ( n50315 , n50307 , n50314 );
not ( n50316 , n50315 );
and ( n50317 , n50303 , n50316 );
not ( n50318 , n50303 );
and ( n50319 , n50318 , n50315 );
nor ( n50320 , n50317 , n50319 );
not ( n50321 , n386020 );
nor ( n50322 , n50320 , n50321 );
nand ( n50323 , n386241 , n386248 );
not ( n50324 , n386040 );
not ( n50325 , n50324 );
not ( n50326 , RI15b448f8_204);
or ( n50327 , n50325 , n50326 );
nand ( n50328 , n50325 , n50309 );
nand ( n50329 , n50327 , n50328 , n50313 );
and ( n50330 , n50323 , n50329 );
not ( n50331 , n50323 );
not ( n50332 , n50329 );
and ( n50333 , n50331 , n50332 );
nor ( n50334 , n50330 , n50333 );
nor ( n50335 , n50334 , n386265 );
buf ( n50336 , n386279 );
and ( n50337 , n50336 , RI15b448f8_204);
not ( n50338 , n50309 );
not ( n50339 , n386278 );
or ( n50340 , n50338 , n50339 );
nand ( n50341 , n50340 , n50313 );
nor ( n50342 , n50337 , n50341 );
not ( n50343 , n50342 );
not ( n50344 , n50343 );
not ( n50345 , n386497 );
or ( n50346 , n50344 , n50345 );
not ( n50347 , n386497 );
nand ( n50348 , n50347 , n50342 );
nand ( n50349 , n50346 , n50348 );
nand ( n50350 , n50349 , n386500 );
buf ( n50351 , n48527 );
nand ( n50352 , n50351 , RI15b4bf90_457);
nand ( n50353 , n50350 , n50352 );
nor ( n50354 , n50322 , n50335 , n50353 );
not ( n50355 , n20637 );
not ( n50356 , n19924 );
or ( n50357 , n50355 , n50356 );
nand ( n50358 , n50357 , n34798 );
and ( n50359 , n50358 , RI15b4b090_425);
or ( n50360 , n34801 , n19924 , RI15b4b090_425);
not ( n50361 , n19951 );
or ( n50362 , n50361 , n22216 );
nand ( n50363 , n50360 , n50362 );
nor ( n50364 , n50359 , n50363 );
nand ( n50365 , n50354 , n50364 );
buf ( n50366 , n50365 );
buf ( n50367 , n386814 );
or ( n50368 , n50367 , n22473 );
nand ( n50369 , n50368 , n386942 );
nand ( n50370 , n50369 , n19625 );
not ( n50371 , n19625 );
nand ( n50372 , n50371 , n45576 , n50367 );
buf ( n50373 , n386965 );
and ( n50374 , n45578 , n50373 );
nor ( n50375 , n50374 , n40140 );
or ( n50376 , n50375 , n386966 );
and ( n50377 , n40145 , RI15b63e10_1273);
or ( n50378 , n34826 , n50373 , RI15b62010_1209);
not ( n50379 , n387026 );
not ( n50380 , RI15b63e10_1273);
and ( n50381 , n50379 , n50380 );
and ( n50382 , n387026 , RI15b63e10_1273);
nor ( n50383 , n50381 , n50382 );
or ( n50384 , n34833 , n50383 );
nand ( n50385 , n50378 , n50384 );
nor ( n50386 , n50377 , n50385 );
nand ( n50387 , n50376 , n50386 );
nand ( n50388 , n50387 , n19201 );
and ( n50389 , n22423 , RI15b63e10_1273);
and ( n50390 , n19599 , RI15b62f10_1241);
nor ( n50391 , n50389 , n50390 , n19513 );
nand ( n50392 , n50370 , n50372 , n50388 , n50391 );
buf ( n50393 , n50392 );
buf ( n50394 , n381490 );
buf ( n50395 , n22404 );
buf ( n50396 , n383174 );
not ( n50397 , n45762 );
not ( n50398 , n50397 );
not ( n50399 , n45120 );
or ( n50400 , n50398 , n50399 );
nand ( n50401 , n50400 , n33584 );
nand ( n50402 , n50401 , n45135 );
nor ( n50403 , n45135 , n33588 );
and ( n50404 , n45137 , n50403 );
and ( n50405 , n383601 , RI15b605d0_1153);
and ( n50406 , n383607 , RI15b5efc8_1106);
nor ( n50407 , n50405 , n50406 );
not ( n50408 , n50407 );
nor ( n50409 , n50404 , n50408 );
nand ( n50410 , n50402 , n50409 );
buf ( n50411 , n50410 );
buf ( n50412 , n19653 );
or ( n50413 , n36238 , n33599 );
not ( n50414 , n33609 );
and ( n50415 , n50414 , RI15b4e8d0_545);
or ( n50416 , n33615 , n32710 );
or ( n50417 , n33597 , n383802 );
or ( n50418 , n33607 , n42402 );
nand ( n50419 , n50416 , n50417 , n50418 );
nor ( n50420 , n50415 , n50419 );
nand ( n50421 , n50413 , n50420 );
buf ( n50422 , n50421 );
buf ( n50423 , n380940 );
buf ( n50424 , n22716 );
buf ( n50425 , n22740 );
buf ( n50426 , n31979 );
buf ( n50427 , n32676 );
or ( n50428 , n39265 , n22083 );
nand ( n50429 , n35525 , RI15b54000_731);
nand ( n50430 , n50428 , n50429 );
buf ( n50431 , n50430 );
and ( n50432 , n379822 , n44787 );
nor ( n50433 , n379834 , n382012 );
nor ( n50434 , n50432 , n50433 );
and ( n50435 , n32747 , RI15b42990_137);
and ( n50436 , n32753 , RI15b416d0_97);
and ( n50437 , n32762 , RI15b41310_89);
nor ( n50438 , n50436 , n50437 );
and ( n50439 , n32755 , RI15b41a90_105);
and ( n50440 , n32759 , RI15b40f50_81);
nor ( n50441 , n50439 , n50440 );
and ( n50442 , n32766 , RI15b434d0_161);
and ( n50443 , n32768 , RI15b43110_153);
nor ( n50444 , n50442 , n50443 );
and ( n50445 , n32771 , RI15b43890_169);
and ( n50446 , n32773 , RI15b42d50_145);
nor ( n50447 , n50445 , n50446 );
nand ( n50448 , n50438 , n50441 , n50444 , n50447 );
and ( n50449 , n46812 , n50448 );
and ( n50450 , n32781 , RI15b40410_57);
nor ( n50451 , n50435 , n50449 , n50450 );
and ( n50452 , n32785 , RI15b425d0_129);
and ( n50453 , n32787 , RI15b42210_121);
nor ( n50454 , n50452 , n50453 );
and ( n50455 , n32792 , RI15b40050_49);
and ( n50456 , n32794 , RI15b41e50_113);
nor ( n50457 , n50455 , n50456 );
and ( n50458 , n32797 , RI15b407d0_65);
and ( n50459 , n32800 , RI15b40b90_73);
nor ( n50460 , n50458 , n50459 );
nand ( n50461 , n50451 , n50454 , n50457 , n50460 );
not ( n50462 , n35456 );
and ( n50463 , n50461 , n50462 );
and ( n50464 , n35335 , RI15b65d78_1340);
not ( n50465 , RI15b489a8_342);
not ( n50466 , n35349 );
not ( n50467 , n50466 );
or ( n50468 , n50465 , n50467 );
or ( n50469 , n50466 , RI15b489a8_342);
nand ( n50470 , n50468 , n50469 );
and ( n50471 , n35363 , n50470 );
nor ( n50472 , n50463 , n50464 , n50471 );
nand ( n50473 , n41726 , RI15b489a8_342);
nand ( n50474 , n50434 , n50472 , n50473 );
buf ( n50475 , n50474 );
buf ( n50476 , n379403 );
buf ( n50477 , n31719 );
buf ( n50478 , n22402 );
buf ( n50479 , n382049 );
buf ( n50480 , n31990 );
nor ( n50481 , n50480 , n382079 );
or ( n50482 , n50481 , n43097 );
nand ( n50483 , n50482 , n42700 );
nor ( n50484 , n32035 , n42700 );
and ( n50485 , n50480 , n50484 );
not ( n50486 , n32962 );
not ( n50487 , n382289 );
buf ( n50488 , n32005 );
not ( n50489 , n50488 );
and ( n50490 , n50487 , n50489 );
and ( n50491 , n382289 , n50488 );
nor ( n50492 , n50490 , n50491 );
or ( n50493 , n50486 , n50492 );
and ( n50494 , n382523 , RI15b4b630_437);
and ( n50495 , n32052 , RI15b45438_228);
nor ( n50496 , n50494 , n50495 );
nand ( n50497 , n50493 , n50496 );
nor ( n50498 , n50485 , n50497 );
nand ( n50499 , n50483 , n50498 );
buf ( n50500 , n50499 );
buf ( n50501 , n381081 );
nand ( n50502 , n31770 , RI15b5c430_1013);
or ( n50503 , n31781 , n31778 );
nand ( n50504 , n50503 , n19423 );
nand ( n50505 , n32386 , n18446 );
nand ( n50506 , n50502 , n50504 , n50505 , n46550 );
buf ( n50507 , n50506 );
buf ( n50508 , n383319 );
not ( n50509 , n44798 );
nor ( n50510 , n50508 , n50509 );
or ( n50511 , n50510 , n381449 );
not ( n50512 , n383294 );
not ( n50513 , n50512 );
nand ( n50514 , n50511 , n50513 );
nand ( n50515 , n50508 , n50512 , n381461 );
and ( n50516 , n381486 , RI15b52a70_685);
nor ( n50517 , n50516 , n46753 );
nand ( n50518 , n50514 , n50515 , n50517 );
buf ( n50519 , n50518 );
buf ( n50520 , n379893 );
or ( n50521 , n31771 , n18440 );
and ( n50522 , n39573 , n19299 );
and ( n50523 , n32386 , n18442 );
and ( n50524 , n31778 , n382582 );
nor ( n50525 , n50522 , n50523 , n50524 );
nand ( n50526 , n50521 , n382602 , n50525 );
buf ( n50527 , n50526 );
buf ( n50528 , n32676 );
not ( n50529 , n36268 );
not ( n50530 , n383138 );
not ( n50531 , n50530 );
or ( n50532 , n50529 , n50531 );
nand ( n50533 , n50532 , n381450 );
nand ( n50534 , n50533 , n383139 );
nor ( n50535 , n50530 , n383139 );
nand ( n50536 , n50535 , n381461 );
nand ( n50537 , n381485 , RI15b52818_680);
nor ( n50538 , n381400 , n384751 );
not ( n50539 , n50538 );
nand ( n50540 , n50534 , n50536 , n50537 , n50539 );
buf ( n50541 , n50540 );
buf ( n50542 , n383174 );
buf ( n50543 , n22408 );
buf ( n50544 , n383345 );
or ( n50545 , n37478 , n38373 );
and ( n50546 , n384983 , n38375 );
or ( n50547 , n38385 , n20398 );
or ( n50548 , n22022 , n38389 );
or ( n50549 , n38383 , n384988 );
nand ( n50550 , n50547 , n50548 , n50549 );
nor ( n50551 , n50546 , n50550 );
nand ( n50552 , n50545 , n50551 );
buf ( n50553 , n50552 );
buf ( n50554 , n381566 );
buf ( n50555 , n32160 );
and ( n50556 , n379822 , RI15b65a30_1333);
and ( n50557 , n379825 , RI15b48660_335);
nor ( n50558 , n50556 , n50557 );
nand ( n50559 , n379832 , RI15b46950_273);
nand ( n50560 , n50558 , n50559 , n49771 );
buf ( n50561 , n50560 );
buf ( n50562 , n22404 );
buf ( n50563 , n32981 );
buf ( n50564 , n35649 );
buf ( n50565 , n17499 );
or ( n50566 , n31149 , n386706 );
and ( n50567 , n31161 , n386718 );
not ( n50568 , RI15b4cf80_491);
or ( n50569 , n386727 , n50568 );
or ( n50570 , n32452 , n386735 );
or ( n50571 , n386725 , n31184 );
nand ( n50572 , n50569 , n50570 , n50571 );
nor ( n50573 , n50567 , n50572 );
nand ( n50574 , n50566 , n50573 );
buf ( n50575 , n50574 );
and ( n50576 , n22646 , RI15b45bb8_244);
and ( n50577 , n22648 , RI15b52020_663);
nor ( n50578 , n50576 , n50577 );
not ( n50579 , n50578 );
buf ( n50580 , n50579 );
or ( n50581 , n384021 , n386963 );
or ( n50582 , n18425 , n386747 );
not ( n50583 , n384033 );
and ( n50584 , n50583 , RI15b61f20_1207);
not ( n50585 , n50583 );
and ( n50586 , n50585 , n386963 );
nor ( n50587 , n50584 , n50586 );
or ( n50588 , n50587 , n384024 );
nand ( n50589 , n50581 , n50582 , n50588 );
buf ( n50590 , n50589 );
buf ( n50591 , n22740 );
buf ( n50592 , n382073 );
buf ( n50593 , n379847 );
not ( n50594 , RI15b65940_1331);
not ( n50595 , n35176 );
or ( n50596 , n50594 , n50595 );
nand ( n50597 , n35187 , RI15b48570_333);
and ( n50598 , n386554 , n32215 );
not ( n50599 , n35195 );
not ( n50600 , RI15b48570_333);
not ( n50601 , n35198 );
or ( n50602 , n50600 , n50601 );
or ( n50603 , n35198 , RI15b48570_333);
nand ( n50604 , n50602 , n50603 );
and ( n50605 , n50599 , n50604 );
nor ( n50606 , n50598 , n50605 );
and ( n50607 , n39235 , n50597 , n50606 );
nand ( n50608 , n50596 , n50607 );
buf ( n50609 , n50608 );
buf ( n50610 , n22404 );
buf ( n50611 , n22738 );
buf ( n50612 , n19653 );
buf ( n50613 , n31033 );
buf ( n50614 , n383174 );
not ( n50615 , n43975 );
not ( n50616 , n43982 );
or ( n50617 , n50615 , n50616 );
or ( n50618 , n43982 , n43975 );
nand ( n50619 , n50617 , n50618 );
not ( n50620 , n34867 );
nand ( n50621 , n50619 , n50620 );
not ( n50622 , n379391 );
buf ( n50623 , n31637 );
not ( n50624 , n50623 );
or ( n50625 , n50622 , n50624 );
nand ( n50626 , n50625 , n31700 );
buf ( n50627 , n31638 );
and ( n50628 , n50626 , n50627 );
or ( n50629 , n31707 , n50623 , n50627 );
and ( n50630 , n379394 , RI15b57a98_856);
and ( n50631 , n379398 , RI15b518a0_647);
nor ( n50632 , n50630 , n50631 );
nand ( n50633 , n50629 , n50632 );
nor ( n50634 , n50628 , n50633 );
nand ( n50635 , n50621 , n50634 );
buf ( n50636 , n50635 );
buf ( n50637 , n385197 );
not ( n50638 , n37774 );
not ( n50639 , n22445 );
and ( n50640 , n50638 , n50639 );
and ( n50641 , n47838 , n19201 );
nor ( n50642 , n50640 , n50641 );
not ( n50643 , n19590 );
and ( n50644 , n50643 , n22427 );
and ( n50645 , n19580 , n22428 );
nor ( n50646 , n50644 , n50645 , n19628 );
nand ( n50647 , n50642 , n50646 );
buf ( n50648 , n50647 );
buf ( n50649 , n19651 );
buf ( n50650 , n32676 );
nor ( n50651 , n49627 , n35049 );
or ( n50652 , n50651 , n49094 );
not ( n50653 , n386538 );
nor ( n50654 , n35184 , n50653 );
nand ( n50655 , n50652 , n50654 );
nand ( n50656 , n50655 , RI15b49308_362);
nor ( n50657 , n49632 , RI15b49308_362);
and ( n50658 , n50651 , n50657 );
nor ( n50659 , n386547 , n22254 );
nor ( n50660 , n50658 , n50659 );
nand ( n50661 , n50656 , n50660 );
buf ( n50662 , n50661 );
buf ( n50663 , n22479 );
buf ( n50664 , n386563 );
or ( n50665 , n381015 , n22241 );
nand ( n50666 , n35327 , RI15b536a0_711);
nand ( n50667 , n50665 , n50666 );
buf ( n50668 , n50667 );
buf ( n50669 , n379895 );
buf ( n50670 , n22655 );
nand ( n50671 , n41173 , n381549 );
nand ( n50672 , n384918 , RI15b5f310_1113);
nand ( n50673 , n37773 , n47530 );
nand ( n50674 , n36535 , n50671 , n50672 , n50673 );
buf ( n50675 , n50674 );
or ( n50676 , n36238 , n40472 );
not ( n50677 , n40480 );
and ( n50678 , n50677 , RI15b4fb90_585);
or ( n50679 , n383802 , n40468 );
or ( n50680 , n48296 , n40485 );
or ( n50681 , n40478 , n42402 );
nand ( n50682 , n50679 , n50680 , n50681 );
nor ( n50683 , n50678 , n50682 );
nand ( n50684 , n50676 , n50683 );
buf ( n50685 , n50684 );
buf ( n50686 , n380942 );
buf ( n50687 , n379802 );
buf ( n50688 , n22408 );
or ( n50689 , n22315 , n36082 );
and ( n50690 , n22326 , n36084 );
not ( n50691 , RI15b41310_89);
or ( n50692 , n36094 , n50691 );
or ( n50693 , n22334 , n36098 );
or ( n50694 , n36092 , n22336 );
nand ( n50695 , n50692 , n50693 , n50694 );
nor ( n50696 , n50690 , n50695 );
nand ( n50697 , n50689 , n50696 );
buf ( n50698 , n50697 );
nor ( n50699 , n38248 , n20637 );
or ( n50700 , n50699 , n20423 );
or ( n50701 , RI15b3fd08_42 , n22216 );
nor ( n50702 , n35876 , n22134 );
or ( n50703 , n50702 , n22298 );
nand ( n50704 , n50700 , n50701 , n50703 );
buf ( n50705 , n50704 );
buf ( n50706 , n33250 );
buf ( n50707 , n382065 );
buf ( n50708 , n382065 );
or ( n50709 , n380968 , n36082 );
and ( n50710 , n380986 , n36084 );
or ( n50711 , n36094 , n20363 );
or ( n50712 , n380994 , n36098 );
or ( n50713 , n36092 , n380996 );
nand ( n50714 , n50711 , n50712 , n50713 );
nor ( n50715 , n50710 , n50714 );
nand ( n50716 , n50709 , n50715 );
buf ( n50717 , n50716 );
buf ( n50718 , n22408 );
buf ( n50719 , n31719 );
and ( n50720 , n36768 , n20501 );
and ( n50721 , n20519 , RI15b3fc18_40);
nor ( n50722 , n50720 , n50721 );
not ( n50723 , n50722 );
buf ( n50724 , n50723 );
buf ( n50725 , n22479 );
or ( n50726 , n383180 , n381530 );
not ( n50727 , n381544 );
and ( n50728 , n50727 , RI15b5bc38_996);
or ( n50729 , n383184 , n381527 );
and ( n50730 , n381556 , n40017 );
and ( n50731 , n40019 , n381553 );
nor ( n50732 , n50730 , n50731 );
nand ( n50733 , n50729 , n50732 );
nor ( n50734 , n50728 , n50733 );
nand ( n50735 , n50726 , n50734 );
buf ( n50736 , n50735 );
buf ( n50737 , n50126 );
or ( n50738 , n42969 , n50737 );
not ( n50739 , n381332 );
nand ( n50740 , n50739 , n381321 );
nand ( n50741 , n381417 , n50740 );
not ( n50742 , n32401 );
not ( n50743 , n50742 );
or ( n50744 , n50743 , n40057 );
nand ( n50745 , n50744 , n381450 );
and ( n50746 , n50745 , n40066 );
and ( n50747 , n381461 , n40069 );
nor ( n50748 , n50746 , n50747 );
and ( n50749 , n50741 , n50748 );
nand ( n50750 , n381486 , RI15b53268_702);
nand ( n50751 , n50738 , n50749 , n50750 );
buf ( n50752 , n50751 );
buf ( n50753 , n380203 );
buf ( n50754 , n22408 );
buf ( n50755 , n385112 );
not ( n50756 , n46960 );
not ( n50757 , n32129 );
or ( n50758 , n50756 , n50757 );
and ( n50759 , n45035 , RI15b43020_151);
or ( n50760 , n32141 , n38377 );
or ( n50761 , n32148 , n38389 );
or ( n50762 , n38383 , n32150 );
nand ( n50763 , n50760 , n50761 , n50762 );
nor ( n50764 , n50759 , n50763 );
nand ( n50765 , n50758 , n50764 );
buf ( n50766 , n50765 );
buf ( n50767 , n381566 );
buf ( n50768 , n381021 );
buf ( n50769 , n380865 );
buf ( n50770 , n385195 );
not ( n50771 , n33387 );
not ( n50772 , n381507 );
or ( n50773 , n50771 , n50772 );
and ( n50774 , n381524 , n33417 );
not ( n50775 , RI15b5b788_986);
or ( n50776 , n33428 , n50775 );
or ( n50777 , n38012 , n33440 );
or ( n50778 , n33426 , n381560 );
nand ( n50779 , n50776 , n50777 , n50778 );
nor ( n50780 , n50774 , n50779 );
nand ( n50781 , n50773 , n50780 );
buf ( n50782 , n50781 );
not ( n50783 , RI15b53718_712);
not ( n50784 , n383170 );
or ( n50785 , n50783 , n50784 );
or ( n50786 , n33454 , n381447 );
nand ( n50787 , n50786 , n33465 );
and ( n50788 , n50787 , n381458 );
and ( n50789 , n33476 , n381463 );
and ( n50790 , n383147 , RI15b52f98_696);
nor ( n50791 , n50788 , n50789 , n50790 );
nand ( n50792 , n50785 , n50791 );
buf ( n50793 , n50792 );
buf ( n50794 , n382067 );
buf ( n50795 , n33382 );
or ( n50796 , n36937 , n48936 );
and ( n50797 , n36946 , n48939 );
not ( n50798 , RI15b4eee8_558);
or ( n50799 , n48948 , n50798 );
or ( n50800 , n39875 , n48953 );
or ( n50801 , n48946 , n36955 );
nand ( n50802 , n50799 , n50800 , n50801 );
nor ( n50803 , n50797 , n50802 );
nand ( n50804 , n50796 , n50803 );
buf ( n50805 , n50804 );
buf ( n50806 , n381707 );
not ( n50807 , RI15b5ffb8_1140);
not ( n50808 , n383601 );
or ( n50809 , n50807 , n50808 );
not ( n50810 , n32306 );
or ( n50811 , n33577 , n50810 );
nand ( n50812 , n50811 , n33584 );
not ( n50813 , n32301 );
and ( n50814 , n50812 , n50813 );
nor ( n50815 , n50813 , n32306 );
and ( n50816 , n40781 , n50815 );
and ( n50817 , n383607 , RI15b5e9b0_1093);
nor ( n50818 , n50814 , n50816 , n50817 );
nand ( n50819 , n50809 , n50818 );
buf ( n50820 , n50819 );
buf ( n50821 , n381021 );
buf ( n50822 , n21800 );
not ( n50823 , RI15b53448_706);
not ( n50824 , n32244 );
or ( n50825 , n50823 , n50824 );
and ( n50826 , n32247 , RI15b64a40_1299);
and ( n50827 , n32249 , RI15b5f8b0_1125);
nor ( n50828 , n50826 , n50827 );
nand ( n50829 , n50825 , n50828 );
buf ( n50830 , n50829 );
buf ( n50831 , n32672 );
buf ( n50832 , n20663 );
not ( n50833 , RI15b4a460_399);
not ( n50834 , n30908 );
or ( n50835 , n50833 , n50834 );
and ( n50836 , n22217 , n19740 );
buf ( n50837 , n19734 );
not ( n50838 , RI15b4a460_399);
and ( n50839 , n50837 , n50838 );
not ( n50840 , n50837 );
and ( n50841 , n50840 , RI15b4a460_399);
nor ( n50842 , n50839 , n50841 );
and ( n50843 , n20637 , n50842 );
nor ( n50844 , n50836 , n50843 );
and ( n50845 , n40215 , n50844 );
nand ( n50846 , n50835 , n50845 );
buf ( n50847 , n50846 );
buf ( n50848 , n22740 );
buf ( n50849 , n19655 );
buf ( n50850 , n386762 );
buf ( n50851 , n19653 );
buf ( n50852 , n32243 );
not ( n50853 , RI15b65b20_1335);
not ( n50854 , n35176 );
or ( n50855 , n50853 , n50854 );
nand ( n50856 , n35187 , RI15b48750_337);
not ( n50857 , n42818 );
and ( n50858 , n386554 , n50857 );
not ( n50859 , RI15b48750_337);
not ( n50860 , n35341 );
or ( n50861 , n50859 , n50860 );
or ( n50862 , n35341 , RI15b48750_337);
nand ( n50863 , n50861 , n50862 );
and ( n50864 , n50599 , n50863 );
nor ( n50865 , n50858 , n50864 );
and ( n50866 , n36927 , n50856 , n50865 );
nand ( n50867 , n50855 , n50866 );
buf ( n50868 , n50867 );
buf ( n50869 , n382052 );
buf ( n50870 , n22343 );
or ( n50871 , n380968 , n36121 );
and ( n50872 , n380986 , n36123 );
or ( n50873 , n36132 , n20341 );
or ( n50874 , n380994 , n36139 );
or ( n50875 , n36130 , n380996 );
nand ( n50876 , n50873 , n50874 , n50875 );
nor ( n50877 , n50872 , n50876 );
nand ( n50878 , n50871 , n50877 );
buf ( n50879 , n50878 );
buf ( n50880 , n379403 );
buf ( n50881 , n18226 );
and ( n50882 , n38047 , RI15b53cb8_724);
and ( n50883 , n35213 , RI15b661b0_1349);
nor ( n50884 , n50882 , n50883 );
not ( n50885 , n50884 );
buf ( n50886 , n50885 );
buf ( n50887 , n22740 );
buf ( n50888 , n19655 );
or ( n50889 , n35333 , n34935 );
and ( n50890 , n35335 , RI15b660c0_1347);
not ( n50891 , n34935 );
not ( n50892 , n35356 );
or ( n50893 , n50891 , n50892 );
or ( n50894 , n35356 , n34935 );
nand ( n50895 , n50893 , n50894 );
and ( n50896 , n50895 , n35363 );
nor ( n50897 , n44278 , n35456 );
nor ( n50898 , n50890 , n50896 , n50897 );
nand ( n50899 , n50889 , n50898 , n48639 );
buf ( n50900 , n50899 );
buf ( n50901 , n381490 );
buf ( n50902 , n380906 );
buf ( n50903 , n381081 );
nand ( n50904 , n32397 , RI15b532e0_703);
not ( n50905 , n48846 );
not ( n50906 , n44645 );
or ( n50907 , n50905 , n50906 );
nand ( n50908 , n50907 , n381450 );
and ( n50909 , n50908 , n48858 );
and ( n50910 , n381461 , n48860 );
nor ( n50911 , n50909 , n50910 );
nand ( n50912 , n386636 , n50904 , n50911 );
buf ( n50913 , n50912 );
buf ( n50914 , n35649 );
not ( n50915 , n35983 );
not ( n50916 , n380703 );
or ( n50917 , n50915 , n50916 );
and ( n50918 , n380719 , n35987 );
not ( n50919 , RI15b5bbc0_995);
or ( n50920 , n35996 , n50919 );
or ( n50921 , n37542 , n36003 );
or ( n50922 , n35994 , n380790 );
nand ( n50923 , n50920 , n50921 , n50922 );
nor ( n50924 , n50918 , n50923 );
nand ( n50925 , n50917 , n50924 );
buf ( n50926 , n50925 );
buf ( n50927 , n21800 );
or ( n50928 , n386588 , n381530 );
and ( n50929 , n386600 , n381528 );
not ( n50930 , RI15b5bcb0_997);
or ( n50931 , n381544 , n50930 );
or ( n50932 , n34706 , n381557 );
or ( n50933 , n381542 , n386627 );
nand ( n50934 , n50931 , n50932 , n50933 );
nor ( n50935 , n50929 , n50934 );
nand ( n50936 , n50928 , n50935 );
buf ( n50937 , n50936 );
buf ( n50938 , n383174 );
or ( n50939 , n42969 , n47758 );
not ( n50940 , n40056 );
not ( n50941 , n38897 );
or ( n50942 , n50940 , n50941 );
nand ( n50943 , n50942 , n381450 );
and ( n50944 , n50943 , n40039 );
nor ( n50945 , n40056 , n40039 );
and ( n50946 , n381461 , n50945 );
nor ( n50947 , n50944 , n50946 );
and ( n50948 , n47761 , n50947 );
nand ( n50949 , n381486 , RI15b531f0_701);
nand ( n50950 , n50939 , n50948 , n50949 );
buf ( n50951 , n50950 );
buf ( n50952 , n381566 );
not ( n50953 , n21862 );
nor ( n50954 , n50953 , n21870 );
and ( n50955 , n21802 , n50954 );
not ( n50956 , n21963 );
not ( n50957 , n21949 );
or ( n50958 , n50956 , n50957 );
nand ( n50959 , n50958 , n21979 );
and ( n50960 , n50959 , RI15b55d10_793);
and ( n50961 , n18150 , RI15b57b10_857);
or ( n50962 , n21982 , n21963 , RI15b55d10_793);
and ( n50963 , n21933 , RI15b57b10_857);
not ( n50964 , n21933 );
and ( n50965 , n50964 , n21934 );
nor ( n50966 , n50963 , n50965 );
or ( n50967 , n21922 , n50966 );
nand ( n50968 , n50962 , n50967 );
nor ( n50969 , n50960 , n50961 , n50968 );
or ( n50970 , n50969 , n18078 );
and ( n50971 , n18177 , RI15b57b10_857);
and ( n50972 , n18219 , RI15b56c10_825);
nor ( n50973 , n50971 , n50972 , n21751 );
nand ( n50974 , n50970 , n50973 );
nor ( n50975 , n50955 , n50974 );
nand ( n50976 , n50953 , n17507 );
not ( n50977 , n50976 );
not ( n50978 , n17565 );
or ( n50979 , n50977 , n50978 );
nand ( n50980 , n50979 , n21870 );
nand ( n50981 , n50975 , n50980 );
buf ( n50982 , n50981 );
buf ( n50983 , n381707 );
buf ( n50984 , n19651 );
not ( n50985 , n22551 );
and ( n50986 , n50985 , n42548 );
or ( n50987 , n381828 , n17520 , RI15b57390_841);
and ( n50988 , n17520 , n384113 );
nor ( n50989 , n50988 , n21791 );
or ( n50990 , n50989 , n17521 );
nand ( n50991 , n50987 , n50990 );
nor ( n50992 , n50986 , n50991 );
nand ( n50993 , n46330 , n50992 );
buf ( n50994 , n50993 );
buf ( n50995 , n382065 );
buf ( n50996 , n19653 );
buf ( n50997 , n22740 );
buf ( n50998 , n386762 );
not ( n50999 , n382044 );
buf ( n51000 , n35351 );
and ( n51001 , n35363 , n51000 );
nor ( n51002 , n51001 , n35186 );
not ( n51003 , n51002 );
nand ( n51004 , n51003 , RI15b48b10_345);
and ( n51005 , n32747 , RI15b42af8_140);
and ( n51006 , n32753 , RI15b41838_100);
and ( n51007 , n32755 , RI15b41bf8_108);
nor ( n51008 , n51006 , n51007 );
and ( n51009 , n32759 , RI15b410b8_84);
and ( n51010 , n32762 , RI15b41478_92);
nor ( n51011 , n51009 , n51010 );
and ( n51012 , n32766 , RI15b43638_164);
and ( n51013 , n32768 , RI15b43278_156);
nor ( n51014 , n51012 , n51013 );
and ( n51015 , n32771 , RI15b439f8_172);
and ( n51016 , n32773 , RI15b42eb8_148);
nor ( n51017 , n51015 , n51016 );
nand ( n51018 , n51008 , n51011 , n51014 , n51017 );
and ( n51019 , n45352 , n51018 );
and ( n51020 , n32781 , RI15b40578_60);
nor ( n51021 , n51005 , n51019 , n51020 );
and ( n51022 , n32785 , RI15b42738_132);
and ( n51023 , n32787 , RI15b42378_124);
nor ( n51024 , n51022 , n51023 );
and ( n51025 , n32792 , RI15b401b8_52);
and ( n51026 , n32794 , RI15b41fb8_116);
nor ( n51027 , n51025 , n51026 );
and ( n51028 , n32797 , RI15b40938_68);
and ( n51029 , n32800 , RI15b40cf8_76);
nor ( n51030 , n51028 , n51029 );
nand ( n51031 , n51021 , n51024 , n51027 , n51030 );
nand ( n51032 , n51031 , n48997 );
and ( n51033 , n35335 , RI15b65ee0_1343);
not ( n51034 , RI15b48a98_344);
or ( n51035 , n51000 , n51034 , RI15b48b10_345);
or ( n51036 , n381950 , RI15b48a98_344);
nand ( n51037 , n51035 , n51036 );
and ( n51038 , n48988 , n51037 );
nor ( n51039 , n51033 , n51038 );
nand ( n51040 , n50999 , n51004 , n51032 , n51039 );
buf ( n51041 , n51040 );
or ( n51042 , n381015 , n22050 );
nand ( n51043 , n35525 , RI15b53e98_728);
nand ( n51044 , n51042 , n51043 );
buf ( n51045 , n51044 );
buf ( n51046 , n380942 );
not ( n51047 , n384058 );
not ( n51048 , n384726 );
or ( n51049 , n51047 , n51048 );
and ( n51050 , n384737 , n384169 );
or ( n51051 , n384182 , n17762 );
or ( n51052 , n39386 , n384190 );
or ( n51053 , n384180 , n384759 );
nand ( n51054 , n51051 , n51052 , n51053 );
nor ( n51055 , n51050 , n51054 );
nand ( n51056 , n51049 , n51055 );
buf ( n51057 , n51056 );
buf ( n51058 , n22402 );
buf ( n51059 , n22653 );
buf ( n51060 , n385112 );
not ( n51061 , n383930 );
not ( n51062 , n39366 );
or ( n51063 , n51061 , n51062 );
and ( n51064 , n384022 , RI15b62088_1210);
not ( n51065 , RI15b62088_1210);
not ( n51066 , n384037 );
or ( n51067 , n51065 , n51066 );
or ( n51068 , n384037 , RI15b62088_1210);
nand ( n51069 , n51067 , n51068 );
and ( n51070 , n384025 , n51069 );
nor ( n51071 , n51064 , n51070 );
nand ( n51072 , n51063 , n51071 );
buf ( n51073 , n51072 );
and ( n51074 , n22646 , RI15b45618_232);
and ( n51075 , n22648 , RI15b51a80_651);
nor ( n51076 , n51074 , n51075 );
not ( n51077 , n51076 );
buf ( n51078 , n51077 );
not ( n51079 , n35784 );
not ( n51080 , n380703 );
or ( n51081 , n51079 , n51080 );
and ( n51082 , n380719 , n35790 );
not ( n51083 , RI15b59dc0_931);
or ( n51084 , n35803 , n51083 );
or ( n51085 , n380782 , n35811 );
or ( n51086 , n35801 , n380790 );
nand ( n51087 , n51084 , n51085 , n51086 );
nor ( n51088 , n51082 , n51087 );
nand ( n51089 , n51081 , n51088 );
buf ( n51090 , n51089 );
or ( n51091 , n382679 , n382654 );
and ( n51092 , n48159 , n386669 );
or ( n51093 , n382691 , n383631 );
and ( n51094 , n382653 , RI15b550e0_767);
not ( n51095 , n382653 );
and ( n51096 , n51095 , n382654 );
nor ( n51097 , n51094 , n51096 );
or ( n51098 , n43699 , n51097 );
nand ( n51099 , n51093 , n51098 , n44873 );
nor ( n51100 , n51092 , n51099 );
nand ( n51101 , n51091 , n51100 );
buf ( n51102 , n51101 );
buf ( n51103 , n385197 );
buf ( n51104 , n22005 );
buf ( n51105 , n22343 );
buf ( n51106 , n32271 );
buf ( n51107 , n383613 );
not ( n51108 , n45106 );
not ( n51109 , n384122 );
or ( n51110 , n51108 , n51109 );
and ( n51111 , n384164 , n40470 );
or ( n51112 , n40480 , n20876 );
or ( n51113 , n33131 , n40485 );
or ( n51114 , n40478 , n384193 );
nand ( n51115 , n51112 , n51113 , n51114 );
nor ( n51116 , n51111 , n51115 );
nand ( n51117 , n51110 , n51116 );
buf ( n51118 , n51117 );
not ( n51119 , RI15b5f040_1107);
not ( n51120 , n384918 );
or ( n51121 , n51119 , n51120 );
and ( n51122 , n32275 , RI15b60d50_1169);
nand ( n51123 , n384906 , n383187 );
not ( n51124 , n51123 );
nor ( n51125 , n51122 , n51124 );
nand ( n51126 , n51121 , n51125 );
buf ( n51127 , n51126 );
buf ( n51128 , n387159 );
not ( n51129 , n38488 );
not ( n51130 , RI15b628f8_1228);
and ( n51131 , n51129 , n51130 );
not ( n51132 , n51129 );
and ( n51133 , n51132 , RI15b628f8_1228);
nor ( n51134 , n51131 , n51133 );
nand ( n51135 , n51134 , n384025 );
and ( n51136 , n384022 , RI15b628f8_1228);
and ( n51137 , n46086 , n386746 );
nor ( n51138 , n51136 , n51137 );
nand ( n51139 , n51135 , n51138 );
buf ( n51140 , n51139 );
buf ( n51141 , n379403 );
or ( n51142 , n36937 , n38825 );
and ( n51143 , n36946 , n38828 );
or ( n51144 , n38837 , n17813 );
or ( n51145 , n41326 , n38841 );
or ( n51146 , n38835 , n36955 );
nand ( n51147 , n51144 , n51145 , n51146 );
nor ( n51148 , n51143 , n51147 );
nand ( n51149 , n51142 , n51148 );
buf ( n51150 , n51149 );
buf ( n51151 , n22716 );
buf ( n51152 , n384199 );
buf ( n51153 , RI15b46ef0_285);
buf ( n51154 , n381006 );
and ( n51155 , n48600 , n37739 );
nor ( n51156 , n46076 , n51155 );
or ( n51157 , n51156 , n45125 );
nor ( n51158 , n46080 , n37739 );
and ( n51159 , n51158 , n45125 );
or ( n51160 , n38817 , n41343 );
or ( n51161 , n380539 , n31052 );
nand ( n51162 , n51160 , n51161 , n37800 );
nor ( n51163 , n51159 , n51162 );
nand ( n51164 , n51157 , n51163 );
buf ( n51165 , n51164 );
buf ( n51166 , n31979 );
or ( n51167 , n31006 , n36242 );
and ( n51168 , n31016 , n43075 );
or ( n51169 , n36250 , n20982 );
or ( n51170 , n40593 , n36254 );
or ( n51171 , n36248 , n31024 );
nand ( n51172 , n51169 , n51170 , n51171 );
nor ( n51173 , n51168 , n51172 );
nand ( n51174 , n51167 , n51173 );
buf ( n51175 , n51174 );
buf ( n51176 , n379895 );
or ( n51177 , n32926 , n32944 );
not ( n51178 , n382080 );
not ( n51179 , n32923 );
not ( n51180 , n51179 );
or ( n51181 , n51178 , n51180 );
nand ( n51182 , n51181 , n46996 );
nand ( n51183 , n51182 , n32944 );
not ( n51184 , n382513 );
not ( n51185 , n32932 );
not ( n51186 , n51185 );
not ( n51187 , n382502 );
or ( n51188 , n51186 , n51187 );
or ( n51189 , n382502 , n51185 );
nand ( n51190 , n51188 , n51189 );
and ( n51191 , n51184 , n51190 );
and ( n51192 , n382523 , RI15b4bea0_455);
and ( n51193 , n32975 , RI15b45ca8_246);
nor ( n51194 , n51191 , n51192 , n51193 );
nand ( n51195 , n51177 , n51183 , n51194 );
buf ( n51196 , n51195 );
buf ( n51197 , n22009 );
buf ( n51198 , n33250 );
buf ( n51199 , n381707 );
buf ( n51200 , n32676 );
buf ( n51201 , n386762 );
or ( n51202 , n34994 , n41015 );
nand ( n51203 , n51202 , n41032 );
nand ( n51204 , n51203 , n35108 );
nand ( n51205 , n41651 , n35119 );
nand ( n51206 , n41582 , RI15b460e0_255);
and ( n51207 , n35459 , n379840 );
and ( n51208 , n35461 , RI15b658c8_1330);
nor ( n51209 , n51207 , n51208 );
nand ( n51210 , n51204 , n51205 , n51206 , n51209 );
buf ( n51211 , n51210 );
buf ( n51212 , n379802 );
buf ( n51213 , n33250 );
buf ( n51214 , n381872 );
not ( n51215 , n33580 );
not ( n51216 , n37809 );
or ( n51217 , n51215 , n51216 );
nand ( n51218 , n51217 , n33584 );
nand ( n51219 , n51218 , n33567 );
nand ( n51220 , n37814 , n40781 );
nand ( n51221 , n383601 , RI15b60288_1146);
nand ( n51222 , n383607 , RI15b5ec80_1099);
nand ( n51223 , n51219 , n51220 , n51221 , n51222 );
buf ( n51224 , n51223 );
buf ( n51225 , n33250 );
not ( n51226 , n33597 );
not ( n51227 , n51226 );
not ( n51228 , n384726 );
or ( n51229 , n51227 , n51228 );
and ( n51230 , n35477 , n33600 );
not ( n51231 , RI15b4ec18_552);
or ( n51232 , n33609 , n51231 );
not ( n51233 , n35490 );
or ( n51234 , n51233 , n33615 );
or ( n51235 , n33607 , n384759 );
nand ( n51236 , n51232 , n51234 , n51235 );
nor ( n51237 , n51230 , n51236 );
nand ( n51238 , n51229 , n51237 );
buf ( n51239 , n51238 );
buf ( n51240 , n384218 );
buf ( n51241 , n381872 );
not ( n51242 , RI15b52bd8_688);
not ( n51243 , n381484 );
or ( n51244 , n51242 , n51243 );
and ( n51245 , n41853 , RI15b548e8_750);
nor ( n51246 , n51245 , n41858 );
nand ( n51247 , n51244 , n51246 );
buf ( n51248 , n51247 );
not ( n51249 , n36276 );
not ( n51250 , n381507 );
or ( n51251 , n51249 , n51250 );
and ( n51252 , n381524 , n36282 );
not ( n51253 , RI15b5c2c8_1010);
or ( n51254 , n36291 , n51253 );
or ( n51255 , n32478 , n36296 );
or ( n51256 , n36289 , n381560 );
nand ( n51257 , n51254 , n51255 , n51256 );
nor ( n51258 , n51252 , n51257 );
nand ( n51259 , n51251 , n51258 );
buf ( n51260 , n51259 );
buf ( n51261 , n22788 );
buf ( n51262 , n386762 );
buf ( n51263 , n381004 );
buf ( n51264 , n22406 );
buf ( n51265 , n387159 );
buf ( n51266 , n18226 );
or ( n51267 , n22102 , n37663 );
and ( n51268 , n22203 , n37666 );
not ( n51269 , RI15b42a08_138);
or ( n51270 , n37675 , n51269 );
or ( n51271 , n22293 , n37679 );
or ( n51272 , n37673 , n22299 );
nand ( n51273 , n51270 , n51271 , n51272 );
nor ( n51274 , n51268 , n51273 );
nand ( n51275 , n51267 , n51274 );
buf ( n51276 , n51275 );
buf ( n51277 , n380906 );
buf ( n51278 , n31030 );
not ( n51279 , n42706 );
nand ( n51280 , n42708 , n51279 );
nor ( n51281 , n51280 , n382079 );
or ( n51282 , n51281 , n32958 );
nand ( n51283 , n51282 , n32016 );
nor ( n51284 , n32924 , n32016 );
and ( n51285 , n51280 , n51284 );
not ( n51286 , n32041 );
not ( n51287 , n382335 );
and ( n51288 , n51286 , n51287 );
and ( n51289 , n32041 , n382335 );
nor ( n51290 , n51288 , n51289 );
or ( n51291 , n382513 , n51290 );
and ( n51292 , n382523 , RI15b4b798_440);
and ( n51293 , n32974 , RI15b455a0_231);
nor ( n51294 , n51292 , n51293 );
nand ( n51295 , n51291 , n51294 );
nor ( n51296 , n51285 , n51295 );
nand ( n51297 , n51283 , n51296 );
buf ( n51298 , n51297 );
buf ( n51299 , n381081 );
buf ( n51300 , n380940 );
buf ( n51301 , n379403 );
buf ( n51302 , n43349 );
buf ( n51303 , n382052 );
or ( n51304 , n384961 , n37663 );
and ( n51305 , n384983 , n37666 );
or ( n51306 , n37675 , n385412 );
or ( n51307 , n22022 , n37679 );
or ( n51308 , n37673 , n384988 );
nand ( n51309 , n51306 , n51307 , n51308 );
nor ( n51310 , n51305 , n51309 );
nand ( n51311 , n51304 , n51310 );
buf ( n51312 , n51311 );
buf ( n51313 , n383174 );
buf ( n51314 , n20663 );
buf ( n51315 , n381004 );
not ( n51316 , n386514 );
or ( n51317 , n51316 , n386099 );
and ( n51318 , n386540 , RI15b43bd8_176);
and ( n51319 , n386549 , n385751 );
and ( n51320 , n386556 , n386099 );
nor ( n51321 , n51318 , n51319 , n51320 );
not ( n51322 , n32230 );
nand ( n51323 , n51317 , n51321 , n51322 );
buf ( n51324 , n51323 );
buf ( n51325 , n379844 );
buf ( n51326 , n32271 );
or ( n51327 , n381015 , n22032 );
nand ( n51328 , n35327 , RI15b53970_717);
nand ( n51329 , n51327 , n51328 );
buf ( n51330 , n51329 );
buf ( n51331 , n380906 );
buf ( n51332 , n22716 );
not ( n51333 , n48980 );
or ( n51334 , n51333 , n35027 );
not ( n51335 , n48974 );
and ( n51336 , n51335 , n35027 );
not ( n51337 , n51335 );
and ( n51338 , n51337 , RI15b49038_356);
nor ( n51339 , n51336 , n51338 );
and ( n51340 , n51339 , n48968 );
not ( n51341 , n37258 );
not ( n51342 , n37230 );
or ( n51343 , n51341 , n51342 );
or ( n51344 , n37230 , n37258 );
nand ( n51345 , n51343 , n51344 );
not ( n51346 , n51345 );
not ( n51347 , n386554 );
or ( n51348 , n51346 , n51347 );
not ( n51349 , RI15b66408_1354);
or ( n51350 , n386547 , n51349 );
nand ( n51351 , n51348 , n51350 );
nor ( n51352 , n51340 , n51351 );
nand ( n51353 , n51334 , n51352 , n41659 );
buf ( n51354 , n51353 );
buf ( n51355 , n384700 );
buf ( n51356 , n382073 );
buf ( n51357 , n31979 );
not ( n51358 , n35473 );
not ( n51359 , n384122 );
or ( n51360 , n51358 , n51359 );
and ( n51361 , n384164 , n35479 );
or ( n51362 , n35488 , n20852 );
or ( n51363 , n46471 , n35497 );
or ( n51364 , n35486 , n384193 );
nand ( n51365 , n51362 , n51363 , n51364 );
nor ( n51366 , n51361 , n51365 );
nand ( n51367 , n51360 , n51366 );
buf ( n51368 , n51367 );
or ( n51369 , n31091 , n31061 );
not ( n51370 , n31790 );
not ( n51371 , n37640 );
and ( n51372 , n51370 , n51371 );
and ( n51373 , n35507 , n18590 );
and ( n51374 , n31060 , n31061 );
not ( n51375 , n31060 );
and ( n51376 , n51375 , RI15b60e40_1171);
nor ( n51377 , n51374 , n51376 );
and ( n51378 , n31078 , n51377 );
nor ( n51379 , n51372 , n51373 , n51378 );
nand ( n51380 , n51369 , n51379 );
buf ( n51381 , n51380 );
buf ( n51382 , n22009 );
buf ( n51383 , n32981 );
buf ( n51384 , RI15b47328_294);
buf ( n51385 , n385195 );
not ( n51386 , n47644 );
not ( n51387 , n37629 );
or ( n51388 , n51386 , n51387 );
and ( n51389 , n37637 , n47649 );
or ( n51390 , n47658 , n18581 );
or ( n51391 , n50080 , n47663 );
or ( n51392 , n47656 , n37646 );
nand ( n51393 , n51390 , n51391 , n51392 );
nor ( n51394 , n51389 , n51393 );
nand ( n51395 , n51388 , n51394 );
buf ( n51396 , n51395 );
buf ( n51397 , n385112 );
buf ( n51398 , n32672 );
or ( n51399 , n22585 , n380001 );
not ( n51400 , n49905 );
or ( n51401 , n51400 , n48429 );
not ( n51402 , n379977 );
and ( n51403 , n51402 , RI15b56238_804);
not ( n51404 , n51402 );
and ( n51405 , n51404 , n22585 );
nor ( n51406 , n51403 , n51405 );
or ( n51407 , n379948 , n51406 );
nand ( n51408 , n51399 , n51401 , n51407 );
buf ( n51409 , n51408 );
buf ( n51410 , n32676 );
not ( n51411 , RI15b53358_704);
not ( n51412 , n383170 );
or ( n51413 , n51411 , n51412 );
and ( n51414 , n33453 , RI15b548e8_750);
and ( n51415 , n383147 , RI15b52bd8_688);
nor ( n51416 , n51414 , n51415 );
nand ( n51417 , n51413 , n51416 );
buf ( n51418 , n51417 );
buf ( n51419 , n35649 );
not ( n51420 , n35983 );
not ( n51421 , n381507 );
or ( n51422 , n51420 , n51421 );
and ( n51423 , n381524 , n35987 );
not ( n51424 , RI15b5bb48_994);
or ( n51425 , n35996 , n51424 );
or ( n51426 , n38012 , n36003 );
or ( n51427 , n35994 , n381560 );
nand ( n51428 , n51425 , n51426 , n51427 );
nor ( n51429 , n51423 , n51428 );
nand ( n51430 , n51422 , n51429 );
buf ( n51431 , n51430 );
or ( n51432 , n36266 , n37443 );
nand ( n51433 , n36269 , RI15b54ac8_754);
and ( n51434 , n37445 , n51433 );
nand ( n51435 , n381486 , RI15b52db8_692);
nand ( n51436 , n51432 , n51434 , n51435 );
buf ( n51437 , n51436 );
not ( n51438 , n36276 );
not ( n51439 , n37629 );
or ( n51440 , n51438 , n51439 );
and ( n51441 , n37637 , n36282 );
not ( n51442 , RI15b5c0e8_1006);
or ( n51443 , n36291 , n51442 );
or ( n51444 , n43001 , n36296 );
or ( n51445 , n36289 , n37646 );
nand ( n51446 , n51443 , n51444 , n51445 );
nor ( n51447 , n51441 , n51446 );
nand ( n51448 , n51440 , n51447 );
buf ( n51449 , n51448 );
buf ( n51450 , n31719 );
buf ( n51451 , n22404 );
buf ( n51452 , n35649 );
not ( n51453 , RI15b55e78_796);
not ( n51454 , n380000 );
or ( n51455 , n51453 , n51454 );
and ( n51456 , n381636 , RI15b4eba0_551);
and ( n51457 , n381639 , RI15b4e7e0_543);
nor ( n51458 , n51456 , n51457 );
and ( n51459 , n381643 , RI15b4ef60_559);
and ( n51460 , n41896 , RI15b4dca0_519);
and ( n51461 , n382852 , RI15b4fe60_591);
nor ( n51462 , n51460 , n51461 );
and ( n51463 , n381661 , RI15b4faa0_583);
and ( n51464 , n381663 , RI15b4f320_567);
nor ( n51465 , n51463 , n51464 );
and ( n51466 , n381667 , RI15b4d520_503);
and ( n51467 , n381669 , RI15b4d8e0_511);
nor ( n51468 , n51466 , n51467 );
and ( n51469 , n381672 , RI15b4e060_527);
and ( n51470 , n381674 , RI15b4f6e0_575);
nor ( n51471 , n51469 , n51470 );
nand ( n51472 , n51462 , n51465 , n51468 , n51471 );
and ( n51473 , n38323 , n51472 );
and ( n51474 , n381680 , RI15b4c9e0_479);
nor ( n51475 , n51459 , n51473 , n51474 );
and ( n51476 , n381684 , RI15b4c620_471);
and ( n51477 , n381686 , RI15b4e420_535);
nor ( n51478 , n51476 , n51477 );
and ( n51479 , n381689 , RI15b4cda0_487);
and ( n51480 , n381691 , RI15b4d160_495);
nor ( n51481 , n51479 , n51480 );
nand ( n51482 , n51458 , n51475 , n51478 , n51481 );
and ( n51483 , n51482 , n381696 );
not ( n51484 , RI15b55e78_796);
not ( n51485 , n379966 );
not ( n51486 , n51485 );
or ( n51487 , n51484 , n51486 );
or ( n51488 , n51485 , RI15b55e78_796);
nand ( n51489 , n51487 , n51488 );
and ( n51490 , n379949 , n51489 );
nor ( n51491 , n51483 , n51490 );
nand ( n51492 , n51455 , n51491 );
buf ( n51493 , n51492 );
buf ( n51494 , n382049 );
buf ( n51495 , n381006 );
not ( n51496 , n381570 );
not ( n51497 , n37629 );
or ( n51498 , n51496 , n51497 );
and ( n51499 , n37637 , n381599 );
or ( n51500 , n381609 , n18997 );
or ( n51501 , n43001 , n381619 );
or ( n51502 , n381607 , n37646 );
nand ( n51503 , n51500 , n51501 , n51502 );
nor ( n51504 , n51499 , n51503 );
nand ( n51505 , n51498 , n51504 );
buf ( n51506 , n51505 );
buf ( n51507 , n382052 );
not ( n51508 , n44317 );
and ( n51509 , n51508 , n34931 );
nor ( n51510 , n51509 , n35114 );
or ( n51511 , n51510 , n35077 );
and ( n51512 , n35118 , n44322 );
and ( n51513 , n20631 , RI15b46248_258);
nor ( n51514 , n51512 , n51513 );
nand ( n51515 , n385213 , RI15b47850_305);
nand ( n51516 , n51511 , n51514 , n51515 );
buf ( n51517 , n51516 );
buf ( n51518 , n35651 );
buf ( n51519 , n32255 );
buf ( n51520 , n382537 );
or ( n51521 , n31053 , n380364 );
not ( n51522 , n384901 );
nand ( n51523 , n384907 , n51522 );
and ( n51524 , n46211 , RI15b61278_1180);
and ( n51525 , n45920 , n31125 );
nor ( n51526 , n31073 , RI15b61278_1180);
and ( n51527 , n40636 , n51526 );
nor ( n51528 , n51524 , n51525 , n51527 );
nand ( n51529 , n51521 , n51523 , n51528 );
buf ( n51530 , n51529 );
buf ( n51531 , n30992 );
or ( n51532 , n36937 , n31151 );
and ( n51533 , n36946 , n31164 );
or ( n51534 , n31175 , n17790 );
or ( n51535 , n36952 , n31182 );
or ( n51536 , n31173 , n36955 );
nand ( n51537 , n51534 , n51535 , n51536 );
nor ( n51538 , n51533 , n51537 );
nand ( n51539 , n51532 , n51538 );
buf ( n51540 , n51539 );
buf ( n51541 , n381006 );
buf ( n51542 , n382073 );
buf ( n51543 , n32255 );
not ( n51544 , n381494 );
not ( n51545 , n37629 );
or ( n51546 , n51544 , n51545 );
and ( n51547 , n37637 , n381528 );
not ( n51548 , RI15b5bd28_998);
or ( n51549 , n381544 , n51548 );
or ( n51550 , n50208 , n381557 );
or ( n51551 , n381542 , n37646 );
nand ( n51552 , n51549 , n51550 , n51551 );
nor ( n51553 , n51547 , n51552 );
nand ( n51554 , n51546 , n51553 );
buf ( n51555 , n51554 );
buf ( n51556 , n384203 );
or ( n51557 , n381407 , n41886 );
or ( n51558 , n50743 , n40055 );
nand ( n51559 , n51558 , n381450 );
and ( n51560 , n51559 , n40046 );
and ( n51561 , n381461 , n50222 );
nor ( n51562 , n51560 , n51561 );
and ( n51563 , n41889 , n51562 );
nand ( n51564 , n381486 , RI15b53178_700);
nand ( n51565 , n51557 , n51563 , n51564 );
buf ( n51566 , n51565 );
not ( n51567 , n22515 );
and ( n51568 , n379897 , n22509 , n51567 );
or ( n51569 , n33298 , n33306 );
buf ( n51570 , n22584 );
and ( n51571 , n51570 , n18086 );
nor ( n51572 , n51571 , n18103 );
or ( n51573 , n22585 , n51572 );
not ( n51574 , n51570 );
and ( n51575 , n51574 , n18198 , n22585 );
or ( n51576 , n18189 , n22617 , RI15b58038_868);
or ( n51577 , n18218 , n22511 );
nand ( n51578 , n51576 , n51577 );
nor ( n51579 , n51575 , n51578 );
nand ( n51580 , n51569 , n51573 , n51579 );
nor ( n51581 , n51568 , n51580 );
not ( n51582 , n17507 );
not ( n51583 , n22509 );
not ( n51584 , n51583 );
or ( n51585 , n51582 , n51584 );
nand ( n51586 , n51585 , n17565 );
nand ( n51587 , n51586 , n22515 );
nand ( n51588 , n51581 , n51587 );
buf ( n51589 , n51588 );
and ( n51590 , n21788 , RI15b56e68_830);
and ( n51591 , n21909 , n33324 );
not ( n51592 , n21903 );
and ( n51593 , n51592 , n17543 );
not ( n51594 , n51592 );
and ( n51595 , n51594 , RI15b56e68_830);
nor ( n51596 , n51593 , n51595 );
and ( n51597 , n51596 , n384127 );
nor ( n51598 , n51590 , n51591 , n51597 );
nand ( n51599 , n36175 , n51598 );
buf ( n51600 , n51599 );
buf ( n51601 , n380865 );
buf ( n51602 , n379893 );
buf ( n51603 , n380906 );
buf ( n51604 , n383613 );
buf ( n51605 , n383174 );
not ( n51606 , RI15b53bc8_722);
not ( n51607 , n383170 );
or ( n51608 , n51606 , n51607 );
or ( n51609 , n383152 , n383110 );
nand ( n51610 , n51609 , n383157 );
and ( n51611 , n51610 , n383102 );
and ( n51612 , n36348 , n383143 );
and ( n51613 , n383147 , RI15b525c0_675);
nor ( n51614 , n51611 , n51612 , n51613 );
nand ( n51615 , n51608 , n51614 );
buf ( n51616 , n51615 );
not ( n51617 , n35145 );
not ( n51618 , n33400 );
or ( n51619 , n51617 , n51618 );
and ( n51620 , n33415 , n35150 );
or ( n51621 , n35160 , n18480 );
or ( n51622 , n36293 , n35166 );
or ( n51623 , n35158 , n33443 );
nand ( n51624 , n51621 , n51622 , n51623 );
nor ( n51625 , n51620 , n51624 );
nand ( n51626 , n51619 , n51625 );
buf ( n51627 , n51626 );
buf ( n51628 , n385197 );
buf ( n51629 , n379895 );
and ( n51630 , n34812 , RI15b63f78_1276);
buf ( n51631 , n386969 );
not ( n51632 , n51631 );
not ( n51633 , n38093 );
or ( n51634 , n51632 , n51633 );
nand ( n51635 , n51634 , n34823 );
and ( n51636 , n51635 , RI15b62178_1212);
or ( n51637 , n34826 , n51631 , RI15b62178_1212);
not ( n51638 , n387030 );
not ( n51639 , RI15b63f78_1276);
and ( n51640 , n51638 , n51639 );
and ( n51641 , n387030 , RI15b63f78_1276);
nor ( n51642 , n51640 , n51641 );
or ( n51643 , n34833 , n51642 );
nand ( n51644 , n51637 , n51643 );
nor ( n51645 , n51630 , n51636 , n51644 );
or ( n51646 , n51645 , n19200 );
not ( n51647 , n386825 );
not ( n51648 , n51647 );
not ( n51649 , n22473 );
and ( n51650 , n51648 , n51649 );
nor ( n51651 , n51650 , n38114 );
or ( n51652 , n386831 , n51651 );
and ( n51653 , n38117 , n51647 , n386831 );
or ( n51654 , n22424 , n379573 );
or ( n51655 , n383446 , n19598 );
nand ( n51656 , n51654 , n51655 , n19512 );
nor ( n51657 , n51653 , n51656 );
nand ( n51658 , n51646 , n51652 , n51657 );
buf ( n51659 , n51658 );
buf ( n51660 , n32672 );
not ( n51661 , n20637 );
not ( n51662 , n19709 );
or ( n51663 , n51661 , n51662 );
nand ( n51664 , n51663 , n34798 );
and ( n51665 , n51664 , RI15b4af28_422);
or ( n51666 , n34801 , n19709 , RI15b4af28_422);
not ( n51667 , n19715 );
or ( n51668 , n51667 , n22216 );
nand ( n51669 , n51666 , n51668 );
nor ( n51670 , n51665 , n51669 );
nand ( n51671 , n46657 , n51670 );
buf ( n51672 , n51671 );
buf ( n51673 , n22404 );
buf ( n51674 , n386563 );
buf ( n51675 , RI15b5d948_1058);
and ( n51676 , n385164 , RI15b508b0_613);
or ( n51677 , n36693 , n21723 );
or ( n51678 , n20696 , n385170 );
or ( n51679 , n21382 , n385178 );
nand ( n51680 , n51677 , n51678 , n51679 );
nor ( n51681 , n51676 , n51680 );
nand ( n51682 , n42546 , n51681 );
buf ( n51683 , n51682 );
buf ( n51684 , n385195 );
buf ( n51685 , n382069 );
not ( n51686 , n47923 );
nor ( n51687 , n47903 , n51686 );
nand ( n51688 , n47916 , n39813 );
or ( n51689 , n51687 , n51688 );
not ( n51690 , n47947 );
nand ( n51691 , n47915 , n51690 );
nor ( n51692 , n47903 , n51691 );
buf ( n51693 , n44379 );
nand ( n51694 , n51693 , n379785 );
not ( n51695 , n51694 );
not ( n51696 , n36494 );
or ( n51697 , n51695 , n51696 );
buf ( n51698 , n44380 );
not ( n51699 , n51698 );
nand ( n51700 , n51697 , n51699 );
not ( n51701 , n51700 );
nor ( n51702 , n51692 , n51701 );
buf ( n51703 , n34249 );
buf ( n51704 , n51693 );
not ( n51705 , n51698 );
nor ( n51706 , n51704 , n51705 );
and ( n51707 , n51703 , n51706 );
and ( n51708 , n379783 , RI15b647e8_1294);
and ( n51709 , n34651 , RI15b5e5f0_1085);
nor ( n51710 , n51708 , n51709 );
not ( n51711 , n51710 );
nor ( n51712 , n51707 , n51711 );
nand ( n51713 , n51689 , n51702 , n51712 );
buf ( n51714 , n51713 );
buf ( n51715 , n22788 );
not ( n51716 , n32629 );
not ( n51717 , n384537 );
and ( n51718 , n51716 , n51717 );
not ( n51719 , n51716 );
and ( n51720 , n51719 , n384537 );
nor ( n51721 , n51718 , n51720 );
and ( n51722 , n51721 , n31960 );
not ( n51723 , n384461 );
not ( n51724 , n51723 );
not ( n51725 , n32644 );
or ( n51726 , n51724 , n51725 );
or ( n51727 , n32644 , n51723 );
nand ( n51728 , n51726 , n51727 );
not ( n51729 , n42099 );
nand ( n51730 , n51728 , n51729 );
and ( n51731 , n384360 , n384370 );
nor ( n51732 , n51731 , n384371 );
not ( n51733 , n51732 );
and ( n51734 , n51733 , n31921 );
and ( n51735 , n19513 , RI15b64428_1286);
nor ( n51736 , n51734 , n51735 );
nand ( n51737 , n51730 , n51736 );
nor ( n51738 , n51722 , n51737 );
and ( n51739 , n31792 , n384537 );
not ( n51740 , n384370 );
or ( n51741 , n51740 , n46430 );
or ( n51742 , n31771 , n384367 );
or ( n51743 , n51723 , n31779 );
nand ( n51744 , n51741 , n51742 , n51743 );
nor ( n51745 , n51739 , n51744 );
nand ( n51746 , n51738 , n51745 );
buf ( n51747 , n51746 );
buf ( n51748 , n32672 );
not ( n51749 , n39643 );
not ( n51750 , n51749 );
not ( n51751 , n39626 );
or ( n51752 , n51750 , n51751 );
not ( n51753 , n39643 );
or ( n51754 , n39626 , n51753 );
nand ( n51755 , n51752 , n51754 );
nand ( n51756 , n51755 , n31602 );
not ( n51757 , n379391 );
buf ( n51758 , n39669 );
not ( n51759 , n51758 );
or ( n51760 , n51757 , n51759 );
nand ( n51761 , n51760 , n31700 );
and ( n51762 , n51761 , n31686 );
or ( n51763 , n51758 , n39678 , n31686 );
and ( n51764 , n379394 , RI15b58308_874);
and ( n51765 , n39683 , RI15b52110_665);
nor ( n51766 , n51764 , n51765 );
nand ( n51767 , n51763 , n51766 );
nor ( n51768 , n51762 , n51767 );
nand ( n51769 , n51756 , n51768 );
buf ( n51770 , n51769 );
or ( n51771 , n37626 , n383436 );
nand ( n51772 , n51771 , n32581 );
and ( n51773 , n51772 , RI15b632d0_1249);
not ( n51774 , n383436 );
or ( n51775 , n384652 , n51774 , RI15b632d0_1249);
or ( n51776 , n386870 , n22775 );
nand ( n51777 , n51775 , n51776 );
nor ( n51778 , n51773 , n51777 );
nand ( n51779 , n37604 , n51778 );
buf ( n51780 , n51779 );
buf ( n51781 , n32981 );
buf ( n51782 , n382537 );
or ( n51783 , n48368 , n382125 );
not ( n51784 , n31806 );
buf ( n51785 , n19987 );
not ( n51786 , n51785 );
or ( n51787 , n51784 , n51786 );
nand ( n51788 , n51787 , n380875 );
nand ( n51789 , n51788 , RI15b49dd0_385);
not ( n51790 , n51785 );
and ( n51791 , n51790 , n32511 , n19988 );
or ( n51792 , n22354 , n48359 , RI15b4bbd0_449);
or ( n51793 , n22390 , n19866 );
nand ( n51794 , n51792 , n51793 );
nor ( n51795 , n51791 , n51794 );
nand ( n51796 , n51789 , n51795 );
buf ( n51797 , n19861 );
not ( n51798 , n19868 );
nor ( n51799 , n51797 , n35305 , n51798 );
nor ( n51800 , n51796 , n51799 );
not ( n51801 , n51797 );
nor ( n51802 , n51801 , n35293 );
or ( n51803 , n51802 , n38940 );
nand ( n51804 , n51803 , n51798 );
nand ( n51805 , n51783 , n51800 , n51804 );
buf ( n51806 , n51805 );
buf ( n51807 , n384700 );
buf ( n51808 , n381872 );
not ( n51809 , n39793 );
not ( n51810 , n51809 );
not ( n51811 , n39798 );
or ( n51812 , n51810 , n51811 );
not ( n51813 , n39823 );
nand ( n51814 , n51812 , n51813 );
nor ( n51815 , n39822 , n39794 );
nand ( n51816 , n36502 , n51815 );
buf ( n51817 , n39805 );
not ( n51818 , n51817 );
and ( n51819 , n51818 , n39803 );
not ( n51820 , n51818 );
and ( n51821 , n51820 , n34488 );
nor ( n51822 , n51819 , n51821 );
and ( n51823 , n51822 , n34646 );
not ( n51824 , RI15b5dee8_1070);
not ( n51825 , n34651 );
or ( n51826 , n51824 , n51825 );
or ( n51827 , n36518 , n379612 );
nand ( n51828 , n51826 , n51827 );
nor ( n51829 , n51823 , n51828 );
nand ( n51830 , n51814 , n51816 , n51829 );
buf ( n51831 , n51830 );
buf ( n51832 , n383498 );
not ( n51833 , n18077 );
not ( n51834 , n40863 );
or ( n51835 , n51833 , n51834 );
and ( n51836 , n39220 , RI15b50fb8_628);
and ( n51837 , n383915 , n18215 );
nor ( n51838 , n51836 , n51837 );
nand ( n51839 , n51835 , n51838 );
buf ( n51840 , n51839 );
buf ( n51841 , n379802 );
buf ( n51842 , n22479 );
buf ( n51843 , n383174 );
buf ( n51844 , n381021 );
buf ( n51845 , n381081 );
not ( n51846 , n383421 );
not ( n51847 , n51846 );
not ( n51848 , n381572 );
or ( n51849 , n51847 , n51848 );
nand ( n51850 , n51849 , n384642 );
nand ( n51851 , n51850 , RI15b63690_1257);
and ( n51852 , n384655 , n383421 , n386774 );
and ( n51853 , n386778 , n19630 );
nor ( n51854 , n51852 , n51853 );
nand ( n51855 , n31744 , n51851 , n51854 );
buf ( n51856 , n51855 );
not ( n51857 , n38988 );
buf ( n51858 , n19808 );
not ( n51859 , n51858 );
or ( n51860 , n51857 , n51859 );
nand ( n51861 , n51860 , n19938 );
not ( n51862 , n19814 );
and ( n51863 , n51861 , n51862 );
or ( n51864 , n38996 , n44582 , RI15b4b810_441);
buf ( n51865 , n19974 );
or ( n51866 , n22362 , n51865 , RI15b49a10_377);
nand ( n51867 , n51864 , n51866 );
nor ( n51868 , n51863 , n51867 );
not ( n51869 , n51862 );
not ( n51870 , n51858 );
nand ( n51871 , n51869 , n383353 , n51870 );
or ( n51872 , n44584 , n20547 );
and ( n51873 , n22378 , n51865 );
nor ( n51874 , n51873 , n22383 );
or ( n51875 , n51874 , n19975 );
nand ( n51876 , n51872 , n51875 );
nand ( n51877 , n51876 , n20501 );
and ( n51878 , n22388 , RI15b4b810_441);
and ( n51879 , n32621 , RI15b4a910_409);
nor ( n51880 , n51878 , n51879 , n383396 );
nand ( n51881 , n51868 , n51871 , n51877 , n51880 );
buf ( n51882 , n51881 );
buf ( n51883 , n380942 );
buf ( n51884 , n22788 );
buf ( n51885 , n380865 );
not ( n51886 , RI15b541e0_735);
nor ( n51887 , n51886 , n383169 );
buf ( n51888 , n51887 );
not ( n51889 , n33220 );
not ( n51890 , n380703 );
or ( n51891 , n51889 , n51890 );
and ( n51892 , n380719 , n33226 );
or ( n51893 , n33237 , n18295 );
or ( n51894 , n48871 , n33241 );
or ( n51895 , n33235 , n380790 );
nand ( n51896 , n51893 , n51894 , n51895 );
nor ( n51897 , n51892 , n51896 );
nand ( n51898 , n51891 , n51897 );
buf ( n51899 , n51898 );
or ( n51900 , n43420 , n32024 );
not ( n51901 , n32909 );
nand ( n51902 , n51900 , n51901 );
not ( n51903 , n33255 );
not ( n51904 , n32035 );
not ( n51905 , n51904 );
or ( n51906 , n51903 , n51905 );
nand ( n51907 , n51906 , n33254 );
and ( n51908 , n51907 , n32909 );
not ( n51909 , n382495 );
nand ( n51910 , n51909 , n32904 );
not ( n51911 , n32915 );
or ( n51912 , n51910 , n51911 );
or ( n51913 , n382129 , n382130 );
nand ( n51914 , n51913 , n51910 , n382142 );
nand ( n51915 , n51912 , n51914 );
or ( n51916 , n44072 , n51915 );
and ( n51917 , n382523 , RI15b4bd38_452);
and ( n51918 , n42720 , RI15b45b40_243);
nor ( n51919 , n51917 , n51918 );
nand ( n51920 , n51916 , n51919 );
nor ( n51921 , n51908 , n51920 );
nand ( n51922 , n51902 , n51921 );
buf ( n51923 , n51922 );
buf ( n51924 , n20665 );
buf ( n51925 , n19653 );
buf ( n51926 , n22714 );
buf ( n51927 , n22716 );
buf ( n51928 , n32255 );
buf ( n51929 , n382073 );
buf ( n51930 , n32271 );
buf ( n51931 , n382065 );
not ( n51932 , n379825 );
not ( n51933 , n50054 );
or ( n51934 , n51932 , n51933 );
nand ( n51935 , n51934 , n41032 );
nand ( n51936 , n51935 , n50058 );
nor ( n51937 , n41036 , n50058 );
and ( n51938 , n50060 , n51937 );
not ( n51939 , RI15b466f8_268);
not ( n51940 , n41581 );
or ( n51941 , n51939 , n51940 );
nand ( n51942 , n51941 , n49638 );
nor ( n51943 , n51938 , n51942 );
nand ( n51944 , n51936 , n51943 );
buf ( n51945 , n51944 );
buf ( n51946 , n386760 );
buf ( n51947 , n380203 );
not ( n51948 , RI15b52548_674);
not ( n51949 , n381485 );
or ( n51950 , n51948 , n51949 );
or ( n51951 , n381423 , n41854 );
nand ( n51952 , n51951 , n381450 );
and ( n51953 , n51952 , n42245 );
and ( n51954 , n42247 , n381461 );
nor ( n51955 , n51953 , n51954 , n44874 );
nand ( n51956 , n51950 , n51955 );
buf ( n51957 , n51956 );
or ( n51958 , n31793 , n384558 );
and ( n51959 , n31770 , RI15b5c958_1024);
or ( n51960 , n39574 , n38910 );
or ( n51961 , n31779 , n384433 );
nand ( n51962 , n51960 , n51961 );
nor ( n51963 , n51959 , n51962 );
nand ( n51964 , n51958 , n38928 , n51963 );
buf ( n51965 , n51964 );
buf ( n51966 , n31719 );
buf ( n51967 , n380865 );
buf ( n51968 , n22655 );
buf ( n51969 , n31979 );
not ( n51970 , n39941 );
not ( n51971 , n50348 );
not ( n51972 , n51971 );
buf ( n51973 , n50336 );
and ( n51974 , n51973 , RI15b44970_205);
nor ( n51975 , n50308 , n50326 );
nand ( n51976 , n51975 , n43641 );
or ( n51977 , n51973 , n51976 );
not ( n51978 , n51975 );
nand ( n51979 , n51978 , RI15b44970_205);
nand ( n51980 , n51977 , n51979 );
nor ( n51981 , n51974 , n51980 );
not ( n51982 , n51981 );
and ( n51983 , n51972 , n51982 );
and ( n51984 , n51971 , n51981 );
nor ( n51985 , n51983 , n51984 );
and ( n51986 , n51970 , n51985 );
not ( n51987 , n51970 );
nand ( n51988 , n50302 , n50316 );
or ( n51989 , n50305 , n43641 );
or ( n51990 , n385943 , n51976 );
nand ( n51991 , n51989 , n51990 , n51979 );
and ( n51992 , n51988 , n51991 );
not ( n51993 , n51988 );
not ( n51994 , n51991 );
and ( n51995 , n51993 , n51994 );
nor ( n51996 , n51992 , n51995 );
and ( n51997 , n51987 , n51996 );
nor ( n51998 , n51986 , n51997 );
buf ( n51999 , n49069 );
nand ( n52000 , n51998 , n51999 );
not ( n52001 , n50323 );
nand ( n52002 , n52001 , n50329 );
and ( n52003 , n50324 , RI15b44970_205);
or ( n52004 , n51976 , n386243 );
nand ( n52005 , n52004 , n51979 );
nor ( n52006 , n52003 , n52005 );
not ( n52007 , n52006 );
and ( n52008 , n52002 , n52007 );
not ( n52009 , n52002 );
and ( n52010 , n52009 , n52006 );
nor ( n52011 , n52008 , n52010 );
or ( n52012 , n52011 , n48511 );
not ( n52013 , n50351 );
not ( n52014 , RI15b4c008_458);
or ( n52015 , n52013 , n52014 );
nand ( n52016 , n52012 , n52015 );
or ( n52017 , n41308 , n51981 );
and ( n52018 , n52007 , n386556 );
and ( n52019 , n386540 , RI15b44970_205);
and ( n52020 , n386549 , n51991 );
nor ( n52021 , n52018 , n52019 , n52020 );
nand ( n52022 , n52017 , n52021 );
nor ( n52023 , n52016 , n52022 );
nand ( n52024 , n52000 , n52023 );
buf ( n52025 , n52024 );
buf ( n52026 , n386563 );
buf ( n52027 , n32676 );
not ( n52028 , RI15b49380_363);
or ( n52029 , n381056 , n52028 );
or ( n52030 , n20248 , n381062 );
or ( n52031 , RI15b49380_363 , n381077 );
nand ( n52032 , n52029 , n52030 , n52031 );
buf ( n52033 , n52032 );
buf ( n52034 , n384700 );
buf ( n52035 , n35651 );
or ( n52036 , n381015 , n22022 );
nand ( n52037 , n381017 , RI15b53628_710);
nand ( n52038 , n52036 , n52037 );
buf ( n52039 , n52038 );
buf ( n52040 , n386563 );
buf ( n52041 , n17499 );
not ( n52042 , RI15b47580_299);
not ( n52043 , n385213 );
or ( n52044 , n52042 , n52043 );
and ( n52045 , n385221 , n381962 );
and ( n52046 , n20631 , RI15b46e00_283);
nor ( n52047 , n52045 , n52046 );
nand ( n52048 , n52044 , n52047 );
buf ( n52049 , n52048 );
buf ( n52050 , n32255 );
buf ( n52051 , n384203 );
buf ( n52052 , n383613 );
not ( n52053 , n381292 );
not ( n52054 , n52053 );
or ( n52055 , n32430 , n52054 );
nand ( n52056 , n381417 , n381296 );
and ( n52057 , n386637 , RI15b54d20_759);
and ( n52058 , n43930 , n386671 );
not ( n52059 , RI15b54d20_759);
not ( n52060 , n382642 );
or ( n52061 , n52059 , n52060 );
or ( n52062 , n382642 , RI15b54d20_759);
nand ( n52063 , n52061 , n52062 );
and ( n52064 , n32439 , n52063 );
nor ( n52065 , n52057 , n52058 , n52064 );
and ( n52066 , n52056 , n52065 );
nand ( n52067 , n52055 , n52066 );
buf ( n52068 , n52067 );
buf ( n52069 , n32271 );
not ( n52070 , n386590 );
not ( n52071 , n380703 );
or ( n52072 , n52070 , n52071 );
and ( n52073 , n380719 , n386603 );
not ( n52074 , RI15b5a180_939);
or ( n52075 , n386612 , n52074 );
or ( n52076 , n380782 , n386624 );
or ( n52077 , n386610 , n380790 );
nand ( n52078 , n52075 , n52076 , n52077 );
nor ( n52079 , n52073 , n52078 );
nand ( n52080 , n52072 , n52079 );
buf ( n52081 , n52080 );
buf ( n52082 , n21800 );
buf ( n52083 , n32271 );
not ( n52084 , RI15b510a8_630);
not ( n52085 , n18078 );
or ( n52086 , n52084 , n52085 );
or ( n52087 , n40876 , n18078 );
nand ( n52088 , n52086 , n52087 );
buf ( n52089 , n52088 );
buf ( n52090 , n386760 );
not ( n52091 , n39170 );
nand ( n52092 , n52091 , n379785 );
not ( n52093 , n52092 );
not ( n52094 , n36574 );
or ( n52095 , n52093 , n52094 );
buf ( n52096 , n39171 );
buf ( n52097 , n52096 );
nand ( n52098 , n52095 , n52097 );
nor ( n52099 , n52091 , n52096 );
nand ( n52100 , n40809 , n52099 );
buf ( n52101 , n39194 );
not ( n52102 , n52101 );
buf ( n52103 , n39195 );
not ( n52104 , n52103 );
and ( n52105 , n52102 , n52104 );
not ( n52106 , n52102 );
and ( n52107 , n52106 , n52103 );
nor ( n52108 , n52105 , n52107 );
and ( n52109 , n52108 , n34646 );
not ( n52110 , RI15b5ddf8_1068);
not ( n52111 , n34651 );
or ( n52112 , n52110 , n52111 );
or ( n52113 , n36518 , n379591 );
nand ( n52114 , n52112 , n52113 );
nor ( n52115 , n52109 , n52114 );
nand ( n52116 , n52098 , n52100 , n52115 );
buf ( n52117 , n52116 );
buf ( n52118 , n31719 );
not ( n52119 , n48936 );
not ( n52120 , n52119 );
not ( n52121 , n384122 );
or ( n52122 , n52120 , n52121 );
and ( n52123 , n384164 , n48939 );
or ( n52124 , n48948 , n20899 );
or ( n52125 , n42970 , n48953 );
or ( n52126 , n48946 , n384193 );
nand ( n52127 , n52124 , n52125 , n52126 );
nor ( n52128 , n52123 , n52127 );
nand ( n52129 , n52122 , n52128 );
buf ( n52130 , n52129 );
buf ( n52131 , n380940 );
not ( n52132 , RI15b5ff40_1139);
not ( n52133 , n383601 );
or ( n52134 , n52132 , n52133 );
and ( n52135 , n50027 , n50810 );
and ( n52136 , n383607 , RI15b5e938_1092);
nor ( n52137 , n52135 , n52136 );
nand ( n52138 , n52134 , n52137 );
buf ( n52139 , n52138 );
buf ( n52140 , n381872 );
and ( n52141 , n41267 , n45618 );
or ( n52142 , n386541 , n385950 );
or ( n52143 , n385946 , n386550 );
or ( n52144 , n386557 , n386234 );
nand ( n52145 , n52142 , n52143 , n52144 );
nor ( n52146 , n52141 , n52145 );
nand ( n52147 , n45625 , n52146 );
buf ( n52148 , n52147 );
buf ( n52149 , n381004 );
buf ( n52150 , n32672 );
buf ( n52151 , n381872 );
buf ( n52152 , n387159 );
buf ( n52153 , n22404 );
buf ( n52154 , n33250 );
not ( n52155 , RI15b47d78_316);
nor ( n52156 , n52155 , n385212 );
buf ( n52157 , n52156 );
buf ( n52158 , n379844 );
buf ( n52159 , n379895 );
buf ( n52160 , n381006 );
and ( n52161 , n22142 , n36120 );
not ( n52162 , n36306 );
nor ( n52163 , n52161 , n52162 );
or ( n52164 , n52163 , n20638 );
or ( n52165 , n22216 , n35932 );
and ( n52166 , n38248 , RI15b3fdf8_44);
and ( n52167 , n381925 , n22109 );
nor ( n52168 , n52166 , n52167 );
nand ( n52169 , n52164 , n52165 , n52168 );
buf ( n52170 , n52169 );
not ( n52171 , n36082 );
not ( n52172 , n52171 );
not ( n52173 , n32129 );
or ( n52174 , n52172 , n52173 );
and ( n52175 , n38230 , RI15b41220_87);
or ( n52176 , n32141 , n36086 );
or ( n52177 , n32148 , n36098 );
or ( n52178 , n36092 , n32150 );
nand ( n52179 , n52176 , n52177 , n52178 );
nor ( n52180 , n52175 , n52179 );
nand ( n52181 , n52174 , n52180 );
buf ( n52182 , n52181 );
buf ( n52183 , n379802 );
buf ( n52184 , n383498 );
buf ( n52185 , n30992 );
buf ( n52186 , n383613 );
buf ( n52187 , RI15b45e88_250);
not ( n52188 , n52171 );
not ( n52189 , n35838 );
or ( n52190 , n52188 , n52189 );
and ( n52191 , n33196 , n36084 );
not ( n52192 , RI15b414f0_93);
or ( n52193 , n36094 , n52192 );
or ( n52194 , n22241 , n36098 );
or ( n52195 , n36092 , n33201 );
nand ( n52196 , n52193 , n52194 , n52195 );
nor ( n52197 , n52191 , n52196 );
nand ( n52198 , n52190 , n52197 );
buf ( n52199 , n52198 );
buf ( n52200 , n381006 );
buf ( n52201 , n380203 );
buf ( n52202 , n31979 );
not ( n52203 , n43203 );
not ( n52204 , n384122 );
or ( n52205 , n52203 , n52204 );
and ( n52206 , n384164 , n385006 );
or ( n52207 , n385019 , n20895 );
or ( n52208 , n33131 , n385023 );
or ( n52209 , n385017 , n384193 );
nand ( n52210 , n52207 , n52208 , n52209 );
nor ( n52211 , n52206 , n52210 );
nand ( n52212 , n52205 , n52211 );
buf ( n52213 , n52212 );
buf ( n52214 , n31030 );
buf ( n52215 , n22009 );
not ( n52216 , n43187 );
not ( n52217 , n379787 );
or ( n52218 , n52216 , n52217 );
or ( n52219 , n43193 , RI15b63a50_1265);
nand ( n52220 , n52218 , n52219 );
buf ( n52221 , n52220 );
buf ( n52222 , n20663 );
buf ( n52223 , n32271 );
or ( n52224 , n382679 , n383021 );
and ( n52225 , n48775 , n386667 );
or ( n52226 , n382691 , n383645 );
not ( n52227 , n382658 );
and ( n52228 , n52227 , RI15b55248_770);
not ( n52229 , n52227 );
and ( n52230 , n52229 , n383021 );
nor ( n52231 , n52228 , n52230 );
or ( n52232 , n52231 , n382625 );
nand ( n52233 , n52226 , n52232 );
nor ( n52234 , n52225 , n52233 , n32410 );
nand ( n52235 , n52224 , n52234 );
buf ( n52236 , n52235 );
not ( n52237 , n35784 );
not ( n52238 , n33400 );
or ( n52239 , n52237 , n52238 );
and ( n52240 , n33415 , n35790 );
or ( n52241 , n35803 , n18475 );
or ( n52242 , n36293 , n35811 );
or ( n52243 , n35801 , n33443 );
nand ( n52244 , n52241 , n52242 , n52243 );
nor ( n52245 , n52240 , n52244 );
nand ( n52246 , n52239 , n52245 );
buf ( n52247 , n52246 );
buf ( n52248 , n380940 );
buf ( n52249 , n22009 );
buf ( n52250 , n22007 );
buf ( n52251 , n381707 );
and ( n52252 , n22515 , n21771 );
not ( n52253 , n37997 );
or ( n52254 , n52253 , RI15b570c0_835);
nand ( n52255 , n52254 , n21790 );
and ( n52256 , n52255 , RI15b57138_836);
nor ( n52257 , n21758 , RI15b57138_836);
and ( n52258 , n21795 , n52257 );
nor ( n52259 , n52252 , n52256 , n52258 );
nand ( n52260 , n33649 , n52259 );
buf ( n52261 , n52260 );
not ( n52262 , n21901 );
nor ( n52263 , n52262 , n21909 );
and ( n52264 , n21802 , n52263 );
and ( n52265 , n21947 , RI15b57d68_862);
not ( n52266 , n21949 );
buf ( n52267 , n21971 );
not ( n52268 , n52267 );
or ( n52269 , n52266 , n52268 );
nand ( n52270 , n52269 , n21979 );
and ( n52271 , n52270 , RI15b55f68_798);
nor ( n52272 , n52265 , n52271 );
or ( n52273 , n52272 , n18078 );
and ( n52274 , n18188 , n21944 , n21986 );
or ( n52275 , n22601 , n52267 , RI15b55f68_798);
and ( n52276 , n18177 , RI15b57d68_862);
and ( n52277 , n18219 , RI15b56e68_830);
nor ( n52278 , n52276 , n52277 , n21751 );
nand ( n52279 , n52275 , n52278 );
nor ( n52280 , n52274 , n52279 );
nand ( n52281 , n52273 , n52280 );
nor ( n52282 , n52264 , n52281 );
not ( n52283 , n17507 );
not ( n52284 , n52262 );
or ( n52285 , n52283 , n52284 );
nand ( n52286 , n52285 , n17565 );
nand ( n52287 , n52286 , n21909 );
nand ( n52288 , n52282 , n52287 );
buf ( n52289 , n52288 );
buf ( n52290 , n381490 );
buf ( n52291 , n381566 );
buf ( n52292 , n385195 );
not ( n52293 , n379363 );
not ( n52294 , n34715 );
or ( n52295 , n52293 , n52294 );
nand ( n52296 , n52295 , n34717 );
buf ( n52297 , n52296 );
not ( n52298 , n32680 );
not ( n52299 , n380703 );
or ( n52300 , n52298 , n52299 );
and ( n52301 , n380719 , n35222 );
or ( n52302 , n32692 , n19017 );
or ( n52303 , n37542 , n32699 );
or ( n52304 , n32690 , n380790 );
nand ( n52305 , n52302 , n52303 , n52304 );
nor ( n52306 , n52301 , n52305 );
nand ( n52307 , n52300 , n52306 );
buf ( n52308 , n52307 );
buf ( n52309 , n384218 );
buf ( n52310 , n22404 );
buf ( n52311 , n384203 );
not ( n52312 , RI15b533d0_705);
not ( n52313 , n383170 );
or ( n52314 , n52312 , n52313 );
and ( n52315 , n33453 , RI15b54960_751);
and ( n52316 , n383147 , RI15b52c50_689);
nor ( n52317 , n52315 , n52316 );
nand ( n52318 , n52314 , n52317 );
buf ( n52319 , n52318 );
not ( n52320 , n35983 );
not ( n52321 , n381589 );
or ( n52322 , n52320 , n52321 );
and ( n52323 , n381596 , n35987 );
or ( n52324 , n35996 , n18712 );
not ( n52325 , n382997 );
or ( n52326 , n52325 , n36003 );
or ( n52327 , n35994 , n381621 );
nand ( n52328 , n52324 , n52326 , n52327 );
nor ( n52329 , n52323 , n52328 );
nand ( n52330 , n52322 , n52329 );
buf ( n52331 , n52330 );
buf ( n52332 , n32676 );
buf ( n52333 , n382052 );
buf ( n52334 , n22479 );
or ( n52335 , n381056 , n32816 );
and ( n52336 , n386555 , RI15b40230_53);
and ( n52337 , n32815 , n32816 );
not ( n52338 , n32815 );
and ( n52339 , n52338 , RI15b496c8_370);
nor ( n52340 , n52337 , n52339 );
and ( n52341 , n36064 , n52340 );
nor ( n52342 , n52336 , n52341 );
nand ( n52343 , n52335 , n52342 );
buf ( n52344 , n52343 );
buf ( n52345 , n32676 );
buf ( n52346 , n381021 );
not ( n52347 , RI15b541e0_735);
not ( n52348 , n32244 );
or ( n52349 , n52347 , n52348 );
and ( n52350 , n32247 , RI15b657d8_1328);
and ( n52351 , n32249 , RI15b60648_1154);
nor ( n52352 , n52350 , n52351 );
nand ( n52353 , n52349 , n52352 );
buf ( n52354 , n52353 );
or ( n52355 , n382512 , n382284 );
and ( n52356 , n382523 , RI15b4b270_429);
and ( n52357 , n382528 , RI15b45078_220);
not ( n52358 , n382160 );
and ( n52359 , n382080 , n52358 );
nor ( n52360 , n52356 , n52357 , n52359 );
nand ( n52361 , n52355 , n52360 );
buf ( n52362 , n52361 );
buf ( n52363 , n19655 );
buf ( n52364 , n383613 );
buf ( n52365 , n33250 );
buf ( n52366 , n32160 );
buf ( n52367 , RI15b5e0c8_1074);
buf ( n52368 , n32160 );
not ( n52369 , n20637 );
not ( n52370 , n19691 );
or ( n52371 , n52369 , n52370 );
nand ( n52372 , n52371 , n34798 );
and ( n52373 , n52372 , RI15b4ad48_418);
or ( n52374 , n34801 , n19691 , RI15b4ad48_418);
not ( n52375 , n19875 );
or ( n52376 , n52375 , n22216 );
nand ( n52377 , n52374 , n52376 );
nor ( n52378 , n52373 , n52377 );
nand ( n52379 , n49028 , n52378 );
buf ( n52380 , n52379 );
buf ( n52381 , n384700 );
buf ( n52382 , n22404 );
buf ( n52383 , n33250 );
and ( n52384 , n34812 , RI15b64158_1280);
buf ( n52385 , n386976 );
not ( n52386 , n52385 );
not ( n52387 , n38093 );
or ( n52388 , n52386 , n52387 );
nand ( n52389 , n52388 , n34823 );
and ( n52390 , n52389 , RI15b62358_1216);
or ( n52391 , n34826 , n52385 , RI15b62358_1216);
not ( n52392 , n387034 );
not ( n52393 , n52392 );
not ( n52394 , RI15b64158_1280);
and ( n52395 , n52393 , n52394 );
and ( n52396 , n52392 , RI15b64158_1280);
nor ( n52397 , n52395 , n52396 );
or ( n52398 , n34833 , n52397 );
nand ( n52399 , n52391 , n52398 );
nor ( n52400 , n52384 , n52390 , n52399 );
or ( n52401 , n52400 , n19200 );
buf ( n52402 , n386853 );
not ( n52403 , n52402 );
not ( n52404 , n22473 );
and ( n52405 , n52403 , n52404 );
nor ( n52406 , n52405 , n386943 );
or ( n52407 , n48387 , n52406 );
and ( n52408 , n38117 , n52402 , n48387 );
or ( n52409 , n22424 , n379431 );
or ( n52410 , n386854 , n19598 );
nand ( n52411 , n52409 , n52410 , n19512 );
nor ( n52412 , n52408 , n52411 );
nand ( n52413 , n52401 , n52407 , n52412 );
buf ( n52414 , n52413 );
buf ( n52415 , n33382 );
buf ( n52416 , n22009 );
not ( n52417 , n385791 );
not ( n52418 , n52417 );
buf ( n52419 , n39952 );
not ( n52420 , n52419 );
or ( n52421 , n52418 , n52420 );
or ( n52422 , n52419 , n52417 );
nand ( n52423 , n52421 , n52422 );
and ( n52424 , n52423 , n386020 );
not ( n52425 , n386172 );
not ( n52426 , n52425 );
not ( n52427 , n39966 );
or ( n52428 , n52426 , n52427 );
or ( n52429 , n39966 , n52425 );
nand ( n52430 , n52428 , n52429 );
nand ( n52431 , n52430 , n39974 );
not ( n52432 , n34733 );
not ( n52433 , n41297 );
or ( n52434 , n52432 , n52433 );
not ( n52435 , n39980 );
nand ( n52436 , n52434 , n52435 );
and ( n52437 , n52436 , n386500 );
and ( n52438 , n39988 , RI15b4b798_440);
nor ( n52439 , n52437 , n52438 );
nand ( n52440 , n52431 , n52439 );
nor ( n52441 , n52424 , n52440 );
and ( n52442 , n49029 , n34733 );
or ( n52443 , n386541 , n385783 );
or ( n52444 , n52417 , n386550 );
or ( n52445 , n52425 , n386557 );
nand ( n52446 , n52443 , n52444 , n52445 );
nor ( n52447 , n52442 , n52446 );
nand ( n52448 , n52441 , n52447 );
buf ( n52449 , n52448 );
buf ( n52450 , n18226 );
buf ( n52451 , n380906 );
buf ( n52452 , n380903 );
not ( n52453 , n31442 );
buf ( n52454 , n31446 );
nand ( n52455 , n52453 , n52454 );
not ( n52456 , n52455 );
not ( n52457 , n49807 );
nor ( n52458 , n52457 , n49805 );
not ( n52459 , n52458 );
and ( n52460 , n52456 , n52459 );
and ( n52461 , n52455 , n52458 );
nor ( n52462 , n52460 , n52461 );
not ( n52463 , n45735 );
or ( n52464 , n52462 , n52463 );
not ( n52465 , n379391 );
nor ( n52466 , n49816 , n379248 );
not ( n52467 , n52466 );
or ( n52468 , n52465 , n52467 );
nand ( n52469 , n52468 , n31700 );
and ( n52470 , n52469 , n31404 );
or ( n52471 , n52466 , n40972 , n31404 );
and ( n52472 , n379394 , RI15b580b0_869);
and ( n52473 , n31712 , RI15b51eb8_660);
nor ( n52474 , n52472 , n52473 );
nand ( n52475 , n52471 , n52474 );
nor ( n52476 , n52470 , n52475 );
nand ( n52477 , n52464 , n52476 );
buf ( n52478 , n52477 );
and ( n52479 , n31792 , n31933 );
or ( n52480 , n31771 , n31835 );
or ( n52481 , n31891 , n37611 );
not ( n52482 , n31841 );
or ( n52483 , n31779 , n52482 );
nand ( n52484 , n52480 , n52481 , n52483 );
nor ( n52485 , n52479 , n52484 );
nand ( n52486 , n45174 , n52485 );
buf ( n52487 , n52486 );
buf ( n52488 , n381081 );
buf ( n52489 , n382537 );
buf ( n52490 , n381004 );
not ( n52491 , n34737 );
not ( n52492 , n39977 );
or ( n52493 , n52491 , n52492 );
not ( n52494 , n34738 );
nand ( n52495 , n52493 , n52494 );
and ( n52496 , n52495 , n386500 );
not ( n52497 , n386174 );
and ( n52498 , n52497 , n386210 );
not ( n52499 , n52497 );
not ( n52500 , n386210 );
and ( n52501 , n52499 , n52500 );
nor ( n52502 , n52498 , n52501 );
not ( n52503 , n386262 );
or ( n52504 , n52502 , n52503 );
not ( n52505 , n385834 );
not ( n52506 , n52505 );
not ( n52507 , n385826 );
or ( n52508 , n52506 , n52507 );
or ( n52509 , n385826 , n52505 );
nand ( n52510 , n52508 , n52509 );
and ( n52511 , n52510 , n30873 );
not ( n52512 , n22396 );
not ( n52513 , n52512 );
and ( n52514 , n52513 , RI15b4b888_442);
nor ( n52515 , n52511 , n52514 );
nand ( n52516 , n52504 , n52515 );
nor ( n52517 , n52496 , n52516 );
and ( n52518 , n41267 , n34737 );
or ( n52519 , n386541 , n385828 );
or ( n52520 , n385834 , n386550 );
or ( n52521 , n52500 , n386557 );
nand ( n52522 , n52519 , n52520 , n52521 );
nor ( n52523 , n52518 , n52522 );
nand ( n52524 , n52517 , n52523 );
buf ( n52525 , n52524 );
buf ( n52526 , n35649 );
buf ( n52527 , n32160 );
buf ( n52528 , n382073 );
or ( n52529 , n36238 , n31163 );
or ( n52530 , n17957 , n31175 );
not ( n52531 , n31182 );
and ( n52532 , n52531 , n32711 );
and ( n52533 , n383803 , n39380 );
and ( n52534 , n36261 , n31180 );
nor ( n52535 , n52532 , n52533 , n52534 );
nand ( n52536 , n52529 , n52530 , n52535 );
buf ( n52537 , n52536 );
buf ( n52538 , n379802 );
or ( n52539 , n31091 , n32281 );
and ( n52540 , n38654 , RI15b5b0f8_972);
and ( n52541 , n39717 , RI15b5ad38_964);
nor ( n52542 , n52540 , n52541 );
and ( n52543 , n39721 , RI15b5a978_956);
and ( n52544 , n39724 , RI15b5a5b8_948);
nor ( n52545 , n52543 , n52544 );
and ( n52546 , n39728 , RI15b5a1f8_940);
and ( n52547 , n39731 , RI15b59e38_932);
nor ( n52548 , n52546 , n52547 );
and ( n52549 , n39735 , RI15b59a78_924);
and ( n52550 , n39738 , RI15b596b8_916);
nor ( n52551 , n52549 , n52550 );
nand ( n52552 , n52542 , n52545 , n52548 , n52551 );
and ( n52553 , n41935 , n52552 );
and ( n52554 , n39746 , RI15b58b78_892);
and ( n52555 , n39751 , RI15b5bff8_1004);
nor ( n52556 , n52553 , n52554 , n52555 );
and ( n52557 , n39756 , RI15b5bc38_996);
and ( n52558 , n39759 , RI15b5b878_988);
nor ( n52559 , n52557 , n52558 );
and ( n52560 , n39763 , RI15b592f8_908);
and ( n52561 , n39765 , RI15b58f38_900);
nor ( n52562 , n52560 , n52561 );
and ( n52563 , n39769 , RI15b587b8_884);
and ( n52564 , n39772 , RI15b5b4b8_980);
nor ( n52565 , n52563 , n52564 );
nand ( n52566 , n52556 , n52559 , n52562 , n52565 );
and ( n52567 , n52566 , n47195 );
not ( n52568 , n380416 );
or ( n52569 , n31052 , n52568 );
not ( n52570 , n41414 );
not ( n52571 , n32281 );
and ( n52572 , n52570 , n52571 );
and ( n52573 , n41414 , n32281 );
nor ( n52574 , n52572 , n52573 );
or ( n52575 , n52574 , n43838 );
nand ( n52576 , n52569 , n52575 , n51123 );
nor ( n52577 , n52567 , n52576 );
nand ( n52578 , n52539 , n52577 );
buf ( n52579 , n52578 );
buf ( n52580 , n35651 );
buf ( n52581 , n381021 );
and ( n52582 , n22646 , RI15b45348_226);
and ( n52583 , n22648 , RI15b517b0_645);
nor ( n52584 , n52582 , n52583 );
not ( n52585 , n52584 );
buf ( n52586 , n52585 );
buf ( n52587 , n384700 );
or ( n52588 , n20640 , n382158 );
and ( n52589 , n22368 , RI15b4a280_395);
nor ( n52590 , n52589 , n20656 );
or ( n52591 , n52590 , n19676 );
or ( n52592 , n19937 , n37053 );
nand ( n52593 , n52592 , n19676 );
and ( n52594 , n20521 , RI15b493f8_364);
not ( n52595 , RI15b493f8_364);
and ( n52596 , n52595 , RI15b49380_363);
and ( n52597 , n52028 , RI15b493f8_364);
nor ( n52598 , n52596 , n52597 );
or ( n52599 , n20529 , n52598 );
or ( n52600 , RI15b4b1f8_428 , n22353 );
or ( n52601 , n36723 , n37048 );
nand ( n52602 , n52599 , n52600 , n52601 );
nor ( n52603 , n52594 , n52602 );
and ( n52604 , n52593 , n52603 );
nand ( n52605 , n52588 , n52591 , n52604 );
buf ( n52606 , n52605 );
buf ( n52607 , n22716 );
buf ( n52608 , n385195 );
and ( n52609 , n37076 , RI15b63ca8_1270);
buf ( n52610 , n386960 );
not ( n52611 , n52610 );
not ( n52612 , n38093 );
or ( n52613 , n52611 , n52612 );
nand ( n52614 , n52613 , n34823 );
and ( n52615 , n52614 , RI15b61ea8_1206);
or ( n52616 , n34826 , n52610 , RI15b61ea8_1206);
not ( n52617 , RI15b63ca8_1270);
and ( n52618 , n37071 , n52617 , RI15b63c30_1269);
nor ( n52619 , n52618 , n379545 );
or ( n52620 , n34833 , n52619 );
nand ( n52621 , n52616 , n52620 );
nor ( n52622 , n52609 , n52615 , n52621 );
or ( n52623 , n52622 , n19200 );
not ( n52624 , n386804 );
not ( n52625 , n52624 );
not ( n52626 , n22473 );
and ( n52627 , n52625 , n52626 );
nor ( n52628 , n52627 , n44568 );
or ( n52629 , n386811 , n52628 );
and ( n52630 , n387011 , n52624 , n386811 );
not ( n52631 , RI15b63ca8_1270);
or ( n52632 , n22424 , n52631 );
or ( n52633 , n386809 , n19598 );
nand ( n52634 , n52632 , n52633 , n19512 );
nor ( n52635 , n52630 , n52634 );
nand ( n52636 , n52623 , n52629 , n52635 );
buf ( n52637 , n52636 );
buf ( n52638 , n22343 );
or ( n52639 , n22315 , n35895 );
and ( n52640 , n22326 , n39462 );
or ( n52641 , n35911 , n46122 );
or ( n52642 , n22334 , n35917 );
or ( n52643 , n35909 , n22336 );
nand ( n52644 , n52641 , n52642 , n52643 );
nor ( n52645 , n52640 , n52644 );
nand ( n52646 , n52639 , n52645 );
buf ( n52647 , n52646 );
or ( n52648 , n22102 , n35869 );
and ( n52649 , n22203 , n35872 );
or ( n52650 , n35884 , n385499 );
or ( n52651 , n22293 , n35888 );
or ( n52652 , n35882 , n22299 );
nand ( n52653 , n52650 , n52651 , n52652 );
nor ( n52654 , n52649 , n52653 );
nand ( n52655 , n52648 , n52654 );
buf ( n52656 , n52655 );
buf ( n52657 , n379403 );
buf ( n52658 , n383498 );
buf ( n52659 , n30992 );
buf ( n52660 , n35649 );
or ( n52661 , n381407 , n32432 );
not ( n52662 , n40054 );
not ( n52663 , n38897 );
or ( n52664 , n52662 , n52663 );
nand ( n52665 , n52664 , n381450 );
and ( n52666 , n52665 , n40052 );
and ( n52667 , n381461 , n43714 );
nor ( n52668 , n52666 , n52667 );
and ( n52669 , n32435 , n52668 );
nand ( n52670 , n381486 , RI15b53100_699);
nand ( n52671 , n52661 , n52669 , n52670 );
buf ( n52672 , n52671 );
not ( n52673 , n381494 );
not ( n52674 , n382912 );
or ( n52675 , n52673 , n52674 );
and ( n52676 , n382931 , n381528 );
not ( n52677 , RI15b5bda0_999);
or ( n52678 , n381544 , n52677 );
or ( n52679 , n35163 , n381557 );
or ( n52680 , n381542 , n382967 );
nand ( n52681 , n52678 , n52679 , n52680 );
nor ( n52682 , n52676 , n52681 );
nand ( n52683 , n52675 , n52682 );
buf ( n52684 , n52683 );
buf ( n52685 , n22404 );
not ( n52686 , n51226 );
not ( n52687 , n384122 );
or ( n52688 , n52686 , n52687 );
and ( n52689 , n384164 , n33600 );
or ( n52690 , n33609 , n20885 );
or ( n52691 , n33131 , n33615 );
or ( n52692 , n33607 , n384193 );
nand ( n52693 , n52690 , n52691 , n52692 );
nor ( n52694 , n52689 , n52693 );
nand ( n52695 , n52688 , n52694 );
buf ( n52696 , n52695 );
buf ( n52697 , n22714 );
buf ( n52698 , n379403 );
nand ( n52699 , n41674 , n40781 );
not ( n52700 , n33580 );
not ( n52701 , n33568 );
or ( n52702 , n52700 , n52701 );
nand ( n52703 , n52702 , n33584 );
nand ( n52704 , n52703 , n41673 );
nand ( n52705 , n383601 , RI15b60300_1147);
nand ( n52706 , n383607 , RI15b5ecf8_1100);
nand ( n52707 , n52699 , n52704 , n52705 , n52706 );
buf ( n52708 , n52707 );
buf ( n52709 , n31979 );
and ( n52710 , n379822 , n41043 );
nor ( n52711 , n379834 , n382000 );
nor ( n52712 , n52710 , n52711 );
nand ( n52713 , n379832 , RI15b46b30_277);
nand ( n52714 , n379825 , RI15b48840_339);
nand ( n52715 , n52712 , n52713 , n52714 );
buf ( n52716 , n52715 );
buf ( n52717 , n19651 );
buf ( n52718 , n380865 );
buf ( n52719 , n382537 );
buf ( n52720 , n383498 );
buf ( n52721 , RI15b5de70_1069);
buf ( n52722 , n35649 );
or ( n52723 , n40340 , n22598 );
not ( n52724 , n382884 );
buf ( n52725 , n48195 );
not ( n52726 , n52725 );
and ( n52727 , n52724 , n52726 );
and ( n52728 , n40348 , n22598 );
nor ( n52729 , n52727 , n52728 );
nand ( n52730 , n52723 , n52729 );
buf ( n52731 , n52730 );
not ( n52732 , n380235 );
not ( n52733 , n382912 );
or ( n52734 , n52732 , n52733 );
and ( n52735 , n382931 , n380745 );
or ( n52736 , n380776 , n19084 );
or ( n52737 , n35805 , n380785 );
or ( n52738 , n380768 , n382967 );
nand ( n52739 , n52736 , n52737 , n52738 );
nor ( n52740 , n52735 , n52739 );
nand ( n52741 , n52734 , n52740 );
buf ( n52742 , n52741 );
buf ( n52743 , n22738 );
buf ( n52744 , n379802 );
or ( n52745 , n385163 , n21091 );
and ( n52746 , n385173 , n21398 );
and ( n52747 , n385177 , n21397 );
nor ( n52748 , n52746 , n52747 );
and ( n52749 , n32368 , n21097 );
nor ( n52750 , n52749 , n35720 );
nand ( n52751 , n52745 , n52748 , n52750 );
buf ( n52752 , n52751 );
buf ( n52753 , n32271 );
buf ( n52754 , n382069 );
and ( n52755 , n33576 , n37775 );
nor ( n52756 , n52755 , n37781 );
or ( n52757 , n33541 , n52756 );
nor ( n52758 , n33576 , n384933 );
nand ( n52759 , n33541 , n52758 );
and ( n52760 , n384918 , RI15b5ee60_1103);
nor ( n52761 , n52760 , n46090 );
nand ( n52762 , n52757 , n52759 , n52761 );
buf ( n52763 , n52762 );
or ( n52764 , n35333 , n38460 );
and ( n52765 , n386554 , n39301 );
and ( n52766 , n35363 , n38460 );
nor ( n52767 , n385202 , n379828 , n35582 );
nor ( n52768 , n52765 , n52766 , n52767 );
nand ( n52769 , n52764 , n52768 );
buf ( n52770 , n52769 );
buf ( n52771 , n31033 );
buf ( n52772 , n21800 );
buf ( n52773 , n380865 );
buf ( n52774 , n381707 );
buf ( n52775 , RI15b5e320_1079);
buf ( n52776 , n381004 );
buf ( n52777 , n383345 );
or ( n52778 , n22102 , n36306 );
and ( n52779 , n22203 , n36309 );
or ( n52780 , n36318 , n385511 );
or ( n52781 , n22293 , n36325 );
or ( n52782 , n36316 , n22299 );
nand ( n52783 , n52780 , n52781 , n52782 );
nor ( n52784 , n52779 , n52783 );
nand ( n52785 , n52778 , n52784 );
buf ( n52786 , n52785 );
buf ( n52787 , n22788 );
buf ( n52788 , n31979 );
buf ( n52789 , n379403 );
buf ( n52790 , n43349 );
or ( n52791 , n381907 , n37663 );
and ( n52792 , n43131 , RI15b42918_136);
or ( n52793 , n381917 , n37665 );
not ( n52794 , n37679 );
and ( n52795 , n52794 , n381923 );
and ( n52796 , n381926 , n37677 );
nor ( n52797 , n52795 , n52796 );
nand ( n52798 , n52793 , n52797 );
nor ( n52799 , n52792 , n52798 );
nand ( n52800 , n52791 , n52799 );
buf ( n52801 , n52800 );
buf ( n52802 , n380903 );
buf ( n52803 , n32981 );
buf ( n52804 , n22005 );
not ( n52805 , n31251 );
not ( n52806 , n379343 );
or ( n52807 , n52805 , n52806 );
not ( n52808 , n47629 );
not ( n52809 , n379383 );
nor ( n52810 , n52809 , n379367 );
not ( n52811 , n52810 );
or ( n52812 , n52808 , n52811 );
or ( n52813 , n52810 , n47629 );
nand ( n52814 , n52812 , n52813 );
and ( n52815 , n52814 , n379391 );
and ( n52816 , n379394 , RI15b577c8_850);
and ( n52817 , n379398 , RI15b515d0_641);
nor ( n52818 , n52815 , n52816 , n52817 );
nand ( n52819 , n52807 , n52818 );
buf ( n52820 , n52819 );
buf ( n52821 , n379847 );
and ( n52822 , n34885 , RI15b60a80_1163);
and ( n52823 , n47614 , RI15b5d8d0_1057);
nor ( n52824 , n52822 , n52823 );
not ( n52825 , n52824 );
buf ( n52826 , n52825 );
buf ( n52827 , n48972 );
and ( n52828 , n52827 , n44504 );
nor ( n52829 , n52828 , n35187 );
or ( n52830 , n52829 , n34969 );
nand ( n52831 , n34969 , RI15b48f48_354);
or ( n52832 , n52827 , n52831 );
or ( n52833 , n34969 , RI15b48f48_354);
nand ( n52834 , n52832 , n52833 );
and ( n52835 , n52834 , n48989 );
and ( n52836 , n44858 , n44495 );
and ( n52837 , n35335 , RI15b66390_1353);
nor ( n52838 , n52835 , n52836 , n52837 );
nand ( n52839 , n52830 , n52838 , n41046 );
buf ( n52840 , n52839 );
buf ( n52841 , n381490 );
buf ( n52842 , n31033 );
buf ( n52843 , n381081 );
buf ( n52844 , n32160 );
and ( n52845 , n381014 , RI15b539e8_718);
and ( n52846 , n35213 , RI15b65ee0_1343);
nor ( n52847 , n52845 , n52846 );
not ( n52848 , n52847 );
buf ( n52849 , n52848 );
buf ( n52850 , n386760 );
buf ( n52851 , n383613 );
or ( n52852 , n35852 , n38065 );
and ( n52853 , n43338 , RI15b42be8_142);
or ( n52854 , n35856 , n38075 );
or ( n52855 , n35582 , n38081 );
or ( n52856 , n38069 , n35858 );
nand ( n52857 , n52854 , n52855 , n52856 );
nor ( n52858 , n52853 , n52857 );
nand ( n52859 , n52852 , n52858 );
buf ( n52860 , n52859 );
buf ( n52861 , n22788 );
buf ( n52862 , n382067 );
buf ( n52863 , n22714 );
or ( n52864 , n36937 , n383845 );
and ( n52865 , n36946 , n383878 );
not ( n52866 , RI15b4f2a8_566);
or ( n52867 , n383903 , n52866 );
or ( n52868 , n39875 , n383911 );
or ( n52869 , n383895 , n36955 );
nand ( n52870 , n52867 , n52868 , n52869 );
nor ( n52871 , n52865 , n52870 );
nand ( n52872 , n52864 , n52871 );
buf ( n52873 , n52872 );
buf ( n52874 , n383613 );
and ( n52875 , n383505 , n383539 );
nor ( n52876 , n52875 , n383577 );
or ( n52877 , n52876 , n383546 );
and ( n52878 , n383601 , RI15b5fbf8_1132);
not ( n52879 , n383546 );
nor ( n52880 , n52879 , n383539 );
and ( n52881 , n383603 , n52880 );
and ( n52882 , n383607 , RI15b5f478_1116);
nor ( n52883 , n52878 , n52881 , n52882 );
nand ( n52884 , n52877 , n52883 );
buf ( n52885 , n52884 );
buf ( n52886 , n31979 );
buf ( n52887 , n386563 );
buf ( n52888 , n384700 );
not ( n52889 , n51031 );
or ( n52890 , n52889 , n36051 );
and ( n52891 , n381055 , RI15b49a10_377);
not ( n52892 , RI15b49a10_377);
not ( n52893 , n36057 );
not ( n52894 , n52893 );
or ( n52895 , n52892 , n52894 );
or ( n52896 , n52893 , RI15b49a10_377);
nand ( n52897 , n52895 , n52896 );
and ( n52898 , n381076 , n52897 );
nor ( n52899 , n52891 , n52898 );
nand ( n52900 , n52890 , n52899 );
buf ( n52901 , n52900 );
buf ( n52902 , n382049 );
buf ( n52903 , n382052 );
not ( n52904 , RI15b53e98_728);
not ( n52905 , n32244 );
or ( n52906 , n52904 , n52905 );
and ( n52907 , n32247 , RI15b65490_1321);
and ( n52908 , n32249 , RI15b60300_1147);
nor ( n52909 , n52907 , n52908 );
nand ( n52910 , n52906 , n52909 );
buf ( n52911 , n52910 );
buf ( n52912 , n383498 );
not ( n52913 , RI15b55b30_789);
not ( n52914 , n380000 );
or ( n52915 , n52913 , n52914 );
and ( n52916 , n380010 , RI15b4c698_472);
not ( n52917 , RI15b55b30_789);
not ( n52918 , n379957 );
not ( n52919 , n52918 );
or ( n52920 , n52917 , n52919 );
or ( n52921 , n52918 , RI15b55b30_789);
nand ( n52922 , n52920 , n52921 );
and ( n52923 , n379949 , n52922 );
nor ( n52924 , n52916 , n52923 );
nand ( n52925 , n52915 , n52924 );
buf ( n52926 , n52925 );
or ( n52927 , n386588 , n36394 );
and ( n52928 , n386600 , n36401 );
or ( n52929 , n36410 , n19150 );
or ( n52930 , n386618 , n36416 );
or ( n52931 , n36408 , n386627 );
nand ( n52932 , n52929 , n52930 , n52931 );
nor ( n52933 , n52928 , n52932 );
nand ( n52934 , n52927 , n52933 );
buf ( n52935 , n52934 );
buf ( n52936 , n383613 );
buf ( n52937 , n382537 );
or ( n52938 , n380968 , n36813 );
and ( n52939 , n380986 , n37013 );
not ( n52940 , RI15b42300_123);
xor ( n52941 , n36824 , n52940 );
xor ( n52942 , n380994 , n36830 );
xor ( n52943 , n36822 , n380996 );
nand ( n52944 , n52941 , n52942 , n52943 );
nor ( n52945 , n52939 , n52944 );
nand ( n52946 , n52938 , n52945 );
buf ( n52947 , n52946 );
buf ( n52948 , n379802 );
buf ( n52949 , n381004 );
buf ( n52950 , n35649 );
buf ( n52951 , n19651 );
or ( n52952 , n36238 , n384168 );
not ( n52953 , n384182 );
and ( n52954 , n52953 , RI15b4cad0_481);
or ( n52955 , n384190 , n32710 );
or ( n52956 , n384057 , n383802 );
or ( n52957 , n384180 , n42402 );
nand ( n52958 , n52955 , n52956 , n52957 );
nor ( n52959 , n52954 , n52958 );
nand ( n52960 , n52952 , n52959 );
buf ( n52961 , n52960 );
buf ( n52962 , n22653 );
buf ( n52963 , n22406 );
buf ( n52964 , n385197 );
not ( n52965 , n41933 );
not ( n52966 , n52566 );
or ( n52967 , n52965 , n52966 );
and ( n52968 , n384022 , RI15b623d0_1217);
not ( n52969 , RI15b623d0_1217);
not ( n52970 , n38477 );
not ( n52971 , n52970 );
or ( n52972 , n52969 , n52971 );
or ( n52973 , n52970 , RI15b623d0_1217);
nand ( n52974 , n52972 , n52973 );
and ( n52975 , n52974 , n384025 );
nor ( n52976 , n52968 , n52975 );
nand ( n52977 , n52967 , n52976 );
buf ( n52978 , n52977 );
buf ( n52979 , n35651 );
buf ( n52980 , n380940 );
buf ( n52981 , n382458 );
nor ( n52982 , n52981 , n382079 );
or ( n52983 , n52982 , n382475 );
buf ( n52984 , n382466 );
nand ( n52985 , n52983 , n52984 );
not ( n52986 , n382478 );
and ( n52987 , n382261 , n47592 );
not ( n52988 , n52987 );
or ( n52989 , n52986 , n52988 );
or ( n52990 , n52987 , n382478 );
nand ( n52991 , n52989 , n52990 );
nand ( n52992 , n32962 , n52991 );
not ( n52993 , n32035 );
not ( n52994 , n52984 );
nand ( n52995 , n52993 , n52981 , n52994 );
and ( n52996 , n382523 , RI15b4b4c8_434);
and ( n52997 , n42153 , RI15b452d0_225);
nor ( n52998 , n52996 , n52997 );
nand ( n52999 , n52985 , n52992 , n52995 , n52998 );
buf ( n53000 , n52999 );
buf ( n53001 , n381490 );
buf ( n53002 , n33250 );
buf ( n53003 , n384199 );
or ( n53004 , n40842 , n18078 );
and ( n53005 , n39220 , RI15b50ec8_626);
or ( n53006 , n21407 , RI15b50dd8_624);
or ( n53007 , n21364 , n37927 );
nand ( n53008 , n53006 , n53007 );
and ( n53009 , n32986 , n53008 );
and ( n53010 , n383915 , n385102 );
nor ( n53011 , n53005 , n53009 , n53010 );
nand ( n53012 , n53004 , n53011 );
buf ( n53013 , n53012 );
buf ( n53014 , n381872 );
buf ( n53015 , n17499 );
buf ( n53016 , n43309 );
not ( n53017 , n53016 );
not ( n53018 , n43308 );
not ( n53019 , n53018 );
or ( n53020 , n53017 , n53019 );
or ( n53021 , n53018 , n53016 );
nand ( n53022 , n53020 , n53021 );
nand ( n53023 , n53022 , n34647 );
not ( n53024 , n36564 );
nand ( n53025 , n53024 , n379785 );
not ( n53026 , n53025 );
not ( n53027 , n39798 );
or ( n53028 , n53026 , n53027 );
nand ( n53029 , n53028 , n36565 );
nor ( n53030 , n53024 , n36565 );
and ( n53031 , n51703 , n53030 );
not ( n53032 , RI15b5dfd8_1072);
not ( n53033 , n34651 );
or ( n53034 , n53032 , n53033 );
or ( n53035 , n36518 , n379632 );
nand ( n53036 , n53034 , n53035 );
nor ( n53037 , n53031 , n53036 );
nand ( n53038 , n53023 , n53029 , n53037 );
buf ( n53039 , n53038 );
buf ( n53040 , n379893 );
buf ( n53041 , n383074 );
not ( n53042 , n38897 );
not ( n53043 , n383142 );
or ( n53044 , n53042 , n53043 );
nand ( n53045 , n53044 , n381450 );
and ( n53046 , n53041 , n53045 );
and ( n53047 , n381484 , RI15b52908_682);
nor ( n53048 , n53046 , n53047 );
nor ( n53049 , n383142 , n381460 );
nand ( n53050 , n383075 , n53049 );
nand ( n53051 , n381401 , n52053 );
nand ( n53052 , n53048 , n53050 , n53051 );
buf ( n53053 , n53052 );
or ( n53054 , n31771 , n18229 );
or ( n53055 , n19308 , n31783 );
and ( n53056 , n32386 , n18451 );
nor ( n53057 , n31779 , n19442 );
nor ( n53058 , n53056 , n36902 , n53057 );
nand ( n53059 , n53054 , n53055 , n53058 );
buf ( n53060 , n53059 );
buf ( n53061 , n22716 );
buf ( n53062 , n382052 );
buf ( n53063 , n32676 );
not ( n53064 , n50461 );
or ( n53065 , n53064 , n36051 );
and ( n53066 , n381055 , RI15b498a8_374);
not ( n53067 , RI15b498a8_374);
not ( n53068 , n32822 );
not ( n53069 , n53068 );
or ( n53070 , n53067 , n53069 );
or ( n53071 , n53068 , RI15b498a8_374);
nand ( n53072 , n53070 , n53071 );
and ( n53073 , n381076 , n53072 );
nor ( n53074 , n53066 , n53073 );
nand ( n53075 , n53065 , n53074 );
buf ( n53076 , n53075 );
buf ( n53077 , n384700 );
buf ( n53078 , n20663 );
not ( n53079 , RI15b54000_731);
not ( n53080 , n32244 );
or ( n53081 , n53079 , n53080 );
and ( n53082 , n32247 , RI15b655f8_1324);
and ( n53083 , n32249 , RI15b60468_1150);
nor ( n53084 , n53082 , n53083 );
nand ( n53085 , n53081 , n53084 );
buf ( n53086 , n53085 );
buf ( n53087 , RI15b47b20_311);
buf ( n53088 , n384700 );
and ( n53089 , n30908 , RI15b4a898_408);
and ( n53090 , n19807 , n22217 );
not ( n53091 , RI15b4a898_408);
not ( n53092 , n19671 );
not ( n53093 , n53092 );
or ( n53094 , n53091 , n53093 );
or ( n53095 , n53092 , RI15b4a898_408);
nand ( n53096 , n53094 , n53095 );
and ( n53097 , n53096 , n20637 );
nor ( n53098 , n53089 , n53090 , n53097 );
nand ( n53099 , n52441 , n53098 );
buf ( n53100 , n53099 );
buf ( n53101 , n382067 );
buf ( n53102 , n32255 );
buf ( n53103 , n19653 );
buf ( n53104 , n386914 );
nor ( n53105 , n53104 , n22473 );
or ( n53106 , n53105 , n386946 );
nand ( n53107 , n53106 , n384650 );
buf ( n53108 , n386992 );
not ( n53109 , n53108 );
nor ( n53110 , n53109 , n387006 );
or ( n53111 , n53110 , n383409 );
nand ( n53112 , n53111 , RI15b62808_1226);
or ( n53113 , n53108 , n383482 , RI15b62808_1226);
buf ( n53114 , n30846 );
or ( n53115 , n53114 , n379445 , RI15b64608_1290);
or ( n53116 , n379446 , RI15b64590_1289);
nand ( n53117 , n53115 , n53116 );
and ( n53118 , n53117 , n22450 );
and ( n53119 , n19599 , RI15b63708_1258);
nor ( n53120 , n53118 , n53119 );
nand ( n53121 , n53113 , n53120 );
and ( n53122 , n53114 , n22450 );
nor ( n53123 , n53122 , n22426 );
nor ( n53124 , n53123 , n379446 );
nor ( n53125 , n53121 , n53124 );
nor ( n53126 , n48004 , n384650 );
nand ( n53127 , n53104 , n53126 );
nand ( n53128 , n53107 , n53112 , n53125 , n53127 );
buf ( n53129 , n53128 );
buf ( n53130 , n381872 );
buf ( n53131 , RI15b47148_290);
or ( n53132 , n22587 , n380001 );
not ( n53133 , n380011 );
not ( n53134 , n380166 );
not ( n53135 , n380140 );
not ( n53136 , n53135 );
or ( n53137 , n53134 , n53136 );
or ( n53138 , n53135 , n380166 );
nand ( n53139 , n53137 , n53138 );
not ( n53140 , n53139 );
or ( n53141 , n53133 , n53140 );
and ( n53142 , n379978 , RI15b562b0_805);
not ( n53143 , n379978 );
and ( n53144 , n53143 , n22587 );
nor ( n53145 , n53142 , n53144 );
or ( n53146 , n379948 , n53145 );
nand ( n53147 , n53132 , n53141 , n53146 );
buf ( n53148 , n53147 );
or ( n53149 , n386588 , n47643 );
and ( n53150 , n386600 , n47649 );
or ( n53151 , n47658 , n19162 );
or ( n53152 , n386618 , n47663 );
or ( n53153 , n47656 , n386627 );
nand ( n53154 , n53151 , n53152 , n53153 );
nor ( n53155 , n53150 , n53154 );
nand ( n53156 , n53149 , n53155 );
buf ( n53157 , n53156 );
buf ( n53158 , n383345 );
buf ( n53159 , n19655 );
buf ( n53160 , n385195 );
and ( n53161 , n43978 , n43981 );
not ( n53162 , n43978 );
not ( n53163 , n43981 );
and ( n53164 , n53162 , n53163 );
nor ( n53165 , n53161 , n53164 );
nand ( n53166 , n53165 , n379393 );
not ( n53167 , n31636 );
not ( n53168 , n31631 );
not ( n53169 , n53168 );
or ( n53170 , n53167 , n53169 );
or ( n53171 , n53168 , n31636 );
nand ( n53172 , n53170 , n53171 );
and ( n53173 , n53172 , n379391 );
and ( n53174 , n379394 , RI15b57a20_855);
and ( n53175 , n41206 , RI15b51828_646);
nor ( n53176 , n53173 , n53174 , n53175 );
nand ( n53177 , n53166 , n53176 );
buf ( n53178 , n53177 );
buf ( n53179 , n379844 );
not ( n53180 , n39050 );
or ( n53181 , n19577 , n22428 );
nand ( n53182 , n53181 , n383597 );
nor ( n53183 , n53180 , n19201 , n53182 , n383607 );
nand ( n53184 , n50642 , n53183 );
buf ( n53185 , n53184 );
buf ( n53186 , n381872 );
or ( n53187 , n31149 , n384057 );
and ( n53188 , n31161 , n384169 );
or ( n53189 , n384182 , n17664 );
or ( n53190 , n32452 , n384190 );
or ( n53191 , n384180 , n31184 );
nand ( n53192 , n53189 , n53190 , n53191 );
nor ( n53193 , n53188 , n53192 );
nand ( n53194 , n53187 , n53193 );
buf ( n53195 , n53194 );
buf ( n53196 , n22406 );
buf ( n53197 , n379844 );
not ( n53198 , n42765 );
not ( n53199 , n31120 );
or ( n53200 , n53198 , n53199 );
and ( n53201 , n384022 , RI15b622e0_1215);
not ( n53202 , n386975 );
not ( n53203 , n38475 );
or ( n53204 , n53202 , n53203 );
or ( n53205 , n38475 , n386975 );
nand ( n53206 , n53204 , n53205 );
and ( n53207 , n384025 , n53206 );
nor ( n53208 , n53201 , n53207 );
nand ( n53209 , n53200 , n53208 );
buf ( n53210 , n53209 );
buf ( n53211 , n31033 );
buf ( n53212 , n22738 );
buf ( n53213 , RI15b47940_307);
buf ( n53214 , n22653 );
and ( n53215 , n30908 , RI15b4a910_409);
and ( n53216 , n51862 , n22217 );
not ( n53217 , n19809 );
and ( n53218 , n53217 , n19673 );
not ( n53219 , n53217 );
and ( n53220 , n53219 , RI15b4a910_409);
nor ( n53221 , n53218 , n53220 );
and ( n53222 , n53221 , n20637 );
nor ( n53223 , n53215 , n53216 , n53222 );
nand ( n53224 , n39991 , n53223 );
buf ( n53225 , n53224 );
buf ( n53226 , n32255 );
buf ( n53227 , n33250 );
not ( n53228 , n19628 );
buf ( n53229 , n386913 );
not ( n53230 , n53229 );
or ( n53231 , n53228 , n53230 );
not ( n53232 , n386945 );
not ( n53233 , n53232 );
not ( n53234 , n53233 );
nand ( n53235 , n53231 , n53234 );
nand ( n53236 , n53235 , n386778 );
buf ( n53237 , n386991 );
nor ( n53238 , n53237 , n387006 );
or ( n53239 , n53238 , n383409 );
nand ( n53240 , n53239 , RI15b62790_1225);
not ( n53241 , n53237 );
nand ( n53242 , n47516 , n48283 );
nor ( n53243 , n53241 , n53242 );
nor ( n53244 , n53123 , n379445 );
or ( n53245 , n53114 , n49459 , RI15b64590_1289);
or ( n53246 , n19598 , n386774 );
nand ( n53247 , n53245 , n53246 );
nor ( n53248 , n53243 , n53244 , n53247 );
not ( n53249 , n53229 );
nor ( n53250 , n48004 , n386778 );
nand ( n53251 , n53249 , n53250 );
nand ( n53252 , n53236 , n53240 , n53248 , n53251 );
buf ( n53253 , n53252 );
buf ( n53254 , n381872 );
or ( n53255 , n32430 , n50737 );
and ( n53256 , n386637 , RI15b54f78_764);
and ( n53257 , n51482 , n32437 );
not ( n53258 , RI15b54f78_764);
not ( n53259 , n382649 );
not ( n53260 , n53259 );
or ( n53261 , n53258 , n53260 );
or ( n53262 , n53259 , RI15b54f78_764);
nand ( n53263 , n53261 , n53262 );
and ( n53264 , n382627 , n53263 );
nor ( n53265 , n53256 , n53257 , n53264 );
and ( n53266 , n50741 , n53265 );
nand ( n53267 , n53255 , n53266 );
buf ( n53268 , n53267 );
not ( n53269 , n386590 );
not ( n53270 , n37629 );
or ( n53271 , n53269 , n53270 );
and ( n53272 , n37637 , n386603 );
not ( n53273 , RI15b59f28_934);
or ( n53274 , n386612 , n53273 );
or ( n53275 , n50208 , n386624 );
or ( n53276 , n386610 , n37646 );
nand ( n53277 , n53274 , n53275 , n53276 );
nor ( n53278 , n53272 , n53277 );
nand ( n53279 , n53271 , n53278 );
buf ( n53280 , n53279 );
buf ( n53281 , n384996 );
buf ( n53282 , n381490 );
buf ( n53283 , n383174 );
nor ( n53284 , n50508 , n383152 );
or ( n53285 , n53284 , n38288 );
nand ( n53286 , n53285 , n50513 );
nand ( n53287 , n50508 , n50512 , n383143 );
and ( n53288 , n383170 , RI15b54078_732);
and ( n53289 , n383147 , RI15b52a70_685);
nor ( n53290 , n53288 , n53289 );
nand ( n53291 , n53286 , n53287 , n53290 );
buf ( n53292 , n53291 );
not ( n53293 , n382976 );
not ( n53294 , n37629 );
or ( n53295 , n53293 , n53294 );
and ( n53296 , n37637 , n382983 );
or ( n53297 , n382995 , n18555 );
or ( n53298 , n37644 , n383001 );
or ( n53299 , n382993 , n37646 );
nand ( n53300 , n53297 , n53298 , n53299 );
nor ( n53301 , n53296 , n53300 );
nand ( n53302 , n53295 , n53301 );
buf ( n53303 , n53302 );
buf ( n53304 , n17499 );
buf ( n53305 , n22343 );
buf ( n53306 , n382071 );
not ( n53307 , RI15b55e00_795);
not ( n53308 , n380000 );
or ( n53309 , n53307 , n53308 );
and ( n53310 , n47789 , n381696 );
not ( n53311 , RI15b55e00_795);
not ( n53312 , n379965 );
or ( n53313 , n53311 , n53312 );
or ( n53314 , n379965 , RI15b55e00_795);
nand ( n53315 , n53313 , n53314 );
and ( n53316 , n379949 , n53315 );
nor ( n53317 , n53310 , n53316 );
nand ( n53318 , n53309 , n53317 );
buf ( n53319 , n53318 );
not ( n53320 , n381570 );
not ( n53321 , n382912 );
or ( n53322 , n53320 , n53321 );
and ( n53323 , n382931 , n381599 );
or ( n53324 , n381609 , n19090 );
or ( n53325 , n40296 , n381619 );
or ( n53326 , n381607 , n382967 );
nand ( n53327 , n53324 , n53325 , n53326 );
nor ( n53328 , n53323 , n53327 );
nand ( n53329 , n53322 , n53328 );
buf ( n53330 , n53329 );
buf ( n53331 , n386760 );
buf ( n53332 , n381490 );
buf ( n53333 , n382067 );
and ( n53334 , n32747 , RI15b42828_134);
and ( n53335 , n32753 , RI15b41568_94);
and ( n53336 , n32762 , RI15b411a8_86);
nor ( n53337 , n53335 , n53336 );
and ( n53338 , n32755 , RI15b41928_102);
and ( n53339 , n32759 , RI15b40de8_78);
nor ( n53340 , n53338 , n53339 );
and ( n53341 , n32771 , RI15b43728_166);
and ( n53342 , n32773 , RI15b42be8_142);
nor ( n53343 , n53341 , n53342 );
and ( n53344 , n32766 , RI15b43368_158);
and ( n53345 , n32768 , RI15b42fa8_150);
nor ( n53346 , n53344 , n53345 );
nand ( n53347 , n53337 , n53340 , n53343 , n53346 );
and ( n53348 , n32750 , n53347 );
and ( n53349 , n32781 , RI15b402a8_54);
nor ( n53350 , n53334 , n53348 , n53349 );
and ( n53351 , n32785 , RI15b42468_126);
and ( n53352 , n32787 , RI15b420a8_118);
nor ( n53353 , n53351 , n53352 );
and ( n53354 , n32792 , RI15b3fee8_46);
and ( n53355 , n32794 , RI15b41ce8_110);
nor ( n53356 , n53354 , n53355 );
and ( n53357 , n32797 , RI15b40668_62);
and ( n53358 , n32800 , RI15b40a28_70);
nor ( n53359 , n53357 , n53358 );
nand ( n53360 , n53350 , n53353 , n53356 , n53359 );
and ( n53361 , n53360 , n41715 );
and ( n53362 , n35335 , RI15b65c10_1337);
not ( n53363 , RI15b48840_339);
not ( n53364 , n35345 );
not ( n53365 , n53364 );
or ( n53366 , n53363 , n53365 );
or ( n53367 , n53364 , RI15b48840_339);
nand ( n53368 , n53366 , n53367 );
and ( n53369 , n35363 , n53368 );
xnor ( n53370 , n53361 , n53362 , n53369 );
nand ( n53371 , n35187 , RI15b48840_339);
and ( n53372 , n52712 , n53370 , n53371 );
buf ( n53373 , n53372 );
buf ( n53374 , n22716 );
buf ( n53375 , n22716 );
buf ( n53376 , n382073 );
or ( n53377 , n381015 , n384945 );
nand ( n53378 , n381017 , RI15b54168_734);
nand ( n53379 , n53377 , n53378 );
not ( n53380 , n53379 );
not ( n53381 , n382061 );
nor ( n53382 , n53381 , n42432 );
buf ( n53383 , n53382 );
buf ( n53384 , n22404 );
buf ( n53385 , n31033 );
buf ( n53386 , n382065 );
buf ( n53387 , n22007 );
buf ( n53388 , n380942 );
nor ( n53389 , n22315 , n35957 );
and ( n53390 , n22326 , n36986 );
or ( n53391 , n35967 , n381058 );
or ( n53392 , n22334 , n35973 );
or ( n53393 , n35965 , n22336 );
nand ( n53394 , n53391 , n53392 , n53393 );
nor ( n53395 , n53390 , n53394 );
nand ( n53396 , n53389 , n53395 );
buf ( n53397 , n53396 );
or ( n53398 , n22102 , n35930 );
and ( n53399 , n22203 , n35935 );
not ( n53400 , RI15b40fc8_82);
or ( n53401 , n35946 , n53400 );
or ( n53402 , n22293 , n35950 );
or ( n53403 , n35944 , n22299 );
nand ( n53404 , n53401 , n53402 , n53403 );
nor ( n53405 , n53399 , n53404 );
nand ( n53406 , n53398 , n53405 );
buf ( n53407 , n53406 );
buf ( n53408 , n384218 );
buf ( n53409 , n22408 );
buf ( n53410 , n22714 );
buf ( n53411 , n22740 );
buf ( n53412 , n22738 );
or ( n53413 , n383814 , n38825 );
and ( n53414 , n383857 , n38828 );
or ( n53415 , n38837 , n21108 );
or ( n53416 , n41182 , n38841 );
or ( n53417 , n38835 , n383917 );
nand ( n53418 , n53415 , n53416 , n53417 );
nor ( n53419 , n53414 , n53418 );
nand ( n53420 , n53413 , n53419 );
buf ( n53421 , n53420 );
buf ( n53422 , n385112 );
not ( n53423 , n387001 );
not ( n53424 , n384025 );
or ( n53425 , n53423 , n53424 );
nand ( n53426 , n53425 , n38494 );
nor ( n53427 , n384024 , RI15b62a60_1231);
nor ( n53428 , n53426 , n53427 );
or ( n53429 , n53428 , n383406 );
nor ( n53430 , n38168 , n387001 , RI15b62ad8_1232);
nand ( n53431 , n38499 , n53430 );
nand ( n53432 , n53429 , n53431 );
buf ( n53433 , n53432 );
buf ( n53434 , n381021 );
buf ( n53435 , RI15b47d00_315);
buf ( n53436 , n22738 );
and ( n53437 , n30908 , RI15b4a820_407);
and ( n53438 , n45189 , n22217 );
and ( n53439 , n19669 , n19670 );
not ( n53440 , n19669 );
and ( n53441 , n53440 , RI15b4a820_407);
nor ( n53442 , n53439 , n53441 );
and ( n53443 , n53442 , n20637 );
nor ( n53444 , n53437 , n53438 , n53443 );
nand ( n53445 , n41306 , n53444 );
buf ( n53446 , n53445 );
buf ( n53447 , n32160 );
buf ( n53448 , n386762 );
buf ( n53449 , n384199 );
not ( n53450 , n386915 );
nor ( n53451 , n53450 , n22473 );
or ( n53452 , n53451 , n386945 );
nand ( n53453 , n53452 , n386771 );
not ( n53454 , n386994 );
nor ( n53455 , n53454 , n387004 );
or ( n53456 , n53455 , n383409 );
nand ( n53457 , n53456 , RI15b62880_1227);
nor ( n53458 , n383482 , RI15b62880_1227);
and ( n53459 , n53454 , n53458 );
not ( n53460 , RI15b64680_1291);
or ( n53461 , n30848 , n49459 );
nand ( n53462 , n53461 , n22425 );
not ( n53463 , n53462 );
or ( n53464 , n53460 , n53463 );
and ( n53465 , n30848 , n22450 , n379448 );
and ( n53466 , n19599 , RI15b63780_1259);
nor ( n53467 , n53465 , n53466 );
nand ( n53468 , n53464 , n53467 );
nor ( n53469 , n53459 , n53468 );
not ( n53470 , n387011 );
nor ( n53471 , n53470 , n386771 );
nand ( n53472 , n53450 , n53471 );
nand ( n53473 , n53453 , n53457 , n53469 , n53472 );
buf ( n53474 , n53473 );
not ( n53475 , n39007 );
and ( n53476 , n53475 , RI15b4b6a8_438);
buf ( n53477 , n19969 );
not ( n53478 , n53477 );
not ( n53479 , n22377 );
or ( n53480 , n53478 , n53479 );
nand ( n53481 , n53480 , n383364 );
and ( n53482 , n53481 , RI15b498a8_374);
or ( n53483 , n22359 , n53477 , RI15b498a8_374);
not ( n53484 , RI15b4b630_437);
and ( n53485 , n53484 , RI15b4b6a8_438);
not ( n53486 , RI15b4b630_437);
nor ( n53487 , n38997 , n53486 , RI15b4b6a8_438);
nor ( n53488 , n53485 , n53487 );
or ( n53489 , n20564 , n53488 );
nand ( n53490 , n53483 , n53489 );
nor ( n53491 , n53476 , n53482 , n53490 );
or ( n53492 , n53491 , n20519 );
not ( n53493 , n19797 );
not ( n53494 , n19789 );
not ( n53495 , n19918 );
and ( n53496 , n53494 , n53495 );
nor ( n53497 , n53496 , n47986 );
or ( n53498 , n53493 , n53497 );
and ( n53499 , n383353 , n19789 , n53493 );
or ( n53500 , n20639 , n382106 );
or ( n53501 , n19790 , n22390 );
nand ( n53502 , n53500 , n53501 , n52512 );
nor ( n53503 , n53499 , n53502 );
nand ( n53504 , n53492 , n53498 , n53503 );
buf ( n53505 , n53504 );
buf ( n53506 , n380865 );
buf ( n53507 , n386563 );
buf ( n53508 , n22716 );
buf ( n53509 , n379893 );
not ( n53510 , n383425 );
not ( n53511 , n381497 );
or ( n53512 , n53510 , n53511 );
nand ( n53513 , n53512 , n384642 );
nand ( n53514 , n53513 , RI15b637f8_1260);
and ( n53515 , n386922 , n19630 );
nor ( n53516 , n383425 , RI15b637f8_1260);
and ( n53517 , n384655 , n53516 );
nor ( n53518 , n53515 , n53517 );
nand ( n53519 , n49850 , n53514 , n53518 );
buf ( n53520 , n53519 );
buf ( n53521 , n380940 );
and ( n53522 , n22646 , RI15b45960_239);
and ( n53523 , n22648 , RI15b51dc8_658);
nor ( n53524 , n53522 , n53523 );
not ( n53525 , n53524 );
buf ( n53526 , n53525 );
or ( n53527 , n22102 , n36200 );
and ( n53528 , n22203 , n36202 );
or ( n53529 , n36212 , n385505 );
or ( n53530 , n22293 , n36217 );
or ( n53531 , n36210 , n22299 );
nand ( n53532 , n53529 , n53530 , n53531 );
nor ( n53533 , n53528 , n53532 );
nand ( n53534 , n53527 , n53533 );
buf ( n53535 , n53534 );
buf ( n53536 , n381566 );
buf ( n53537 , n22788 );
buf ( n53538 , n22714 );
buf ( n53539 , n386563 );
not ( n53540 , RI15b49d58_384);
or ( n53541 , n381056 , n53540 );
or ( n53542 , n32807 , n35454 );
not ( n53543 , n37124 );
and ( n53544 , n53543 , RI15b49d58_384);
not ( n53545 , n53543 );
and ( n53546 , n53545 , n53540 );
nor ( n53547 , n53544 , n53546 );
or ( n53548 , n42690 , n53547 );
nand ( n53549 , n53541 , n53542 , n53548 );
buf ( n53550 , n53549 );
buf ( n53551 , n22479 );
buf ( n53552 , n19655 );
buf ( n53553 , n380906 );
not ( n53554 , RI15b53b50_721);
not ( n53555 , n32244 );
or ( n53556 , n53554 , n53555 );
and ( n53557 , n32247 , RI15b65148_1314);
and ( n53558 , n32249 , RI15b5ffb8_1140);
nor ( n53559 , n53557 , n53558 );
nand ( n53560 , n53556 , n53559 );
buf ( n53561 , n53560 );
buf ( n53562 , n31719 );
buf ( n53563 , n381081 );
or ( n53564 , n381056 , n52595 );
not ( n53565 , n381075 );
not ( n53566 , n53565 );
not ( n53567 , n52598 );
and ( n53568 , n53566 , n53567 );
and ( n53569 , n386555 , RI15b3ff60_47);
nor ( n53570 , n53568 , n53569 );
nand ( n53571 , n53564 , n53570 );
buf ( n53572 , n53571 );
buf ( n53573 , n22738 );
buf ( n53574 , n22402 );
or ( n53575 , n39265 , n22020 );
nand ( n53576 , n35525 , RI15b535b0_709);
nand ( n53577 , n53575 , n53576 );
buf ( n53578 , n53577 );
and ( n53579 , n385164 , RI15b50c70_621);
or ( n53580 , n33651 , n36677 );
or ( n53581 , n36658 , n385170 );
or ( n53582 , n36624 , n385178 );
nand ( n53583 , n53580 , n53581 , n53582 );
nor ( n53584 , n53579 , n53583 );
nand ( n53585 , n47271 , n53584 );
buf ( n53586 , n53585 );
buf ( n53587 , n22408 );
buf ( n53588 , n381006 );
not ( n53589 , n46282 );
nand ( n53590 , n53589 , n379785 );
not ( n53591 , n53590 );
not ( n53592 , n46287 );
or ( n53593 , n53591 , n53592 );
buf ( n53594 , n46283 );
buf ( n53595 , n53594 );
nand ( n53596 , n53593 , n53595 );
nor ( n53597 , n53589 , n53594 );
nand ( n53598 , n36580 , n53597 );
and ( n53599 , n34529 , n34543 );
not ( n53600 , n34529 );
not ( n53601 , n34543 );
and ( n53602 , n53600 , n53601 );
nor ( n53603 , n53599 , n53602 );
and ( n53604 , n53603 , n46302 );
not ( n53605 , RI15b5e230_1077);
not ( n53606 , n34651 );
or ( n53607 , n53605 , n53606 );
or ( n53608 , n36518 , n379440 );
nand ( n53609 , n53607 , n53608 );
nor ( n53610 , n53604 , n53609 );
nand ( n53611 , n53596 , n53598 , n53610 );
buf ( n53612 , n53611 );
buf ( n53613 , n379802 );
or ( n53614 , n380968 , n38373 );
and ( n53615 , n380986 , n38375 );
or ( n53616 , n38385 , n20337 );
or ( n53617 , n380994 , n38389 );
or ( n53618 , n38383 , n380996 );
nand ( n53619 , n53616 , n53617 , n53618 );
nor ( n53620 , n53615 , n53619 );
nand ( n53621 , n53614 , n53620 );
buf ( n53622 , n53621 );
buf ( n53623 , n379847 );
buf ( n53624 , n18226 );
buf ( n53625 , n22653 );
buf ( n53626 , RI15b5dc18_1064);
or ( n53627 , n36937 , n386706 );
and ( n53628 , n36946 , n386718 );
not ( n53629 , RI15b4d0e8_494);
or ( n53630 , n386727 , n53629 );
or ( n53631 , n39875 , n386735 );
or ( n53632 , n386725 , n36955 );
nand ( n53633 , n53630 , n53631 , n53632 );
nor ( n53634 , n53628 , n53633 );
nand ( n53635 , n53627 , n53634 );
buf ( n53636 , n53635 );
buf ( n53637 , n381707 );
buf ( n53638 , n386760 );
or ( n53639 , n384021 , n386958 );
or ( n53640 , n19084 , n386747 );
not ( n53641 , n384029 );
and ( n53642 , n53641 , RI15b61db8_1204);
not ( n53643 , n53641 );
and ( n53644 , n53643 , n386958 );
nor ( n53645 , n53642 , n53644 );
or ( n53646 , n53645 , n384024 );
nand ( n53647 , n53639 , n53640 , n53646 );
buf ( n53648 , n53647 );
buf ( n53649 , n384199 );
or ( n53650 , n41015 , n381949 );
nand ( n53651 , n379832 , RI15b46c98_280);
nand ( n53652 , n53650 , n50434 , n53651 );
buf ( n53653 , n53652 );
buf ( n53654 , n22402 );
buf ( n53655 , n32255 );
buf ( n53656 , n17499 );
buf ( n53657 , n382071 );
not ( n53658 , n32610 );
and ( n53659 , n53658 , RI15b4b978_444);
not ( n53660 , n22377 );
buf ( n53661 , n19979 );
not ( n53662 , n53661 );
or ( n53663 , n53660 , n53662 );
nand ( n53664 , n53663 , n383364 );
and ( n53665 , n53664 , RI15b49b78_380);
or ( n53666 , n53661 , n22359 , RI15b49b78_380);
and ( n53667 , n382114 , RI15b4b978_444);
nor ( n53668 , n20549 , n382114 , RI15b4b978_444);
nor ( n53669 , n53667 , n53668 );
or ( n53670 , n20564 , n53669 );
nand ( n53671 , n53666 , n53670 );
nor ( n53672 , n53659 , n53665 , n53671 );
or ( n53673 , n53672 , n20519 );
buf ( n53674 , n19721 );
not ( n53675 , n19831 );
not ( n53676 , n53675 );
not ( n53677 , n19918 );
and ( n53678 , n53676 , n53677 );
nor ( n53679 , n53678 , n384684 );
or ( n53680 , n53674 , n53679 );
and ( n53681 , n383353 , n53674 , n53675 );
or ( n53682 , n20639 , n382115 );
or ( n53683 , n19717 , n22390 );
nand ( n53684 , n53682 , n53683 , n384692 );
nor ( n53685 , n53681 , n53684 );
nand ( n53686 , n53673 , n53680 , n53685 );
buf ( n53687 , n53686 );
buf ( n53688 , n382537 );
buf ( n53689 , n22402 );
buf ( n53690 , n384700 );
buf ( n53691 , n380203 );
and ( n53692 , n384641 , RI15b63528_1254);
and ( n53693 , n386905 , n19630 );
and ( n53694 , n384655 , n386902 );
nor ( n53695 , n53692 , n53693 , n53694 );
nand ( n53696 , n51738 , n53695 );
buf ( n53697 , n53696 );
buf ( n53698 , n32981 );
buf ( n53699 , n21800 );
not ( n53700 , RI15b473a0_295);
not ( n53701 , n385213 );
or ( n53702 , n53700 , n53701 );
and ( n53703 , n385221 , RI15b48930_341);
and ( n53704 , n20631 , RI15b46c20_279);
nor ( n53705 , n53703 , n53704 );
nand ( n53706 , n53702 , n53705 );
buf ( n53707 , n53706 );
buf ( n53708 , n379844 );
buf ( n53709 , n22653 );
buf ( n53710 , n382065 );
buf ( n53711 , RI15b47760_303);
buf ( n53712 , n381021 );
and ( n53713 , n30908 , RI15b4a988_410);
or ( n53714 , n44601 , n22216 );
not ( n53715 , n19816 );
and ( n53716 , n53715 , RI15b4a988_410);
not ( n53717 , n53715 );
and ( n53718 , n53717 , n19820 );
nor ( n53719 , n53716 , n53718 );
or ( n53720 , n53719 , n20638 );
nand ( n53721 , n53714 , n53720 );
nor ( n53722 , n53713 , n53721 );
nand ( n53723 , n52517 , n53722 );
buf ( n53724 , n53723 );
buf ( n53725 , n382049 );
buf ( n53726 , n31030 );
not ( n53727 , n387005 );
buf ( n53728 , n386989 );
not ( n53729 , n53728 );
or ( n53730 , n53727 , n53729 );
nand ( n53731 , n53730 , n383408 );
and ( n53732 , n53731 , RI15b62718_1224);
or ( n53733 , n53728 , n383482 , RI15b62718_1224);
not ( n53734 , n30844 );
or ( n53735 , n53734 , n379708 , RI15b64518_1288);
or ( n53736 , n379711 , RI15b644a0_1287);
nand ( n53737 , n53735 , n53736 );
and ( n53738 , n53737 , n22450 );
and ( n53739 , n19599 , RI15b63618_1256);
nor ( n53740 , n53738 , n53739 );
nand ( n53741 , n53733 , n53740 );
nor ( n53742 , n53732 , n53741 );
buf ( n53743 , n386907 );
nor ( n53744 , n53743 , n22473 );
or ( n53745 , n53744 , n53233 );
nand ( n53746 , n53745 , n386912 );
not ( n53747 , n386912 );
nand ( n53748 , n53747 , n53743 , n48005 );
and ( n53749 , n22450 , n53734 );
nor ( n53750 , n53749 , n22426 );
not ( n53751 , n53750 );
nand ( n53752 , n53751 , RI15b64518_1288);
nand ( n53753 , n53742 , n53746 , n53748 , n53752 );
buf ( n53754 , n53753 );
buf ( n53755 , n35649 );
not ( n53756 , RI15b53448_706);
not ( n53757 , n383170 );
or ( n53758 , n53756 , n53757 );
and ( n53759 , n33453 , RI15b549d8_752);
and ( n53760 , n383147 , RI15b52cc8_690);
nor ( n53761 , n53759 , n53760 );
nand ( n53762 , n53758 , n53761 );
buf ( n53763 , n53762 );
not ( n53764 , n35983 );
not ( n53765 , n33400 );
or ( n53766 , n53764 , n53765 );
and ( n53767 , n33415 , n35987 );
or ( n53768 , n35996 , n18504 );
or ( n53769 , n36293 , n36003 );
or ( n53770 , n35994 , n33443 );
nand ( n53771 , n53768 , n53769 , n53770 );
nor ( n53772 , n53767 , n53771 );
nand ( n53773 , n53766 , n53772 );
buf ( n53774 , n53773 );
buf ( n53775 , n19655 );
buf ( n53776 , RI15b5e578_1084);
or ( n53777 , n31149 , n36242 );
and ( n53778 , n31161 , n43075 );
not ( n53779 , RI15b4d340_499);
or ( n53780 , n36250 , n53779 );
or ( n53781 , n32452 , n36254 );
or ( n53782 , n36248 , n31184 );
nand ( n53783 , n53780 , n53781 , n53782 );
nor ( n53784 , n53778 , n53783 );
nand ( n53785 , n53777 , n53784 );
buf ( n53786 , n53785 );
buf ( n53787 , n381021 );
buf ( n53788 , n381006 );
not ( n53789 , n45125 );
not ( n53790 , n48601 );
not ( n53791 , n53790 );
or ( n53792 , n53789 , n53791 );
nand ( n53793 , n53792 , n51156 );
not ( n53794 , n53793 );
or ( n53795 , n53794 , n45131 );
and ( n53796 , n51158 , n45131 , RI15b61ae8_1198);
not ( n53797 , n38783 );
nor ( n53798 , n53797 , n38813 );
not ( n53799 , n53798 );
and ( n53800 , n38502 , RI15b59dc0_931);
and ( n53801 , n38506 , RI15b5bf80_1003);
nor ( n53802 , n53800 , n53801 );
and ( n53803 , n38509 , RI15b5a180_939);
and ( n53804 , n38512 , RI15b5bbc0_995);
nor ( n53805 , n53803 , n53804 );
and ( n53806 , n38515 , RI15b5a540_947);
and ( n53807 , n38517 , RI15b5acc0_963);
nor ( n53808 , n53806 , n53807 );
and ( n53809 , n38794 , RI15b5b440_979);
and ( n53810 , n38525 , RI15b5c340_1011);
nor ( n53811 , n53809 , n53810 );
nand ( n53812 , n53802 , n53805 , n53808 , n53811 );
and ( n53813 , n38529 , RI15b5b800_987);
and ( n53814 , n38531 , RI15b5b080_971);
nor ( n53815 , n53813 , n53814 );
and ( n53816 , n38534 , RI15b59a00_923);
and ( n53817 , n38536 , RI15b5a900_955);
nor ( n53818 , n53816 , n53817 );
and ( n53819 , n38539 , RI15b58b00_891);
and ( n53820 , n38541 , RI15b59640_915);
nor ( n53821 , n53819 , n53820 );
and ( n53822 , n38544 , RI15b58ec0_899);
and ( n53823 , n38809 , RI15b59280_907);
nor ( n53824 , n53822 , n53823 );
nand ( n53825 , n53815 , n53818 , n53821 , n53824 );
nor ( n53826 , n53812 , n53825 );
not ( n53827 , n53826 );
and ( n53828 , n53799 , n53827 );
and ( n53829 , n53798 , n53826 );
nor ( n53830 , n53828 , n53829 );
or ( n53831 , n53830 , n46087 );
or ( n53832 , n380562 , n31052 );
nand ( n53833 , n53831 , n53832 , n45144 );
nor ( n53834 , n53796 , n53833 );
nand ( n53835 , n53795 , n53834 );
buf ( n53836 , n53835 );
buf ( n53837 , n18226 );
buf ( n53838 , n30992 );
not ( n53839 , n52119 );
not ( n53840 , n384726 );
or ( n53841 , n53839 , n53840 );
and ( n53842 , n35477 , n48939 );
or ( n53843 , n48948 , n20786 );
or ( n53844 , n51233 , n48953 );
or ( n53845 , n48946 , n384759 );
nand ( n53846 , n53843 , n53844 , n53845 );
nor ( n53847 , n53842 , n53846 );
nand ( n53848 , n53841 , n53847 );
buf ( n53849 , n53848 );
buf ( n53850 , n380942 );
nor ( n53851 , n45668 , n45676 );
and ( n53852 , n383505 , n53851 );
nor ( n53853 , n53852 , n383577 );
or ( n53854 , n32291 , n383523 );
and ( n53855 , n53854 , RI15b61458_1184);
not ( n53856 , n53854 );
and ( n53857 , n53856 , n32280 );
nor ( n53858 , n53855 , n53857 );
or ( n53859 , n53853 , n53858 );
and ( n53860 , n383601 , RI15b5fec8_1138);
not ( n53861 , n53858 );
nor ( n53862 , n53861 , n53851 );
and ( n53863 , n383603 , n53862 );
and ( n53864 , n383607 , RI15b5f748_1122);
nor ( n53865 , n53860 , n53863 , n53864 );
nand ( n53866 , n53859 , n53865 );
buf ( n53867 , n53866 );
buf ( n53868 , n30992 );
buf ( n53869 , n32981 );
buf ( n53870 , n32255 );
not ( n53871 , n46036 );
not ( n53872 , n34930 );
and ( n53873 , n53871 , n53872 );
nor ( n53874 , n53873 , n35114 );
or ( n53875 , n53874 , n35088 );
and ( n53876 , n35118 , n46040 );
and ( n53877 , n20631 , RI15b461d0_257);
nor ( n53878 , n53876 , n53877 );
nand ( n53879 , n385213 , RI15b477d8_304);
nand ( n53880 , n53875 , n53878 , n53879 );
buf ( n53881 , n53880 );
buf ( n53882 , n33382 );
buf ( n53883 , n380203 );
or ( n53884 , n386705 , n35622 );
and ( n53885 , n386716 , n35625 );
not ( n53886 , RI15b4f5f0_573);
or ( n53887 , n35635 , n53886 );
or ( n53888 , n386732 , n35640 );
or ( n53889 , n35633 , n386738 );
nand ( n53890 , n53887 , n53888 , n53889 );
nor ( n53891 , n53885 , n53890 );
nand ( n53892 , n53884 , n53891 );
buf ( n53893 , n53892 );
buf ( n53894 , n22714 );
buf ( n53895 , n384996 );
not ( n53896 , RI15b5f8b0_1125);
not ( n53897 , n383601 );
or ( n53898 , n53896 , n53897 );
and ( n53899 , n383505 , RI15b60e40_1171);
and ( n53900 , n383607 , RI15b5f130_1109);
nor ( n53901 , n53899 , n53900 );
nand ( n53902 , n53898 , n53901 );
buf ( n53903 , n53902 );
buf ( n53904 , n36704 );
or ( n53905 , n383814 , n35622 );
and ( n53906 , n383857 , n35625 );
or ( n53907 , n35635 , n21158 );
or ( n53908 , n41182 , n35640 );
or ( n53909 , n35633 , n383917 );
nand ( n53910 , n53907 , n53908 , n53909 );
nor ( n53911 , n53906 , n53910 );
nand ( n53912 , n53905 , n53911 );
buf ( n53913 , n53912 );
buf ( n53914 , n36704 );
buf ( n53915 , n22343 );
not ( n53916 , RI15b5fa18_1128);
not ( n53917 , n383601 );
or ( n53918 , n53916 , n53917 );
and ( n53919 , n383505 , RI15b60fa8_1174);
and ( n53920 , n383607 , RI15b5f298_1112);
nor ( n53921 , n53919 , n53920 );
nand ( n53922 , n53918 , n53921 );
buf ( n53923 , n53922 );
buf ( n53924 , n387159 );
and ( n53925 , n22646 , RI15b45c30_245);
and ( n53926 , n22648 , RI15b52098_664);
nor ( n53927 , n53925 , n53926 );
not ( n53928 , n53927 );
buf ( n53929 , n53928 );
buf ( n53930 , n32271 );
not ( n53931 , n39103 );
or ( n53932 , n53931 , RI15b56760_815);
or ( n53933 , n21788 , n36237 );
nand ( n53934 , n53933 , RI15b56760_815);
not ( n53935 , n37718 );
not ( n53936 , n21401 );
and ( n53937 , n53936 , n21402 );
or ( n53938 , n32096 , n21364 );
nand ( n53939 , n53938 , n21409 );
nor ( n53940 , n53937 , n53939 );
not ( n53941 , n53940 );
or ( n53942 , n53935 , n53941 );
or ( n53943 , n53940 , n37718 );
nand ( n53944 , n53942 , n53943 );
and ( n53945 , n21559 , n53944 );
not ( n53946 , n37721 );
not ( n53947 , n53940 );
not ( n53948 , n53947 );
or ( n53949 , n53946 , n53948 );
or ( n53950 , n53947 , n37721 );
nand ( n53951 , n53949 , n53950 );
and ( n53952 , n21740 , n53951 );
and ( n53953 , n21751 , RI15b57660_847);
nor ( n53954 , n53945 , n53952 , n53953 );
nand ( n53955 , n53932 , n53934 , n53954 );
buf ( n53956 , n53955 );
and ( n53957 , n35684 , RI15b58740_883);
buf ( n53958 , n53957 );
buf ( n53959 , n32672 );
buf ( n53960 , n22343 );
buf ( n53961 , n22005 );
not ( n53962 , n379870 );
not ( n53963 , n381481 );
and ( n53964 , n53962 , n53963 );
nor ( n53965 , n53964 , n37707 );
not ( n53966 , n53965 );
not ( n53967 , n381475 );
or ( n53968 , n53966 , n53967 );
nand ( n53969 , n53968 , RI15b54348_738);
and ( n53970 , n33211 , n381477 );
not ( n53971 , n383165 );
nor ( n53972 , n53970 , n50742 , n53971 );
nand ( n53973 , n53969 , n53972 );
buf ( n53974 , n53973 );
not ( n53975 , n33220 );
not ( n53976 , n33400 );
or ( n53977 , n53975 , n53976 );
and ( n53978 , n33415 , n33226 );
or ( n53979 , n33237 , n18471 );
or ( n53980 , n36293 , n33241 );
or ( n53981 , n33235 , n33443 );
nand ( n53982 , n53979 , n53980 , n53981 );
nor ( n53983 , n53978 , n53982 );
nand ( n53984 , n53977 , n53983 );
buf ( n53985 , n53984 );
buf ( n53986 , n17499 );
buf ( n53987 , n33382 );
not ( n53988 , RI15b46068_254);
not ( n53989 , n379832 );
or ( n53990 , n53988 , n53989 );
not ( n53991 , n41015 );
not ( n53992 , n34964 );
and ( n53993 , n53991 , n53992 );
nor ( n53994 , n53993 , n35583 );
nand ( n53995 , n53990 , n53994 );
buf ( n53996 , n53995 );
buf ( n53997 , n21800 );
buf ( n53998 , n22343 );
buf ( n53999 , n382073 );
buf ( n54000 , n31719 );
buf ( n54001 , n380940 );
buf ( n54002 , n381004 );
or ( n54003 , n380968 , n37495 );
and ( n54004 , n380986 , n37498 );
not ( n54005 , RI15b426c0_131);
or ( n54006 , n37507 , n54005 );
or ( n54007 , n380994 , n37512 );
or ( n54008 , n37505 , n380996 );
nand ( n54009 , n54006 , n54007 , n54008 );
nor ( n54010 , n54004 , n54009 );
nand ( n54011 , n54003 , n54010 );
buf ( n54012 , n54011 );
buf ( n54013 , n22007 );
buf ( n54014 , n382073 );
buf ( n54015 , n380203 );
and ( n54016 , n18168 , n35244 );
not ( n54017 , n18164 );
and ( n54018 , n54017 , n18072 );
nor ( n54019 , n54016 , n54018 , n17507 );
nand ( n54020 , n44800 , n54019 );
buf ( n54021 , n54020 );
buf ( n54022 , n381566 );
not ( n54023 , n36558 );
nand ( n54024 , n54023 , n379785 );
not ( n54025 , n54024 );
not ( n54026 , n36574 );
or ( n54027 , n54025 , n54026 );
buf ( n54028 , n36559 );
buf ( n54029 , n54028 );
nand ( n54030 , n54027 , n54029 );
nor ( n54031 , n54023 , n54028 );
nand ( n54032 , n40809 , n54031 );
not ( n54033 , n39191 );
not ( n54034 , n39190 );
not ( n54035 , n54034 );
or ( n54036 , n54033 , n54035 );
or ( n54037 , n54034 , n39191 );
nand ( n54038 , n54036 , n54037 );
and ( n54039 , n54038 , n46302 );
not ( n54040 , RI15b5dd08_1066);
not ( n54041 , n34651 );
or ( n54042 , n54040 , n54041 );
not ( n54043 , RI15b63f00_1275);
or ( n54044 , n36518 , n54043 );
nand ( n54045 , n54042 , n54044 );
nor ( n54046 , n54039 , n54045 );
nand ( n54047 , n54030 , n54032 , n54046 );
buf ( n54048 , n54047 );
not ( n54049 , n35471 );
or ( n54050 , n383814 , n54049 );
and ( n54051 , n383857 , n35479 );
or ( n54052 , n35488 , n21102 );
or ( n54053 , n383908 , n35497 );
or ( n54054 , n35486 , n383917 );
nand ( n54055 , n54052 , n54053 , n54054 );
nor ( n54056 , n54051 , n54055 );
nand ( n54057 , n54050 , n54056 );
buf ( n54058 , n54057 );
buf ( n54059 , n380906 );
buf ( n54060 , n384218 );
or ( n54061 , n31053 , n48871 );
and ( n54062 , n36536 , RI15b61098_1176);
and ( n54063 , n36538 , n18366 );
not ( n54064 , RI15b61098_1176);
not ( n54065 , n31067 );
or ( n54066 , n54064 , n54065 );
or ( n54067 , n31067 , RI15b61098_1176);
nand ( n54068 , n54066 , n54067 );
and ( n54069 , n36541 , n54068 );
nor ( n54070 , n54062 , n54063 , n54069 );
nand ( n54071 , n54061 , n384909 , n54070 );
buf ( n54072 , n54071 );
buf ( n54073 , n382071 );
or ( n54074 , n40390 , n386414 );
not ( n54075 , n39949 );
not ( n54076 , n39939 );
and ( n54077 , n54075 , n54076 );
and ( n54078 , n39949 , n39939 );
nor ( n54079 , n54077 , n54078 );
not ( n54080 , n386018 );
nor ( n54081 , n54079 , n54080 );
not ( n54082 , n386158 );
and ( n54083 , n39963 , n54082 );
nor ( n54084 , n39963 , n54082 );
nor ( n54085 , n54083 , n54084 );
or ( n54086 , n54085 , n386263 );
or ( n54087 , n44685 , n386414 );
nand ( n54088 , n54087 , n41292 );
and ( n54089 , n54088 , n386500 );
and ( n54090 , n22398 , RI15b4b6a8_438);
nor ( n54091 , n54089 , n54090 );
nand ( n54092 , n54086 , n54091 );
nor ( n54093 , n54081 , n54092 );
and ( n54094 , n386540 , RI15b44010_185);
and ( n54095 , n386549 , n385815 );
and ( n54096 , n386556 , n54082 );
nor ( n54097 , n54094 , n54095 , n54096 );
nand ( n54098 , n54074 , n54093 , n54097 );
buf ( n54099 , n54098 );
buf ( n54100 , n22655 );
buf ( n54101 , n385197 );
buf ( n54102 , n22007 );
buf ( n54103 , n386563 );
buf ( n54104 , n379844 );
or ( n54105 , n32259 , n36121 );
and ( n54106 , n384983 , n36123 );
or ( n54107 , n36132 , n385405 );
or ( n54108 , n22022 , n36139 );
or ( n54109 , n36130 , n384988 );
nand ( n54110 , n54107 , n54108 , n54109 );
nor ( n54111 , n54106 , n54110 );
nand ( n54112 , n54105 , n54111 );
buf ( n54113 , n54112 );
buf ( n54114 , n384996 );
buf ( n54115 , n32271 );
buf ( n54116 , n32981 );
buf ( n54117 , n22788 );
buf ( n54118 , n44220 );
or ( n54119 , n381407 , n54118 );
nand ( n54120 , n381417 , n381290 );
or ( n54121 , n381424 , n33463 );
nand ( n54122 , n54121 , n381450 );
and ( n54123 , n54122 , n33474 );
and ( n54124 , n381461 , n33478 );
nor ( n54125 , n54123 , n54124 );
and ( n54126 , n54120 , n54125 );
nand ( n54127 , n381486 , RI15b53088_698);
nand ( n54128 , n54119 , n54126 , n54127 );
buf ( n54129 , n54128 );
not ( n54130 , n381494 );
not ( n54131 , n33400 );
or ( n54132 , n54130 , n54131 );
and ( n54133 , n33415 , n381528 );
or ( n54134 , n381544 , n18453 );
or ( n54135 , n36293 , n381557 );
or ( n54136 , n381542 , n33443 );
nand ( n54137 , n54134 , n54135 , n54136 );
nor ( n54138 , n54133 , n54137 );
nand ( n54139 , n54132 , n54138 );
buf ( n54140 , n54139 );
buf ( n54141 , n21800 );
and ( n54142 , n22646 , RI15b45690_233);
and ( n54143 , n22648 , RI15b51af8_652);
nor ( n54144 , n54142 , n54143 );
not ( n54145 , n54144 );
buf ( n54146 , n54145 );
buf ( n54147 , n379893 );
not ( n54148 , n45544 );
and ( n54149 , n21788 , RI15b568c8_818);
and ( n54150 , n21767 , n21825 );
buf ( n54151 , n21818 );
not ( n54152 , RI15b568c8_818);
and ( n54153 , n54151 , n54152 );
not ( n54154 , n54151 );
and ( n54155 , n54154 , RI15b568c8_818);
nor ( n54156 , n54153 , n54155 );
and ( n54157 , n21794 , n54156 );
nor ( n54158 , n54149 , n54150 , n54157 );
nand ( n54159 , n54148 , n54158 );
buf ( n54160 , n54159 );
nor ( n54161 , n35684 , n19640 );
or ( n54162 , n54161 , n19261 );
or ( n54163 , RI15b585d8_880 , n22775 );
not ( n54164 , n35154 );
nor ( n54165 , n54164 , n380737 );
or ( n54166 , n54165 , n380788 );
nand ( n54167 , n54162 , n54163 , n54166 );
buf ( n54168 , n54167 );
buf ( n54169 , n22738 );
buf ( n54170 , n380942 );
buf ( n54171 , n32676 );
buf ( n54172 , n20665 );
nor ( n54173 , n32950 , n32938 , n32944 );
nand ( n54174 , n51179 , n54173 );
or ( n54175 , n54174 , n382079 );
not ( n54176 , n43099 );
nand ( n54177 , n54175 , n54176 );
or ( n54178 , n382473 , n32967 );
nand ( n54179 , n54178 , n22725 );
nand ( n54180 , n54177 , n54179 );
not ( n54181 , n32929 );
nor ( n54182 , n54181 , n54179 );
and ( n54183 , n54174 , n54182 );
not ( n54184 , RI15b45e10_249);
not ( n54185 , n32975 );
or ( n54186 , n54184 , n54185 );
not ( n54187 , n46999 );
nand ( n54188 , n54186 , n54187 );
nor ( n54189 , n54183 , n54188 );
nand ( n54190 , n54180 , n54189 );
buf ( n54191 , n54190 );
buf ( n54192 , n31979 );
buf ( n54193 , n22714 );
buf ( n54194 , n31719 );
not ( n54195 , RI15b4a0a0_391);
not ( n54196 , n37135 );
or ( n54197 , n54195 , n54196 );
not ( n54198 , n48996 );
not ( n54199 , n54198 );
not ( n54200 , n48911 );
not ( n54201 , n54200 );
and ( n54202 , n54199 , n54201 );
and ( n54203 , n37422 , n37136 );
nor ( n54204 , n54202 , n54203 );
nand ( n54205 , n54197 , n54204 );
buf ( n54206 , n54205 );
buf ( n54207 , n381490 );
buf ( n54208 , n32255 );
buf ( n54209 , n386563 );
not ( n54210 , RI15b53808_714);
not ( n54211 , n32244 );
or ( n54212 , n54210 , n54211 );
and ( n54213 , n32247 , RI15b64e00_1307);
and ( n54214 , n32249 , RI15b5fc70_1133);
nor ( n54215 , n54213 , n54214 );
nand ( n54216 , n54212 , n54215 );
buf ( n54217 , n54216 );
or ( n54218 , n381056 , n19983 );
not ( n54219 , n46126 );
or ( n54220 , n45380 , n54219 );
not ( n54221 , n37122 );
and ( n54222 , n54221 , RI15b49c68_382);
not ( n54223 , n54221 );
and ( n54224 , n54223 , n19983 );
nor ( n54225 , n54222 , n54224 );
or ( n54226 , n37110 , n54225 );
nand ( n54227 , n54218 , n54220 , n54226 );
buf ( n54228 , n54227 );
buf ( n54229 , n22402 );
buf ( n54230 , n19655 );
buf ( n54231 , n382049 );
buf ( n54232 , n32981 );
not ( n54233 , RI15b53c40_723);
not ( n54234 , n32244 );
or ( n54235 , n54233 , n54234 );
and ( n54236 , n32247 , RI15b65238_1316);
and ( n54237 , n32249 , RI15b600a8_1142);
nor ( n54238 , n54236 , n54237 );
nand ( n54239 , n54235 , n54238 );
buf ( n54240 , n54239 );
buf ( n54241 , n382049 );
and ( n54242 , n30908 , RI15b4a7a8_406);
or ( n54243 , n53493 , n22216 );
and ( n54244 , n19792 , RI15b4a7a8_406);
not ( n54245 , n19792 );
and ( n54246 , n54245 , n19790 );
nor ( n54247 , n54244 , n54246 );
or ( n54248 , n54247 , n20638 );
nand ( n54249 , n54243 , n54248 );
nor ( n54250 , n54242 , n54249 );
nand ( n54251 , n54093 , n54250 );
buf ( n54252 , n54251 );
buf ( n54253 , n35651 );
buf ( n54254 , n382049 );
buf ( n54255 , n19653 );
buf ( n54256 , n386916 );
nor ( n54257 , n54256 , n22473 );
or ( n54258 , n54257 , n386945 );
nand ( n54259 , n54258 , n386922 );
buf ( n54260 , n386996 );
not ( n54261 , n387004 );
not ( n54262 , n54261 );
nor ( n54263 , n54260 , n54262 );
or ( n54264 , n54263 , n383409 );
nand ( n54265 , n54264 , RI15b628f8_1228);
nor ( n54266 , n53470 , n386922 );
nand ( n54267 , n54256 , n54266 );
nor ( n54268 , n383482 , RI15b628f8_1228);
and ( n54269 , n54260 , n54268 );
not ( n54270 , RI15b646f8_1292);
not ( n54271 , n53462 );
or ( n54272 , n54270 , n54271 );
not ( n54273 , RI15b646f8_1292);
not ( n54274 , n379448 );
or ( n54275 , n54273 , n54274 );
nand ( n54276 , n30848 , n379720 , RI15b64680_1291);
nand ( n54277 , n54275 , n54276 );
and ( n54278 , n54277 , n22450 );
and ( n54279 , n19599 , RI15b637f8_1260);
nor ( n54280 , n54278 , n54279 );
nand ( n54281 , n54272 , n54280 );
nor ( n54282 , n54269 , n54281 );
nand ( n54283 , n54259 , n54265 , n54267 , n54282 );
buf ( n54284 , n54283 );
not ( n54285 , n34740 );
nor ( n54286 , n54285 , n386404 );
not ( n54287 , n54286 );
not ( n54288 , n44906 );
nand ( n54289 , n54287 , n54288 );
nand ( n54290 , n54289 , n386500 );
not ( n54291 , n34755 );
and ( n54292 , n54291 , n386194 );
not ( n54293 , n54291 );
and ( n54294 , n54293 , n34756 );
nor ( n54295 , n54292 , n54294 );
and ( n54296 , n54295 , n39973 );
buf ( n54297 , n34770 );
not ( n54298 , n385891 );
and ( n54299 , n54297 , n54298 );
not ( n54300 , n54297 );
and ( n54301 , n54300 , n385891 );
nor ( n54302 , n54299 , n54301 );
not ( n54303 , n386018 );
or ( n54304 , n54302 , n54303 );
nand ( n54305 , n41301 , RI15b4b978_444);
nand ( n54306 , n54304 , n54305 );
nor ( n54307 , n54296 , n54306 );
nand ( n54308 , n54290 , n54307 );
not ( n54309 , n54308 );
and ( n54310 , n40389 , n34741 );
or ( n54311 , n386541 , n385880 );
or ( n54312 , n385891 , n386550 );
or ( n54313 , n386194 , n386557 );
nand ( n54314 , n54311 , n54312 , n54313 );
nor ( n54315 , n54310 , n54314 );
nand ( n54316 , n54309 , n54315 );
buf ( n54317 , n54316 );
buf ( n54318 , n19655 );
buf ( n54319 , n22655 );
buf ( n54320 , n379895 );
buf ( n54321 , n382067 );
buf ( n54322 , n385197 );
buf ( n54323 , n381566 );
or ( n54324 , n380968 , n38065 );
and ( n54325 , n380986 , n38067 );
or ( n54326 , n38077 , n20334 );
or ( n54327 , n380994 , n38081 );
or ( n54328 , n38075 , n380996 );
nand ( n54329 , n54326 , n54327 , n54328 );
nor ( n54330 , n54325 , n54329 );
nand ( n54331 , n54324 , n54330 );
buf ( n54332 , n54331 );
buf ( n54333 , n384203 );
buf ( n54334 , n381872 );
buf ( n54335 , n384203 );
not ( n54336 , RI15b55950_785);
not ( n54337 , n380000 );
or ( n54338 , n54336 , n54337 );
and ( n54339 , n36384 , RI15b4c4b8_468);
not ( n54340 , RI15b55950_785);
not ( n54341 , n379952 );
not ( n54342 , n54341 );
or ( n54343 , n54340 , n54342 );
or ( n54344 , n54341 , RI15b55950_785);
nand ( n54345 , n54343 , n54344 );
and ( n54346 , n379949 , n54345 );
nor ( n54347 , n54339 , n54346 );
nand ( n54348 , n54338 , n54347 );
buf ( n54349 , n54348 );
not ( n54350 , n36395 );
not ( n54351 , n381589 );
or ( n54352 , n54350 , n54351 );
and ( n54353 , n381596 , n36401 );
or ( n54354 , n36410 , n18724 );
or ( n54355 , n381616 , n36416 );
or ( n54356 , n36408 , n381621 );
nand ( n54357 , n54354 , n54355 , n54356 );
nor ( n54358 , n54353 , n54357 );
nand ( n54359 , n54352 , n54358 );
buf ( n54360 , n54359 );
buf ( n54361 , n380940 );
buf ( n54362 , n17499 );
buf ( n54363 , n379893 );
not ( n54364 , RI15b522f0_669);
not ( n54365 , n379397 );
or ( n54366 , n54364 , n54365 );
or ( n54367 , n43293 , RI15b542d0_737);
nand ( n54368 , n54366 , n54367 );
buf ( n54369 , n54368 );
nor ( n54370 , n37581 , n384267 );
not ( n54371 , n54370 );
nand ( n54372 , n54371 , n32543 );
nand ( n54373 , n54372 , n49833 );
nand ( n54374 , n37585 , n384582 );
not ( n54375 , n384577 );
and ( n54376 , n54374 , n54375 );
not ( n54377 , n54374 );
and ( n54378 , n54377 , n384577 );
nor ( n54379 , n54376 , n54378 );
and ( n54380 , n54379 , n49846 );
not ( n54381 , n32567 );
not ( n54382 , n384470 );
not ( n54383 , n54382 );
and ( n54384 , n54381 , n54383 );
and ( n54385 , n32567 , n54382 );
nor ( n54386 , n54384 , n54385 );
or ( n54387 , n54386 , n38921 );
or ( n54388 , n19512 , n379662 );
nand ( n54389 , n54387 , n54388 );
nor ( n54390 , n54380 , n54389 );
nand ( n54391 , n54373 , n54390 );
not ( n54392 , n54391 );
and ( n54393 , n31792 , n384577 );
or ( n54394 , n31771 , n384265 );
or ( n54395 , n384267 , n32378 );
or ( n54396 , n54382 , n31779 );
nand ( n54397 , n54394 , n54395 , n54396 );
nor ( n54398 , n54393 , n54397 );
nand ( n54399 , n54392 , n54398 );
buf ( n54400 , n54399 );
buf ( n54401 , n384700 );
buf ( n54402 , n381566 );
buf ( n54403 , n384700 );
not ( n54404 , n44064 );
not ( n54405 , n32851 );
nand ( n54406 , n54404 , n54405 );
nor ( n54407 , n54406 , n382079 );
or ( n54408 , n54407 , n32958 );
nand ( n54409 , n54408 , n32845 );
nor ( n54410 , n54181 , n32845 );
and ( n54411 , n54406 , n54410 );
not ( n54412 , n32841 );
nor ( n54413 , n54412 , n44073 );
not ( n54414 , n54413 );
not ( n54415 , n32878 );
and ( n54416 , n54414 , n54415 );
and ( n54417 , n54413 , n32878 );
nor ( n54418 , n54416 , n54417 );
or ( n54419 , n43107 , n54418 );
and ( n54420 , n382523 , RI15b4b9f0_445);
and ( n54421 , n43116 , RI15b457f8_236);
nor ( n54422 , n54420 , n54421 );
nand ( n54423 , n54419 , n54422 );
nor ( n54424 , n54411 , n54423 );
nand ( n54425 , n54409 , n54424 );
buf ( n54426 , n54425 );
buf ( n54427 , n382067 );
buf ( n54428 , n382073 );
buf ( n54429 , n20663 );
not ( n54430 , RI15b47238_292);
not ( n54431 , n385213 );
or ( n54432 , n54430 , n54431 );
and ( n54433 , n385221 , RI15b487c8_338);
and ( n54434 , n20631 , RI15b46ab8_276);
nor ( n54435 , n54433 , n54434 );
nand ( n54436 , n54432 , n54435 );
buf ( n54437 , n54436 );
buf ( n54438 , n380865 );
buf ( n54439 , n43349 );
buf ( n54440 , n22788 );
buf ( n54441 , n379895 );
buf ( n54442 , n381707 );
and ( n54443 , n22544 , n21770 );
not ( n54444 , n384113 );
or ( n54445 , n54444 , n17519 );
nand ( n54446 , n54445 , n21790 );
and ( n54447 , n54446 , RI15b57318_840);
and ( n54448 , n17519 , n22540 );
and ( n54449 , n21795 , n54448 );
nor ( n54450 , n54443 , n54447 , n54449 );
nand ( n54451 , n36470 , n54450 );
buf ( n54452 , n54451 );
nor ( n54453 , n21871 , n45272 );
and ( n54454 , n21802 , n54453 );
and ( n54455 , n381844 , RI15b57b88_858);
not ( n54456 , n21965 );
not ( n54457 , n54456 );
not ( n54458 , n21949 );
or ( n54459 , n54457 , n54458 );
nand ( n54460 , n54459 , n21979 );
and ( n54461 , n54460 , RI15b55d88_794);
nor ( n54462 , n54455 , n54461 );
or ( n54463 , n54462 , n18078 );
and ( n54464 , n18188 , n381842 , n21936 );
or ( n54465 , n22601 , n54456 , RI15b55d88_794);
and ( n54466 , n18177 , RI15b57b88_858);
and ( n54467 , n18219 , RI15b56c88_826);
nor ( n54468 , n54466 , n54467 , n21751 );
nand ( n54469 , n54465 , n54468 );
nor ( n54470 , n54464 , n54469 );
nand ( n54471 , n54463 , n54470 );
nor ( n54472 , n54454 , n54471 );
not ( n54473 , n17507 );
not ( n54474 , n21871 );
or ( n54475 , n54473 , n54474 );
nand ( n54476 , n54475 , n17565 );
nand ( n54477 , n54476 , n45272 );
nand ( n54478 , n54472 , n54477 );
buf ( n54479 , n54478 );
buf ( n54480 , n32676 );
buf ( n54481 , n384218 );
buf ( n54482 , n381081 );
buf ( n54483 , n379802 );
not ( n54484 , n32924 );
not ( n54485 , n32891 );
nand ( n54486 , n54484 , n54485 );
or ( n54487 , n43102 , n54486 );
nor ( n54488 , n54485 , n32884 , n382079 );
nand ( n54489 , n43102 , n54488 );
xor ( n54490 , n44180 , n44181 );
and ( n54491 , n32963 , n54490 );
nand ( n54492 , n54485 , n32884 );
nor ( n54493 , n32928 , n54492 );
or ( n54494 , n46720 , n54485 );
and ( n54495 , n382523 , RI15b4bae0_447);
and ( n54496 , n32052 , RI15b458e8_238);
nor ( n54497 , n54495 , n54496 );
nand ( n54498 , n54494 , n54497 );
nor ( n54499 , n54491 , n54493 , n54498 );
nand ( n54500 , n54487 , n54489 , n54499 );
buf ( n54501 , n54500 );
buf ( n54502 , n19653 );
buf ( n54503 , n382071 );
not ( n54504 , n41979 );
not ( n54505 , n384122 );
or ( n54506 , n54504 , n54505 );
and ( n54507 , n384164 , n39694 );
or ( n54508 , n39703 , n17897 );
or ( n54509 , n33131 , n39707 );
or ( n54510 , n39701 , n384193 );
nand ( n54511 , n54508 , n54509 , n54510 );
nor ( n54512 , n54507 , n54511 );
nand ( n54513 , n54506 , n54512 );
buf ( n54514 , n54513 );
buf ( n54515 , n384199 );
buf ( n54516 , n380942 );
buf ( n54517 , n385112 );
or ( n54518 , n47223 , n41932 );
or ( n54519 , n40142 , n384021 );
not ( n54520 , n38479 );
and ( n54521 , n54520 , RI15b624c0_1219);
not ( n54522 , n54520 );
and ( n54523 , n54522 , n40142 );
nor ( n54524 , n54521 , n54523 );
or ( n54525 , n384024 , n54524 );
nand ( n54526 , n54518 , n54519 , n54525 );
buf ( n54527 , n54526 );
buf ( n54528 , n22402 );
buf ( n54529 , n382052 );
or ( n54530 , n381056 , n19990 );
not ( n54531 , n37169 );
not ( n54532 , n37200 );
and ( n54533 , n54531 , n54532 );
and ( n54534 , n37169 , n37200 );
nor ( n54535 , n54533 , n54534 );
or ( n54536 , n381062 , n54535 );
not ( n54537 , n37126 );
and ( n54538 , n54537 , RI15b49e48_386);
not ( n54539 , n54537 );
and ( n54540 , n54539 , n19990 );
nor ( n54541 , n54538 , n54540 );
or ( n54542 , n54541 , n42690 );
nand ( n54543 , n54530 , n54536 , n54542 );
buf ( n54544 , n54543 );
buf ( n54545 , n22716 );
buf ( n54546 , n32255 );
buf ( n54547 , n31033 );
not ( n54548 , RI15b53a60_719);
not ( n54549 , n32244 );
or ( n54550 , n54548 , n54549 );
and ( n54551 , n32247 , RI15b65058_1312);
and ( n54552 , n32249 , RI15b5fec8_1138);
nor ( n54553 , n54551 , n54552 );
nand ( n54554 , n54550 , n54553 );
buf ( n54555 , n54554 );
buf ( n54556 , n18226 );
not ( n54557 , RI15b557e8_782);
not ( n54558 , n380000 );
or ( n54559 , n54557 , n54558 );
and ( n54560 , n380010 , RI15b4c350_465);
and ( n54561 , n379949 , n385097 );
nor ( n54562 , n54560 , n54561 );
nand ( n54563 , n54559 , n54562 );
buf ( n54564 , n54563 );
or ( n54565 , n383180 , n382936 );
not ( n54566 , n382949 );
and ( n54567 , n54566 , RI15b596b8_916);
or ( n54568 , n383184 , n382933 );
and ( n54569 , n382964 , n41701 );
and ( n54570 , n40019 , n382961 );
nor ( n54571 , n54569 , n54570 );
nand ( n54572 , n54568 , n54571 );
nor ( n54573 , n54567 , n54572 );
nand ( n54574 , n54565 , n54573 );
buf ( n54575 , n54574 );
buf ( n54576 , n383613 );
buf ( n54577 , n22009 );
or ( n54578 , n36937 , n33597 );
and ( n54579 , n36946 , n33600 );
not ( n54580 , RI15b4eb28_550);
or ( n54581 , n33609 , n54580 );
or ( n54582 , n41326 , n33615 );
or ( n54583 , n33607 , n36955 );
nand ( n54584 , n54581 , n54582 , n54583 );
nor ( n54585 , n54579 , n54584 );
nand ( n54586 , n54578 , n54585 );
buf ( n54587 , n54586 );
buf ( n54588 , n31979 );
buf ( n54589 , n379403 );
not ( n54590 , n33581 );
not ( n54591 , n45552 );
or ( n54592 , n54590 , n54591 );
nand ( n54593 , n54592 , n33584 );
nand ( n54594 , n54593 , n33573 );
not ( n54595 , n45552 );
nor ( n54596 , n33573 , n33588 );
and ( n54597 , n54595 , n54596 );
and ( n54598 , n383607 , RI15b5ed70_1101);
and ( n54599 , n383601 , RI15b60378_1148);
nor ( n54600 , n54597 , n54598 , n54599 );
nand ( n54601 , n54594 , n54600 );
buf ( n54602 , n54601 );
buf ( n54603 , n30992 );
buf ( n54604 , n33250 );
not ( n54605 , n33112 );
not ( n54606 , n384726 );
or ( n54607 , n54605 , n54606 );
and ( n54608 , n384737 , n33117 );
or ( n54609 , n33128 , n20792 );
or ( n54610 , n51233 , n33134 );
or ( n54611 , n33126 , n384759 );
nand ( n54612 , n54609 , n54610 , n54611 );
nor ( n54613 , n54608 , n54612 );
nand ( n54614 , n54607 , n54613 );
buf ( n54615 , n54614 );
buf ( n54616 , n380940 );
not ( n54617 , RI15b60648_1154);
nor ( n54618 , n54617 , n383600 );
buf ( n54619 , n54618 );
buf ( n54620 , n384203 );
buf ( n54621 , n22479 );
buf ( n54622 , RI15b47580_299);
buf ( n54623 , n20663 );
not ( n54624 , n34796 );
and ( n54625 , n54624 , RI15b4aa00_411);
and ( n54626 , n19830 , n22217 );
not ( n54627 , n34797 );
and ( n54628 , n34793 , n54627 );
nor ( n54629 , n54625 , n54626 , n54628 );
nand ( n54630 , n41499 , n54629 );
buf ( n54631 , n54630 );
buf ( n54632 , n381490 );
buf ( n54633 , n31030 );
or ( n54634 , n53750 , n379708 );
not ( n54635 , n386987 );
or ( n54636 , n54635 , n387004 );
nand ( n54637 , n54636 , n383408 );
nand ( n54638 , n54637 , RI15b626a0_1223);
and ( n54639 , n54635 , n47516 , n386988 );
or ( n54640 , n49459 , n53734 , RI15b644a0_1287);
or ( n54641 , n19598 , n386781 );
nand ( n54642 , n54640 , n54641 );
nor ( n54643 , n54639 , n54642 );
not ( n54644 , n386785 );
not ( n54645 , n386906 );
nand ( n54646 , n54644 , n54645 , n34844 );
and ( n54647 , n54638 , n54643 , n54646 );
or ( n54648 , n54645 , n22473 );
nand ( n54649 , n54648 , n53232 );
nand ( n54650 , n54649 , n386785 );
nand ( n54651 , n54634 , n54647 , n54650 );
buf ( n54652 , n54651 );
not ( n54653 , n385218 );
nand ( n54654 , n382509 , RI15b48318_328);
nand ( n54655 , n54653 , n54654 );
and ( n54656 , n54655 , RI15b3fab0_37);
and ( n54657 , n43961 , n40007 );
nor ( n54658 , n54657 , n19913 );
nor ( n54659 , n54656 , n54658 , n43964 );
not ( n54660 , n54659 );
buf ( n54661 , n54660 );
buf ( n54662 , n22406 );
buf ( n54663 , n31719 );
buf ( n54664 , n385197 );
buf ( n54665 , n385195 );
buf ( n54666 , n22740 );
buf ( n54667 , n32255 );
not ( n54668 , RI15b46770_269);
not ( n54669 , n379832 );
or ( n54670 , n54668 , n54669 );
and ( n54671 , n379825 , RI15b48480_331);
nor ( n54672 , n54671 , n35583 );
nand ( n54673 , n54670 , n54672 );
buf ( n54674 , n54673 );
buf ( n54675 , n379802 );
buf ( n54676 , n35649 );
buf ( n54677 , n32676 );
not ( n54678 , RI15b4a3e8_398);
not ( n54679 , n30908 );
or ( n54680 , n54678 , n54679 );
or ( n54681 , n22216 , n19727 );
not ( n54682 , RI15b4a3e8_398);
and ( n54683 , n54682 , RI15b4a370_397);
and ( n54684 , n32195 , RI15b4a3e8_398);
nor ( n54685 , n54683 , n54684 );
or ( n54686 , n54685 , n20638 );
not ( n54687 , n40183 );
and ( n54688 , n386333 , n54687 );
not ( n54689 , n386333 );
and ( n54690 , n32203 , n40182 );
not ( n54691 , n386307 );
nor ( n54692 , n54690 , n54691 );
and ( n54693 , n54689 , n54692 );
nor ( n54694 , n54688 , n54693 );
not ( n54695 , n35191 );
and ( n54696 , n54694 , n54695 );
not ( n54697 , n54694 );
and ( n54698 , n54697 , n35191 );
nor ( n54699 , n54696 , n54698 );
and ( n54700 , n386500 , n54699 );
not ( n54701 , n385753 );
not ( n54702 , n54701 );
not ( n54703 , n385558 );
not ( n54704 , n35189 );
not ( n54705 , n54704 );
or ( n54706 , n54703 , n54705 );
or ( n54707 , n35190 , n385558 );
nand ( n54708 , n54706 , n54707 );
not ( n54709 , n54708 );
and ( n54710 , n54702 , n54709 );
and ( n54711 , n54701 , n54708 );
nor ( n54712 , n54710 , n54711 );
or ( n54713 , n386013 , n54712 );
xor ( n54714 , n386094 , n385591 );
xor ( n54715 , n54714 , n386117 );
and ( n54716 , n386258 , n54715 );
and ( n54717 , n22393 , RI15b4b2e8_430);
nor ( n54718 , n54716 , n54717 );
nand ( n54719 , n54713 , n54718 );
nor ( n54720 , n54700 , n54719 );
nand ( n54721 , n54681 , n54686 , n54720 );
not ( n54722 , n54721 );
nand ( n54723 , n54680 , n54722 );
buf ( n54724 , n54723 );
buf ( n54725 , n386563 );
buf ( n54726 , n32672 );
buf ( n54727 , n22402 );
not ( n54728 , RI15b534c0_707);
not ( n54729 , n32244 );
or ( n54730 , n54728 , n54729 );
and ( n54731 , n32247 , RI15b64ab8_1300);
and ( n54732 , n32249 , RI15b5f928_1126);
nor ( n54733 , n54731 , n54732 );
nand ( n54734 , n54730 , n54733 );
buf ( n54735 , n54734 );
and ( n54736 , n385164 , RI15b50b08_618);
not ( n54737 , n36473 );
or ( n54738 , n54737 , n381816 );
or ( n54739 , n381784 , n385170 );
or ( n54740 , n381726 , n385178 );
nand ( n54741 , n54738 , n54739 , n54740 );
nor ( n54742 , n54736 , n54741 );
nand ( n54743 , n381825 , n54742 );
buf ( n54744 , n54743 );
buf ( n54745 , n18226 );
buf ( n54746 , n379802 );
and ( n54747 , n36490 , n33995 );
nand ( n54748 , n54747 , n379785 );
not ( n54749 , n54748 );
not ( n54750 , n46287 );
or ( n54751 , n54749 , n54750 );
not ( n54752 , n33984 );
nand ( n54753 , n54751 , n54752 );
nor ( n54754 , n54747 , n54752 );
nand ( n54755 , n40809 , n54754 );
buf ( n54756 , n34568 );
not ( n54757 , n54756 );
not ( n54758 , n34588 );
and ( n54759 , n54757 , n54758 );
not ( n54760 , n54757 );
and ( n54761 , n54760 , n34588 );
nor ( n54762 , n54759 , n54761 );
and ( n54763 , n54762 , n36513 );
not ( n54764 , RI15b5e398_1080);
not ( n54765 , n34651 );
or ( n54766 , n54764 , n54765 );
or ( n54767 , n36518 , n379445 );
nand ( n54768 , n54766 , n54767 );
nor ( n54769 , n54763 , n54768 );
nand ( n54770 , n54753 , n54755 , n54769 );
buf ( n54771 , n54770 );
buf ( n54772 , n31719 );
buf ( n54773 , n386760 );
not ( n54774 , n37114 );
nor ( n54775 , n54774 , RI15b4a190_393);
nor ( n54776 , n37138 , n54775 );
or ( n54777 , n54776 , n20528 );
nor ( n54778 , n37140 , n37107 , RI15b4a208_394);
nand ( n54779 , n37426 , n54778 );
nand ( n54780 , n54777 , n54779 );
buf ( n54781 , n54780 );
buf ( n54782 , n22716 );
buf ( n54783 , n20663 );
not ( n54784 , RI15b536a0_711);
not ( n54785 , n32244 );
or ( n54786 , n54784 , n54785 );
and ( n54787 , n32247 , RI15b64c98_1304);
and ( n54788 , n32249 , RI15b5fb08_1130);
nor ( n54789 , n54787 , n54788 );
nand ( n54790 , n54786 , n54789 );
buf ( n54791 , n54790 );
buf ( n54792 , n382071 );
or ( n54793 , n31006 , n384704 );
and ( n54794 , n31016 , n384739 );
or ( n54795 , n384749 , n17729 );
or ( n54796 , n40593 , n384757 );
or ( n54797 , n384747 , n31024 );
nand ( n54798 , n54795 , n54796 , n54797 );
nor ( n54799 , n54794 , n54798 );
nand ( n54800 , n54793 , n54799 );
buf ( n54801 , n54800 );
buf ( n54802 , n384996 );
nand ( n54803 , n384914 , n384897 );
nand ( n54804 , n384918 , RI15b5f568_1118);
and ( n54805 , n384922 , n44092 );
nor ( n54806 , n54805 , n32342 );
not ( n54807 , n54806 );
not ( n54808 , n383565 );
and ( n54809 , n54807 , n54808 );
and ( n54810 , n384934 , n44098 );
nor ( n54811 , n54809 , n54810 );
nand ( n54812 , n51523 , n54803 , n54804 , n54811 );
buf ( n54813 , n54812 );
buf ( n54814 , n386563 );
or ( n54815 , n52829 , n34967 );
not ( n54816 , n52827 );
and ( n54817 , n54816 , n48968 , n34967 );
or ( n54818 , n49099 , n54535 );
or ( n54819 , n386547 , n22059 );
nand ( n54820 , n54818 , n54819 );
nor ( n54821 , n54817 , n54820 );
nand ( n54822 , n54815 , n54821 , n41021 );
buf ( n54823 , n54822 );
buf ( n54824 , n386762 );
buf ( n54825 , n31033 );
buf ( n54826 , n22738 );
buf ( n54827 , n22402 );
or ( n54828 , n44431 , n22035 );
nand ( n54829 , n35525 , RI15b53a60_719);
nand ( n54830 , n54828 , n54829 );
buf ( n54831 , n54830 );
buf ( n54832 , n35651 );
not ( n54833 , RI15b53790_713);
not ( n54834 , n383170 );
or ( n54835 , n54833 , n54834 );
not ( n54836 , n33455 );
not ( n54837 , n33453 );
or ( n54838 , n54836 , n54837 );
nand ( n54839 , n54838 , n33465 );
not ( n54840 , n33462 );
and ( n54841 , n54839 , n54840 );
nor ( n54842 , n33455 , n54840 );
and ( n54843 , n33476 , n54842 );
and ( n54844 , n383147 , RI15b53010_697);
nor ( n54845 , n54841 , n54843 , n54844 );
nand ( n54846 , n54835 , n54845 );
buf ( n54847 , n54846 );
not ( n54848 , n33387 );
not ( n54849 , n381589 );
or ( n54850 , n54848 , n54849 );
and ( n54851 , n381596 , n33417 );
not ( n54852 , RI15b5b710_985);
or ( n54853 , n33428 , n54852 );
or ( n54854 , n42258 , n33440 );
or ( n54855 , n33426 , n381621 );
nand ( n54856 , n54853 , n54854 , n54855 );
nor ( n54857 , n54851 , n54856 );
nand ( n54858 , n54850 , n54857 );
buf ( n54859 , n54858 );
buf ( n54860 , n382537 );
buf ( n54861 , n20665 );
buf ( n54862 , n386760 );
or ( n54863 , n37478 , n35957 );
and ( n54864 , n384983 , n36986 );
or ( n54865 , n35967 , n20409 );
or ( n54866 , n22022 , n35973 );
or ( n54867 , n35965 , n384988 );
nand ( n54868 , n54865 , n54866 , n54867 );
nor ( n54869 , n54864 , n54868 );
nand ( n54870 , n54863 , n54869 );
buf ( n54871 , n54870 );
not ( n54872 , n35930 );
not ( n54873 , n54872 );
not ( n54874 , n32129 );
or ( n54875 , n54873 , n54874 );
and ( n54876 , n36974 , RI15b40e60_79);
or ( n54877 , n32141 , n35934 );
or ( n54878 , n32148 , n35950 );
or ( n54879 , n35944 , n32150 );
nand ( n54880 , n54877 , n54878 , n54879 );
nor ( n54881 , n54876 , n54880 );
nand ( n54882 , n54875 , n54881 );
buf ( n54883 , n54882 );
buf ( n54884 , n383498 );
buf ( n54885 , n32981 );
buf ( n54886 , n381490 );
and ( n54887 , n49030 , n50343 );
or ( n54888 , n386541 , n50326 );
or ( n54889 , n50315 , n386550 );
or ( n54890 , n386557 , n50332 );
nand ( n54891 , n54888 , n54889 , n54890 );
nor ( n54892 , n54887 , n54891 );
nand ( n54893 , n50354 , n54892 );
buf ( n54894 , n54893 );
buf ( n54895 , n22655 );
buf ( n54896 , n31719 );
buf ( n54897 , n35651 );
buf ( n54898 , n384199 );
or ( n54899 , n386705 , n384057 );
and ( n54900 , n386716 , n384169 );
or ( n54901 , n384182 , n17862 );
or ( n54902 , n37443 , n384190 );
or ( n54903 , n384180 , n386738 );
nand ( n54904 , n54901 , n54902 , n54903 );
nor ( n54905 , n54900 , n54904 );
nand ( n54906 , n54899 , n54905 );
buf ( n54907 , n54906 );
and ( n54908 , n22646 , RI15b45078_220);
and ( n54909 , n22648 , RI15b514e0_639);
nor ( n54910 , n54908 , n54909 );
not ( n54911 , n54910 );
buf ( n54912 , n54911 );
buf ( n54913 , n383345 );
and ( n54914 , n46239 , n383930 );
and ( n54915 , n45927 , RI15b621f0_1213);
or ( n54916 , n45923 , n386970 , RI15b621f0_1213);
or ( n54917 , n386972 , RI15b62178_1212);
nand ( n54918 , n54916 , n54917 );
and ( n54919 , n384025 , n54918 );
nor ( n54920 , n54914 , n54915 , n54919 );
not ( n54921 , n54920 );
buf ( n54922 , n54921 );
buf ( n54923 , n31033 );
or ( n54924 , n40166 , n386325 );
not ( n54925 , n42859 );
and ( n54926 , n386540 , RI15b43db8_180);
and ( n54927 , n386549 , n385432 );
and ( n54928 , n386556 , n386131 );
nor ( n54929 , n54926 , n54927 , n54928 );
nand ( n54930 , n54924 , n54925 , n54929 );
buf ( n54931 , n54930 );
buf ( n54932 , n22655 );
buf ( n54933 , n385197 );
buf ( n54934 , n22007 );
buf ( n54935 , n32160 );
or ( n54936 , n383814 , n39691 );
and ( n54937 , n383857 , n39694 );
or ( n54938 , n39703 , n21111 );
or ( n54939 , n41099 , n39707 );
or ( n54940 , n39701 , n383917 );
nand ( n54941 , n54938 , n54939 , n54940 );
nor ( n54942 , n54937 , n54941 );
nand ( n54943 , n54936 , n54942 );
buf ( n54944 , n54943 );
buf ( n54945 , n22653 );
buf ( n54946 , n19655 );
buf ( n54947 , n379847 );
or ( n54948 , n386990 , n384021 );
or ( n54949 , n386747 , n41436 );
and ( n54950 , n38484 , RI15b62718_1224);
not ( n54951 , n38484 );
and ( n54952 , n54951 , n386990 );
nor ( n54953 , n54950 , n54952 );
or ( n54954 , n384024 , n54953 );
nand ( n54955 , n54948 , n54949 , n54954 );
buf ( n54956 , n54955 );
buf ( n54957 , n382052 );
or ( n54958 , n386705 , n35472 );
and ( n54959 , n386716 , n35479 );
not ( n54960 , RI15b4df70_525);
or ( n54961 , n35488 , n54960 );
or ( n54962 , n45435 , n35497 );
or ( n54963 , n35486 , n386738 );
nand ( n54964 , n54961 , n54962 , n54963 );
nor ( n54965 , n54959 , n54964 );
nand ( n54966 , n54958 , n54965 );
buf ( n54967 , n54966 );
buf ( n54968 , n22714 );
buf ( n54969 , n22343 );
or ( n54970 , n31053 , n36293 );
nand ( n54971 , n384907 , n384860 );
and ( n54972 , n41338 , RI15b60f30_1173);
and ( n54973 , n36538 , n36869 );
not ( n54974 , RI15b60eb8_1172);
or ( n54975 , n41341 , n54974 , RI15b60f30_1173);
not ( n54976 , RI15b60f30_1173);
or ( n54977 , n54976 , RI15b60eb8_1172);
nand ( n54978 , n54975 , n54977 );
and ( n54979 , n36541 , n54978 );
nor ( n54980 , n54972 , n54973 , n54979 );
nand ( n54981 , n54970 , n54971 , n54980 );
buf ( n54982 , n54981 );
buf ( n54983 , n19651 );
buf ( n54984 , n381006 );
not ( n54985 , n36200 );
not ( n54986 , n54985 );
not ( n54987 , n33174 );
or ( n54988 , n54986 , n54987 );
and ( n54989 , n33196 , n36202 );
or ( n54990 , n36212 , n385311 );
or ( n54991 , n22241 , n36217 );
or ( n54992 , n36210 , n33201 );
nand ( n54993 , n54990 , n54991 , n54992 );
nor ( n54994 , n54989 , n54993 );
nand ( n54995 , n54988 , n54994 );
buf ( n54996 , n54995 );
buf ( n54997 , RI15b5d9c0_1059);
buf ( n54998 , n382069 );
buf ( n54999 , n22788 );
buf ( n55000 , n22714 );
buf ( n55001 , n21800 );
buf ( n55002 , n31033 );
or ( n55003 , n35333 , n34979 );
and ( n55004 , n35373 , RI15b433e0_159);
and ( n55005 , n35376 , RI15b437a0_167);
and ( n55006 , n35537 , RI15b43020_151);
and ( n55007 , n35384 , RI15b42c60_143);
nor ( n55008 , n55006 , n55007 );
and ( n55009 , n35541 , RI15b41220_87);
and ( n55010 , n35543 , RI15b40e60_79);
nor ( n55011 , n55009 , n55010 );
and ( n55012 , n35546 , RI15b419a0_103);
and ( n55013 , n35548 , RI15b415e0_95);
nor ( n55014 , n55012 , n55013 );
and ( n55015 , n35391 , RI15b42120_119);
and ( n55016 , n35396 , RI15b424e0_127);
and ( n55017 , n35401 , RI15b3ff60_47);
and ( n55018 , n35407 , RI15b40320_55);
nor ( n55019 , n55016 , n55017 , n55018 );
and ( n55020 , n35410 , RI15b40aa0_71);
and ( n55021 , n35412 , RI15b41d60_111);
nor ( n55022 , n55020 , n55021 );
and ( n55023 , n35415 , RI15b428a0_135);
and ( n55024 , n383378 , RI15b406e0_63);
nor ( n55025 , n55023 , n55024 );
and ( n55026 , n55019 , n55022 , n55025 );
nor ( n55027 , n55026 , n381047 );
nor ( n55028 , n55015 , n55027 );
and ( n55029 , n55011 , n55014 , n55028 );
nand ( n55030 , n55008 , n55029 );
nor ( n55031 , n55004 , n55005 , n55030 );
not ( n55032 , n55031 );
and ( n55033 , n55032 , n41715 );
and ( n55034 , n35335 , RI15b66048_1346);
and ( n55035 , n35355 , n34979 );
not ( n55036 , n35355 );
and ( n55037 , n55036 , RI15b48c78_348);
nor ( n55038 , n55035 , n55037 );
and ( n55039 , n55038 , n35580 );
nor ( n55040 , n55033 , n55034 , n55039 );
nand ( n55041 , n55003 , n55040 , n51209 );
buf ( n55042 , n55041 );
buf ( n55043 , n381490 );
buf ( n55044 , n381021 );
or ( n55045 , n381017 , n22044 );
nand ( n55046 , n35525 , RI15b53d30_725);
nand ( n55047 , n55045 , n55046 );
buf ( n55048 , n55047 );
buf ( n55049 , n19856 );
not ( n55050 , n35293 );
and ( n55051 , n55049 , n55050 );
nor ( n55052 , n55051 , n38940 );
or ( n55053 , n55052 , n19860 );
or ( n55054 , n382122 , n32526 );
not ( n55055 , n19860 );
nor ( n55056 , n55055 , n380868 );
not ( n55057 , n55049 );
and ( n55058 , n55056 , n55057 );
not ( n55059 , n31806 );
not ( n55060 , n19986 );
not ( n55061 , n55060 );
or ( n55062 , n55059 , n55061 );
nand ( n55063 , n55062 , n380875 );
and ( n55064 , n55063 , RI15b49d58_384);
or ( n55065 , n55060 , n20529 , RI15b49d58_384);
or ( n55066 , n20553 , n382120 , RI15b4bb58_448);
or ( n55067 , n382122 , RI15b4bae0_447);
nand ( n55068 , n55066 , n55067 );
and ( n55069 , n20566 , n55068 );
and ( n55070 , n22388 , RI15b4bb58_448);
and ( n55071 , n42325 , RI15b4ac58_416);
nor ( n55072 , n55069 , n55070 , n55071 );
nand ( n55073 , n55065 , n55072 );
nor ( n55074 , n55058 , n55064 , n55073 );
nand ( n55075 , n55053 , n55054 , n55074 );
buf ( n55076 , n55075 );
buf ( n55077 , n382537 );
buf ( n55078 , n22740 );
buf ( n55079 , n381490 );
buf ( n55080 , n22005 );
or ( n55081 , n380716 , n383437 );
nand ( n55082 , n55081 , n32582 );
and ( n55083 , n55082 , RI15b63348_1250);
not ( n55084 , n383437 );
or ( n55085 , n384652 , n55084 , RI15b63348_1250);
or ( n55086 , n386878 , n22775 );
nand ( n55087 , n55085 , n55086 );
nor ( n55088 , n55083 , n55087 );
nand ( n55089 , n54392 , n55088 );
buf ( n55090 , n55089 );
buf ( n55091 , n22738 );
and ( n55092 , n30908 , RI15b4a730_405);
and ( n55093 , n38994 , n22217 );
not ( n55094 , n19782 );
and ( n55095 , n55094 , n19786 );
not ( n55096 , n55094 );
and ( n55097 , n55096 , RI15b4a730_405);
nor ( n55098 , n55095 , n55097 );
and ( n55099 , n55098 , n20637 );
nor ( n55100 , n55092 , n55093 , n55099 );
nand ( n55101 , n44691 , n55100 );
buf ( n55102 , n55101 );
buf ( n55103 , n32981 );
buf ( n55104 , n21800 );
buf ( n55105 , n384199 );
not ( n55106 , n386923 );
nor ( n55107 , n55106 , n22473 );
or ( n55108 , n55107 , n386945 );
nand ( n55109 , n55108 , n386930 );
not ( n55110 , n383408 );
buf ( n55111 , n386997 );
not ( n55112 , n387004 );
nand ( n55113 , n55111 , n55112 );
not ( n55114 , n55113 );
or ( n55115 , n55110 , n55114 );
nand ( n55116 , n55115 , RI15b62970_1229);
not ( n55117 , n34844 );
nor ( n55118 , n55117 , n386930 );
nand ( n55119 , n55106 , n55118 );
not ( n55120 , n55111 );
nor ( n55121 , n383482 , RI15b62970_1229);
and ( n55122 , n55120 , n55121 );
nand ( n55123 , n30850 , n22450 );
nand ( n55124 , n55123 , n22425 );
nand ( n55125 , n55124 , RI15b64770_1293);
and ( n55126 , n30851 , n22450 , n33958 );
and ( n55127 , n19599 , RI15b63870_1261);
nor ( n55128 , n55126 , n55127 );
nand ( n55129 , n55125 , n55128 );
nor ( n55130 , n55122 , n55129 );
nand ( n55131 , n55109 , n55116 , n55119 , n55130 );
buf ( n55132 , n55131 );
or ( n55133 , n383814 , n384704 );
and ( n55134 , n383857 , n384739 );
or ( n55135 , n384749 , n21155 );
or ( n55136 , n41182 , n384757 );
or ( n55137 , n384747 , n383917 );
nand ( n55138 , n55135 , n55136 , n55137 );
nor ( n55139 , n55134 , n55138 );
nand ( n55140 , n55133 , n55139 );
buf ( n55141 , n55140 );
buf ( n55142 , n379895 );
buf ( n55143 , n22343 );
nand ( n55144 , n44037 , n40602 );
nand ( n55145 , n384918 , RI15b5f658_1120);
and ( n55146 , n384922 , n383575 );
nor ( n55147 , n55146 , n32342 );
not ( n55148 , n55147 );
not ( n55149 , n383586 );
and ( n55150 , n55148 , n55149 );
and ( n55151 , n384934 , n383605 );
nor ( n55152 , n55150 , n55151 );
nand ( n55153 , n40606 , n55144 , n55145 , n55152 );
buf ( n55154 , n55153 );
buf ( n55155 , n35651 );
buf ( n55156 , n380865 );
and ( n55157 , n379822 , RI15b65aa8_1334);
and ( n55158 , n379825 , RI15b486d8_336);
nor ( n55159 , n55157 , n55158 );
nand ( n55160 , n379832 , RI15b469c8_274);
nand ( n55161 , n55159 , n55160 , n35591 );
buf ( n55162 , n55161 );
buf ( n55163 , n22402 );
buf ( n55164 , n383345 );
buf ( n55165 , n32271 );
buf ( n55166 , n384203 );
or ( n55167 , n32430 , n54118 );
and ( n55168 , n386637 , RI15b54d98_760);
and ( n55169 , n38346 , n386671 );
not ( n55170 , RI15b54d98_760);
not ( n55171 , n382644 );
not ( n55172 , n55171 );
or ( n55173 , n55170 , n55172 );
or ( n55174 , n55171 , RI15b54d98_760);
nand ( n55175 , n55173 , n55174 );
and ( n55176 , n37449 , n55175 );
nor ( n55177 , n55168 , n55169 , n55176 );
and ( n55178 , n54120 , n55177 );
nand ( n55179 , n55167 , n55178 );
buf ( n55180 , n55179 );
not ( n55181 , n386590 );
not ( n55182 , n381507 );
or ( n55183 , n55181 , n55182 );
and ( n55184 , n381524 , n386603 );
not ( n55185 , RI15b5a108_938);
or ( n55186 , n386612 , n55185 );
or ( n55187 , n47660 , n386624 );
or ( n55188 , n386610 , n381560 );
nand ( n55189 , n55186 , n55187 , n55188 );
nor ( n55190 , n55184 , n55189 );
nand ( n55191 , n55183 , n55190 );
buf ( n55192 , n55191 );
buf ( n55193 , n384996 );
buf ( n55194 , n386762 );
buf ( n55195 , n379895 );
buf ( n55196 , RI15b46f68_286);
or ( n55197 , n47344 , n380001 );
or ( n55198 , n51400 , n45835 );
not ( n55199 , n379979 );
and ( n55200 , n55199 , RI15b56328_806);
not ( n55201 , n55199 );
and ( n55202 , n55201 , n47344 );
nor ( n55203 , n55200 , n55202 );
or ( n55204 , n379948 , n55203 );
nand ( n55205 , n55197 , n55198 , n55204 );
buf ( n55206 , n55205 );
or ( n55207 , n383180 , n47643 );
not ( n55208 , n47658 );
and ( n55209 , n55208 , RI15b58b78_892);
or ( n55210 , n383184 , n47648 );
or ( n55211 , n383189 , n47663 );
or ( n55212 , n47656 , n383192 );
nand ( n55213 , n55210 , n55211 , n55212 );
nor ( n55214 , n55209 , n55213 );
and ( n55215 , n55207 , n55214 );
buf ( n55216 , n55215 );
buf ( n55217 , n385112 );
buf ( n55218 , n22738 );
and ( n55219 , n385164 , RI15b50928_614);
not ( n55220 , n21735 );
or ( n55221 , n36694 , n55220 );
or ( n55222 , n21329 , n385170 );
or ( n55223 , n21542 , n385178 );
nand ( n55224 , n55221 , n55222 , n55223 );
nor ( n55225 , n55219 , n55224 );
nand ( n55226 , n21755 , n55225 );
buf ( n55227 , n55226 );
buf ( n55228 , n22005 );
buf ( n55229 , n382069 );
not ( n55230 , n47923 );
not ( n55231 , n34645 );
nand ( n55232 , n55230 , n55231 );
nor ( n55233 , n47903 , n55232 );
buf ( n55234 , n44377 );
nand ( n55235 , n55234 , n379785 );
not ( n55236 , n55235 );
not ( n55237 , n36494 );
or ( n55238 , n55236 , n55237 );
buf ( n55239 , n44378 );
not ( n55240 , n55239 );
nand ( n55241 , n55238 , n55240 );
not ( n55242 , n55241 );
nor ( n55243 , n55233 , n55242 );
not ( n55244 , n51690 );
not ( n55245 , n47903 );
or ( n55246 , n55244 , n55245 );
not ( n55247 , n55239 );
nor ( n55248 , n55234 , n55247 );
not ( n55249 , n55248 );
not ( n55250 , n34249 );
or ( n55251 , n55249 , n55250 );
and ( n55252 , n379783 , RI15b64770_1293);
and ( n55253 , n34651 , RI15b5e578_1084);
nor ( n55254 , n55252 , n55253 );
nand ( n55255 , n55251 , n55254 );
not ( n55256 , n55255 );
nand ( n55257 , n55246 , n55256 );
not ( n55258 , n55257 );
nand ( n55259 , n55243 , n55258 );
not ( n55260 , n55259 );
not ( n55261 , n35651 );
not ( n55262 , n35651 );
not ( n55263 , n21276 );
not ( n55264 , n45249 );
or ( n55265 , n55263 , n55264 );
or ( n55266 , n45249 , n21276 );
nand ( n55267 , n55265 , n55266 );
and ( n55268 , n55267 , n21357 );
not ( n55269 , n45259 );
not ( n55270 , n55269 );
not ( n55271 , n45260 );
and ( n55272 , n55270 , n55271 );
and ( n55273 , n55269 , n45260 );
nor ( n55274 , n55272 , n55273 );
or ( n55275 , n55274 , n21561 );
or ( n55276 , n21750 , n21934 );
nand ( n55277 , n55275 , n55276 );
nor ( n55278 , n55268 , n55277 );
not ( n55279 , n21679 );
not ( n55280 , n44730 );
not ( n55281 , n55280 );
or ( n55282 , n55279 , n55281 );
nand ( n55283 , n55282 , n45241 );
nand ( n55284 , n55283 , n21746 );
nand ( n55285 , n55278 , n55284 );
not ( n55286 , n55285 );
and ( n55287 , n21788 , RI15b56c10_825);
and ( n55288 , n21870 , n21768 );
buf ( n55289 , n21864 );
and ( n55290 , n55289 , n17536 );
not ( n55291 , n55289 );
and ( n55292 , n55291 , RI15b56c10_825);
nor ( n55293 , n55290 , n55292 );
and ( n55294 , n55293 , n384113 );
nor ( n55295 , n55287 , n55288 , n55294 );
nand ( n55296 , n55286 , n55295 );
buf ( n55297 , n55296 );
not ( n55298 , n22545 );
nor ( n55299 , n55298 , n17506 );
or ( n55300 , n55299 , n379905 );
nand ( n55301 , n55300 , n50985 );
buf ( n55302 , n22593 );
nor ( n55303 , n55302 , n18079 );
or ( n55304 , n55303 , n18103 );
nand ( n55305 , n55304 , RI15b56490_809);
nor ( n55306 , n18197 , RI15b56490_809);
and ( n55307 , n55302 , n55306 );
or ( n55308 , n45231 , n379309 );
not ( n55309 , n22620 );
or ( n55310 , n55309 , n22839 , RI15b58290_873);
or ( n55311 , n379309 , RI15b58218_872);
nand ( n55312 , n55310 , n55311 );
and ( n55313 , n55312 , n18188 );
and ( n55314 , n18219 , RI15b57390_841);
nor ( n55315 , n55313 , n55314 );
nand ( n55316 , n55308 , n55315 );
nor ( n55317 , n55307 , n55316 );
nor ( n55318 , n17577 , n50985 );
nand ( n55319 , n55298 , n55318 );
nand ( n55320 , n55301 , n55305 , n55317 , n55319 );
buf ( n55321 , n55320 );
buf ( n55322 , n22479 );
buf ( n55323 , n22406 );
buf ( n55324 , n382069 );
buf ( n55325 , n383345 );
or ( n55326 , n35852 , n35957 );
and ( n55327 , n35968 , RI15b3fee8_46);
or ( n55328 , n35582 , n35973 );
or ( n55329 , n35856 , n35965 );
or ( n55330 , n35959 , n35858 );
nand ( n55331 , n55328 , n55329 , n55330 );
nor ( n55332 , n55327 , n55331 );
nand ( n55333 , n55326 , n55332 );
buf ( n55334 , n55333 );
not ( n55335 , n54872 );
not ( n55336 , n39319 );
or ( n55337 , n55335 , n55336 );
and ( n55338 , n33196 , n35935 );
not ( n55339 , RI15b41130_85);
or ( n55340 , n35946 , n55339 );
or ( n55341 , n22241 , n35950 );
or ( n55342 , n35944 , n33201 );
nand ( n55343 , n55340 , n55341 , n55342 );
nor ( n55344 , n55338 , n55343 );
nand ( n55345 , n55337 , n55344 );
buf ( n55346 , n55345 );
buf ( n55347 , n22007 );
buf ( n55348 , n382067 );
buf ( n55349 , n380903 );
buf ( n55350 , n31591 );
not ( n55351 , n55350 );
buf ( n55352 , n31583 );
not ( n55353 , n55352 );
and ( n55354 , n55351 , n55353 );
not ( n55355 , n55351 );
and ( n55356 , n55355 , n55352 );
nor ( n55357 , n55354 , n55356 );
or ( n55358 , n55357 , n52463 );
buf ( n55359 , n31659 );
not ( n55360 , n55359 );
or ( n55361 , n55360 , n31667 );
nand ( n55362 , n55361 , n31700 );
and ( n55363 , n55362 , n31663 );
or ( n55364 , n55359 , n40972 , n31663 );
and ( n55365 , n379394 , RI15b58128_870);
and ( n55366 , n47038 , RI15b51f30_661);
nor ( n55367 , n55365 , n55366 );
nand ( n55368 , n55364 , n55367 );
nor ( n55369 , n55363 , n55368 );
nand ( n55370 , n55358 , n55369 );
buf ( n55371 , n55370 );
and ( n55372 , n31792 , n384612 );
not ( n55373 , RI15b5cf70_1037);
not ( n55374 , n31770 );
or ( n55375 , n55373 , n55374 );
and ( n55376 , n49122 , n384250 );
and ( n55377 , n384489 , n31778 );
nor ( n55378 , n55376 , n55377 );
nand ( n55379 , n55375 , n55378 );
nor ( n55380 , n55372 , n55379 );
nand ( n55381 , n384621 , n55380 );
buf ( n55382 , n55381 );
buf ( n55383 , n32672 );
buf ( n55384 , n384199 );
or ( n55385 , n383814 , n31151 );
and ( n55386 , n383857 , n31164 );
or ( n55387 , n31175 , n21151 );
or ( n55388 , n41458 , n31182 );
or ( n55389 , n31173 , n383917 );
nand ( n55390 , n55387 , n55388 , n55389 );
nor ( n55391 , n55386 , n55390 );
nand ( n55392 , n55385 , n55391 );
buf ( n55393 , n55392 );
buf ( n55394 , n22009 );
and ( n55395 , n36536 , RI15b61458_1184);
not ( n55396 , n384903 );
and ( n55397 , n55396 , n384774 );
nor ( n55398 , n55397 , n384912 );
not ( n55399 , n41080 );
or ( n55400 , n55399 , n31122 );
not ( n55401 , n384772 );
or ( n55402 , n55401 , n31052 );
not ( n55403 , n41413 );
not ( n55404 , RI15b61458_1184);
and ( n55405 , n55403 , n55404 );
and ( n55406 , n41413 , RI15b61458_1184);
nor ( n55407 , n55405 , n55406 );
or ( n55408 , n55407 , n41336 );
nand ( n55409 , n55400 , n55402 , n55408 );
nor ( n55410 , n55395 , n55398 , n55409 );
not ( n55411 , n55410 );
buf ( n55412 , n55411 );
buf ( n55413 , n22408 );
buf ( n55414 , n22343 );
or ( n55415 , n381907 , n37495 );
and ( n55416 , n44521 , RI15b42558_128);
or ( n55417 , n381917 , n37497 );
not ( n55418 , n37512 );
and ( n55419 , n55418 , n381923 );
and ( n55420 , n381926 , n37510 );
nor ( n55421 , n55419 , n55420 );
nand ( n55422 , n55417 , n55421 );
nor ( n55423 , n55416 , n55422 );
nand ( n55424 , n55415 , n55423 );
buf ( n55425 , n55424 );
buf ( n55426 , n379802 );
buf ( n55427 , n22788 );
buf ( n55428 , n22402 );
not ( n55429 , n54985 );
not ( n55430 , n32129 );
or ( n55431 , n55429 , n55430 );
and ( n55432 , n42409 , RI15b415e0_95);
or ( n55433 , n32141 , n36204 );
or ( n55434 , n32148 , n36217 );
or ( n55435 , n36210 , n32150 );
nand ( n55436 , n55433 , n55434 , n55435 );
nor ( n55437 , n55432 , n55436 );
nand ( n55438 , n55431 , n55437 );
buf ( n55439 , n55438 );
buf ( n55440 , n381006 );
buf ( n55441 , n384218 );
and ( n55442 , n22646 , RI15b453c0_227);
and ( n55443 , n22648 , RI15b51828_646);
nor ( n55444 , n55442 , n55443 );
not ( n55445 , n55444 );
buf ( n55446 , n55445 );
buf ( n55447 , n22007 );
buf ( n55448 , n22714 );
buf ( n55449 , n384203 );
not ( n55450 , RI15b534c0_707);
not ( n55451 , n383170 );
or ( n55452 , n55450 , n55451 );
and ( n55453 , n33453 , RI15b54a50_753);
and ( n55454 , n383147 , RI15b52d40_691);
nor ( n55455 , n55453 , n55454 );
nand ( n55456 , n55452 , n55455 );
buf ( n55457 , n55456 );
not ( n55458 , n35983 );
not ( n55459 , n382912 );
or ( n55460 , n55458 , n55459 );
and ( n55461 , n382931 , n35987 );
not ( n55462 , RI15b5b9e0_991);
or ( n55463 , n35996 , n55462 );
or ( n55464 , n40296 , n36003 );
or ( n55465 , n35994 , n382967 );
nand ( n55466 , n55463 , n55464 , n55465 );
nor ( n55467 , n55461 , n55466 );
nand ( n55468 , n55460 , n55467 );
buf ( n55469 , n55468 );
buf ( n55470 , n384700 );
buf ( n55471 , n380203 );
not ( n55472 , RI15b55d88_794);
not ( n55473 , n380000 );
or ( n55474 , n55472 , n55473 );
and ( n55475 , n41919 , n381696 );
not ( n55476 , RI15b55d88_794);
not ( n55477 , n379964 );
not ( n55478 , n55477 );
or ( n55479 , n55476 , n55478 );
or ( n55480 , n55477 , RI15b55d88_794);
nand ( n55481 , n55479 , n55480 );
and ( n55482 , n379949 , n55481 );
nor ( n55483 , n55475 , n55482 );
nand ( n55484 , n55474 , n55483 );
buf ( n55485 , n55484 );
not ( n55486 , n381570 );
not ( n55487 , n33400 );
or ( n55488 , n55486 , n55487 );
and ( n55489 , n33415 , n381599 );
or ( n55490 , n381609 , n18461 );
or ( n55491 , n36293 , n381619 );
or ( n55492 , n381607 , n33443 );
nand ( n55493 , n55490 , n55491 , n55492 );
nor ( n55494 , n55489 , n55493 );
nand ( n55495 , n55488 , n55494 );
buf ( n55496 , n55495 );
buf ( n55497 , n22009 );
buf ( n55498 , n32672 );
buf ( n55499 , n380903 );
and ( n55500 , RI15b52458_672 , RI15b54780_747);
nor ( n55501 , n55500 , n45856 );
not ( n55502 , n55501 );
buf ( n55503 , n55502 );
and ( n55504 , n31770 , RI15b5ca48_1026);
or ( n55505 , n32378 , n384318 );
or ( n55506 , n31779 , n384441 );
nand ( n55507 , n55505 , n55506 );
nor ( n55508 , n31793 , n384565 );
nor ( n55509 , n55504 , n55507 , n55508 );
nand ( n55510 , n45095 , n55509 );
buf ( n55511 , n55510 );
buf ( n55512 , n386760 );
not ( n55513 , n41308 );
not ( n55514 , n386465 );
and ( n55515 , n55513 , n55514 );
or ( n55516 , n386541 , n385849 );
or ( n55517 , n48517 , n386550 );
or ( n55518 , n48504 , n386557 );
nand ( n55519 , n55516 , n55517 , n55518 );
nor ( n55520 , n55515 , n55519 );
nand ( n55521 , n48531 , n55520 );
buf ( n55522 , n55521 );
buf ( n55523 , n382537 );
buf ( n55524 , n381004 );
buf ( n55525 , n381872 );
buf ( n55526 , n31033 );
not ( n55527 , RI15b50478_604);
not ( n55528 , n385164 );
or ( n55529 , n55527 , n55528 );
and ( n55530 , n36473 , n21679 );
or ( n55531 , n385170 , n21276 );
or ( n55532 , n385178 , n45260 );
nand ( n55533 , n55531 , n55532 );
nor ( n55534 , n55530 , n55533 );
nand ( n55535 , n55529 , n55534 );
nor ( n55536 , n55285 , n55535 );
not ( n55537 , n55536 );
buf ( n55538 , n55537 );
buf ( n55539 , n22005 );
buf ( n55540 , n381004 );
not ( n55541 , RI15b5ea28_1094);
not ( n55542 , n384918 );
or ( n55543 , n55541 , n55542 );
and ( n55544 , n49762 , n384934 );
not ( n55545 , n384920 );
or ( n55546 , n32307 , n55545 );
nand ( n55547 , n55546 , n384925 );
and ( n55548 , n55547 , n32289 );
nor ( n55549 , n55544 , n55548 , n40496 );
nand ( n55550 , n55543 , n55549 );
buf ( n55551 , n55550 );
not ( n55552 , RI15b49470_365);
or ( n55553 , n381056 , n55552 );
and ( n55554 , n386555 , RI15b3ffd8_48);
not ( n55555 , RI15b49470_365);
and ( n55556 , n381064 , n55555 );
not ( n55557 , n381064 );
and ( n55558 , n55557 , RI15b49470_365);
nor ( n55559 , n55556 , n55558 );
and ( n55560 , n36064 , n55559 );
nor ( n55561 , n55554 , n55560 );
nand ( n55562 , n55553 , n55561 );
buf ( n55563 , n55562 );
buf ( n55564 , n33250 );
buf ( n55565 , n22404 );
buf ( n55566 , n384700 );
buf ( n55567 , n381872 );
or ( n55568 , n44431 , n22289 );
nand ( n55569 , n35525 , RI15b53538_708);
nand ( n55570 , n55568 , n55569 );
buf ( n55571 , n55570 );
and ( n55572 , n40008 , RI15b48228_326);
and ( n55573 , n54654 , n385219 );
nor ( n55574 , n55573 , RI15b3fab0_37);
nor ( n55575 , n55572 , n55574 );
not ( n55576 , n55575 );
buf ( n55577 , n55576 );
buf ( n55578 , n21800 );
buf ( n55579 , n380906 );
buf ( n55580 , n382065 );
buf ( n55581 , n30992 );
buf ( n55582 , n380942 );
buf ( n55583 , n382441 );
and ( n55584 , n42129 , n55583 );
nand ( n55585 , n382080 , n382160 );
nand ( n55586 , n382474 , n55585 );
nor ( n55587 , n55584 , n55586 );
or ( n55588 , n55587 , n382284 );
or ( n55589 , n382487 , n382160 );
or ( n55590 , n382512 , n55583 );
nand ( n55591 , n55589 , n55590 );
nand ( n55592 , n55591 , n382284 );
and ( n55593 , n382510 , n382445 );
and ( n55594 , n42153 , RI15b450f0_221);
nor ( n55595 , n55593 , n55594 );
nand ( n55596 , n55588 , n55592 , n55595 );
buf ( n55597 , n55596 );
buf ( n55598 , n21800 );
buf ( n55599 , n22714 );
buf ( n55600 , n386563 );
buf ( n55601 , n32271 );
or ( n55602 , n31149 , n40468 );
and ( n55603 , n31161 , n40470 );
not ( n55604 , RI15b4fc80_587);
or ( n55605 , n40480 , n55604 );
or ( n55606 , n32452 , n40485 );
or ( n55607 , n40478 , n31184 );
nand ( n55608 , n55605 , n55606 , n55607 );
nor ( n55609 , n55603 , n55608 );
nand ( n55610 , n55602 , n55609 );
buf ( n55611 , n55610 );
buf ( n55612 , n22343 );
nand ( n55613 , n41173 , n33433 );
nand ( n55614 , n384918 , RI15b5f220_1111);
nand ( n55615 , n37773 , RI15b60f30_1173);
nand ( n55616 , n54971 , n55613 , n55614 , n55615 );
buf ( n55617 , n55616 );
buf ( n55618 , n380903 );
nand ( n55619 , n381406 , n33611 );
nand ( n55620 , n381486 , RI15b52d40_691);
nand ( n55621 , n41992 , RI15b54a50_753);
nand ( n55622 , n55619 , n34895 , n55620 , n55621 );
buf ( n55623 , n55622 );
not ( n55624 , n36276 );
not ( n55625 , n382912 );
or ( n55626 , n55624 , n55625 );
and ( n55627 , n382931 , n36282 );
not ( n55628 , RI15b5c160_1007);
or ( n55629 , n36291 , n55628 );
or ( n55630 , n38307 , n36296 );
or ( n55631 , n36289 , n382967 );
nand ( n55632 , n55629 , n55630 , n55631 );
nor ( n55633 , n55627 , n55632 );
nand ( n55634 , n55626 , n55633 );
buf ( n55635 , n55634 );
buf ( n55636 , n382049 );
buf ( n55637 , n383498 );
and ( n55638 , n385164 , RI15b504f0_605);
or ( n55639 , n54737 , n21668 );
or ( n55640 , n21270 , n385170 );
or ( n55641 , n45257 , n385178 );
nand ( n55642 , n55639 , n55640 , n55641 );
nor ( n55643 , n55638 , n55642 );
nand ( n55644 , n45270 , n55643 );
buf ( n55645 , n55644 );
buf ( n55646 , n382069 );
not ( n55647 , RI15b5e9b0_1093);
not ( n55648 , n384918 );
or ( n55649 , n55647 , n55648 );
or ( n55650 , n384921 , n50810 );
nand ( n55651 , n55650 , n384925 );
and ( n55652 , n55651 , n50813 );
not ( n55653 , n384934 );
not ( n55654 , n50815 );
or ( n55655 , n55653 , n55654 );
nand ( n55656 , n55655 , n49953 );
nor ( n55657 , n55652 , n55656 );
nand ( n55658 , n55649 , n55657 );
buf ( n55659 , n55658 );
buf ( n55660 , n35651 );
or ( n55661 , n34720 , n34716 );
nor ( n55662 , n34716 , RI15b54618_744);
or ( n55663 , n55662 , n43011 );
nand ( n55664 , n55663 , n34715 );
nand ( n55665 , n55661 , n55664 );
buf ( n55666 , n55665 );
or ( n55667 , n383180 , n33219 );
not ( n55668 , n33237 );
and ( n55669 , n55668 , RI15b5a978_956);
or ( n55670 , n383184 , n33225 );
or ( n55671 , n32696 , n33241 );
or ( n55672 , n33235 , n383192 );
nand ( n55673 , n55670 , n55671 , n55672 );
nor ( n55674 , n55669 , n55673 );
nand ( n55675 , n55667 , n55674 );
buf ( n55676 , n55675 );
buf ( n55677 , n381006 );
buf ( n55678 , n32672 );
buf ( n55679 , n381004 );
buf ( n55680 , n382065 );
not ( n55681 , n43089 );
nor ( n55682 , n55681 , n382079 );
or ( n55683 , n55682 , n32024 );
nand ( n55684 , n55683 , n32855 );
nor ( n55685 , n32035 , n32855 );
not ( n55686 , n55685 );
not ( n55687 , n55681 );
or ( n55688 , n55686 , n55687 );
not ( n55689 , n42129 );
not ( n55690 , n55689 );
not ( n55691 , n382347 );
not ( n55692 , n32847 );
and ( n55693 , n55691 , n55692 );
and ( n55694 , n382347 , n32847 );
nor ( n55695 , n55693 , n55694 );
not ( n55696 , n55695 );
and ( n55697 , n55690 , n55696 );
not ( n55698 , RI15b45708_234);
not ( n55699 , n33159 );
or ( n55700 , n55698 , n55699 );
or ( n55701 , n43048 , n382114 );
nand ( n55702 , n55700 , n55701 );
nor ( n55703 , n55697 , n55702 );
nand ( n55704 , n55688 , n55703 );
not ( n55705 , n55704 );
nand ( n55706 , n55684 , n55705 );
buf ( n55707 , n55706 );
buf ( n55708 , n33250 );
buf ( n55709 , n19653 );
buf ( n55710 , n379893 );
buf ( n55711 , n35651 );
not ( n55712 , n21745 );
not ( n55713 , n55712 );
not ( n55714 , n44728 );
nand ( n55715 , n46002 , n21691 );
nand ( n55716 , n55714 , n55715 );
not ( n55717 , n55716 );
or ( n55718 , n55713 , n55717 );
not ( n55719 , n21248 );
not ( n55720 , n55719 );
not ( n55721 , n21254 );
nor ( n55722 , n46005 , n55721 );
not ( n55723 , n55722 );
and ( n55724 , n55720 , n55723 );
and ( n55725 , n55722 , n55719 );
and ( n55726 , n55724 , n55725 );
not ( n55727 , n44740 );
and ( n55728 , n55726 , n55727 );
not ( n55729 , n21472 );
not ( n55730 , n21478 );
not ( n55731 , n55730 );
and ( n55732 , n55729 , n55731 );
and ( n55733 , n21472 , n55730 );
nor ( n55734 , n55732 , n55733 );
or ( n55735 , n55734 , n45531 );
or ( n55736 , n21750 , n379136 );
nand ( n55737 , n55735 , n55736 );
nor ( n55738 , n55728 , n55737 );
nand ( n55739 , n55718 , n55738 );
not ( n55740 , n55739 );
and ( n55741 , n21788 , RI15b56b20_823);
and ( n55742 , n44330 , n21768 );
not ( n55743 , n21848 );
and ( n55744 , n55743 , n17533 );
not ( n55745 , n55743 );
and ( n55746 , n55745 , RI15b56b20_823);
nor ( n55747 , n55744 , n55746 );
and ( n55748 , n55747 , n384112 );
nor ( n55749 , n55741 , n55742 , n55748 );
nand ( n55750 , n55740 , n55749 );
buf ( n55751 , n55750 );
or ( n55752 , n22596 , n18079 );
nand ( n55753 , n55752 , n18104 );
and ( n55754 , n55753 , RI15b56580_811);
nor ( n55755 , n17576 , n22564 );
and ( n55756 , n22559 , n55755 );
nor ( n55757 , n18197 , RI15b56580_811);
not ( n55758 , n55757 );
not ( n55759 , n22596 );
or ( n55760 , n55758 , n55759 );
and ( n55761 , n44714 , RI15b58380_875);
or ( n55762 , n22621 , n22622 , RI15b58380_875);
or ( n55763 , n22623 , RI15b58308_874);
nand ( n55764 , n55762 , n55763 );
and ( n55765 , n55764 , n18188 );
and ( n55766 , n18219 , RI15b57480_843);
nor ( n55767 , n55761 , n55765 , n55766 );
nand ( n55768 , n55760 , n55767 );
nor ( n55769 , n55754 , n55756 , n55768 );
nor ( n55770 , n22559 , n17506 );
or ( n55771 , n55770 , n379905 );
nand ( n55772 , n55771 , n22564 );
nand ( n55773 , n55769 , n55772 );
buf ( n55774 , n55773 );
buf ( n55775 , n384700 );
buf ( n55776 , n22655 );
buf ( n55777 , n379895 );
or ( n55778 , n36937 , n384704 );
and ( n55779 , n36946 , n384739 );
not ( n55780 , RI15b4fa28_582);
or ( n55781 , n384749 , n55780 );
or ( n55782 , n38403 , n384757 );
or ( n55783 , n384747 , n36955 );
nand ( n55784 , n55781 , n55782 , n55783 );
nor ( n55785 , n55779 , n55784 );
nand ( n55786 , n55778 , n55785 );
buf ( n55787 , n55786 );
buf ( n55788 , n22655 );
nand ( n55789 , n44037 , n39334 );
nand ( n55790 , n384918 , RI15b5f478_1116);
and ( n55791 , n384922 , n383539 );
nor ( n55792 , n55791 , n384927 );
not ( n55793 , n55792 );
not ( n55794 , n383546 );
and ( n55795 , n55793 , n55794 );
and ( n55796 , n384934 , n52880 );
nor ( n55797 , n55795 , n55796 );
nand ( n55798 , n39338 , n55789 , n55790 , n55797 );
buf ( n55799 , n55798 );
or ( n55800 , n385163 , n21280 );
and ( n55801 , n37878 , n21685 );
and ( n55802 , n32368 , n44735 );
and ( n55803 , n385177 , n21494 );
nor ( n55804 , n55801 , n55802 , n55803 );
nand ( n55805 , n55800 , n44754 , n55804 );
buf ( n55806 , n55805 );
buf ( n55807 , n35649 );
buf ( n55808 , n381004 );
not ( n55809 , RI15b5eaa0_1095);
not ( n55810 , n384918 );
or ( n55811 , n55809 , n55810 );
or ( n55812 , n49159 , n384921 );
nand ( n55813 , n55812 , n384925 );
and ( n55814 , n55813 , n49162 );
not ( n55815 , n384934 );
not ( n55816 , n49165 );
or ( n55817 , n55815 , n55816 );
nand ( n55818 , n55817 , n45462 );
nor ( n55819 , n55814 , n55818 );
nand ( n55820 , n55811 , n55819 );
buf ( n55821 , n55820 );
buf ( n55822 , n22007 );
and ( n55823 , n40674 , RI15b54528_742);
and ( n55824 , n47549 , RI15b513f0_637);
nor ( n55825 , n55823 , n55824 );
not ( n55826 , n55825 );
buf ( n55827 , n55826 );
buf ( n55828 , n385197 );
not ( n55829 , n40651 );
and ( n55830 , n40650 , n55829 );
not ( n55831 , n40650 );
not ( n55832 , n55829 );
and ( n55833 , n55831 , n55832 );
nor ( n55834 , n55830 , n55833 );
or ( n55835 , n55834 , n385039 );
buf ( n55836 , n34304 );
not ( n55837 , n55836 );
buf ( n55838 , n34310 );
not ( n55839 , n55838 );
or ( n55840 , n55837 , n55839 );
or ( n55841 , n55838 , n55836 );
nand ( n55842 , n55840 , n55841 );
and ( n55843 , n55842 , n22440 );
not ( n55844 , RI15b5dab0_1061);
not ( n55845 , n379796 );
or ( n55846 , n55844 , n55845 );
not ( n55847 , RI15b63ca8_1270);
or ( n55848 , n36518 , n55847 );
nand ( n55849 , n55846 , n55848 );
nor ( n55850 , n55843 , n55849 );
nand ( n55851 , n55835 , n55850 );
buf ( n55852 , n55851 );
buf ( n55853 , n380903 );
or ( n55854 , n42969 , n52054 );
not ( n55855 , n33455 );
not ( n55856 , n36268 );
or ( n55857 , n55855 , n55856 );
nand ( n55858 , n55857 , n381450 );
and ( n55859 , n55858 , n54840 );
and ( n55860 , n381461 , n54842 );
nor ( n55861 , n55859 , n55860 );
and ( n55862 , n52056 , n55861 );
nand ( n55863 , n381486 , RI15b53010_697);
nand ( n55864 , n55854 , n55862 , n55863 );
buf ( n55865 , n55864 );
not ( n55866 , n381494 );
not ( n55867 , n381589 );
or ( n55868 , n55866 , n55867 );
and ( n55869 , n381596 , n381528 );
or ( n55870 , n381544 , n18694 );
or ( n55871 , n42258 , n381557 );
or ( n55872 , n381542 , n381621 );
nand ( n55873 , n55870 , n55871 , n55872 );
nor ( n55874 , n55869 , n55873 );
nand ( n55875 , n55868 , n55874 );
buf ( n55876 , n55875 );
buf ( n55877 , n22406 );
buf ( n55878 , n379847 );
buf ( n55879 , n381566 );
or ( n55880 , n35852 , n38373 );
and ( n55881 , n45035 , RI15b42fa8_150);
or ( n55882 , n35856 , n38383 );
or ( n55883 , n35582 , n38389 );
or ( n55884 , n38377 , n35858 );
nand ( n55885 , n55882 , n55883 , n55884 );
nor ( n55886 , n55881 , n55885 );
nand ( n55887 , n55880 , n55886 );
buf ( n55888 , n55887 );
buf ( n55889 , n22408 );
buf ( n55890 , n387159 );
buf ( n55891 , n21800 );
buf ( n55892 , RI15b473a0_295);
buf ( n55893 , n32160 );
not ( n55894 , n34798 );
and ( n55895 , n55894 , RI15b4aa78_412);
or ( n55896 , n53674 , n22216 );
or ( n55897 , n34801 , RI15b4aa78_412);
nand ( n55898 , n55896 , n55897 );
nor ( n55899 , n55895 , n55898 );
nand ( n55900 , n54309 , n55899 );
buf ( n55901 , n55900 );
buf ( n55902 , n32255 );
buf ( n55903 , n30992 );
buf ( n55904 , n386898 );
not ( n55905 , n55904 );
and ( n55906 , n55905 , n19628 );
nor ( n55907 , n55906 , n386945 );
or ( n55908 , n55907 , n386904 );
and ( n55909 , n55904 , n45576 , n386904 );
and ( n55910 , n22450 , n30842 );
nor ( n55911 , n55910 , n383413 );
nor ( n55912 , n55911 , n379440 );
nor ( n55913 , n55909 , n55912 );
buf ( n55914 , n386986 );
or ( n55915 , n55914 , n387003 );
nand ( n55916 , n55915 , n383408 );
nand ( n55917 , n55916 , RI15b62628_1222);
nand ( n55918 , n55914 , n47516 , n38482 );
or ( n55919 , n30842 , n379439 , RI15b64428_1286);
or ( n55920 , n379440 , RI15b643b0_1285);
nand ( n55921 , n55919 , n55920 );
and ( n55922 , n22450 , n55921 );
and ( n55923 , n22423 , RI15b64428_1286);
and ( n55924 , n19599 , RI15b63528_1254);
nor ( n55925 , n55922 , n55923 , n55924 );
and ( n55926 , n55913 , n55917 , n55918 , n55925 );
nand ( n55927 , n55908 , n55926 );
buf ( n55928 , n55927 );
or ( n55929 , n36238 , n383877 );
not ( n55930 , RI15b4f050_561);
or ( n55931 , n55930 , n383903 );
not ( n55932 , n383911 );
and ( n55933 , n55932 , n36257 );
and ( n55934 , n383803 , n40519 );
and ( n55935 , n36261 , n383909 );
nor ( n55936 , n55933 , n55934 , n55935 );
nand ( n55937 , n55929 , n55931 , n55936 );
buf ( n55938 , n55937 );
buf ( n55939 , n380906 );
buf ( n55940 , n380942 );
not ( n55941 , n38974 );
not ( n55942 , n45668 );
and ( n55943 , n55941 , n55942 );
nor ( n55944 , n55943 , n383577 );
or ( n55945 , n55944 , n45678 );
and ( n55946 , n383601 , RI15b5fe50_1137);
and ( n55947 , n383603 , n45679 );
and ( n55948 , n383607 , RI15b5f6d0_1121);
nor ( n55949 , n55946 , n55947 , n55948 );
nand ( n55950 , n55945 , n55949 );
buf ( n55951 , n55950 );
buf ( n55952 , n379893 );
buf ( n55953 , n32271 );
not ( n55954 , RI15b53970_717);
not ( n55955 , n383170 );
or ( n55956 , n55954 , n55955 );
not ( n55957 , n40056 );
not ( n55958 , n33453 );
or ( n55959 , n55957 , n55958 );
nand ( n55960 , n55959 , n33465 );
and ( n55961 , n55960 , n40039 );
and ( n55962 , n33476 , n50945 );
and ( n55963 , n383147 , RI15b531f0_701);
nor ( n55964 , n55961 , n55962 , n55963 );
nand ( n55965 , n55956 , n55964 );
buf ( n55966 , n55965 );
or ( n55967 , n386588 , n33419 );
and ( n55968 , n386600 , n33417 );
not ( n55969 , RI15b5b530_981);
or ( n55970 , n33428 , n55969 );
or ( n55971 , n34706 , n33440 );
or ( n55972 , n33426 , n386627 );
nand ( n55973 , n55970 , n55971 , n55972 );
nor ( n55974 , n55968 , n55973 );
nand ( n55975 , n55967 , n55974 );
buf ( n55976 , n55975 );
buf ( n55977 , n22738 );
buf ( n55978 , n383613 );
buf ( n55979 , n385197 );
or ( n55980 , n36119 , n37663 );
and ( n55981 , n43131 , RI15b42828_134);
or ( n55982 , n35856 , n37673 );
or ( n55983 , n35582 , n37679 );
or ( n55984 , n37665 , n35858 );
nand ( n55985 , n55982 , n55983 , n55984 );
nor ( n55986 , n55981 , n55985 );
nand ( n55987 , n55980 , n55986 );
buf ( n55988 , n55987 );
buf ( n55989 , n385195 );
buf ( n55990 , n19651 );
and ( n55991 , n385164 , RI15b50dd8_624);
not ( n55992 , n33652 );
and ( n55993 , n55992 , n37947 );
not ( n55994 , n385170 );
and ( n55995 , n55994 , n37935 );
and ( n55996 , n385177 , n37978 );
nor ( n55997 , n55993 , n55995 , n55996 );
not ( n55998 , n55997 );
nor ( n55999 , n55991 , n55998 );
nand ( n56000 , n37961 , n37985 , n55999 );
buf ( n56001 , n56000 );
buf ( n56002 , n22408 );
buf ( n56003 , n383345 );
nor ( n56004 , n43310 , n43312 );
not ( n56005 , n56004 );
not ( n56006 , n34426 );
not ( n56007 , n56006 );
and ( n56008 , n56005 , n56007 );
and ( n56009 , n56004 , n56006 );
nor ( n56010 , n56008 , n56009 );
or ( n56011 , n56010 , n43241 );
buf ( n56012 , n34110 );
not ( n56013 , n56012 );
not ( n56014 , n43321 );
not ( n56015 , n36566 );
or ( n56016 , n56014 , n56015 );
buf ( n56017 , n34248 );
nand ( n56018 , n56016 , n56017 );
not ( n56019 , n56018 );
or ( n56020 , n56013 , n56019 );
or ( n56021 , n56018 , n56012 );
nand ( n56022 , n56020 , n56021 );
and ( n56023 , n56022 , n379785 );
not ( n56024 , RI15b5e0c8_1074);
not ( n56025 , n34651 );
or ( n56026 , n56024 , n56025 );
or ( n56027 , n36518 , n379436 );
nand ( n56028 , n56026 , n56027 );
nor ( n56029 , n56023 , n56028 );
nand ( n56030 , n56011 , n56029 );
buf ( n56031 , n56030 );
buf ( n56032 , n22408 );
or ( n56033 , n45830 , n382665 );
and ( n56034 , n382664 , n382665 , RI15b55428_774);
and ( n56035 , n382666 , RI15b554a0_775);
nor ( n56036 , n56034 , n56035 );
or ( n56037 , n382629 , n56036 );
and ( n56038 , n382885 , n380197 );
or ( n56039 , n382691 , n383675 );
nand ( n56040 , n56039 , n53051 );
nor ( n56041 , n56038 , n56040 );
nand ( n56042 , n56033 , n56037 , n56041 );
buf ( n56043 , n56042 );
not ( n56044 , n382898 );
not ( n56045 , n380703 );
or ( n56046 , n56044 , n56045 );
and ( n56047 , n380719 , n382934 );
not ( n56048 , RI15b59a00_923);
or ( n56049 , n382949 , n56048 );
or ( n56050 , n380782 , n382965 );
or ( n56051 , n382947 , n380790 );
nand ( n56052 , n56049 , n56050 , n56051 );
nor ( n56053 , n56047 , n56052 );
nand ( n56054 , n56046 , n56053 );
buf ( n56055 , n56054 );
buf ( n56056 , n382069 );
buf ( n56057 , n379403 );
buf ( n56058 , n385195 );
not ( n56059 , RI15b53ad8_720);
not ( n56060 , n383170 );
nor ( n56061 , n56059 , n56060 );
or ( n56062 , n383153 , n41854 );
and ( n56063 , n383147 , RI15b524d0_673);
nor ( n56064 , n56062 , n56063 );
nand ( n56065 , n56061 , n56064 );
buf ( n56066 , n56065 );
not ( n56067 , n35145 );
not ( n56068 , n381507 );
or ( n56069 , n56067 , n56068 );
and ( n56070 , n381524 , n35150 );
or ( n56071 , n35160 , n18388 );
or ( n56072 , n36413 , n35166 );
or ( n56073 , n35158 , n381560 );
nand ( n56074 , n56071 , n56072 , n56073 );
nor ( n56075 , n56070 , n56074 );
nand ( n56076 , n56069 , n56075 );
buf ( n56077 , n56076 );
buf ( n56078 , n382069 );
nor ( n56079 , n32035 , n44172 );
nor ( n56080 , n44169 , n56079 );
or ( n56081 , n56080 , n46994 );
not ( n56082 , n46992 );
nor ( n56083 , n44167 , n56082 );
or ( n56084 , n56083 , n43098 );
nand ( n56085 , n56084 , n46994 );
not ( n56086 , n32870 );
not ( n56087 , n382414 );
or ( n56088 , n56086 , n56087 );
or ( n56089 , n382414 , n32870 );
nand ( n56090 , n56088 , n56089 );
and ( n56091 , n51184 , n56090 );
and ( n56092 , n382523 , RI15b4bbd0_449);
and ( n56093 , n42720 , RI15b459d8_240);
nor ( n56094 , n56092 , n56093 );
not ( n56095 , n56094 );
nor ( n56096 , n56091 , n56095 );
nand ( n56097 , n56081 , n56085 , n56096 );
buf ( n56098 , n56097 );
buf ( n56099 , n381490 );
buf ( n56100 , n383613 );
buf ( n56101 , n384199 );
buf ( n56102 , n387159 );
buf ( n56103 , n31030 );
or ( n56104 , n31006 , n33111 );
and ( n56105 , n31016 , n33117 );
or ( n56106 , n33128 , n21013 );
or ( n56107 , n33612 , n33134 );
or ( n56108 , n33126 , n31024 );
nand ( n56109 , n56106 , n56107 , n56108 );
nor ( n56110 , n56105 , n56109 );
nand ( n56111 , n56104 , n56110 );
buf ( n56112 , n56111 );
buf ( n56113 , n20665 );
and ( n56114 , n19549 , n19201 );
nor ( n56115 , n56114 , n40503 );
or ( n56116 , n56115 , n385189 );
and ( n56117 , n22431 , n22462 );
not ( n56118 , n380773 );
nor ( n56119 , n56117 , n384922 , n56118 );
nand ( n56120 , n56116 , n56119 );
buf ( n56121 , n56120 );
buf ( n56122 , n31979 );
buf ( n56123 , n379847 );
buf ( n56124 , n381566 );
or ( n56125 , n381907 , n38065 );
and ( n56126 , n43338 , RI15b42cd8_144);
or ( n56127 , n381917 , n38069 );
not ( n56128 , n38081 );
and ( n56129 , n56128 , n381923 );
and ( n56130 , n381926 , n38079 );
nor ( n56131 , n56129 , n56130 );
nand ( n56132 , n56127 , n56131 );
nor ( n56133 , n56126 , n56132 );
nand ( n56134 , n56125 , n56133 );
buf ( n56135 , n56134 );
buf ( n56136 , n384203 );
buf ( n56137 , n382067 );
buf ( n56138 , n22343 );
buf ( n56139 , n20665 );
or ( n56140 , n381907 , n35895 );
and ( n56141 , n35912 , RI15b40398_56);
or ( n56142 , n381917 , n35900 );
not ( n56143 , n35917 );
and ( n56144 , n56143 , n381923 );
and ( n56145 , n381926 , n35915 );
nor ( n56146 , n56144 , n56145 );
nand ( n56147 , n56142 , n56146 );
nor ( n56148 , n56141 , n56147 );
nand ( n56149 , n56140 , n56148 );
buf ( n56150 , n56149 );
or ( n56151 , n380968 , n35869 );
and ( n56152 , n380986 , n35872 );
or ( n56153 , n35884 , n385446 );
or ( n56154 , n380994 , n35888 );
or ( n56155 , n35882 , n380996 );
nand ( n56156 , n56153 , n56154 , n56155 );
nor ( n56157 , n56152 , n56156 );
nand ( n56158 , n56151 , n56157 );
buf ( n56159 , n56158 );
buf ( n56160 , n380203 );
buf ( n56161 , n30992 );
not ( n56162 , n31485 );
nand ( n56163 , n56162 , n34860 );
not ( n56164 , n31493 );
and ( n56165 , n56163 , n56164 );
not ( n56166 , n56163 );
and ( n56167 , n56166 , n31493 );
nor ( n56168 , n56165 , n56167 );
nand ( n56169 , n56168 , n31599 );
not ( n56170 , n31609 );
not ( n56171 , n31630 );
or ( n56172 , n56170 , n56171 );
or ( n56173 , n31630 , n31609 );
nand ( n56174 , n56172 , n56173 );
and ( n56175 , n56174 , n379391 );
and ( n56176 , n379394 , RI15b579a8_854);
and ( n56177 , n41206 , RI15b517b0_645);
nor ( n56178 , n56175 , n56176 , n56177 );
nand ( n56179 , n56169 , n56178 );
buf ( n56180 , n56179 );
buf ( n56181 , n385195 );
buf ( n56182 , n385197 );
buf ( n56183 , n19596 );
buf ( n56184 , n381872 );
not ( n56185 , n21716 );
not ( n56186 , n56185 );
not ( n56187 , n45244 );
not ( n56188 , n56187 );
or ( n56189 , n56186 , n56188 );
nand ( n56190 , n56189 , n47364 );
and ( n56191 , n56190 , n21748 );
not ( n56192 , n47371 );
not ( n56193 , n21290 );
and ( n56194 , n56192 , n56193 );
and ( n56195 , n47371 , n21290 );
nor ( n56196 , n56194 , n56195 );
or ( n56197 , n56196 , n21359 );
not ( n56198 , n21503 );
not ( n56199 , n47378 );
or ( n56200 , n56198 , n56199 );
or ( n56201 , n47378 , n21503 );
nand ( n56202 , n56200 , n56201 );
and ( n56203 , n56202 , n36442 );
and ( n56204 , n21751 , RI15b57c00_859);
nor ( n56205 , n56203 , n56204 );
nand ( n56206 , n56197 , n56205 );
nor ( n56207 , n56191 , n56206 );
and ( n56208 , n385164 , RI15b50568_606);
or ( n56209 , n33651 , n21716 );
or ( n56210 , n21290 , n385170 );
or ( n56211 , n21503 , n385178 );
nand ( n56212 , n56209 , n56210 , n56211 );
nor ( n56213 , n56208 , n56212 );
nand ( n56214 , n56207 , n56213 );
buf ( n56215 , n56214 );
buf ( n56216 , n381566 );
not ( n56217 , RI15b5e938_1092);
not ( n56218 , n384918 );
or ( n56219 , n56217 , n56218 );
and ( n56220 , n32275 , n50810 );
nor ( n56221 , n56220 , n51124 );
nand ( n56222 , n56219 , n56221 );
buf ( n56223 , n56222 );
not ( n56224 , n39923 );
not ( n56225 , n384122 );
or ( n56226 , n56224 , n56225 );
and ( n56227 , n384164 , n38828 );
or ( n56228 , n38837 , n17904 );
or ( n56229 , n42970 , n38841 );
or ( n56230 , n38835 , n384193 );
nand ( n56231 , n56228 , n56229 , n56230 );
nor ( n56232 , n56227 , n56231 );
nand ( n56233 , n56226 , n56232 );
buf ( n56234 , n56233 );
buf ( n56235 , n382071 );
buf ( n56236 , n380940 );
buf ( n56237 , n379403 );
and ( n56238 , n38487 , n386995 );
not ( n56239 , n38487 );
and ( n56240 , n56239 , RI15b62880_1227);
nor ( n56241 , n56238 , n56240 );
nand ( n56242 , n56241 , n384025 );
and ( n56243 , n384022 , RI15b62880_1227);
not ( n56244 , n44464 );
and ( n56245 , n386746 , n56244 );
nor ( n56246 , n56243 , n56245 );
nand ( n56247 , n56242 , n56246 );
buf ( n56248 , n56247 );
buf ( n56249 , n22402 );
buf ( n56250 , n17499 );
or ( n56251 , n22315 , n36306 );
and ( n56252 , n22326 , n36309 );
not ( n56253 , RI15b41a90_105);
or ( n56254 , n36318 , n56253 );
or ( n56255 , n22334 , n36325 );
or ( n56256 , n36316 , n22336 );
nand ( n56257 , n56254 , n56255 , n56256 );
nor ( n56258 , n56252 , n56257 );
nand ( n56259 , n56251 , n56258 );
buf ( n56260 , n56259 );
buf ( n56261 , RI15b5e140_1075);
buf ( n56262 , n384996 );
buf ( n56263 , n22788 );
buf ( n56264 , n22653 );
buf ( n56265 , n384203 );
not ( n56266 , n382670 );
and ( n56267 , n56266 , n383203 );
not ( n56268 , n56266 );
and ( n56269 , n56268 , RI15b55590_777);
nor ( n56270 , n56267 , n56269 );
not ( n56271 , n39526 );
nand ( n56272 , n56270 , n56271 );
and ( n56273 , n386637 , RI15b55590_777);
or ( n56274 , n382886 , n43545 );
or ( n56275 , n383686 , n382691 );
nor ( n56276 , n381400 , n32431 );
not ( n56277 , n56276 );
nand ( n56278 , n56274 , n56275 , n56277 );
nor ( n56279 , n56273 , n56278 );
nand ( n56280 , n56272 , n56279 );
buf ( n56281 , n56280 );
not ( n56282 , n382898 );
not ( n56283 , n381589 );
or ( n56284 , n56282 , n56283 );
and ( n56285 , n381596 , n382934 );
not ( n56286 , RI15b59910_921);
or ( n56287 , n382949 , n56286 );
or ( n56288 , n52325 , n382965 );
or ( n56289 , n382947 , n381621 );
nand ( n56290 , n56287 , n56288 , n56289 );
nor ( n56291 , n56285 , n56290 );
nand ( n56292 , n56284 , n56291 );
buf ( n56293 , n56292 );
buf ( n56294 , n22655 );
buf ( n56295 , n380940 );
or ( n56296 , n381056 , n19980 );
or ( n56297 , n32805 , n55031 );
not ( n56298 , n37119 );
and ( n56299 , n56298 , RI15b49b78_380);
not ( n56300 , n56298 );
and ( n56301 , n56300 , n19980 );
nor ( n56302 , n56299 , n56301 );
or ( n56303 , n43461 , n56302 );
nand ( n56304 , n56296 , n56297 , n56303 );
buf ( n56305 , n56304 );
buf ( n56306 , n32981 );
buf ( n56307 , n22479 );
buf ( n56308 , n32676 );
buf ( n56309 , n22653 );
not ( n56310 , RI15b53d30_725);
not ( n56311 , n32244 );
or ( n56312 , n56310 , n56311 );
and ( n56313 , n32247 , RI15b65328_1318);
and ( n56314 , n32249 , RI15b60198_1144);
nor ( n56315 , n56313 , n56314 );
nand ( n56316 , n56312 , n56315 );
buf ( n56317 , n56316 );
not ( n56318 , n39380 );
not ( n56319 , n384122 );
or ( n56320 , n56318 , n56319 );
and ( n56321 , n384164 , n31164 );
or ( n56322 , n31175 , n17883 );
or ( n56323 , n46471 , n31182 );
or ( n56324 , n31173 , n384193 );
nand ( n56325 , n56322 , n56323 , n56324 );
nor ( n56326 , n56321 , n56325 );
nand ( n56327 , n56320 , n56326 );
buf ( n56328 , n56327 );
buf ( n56329 , n33250 );
buf ( n56330 , n381006 );
not ( n56331 , n44290 );
or ( n56332 , n31053 , n56331 );
and ( n56333 , n36536 , RI15b61200_1179);
and ( n56334 , n384002 , n39368 );
not ( n56335 , RI15b61200_1179);
not ( n56336 , n31071 );
or ( n56337 , n56335 , n56336 );
or ( n56338 , n31071 , RI15b61200_1179);
nand ( n56339 , n56337 , n56338 );
and ( n56340 , n47154 , n56339 );
nor ( n56341 , n56333 , n56334 , n56340 );
nand ( n56342 , n56332 , n44288 , n56341 );
buf ( n56343 , n56342 );
buf ( n56344 , n30992 );
buf ( n56345 , n22007 );
or ( n56346 , n36937 , n40468 );
and ( n56347 , n36946 , n40470 );
not ( n56348 , RI15b4fde8_590);
or ( n56349 , n40480 , n56348 );
or ( n56350 , n36952 , n40485 );
or ( n56351 , n40478 , n36955 );
nand ( n56352 , n56349 , n56350 , n56351 );
nor ( n56353 , n56347 , n56352 );
nand ( n56354 , n56346 , n56353 );
buf ( n56355 , n56354 );
buf ( n56356 , n380940 );
not ( n56357 , RI15b5f0b8_1108);
not ( n56358 , n384918 );
or ( n56359 , n56357 , n56358 );
or ( n56360 , n384921 , RI15b60d50_1169);
nand ( n56361 , n56360 , n384925 , n384933 );
and ( n56362 , n56361 , RI15b60dc8_1170);
not ( n56363 , n49953 );
nor ( n56364 , n56362 , n56363 );
nand ( n56365 , n56359 , n56364 );
buf ( n56366 , n56365 );
and ( n56367 , n385164 , RI15b50388_602);
not ( n56368 , n21691 );
not ( n56369 , n36472 );
or ( n56370 , n56368 , n56369 );
and ( n56371 , n32368 , n21248 );
and ( n56372 , n385177 , n55730 );
nor ( n56373 , n56371 , n56372 );
nand ( n56374 , n56370 , n56373 );
nor ( n56375 , n56367 , n55739 , n56374 );
not ( n56376 , n56375 );
buf ( n56377 , n56376 );
buf ( n56378 , n379893 );
buf ( n56379 , n384996 );
not ( n56380 , RI15b5eb18_1096);
not ( n56381 , n384918 );
or ( n56382 , n56380 , n56381 );
not ( n56383 , n48928 );
and ( n56384 , n56383 , n384934 );
or ( n56385 , n48922 , n55545 );
nand ( n56386 , n56385 , n384925 );
and ( n56387 , n56386 , n32327 );
nor ( n56388 , n56384 , n56387 , n43842 );
nand ( n56389 , n56382 , n56388 );
buf ( n56390 , n56389 );
or ( n56391 , n19693 , n20638 );
nand ( n56392 , n56391 , n34798 );
nand ( n56393 , n56392 , RI15b4adc0_419);
and ( n56394 , n45068 , n22217 );
not ( n56395 , n34801 );
and ( n56396 , n56395 , n19693 , n19880 );
nor ( n56397 , n56394 , n56396 );
nand ( n56398 , n41265 , n56393 , n56397 );
buf ( n56399 , n56398 );
buf ( n56400 , n32672 );
buf ( n56401 , RI15b5dee8_1070);
buf ( n56402 , n382067 );
buf ( n56403 , n386762 );
buf ( n56404 , n379895 );
not ( n56405 , n386845 );
or ( n56406 , n56405 , n22473 );
nand ( n56407 , n56406 , n383474 );
nand ( n56408 , n56407 , n45100 );
not ( n56409 , n45100 );
nand ( n56410 , n56409 , n37068 , n56405 );
buf ( n56411 , n386974 );
nand ( n56412 , n43748 , n56411 );
or ( n56413 , n56412 , n40140 );
or ( n56414 , n56413 , n386975 );
not ( n56415 , n40144 );
and ( n56416 , n56415 , RI15b640e0_1279);
or ( n56417 , n34826 , n56411 , RI15b622e0_1215);
not ( n56418 , n387033 );
not ( n56419 , RI15b640e0_1279);
and ( n56420 , n56418 , n56419 );
and ( n56421 , n387033 , RI15b640e0_1279);
nor ( n56422 , n56420 , n56421 );
or ( n56423 , n34833 , n56422 );
nand ( n56424 , n56417 , n56423 );
nor ( n56425 , n56416 , n56424 );
nand ( n56426 , n56414 , n56425 );
nand ( n56427 , n56426 , n19201 );
and ( n56428 , n22423 , RI15b640e0_1279);
and ( n56429 , n19599 , RI15b631e0_1247);
nor ( n56430 , n56428 , n56429 , n19513 );
nand ( n56431 , n56408 , n56410 , n56427 , n56430 );
buf ( n56432 , n56431 );
buf ( n56433 , n387159 );
or ( n56434 , n36238 , n33116 );
not ( n56435 , n33128 );
and ( n56436 , n56435 , RI15b4e510_537);
or ( n56437 , n33134 , n32710 );
or ( n56438 , n33111 , n383802 );
or ( n56439 , n33126 , n42402 );
nand ( n56440 , n56437 , n56438 , n56439 );
nor ( n56441 , n56436 , n56440 );
nand ( n56442 , n56434 , n56441 );
buf ( n56443 , n56442 );
buf ( n56444 , n381004 );
nand ( n56445 , n52219 , n43197 );
buf ( n56446 , n56445 );
buf ( n56447 , n22402 );
or ( n56448 , n40166 , n386333 );
and ( n56449 , n386540 , RI15b43c50_177);
and ( n56450 , n386549 , n385558 );
and ( n56451 , n386556 , n386094 );
nor ( n56452 , n56449 , n56450 , n56451 );
nand ( n56453 , n56448 , n56452 , n54720 );
buf ( n56454 , n56453 );
buf ( n56455 , n33382 );
buf ( n56456 , n382537 );
buf ( n56457 , n382071 );
buf ( n56458 , n19651 );
not ( n56459 , n48629 );
and ( n56460 , n56459 , n34931 );
nor ( n56461 , n56460 , n35114 );
or ( n56462 , n56461 , n35098 );
and ( n56463 , n35118 , n48634 );
and ( n56464 , n20631 , RI15b46158_256);
nor ( n56465 , n56463 , n56464 );
nand ( n56466 , n385213 , RI15b47760_303);
nand ( n56467 , n56462 , n56465 , n56466 );
buf ( n56468 , n56467 );
buf ( n56469 , n382052 );
buf ( n56470 , n379844 );
buf ( n56471 , n385197 );
buf ( n56472 , n22788 );
buf ( n56473 , n382071 );
buf ( n56474 , n22653 );
and ( n56475 , n21788 , RI15b56d00_827);
and ( n56476 , n21885 , n42917 );
not ( n56477 , n17538 );
and ( n56478 , n56477 , n21881 );
not ( n56479 , n56477 );
and ( n56480 , n56479 , RI15b56d00_827);
nor ( n56481 , n56478 , n56480 );
and ( n56482 , n56481 , n37989 );
nor ( n56483 , n56475 , n56476 , n56482 );
nand ( n56484 , n56207 , n56483 );
buf ( n56485 , n56484 );
buf ( n56486 , n22530 );
nor ( n56487 , n56486 , n381826 );
and ( n56488 , n379855 , n56487 );
not ( n56489 , n22589 );
nor ( n56490 , n56489 , n18079 );
or ( n56491 , n56490 , n18103 );
nand ( n56492 , n56491 , RI15b563a0_807);
nor ( n56493 , n18197 , RI15b563a0_807);
and ( n56494 , n56489 , n56493 );
or ( n56495 , n47349 , n22838 );
or ( n56496 , n47347 , n22836 , RI15b581a0_871);
or ( n56497 , n22838 , RI15b58128_870);
nand ( n56498 , n56496 , n56497 );
and ( n56499 , n18188 , n56498 );
and ( n56500 , n18219 , RI15b572a0_839);
nor ( n56501 , n56499 , n56500 );
nand ( n56502 , n56495 , n56501 );
nor ( n56503 , n56494 , n56502 );
nand ( n56504 , n56492 , n56503 );
nor ( n56505 , n56488 , n56504 );
nand ( n56506 , n56486 , n17507 );
not ( n56507 , n56506 );
not ( n56508 , n17565 );
or ( n56509 , n56507 , n56508 );
nand ( n56510 , n56509 , n381826 );
nand ( n56511 , n56505 , n56510 );
buf ( n56512 , n56511 );
buf ( n56513 , n22404 );
buf ( n56514 , n20665 );
buf ( n56515 , n379893 );
xor ( n56516 , n39644 , n39619 );
not ( n56517 , n39662 );
or ( n56518 , n56516 , n56517 );
not ( n56519 , n379391 );
not ( n56520 , n39670 );
not ( n56521 , n56520 );
or ( n56522 , n56519 , n56521 );
nand ( n56523 , n56522 , n31700 );
and ( n56524 , n56523 , n31672 );
not ( n56525 , n31672 );
nand ( n56526 , n56525 , n39679 );
or ( n56527 , n56520 , n56526 );
and ( n56528 , n379394 , RI15b58380_875);
and ( n56529 , n39683 , RI15b52188_666);
nor ( n56530 , n56528 , n56529 );
nand ( n56531 , n56527 , n56530 );
nor ( n56532 , n56524 , n56531 );
nand ( n56533 , n56518 , n56532 );
buf ( n56534 , n56533 );
and ( n56535 , n31792 , n384543 );
or ( n56536 , n31771 , n384237 );
or ( n56537 , n48247 , n37611 );
or ( n56538 , n32643 , n31779 );
nand ( n56539 , n56536 , n56537 , n56538 );
nor ( n56540 , n56535 , n56539 );
nand ( n56541 , n48265 , n56540 );
buf ( n56542 , n56541 );
buf ( n56543 , n381081 );
buf ( n56544 , n380940 );
or ( n56545 , n32259 , n36813 );
and ( n56546 , n384983 , n37013 );
not ( n56547 , RI15b42378_124);
or ( n56548 , n36824 , n56547 );
or ( n56549 , n22022 , n36830 );
or ( n56550 , n36822 , n384988 );
nand ( n56551 , n56548 , n56549 , n56550 );
nor ( n56552 , n56546 , n56551 );
nand ( n56553 , n56545 , n56552 );
buf ( n56554 , n56553 );
buf ( n56555 , n383345 );
buf ( n56556 , n35649 );
buf ( n56557 , n381021 );
buf ( n56558 , n382071 );
or ( n56559 , n385173 , n385177 );
nand ( n56560 , n56559 , n21408 );
nand ( n56561 , n385164 , RI15b4ffc8_594);
nand ( n56562 , n32368 , n21093 );
nand ( n56563 , n56560 , n56561 , n56562 , n53954 );
buf ( n56564 , n56563 );
buf ( n56565 , n383613 );
and ( n56566 , n40778 , n40773 , n384934 );
not ( n56567 , RI15b5eed8_1104);
not ( n56568 , n384918 );
or ( n56569 , n56567 , n56568 );
nand ( n56570 , n56569 , n48610 );
nor ( n56571 , n56566 , n56570 );
nor ( n56572 , n40773 , n37776 );
or ( n56573 , n56572 , n37782 );
nand ( n56574 , n56573 , n40779 );
nand ( n56575 , n56571 , n56574 );
buf ( n56576 , n56575 );
buf ( n56577 , n386762 );
and ( n56578 , n43516 , RI15b47e68_318 , RI15b48318_328);
and ( n56579 , n385032 , RI15b48318_328);
not ( n56580 , n382509 );
nor ( n56581 , n56579 , n56580 );
nor ( n56582 , n56578 , n56581 );
nand ( n56583 , n56582 , n43514 , n385219 );
buf ( n56584 , n56583 );
buf ( n56585 , n380906 );
buf ( n56586 , n36854 );
buf ( n56587 , n30992 );
buf ( n56588 , n20663 );
buf ( n56589 , n32255 );
not ( n56590 , RI15b47508_298);
not ( n56591 , n385213 );
or ( n56592 , n56590 , n56591 );
and ( n56593 , n385221 , RI15b48a98_344);
and ( n56594 , n20631 , RI15b46d88_282);
nor ( n56595 , n56593 , n56594 );
nand ( n56596 , n56592 , n56595 );
buf ( n56597 , n56596 );
buf ( n56598 , n385197 );
buf ( n56599 , n383174 );
buf ( n56600 , n32255 );
not ( n56601 , RI15b46ef0_285);
not ( n56602 , n385213 );
or ( n56603 , n56601 , n56602 );
and ( n56604 , n385221 , RI15b48480_331);
and ( n56605 , n20631 , RI15b46770_269);
nor ( n56606 , n56604 , n56605 );
nand ( n56607 , n56603 , n56606 );
buf ( n56608 , n56607 );
buf ( n56609 , n382073 );
buf ( n56610 , n17499 );
buf ( n56611 , n22788 );
buf ( n56612 , n383498 );
buf ( n56613 , n18226 );
and ( n56614 , n21788 , RI15b56f58_832);
and ( n56615 , n22498 , n42917 );
buf ( n56616 , n22492 );
and ( n56617 , n56616 , n17546 );
not ( n56618 , n56616 );
and ( n56619 , n56618 , RI15b56f58_832);
nor ( n56620 , n56617 , n56619 );
and ( n56621 , n56620 , n37989 );
nor ( n56622 , n56614 , n56615 , n56621 );
nand ( n56623 , n44421 , n56622 );
buf ( n56624 , n56623 );
not ( n56625 , n22500 );
nor ( n56626 , n56625 , n22507 );
and ( n56627 , n379855 , n56626 );
buf ( n56628 , n22581 );
and ( n56629 , n56628 , n18086 );
nor ( n56630 , n56629 , n18103 );
or ( n56631 , n56630 , n22582 );
and ( n56632 , n18219 , RI15b57048_834);
nor ( n56633 , n56628 , n18197 , RI15b56148_802);
nor ( n56634 , n18189 , n42887 , RI15b57f48_866);
nor ( n56635 , n56632 , n56633 , n56634 );
not ( n56636 , n18178 );
not ( n56637 , n42889 );
or ( n56638 , n56636 , n56637 );
nand ( n56639 , n56638 , RI15b57f48_866);
nand ( n56640 , n56631 , n56635 , n56639 );
nor ( n56641 , n56627 , n56640 );
not ( n56642 , n17507 );
not ( n56643 , n56625 );
or ( n56644 , n56642 , n56643 );
nand ( n56645 , n56644 , n17565 );
nand ( n56646 , n56645 , n22507 );
nand ( n56647 , n56641 , n56646 );
buf ( n56648 , n56647 );
buf ( n56649 , n382049 );
buf ( n56650 , n383613 );
buf ( n56651 , n387159 );
and ( n56652 , n22646 , RI15b459d8_240);
and ( n56653 , n22648 , RI15b51e40_659);
nor ( n56654 , n56652 , n56653 );
not ( n56655 , n56654 );
buf ( n56656 , n56655 );
or ( n56657 , n383814 , n386706 );
and ( n56658 , n383857 , n386718 );
or ( n56659 , n386727 , n21135 );
or ( n56660 , n41099 , n386735 );
or ( n56661 , n386725 , n383917 );
nand ( n56662 , n56659 , n56660 , n56661 );
nor ( n56663 , n56658 , n56662 );
nand ( n56664 , n56657 , n56663 );
buf ( n56665 , n56664 );
buf ( n56666 , n379847 );
or ( n56667 , n384021 , n384035 );
and ( n56668 , n386746 , RI15b58b00_891);
and ( n56669 , n384034 , n384035 );
not ( n56670 , n384034 );
and ( n56671 , n56670 , RI15b61f98_1208);
nor ( n56672 , n56669 , n56671 );
and ( n56673 , n384025 , n56672 );
nor ( n56674 , n56668 , n56673 );
nand ( n56675 , n56667 , n56674 );
buf ( n56676 , n56675 );
buf ( n56677 , n381021 );
buf ( n56678 , n22406 );
buf ( n56679 , n22479 );
not ( n56680 , n42701 );
nor ( n56681 , n56680 , n382079 );
or ( n56682 , n56681 , n32024 );
nand ( n56683 , n56682 , n32009 );
and ( n56684 , n56680 , n51904 , n42702 );
not ( n56685 , n382289 );
nand ( n56686 , n56685 , n50488 );
not ( n56687 , n56686 );
buf ( n56688 , n31997 );
not ( n56689 , n56688 );
and ( n56690 , n56687 , n56689 );
and ( n56691 , n56686 , n56688 );
nor ( n56692 , n56690 , n56691 );
or ( n56693 , n382513 , n56692 );
and ( n56694 , n382523 , RI15b4b6a8_438);
and ( n56695 , n33159 , RI15b454b0_229);
nor ( n56696 , n56694 , n56695 );
nand ( n56697 , n56693 , n56696 );
nor ( n56698 , n56684 , n56697 );
nand ( n56699 , n56683 , n56698 );
buf ( n56700 , n56699 );
buf ( n56701 , n387159 );
buf ( n56702 , n384199 );
buf ( n56703 , n35651 );
buf ( n56704 , n32672 );
not ( n56705 , n385801 );
not ( n56706 , n56705 );
nor ( n56707 , n30868 , n49405 );
not ( n56708 , n56707 );
or ( n56709 , n56706 , n56708 );
or ( n56710 , n56707 , n56705 );
nand ( n56711 , n56709 , n56710 );
and ( n56712 , n56711 , n386018 );
not ( n56713 , n386140 );
not ( n56714 , n386146 );
not ( n56715 , n56714 );
and ( n56716 , n56713 , n56715 );
and ( n56717 , n386140 , n56714 );
nor ( n56718 , n56716 , n56717 );
or ( n56719 , n56718 , n386261 );
or ( n56720 , n30891 , n386425 );
nand ( n56721 , n56720 , n44683 );
and ( n56722 , n56721 , n386500 );
and ( n56723 , n41300 , RI15b4b5b8_436);
nor ( n56724 , n56722 , n56723 );
nand ( n56725 , n56719 , n56724 );
nor ( n56726 , n56712 , n56725 );
and ( n56727 , n30908 , RI15b4a6b8_404);
or ( n56728 , n19780 , n22216 );
not ( n56729 , n19775 );
and ( n56730 , n56729 , RI15b4a6b8_404);
not ( n56731 , n56729 );
and ( n56732 , n56731 , n19666 );
nor ( n56733 , n56730 , n56732 );
or ( n56734 , n56733 , n20638 );
nand ( n56735 , n56728 , n56734 );
or ( n56736 , n56727 , n56735 );
and ( n56737 , n56726 , n56736 );
not ( n56738 , n56737 );
buf ( n56739 , n21800 );
buf ( n56740 , n384199 );
nor ( n56741 , n55117 , n386938 );
and ( n56742 , n386932 , n56741 );
not ( n56743 , n55112 );
or ( n56744 , n386999 , n56743 );
nand ( n56745 , n56744 , n383408 );
and ( n56746 , n56745 , RI15b629e8_1230);
nand ( n56747 , n47516 , n387001 );
or ( n56748 , n387000 , n56747 );
nand ( n56749 , n379451 , RI15b64770_1293);
or ( n56750 , n30850 , n56749 );
or ( n56751 , n379451 , RI15b64770_1293);
nand ( n56752 , n56750 , n56751 );
and ( n56753 , n56752 , n22450 );
and ( n56754 , n19599 , RI15b638e8_1262);
nor ( n56755 , n56753 , n56754 );
nand ( n56756 , n55124 , RI15b647e8_1294);
and ( n56757 , n56755 , n56756 );
nand ( n56758 , n56748 , n56757 );
nor ( n56759 , n56742 , n56746 , n56758 );
nor ( n56760 , n386932 , n22473 );
or ( n56761 , n56760 , n386946 );
nand ( n56762 , n56761 , n386938 );
nand ( n56763 , n56759 , n56762 );
buf ( n56764 , n56763 );
buf ( n56765 , n33250 );
or ( n56766 , n386705 , n33597 );
and ( n56767 , n386716 , n33600 );
not ( n56768 , RI15b4eab0_549);
or ( n56769 , n33609 , n56768 );
or ( n56770 , n44306 , n33615 );
or ( n56771 , n33607 , n386738 );
nand ( n56772 , n56769 , n56770 , n56771 );
nor ( n56773 , n56767 , n56772 );
nand ( n56774 , n56766 , n56773 );
buf ( n56775 , n56774 );
buf ( n56776 , n380942 );
not ( n56777 , n33581 );
not ( n56778 , n33574 );
or ( n56779 , n56777 , n56778 );
nand ( n56780 , n56779 , n33584 );
nand ( n56781 , n56780 , n49176 );
nand ( n56782 , n49175 , n49178 , n40781 );
and ( n56783 , n383601 , RI15b603f0_1149);
and ( n56784 , n383607 , RI15b5ede8_1102);
nor ( n56785 , n56783 , n56784 );
nand ( n56786 , n56781 , n56782 , n56785 );
buf ( n56787 , n56786 );
buf ( n56788 , n379895 );
buf ( n56789 , n381490 );
buf ( n56790 , n387159 );
not ( n56791 , RI15b46fe0_287);
not ( n56792 , n385213 );
or ( n56793 , n56791 , n56792 );
and ( n56794 , n385221 , RI15b48570_333);
and ( n56795 , n20631 , RI15b46860_271);
nor ( n56796 , n56794 , n56795 );
nand ( n56797 , n56793 , n56796 );
buf ( n56798 , n56797 );
buf ( n56799 , n381004 );
buf ( n56800 , n35651 );
buf ( n56801 , n31979 );
buf ( n56802 , RI15b5e398_1080);
or ( n56803 , n383814 , n36242 );
and ( n56804 , n383857 , n43075 );
or ( n56805 , n36250 , n21116 );
or ( n56806 , n41099 , n36254 );
or ( n56807 , n36248 , n383917 );
nand ( n56808 , n56805 , n56806 , n56807 );
nor ( n56809 , n56804 , n56808 );
nand ( n56810 , n56803 , n56809 );
buf ( n56811 , n56810 );
buf ( n56812 , n383345 );
not ( n56813 , n53790 );
nor ( n56814 , n56813 , RI15b61b60_1199);
nor ( n56815 , n53793 , n56814 );
or ( n56816 , n56815 , n383523 );
and ( n56817 , n31051 , n380713 );
nor ( n56818 , n45131 , n45125 , RI15b61bd8_1200);
and ( n56819 , n51158 , n56818 );
nor ( n56820 , n56817 , n56819 );
nand ( n56821 , n56816 , n56820 );
buf ( n56822 , n56821 );
buf ( n56823 , n31719 );
buf ( n56824 , n22716 );
buf ( n56825 , n382067 );
or ( n56826 , n51002 , n51034 );
and ( n56827 , n45378 , n44495 );
or ( n56828 , n35195 , n51000 , RI15b48a98_344);
not ( n56829 , n386548 );
or ( n56830 , n56829 , n22032 );
nand ( n56831 , n56828 , n56830 );
nor ( n56832 , n56827 , n56831 );
nand ( n56833 , n56826 , n56832 );
buf ( n56834 , n56833 );
buf ( n56835 , n384700 );
buf ( n56836 , n384199 );
not ( n56837 , RI15b66408_1354);
or ( n56838 , n381015 , n56837 );
nand ( n56839 , n35327 , RI15b53f10_729);
nand ( n56840 , n56838 , n56839 );
buf ( n56841 , n56840 );
not ( n56842 , n53360 );
or ( n56843 , n56842 , n45380 );
and ( n56844 , n381055 , RI15b49740_371);
not ( n56845 , RI15b49740_371);
not ( n56846 , n32817 );
not ( n56847 , n56846 );
or ( n56848 , n56845 , n56847 );
or ( n56849 , n56846 , RI15b49740_371);
nand ( n56850 , n56848 , n56849 );
and ( n56851 , n381076 , n56850 );
nor ( n56852 , n56844 , n56851 );
nand ( n56853 , n56843 , n56852 );
buf ( n56854 , n56853 );
buf ( n56855 , n20663 );
buf ( n56856 , n22479 );
buf ( n56857 , n386760 );
buf ( n56858 , n386563 );
not ( n56859 , RI15b54168_734);
not ( n56860 , n32244 );
or ( n56861 , n56859 , n56860 );
and ( n56862 , n32247 , RI15b65760_1327);
and ( n56863 , n32249 , RI15b605d0_1153);
nor ( n56864 , n56862 , n56863 );
nand ( n56865 , n56861 , n56864 );
buf ( n56866 , n56865 );
buf ( n56867 , n35651 );
not ( n56868 , n37129 );
and ( n56869 , n56868 , n19993 );
not ( n56870 , n56868 );
and ( n56871 , n56870 , RI15b49f38_388);
nor ( n56872 , n56869 , n56871 );
nand ( n56873 , n56872 , n37113 );
and ( n56874 , n381055 , RI15b49f38_388);
and ( n56875 , n386555 , n51345 );
nor ( n56876 , n56874 , n56875 );
nand ( n56877 , n56873 , n56876 );
buf ( n56878 , n56877 );
buf ( n56879 , n19655 );
buf ( n56880 , n32676 );
buf ( n56881 , n380906 );
not ( n56882 , RI15b53970_717);
not ( n56883 , n32244 );
or ( n56884 , n56882 , n56883 );
and ( n56885 , n32247 , RI15b64f68_1310);
and ( n56886 , n32249 , RI15b5fdd8_1136);
nor ( n56887 , n56885 , n56886 );
nand ( n56888 , n56884 , n56887 );
buf ( n56889 , n56888 );
buf ( n56890 , n20665 );
and ( n56891 , RI15b45ff0_253 , RI15b48318_328);
nor ( n56892 , n56891 , n54655 );
not ( n56893 , n56892 );
buf ( n56894 , n56893 );
buf ( n56895 , n21800 );
buf ( n56896 , n382073 );
buf ( n56897 , n33250 );
buf ( n56898 , n385195 );
not ( n56899 , n41992 );
not ( n56900 , n383327 );
or ( n56901 , n56899 , n56900 );
nand ( n56902 , n56901 , n381450 );
nand ( n56903 , n56902 , n383213 );
nor ( n56904 , n383213 , n381460 );
not ( n56905 , n56904 );
not ( n56906 , n383335 );
or ( n56907 , n56905 , n56906 );
and ( n56908 , n381486 , RI15b52b60_687);
nor ( n56909 , n56908 , n50127 );
nand ( n56910 , n56907 , n56909 );
not ( n56911 , n56910 );
nand ( n56912 , n56903 , n56911 );
buf ( n56913 , n56912 );
not ( n56914 , n36276 );
not ( n56915 , n380703 );
or ( n56916 , n56914 , n56915 );
and ( n56917 , n380719 , n36282 );
not ( n56918 , RI15b5c340_1011);
or ( n56919 , n36291 , n56918 );
or ( n56920 , n48871 , n36296 );
or ( n56921 , n36289 , n380790 );
nand ( n56922 , n56919 , n56920 , n56921 );
nor ( n56923 , n56917 , n56922 );
nand ( n56924 , n56916 , n56923 );
buf ( n56925 , n56924 );
buf ( n56926 , n380942 );
buf ( n56927 , n22716 );
buf ( n56928 , n31033 );
and ( n56929 , n42686 , n44495 );
and ( n56930 , n35335 , RI15b662a0_1351);
and ( n56931 , n48970 , RI15b48ed0_353);
not ( n56932 , n48970 );
not ( n56933 , RI15b48ed0_353);
and ( n56934 , n56932 , n56933 );
nor ( n56935 , n56931 , n56934 );
not ( n56936 , n48988 );
nor ( n56937 , n56935 , n56936 );
nor ( n56938 , n56929 , n56930 , n56937 );
nand ( n56939 , n48979 , RI15b48ed0_353);
nand ( n56940 , n56938 , n56939 , n41586 );
buf ( n56941 , n56940 );
buf ( n56942 , n382049 );
buf ( n56943 , n19651 );
or ( n56944 , n381015 , n22036 );
nand ( n56945 , n35525 , RI15b53ad8_720);
nand ( n56946 , n56944 , n56945 );
buf ( n56947 , n56946 );
or ( n56948 , n44669 , n386425 );
and ( n56949 , n386540 , RI15b43f20_183);
and ( n56950 , n386549 , n385801 );
and ( n56951 , n386556 , n56714 );
nor ( n56952 , n56949 , n56950 , n56951 );
nand ( n56953 , n56948 , n56726 , n56952 );
buf ( n56954 , n56953 );
buf ( n56955 , n33382 );
buf ( n56956 , n19655 );
buf ( n56957 , n20663 );
buf ( n56958 , n31033 );
or ( n56959 , n31149 , n38825 );
and ( n56960 , n31161 , n38828 );
or ( n56961 , n38837 , n17660 );
or ( n56962 , n31179 , n38841 );
or ( n56963 , n38835 , n31184 );
nand ( n56964 , n56961 , n56962 , n56963 );
nor ( n56965 , n56960 , n56964 );
nand ( n56966 , n56959 , n56965 );
buf ( n56967 , n56966 );
buf ( n56968 , n22402 );
buf ( n56969 , n382537 );
buf ( n56970 , n385112 );
not ( n56971 , n53426 );
or ( n56972 , n56971 , n38168 );
not ( n56973 , n53830 );
not ( n56974 , n386747 );
and ( n56975 , n56973 , n56974 );
nor ( n56976 , n387001 , RI15b62a60_1231);
and ( n56977 , n38499 , n56976 );
nor ( n56978 , n56975 , n56977 );
nand ( n56979 , n56972 , n56978 );
buf ( n56980 , n56979 );
buf ( n56981 , n19651 );
buf ( n56982 , n380865 );
and ( n56983 , n19926 , n20637 );
nor ( n56984 , n56983 , n55894 );
or ( n56985 , n56984 , n19931 );
or ( n56986 , n34801 , n19926 , RI15b4b108_426);
or ( n56987 , n19933 , n22215 );
nand ( n56988 , n56986 , n56987 );
nor ( n56989 , n41828 , n56988 );
nand ( n56990 , n56985 , n56989 );
nor ( n56991 , n52016 , n56990 );
nand ( n56992 , n52000 , n56991 );
buf ( n56993 , n56992 );
buf ( n56994 , n382067 );
and ( n56995 , n22646 , RI15b45708_234);
and ( n56996 , n22648 , RI15b51b70_653);
nor ( n56997 , n56995 , n56996 );
not ( n56998 , n56997 );
buf ( n56999 , n56998 );
buf ( n57000 , n386762 );
buf ( n57001 , n379895 );
or ( n57002 , n34815 , n386964 );
nand ( n57003 , n57002 , n34823 );
and ( n57004 , n57003 , RI15b61f98_1208);
and ( n57005 , n34812 , RI15b63d98_1272);
not ( n57006 , n386964 );
or ( n57007 , n34826 , n57006 , RI15b61f98_1208);
not ( n57008 , n387025 );
not ( n57009 , n57008 );
not ( n57010 , RI15b63d98_1272);
and ( n57011 , n57009 , n57010 );
and ( n57012 , n57008 , RI15b63d98_1272);
nor ( n57013 , n57011 , n57012 );
or ( n57014 , n34833 , n57013 );
nand ( n57015 , n57007 , n57014 );
nor ( n57016 , n57004 , n57005 , n57015 );
or ( n57017 , n57016 , n19200 );
not ( n57018 , n386813 );
not ( n57019 , n57018 );
not ( n57020 , n22473 );
and ( n57021 , n57019 , n57020 );
nor ( n57022 , n57021 , n38114 );
or ( n57023 , n22774 , n57022 );
and ( n57024 , n387011 , n57018 , n22774 );
or ( n57025 , n22424 , n379530 );
or ( n57026 , n22772 , n19598 );
nand ( n57027 , n57025 , n57026 , n19512 );
nor ( n57028 , n57024 , n57027 );
nand ( n57029 , n57017 , n57023 , n57028 );
buf ( n57030 , n57029 );
buf ( n57031 , n385197 );
buf ( n57032 , n383613 );
or ( n57033 , n22102 , n38373 );
and ( n57034 , n22203 , n38375 );
or ( n57035 , n38385 , n20276 );
or ( n57036 , n22293 , n38389 );
or ( n57037 , n38383 , n22299 );
nand ( n57038 , n57035 , n57036 , n57037 );
nor ( n57039 , n57034 , n57038 );
nand ( n57040 , n57033 , n57039 );
buf ( n57041 , n57040 );
buf ( n57042 , n380903 );
buf ( n57043 , n22653 );
buf ( n57044 , n379895 );
and ( n57045 , n385164 , RI15b505e0_607);
or ( n57046 , n36693 , n21710 );
or ( n57047 , n21264 , n385170 );
or ( n57048 , n21499 , n385178 );
nand ( n57049 , n57046 , n57047 , n57048 );
nor ( n57050 , n57045 , n57049 );
nand ( n57051 , n47389 , n57050 );
buf ( n57052 , n57051 );
buf ( n57053 , n382065 );
and ( n57054 , RI15b5e8c0_1091 , RI15b60be8_1166);
nor ( n57055 , n57054 , n33102 );
not ( n57056 , n57055 );
buf ( n57057 , n57056 );
buf ( n57058 , n385195 );
and ( n57059 , n50535 , n383143 );
and ( n57060 , n383147 , RI15b52818_680);
nor ( n57061 , n57059 , n57060 );
nand ( n57062 , n383170 , RI15b53e20_727);
not ( n57063 , n383153 );
not ( n57064 , n50530 );
or ( n57065 , n57063 , n57064 );
nand ( n57066 , n57065 , n383157 );
nand ( n57067 , n57066 , n383139 );
nand ( n57068 , n57061 , n57062 , n57067 );
buf ( n57069 , n57068 );
not ( n57070 , n382976 );
not ( n57071 , n380703 );
or ( n57072 , n57070 , n57071 );
and ( n57073 , n380719 , n382983 );
or ( n57074 , n382995 , n19014 );
or ( n57075 , n37542 , n383001 );
or ( n57076 , n382993 , n380790 );
nand ( n57077 , n57074 , n57075 , n57076 );
nor ( n57078 , n57073 , n57077 );
nand ( n57079 , n57072 , n57078 );
buf ( n57080 , n57079 );
buf ( n57081 , n385197 );
buf ( n57082 , n22406 );
buf ( n57083 , n381081 );
and ( n57084 , n41267 , n386478 );
not ( n57085 , RI15b446a0_199);
or ( n57086 , n386541 , n57085 );
or ( n57087 , n385935 , n386550 );
or ( n57088 , n386557 , n386049 );
nand ( n57089 , n57086 , n57087 , n57088 );
nor ( n57090 , n57084 , n57089 );
nand ( n57091 , n38151 , n57090 );
buf ( n57092 , n57091 );
buf ( n57093 , n22343 );
buf ( n57094 , n31719 );
buf ( n57095 , n382052 );
buf ( n57096 , n22005 );
and ( n57097 , n382885 , n53139 );
not ( n57098 , RI15b553b0_773);
not ( n57099 , n382663 );
not ( n57100 , n57099 );
or ( n57101 , n57098 , n57100 );
or ( n57102 , n57099 , RI15b553b0_773);
nand ( n57103 , n57101 , n57102 );
and ( n57104 , n57103 , n32459 );
nor ( n57105 , n57097 , n57104 );
nand ( n57106 , n386637 , RI15b553b0_773);
and ( n57107 , n382692 , n383688 );
nor ( n57108 , n57107 , n50538 );
nand ( n57109 , n57105 , n57106 , n57108 );
buf ( n57110 , n57109 );
or ( n57111 , n386588 , n35792 );
and ( n57112 , n386600 , n35790 );
or ( n57113 , n35803 , n18622 );
or ( n57114 , n386618 , n35811 );
or ( n57115 , n35801 , n386627 );
nand ( n57116 , n57113 , n57114 , n57115 );
nor ( n57117 , n57112 , n57116 );
nand ( n57118 , n57111 , n57117 );
buf ( n57119 , n57118 );
buf ( n57120 , n22406 );
buf ( n57121 , n22655 );
not ( n57122 , n20637 );
not ( n57123 , n19698 );
or ( n57124 , n57122 , n57123 );
nand ( n57125 , n57124 , n34798 );
and ( n57126 , n57125 , RI15b4afa0_423);
or ( n57127 , n34801 , n19698 , RI15b4afa0_423);
not ( n57128 , n19905 );
or ( n57129 , n57128 , n22216 );
nand ( n57130 , n57127 , n57129 );
nor ( n57131 , n57126 , n57130 );
nand ( n57132 , n40763 , n57131 );
buf ( n57133 , n57132 );
buf ( n57134 , n381081 );
and ( n57135 , n22646 , RI15b45ca8_246);
and ( n57136 , n22648 , RI15b52110_665);
nor ( n57137 , n57135 , n57136 );
not ( n57138 , n57137 );
buf ( n57139 , n57138 );
buf ( n57140 , n382052 );
buf ( n57141 , n381081 );
buf ( n57142 , n35649 );
buf ( n57143 , n386816 );
or ( n57144 , n57143 , n22473 );
nand ( n57145 , n57144 , n386942 );
nand ( n57146 , n57145 , n386824 );
not ( n57147 , n386824 );
nand ( n57148 , n57147 , n45576 , n57143 );
not ( n57149 , n386968 );
and ( n57150 , n43748 , n57149 );
nor ( n57151 , n57150 , n40140 );
not ( n57152 , RI15b62100_1211);
or ( n57153 , n57151 , n57152 );
and ( n57154 , n56415 , RI15b63f00_1275);
or ( n57155 , n34826 , n57149 , RI15b62100_1211);
not ( n57156 , n387028 );
not ( n57157 , RI15b63f00_1275);
and ( n57158 , n57156 , n57157 );
and ( n57159 , n387028 , RI15b63f00_1275);
nor ( n57160 , n57158 , n57159 );
or ( n57161 , n34833 , n57160 );
nand ( n57162 , n57155 , n57161 );
nor ( n57163 , n57154 , n57162 );
nand ( n57164 , n57153 , n57163 );
nand ( n57165 , n57164 , n19201 );
and ( n57166 , n22423 , RI15b63f00_1275);
and ( n57167 , n19599 , RI15b63000_1243);
nor ( n57168 , n57166 , n57167 , n19513 );
nand ( n57169 , n57146 , n57148 , n57165 , n57168 );
buf ( n57170 , n57169 );
buf ( n57171 , n379893 );
buf ( n57172 , RI15b5dc90_1065);
not ( n57173 , n40341 );
or ( n57174 , n57173 , n40349 );
not ( n57175 , n50123 );
not ( n57176 , n52725 );
and ( n57177 , n57175 , n57176 );
nor ( n57178 , n22598 , RI15b565f8_812);
and ( n57179 , n40348 , n57178 );
nor ( n57180 , n57177 , n57179 );
nand ( n57181 , n57174 , n57180 );
buf ( n57182 , n57181 );
not ( n57183 , n380235 );
not ( n57184 , n37629 );
or ( n57185 , n57183 , n57184 );
and ( n57186 , n37637 , n380745 );
or ( n57187 , n380776 , n18992 );
or ( n57188 , n50080 , n380785 );
or ( n57189 , n380768 , n37646 );
nand ( n57190 , n57187 , n57188 , n57189 );
nor ( n57191 , n57186 , n57190 );
nand ( n57192 , n57185 , n57191 );
buf ( n57193 , n57192 );
buf ( n57194 , n382537 );
buf ( n57195 , n381006 );
or ( n57196 , n386705 , n39691 );
and ( n57197 , n386716 , n39694 );
not ( n57198 , RI15b4c8f0_477);
or ( n57199 , n39703 , n57198 );
or ( n57200 , n44306 , n39707 );
or ( n57201 , n39701 , n386738 );
nand ( n57202 , n57199 , n57200 , n57201 );
nor ( n57203 , n57197 , n57202 );
nand ( n57204 , n57196 , n57203 );
buf ( n57205 , n57204 );
buf ( n57206 , n31979 );
buf ( n57207 , n382537 );
buf ( n57208 , n381004 );
or ( n57209 , n44987 , n386985 );
and ( n57210 , n43831 , n42765 );
or ( n57211 , n44985 , n386983 , RI15b625b0_1221);
or ( n57212 , n386985 , RI15b62538_1220);
nand ( n57213 , n57211 , n57212 );
and ( n57214 , n57213 , n384025 );
nor ( n57215 , n57210 , n57214 );
nand ( n57216 , n57209 , n57215 );
buf ( n57217 , n57216 );
buf ( n57218 , n35651 );
buf ( n57219 , n379893 );
nor ( n57220 , n38286 , n41991 );
or ( n57221 , n57220 , n381449 );
not ( n57222 , n38290 );
nand ( n57223 , n57221 , n57222 );
nand ( n57224 , n38290 , n38286 , n381461 );
and ( n57225 , n32397 , RI15b529f8_684);
nor ( n57226 , n57225 , n56276 );
nand ( n57227 , n57223 , n57224 , n57226 );
buf ( n57228 , n57227 );
or ( n57229 , n31771 , n18593 );
or ( n57230 , n19328 , n44202 );
and ( n57231 , n32386 , n18595 );
and ( n57232 , n31778 , n19328 );
nor ( n57233 , n57231 , n57232 , n43602 );
nand ( n57234 , n57229 , n57230 , n57233 );
buf ( n57235 , n57234 );
buf ( n57236 , n22404 );
buf ( n57237 , n31719 );
nand ( n57238 , n40887 , RI15b51288_634);
or ( n57239 , n40881 , n57238 );
nand ( n57240 , n57239 , n18157 );
buf ( n57241 , n57240 );
buf ( n57242 , n385197 );
and ( n57243 , n44814 , n44816 );
not ( n57244 , n44814 );
not ( n57245 , n44816 );
and ( n57246 , n57244 , n57245 );
nor ( n57247 , n57243 , n57246 );
nand ( n57248 , n57247 , n22440 );
buf ( n57249 , n36555 );
and ( n57250 , n34282 , n57249 );
not ( n57251 , n34282 );
not ( n57252 , n57249 );
and ( n57253 , n57251 , n57252 );
nor ( n57254 , n57250 , n57253 );
nand ( n57255 , n57254 , n379785 );
and ( n57256 , n379783 , RI15b63e10_1273);
and ( n57257 , n34650 , RI15b5dc18_1064);
nor ( n57258 , n57256 , n57257 );
nand ( n57259 , n57248 , n57255 , n57258 );
buf ( n57260 , n57259 );
not ( n57261 , n47542 );
not ( n57262 , n384726 );
or ( n57263 , n57261 , n57262 );
and ( n57264 , n384737 , n35625 );
or ( n57265 , n35635 , n20806 );
or ( n57266 , n384754 , n35640 );
or ( n57267 , n35633 , n384759 );
nand ( n57268 , n57265 , n57266 , n57267 );
nor ( n57269 , n57264 , n57268 );
nand ( n57270 , n57263 , n57269 );
buf ( n57271 , n57270 );
buf ( n57272 , n22007 );
buf ( n57273 , n379403 );
not ( n57274 , n55398 );
and ( n57275 , n384918 , RI15b5f748_1122);
not ( n57276 , n53862 );
not ( n57277 , n384934 );
or ( n57278 , n57276 , n57277 );
and ( n57279 , n32274 , n53851 );
not ( n57280 , n384925 );
nor ( n57281 , n57279 , n57280 );
or ( n57282 , n57281 , n53858 );
nand ( n57283 , n57278 , n57282 );
nor ( n57284 , n57275 , n57283 );
nand ( n57285 , n57274 , n57284 );
buf ( n57286 , n57285 );
buf ( n57287 , n35649 );
and ( n57288 , n41309 , n34748 );
or ( n57289 , n386541 , n385843 );
or ( n57290 , n385906 , n386550 );
or ( n57291 , n386198 , n386557 );
nand ( n57292 , n57289 , n57290 , n57291 );
nor ( n57293 , n57288 , n57292 );
nand ( n57294 , n34790 , n57293 );
buf ( n57295 , n57294 );
buf ( n57296 , n22738 );
buf ( n57297 , n22655 );
buf ( n57298 , n381707 );
buf ( n57299 , n31033 );
buf ( n57300 , n32255 );
buf ( n57301 , n31033 );
and ( n57302 , n46838 , n50462 );
and ( n57303 , n35335 , RI15b65d00_1339);
not ( n57304 , RI15b48930_341);
not ( n57305 , n35348 );
not ( n57306 , n57305 );
or ( n57307 , n57304 , n57306 );
or ( n57308 , n57305 , RI15b48930_341);
nand ( n57309 , n57307 , n57308 );
and ( n57310 , n35363 , n57309 );
nor ( n57311 , n57302 , n57303 , n57310 );
nand ( n57312 , n41726 , RI15b48930_341);
nand ( n57313 , n45689 , n57311 , n57312 );
buf ( n57314 , n57313 );
buf ( n57315 , n382065 );
buf ( n57316 , n22714 );
or ( n57317 , n44431 , n22098 );
nand ( n57318 , n381017 , RI15b54078_732);
nand ( n57319 , n57317 , n57318 );
buf ( n57320 , n57319 );
not ( n57321 , n40519 );
not ( n57322 , n384122 );
or ( n57323 , n57321 , n57322 );
and ( n57324 , n384164 , n383878 );
or ( n57325 , n383903 , n20892 );
or ( n57326 , n46471 , n383911 );
or ( n57327 , n383895 , n384193 );
nand ( n57328 , n57325 , n57326 , n57327 );
nor ( n57329 , n57324 , n57328 );
nand ( n57330 , n57323 , n57329 );
buf ( n57331 , n57330 );
buf ( n57332 , n31719 );
buf ( n57333 , n383613 );
not ( n57334 , n38974 );
not ( n57335 , n46483 );
and ( n57336 , n57334 , n57335 );
nor ( n57337 , n57336 , n383577 );
or ( n57338 , n57337 , n383538 );
and ( n57339 , n383601 , RI15b5fb80_1131);
and ( n57340 , n383603 , n46488 );
and ( n57341 , n383607 , RI15b5f400_1115);
nor ( n57342 , n57339 , n57340 , n57341 );
nand ( n57343 , n57338 , n57342 );
buf ( n57344 , n57343 );
buf ( n57345 , n22740 );
buf ( n57346 , n382069 );
nor ( n57347 , n43421 , n43424 );
or ( n57348 , n57347 , n32958 );
buf ( n57349 , n43434 );
nand ( n57350 , n57348 , n57349 );
not ( n57351 , n43424 );
not ( n57352 , n54484 );
or ( n57353 , n57351 , n57352 );
not ( n57354 , n43430 );
nand ( n57355 , n57353 , n57354 );
not ( n57356 , n57349 );
and ( n57357 , n57355 , n57356 );
not ( n57358 , n382499 );
buf ( n57359 , n32943 );
not ( n57360 , n57359 );
and ( n57361 , n57358 , n57360 );
and ( n57362 , n382499 , n57359 );
nor ( n57363 , n57361 , n57362 );
or ( n57364 , n32964 , n57363 );
and ( n57365 , n382523 , RI15b4be28_454);
and ( n57366 , n43116 , RI15b45c30_245);
nor ( n57367 , n57365 , n57366 );
nand ( n57368 , n57364 , n57367 );
nor ( n57369 , n57357 , n57368 );
nand ( n57370 , n57350 , n57369 );
buf ( n57371 , n57370 );
buf ( n57372 , n22716 );
buf ( n57373 , n20663 );
buf ( n57374 , n33250 );
buf ( n57375 , n31033 );
or ( n57376 , n32525 , n385208 );
nand ( n57377 , n57376 , RI15b47e68_318);
or ( n57378 , n20516 , n19913 );
nand ( n57379 , n57378 , n379825 );
or ( n57380 , n39294 , n37554 );
not ( n57381 , n379824 );
or ( n57382 , n20579 , n57381 );
not ( n57383 , RI15b47e68_318);
or ( n57384 , n57383 , n20630 );
nand ( n57385 , n57380 , n57382 , n57384 );
nand ( n57386 , n57385 , n20492 );
and ( n57387 , n379824 , n36800 , n20516 );
nor ( n57388 , n57387 , n385207 );
nand ( n57389 , n57377 , n57379 , n57386 , n57388 );
buf ( n57390 , n57389 );
buf ( n57391 , n21800 );
buf ( n57392 , n383345 );
buf ( n57393 , n35649 );
buf ( n57394 , n22408 );
or ( n57395 , n382679 , n383018 );
and ( n57396 , n47697 , n386669 );
or ( n57397 , n382691 , n383641 );
not ( n57398 , n382655 );
and ( n57399 , n57398 , RI15b55158_768);
not ( n57400 , n57398 );
and ( n57401 , n57400 , n383018 );
nor ( n57402 , n57399 , n57401 );
or ( n57403 , n43699 , n57402 );
nand ( n57404 , n57397 , n57403 , n36351 );
nor ( n57405 , n57396 , n57404 );
nand ( n57406 , n57395 , n57405 );
buf ( n57407 , n57406 );
not ( n57408 , n35784 );
not ( n57409 , n381507 );
or ( n57410 , n57408 , n57409 );
and ( n57411 , n381524 , n35790 );
not ( n57412 , RI15b59d48_930);
or ( n57413 , n35803 , n57412 );
or ( n57414 , n38012 , n35811 );
or ( n57415 , n35801 , n381560 );
nand ( n57416 , n57413 , n57414 , n57415 );
nor ( n57417 , n57411 , n57416 );
and ( n57418 , n57410 , n57417 );
buf ( n57419 , n57418 );
buf ( n57420 , n379403 );
buf ( n57421 , n383345 );
or ( n57422 , n385163 , n21250 );
and ( n57423 , n385173 , n21662 );
and ( n57424 , n32368 , n21254 );
and ( n57425 , n385177 , n21471 );
nor ( n57426 , n57423 , n57424 , n57425 );
nand ( n57427 , n57422 , n57426 , n46022 );
buf ( n57428 , n57427 );
buf ( n57429 , n32271 );
buf ( n57430 , n384996 );
and ( n57431 , n49338 , n384922 );
nor ( n57432 , n57431 , n57280 );
or ( n57433 , n57432 , n32337 );
and ( n57434 , n49343 , n384934 );
nor ( n57435 , n57434 , n42643 );
nand ( n57436 , n384918 , RI15b5eb90_1097);
nand ( n57437 , n57433 , n57435 , n57436 );
buf ( n57438 , n57437 );
or ( n57439 , n20638 , RI15b4aa78_412);
nand ( n57440 , n57439 , n34798 );
and ( n57441 , n57440 , RI15b4aaf0_413);
or ( n57442 , n34801 , n19717 , RI15b4aaf0_413);
not ( n57443 , n19838 );
or ( n57444 , n57443 , n22216 );
nand ( n57445 , n57442 , n57444 );
nor ( n57446 , n57441 , n57445 );
nand ( n57447 , n44931 , n57446 );
buf ( n57448 , n57447 );
buf ( n57449 , n382065 );
buf ( n57450 , RI15b471c0_291);
buf ( n57451 , n32160 );
buf ( n57452 , n32255 );
buf ( n57453 , n31979 );
buf ( n57454 , n386984 );
and ( n57455 , n57454 , n54261 );
nor ( n57456 , n57455 , n383409 );
or ( n57457 , n57456 , n386985 );
nand ( n57458 , n55911 , n22424 );
and ( n57459 , n57458 , RI15b643b0_1285);
not ( n57460 , n386893 );
or ( n57461 , n57460 , n22473 );
nand ( n57462 , n57461 , n40133 );
not ( n57463 , n386897 );
and ( n57464 , n57462 , n57463 );
nor ( n57465 , n57459 , n57464 );
and ( n57466 , n57460 , n387011 , n386897 );
or ( n57467 , n57454 , n383482 , RI15b625b0_1221);
nor ( n57468 , n30842 , RI15b643b0_1285);
and ( n57469 , n22450 , n57468 );
and ( n57470 , n19599 , RI15b634b0_1253);
nor ( n57471 , n57469 , n57470 );
nand ( n57472 , n57467 , n57471 );
nor ( n57473 , n57466 , n57472 );
nand ( n57474 , n57457 , n57465 , n57473 );
buf ( n57475 , n57474 );
buf ( n57476 , n22408 );
or ( n57477 , n380001 , n379956 );
and ( n57478 , n380010 , RI15b4c620_471);
and ( n57479 , n379955 , n379956 );
not ( n57480 , n379955 );
and ( n57481 , n57480 , RI15b55ab8_788);
nor ( n57482 , n57479 , n57481 );
and ( n57483 , n379949 , n57482 );
nor ( n57484 , n57478 , n57483 );
nand ( n57485 , n57477 , n57484 );
buf ( n57486 , n57485 );
not ( n57487 , n36395 );
not ( n57488 , n37629 );
or ( n57489 , n57487 , n57488 );
and ( n57490 , n37637 , n36401 );
or ( n57491 , n36410 , n18990 );
or ( n57492 , n50080 , n36416 );
or ( n57493 , n36408 , n37646 );
nand ( n57494 , n57491 , n57492 , n57493 );
nor ( n57495 , n57490 , n57494 );
nand ( n57496 , n57489 , n57495 );
buf ( n57497 , n57496 );
buf ( n57498 , n379403 );
buf ( n57499 , n385112 );
not ( n57500 , n39150 );
not ( n57501 , n33370 );
or ( n57502 , n57500 , n57501 );
and ( n57503 , n33196 , n36123 );
or ( n57504 , n36132 , n20127 );
or ( n57505 , n22241 , n36139 );
or ( n57506 , n36130 , n33201 );
nand ( n57507 , n57504 , n57505 , n57506 );
nor ( n57508 , n57503 , n57507 );
nand ( n57509 , n57502 , n57508 );
buf ( n57510 , n57509 );
buf ( n57511 , n33382 );
buf ( n57512 , n379847 );
buf ( n57513 , n32271 );
buf ( n57514 , n382052 );
buf ( n57515 , n22788 );
not ( n57516 , RI15b53538_708);
not ( n57517 , n383170 );
or ( n57518 , n57516 , n57517 );
and ( n57519 , n33453 , RI15b54ac8_754);
and ( n57520 , n383147 , RI15b52db8_692);
nor ( n57521 , n57519 , n57520 );
nand ( n57522 , n57518 , n57521 );
buf ( n57523 , n57522 );
not ( n57524 , n35983 );
not ( n57525 , n37629 );
or ( n57526 , n57524 , n57525 );
and ( n57527 , n37637 , n35987 );
or ( n57528 , n35996 , n18566 );
or ( n57529 , n50208 , n36003 );
or ( n57530 , n35994 , n37646 );
nand ( n57531 , n57528 , n57529 , n57530 );
nor ( n57532 , n57527 , n57531 );
nand ( n57533 , n57526 , n57532 );
buf ( n57534 , n57533 );
buf ( n57535 , n22738 );
buf ( n57536 , n22788 );
not ( n57537 , RI15b53d30_725);
not ( n57538 , n383170 );
or ( n57539 , n57537 , n57538 );
or ( n57540 , n49133 , n383152 );
nand ( n57541 , n57540 , n383157 );
and ( n57542 , n57541 , n383128 );
and ( n57543 , n49138 , n383143 );
and ( n57544 , n383147 , RI15b52728_678);
nor ( n57545 , n57542 , n57543 , n57544 );
nand ( n57546 , n57539 , n57545 );
buf ( n57547 , n57546 );
or ( n57548 , n386588 , n35144 );
and ( n57549 , n386600 , n35150 );
not ( n57550 , RI15b5b170_973);
or ( n57551 , n35160 , n57550 );
or ( n57552 , n34706 , n35166 );
or ( n57553 , n35158 , n386627 );
nand ( n57554 , n57551 , n57552 , n57553 );
nor ( n57555 , n57549 , n57554 );
nand ( n57556 , n57548 , n57555 );
buf ( n57557 , n57556 );
buf ( n57558 , n17499 );
and ( C0 , n17501 , RI15b51198_632 );
endmodule

