//NOTE: no-implementation module stub

module REG12L (
    input wire DSPCLK,
    input wire IDR_enb,
    input wire IDR_we,
    input wire [11:0] IDR_di,
    output reg [11:0] IDR
);

endmodule
