//NOTE: no-implementation module stub

module GTECH_NOT (
    input wire A,
    output wire Z
);

endmodule
