//NOTE: no-implementation module stub

module REG8LCI (
    input wire DSPCLK,
    input wire MMR_web,
    input wire WSCR_ext_we,
    input wire [7:0] DMD,
    output reg [7:0] WSCR_ext,
    input wire RST
);

endmodule
