//NOTE: no-implementation module stub

module REG2D16L (
    input wire DSPCLK,
    input wire CLKMXOPenb,
    input wire MXOPwe,
    input wire [15:0] R_in_D,
    output reg [15:0] MXOPDI2,
    output reg [15:0] MXOP_E,
    input wire SCAN_TEST
);

endmodule
