// IWLS benchmark module "MinMax9b" printed on Wed May 29 22:12:27 2002
module MinMax9b(\1 , \2 , \3 , \4 , \5 , \6 , \7 , \8 , \9 , \10 , \11 , \12 , \39 , \40 , \41 , \42 , \43 , \44 , \45 , \46 , \47 );
input
  \1 ,
  \2 ,
  \3 ,
  \4 ,
  \5 ,
  \6 ,
  \7 ,
  \8 ,
  \9 ,
  \10 ,
  \11 ,
  \12 ;
output
  \39 ,
  \40 ,
  \41 ,
  \42 ,
  \43 ,
  \44 ,
  \45 ,
  \46 ,
  \47 ;
reg
  \13 ,
  \14 ,
  \15 ,
  \16 ,
  \17 ,
  \18 ,
  \19 ,
  \20 ,
  \21 ,
  \22 ,
  \23 ,
  \24 ,
  \25 ,
  \26 ,
  \27 ,
  \28 ,
  \29 ,
  \30 ,
  \31 ,
  \32 ,
  \33 ,
  \34 ,
  \35 ,
  \36 ,
  \37 ,
  \38 ;
wire
  \57 ,
  \58 ,
  \59 ,
  \60 ,
  \61 ,
  \62 ,
  \63 ,
  \64 ,
  \81 ,
  \83 ,
  \85 ,
  \87 ,
  \89 ,
  \91 ,
  \93 ,
  \95 ,
  \97 ,
  \99 ,
  \101 ,
  \105 ,
  \107 ,
  \109 ,
  \111 ,
  \113 ,
  \115 ,
  \117 ,
  \119 ,
  \121 ,
  \233 ,
  \260 ,
  \325 ,
  \326 ,
  \327 ,
  \328 ,
  \329 ,
  \330 ,
  \331 ,
  \332 ,
  \333 ,
  \365 ,
  \368 ,
  \371 ,
  \374 ,
  \377 ,
  \380 ,
  \383 ,
  \386 ,
  \389 ,
  \392 ,
  \395 ,
  \398 ,
  \401 ,
  \404 ,
  \407 ,
  \408 ,
  \409 ,
  \410 ,
  \411 ,
  \412 ,
  \413 ,
  \414 ,
  \415 ,
  \416 ,
  \417 ,
  \418 ,
  \419 ,
  \420 ,
  \421 ,
  \422 ,
  \423 ,
  \424 ,
  \425 ,
  \426 ,
  \427 ,
  \428 ,
  \430 ,
  \431 ,
  \432 ,
  \433 ,
  \434 ,
  \435 ,
  \436 ,
  \437 ,
  \438 ,
  \439 ,
  \440 ,
  \441 ,
  \442 ,
  \443 ,
  \444 ,
  \445 ,
  \446 ,
  \447 ,
  \448 ,
  \449 ,
  \450 ,
  \451 ,
  \452 ,
  \453 ,
  \454 ,
  \455 ,
  \456 ,
  \457 ,
  \458 ,
  \459 ,
  \460 ,
  \461 ,
  \462 ,
  \464 ,
  \465 ,
  \466 ,
  \467 ,
  \468 ,
  \469 ,
  \470 ,
  \472 ,
  \473 ,
  \474 ,
  \475 ,
  \476 ,
  \477 ,
  \478 ,
  \480 ,
  \481 ,
  \482 ,
  \483 ,
  \484 ,
  \485 ,
  \486 ,
  \488 ,
  \489 ,
  \490 ,
  \491 ,
  \492 ,
  \493 ,
  \494 ,
  \496 ,
  \497 ,
  \498 ,
  \499 ,
  \500 ,
  \501 ,
  \502 ,
  \504 ,
  \505 ,
  \506 ,
  \507 ,
  \508 ,
  \509 ,
  \510 ,
  \512 ,
  \513 ,
  \514 ,
  \515 ,
  \516 ,
  \517 ,
  \518 ,
  \520 ,
  \521 ,
  \522 ,
  \523 ,
  \524 ,
  \525 ,
  \526 ,
  \528 ,
  \529 ,
  \530 ,
  \531 ,
  \533 ,
  \534 ,
  \535 ,
  \536 ,
  \538 ,
  \539 ,
  \540 ,
  \541 ,
  \543 ,
  \544 ,
  \545 ,
  \546 ,
  \548 ,
  \549 ,
  \550 ,
  \551 ,
  \553 ,
  \554 ,
  \555 ,
  \556 ,
  \558 ,
  \559 ,
  \560 ,
  \561 ,
  \563 ,
  \564 ,
  \565 ,
  \566 ,
  \568 ,
  \569 ,
  \570 ,
  \571 ,
  \573 ,
  \575 ,
  \576 ,
  \578 ,
  \579 ,
  \581 ,
  \583 ,
  \584 ,
  \586 ,
  \587 ,
  \589 ,
  \591 ,
  \592 ,
  \594 ,
  \595 ,
  \597 ,
  \599 ,
  \[35] ,
  \[36] ,
  \600 ,
  \602 ,
  \603 ,
  \605 ,
  \607 ,
  \608 ,
  \[37] ,
  \610 ,
  \611 ,
  \613 ,
  \615 ,
  \616 ,
  \618 ,
  \619 ,
  \[38] ,
  \621 ,
  \623 ,
  \624 ,
  \626 ,
  \627 ,
  \629 ,
  \[39] ,
  \631 ,
  \632 ,
  \634 ,
  \635 ,
  \637 ,
  \640 ,
  \643 ,
  \645 ,
  \648 ,
  \651 ,
  \653 ,
  \656 ,
  \659 ,
  \661 ,
  \664 ,
  \667 ,
  \669 ,
  \672 ,
  \675 ,
  \677 ,
  \680 ,
  \683 ,
  \685 ,
  \688 ,
  \691 ,
  \693 ,
  \696 ,
  \699 ,
  \[40] ,
  \[41] ,
  \[42] ,
  \[43] ,
  \[44] ,
  \[45] ,
  \[46] ,
  \701 ,
  \702 ,
  \703 ,
  \704 ,
  \705 ,
  \706 ,
  \707 ,
  \708 ,
  \709 ,
  \[47] ,
  \710 ,
  \712 ,
  \713 ,
  \714 ,
  \715 ,
  \716 ,
  \717 ,
  \718 ,
  \719 ,
  \[48] ,
  \720 ,
  \721 ,
  \722 ,
  \723 ,
  \724 ,
  \725 ,
  \726 ,
  \727 ,
  \728 ,
  \729 ,
  \[49] ,
  \730 ,
  \731 ,
  \732 ,
  \733 ,
  \734 ,
  \735 ,
  \736 ,
  \737 ,
  \738 ,
  \739 ,
  \740 ,
  \741 ,
  \742 ,
  \743 ,
  \744 ,
  \745 ,
  \746 ,
  \747 ,
  \748 ,
  \749 ,
  \750 ,
  \751 ,
  \752 ,
  \753 ,
  \754 ,
  \755 ,
  \756 ,
  \757 ,
  \758 ,
  \759 ,
  \760 ,
  \761 ,
  \762 ,
  \763 ,
  \764 ,
  \765 ,
  \766 ,
  \767 ,
  \768 ,
  \769 ,
  \770 ,
  \771 ,
  \772 ,
  \773 ,
  \774 ,
  \775 ,
  \776 ,
  \777 ,
  \778 ,
  \779 ,
  \780 ,
  \781 ,
  \782 ,
  \783 ,
  \784 ,
  \785 ,
  \786 ,
  \787 ,
  \788 ,
  \789 ,
  \790 ,
  \791 ,
  \792 ,
  \793 ,
  \794 ,
  \795 ,
  \796 ,
  \797 ,
  \798 ,
  \799 ,
  \[50] ,
  \[51] ,
  \[52] ,
  \[53] ,
  \[54] ,
  \[55] ,
  \[56] ,
  \800 ,
  \801 ,
  \803 ,
  \805 ,
  \806 ,
  \807 ,
  \808 ,
  \809 ,
  \[57] ,
  \810 ,
  \811 ,
  \812 ,
  \813 ,
  \814 ,
  \815 ,
  \816 ,
  \817 ,
  \818 ,
  \819 ,
  \[58] ,
  \820 ,
  \821 ,
  \822 ,
  \823 ,
  \824 ,
  \825 ,
  \826 ,
  \827 ,
  \828 ,
  \829 ,
  \[59] ,
  \830 ,
  \831 ,
  \833 ,
  \834 ,
  \835 ,
  \836 ,
  \838 ,
  \839 ,
  \840 ,
  \841 ,
  \843 ,
  \844 ,
  \845 ,
  \846 ,
  \848 ,
  \849 ,
  \850 ,
  \851 ,
  \853 ,
  \854 ,
  \855 ,
  \856 ,
  \858 ,
  \859 ,
  \860 ,
  \861 ,
  \863 ,
  \864 ,
  \865 ,
  \866 ,
  \868 ,
  \869 ,
  \870 ,
  \871 ,
  \873 ,
  \874 ,
  \875 ,
  \877 ,
  \879 ,
  \880 ,
  \881 ,
  \882 ,
  \883 ,
  \884 ,
  \885 ,
  \886 ,
  \887 ,
  \888 ,
  \889 ,
  \890 ,
  \891 ,
  \892 ,
  \893 ,
  \894 ,
  \895 ,
  \896 ,
  \897 ,
  \898 ,
  \899 ,
  \[60] ,
  \900 ,
  \901 ,
  \902 ,
  \903 ,
  \904 ,
  \905 ,
  \908 ,
  \909 ,
  \910 ,
  \913 ,
  \914 ,
  \915 ,
  \918 ,
  \919 ,
  \920 ,
  \923 ,
  \924 ,
  \925 ,
  \928 ,
  \929 ,
  \930 ,
  \933 ,
  \934 ,
  \935 ,
  \938 ,
  \939 ,
  \940 ,
  \943 ,
  \944 ,
  \945 ,
  \948 ,
  \949 ,
  \953 ,
  \954 ;
assign
  \39  = \462 ,
  \40  = \470 ,
  \41  = \478 ,
  \42  = \486 ,
  \43  = \494 ,
  \44  = \502 ,
  \45  = \510 ,
  \46  = \518 ,
  \47  = \526 ,
  \57  = \579  | \1 ,
  \58  = \587  | \1 ,
  \59  = \595  | \1 ,
  \60  = \603  | \1 ,
  \61  = \611  | \1 ,
  \62  = \619  | \1 ,
  \63  = \627  | \1 ,
  \64  = \635  | \1 ,
  \81  = \404  & \22 ,
  \83  = \408  & \407 ,
  \85  = (~\409  & \12 ) | (\409  & ~\12 ),
  \87  = (~\410  & \11 ) | (\410  & ~\11 ),
  \89  = (~\411  & \10 ) | (\411  & ~\10 ),
  \91  = (~\412  & \9 ) | (\412  & ~\9 ),
  \93  = (~\413  & \8 ) | (\413  & ~\8 ),
  \95  = (~\414  & \7 ) | (\414  & ~\7 ),
  \97  = (~\415  & \6 ) | (\415  & ~\6 ),
  \99  = (~\416  & \5 ) | (\416  & ~\5 ),
  \101  = (~\417  & \4 ) | (\417  & ~\4 ),
  \105  = (~\419  & \12 ) | (\419  & ~\12 ),
  \107  = (~\420  & \11 ) | (\420  & ~\11 ),
  \109  = (~\421  & \10 ) | (\421  & ~\10 ),
  \111  = (~\422  & \9 ) | (\422  & ~\9 ),
  \113  = (~\423  & \8 ) | (\423  & ~\8 ),
  \115  = (~\424  & \7 ) | (\424  & ~\7 ),
  \117  = (~\425  & \6 ) | (\425  & ~\6 ),
  \119  = (~\426  & \5 ) | (\426  & ~\5 ),
  \121  = (~\427  & \4 ) | (\427  & ~\4 ),
  \233  = \21  & \38 ,
  \260  = \21  | \38 ,
  \325  = (\455  & \454 ) | ((\455  & \453 ) | (\454  & \453 )),
  \326  = (~\434  & (~\433  & \432 )) | ((~\434  & (\433  & ~\432 )) | ((\434  & (~\433  & ~\432 )) | (\434  & (\433  & \432 )))),
  \327  = (~\437  & (~\436  & \435 )) | ((~\437  & (\436  & ~\435 )) | ((\437  & (~\436  & ~\435 )) | (\437  & (\436  & \435 )))),
  \328  = (~\440  & (~\439  & \438 )) | ((~\440  & (\439  & ~\438 )) | ((\440  & (~\439  & ~\438 )) | (\440  & (\439  & \438 )))),
  \329  = (~\443  & (~\442  & \441 )) | ((~\443  & (\442  & ~\441 )) | ((\443  & (~\442  & ~\441 )) | (\443  & (\442  & \441 )))),
  \330  = (~\446  & (~\445  & \444 )) | ((~\446  & (\445  & ~\444 )) | ((\446  & (~\445  & ~\444 )) | (\446  & (\445  & \444 )))),
  \331  = (~\449  & (~\448  & \447 )) | ((~\449  & (\448  & ~\447 )) | ((\449  & (~\448  & ~\447 )) | (\449  & (\448  & \447 )))),
  \332  = (~\452  & (~\451  & \450 )) | ((~\452  & (\451  & ~\450 )) | ((\452  & (~\451  & ~\450 )) | (\452  & (\451  & \450 )))),
  \333  = (~\455  & (~\454  & \453 )) | ((~\455  & (\454  & ~\453 )) | ((\455  & (~\454  & ~\453 )) | (\455  & (\454  & \453 )))),
  \365  = ~\37  & ~\36 ,
  \368  = \365  & ~\35 ,
  \371  = \368  & ~\34 ,
  \374  = \371  & ~\33 ,
  \377  = \374  & ~\32 ,
  \380  = \377  & ~\31 ,
  \383  = \380  & ~\30 ,
  \386  = \383  & \29 ,
  \389  = \386  & \28 ,
  \392  = \389  & \27 ,
  \395  = \392  & \26 ,
  \398  = \395  & \25 ,
  \401  = \398  & \24 ,
  \404  = \401  & \23 ,
  \407  = (~\21  & ~\38 ) | (\21  & \38 ),
  \408  = \954  & \81 ,
  \409  = \945  & \949 ,
  \410  = \940  & \944 ,
  \411  = \935  & \939 ,
  \412  = \930  & \934 ,
  \413  = \925  & \929 ,
  \414  = \920  & \924 ,
  \415  = \915  & \919 ,
  \416  = \910  & \914 ,
  \417  = \905  & \909 ,
  \418  = \904  & \902 ,
  \419  = \875  & \873 ,
  \420  = \870  & \868 ,
  \421  = \865  & \863 ,
  \422  = \860  & \858 ,
  \423  = \855  & \853 ,
  \424  = \850  & \848 ,
  \425  = \845  & \843 ,
  \426  = \840  & \838 ,
  \427  = \835  & \833 ,
  \428  = \830  & \828 ,
  \430  = \801  & \799 ,
  \431  = \796  & \794 ,
  \432  = \431  & \430 ,
  \433  = \791  & \789 ,
  \434  = \786  & \784 ,
  \435  = (\434  & \433 ) | ((\434  & \432 ) | (\433  & \432 )),
  \436  = \781  & \779 ,
  \437  = \776  & \774 ,
  \438  = (\437  & \436 ) | ((\437  & \435 ) | (\436  & \435 )),
  \439  = \771  & \769 ,
  \440  = \766  & \764 ,
  \441  = (\440  & \439 ) | ((\440  & \438 ) | (\439  & \438 )),
  \442  = \761  & \759 ,
  \443  = \756  & \754 ,
  \444  = (\443  & \442 ) | ((\443  & \441 ) | (\442  & \441 )),
  \445  = \751  & \749 ,
  \446  = \746  & \744 ,
  \447  = (\446  & \445 ) | ((\446  & \444 ) | (\445  & \444 )),
  \448  = \741  & \739 ,
  \449  = \736  & \734 ,
  \450  = (\449  & \448 ) | ((\449  & \447 ) | (\448  & \447 )),
  \451  = \731  & \729 ,
  \452  = \726  & \724 ,
  \453  = (\452  & \451 ) | ((\452  & \450 ) | (\451  & \450 )),
  \454  = \721  & \719 ,
  \455  = \716  & \714 ,
  \456  = \326  & ~\3 ,
  \457  = \4  & \3 ,
  \458  = \457  | \456 ,
  \459  = \458  & \2 ,
  \460  = \13  & ~\2 ,
  \461  = \460  | \459 ,
  \462  = \461  & ~\1 ,
  \464  = \327  & ~\3 ,
  \465  = \5  & \3 ,
  \466  = \465  | \464 ,
  \467  = \466  & \2 ,
  \468  = \14  & ~\2 ,
  \469  = \468  | \467 ,
  \470  = \469  & ~\1 ,
  \472  = \328  & ~\3 ,
  \473  = \6  & \3 ,
  \474  = \473  | \472 ,
  \475  = \474  & \2 ,
  \476  = \15  & ~\2 ,
  \477  = \476  | \475 ,
  \478  = \477  & ~\1 ,
  \480  = \329  & ~\3 ,
  \481  = \7  & \3 ,
  \482  = \481  | \480 ,
  \483  = \482  & \2 ,
  \484  = \16  & ~\2 ,
  \485  = \484  | \483 ,
  \486  = \485  & ~\1 ,
  \488  = \330  & ~\3 ,
  \489  = \8  & \3 ,
  \490  = \489  | \488 ,
  \491  = \490  & \2 ,
  \492  = \17  & ~\2 ,
  \493  = \492  | \491 ,
  \494  = \493  & ~\1 ,
  \496  = \331  & ~\3 ,
  \497  = \9  & \3 ,
  \498  = \497  | \496 ,
  \499  = \498  & \2 ,
  \500  = \18  & ~\2 ,
  \501  = \500  | \499 ,
  \502  = \501  & ~\1 ,
  \504  = \332  & ~\3 ,
  \505  = \10  & \3 ,
  \506  = \505  | \504 ,
  \507  = \506  & \2 ,
  \508  = \19  & ~\2 ,
  \509  = \508  | \507 ,
  \510  = \509  & ~\1 ,
  \512  = \333  & ~\3 ,
  \513  = \11  & \3 ,
  \514  = \513  | \512 ,
  \515  = \514  & \2 ,
  \516  = \20  & ~\2 ,
  \517  = \516  | \515 ,
  \518  = \517  & ~\1 ,
  \520  = \325  & ~\3 ,
  \521  = \12  & \3 ,
  \522  = \521  | \520 ,
  \523  = \522  & \2 ,
  \524  = \21  & ~\2 ,
  \525  = \524  | \523 ,
  \526  = \525  & ~\1 ,
  \528  = \4  & \2 ,
  \529  = \13  & ~\2 ,
  \530  = \529  | \528 ,
  \531  = \530  & ~\1 ,
  \533  = \5  & \2 ,
  \534  = \14  & ~\2 ,
  \535  = \534  | \533 ,
  \536  = \535  & ~\1 ,
  \538  = \6  & \2 ,
  \539  = \15  & ~\2 ,
  \540  = \539  | \538 ,
  \541  = \540  & ~\1 ,
  \543  = \7  & \2 ,
  \544  = \16  & ~\2 ,
  \545  = \544  | \543 ,
  \546  = \545  & ~\1 ,
  \548  = \8  & \2 ,
  \549  = \17  & ~\2 ,
  \550  = \549  | \548 ,
  \551  = \550  & ~\1 ,
  \553  = \9  & \2 ,
  \554  = \18  & ~\2 ,
  \555  = \554  | \553 ,
  \556  = \555  & ~\1 ,
  \558  = \10  & \2 ,
  \559  = \19  & ~\2 ,
  \560  = \559  | \558 ,
  \561  = \560  & ~\1 ,
  \563  = \11  & \2 ,
  \564  = \20  & ~\2 ,
  \565  = \564  | \563 ,
  \566  = \565  & ~\1 ,
  \568  = \12  & \2 ,
  \569  = \21  & ~\2 ,
  \570  = \569  | \568 ,
  \571  = \570  & ~\1 ,
  \573  = \431  & ~\3 ,
  \575  = \573  | \3 ,
  \576  = \575  & \2 ,
  \578  = \576  | ~\2 ,
  \579  = \578  & ~\1 ,
  \581  = \434  & ~\3 ,
  \583  = \581  | \3 ,
  \584  = \583  & \2 ,
  \586  = \584  | ~\2 ,
  \587  = \586  & ~\1 ,
  \589  = \437  & ~\3 ,
  \591  = \589  | \3 ,
  \592  = \591  & \2 ,
  \594  = \592  | ~\2 ,
  \595  = \594  & ~\1 ,
  \597  = \440  & ~\3 ,
  \599  = \597  | \3 ,
  \[35]  = \531 ,
  \[36]  = \536 ,
  \600  = \599  & \2 ,
  \602  = \600  | ~\2 ,
  \603  = \602  & ~\1 ,
  \605  = \443  & ~\3 ,
  \607  = \605  | \3 ,
  \608  = \607  & \2 ,
  \[37]  = \541 ,
  \610  = \608  | ~\2 ,
  \611  = \610  & ~\1 ,
  \613  = \446  & ~\3 ,
  \615  = \613  | \3 ,
  \616  = \615  & \2 ,
  \618  = \616  | ~\2 ,
  \619  = \618  & ~\1 ,
  \[38]  = \546 ,
  \621  = \449  & ~\3 ,
  \623  = \621  | \3 ,
  \624  = \623  & \2 ,
  \626  = \624  | ~\2 ,
  \627  = \626  & ~\1 ,
  \629  = \452  & ~\3 ,
  \[39]  = \551 ,
  \631  = \629  | \3 ,
  \632  = \631  & \2 ,
  \634  = \632  | ~\2 ,
  \635  = \634  & ~\1 ,
  \637  = \430  & ~\3 ,
  \640  = \637  & \2 ,
  \643  = \640  & ~\1 ,
  \645  = \433  & ~\3 ,
  \648  = \645  & \2 ,
  \651  = \648  & ~\1 ,
  \653  = \436  & ~\3 ,
  \656  = \653  & \2 ,
  \659  = \656  & ~\1 ,
  \661  = \439  & ~\3 ,
  \664  = \661  & \2 ,
  \667  = \664  & ~\1 ,
  \669  = \442  & ~\3 ,
  \672  = \669  & \2 ,
  \675  = \672  & ~\1 ,
  \677  = \445  & ~\3 ,
  \680  = \677  & \2 ,
  \683  = \680  & ~\1 ,
  \685  = \448  & ~\3 ,
  \688  = \685  & \2 ,
  \691  = \688  & ~\1 ,
  \693  = \451  & ~\3 ,
  \696  = \693  & \2 ,
  \699  = \696  & ~\1 ,
  \[40]  = \556 ,
  \[41]  = \561 ,
  \[42]  = \566 ,
  \[43]  = \571 ,
  \[44]  = \57 ,
  \[45]  = \58 ,
  \[46]  = \59 ,
  \701  = \455  & \12 ,
  \702  = \454  & ~\12 ,
  \703  = \702  | \701 ,
  \704  = \703  & ~\3 ,
  \705  = \12  & \3 ,
  \706  = \705  | \704 ,
  \707  = \706  & \2 ,
  \708  = \21  & ~\2 ,
  \709  = \708  | \707 ,
  \[47]  = \60 ,
  \710  = \709  & ~\1 ,
  \712  = ~\428  & \12 ,
  \713  = \428  & \419 ,
  \714  = \713  | \712 ,
  \715  = ~\3  & \2 ,
  \716  = \715  & ~\1 ,
  \717  = ~\418  & \409 ,
  \718  = \418  & \12 ,
  \719  = \718  | \717 ,
  \[48]  = \61 ,
  \720  = ~\3  & \2 ,
  \721  = \720  & ~\1 ,
  \722  = ~\428  & \11 ,
  \723  = \428  & \420 ,
  \724  = \723  | \722 ,
  \725  = ~\3  & \2 ,
  \726  = \725  & ~\1 ,
  \727  = ~\418  & \410 ,
  \728  = \418  & \11 ,
  \729  = \728  | \727 ,
  \[49]  = \62 ,
  \730  = ~\3  & \2 ,
  \731  = \730  & ~\1 ,
  \732  = ~\428  & \10 ,
  \733  = \428  & \421 ,
  \734  = \733  | \732 ,
  \735  = ~\3  & \2 ,
  \736  = \735  & ~\1 ,
  \737  = ~\418  & \411 ,
  \738  = \418  & \10 ,
  \739  = \738  | \737 ,
  \740  = ~\3  & \2 ,
  \741  = \740  & ~\1 ,
  \742  = ~\428  & \9 ,
  \743  = \428  & \422 ,
  \744  = \743  | \742 ,
  \745  = ~\3  & \2 ,
  \746  = \745  & ~\1 ,
  \747  = ~\418  & \412 ,
  \748  = \418  & \9 ,
  \749  = \748  | \747 ,
  \750  = ~\3  & \2 ,
  \751  = \750  & ~\1 ,
  \752  = ~\428  & \8 ,
  \753  = \428  & \423 ,
  \754  = \753  | \752 ,
  \755  = ~\3  & \2 ,
  \756  = \755  & ~\1 ,
  \757  = ~\418  & \413 ,
  \758  = \418  & \8 ,
  \759  = \758  | \757 ,
  \760  = ~\3  & \2 ,
  \761  = \760  & ~\1 ,
  \762  = ~\428  & \7 ,
  \763  = \428  & \424 ,
  \764  = \763  | \762 ,
  \765  = ~\3  & \2 ,
  \766  = \765  & ~\1 ,
  \767  = ~\418  & \414 ,
  \768  = \418  & \7 ,
  \769  = \768  | \767 ,
  \770  = ~\3  & \2 ,
  \771  = \770  & ~\1 ,
  \772  = ~\428  & \6 ,
  \773  = \428  & \425 ,
  \774  = \773  | \772 ,
  \775  = ~\3  & \2 ,
  \776  = \775  & ~\1 ,
  \777  = ~\418  & \415 ,
  \778  = \418  & \6 ,
  \779  = \778  | \777 ,
  \780  = ~\3  & \2 ,
  \781  = \780  & ~\1 ,
  \782  = ~\428  & \5 ,
  \783  = \428  & \426 ,
  \784  = \783  | \782 ,
  \785  = ~\3  & \2 ,
  \786  = \785  & ~\1 ,
  \787  = ~\418  & \416 ,
  \788  = \418  & \5 ,
  \789  = \788  | \787 ,
  \790  = ~\3  & \2 ,
  \791  = \790  & ~\1 ,
  \792  = ~\428  & \4 ,
  \793  = \428  & \427 ,
  \794  = \793  | \792 ,
  \795  = ~\3  & \2 ,
  \796  = \795  & ~\1 ,
  \797  = ~\418  & \417 ,
  \798  = \418  & \4 ,
  \799  = \798  | \797 ,
  \[50]  = \63 ,
  \[51]  = \64 ,
  \[52]  = \643 ,
  \[53]  = \651 ,
  \[54]  = \659 ,
  \[55]  = \667 ,
  \[56]  = \675 ,
  \800  = ~\3  & \2 ,
  \801  = \800  & ~\1 ,
  \803  = \121  & \4 ,
  \805  = \803  & ~\119 ,
  \806  = \119  & \5 ,
  \807  = \806  | \805 ,
  \808  = \807  & ~\117 ,
  \809  = \117  & \6 ,
  \[57]  = \683 ,
  \810  = \809  | \808 ,
  \811  = \810  & ~\115 ,
  \812  = \115  & \7 ,
  \813  = \812  | \811 ,
  \814  = \813  & ~\113 ,
  \815  = \113  & \8 ,
  \816  = \815  | \814 ,
  \817  = \816  & ~\111 ,
  \818  = \111  & \9 ,
  \819  = \818  | \817 ,
  \[58]  = \691 ,
  \820  = \819  & ~\109 ,
  \821  = \109  & \10 ,
  \822  = \821  | \820 ,
  \823  = \822  & ~\107 ,
  \824  = \107  & \11 ,
  \825  = \824  | \823 ,
  \826  = \825  & ~\105 ,
  \827  = \105  & \12 ,
  \828  = \827  | \826 ,
  \829  = ~\3  & \2 ,
  \[59]  = \699 ,
  \830  = \829  & ~\1 ,
  \831  = ~\83  & \22 ,
  \833  = \831  | \83 ,
  \834  = ~\3  & \2 ,
  \835  = \834  & ~\1 ,
  \836  = ~\83  & \23 ,
  \838  = \836  | \83 ,
  \839  = ~\3  & \2 ,
  \840  = \839  & ~\1 ,
  \841  = ~\83  & \24 ,
  \843  = \841  | \83 ,
  \844  = ~\3  & \2 ,
  \845  = \844  & ~\1 ,
  \846  = ~\83  & \25 ,
  \848  = \846  | \83 ,
  \849  = ~\3  & \2 ,
  \850  = \849  & ~\1 ,
  \851  = ~\83  & \26 ,
  \853  = \851  | \83 ,
  \854  = ~\3  & \2 ,
  \855  = \854  & ~\1 ,
  \856  = ~\83  & \27 ,
  \858  = \856  | \83 ,
  \859  = ~\3  & \2 ,
  \860  = \859  & ~\1 ,
  \861  = ~\83  & \28 ,
  \863  = \861  | \83 ,
  \864  = ~\3  & \2 ,
  \865  = \864  & ~\1 ,
  \866  = ~\83  & \29 ,
  \868  = \866  | \83 ,
  \869  = ~\3  & \2 ,
  \870  = \869  & ~\1 ,
  \871  = \233  & ~\83 ,
  \873  = \871  | \83 ,
  \874  = ~\3  & \2 ,
  \875  = \874  & ~\1 ,
  \877  = \101  & \4 ,
  \879  = \877  & ~\99 ,
  \880  = \99  & \5 ,
  \881  = \880  | \879 ,
  \882  = \881  & ~\97 ,
  \883  = \97  & \6 ,
  \884  = \883  | \882 ,
  \885  = \884  & ~\95 ,
  \886  = \95  & \7 ,
  \887  = \886  | \885 ,
  \888  = \887  & ~\93 ,
  \889  = \93  & \8 ,
  \890  = \889  | \888 ,
  \891  = \890  & ~\91 ,
  \892  = \91  & \9 ,
  \893  = \892  | \891 ,
  \894  = \893  & ~\89 ,
  \895  = \89  & \10 ,
  \896  = \895  | \894 ,
  \897  = \896  & ~\87 ,
  \898  = \87  & \11 ,
  \899  = \898  | \897 ,
  \[60]  = \710 ,
  \900  = \899  & ~\85 ,
  \901  = \85  & \12 ,
  \902  = \901  | \900 ,
  \903  = ~\3  & \2 ,
  \904  = \903  & ~\1 ,
  \905  = ~\83  & \30 ,
  \908  = ~\3  & \2 ,
  \909  = \908  & ~\1 ,
  \910  = ~\83  & \31 ,
  \913  = ~\3  & \2 ,
  \914  = \913  & ~\1 ,
  \915  = ~\83  & \32 ,
  \918  = ~\3  & \2 ,
  \919  = \918  & ~\1 ,
  \920  = ~\83  & \33 ,
  \923  = ~\3  & \2 ,
  \924  = \923  & ~\1 ,
  \925  = ~\83  & \34 ,
  \928  = ~\3  & \2 ,
  \929  = \928  & ~\1 ,
  \930  = ~\83  & \35 ,
  \933  = ~\3  & \2 ,
  \934  = \933  & ~\1 ,
  \935  = ~\83  & \36 ,
  \938  = ~\3  & \2 ,
  \939  = \938  & ~\1 ,
  \940  = ~\83  & \37 ,
  \943  = ~\3  & \2 ,
  \944  = \943  & ~\1 ,
  \945  = \260  & ~\83 ,
  \948  = ~\3  & \2 ,
  \949  = \948  & ~\1 ,
  \953  = ~\3  & \2 ,
  \954  = \953  & ~\1 ;
always begin
  \13  = \[35] ;
  \14  = \[36] ;
  \15  = \[37] ;
  \16  = \[38] ;
  \17  = \[39] ;
  \18  = \[40] ;
  \19  = \[41] ;
  \20  = \[42] ;
  \21  = \[43] ;
  \22  = \[44] ;
  \23  = \[45] ;
  \24  = \[46] ;
  \25  = \[47] ;
  \26  = \[48] ;
  \27  = \[49] ;
  \28  = \[50] ;
  \29  = \[51] ;
  \30  = \[52] ;
  \31  = \[53] ;
  \32  = \[54] ;
  \33  = \[55] ;
  \34  = \[56] ;
  \35  = \[57] ;
  \36  = \[58] ;
  \37  = \[59] ;
  \38  = \[60] ;
end
initial begin
  \13  = 0;
  \14  = 0;
  \15  = 0;
  \16  = 0;
  \17  = 0;
  \18  = 0;
  \19  = 0;
  \20  = 0;
  \21  = 0;
  \22  = 1;
  \23  = 1;
  \24  = 1;
  \25  = 1;
  \26  = 1;
  \27  = 1;
  \28  = 1;
  \29  = 1;
  \30  = 0;
  \31  = 0;
  \32  = 0;
  \33  = 0;
  \34  = 0;
  \35  = 0;
  \36  = 0;
  \37  = 0;
  \38  = 0;
end
endmodule

