//NOTE: no-implementation module stub

module PSQ (
    input T_RST,
    input DSPCLK,
    input X_PWDn,
    input X_IRQ2n,
    input X_IRQL1n,
    input X_IRQL0n,
    input X_IRQE1n,
    input X_IRQE0n,
    input X_IRQ1n,
    input X_IRQ0n,
    input T_IST0,
    input T_ISR0,
    input T_IST1,
    input T_ISR1,
    input T_ITMR,
    input [17:4] IR,
    input [15:0] DMDix,
    input RSTtext_h,
    input Awake,
    input enTRAP_RL,
    input STBY,
    input [19:0] IRE,
    input EX_en,
    input Dummy_R,
    input dBR_R,
    input idBR_R,
    input RET_R,
    input DU_Eg,
    input Call_Ed,
    input RTI_Ed,
    input BR_Ed,
    input EXIT_E,
    input RET_Ed,
    input Nseq_Ed,
    input IDLE_Eg,
    input MACdep_Eg,
    input LDaST_Eg,
    input MTCNTR_Eg,
    input MTOWRCNTR_Eg,
    input MTtoppcs_Eg,
    input MTIMASK_Eg,
    input MTICNTL_Eg,
    input MTIFC_Eg,
    input MTMSTAT_Eg,
    input MFPSQ_E,
    input MFtoppcs_E,
    input MFIMASK_E,
    input MFICNTL_E,
    input MFSSTAT_E,
    input MFMSTAT_E,
    input MFCNTR_E,
    input Stkctl_Eg,
    input Modctl_Eg,
    input MpopLP_Eg,
    input imm16_E,
    input imm14_E,
    input MFIDR_E,
    input Long_Eg,
    input Nrti_Ed,
    input MTPMOVL_E,
    input MTDMOVL_E,
    input MFPMOVL_E,
    input MFDMOVL_E,
    input accCM_R,
    input accCM_E,
    input [13:0] Bt_I,
    input BTaken_I,
    input RTaken_I,
    input PTaken_R,
    input PTaken_E,
    input [13:0] PMA_R,
    input Ctrue,
    input Ttrue,
    input [7:0] ASTAT,
    input SP1_EN,
    input X_BRn,
    input eRDY,
    input EXTC_Eg,
    input STI_Cg,
    input BOOT,
    input STEAL,
    input SREQ,
    input [13:0] DCTL,
    input DSreqx,
    input GO_Fx,
    input GO_Ex,
    input GO_Cx,
    input [13:0] IRR,
    input [15:0] IDR,
    input HALT_Eg,
    input GOICE_syn,
    input PDFORCE,
    input [13:0] BIAD,
    input T_BDMA,
    input BSreqx,
    `ifdef FD_DFT
    input SCAN_TEST,
    `endif
    input GO_F,
    input GO_D,
    input GO_E,
    input GO_C,
    input PPclr_h,
    input [6:0] MSTAT,
    input ICE_ST_h,
    input ICE_ST,
    input IDLE_ST_h,
    input IDLE_ST,
    input TRAP_Eg,
    input redoM_h,
    input redoSTI_h,
    input redoLD_h,
    input redoEX_h,
    input TRAP_R,
    input TRAP_R_L,
    input Prderr_Eg,
    input Bterr_E,
    input [13:0] Taddr_E,
    input [4:0] IFA_nx,
    input CE,
    input VpopST_Eg,
    input [7:0] popASTATo,
    input [3:0] Term,
    input GO_MAC,
    input BGn,
    input [13:0] IFA,
    input [7:0] PMOVL,
    input [3:0] DMOVL,
    input redoIF_h,
    input GO_EC,
    input ECYC,
    input [13:0] CMAin,
    input HALTclr_h,
    input GOICEclr_h,
    input GOICEdis,
    input [13:0] DRA,
    input [13:0] EXA,
    output [15:0] psqDMD_do
);

endmodule
