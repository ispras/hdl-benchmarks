// IWLS benchmark module "cordic" printed on Wed May 29 16:31:29 2002
module cordic(a6, a4, a3, a2, a5, v, x0, x1, x2, x3, y0, y1, y2, y3, z0, z1, z2, ex0, ex1, ex2, ey0, ey1, ey2, d, dn);
input
  z0,
  z1,
  z2,
  v,
  ex0,
  ex1,
  ex2,
  ey0,
  ey1,
  ey2,
  a2,
  a3,
  a4,
  a5,
  a6,
  x0,
  x1,
  x2,
  x3,
  y0,
  y1,
  y2,
  y3;
output
  dn,
  d;
wire
  \[368] ,
  \[375] ,
  \[8] ,
  \[157] ,
  \[376] ,
  \[0] ,
  \[505] ,
  \[1] ,
  \[511] ,
  \[367] ,
  \[6] ;
assign
  \[368]  = (~x3 & x2) | (x3 & ~x2),
  \[375]  = (~y1 & ~y0) | (y1 & y0),
  \[8]  = (~z2 & (~z1 & z0)) | ((z2 & (z1 & ~z0)) | ((~\[376]  & ~\[375] ) | ((\[376]  & \[375] ) | ((~\[368]  & ~\[367] ) | (\[368]  & \[367] ))))),
  \[157]  = (~ey2 & (~ey1 & (~ey0 & (~ex2 & (~ex1 & ~ex0))))) | ((~ey2 & (~ey1 & (~ey0 & (ex2 & (ex1 & ex0))))) | ((ey2 & (ey1 & (ey0 & (~ex2 & (~ex1 & ~ex0))))) | (ey2 & (ey1 & (ey0 & (ex2 & (ex1 & ex0))))))),
  \[376]  = (~y3 & y2) | (y3 & ~y2),
  dn = \[1] ,
  \[0]  = (\[6]  & (~\[157]  & \[505] )) | ~\[1] ,
  \[505]  = a2 | (a3 | (~a4 | ~a6)),
  d = \[0] ,
  \[1]  = (~\[8]  & (\[157]  & ~v)) | ((\[6]  & ~v) | ~\[511] ),
  \[511]  = a5 | (a2 | (a3 | (a4 | a6))),
  \[367]  = (~x1 & ~x0) | (x1 & x0),
  \[6]  = (~a2 & (a3 & (~a4 & a6))) | ~\[505] ;
endmodule

