//NOTE: no-implementation module stub

module GTECH_MUX8 (
    input wire [2:0] S,
    input wire A,
    input wire B,
    input wire C,
    input wire D0,
    input wire D1,
    input wire D2,
    input wire D3,
    input wire D4,
    input wire D5,
    input wire D6,
    input wire D7,
    output wire Z
);

endmodule
