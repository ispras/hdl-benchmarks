

































































`define DMA_MAX_CHNO 8 
`define DMA_HAVE_CH0 
`define DMA_HAVE_CH1 
`define DMA_HAVE_CH2 
`define DMA_HAVE_CH3 
`define DMA_HAVE_CH4 
`define DMA_HAVE_CH5 
`define DMA_HAVE_CH6 
`define DMA_HAVE_CH7 


`define DMA_HAVE_BRIDGE 


`define DMA_HAVE_AHB1 


`define DMA_HAVE_LINKLIST 



`define DMA_FF_TH 8 
`define DMA_FF_ADD_WIDTH 3 
`include "DMA_FIX_DEFINE.vh" 
